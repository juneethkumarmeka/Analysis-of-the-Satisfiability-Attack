module basic_3000_30000_3500_150_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_653,In_1408);
and U1 (N_1,In_2503,In_2876);
nor U2 (N_2,In_1361,In_2401);
nand U3 (N_3,In_1466,In_1106);
nor U4 (N_4,In_709,In_1428);
xnor U5 (N_5,In_1798,In_2245);
or U6 (N_6,In_2691,In_1663);
and U7 (N_7,In_2649,In_2175);
nand U8 (N_8,In_1620,In_2229);
nand U9 (N_9,In_1727,In_307);
nand U10 (N_10,In_1149,In_1314);
nand U11 (N_11,In_324,In_2594);
nor U12 (N_12,In_447,In_88);
and U13 (N_13,In_2798,In_1771);
nand U14 (N_14,In_2886,In_822);
xor U15 (N_15,In_710,In_334);
and U16 (N_16,In_2903,In_1407);
nor U17 (N_17,In_588,In_2641);
nor U18 (N_18,In_490,In_605);
and U19 (N_19,In_789,In_715);
nand U20 (N_20,In_1604,In_2607);
nand U21 (N_21,In_1935,In_997);
nand U22 (N_22,In_2666,In_2900);
nand U23 (N_23,In_2013,In_949);
xor U24 (N_24,In_1923,In_1014);
and U25 (N_25,In_589,In_555);
xor U26 (N_26,In_2249,In_990);
xor U27 (N_27,In_1778,In_1949);
and U28 (N_28,In_2687,In_941);
or U29 (N_29,In_2655,In_2343);
nor U30 (N_30,In_1285,In_2370);
nor U31 (N_31,In_1215,In_2162);
or U32 (N_32,In_1198,In_1832);
xor U33 (N_33,In_873,In_1510);
nor U34 (N_34,In_2638,In_115);
nor U35 (N_35,In_2684,In_1824);
xor U36 (N_36,In_2730,In_1556);
and U37 (N_37,In_1977,In_207);
or U38 (N_38,In_2048,In_425);
and U39 (N_39,In_2880,In_1305);
nor U40 (N_40,In_638,In_1288);
or U41 (N_41,In_2458,In_482);
or U42 (N_42,In_360,In_2637);
xnor U43 (N_43,In_198,In_2344);
nor U44 (N_44,In_2979,In_1060);
or U45 (N_45,In_1272,In_811);
xor U46 (N_46,In_2051,In_1256);
and U47 (N_47,In_2211,In_861);
or U48 (N_48,In_1787,In_1085);
xnor U49 (N_49,In_1374,In_2827);
nor U50 (N_50,In_714,In_2188);
or U51 (N_51,In_1377,In_84);
or U52 (N_52,In_2824,In_2657);
and U53 (N_53,In_2285,In_1416);
or U54 (N_54,In_1677,In_1793);
or U55 (N_55,In_1699,In_366);
and U56 (N_56,In_1839,In_572);
xor U57 (N_57,In_126,In_2072);
or U58 (N_58,In_2368,In_2003);
nand U59 (N_59,In_1298,In_1701);
or U60 (N_60,In_2681,In_2036);
nand U61 (N_61,In_1204,In_1094);
nor U62 (N_62,In_1858,In_2017);
nor U63 (N_63,In_2189,In_2236);
nand U64 (N_64,In_568,In_2970);
and U65 (N_65,In_991,In_687);
xor U66 (N_66,In_7,In_1647);
or U67 (N_67,In_2582,In_202);
nor U68 (N_68,In_1841,In_2144);
and U69 (N_69,In_1936,In_1296);
xor U70 (N_70,In_2323,In_2595);
or U71 (N_71,In_278,In_1584);
or U72 (N_72,In_1736,In_2842);
xor U73 (N_73,In_2535,In_368);
xor U74 (N_74,In_1483,In_61);
nor U75 (N_75,In_1718,In_1872);
nor U76 (N_76,In_1074,In_2800);
nor U77 (N_77,In_1000,In_59);
nor U78 (N_78,In_2152,In_648);
and U79 (N_79,In_182,In_1375);
or U80 (N_80,In_1698,In_1570);
nand U81 (N_81,In_64,In_580);
nor U82 (N_82,In_1174,In_2084);
and U83 (N_83,In_2895,In_2784);
xor U84 (N_84,In_2635,In_1214);
nand U85 (N_85,In_1444,In_890);
nor U86 (N_86,In_684,In_987);
nand U87 (N_87,In_2546,In_1630);
and U88 (N_88,In_2751,In_1997);
or U89 (N_89,In_1911,In_1527);
and U90 (N_90,In_650,In_2106);
xnor U91 (N_91,In_2685,In_2530);
nor U92 (N_92,In_1291,In_1598);
nand U93 (N_93,In_1823,In_1354);
nor U94 (N_94,In_2678,In_1413);
nand U95 (N_95,In_2563,In_1742);
and U96 (N_96,In_1397,In_578);
or U97 (N_97,In_475,In_1726);
nand U98 (N_98,In_336,In_36);
xor U99 (N_99,In_1998,In_1730);
nor U100 (N_100,In_807,In_901);
nand U101 (N_101,In_2142,In_1062);
xor U102 (N_102,In_2041,In_2485);
nand U103 (N_103,In_924,In_1825);
nand U104 (N_104,In_2606,In_2772);
and U105 (N_105,In_184,In_2555);
nand U106 (N_106,In_358,In_850);
nand U107 (N_107,In_2472,In_1147);
nor U108 (N_108,In_2569,In_2646);
and U109 (N_109,In_905,In_1897);
xnor U110 (N_110,In_737,In_1007);
xnor U111 (N_111,In_1142,In_2576);
nand U112 (N_112,In_1696,In_522);
or U113 (N_113,In_1469,In_1477);
xnor U114 (N_114,In_2651,In_1208);
or U115 (N_115,In_1864,In_611);
nand U116 (N_116,In_621,In_1667);
and U117 (N_117,In_1226,In_466);
or U118 (N_118,In_593,In_49);
xnor U119 (N_119,In_1980,In_2961);
xor U120 (N_120,In_2934,In_893);
or U121 (N_121,In_9,In_1020);
nand U122 (N_122,In_478,In_1616);
nor U123 (N_123,In_2132,In_1826);
or U124 (N_124,In_2000,In_998);
or U125 (N_125,In_66,In_2686);
or U126 (N_126,In_1355,In_1964);
xnor U127 (N_127,In_1645,In_2930);
or U128 (N_128,In_34,In_2513);
and U129 (N_129,In_678,In_586);
or U130 (N_130,In_2831,In_22);
xor U131 (N_131,In_62,In_2781);
nor U132 (N_132,In_1888,In_20);
xor U133 (N_133,In_1286,In_888);
nor U134 (N_134,In_1763,In_2562);
xnor U135 (N_135,In_1751,In_2139);
xnor U136 (N_136,In_614,In_1329);
or U137 (N_137,In_628,In_966);
xnor U138 (N_138,In_544,In_2253);
and U139 (N_139,In_1788,In_2810);
xnor U140 (N_140,In_1536,In_1830);
nand U141 (N_141,In_17,In_2622);
xor U142 (N_142,In_2160,In_428);
nand U143 (N_143,In_866,In_2969);
nand U144 (N_144,In_1780,In_1302);
and U145 (N_145,In_1590,In_1404);
xor U146 (N_146,In_2461,In_2644);
or U147 (N_147,In_19,In_1603);
and U148 (N_148,In_756,In_1947);
or U149 (N_149,In_1595,In_102);
nor U150 (N_150,In_2719,In_782);
nor U151 (N_151,In_733,In_86);
and U152 (N_152,In_1072,In_1225);
and U153 (N_153,In_192,In_1546);
xor U154 (N_154,In_2235,In_2814);
xnor U155 (N_155,In_2990,In_1126);
xnor U156 (N_156,In_1899,In_1114);
and U157 (N_157,In_2349,In_2418);
xor U158 (N_158,In_537,In_189);
or U159 (N_159,In_379,In_2373);
and U160 (N_160,In_2664,In_1379);
nor U161 (N_161,In_1955,In_796);
nor U162 (N_162,In_985,In_1187);
or U163 (N_163,In_1414,In_2426);
nor U164 (N_164,In_2325,In_690);
xor U165 (N_165,In_2540,In_2987);
xor U166 (N_166,In_2296,In_331);
xnor U167 (N_167,In_1593,In_500);
or U168 (N_168,In_1451,In_1756);
and U169 (N_169,In_2611,In_1229);
and U170 (N_170,In_2700,In_1674);
xnor U171 (N_171,In_1574,In_30);
nor U172 (N_172,In_57,In_1680);
and U173 (N_173,In_864,In_2670);
and U174 (N_174,In_180,In_1326);
nand U175 (N_175,In_453,In_1464);
and U176 (N_176,In_2591,In_1580);
nand U177 (N_177,In_2140,In_105);
or U178 (N_178,In_892,In_932);
nor U179 (N_179,In_1626,In_2650);
xor U180 (N_180,In_881,In_210);
xor U181 (N_181,In_1242,In_2436);
nand U182 (N_182,In_1112,In_625);
xor U183 (N_183,In_2532,In_2740);
or U184 (N_184,In_2858,In_2980);
and U185 (N_185,In_567,In_1009);
xnor U186 (N_186,In_146,In_2374);
xnor U187 (N_187,In_814,In_217);
and U188 (N_188,In_1493,In_1656);
nand U189 (N_189,In_2494,In_96);
or U190 (N_190,In_1925,In_2257);
and U191 (N_191,In_2796,In_1282);
xor U192 (N_192,In_1765,In_2094);
nand U193 (N_193,In_1902,In_2205);
and U194 (N_194,In_1708,In_1212);
xnor U195 (N_195,In_536,In_325);
or U196 (N_196,In_2214,In_2981);
and U197 (N_197,In_792,In_1153);
and U198 (N_198,In_1439,In_2272);
nand U199 (N_199,In_2108,In_2081);
nor U200 (N_200,In_2887,In_1158);
nand U201 (N_201,In_1188,In_2720);
and U202 (N_202,In_2748,In_1492);
xnor U203 (N_203,In_196,In_664);
and U204 (N_204,In_1786,In_2742);
nand U205 (N_205,In_349,In_2250);
and U206 (N_206,In_1065,In_1873);
and U207 (N_207,In_1422,In_1213);
or U208 (N_208,In_1795,In_1359);
and U209 (N_209,N_30,N_190);
and U210 (N_210,In_2931,In_332);
or U211 (N_211,N_198,In_157);
nand U212 (N_212,In_1983,In_1392);
xnor U213 (N_213,In_1032,N_82);
nand U214 (N_214,In_1643,In_2419);
xor U215 (N_215,In_2406,In_2303);
and U216 (N_216,In_1043,In_896);
xnor U217 (N_217,In_2092,In_199);
nor U218 (N_218,In_2093,In_1034);
or U219 (N_219,In_2201,In_175);
nand U220 (N_220,In_251,In_78);
xor U221 (N_221,In_242,In_290);
and U222 (N_222,In_2804,In_2445);
and U223 (N_223,In_2805,In_298);
nor U224 (N_224,In_11,In_1356);
nor U225 (N_225,In_506,N_111);
xor U226 (N_226,In_1211,In_1253);
xor U227 (N_227,In_1050,In_1070);
xnor U228 (N_228,In_44,In_601);
and U229 (N_229,N_2,In_793);
nor U230 (N_230,In_582,In_933);
and U231 (N_231,In_2277,In_1912);
nor U232 (N_232,In_765,In_361);
xnor U233 (N_233,In_1898,N_35);
nor U234 (N_234,In_1679,In_2791);
nand U235 (N_235,In_1908,In_398);
nand U236 (N_236,In_350,In_415);
or U237 (N_237,In_778,In_2806);
or U238 (N_238,In_620,In_419);
nor U239 (N_239,In_2807,In_2902);
nor U240 (N_240,In_618,In_156);
nor U241 (N_241,In_381,In_2975);
xor U242 (N_242,In_1185,In_1886);
and U243 (N_243,In_2669,In_2982);
xnor U244 (N_244,In_2451,In_590);
nand U245 (N_245,In_333,In_2258);
nand U246 (N_246,In_676,In_1423);
and U247 (N_247,In_812,In_56);
or U248 (N_248,In_449,In_173);
nor U249 (N_249,In_1715,In_2398);
or U250 (N_250,In_1722,In_2482);
nand U251 (N_251,In_285,In_1884);
nor U252 (N_252,In_2034,In_2575);
xnor U253 (N_253,In_227,In_1999);
xor U254 (N_254,In_2116,In_2709);
and U255 (N_255,In_777,In_695);
nand U256 (N_256,In_732,In_1497);
xnor U257 (N_257,In_2598,In_1137);
nand U258 (N_258,N_123,In_1491);
nand U259 (N_259,In_2099,In_1564);
xnor U260 (N_260,N_154,In_2518);
or U261 (N_261,In_2935,N_127);
nand U262 (N_262,In_2290,In_2002);
nand U263 (N_263,In_230,In_2376);
nand U264 (N_264,In_1460,In_2115);
nor U265 (N_265,In_1967,In_1022);
and U266 (N_266,In_1867,In_2531);
xor U267 (N_267,In_2843,In_370);
or U268 (N_268,In_2021,In_2399);
and U269 (N_269,In_768,In_255);
and U270 (N_270,In_417,In_2878);
xor U271 (N_271,In_2945,In_1498);
nor U272 (N_272,In_2788,In_2988);
or U273 (N_273,In_2404,N_192);
nand U274 (N_274,In_2022,In_233);
or U275 (N_275,N_26,In_471);
or U276 (N_276,In_1853,In_1535);
and U277 (N_277,In_2917,In_713);
or U278 (N_278,In_1711,In_1686);
or U279 (N_279,In_2244,In_511);
nand U280 (N_280,In_984,N_163);
nand U281 (N_281,In_293,In_1928);
xor U282 (N_282,N_18,In_579);
or U283 (N_283,In_619,In_2424);
and U284 (N_284,In_2318,In_2570);
and U285 (N_285,In_749,In_137);
nor U286 (N_286,In_762,In_2083);
nand U287 (N_287,In_2006,In_2243);
nand U288 (N_288,In_2141,In_2762);
and U289 (N_289,In_1266,In_372);
nor U290 (N_290,In_2568,In_718);
or U291 (N_291,In_657,In_2809);
nor U292 (N_292,N_38,In_2486);
nand U293 (N_293,In_1611,In_1077);
xnor U294 (N_294,In_2763,In_1505);
xnor U295 (N_295,In_90,In_218);
nor U296 (N_296,In_1357,In_688);
and U297 (N_297,In_805,In_1878);
xor U298 (N_298,In_1910,In_426);
nand U299 (N_299,In_441,In_2792);
nor U300 (N_300,In_716,In_1136);
or U301 (N_301,In_480,In_2996);
or U302 (N_302,In_2653,In_2114);
nand U303 (N_303,In_1642,In_267);
xor U304 (N_304,In_772,In_1594);
nor U305 (N_305,In_1271,In_1487);
xor U306 (N_306,In_47,In_1154);
nor U307 (N_307,In_1588,N_158);
or U308 (N_308,In_2501,In_378);
or U309 (N_309,In_1612,In_951);
xor U310 (N_310,In_2832,In_2713);
and U311 (N_311,In_1243,In_651);
nand U312 (N_312,In_2924,In_2884);
or U313 (N_313,In_2916,In_1311);
xor U314 (N_314,In_1338,N_184);
or U315 (N_315,In_935,In_469);
nor U316 (N_316,In_2328,In_1929);
nand U317 (N_317,In_162,In_122);
or U318 (N_318,In_2705,In_248);
and U319 (N_319,In_1175,In_2589);
or U320 (N_320,In_2079,N_3);
or U321 (N_321,In_314,In_1462);
and U322 (N_322,In_2549,In_725);
nor U323 (N_323,In_1465,N_41);
xor U324 (N_324,In_1761,In_830);
xnor U325 (N_325,In_114,In_271);
and U326 (N_326,In_685,In_2830);
nand U327 (N_327,In_1053,In_2283);
nand U328 (N_328,In_2271,In_817);
nor U329 (N_329,In_1167,In_1633);
xnor U330 (N_330,In_2602,In_654);
or U331 (N_331,In_2457,In_234);
xor U332 (N_332,In_2951,In_1161);
or U333 (N_333,In_1219,In_2206);
nand U334 (N_334,In_439,In_2624);
nor U335 (N_335,In_1945,In_2487);
or U336 (N_336,In_2993,In_2186);
nor U337 (N_337,In_891,In_2163);
nor U338 (N_338,In_1415,In_1320);
or U339 (N_339,In_239,In_829);
nand U340 (N_340,In_655,In_297);
xor U341 (N_341,In_1012,In_2356);
nor U342 (N_342,In_2011,In_529);
nor U343 (N_343,In_723,In_1639);
or U344 (N_344,In_2053,In_394);
or U345 (N_345,In_2262,N_47);
nor U346 (N_346,In_919,In_1655);
xnor U347 (N_347,In_166,In_1476);
nor U348 (N_348,In_2545,In_993);
nor U349 (N_349,In_2914,In_364);
xor U350 (N_350,In_1261,In_1729);
nor U351 (N_351,In_2915,In_2219);
nor U352 (N_352,In_1533,In_2933);
or U353 (N_353,In_77,In_538);
and U354 (N_354,In_2161,In_2642);
nor U355 (N_355,In_1249,In_1485);
xnor U356 (N_356,In_1484,In_483);
xor U357 (N_357,In_1479,In_2320);
nand U358 (N_358,In_2780,In_1482);
nor U359 (N_359,In_771,In_2107);
nor U360 (N_360,In_1087,In_1892);
and U361 (N_361,In_2965,In_2413);
xor U362 (N_362,In_1712,In_2009);
nand U363 (N_363,In_2688,N_21);
or U364 (N_364,In_1090,In_2874);
nor U365 (N_365,In_1164,N_25);
nand U366 (N_366,In_1720,In_2778);
xor U367 (N_367,In_2191,In_1963);
or U368 (N_368,In_308,In_2440);
nand U369 (N_369,In_865,In_326);
xor U370 (N_370,In_971,In_1644);
xor U371 (N_371,In_244,N_139);
and U372 (N_372,In_948,In_565);
nor U373 (N_373,In_2365,N_137);
and U374 (N_374,In_942,In_343);
or U375 (N_375,In_1301,In_2336);
or U376 (N_376,In_2408,In_1001);
xnor U377 (N_377,In_375,In_1016);
nor U378 (N_378,In_2516,In_2870);
nor U379 (N_379,In_424,In_1152);
xor U380 (N_380,In_2668,In_2825);
nand U381 (N_381,In_1767,In_508);
xnor U382 (N_382,In_459,In_2279);
or U383 (N_383,In_299,In_2695);
nand U384 (N_384,In_1394,In_2118);
and U385 (N_385,N_100,In_1337);
nor U386 (N_386,In_1489,N_186);
xor U387 (N_387,In_1969,In_1917);
and U388 (N_388,In_722,In_1019);
nand U389 (N_389,In_2717,In_2171);
or U390 (N_390,In_2226,In_10);
nor U391 (N_391,In_2131,In_1985);
and U392 (N_392,In_2468,In_1033);
nor U393 (N_393,In_2621,In_953);
or U394 (N_394,In_412,In_1614);
or U395 (N_395,In_2659,In_849);
nand U396 (N_396,In_2848,In_1443);
and U397 (N_397,In_28,In_2489);
nand U398 (N_398,In_2039,In_904);
xnor U399 (N_399,In_1182,In_1124);
xnor U400 (N_400,In_683,In_945);
xor U401 (N_401,In_1666,In_983);
nor U402 (N_402,In_2001,N_19);
nor U403 (N_403,In_1036,In_2429);
or U404 (N_404,In_2819,N_94);
or U405 (N_405,In_1657,In_663);
nor U406 (N_406,In_74,In_2231);
and U407 (N_407,In_2797,In_1100);
nor U408 (N_408,In_279,In_721);
nand U409 (N_409,N_249,In_2337);
and U410 (N_410,In_1123,In_875);
or U411 (N_411,In_930,N_171);
xnor U412 (N_412,In_834,In_699);
and U413 (N_413,In_1209,In_1058);
xor U414 (N_414,In_2726,N_113);
nand U415 (N_415,In_2444,In_2833);
or U416 (N_416,In_2101,N_8);
nor U417 (N_417,In_1192,In_2075);
xor U418 (N_418,In_1403,In_2417);
and U419 (N_419,In_2218,N_360);
or U420 (N_420,In_2178,In_1926);
and U421 (N_421,In_940,In_534);
and U422 (N_422,N_337,N_44);
nor U423 (N_423,In_1622,N_187);
or U424 (N_424,In_2850,In_1168);
xnor U425 (N_425,In_1807,In_1779);
and U426 (N_426,In_416,In_2431);
nand U427 (N_427,In_1488,In_1957);
nor U428 (N_428,N_268,In_2939);
xnor U429 (N_429,In_2,In_2708);
xor U430 (N_430,N_277,In_1968);
xnor U431 (N_431,In_1181,In_71);
nand U432 (N_432,In_2599,In_2732);
nand U433 (N_433,N_282,In_1875);
or U434 (N_434,In_235,In_1907);
xor U435 (N_435,In_2922,In_1648);
or U436 (N_436,In_868,In_2452);
and U437 (N_437,In_2603,In_2280);
or U438 (N_438,In_745,In_839);
xor U439 (N_439,In_1195,In_435);
xor U440 (N_440,In_400,In_2380);
or U441 (N_441,In_2510,In_1901);
or U442 (N_442,In_286,In_1409);
xnor U443 (N_443,In_1669,N_310);
xnor U444 (N_444,In_2834,In_2753);
and U445 (N_445,N_27,In_776);
and U446 (N_446,In_2663,In_1659);
nand U447 (N_447,In_2331,N_57);
and U448 (N_448,N_276,In_1855);
or U449 (N_449,In_377,In_2561);
or U450 (N_450,In_2129,N_63);
or U451 (N_451,In_269,In_236);
xnor U452 (N_452,In_2307,In_2018);
or U453 (N_453,In_2088,In_1852);
nor U454 (N_454,N_220,In_273);
or U455 (N_455,N_221,In_1324);
nor U456 (N_456,In_2335,In_2565);
xnor U457 (N_457,In_402,In_2112);
nor U458 (N_458,In_514,In_455);
nor U459 (N_459,In_2706,In_1171);
and U460 (N_460,In_697,In_2427);
xnor U461 (N_461,In_2077,In_1148);
and U462 (N_462,In_1134,N_16);
xnor U463 (N_463,N_0,N_233);
nand U464 (N_464,In_91,In_1738);
nor U465 (N_465,In_2768,In_836);
or U466 (N_466,In_413,In_1131);
nor U467 (N_467,In_194,In_1135);
nor U468 (N_468,N_228,In_2693);
nor U469 (N_469,In_857,In_323);
or U470 (N_470,In_952,N_23);
nand U471 (N_471,In_371,In_802);
xnor U472 (N_472,In_2420,In_2514);
and U473 (N_473,In_519,In_2375);
xnor U474 (N_474,In_2964,In_2696);
and U475 (N_475,In_2221,In_127);
nand U476 (N_476,In_1694,In_2090);
and U477 (N_477,N_114,In_1003);
or U478 (N_478,In_1141,In_125);
and U479 (N_479,In_1608,N_29);
nand U480 (N_480,In_717,In_943);
xor U481 (N_481,In_862,In_452);
xor U482 (N_482,In_329,In_2350);
nor U483 (N_483,In_2478,In_1046);
and U484 (N_484,In_2704,In_2471);
or U485 (N_485,In_467,In_2973);
or U486 (N_486,In_1806,In_1317);
xnor U487 (N_487,In_69,N_236);
nor U488 (N_488,In_2287,In_1775);
nand U489 (N_489,In_844,N_152);
or U490 (N_490,In_1794,In_2415);
nor U491 (N_491,In_226,In_1405);
xnor U492 (N_492,In_1410,In_1071);
nor U493 (N_493,In_1772,N_5);
nor U494 (N_494,In_869,In_1640);
nand U495 (N_495,In_1467,In_1067);
or U496 (N_496,In_2701,In_1078);
nand U497 (N_497,In_120,In_2387);
and U498 (N_498,In_1760,In_743);
nor U499 (N_499,In_1490,In_107);
xor U500 (N_500,In_1006,In_1511);
nand U501 (N_501,N_376,In_2937);
and U502 (N_502,In_2794,In_2263);
or U503 (N_503,In_265,In_2405);
and U504 (N_504,In_2153,In_532);
xnor U505 (N_505,In_2492,In_135);
or U506 (N_506,In_302,In_2136);
or U507 (N_507,In_1323,In_284);
xor U508 (N_508,In_53,In_1764);
or U509 (N_509,In_359,N_130);
or U510 (N_510,In_2847,In_2995);
nand U511 (N_511,In_1922,In_1457);
xnor U512 (N_512,In_798,In_2941);
and U513 (N_513,N_170,In_2459);
xnor U514 (N_514,In_2216,N_314);
nor U515 (N_515,In_1526,In_1025);
and U516 (N_516,N_80,In_2448);
or U517 (N_517,In_1294,In_701);
or U518 (N_518,In_352,In_2035);
and U519 (N_519,In_962,In_2465);
nor U520 (N_520,N_126,In_1857);
xnor U521 (N_521,In_1524,In_1336);
and U522 (N_522,In_1024,In_2923);
nor U523 (N_523,In_956,In_2811);
or U524 (N_524,In_1449,In_1335);
nor U525 (N_525,In_1944,In_1769);
or U526 (N_526,In_165,In_1774);
and U527 (N_527,N_350,N_211);
and U528 (N_528,In_2752,In_769);
and U529 (N_529,In_1102,In_2725);
nand U530 (N_530,In_32,In_2647);
nand U531 (N_531,In_2396,In_1235);
or U532 (N_532,In_1066,In_405);
nand U533 (N_533,In_1269,In_288);
nor U534 (N_534,In_734,In_1352);
nor U535 (N_535,In_2292,In_178);
xor U536 (N_536,In_1933,In_2528);
and U537 (N_537,In_1501,In_1319);
nand U538 (N_538,In_980,In_1713);
or U539 (N_539,N_125,In_583);
nand U540 (N_540,In_766,N_283);
and U541 (N_541,In_395,In_304);
nor U542 (N_542,In_465,In_1382);
or U543 (N_543,N_185,In_60);
nand U544 (N_544,N_374,In_944);
or U545 (N_545,In_1005,In_121);
xor U546 (N_546,In_2905,N_331);
or U547 (N_547,In_383,In_1459);
nand U548 (N_548,N_39,In_1592);
nor U549 (N_549,In_2286,In_247);
or U550 (N_550,In_2826,In_622);
and U551 (N_551,In_2348,In_1973);
and U552 (N_552,In_2062,N_182);
and U553 (N_553,In_2845,In_1);
nand U554 (N_554,N_252,N_115);
nand U555 (N_555,In_2467,In_2063);
xnor U556 (N_556,In_1373,In_540);
nor U557 (N_557,In_2853,In_1049);
or U558 (N_558,In_2852,N_74);
or U559 (N_559,In_978,In_33);
xnor U560 (N_560,In_2352,In_2749);
xor U561 (N_561,In_252,In_2470);
xor U562 (N_562,In_1813,In_1013);
xnor U563 (N_563,In_2080,In_1119);
nor U564 (N_564,In_2126,In_2342);
xnor U565 (N_565,In_1241,In_213);
or U566 (N_566,In_2672,In_644);
nand U567 (N_567,N_271,In_2447);
nand U568 (N_568,In_222,In_2908);
and U569 (N_569,In_1804,In_444);
nor U570 (N_570,N_383,N_109);
nor U571 (N_571,In_1531,In_2572);
nand U572 (N_572,In_975,In_2439);
xor U573 (N_573,N_45,In_1206);
nand U574 (N_574,N_58,In_1417);
xor U575 (N_575,In_637,N_306);
and U576 (N_576,In_2488,N_129);
nor U577 (N_577,In_1486,In_296);
nand U578 (N_578,In_153,In_1105);
and U579 (N_579,In_1831,N_224);
nor U580 (N_580,In_2495,In_1808);
nor U581 (N_581,N_355,In_403);
and U582 (N_582,In_1846,In_1514);
xnor U583 (N_583,In_1231,N_375);
or U584 (N_584,In_1306,In_2976);
and U585 (N_585,N_342,In_2203);
nand U586 (N_586,In_2295,In_14);
and U587 (N_587,In_1127,In_1561);
nor U588 (N_588,In_1842,In_3);
or U589 (N_589,In_1029,In_437);
nand U590 (N_590,In_740,In_2176);
nand U591 (N_591,In_630,In_2871);
xor U592 (N_592,In_575,In_2985);
xnor U593 (N_593,In_1637,In_2082);
nor U594 (N_594,In_2633,In_1156);
and U595 (N_595,In_600,In_168);
and U596 (N_596,In_1387,In_2247);
nor U597 (N_597,In_2673,In_55);
nor U598 (N_598,In_1811,In_2507);
nand U599 (N_599,In_2050,In_1447);
nor U600 (N_600,In_1179,In_1566);
or U601 (N_601,N_327,In_1571);
nor U602 (N_602,In_1553,In_526);
xor U603 (N_603,N_259,In_2268);
nand U604 (N_604,In_363,In_65);
and U605 (N_605,N_308,N_367);
and U606 (N_606,N_61,N_104);
nand U607 (N_607,In_577,In_2731);
nand U608 (N_608,In_305,In_2384);
nand U609 (N_609,In_1234,In_1707);
xor U610 (N_610,In_946,In_1055);
xnor U611 (N_611,In_553,In_2593);
nand U612 (N_612,In_1045,N_359);
nor U613 (N_613,In_2782,N_312);
and U614 (N_614,In_970,In_97);
nand U615 (N_615,In_855,N_215);
and U616 (N_616,In_2581,In_151);
nand U617 (N_617,In_1297,In_2512);
and U618 (N_618,In_2037,In_2180);
and U619 (N_619,In_2409,In_2148);
xor U620 (N_620,In_2275,In_505);
nor U621 (N_621,N_580,In_1733);
nand U622 (N_622,In_150,In_2181);
and U623 (N_623,In_2390,In_1452);
or U624 (N_624,In_2197,N_150);
nor U625 (N_625,In_1155,N_551);
nand U626 (N_626,In_1445,In_1370);
nand U627 (N_627,In_1412,In_2894);
xor U628 (N_628,In_1191,In_1481);
and U629 (N_629,In_2097,In_604);
xnor U630 (N_630,N_499,N_213);
or U631 (N_631,In_98,N_112);
and U632 (N_632,N_32,N_561);
nand U633 (N_633,N_444,In_427);
nand U634 (N_634,In_355,N_322);
xnor U635 (N_635,N_101,In_489);
nand U636 (N_636,In_1685,In_1581);
nor U637 (N_637,In_1966,In_900);
or U638 (N_638,In_2983,In_174);
nor U639 (N_639,In_719,N_409);
and U640 (N_640,In_1618,N_281);
and U641 (N_641,In_741,In_2276);
xor U642 (N_642,In_2223,In_1376);
or U643 (N_643,In_1429,In_2110);
xnor U644 (N_644,In_2840,In_2737);
nor U645 (N_645,N_324,In_1166);
nand U646 (N_646,N_77,In_409);
and U647 (N_647,In_223,In_1890);
nand U648 (N_648,In_939,In_39);
nor U649 (N_649,In_1965,N_378);
xor U650 (N_650,N_34,In_1752);
nand U651 (N_651,In_969,In_388);
nand U652 (N_652,In_2927,In_2573);
xor U653 (N_653,In_376,In_761);
nor U654 (N_654,In_1658,In_2626);
nand U655 (N_655,In_221,In_2554);
nor U656 (N_656,In_1461,In_277);
xnor U657 (N_657,N_386,In_2149);
or U658 (N_658,In_828,In_731);
nor U659 (N_659,In_1914,In_2754);
nand U660 (N_660,N_218,In_518);
nor U661 (N_661,In_2055,In_1757);
nor U662 (N_662,In_1606,N_140);
nand U663 (N_663,N_10,In_2463);
xor U664 (N_664,In_1959,In_1368);
xnor U665 (N_665,In_2616,N_189);
nor U666 (N_666,In_2379,In_2547);
nand U667 (N_667,In_472,In_2636);
nand U668 (N_668,N_470,In_1129);
or U669 (N_669,In_640,In_2795);
nand U670 (N_670,In_1879,In_835);
or U671 (N_671,N_301,N_73);
and U672 (N_672,In_758,N_575);
and U673 (N_673,N_505,In_2891);
or U674 (N_674,In_2434,N_398);
nor U675 (N_675,In_602,In_2943);
and U676 (N_676,In_1117,In_2259);
nor U677 (N_677,In_1237,In_2998);
and U678 (N_678,In_2207,In_2143);
or U679 (N_679,In_1230,In_1178);
or U680 (N_680,In_40,In_658);
nor U681 (N_681,In_496,In_2950);
nand U682 (N_682,In_556,N_181);
and U683 (N_683,In_330,In_2948);
nor U684 (N_684,N_153,In_473);
xor U685 (N_685,N_460,In_562);
nor U686 (N_686,In_1363,In_380);
xnor U687 (N_687,In_2113,In_2893);
nand U688 (N_688,In_2085,In_750);
or U689 (N_689,N_379,In_2680);
nor U690 (N_690,In_2984,In_754);
nand U691 (N_691,In_2517,In_1339);
nor U692 (N_692,N_486,In_1202);
xor U693 (N_693,In_2430,In_87);
or U694 (N_694,In_774,In_1918);
or U695 (N_695,In_2313,N_201);
and U696 (N_696,In_936,In_1193);
nor U697 (N_697,In_2182,In_2288);
nor U698 (N_698,N_33,In_816);
xnor U699 (N_699,In_1424,In_1035);
and U700 (N_700,In_103,In_1086);
nor U701 (N_701,In_1953,In_700);
nor U702 (N_702,In_1063,In_2767);
and U703 (N_703,In_2255,In_2422);
and U704 (N_704,In_513,In_1480);
and U705 (N_705,In_313,N_287);
nor U706 (N_706,In_2237,In_2926);
nand U707 (N_707,In_429,N_90);
xnor U708 (N_708,In_2873,In_2533);
xor U709 (N_709,In_1173,In_238);
nor U710 (N_710,In_1854,In_594);
nor U711 (N_711,In_393,In_1530);
nand U712 (N_712,N_382,In_2758);
nor U713 (N_713,In_2785,N_138);
xor U714 (N_714,In_356,In_1847);
xor U715 (N_715,In_280,N_89);
and U716 (N_716,In_1280,In_484);
and U717 (N_717,In_2392,In_2580);
nor U718 (N_718,N_368,In_592);
nand U719 (N_719,In_831,In_584);
and U720 (N_720,In_1613,N_43);
or U721 (N_721,In_2643,N_530);
nor U722 (N_722,In_1434,In_2046);
or U723 (N_723,In_2585,In_2604);
xnor U724 (N_724,In_205,In_2958);
and U725 (N_725,N_162,In_1040);
nor U726 (N_726,In_2187,In_609);
nor U727 (N_727,In_2388,In_2213);
and U728 (N_728,N_148,In_2274);
nor U729 (N_729,In_436,In_309);
xor U730 (N_730,In_2435,N_535);
xnor U731 (N_731,In_510,In_464);
nand U732 (N_732,In_2252,N_103);
and U733 (N_733,In_1133,In_2920);
xor U734 (N_734,In_262,In_2460);
nor U735 (N_735,In_1441,In_2660);
nand U736 (N_736,N_40,N_231);
nor U737 (N_737,N_265,In_1971);
nand U738 (N_738,N_387,In_1220);
and U739 (N_739,N_543,In_2543);
and U740 (N_740,In_434,In_595);
and U741 (N_741,In_1262,In_1509);
and U742 (N_742,In_1731,In_982);
nor U743 (N_743,In_2265,In_1503);
xnor U744 (N_744,In_515,In_548);
or U745 (N_745,N_363,In_1216);
or U746 (N_746,In_2583,In_1259);
or U747 (N_747,In_1162,In_2499);
or U748 (N_748,N_267,In_35);
and U749 (N_749,In_1869,In_16);
xor U750 (N_750,In_2857,In_917);
or U751 (N_751,In_479,In_351);
nor U752 (N_752,In_1506,In_906);
and U753 (N_753,N_484,In_1010);
and U754 (N_754,In_1454,In_977);
and U755 (N_755,N_258,In_665);
nand U756 (N_756,In_2442,In_1223);
xor U757 (N_757,In_474,In_520);
or U758 (N_758,In_1183,In_1236);
or U759 (N_759,In_300,In_2525);
nand U760 (N_760,N_559,In_1913);
or U761 (N_761,In_2828,In_229);
and U762 (N_762,N_11,In_2266);
xor U763 (N_763,N_582,In_2185);
and U764 (N_764,In_2294,In_624);
and U765 (N_765,In_2065,In_616);
nand U766 (N_766,N_289,In_1638);
nor U767 (N_767,In_295,In_530);
or U768 (N_768,In_1310,In_2617);
nand U769 (N_769,In_527,In_1709);
nor U770 (N_770,N_59,In_1889);
xor U771 (N_771,In_1838,In_2722);
or U772 (N_772,In_2056,In_1732);
nand U773 (N_773,N_515,In_1996);
nor U774 (N_774,N_333,In_1596);
or U775 (N_775,N_442,In_1218);
nor U776 (N_776,In_2959,In_1800);
or U777 (N_777,In_1199,N_169);
or U778 (N_778,In_2770,In_1827);
xnor U779 (N_779,In_1791,In_1522);
xor U780 (N_780,In_2724,In_1625);
and U781 (N_781,In_591,In_2166);
or U782 (N_782,In_1876,In_1008);
nor U783 (N_783,In_2071,In_920);
and U784 (N_784,In_1264,In_2579);
or U785 (N_785,N_116,In_2366);
xnor U786 (N_786,In_1583,In_642);
nand U787 (N_787,In_382,In_281);
xnor U788 (N_788,In_52,In_2446);
or U789 (N_789,N_573,In_495);
or U790 (N_790,N_452,In_2222);
or U791 (N_791,In_2326,In_1426);
xor U792 (N_792,In_2338,In_1573);
and U793 (N_793,N_412,In_111);
nor U794 (N_794,In_2801,N_7);
xor U795 (N_795,In_927,N_161);
nor U796 (N_796,In_1499,In_2150);
or U797 (N_797,N_568,In_2319);
nand U798 (N_798,N_401,In_1250);
xor U799 (N_799,In_1122,N_569);
nor U800 (N_800,In_550,N_36);
nand U801 (N_801,In_1790,In_1081);
and U802 (N_802,In_491,N_413);
xor U803 (N_803,N_210,In_559);
or U804 (N_804,In_1568,In_72);
nand U805 (N_805,N_542,In_2904);
nand U806 (N_806,In_2232,In_1805);
xnor U807 (N_807,N_473,In_2771);
xor U808 (N_808,In_2615,In_408);
or U809 (N_809,In_2070,N_274);
nor U810 (N_810,In_2962,In_746);
xor U811 (N_811,In_1746,In_2665);
and U812 (N_812,N_661,In_268);
xnor U813 (N_813,In_209,In_1247);
nor U814 (N_814,In_923,In_270);
nor U815 (N_815,N_288,N_159);
and U816 (N_816,N_426,In_54);
and U817 (N_817,In_2230,N_673);
and U818 (N_818,N_617,In_2103);
and U819 (N_819,N_157,N_145);
or U820 (N_820,N_416,N_136);
xor U821 (N_821,N_780,In_160);
nor U822 (N_822,In_791,In_738);
xnor U823 (N_823,In_2278,N_443);
nor U824 (N_824,N_453,In_2078);
nand U825 (N_825,In_2837,In_1084);
xor U826 (N_826,In_974,In_788);
or U827 (N_827,In_2109,In_2946);
nand U828 (N_828,N_421,N_712);
and U829 (N_829,In_319,In_2736);
and U830 (N_830,In_1120,In_1961);
nor U831 (N_831,In_1621,N_584);
xor U832 (N_832,In_457,N_253);
nand U833 (N_833,In_2019,N_472);
xor U834 (N_834,In_2864,N_595);
or U835 (N_835,In_200,In_470);
xor U836 (N_836,N_776,N_381);
xnor U837 (N_837,In_2899,In_2484);
or U838 (N_838,In_241,N_631);
or U839 (N_839,N_740,In_414);
xor U840 (N_840,In_1369,N_165);
and U841 (N_841,N_419,N_475);
nand U842 (N_842,In_918,In_2483);
nand U843 (N_843,In_2808,In_1602);
xor U844 (N_844,In_159,In_2212);
and U845 (N_845,In_1273,In_2127);
or U846 (N_846,In_163,N_430);
nor U847 (N_847,In_2534,In_854);
nand U848 (N_848,In_2667,In_2412);
nor U849 (N_849,In_2608,In_339);
nand U850 (N_850,In_1322,In_2068);
xnor U851 (N_851,In_1468,In_1819);
or U852 (N_852,N_464,In_573);
or U853 (N_853,In_2625,N_279);
or U854 (N_854,N_678,In_1307);
nand U855 (N_855,In_925,N_554);
or U856 (N_856,In_2817,In_2759);
nand U857 (N_857,In_1817,In_220);
nor U858 (N_858,In_1248,In_2527);
and U859 (N_859,In_1455,In_2128);
or U860 (N_860,In_2912,In_610);
or U861 (N_861,In_1894,N_710);
and U862 (N_862,In_2815,In_1740);
nor U863 (N_863,N_696,In_894);
and U864 (N_864,In_2367,N_133);
nor U865 (N_865,In_2925,In_254);
and U866 (N_866,In_291,In_2008);
xnor U867 (N_867,N_235,N_407);
nand U868 (N_868,In_1950,In_2846);
or U869 (N_869,In_2816,In_972);
xnor U870 (N_870,N_315,In_2052);
xnor U871 (N_871,In_1650,In_521);
nand U872 (N_872,In_487,In_2955);
nand U873 (N_873,In_1346,N_686);
xnor U874 (N_874,N_128,In_2381);
and U875 (N_875,N_320,In_1309);
xor U876 (N_876,N_86,In_1186);
and U877 (N_877,In_2560,N_238);
nor U878 (N_878,In_1683,In_1803);
or U879 (N_879,In_185,N_305);
xor U880 (N_880,In_2493,In_581);
xor U881 (N_881,N_295,In_1239);
or U882 (N_882,N_732,In_224);
nand U883 (N_883,In_446,In_1828);
nand U884 (N_884,In_2938,In_1205);
xor U885 (N_885,In_2882,N_70);
xnor U886 (N_886,N_798,In_2612);
and U887 (N_887,N_723,N_615);
nand U888 (N_888,N_650,In_303);
nand U889 (N_889,In_1472,In_742);
xnor U890 (N_890,In_1755,N_762);
or U891 (N_891,In_1159,N_50);
xor U892 (N_892,In_214,In_2026);
or U893 (N_893,In_1859,In_1627);
or U894 (N_894,In_1916,N_777);
nand U895 (N_895,N_733,In_1903);
xnor U896 (N_896,N_664,N_175);
nor U897 (N_897,In_1276,In_2812);
xnor U898 (N_898,In_1442,In_1781);
nand U899 (N_899,In_1802,In_2727);
nor U900 (N_900,In_783,In_1861);
nand U901 (N_901,In_1145,N_744);
nor U902 (N_902,In_2100,In_2209);
nor U903 (N_903,In_2538,In_1270);
xor U904 (N_904,In_433,In_1665);
nand U905 (N_905,In_1128,N_448);
xor U906 (N_906,In_1744,N_22);
xnor U907 (N_907,N_621,In_1871);
or U908 (N_908,In_253,In_512);
and U909 (N_909,In_846,In_1974);
nor U910 (N_910,In_606,In_1610);
or U911 (N_911,In_833,In_959);
or U912 (N_912,In_673,In_2023);
xor U913 (N_913,In_310,In_517);
xor U914 (N_914,In_337,In_1849);
nand U915 (N_915,In_1704,In_167);
nor U916 (N_916,N_778,In_1684);
nor U917 (N_917,In_851,In_1587);
nor U918 (N_918,In_585,In_499);
xnor U919 (N_919,N_704,N_49);
nand U920 (N_920,N_24,N_461);
xor U921 (N_921,N_309,In_2628);
nor U922 (N_922,In_391,In_2587);
xnor U923 (N_923,In_76,In_2679);
and U924 (N_924,N_513,In_2410);
and U925 (N_925,In_679,N_578);
and U926 (N_926,In_2859,In_1366);
and U927 (N_927,In_837,N_591);
nand U928 (N_928,In_1938,In_633);
nor U929 (N_929,In_2240,In_2885);
xnor U930 (N_930,In_2363,In_1396);
and U931 (N_931,In_1496,N_270);
nand U932 (N_932,In_2577,In_886);
and U933 (N_933,In_2031,In_1822);
and U934 (N_934,N_414,N_611);
nor U935 (N_935,N_758,In_497);
and U936 (N_936,In_1934,In_1563);
nor U937 (N_937,In_531,N_438);
and U938 (N_938,In_385,In_661);
nor U939 (N_939,In_1165,In_1930);
and U940 (N_940,In_2918,N_76);
nand U941 (N_941,In_2242,In_1289);
nand U942 (N_942,N_726,In_1378);
nor U943 (N_943,In_1754,In_2264);
xnor U944 (N_944,In_660,In_634);
nor U945 (N_945,In_1773,In_1098);
nor U946 (N_946,In_2155,N_106);
or U947 (N_947,In_2786,In_1096);
and U948 (N_948,In_818,In_813);
nand U949 (N_949,N_147,N_394);
nor U950 (N_950,In_804,In_693);
and U951 (N_951,In_2104,In_2172);
and U952 (N_952,N_498,In_389);
nand U953 (N_953,In_1544,In_2789);
and U954 (N_954,In_154,N_338);
xor U955 (N_955,In_2714,In_2862);
or U956 (N_956,In_2605,In_988);
and U957 (N_957,In_2045,N_263);
or U958 (N_958,In_524,N_716);
xor U959 (N_959,N_771,In_2005);
xnor U960 (N_960,In_2803,In_667);
nor U961 (N_961,N_456,In_190);
xor U962 (N_962,In_2793,N_793);
or U963 (N_963,In_2813,In_2896);
or U964 (N_964,N_656,In_113);
or U965 (N_965,In_2233,N_735);
or U966 (N_966,N_449,N_247);
or U967 (N_967,In_1814,In_1089);
or U968 (N_968,N_600,In_100);
or U969 (N_969,In_2480,In_2597);
nand U970 (N_970,In_1636,In_2855);
nor U971 (N_971,In_1952,In_1782);
or U972 (N_972,N_257,In_1874);
and U973 (N_973,N_286,N_300);
xnor U974 (N_974,N_676,In_1265);
nand U975 (N_975,In_2389,In_1143);
xnor U976 (N_976,In_1453,In_963);
or U977 (N_977,In_1597,N_269);
xor U978 (N_978,In_2299,In_2504);
xor U979 (N_979,In_1051,In_327);
and U980 (N_980,In_2716,N_790);
nor U981 (N_981,In_2783,In_1628);
nor U982 (N_982,In_2897,In_481);
nor U983 (N_983,In_2317,In_539);
or U984 (N_984,N_200,In_171);
and U985 (N_985,In_2192,In_468);
xnor U986 (N_986,In_698,N_779);
nor U987 (N_987,N_623,In_2690);
nor U988 (N_988,N_766,In_1516);
and U989 (N_989,N_606,In_1577);
nor U990 (N_990,In_477,In_2042);
and U991 (N_991,In_2270,In_826);
or U992 (N_992,N_658,In_691);
and U993 (N_993,In_808,In_2407);
or U994 (N_994,In_2536,In_2450);
xnor U995 (N_995,In_744,In_2333);
or U996 (N_996,N_772,N_640);
or U997 (N_997,In_1877,In_914);
nand U998 (N_998,N_589,In_2456);
or U999 (N_999,In_785,N_352);
nor U1000 (N_1000,In_2548,N_755);
xnor U1001 (N_1001,In_1002,In_134);
or U1002 (N_1002,In_1140,In_724);
nor U1003 (N_1003,In_2712,N_995);
or U1004 (N_1004,In_231,In_2310);
and U1005 (N_1005,N_46,N_53);
or U1006 (N_1006,In_1508,In_2854);
xnor U1007 (N_1007,In_2173,In_1975);
nand U1008 (N_1008,In_1706,In_1438);
or U1009 (N_1009,N_826,In_203);
or U1010 (N_1010,N_662,N_985);
nand U1011 (N_1011,In_1979,In_915);
nand U1012 (N_1012,In_1909,In_1844);
xor U1013 (N_1013,In_1299,In_228);
and U1014 (N_1014,N_435,In_132);
or U1015 (N_1015,In_1543,In_1690);
nor U1016 (N_1016,N_117,In_759);
nor U1017 (N_1017,In_730,N_402);
xor U1018 (N_1018,In_2322,In_2932);
nor U1019 (N_1019,N_945,N_155);
nor U1020 (N_1020,N_358,In_929);
or U1021 (N_1021,In_2477,In_934);
nor U1022 (N_1022,In_2954,In_760);
nor U1023 (N_1023,N_537,N_692);
and U1024 (N_1024,In_2462,In_1091);
and U1025 (N_1025,In_626,In_1988);
nand U1026 (N_1026,In_2866,N_81);
nand U1027 (N_1027,In_2773,In_907);
nand U1028 (N_1028,In_1418,N_225);
or U1029 (N_1029,N_98,In_842);
nor U1030 (N_1030,N_97,In_1896);
nor U1031 (N_1031,N_567,In_2526);
nand U1032 (N_1032,In_1224,N_845);
xor U1033 (N_1033,N_37,In_225);
nor U1034 (N_1034,In_1735,In_887);
or U1035 (N_1035,N_441,In_2648);
nor U1036 (N_1036,In_2699,In_1330);
nand U1037 (N_1037,In_1562,In_752);
nand U1038 (N_1038,In_2032,In_1848);
nand U1039 (N_1039,N_348,In_2341);
and U1040 (N_1040,In_1989,N_328);
nor U1041 (N_1041,In_2991,In_2061);
nand U1042 (N_1042,N_729,N_550);
and U1043 (N_1043,In_118,In_675);
xor U1044 (N_1044,In_1724,In_1710);
nand U1045 (N_1045,In_131,N_361);
xnor U1046 (N_1046,In_2868,In_2098);
xor U1047 (N_1047,N_690,In_2956);
and U1048 (N_1048,In_2747,In_2521);
xor U1049 (N_1049,N_146,In_353);
nand U1050 (N_1050,N_205,In_2200);
nor U1051 (N_1051,In_406,In_1768);
or U1052 (N_1052,In_1190,In_1812);
and U1053 (N_1053,N_294,N_199);
and U1054 (N_1054,In_2321,N_871);
xor U1055 (N_1055,In_140,N_655);
nand U1056 (N_1056,In_608,In_1654);
nand U1057 (N_1057,N_212,In_2227);
or U1058 (N_1058,In_249,In_542);
nor U1059 (N_1059,In_2502,In_2117);
nand U1060 (N_1060,N_781,In_2054);
xor U1061 (N_1061,N_626,In_1865);
xor U1062 (N_1062,In_961,In_704);
nand U1063 (N_1063,In_2087,In_2697);
nand U1064 (N_1064,In_1047,In_2309);
nor U1065 (N_1065,N_429,In_739);
or U1066 (N_1066,In_2137,In_1196);
and U1067 (N_1067,In_1820,N_657);
and U1068 (N_1068,N_903,In_790);
nand U1069 (N_1069,In_1277,In_2040);
nand U1070 (N_1070,In_2557,In_1292);
and U1071 (N_1071,N_956,In_186);
xnor U1072 (N_1072,N_298,In_50);
nor U1073 (N_1073,N_149,In_79);
xnor U1074 (N_1074,In_1515,N_959);
nand U1075 (N_1075,N_581,In_1904);
xnor U1076 (N_1076,N_822,In_1388);
nor U1077 (N_1077,In_2133,In_1513);
or U1078 (N_1078,N_119,In_2130);
or U1079 (N_1079,In_2662,In_535);
xor U1080 (N_1080,In_1681,N_285);
nand U1081 (N_1081,N_697,In_2971);
xnor U1082 (N_1082,N_869,In_256);
or U1083 (N_1083,In_2721,N_888);
nor U1084 (N_1084,In_13,In_2179);
nor U1085 (N_1085,N_440,N_641);
nor U1086 (N_1086,In_2334,In_1365);
or U1087 (N_1087,In_1920,In_801);
and U1088 (N_1088,N_17,In_1115);
or U1089 (N_1089,In_809,In_1018);
or U1090 (N_1090,N_701,In_2135);
xor U1091 (N_1091,N_986,N_492);
or U1092 (N_1092,N_434,In_1398);
and U1093 (N_1093,In_1221,N_639);
and U1094 (N_1094,In_1151,In_1079);
xnor U1095 (N_1095,In_2919,N_770);
nor U1096 (N_1096,N_739,In_596);
and U1097 (N_1097,In_613,N_278);
nand U1098 (N_1098,In_672,In_2165);
or U1099 (N_1099,In_1519,In_1843);
or U1100 (N_1100,In_825,N_761);
xnor U1101 (N_1101,In_1668,N_998);
nor U1102 (N_1102,In_158,In_2393);
xor U1103 (N_1103,In_2694,N_748);
or U1104 (N_1104,In_563,N_721);
nand U1105 (N_1105,N_354,In_2190);
nor U1106 (N_1106,N_613,N_67);
and U1107 (N_1107,In_2907,In_1343);
nand U1108 (N_1108,In_89,N_240);
or U1109 (N_1109,In_357,N_932);
nand U1110 (N_1110,N_944,In_2386);
nor U1111 (N_1111,N_370,In_631);
and U1112 (N_1112,N_183,In_2208);
and U1113 (N_1113,N_334,N_773);
nor U1114 (N_1114,In_2989,N_420);
and U1115 (N_1115,N_968,N_994);
or U1116 (N_1116,N_722,In_139);
and U1117 (N_1117,N_528,In_1634);
nand U1118 (N_1118,N_713,N_79);
xor U1119 (N_1119,In_164,In_2872);
xnor U1120 (N_1120,N_256,In_1017);
nand U1121 (N_1121,In_2073,N_255);
nand U1122 (N_1122,N_993,N_891);
nor U1123 (N_1123,In_2416,N_297);
nor U1124 (N_1124,N_823,In_2154);
and U1125 (N_1125,In_386,In_133);
nand U1126 (N_1126,In_1358,N_272);
and U1127 (N_1127,In_2194,N_605);
and U1128 (N_1128,In_2305,N_536);
and U1129 (N_1129,N_803,In_2059);
nor U1130 (N_1130,In_2433,In_276);
and U1131 (N_1131,In_636,In_860);
and U1132 (N_1132,N_326,N_990);
and U1133 (N_1133,In_612,N_132);
and U1134 (N_1134,N_51,In_1400);
xor U1135 (N_1135,In_1984,N_418);
nor U1136 (N_1136,In_898,In_191);
or U1137 (N_1137,N_964,In_882);
or U1138 (N_1138,N_347,N_981);
and U1139 (N_1139,In_1268,N_763);
nand U1140 (N_1140,N_390,In_2974);
nor U1141 (N_1141,In_1180,N_511);
or U1142 (N_1142,In_1390,In_2677);
nor U1143 (N_1143,N_565,In_571);
xnor U1144 (N_1144,N_431,N_174);
nor U1145 (N_1145,In_1576,N_476);
and U1146 (N_1146,In_1395,N_178);
and U1147 (N_1147,In_392,N_560);
nand U1148 (N_1148,In_670,In_705);
and U1149 (N_1149,In_2193,N_622);
xor U1150 (N_1150,In_2498,N_899);
nor U1151 (N_1151,In_206,N_217);
nor U1152 (N_1152,In_1194,In_2999);
and U1153 (N_1153,In_1367,In_169);
nor U1154 (N_1154,N_970,In_407);
xnor U1155 (N_1155,In_872,N_107);
or U1156 (N_1156,N_675,N_56);
nor U1157 (N_1157,In_2777,N_245);
or U1158 (N_1158,In_2745,In_1835);
nor U1159 (N_1159,In_1672,In_2491);
nor U1160 (N_1160,N_592,N_574);
nor U1161 (N_1161,In_832,In_176);
nor U1162 (N_1162,In_488,In_910);
nand U1163 (N_1163,N_479,In_2775);
xor U1164 (N_1164,N_275,In_1815);
or U1165 (N_1165,N_93,N_843);
xor U1166 (N_1166,In_149,In_2183);
nand U1167 (N_1167,In_1572,In_2198);
nor U1168 (N_1168,In_2623,In_2829);
or U1169 (N_1169,N_404,In_2790);
nor U1170 (N_1170,N_760,In_2566);
xnor U1171 (N_1171,N_66,In_130);
nor U1172 (N_1172,N_556,In_1384);
and U1173 (N_1173,N_585,In_1883);
xnor U1174 (N_1174,N_931,In_2844);
nand U1175 (N_1175,In_1885,In_773);
nor U1176 (N_1176,N_901,In_282);
and U1177 (N_1177,N_135,In_1651);
xnor U1178 (N_1178,In_502,In_2358);
or U1179 (N_1179,In_422,N_457);
xor U1180 (N_1180,In_677,In_123);
or U1181 (N_1181,In_703,In_250);
nand U1182 (N_1182,N_877,N_693);
xor U1183 (N_1183,N_459,In_1433);
nor U1184 (N_1184,In_1427,N_737);
nor U1185 (N_1185,In_301,In_2715);
xnor U1186 (N_1186,In_2156,In_2821);
xor U1187 (N_1187,N_424,In_570);
xnor U1188 (N_1188,In_2571,In_2076);
nor U1189 (N_1189,In_2755,N_923);
nor U1190 (N_1190,In_2556,N_494);
and U1191 (N_1191,In_560,In_1691);
nand U1192 (N_1192,In_432,In_645);
nand U1193 (N_1193,In_117,In_1172);
or U1194 (N_1194,In_1990,In_2947);
xnor U1195 (N_1195,In_1244,In_1747);
or U1196 (N_1196,In_781,In_237);
and U1197 (N_1197,N_915,In_764);
xnor U1198 (N_1198,In_1881,In_2298);
xnor U1199 (N_1199,N_329,N_193);
and U1200 (N_1200,N_1110,N_6);
nor U1201 (N_1201,In_1430,N_408);
and U1202 (N_1202,N_251,In_2707);
nand U1203 (N_1203,N_828,N_1050);
xor U1204 (N_1204,N_689,N_850);
nor U1205 (N_1205,N_48,N_516);
and U1206 (N_1206,In_2125,N_356);
nor U1207 (N_1207,In_1565,N_1097);
nor U1208 (N_1208,N_466,In_1792);
and U1209 (N_1209,In_2613,In_1279);
nand U1210 (N_1210,In_2949,N_313);
or U1211 (N_1211,N_495,In_2067);
or U1212 (N_1212,In_2038,In_1629);
or U1213 (N_1213,In_272,In_1703);
and U1214 (N_1214,In_2537,In_2345);
and U1215 (N_1215,N_714,N_563);
xnor U1216 (N_1216,In_1725,N_680);
xnor U1217 (N_1217,N_745,In_2552);
xor U1218 (N_1218,N_173,In_2473);
and U1219 (N_1219,In_181,In_2364);
nor U1220 (N_1220,In_767,In_840);
xnor U1221 (N_1221,N_756,N_1078);
xnor U1222 (N_1222,In_1088,In_1342);
nand U1223 (N_1223,N_1139,N_980);
and U1224 (N_1224,In_1421,In_1189);
and U1225 (N_1225,N_502,In_442);
and U1226 (N_1226,In_1693,N_805);
nor U1227 (N_1227,In_1437,In_2353);
or U1228 (N_1228,N_250,N_610);
and U1229 (N_1229,N_711,In_2437);
nand U1230 (N_1230,In_2202,In_552);
and U1231 (N_1231,N_751,N_936);
xnor U1232 (N_1232,In_1960,N_1018);
nor U1233 (N_1233,In_1295,In_903);
or U1234 (N_1234,In_1099,N_503);
and U1235 (N_1235,N_1121,N_1129);
nor U1236 (N_1236,In_1721,N_1100);
xnor U1237 (N_1237,In_1558,In_1015);
and U1238 (N_1238,In_2102,N_364);
or U1239 (N_1239,In_2692,N_1000);
nor U1240 (N_1240,In_1139,N_812);
nand U1241 (N_1241,N_728,N_609);
nor U1242 (N_1242,N_765,In_2248);
and U1243 (N_1243,N_1181,In_1783);
xor U1244 (N_1244,N_458,In_145);
xnor U1245 (N_1245,N_806,N_1015);
nand U1246 (N_1246,N_1021,In_1785);
and U1247 (N_1247,N_596,In_728);
nand U1248 (N_1248,In_1399,In_895);
xnor U1249 (N_1249,In_410,In_992);
or U1250 (N_1250,N_4,In_662);
nor U1251 (N_1251,In_2015,In_2301);
nand U1252 (N_1252,N_517,N_369);
and U1253 (N_1253,In_2260,In_2340);
xnor U1254 (N_1254,N_950,N_972);
nor U1255 (N_1255,N_996,In_2630);
or U1256 (N_1256,N_852,In_152);
nor U1257 (N_1257,In_1927,N_1094);
nor U1258 (N_1258,N_886,In_2033);
xnor U1259 (N_1259,In_1101,In_1591);
xnor U1260 (N_1260,In_666,In_960);
and U1261 (N_1261,In_294,In_999);
or U1262 (N_1262,In_2119,In_1290);
and U1263 (N_1263,N_496,N_1164);
nand U1264 (N_1264,N_1082,In_2254);
nand U1265 (N_1265,In_2124,In_2147);
xor U1266 (N_1266,In_504,In_1328);
or U1267 (N_1267,N_1077,N_824);
and U1268 (N_1268,In_1321,N_280);
or U1269 (N_1269,N_1099,In_1389);
nor U1270 (N_1270,In_2414,N_887);
xor U1271 (N_1271,In_1554,In_1799);
nor U1272 (N_1272,In_201,N_1143);
or U1273 (N_1273,N_570,In_1937);
and U1274 (N_1274,In_2145,N_918);
xnor U1275 (N_1275,In_1682,N_1103);
xnor U1276 (N_1276,In_1759,In_876);
xnor U1277 (N_1277,In_845,In_240);
or U1278 (N_1278,N_642,In_2158);
nand U1279 (N_1279,In_1891,In_708);
nor U1280 (N_1280,In_2901,N_612);
or U1281 (N_1281,In_1064,N_924);
nor U1282 (N_1282,In_2574,In_369);
or U1283 (N_1283,N_749,In_51);
and U1284 (N_1284,N_427,In_847);
xor U1285 (N_1285,N_1131,In_806);
nand U1286 (N_1286,N_1151,N_841);
nor U1287 (N_1287,In_2315,In_1631);
or U1288 (N_1288,In_2652,N_1061);
and U1289 (N_1289,N_873,N_1136);
xnor U1290 (N_1290,N_332,N_1132);
nand U1291 (N_1291,In_2411,In_2096);
nand U1292 (N_1292,In_2977,In_2761);
and U1293 (N_1293,In_1517,In_1887);
or U1294 (N_1294,In_2744,N_1059);
nor U1295 (N_1295,In_2711,N_651);
or U1296 (N_1296,In_671,In_274);
nand U1297 (N_1297,N_141,In_1697);
nand U1298 (N_1298,In_2841,In_2509);
or U1299 (N_1299,N_789,In_2196);
xnor U1300 (N_1300,In_2698,N_317);
and U1301 (N_1301,N_436,In_445);
and U1302 (N_1302,In_2169,N_727);
xnor U1303 (N_1303,In_1993,In_2297);
xor U1304 (N_1304,N_1072,In_2551);
nand U1305 (N_1305,In_1605,In_1304);
and U1306 (N_1306,N_791,N_1149);
nand U1307 (N_1307,N_853,In_726);
nand U1308 (N_1308,N_1062,In_2558);
or U1309 (N_1309,N_648,N_666);
xnor U1310 (N_1310,N_685,N_669);
xnor U1311 (N_1311,In_2007,In_2164);
nor U1312 (N_1312,N_562,N_223);
xor U1313 (N_1313,In_2682,In_43);
nand U1314 (N_1314,In_109,N_1054);
xnor U1315 (N_1315,N_14,In_1093);
and U1316 (N_1316,N_699,In_2564);
or U1317 (N_1317,N_468,N_999);
or U1318 (N_1318,N_311,N_1193);
or U1319 (N_1319,N_679,In_1254);
nand U1320 (N_1320,N_741,In_148);
xnor U1321 (N_1321,In_784,In_780);
and U1322 (N_1322,N_195,In_2423);
xor U1323 (N_1323,N_1083,In_1956);
and U1324 (N_1324,N_821,In_492);
and U1325 (N_1325,In_1251,In_913);
or U1326 (N_1326,In_2159,In_2851);
nand U1327 (N_1327,In_322,N_1071);
or U1328 (N_1328,N_237,N_965);
or U1329 (N_1329,N_786,In_2028);
or U1330 (N_1330,N_491,In_2733);
and U1331 (N_1331,In_853,In_1845);
xnor U1332 (N_1332,In_311,In_643);
and U1333 (N_1333,In_321,N_652);
nand U1334 (N_1334,In_1548,In_1163);
nor U1335 (N_1335,In_67,N_105);
nand U1336 (N_1336,In_2723,N_177);
xnor U1337 (N_1337,In_2879,N_1126);
xnor U1338 (N_1338,In_2936,In_1777);
nand U1339 (N_1339,In_29,In_879);
nand U1340 (N_1340,In_2300,N_1197);
or U1341 (N_1341,In_558,In_706);
nor U1342 (N_1342,In_884,N_1048);
nand U1343 (N_1343,In_2047,N_1135);
xor U1344 (N_1344,In_24,In_2541);
nand U1345 (N_1345,N_527,In_346);
or U1346 (N_1346,In_15,In_485);
and U1347 (N_1347,N_634,In_1549);
nor U1348 (N_1348,In_528,N_720);
or U1349 (N_1349,In_136,In_1578);
or U1350 (N_1350,In_1203,N_840);
nand U1351 (N_1351,In_994,N_601);
and U1352 (N_1352,In_827,N_1014);
and U1353 (N_1353,In_2004,In_2968);
nor U1354 (N_1354,N_522,In_2371);
nor U1355 (N_1355,In_2756,In_2929);
or U1356 (N_1356,N_1134,In_2601);
nand U1357 (N_1357,In_909,N_292);
nand U1358 (N_1358,N_510,In_1541);
and U1359 (N_1359,In_549,In_1982);
xor U1360 (N_1360,In_2728,In_420);
nor U1361 (N_1361,N_1024,N_734);
and U1362 (N_1362,In_1635,N_860);
or U1363 (N_1363,In_2972,N_638);
xor U1364 (N_1364,In_399,In_871);
nor U1365 (N_1365,N_817,In_1316);
and U1366 (N_1366,N_784,In_1312);
nor U1367 (N_1367,N_1069,In_501);
xnor U1368 (N_1368,In_1027,N_229);
and U1369 (N_1369,In_1652,N_928);
or U1370 (N_1370,N_54,In_2454);
nor U1371 (N_1371,In_2238,In_1284);
or U1372 (N_1372,N_677,In_143);
xnor U1373 (N_1373,In_1987,N_1175);
nor U1374 (N_1374,N_795,In_1362);
nand U1375 (N_1375,In_1567,In_1750);
nor U1376 (N_1376,In_1579,N_810);
xnor U1377 (N_1377,In_1108,In_1776);
nor U1378 (N_1378,N_538,In_2224);
and U1379 (N_1379,N_671,In_2312);
and U1380 (N_1380,N_757,In_1381);
nor U1381 (N_1381,In_639,In_128);
nand U1382 (N_1382,In_8,N_91);
and U1383 (N_1383,In_1258,In_374);
nor U1384 (N_1384,N_500,In_712);
and U1385 (N_1385,In_2086,In_786);
xnor U1386 (N_1386,In_259,In_681);
xor U1387 (N_1387,N_230,In_680);
or U1388 (N_1388,N_507,In_365);
nor U1389 (N_1389,In_1829,In_1675);
xor U1390 (N_1390,In_2506,In_908);
nor U1391 (N_1391,N_227,N_935);
nand U1392 (N_1392,In_1502,In_1745);
nor U1393 (N_1393,In_2351,In_1097);
nor U1394 (N_1394,N_889,In_1075);
xor U1395 (N_1395,N_160,N_880);
nand U1396 (N_1396,In_916,In_2835);
xor U1397 (N_1397,In_1700,In_283);
and U1398 (N_1398,In_94,In_418);
and U1399 (N_1399,In_1308,In_2060);
or U1400 (N_1400,In_1695,In_1340);
or U1401 (N_1401,In_1082,In_1948);
xnor U1402 (N_1402,N_830,In_2316);
nand U1403 (N_1403,In_2293,N_1399);
and U1404 (N_1404,In_757,N_644);
nor U1405 (N_1405,N_1101,In_2640);
or U1406 (N_1406,N_1382,In_546);
xor U1407 (N_1407,N_545,N_1258);
or U1408 (N_1408,N_804,In_421);
nand U1409 (N_1409,N_260,N_813);
xor U1410 (N_1410,In_2025,N_951);
xnor U1411 (N_1411,N_242,N_643);
nand U1412 (N_1412,N_1241,In_18);
xor U1413 (N_1413,In_1217,N_1378);
and U1414 (N_1414,In_1353,N_380);
xor U1415 (N_1415,N_188,N_325);
xor U1416 (N_1416,In_1207,N_940);
nor U1417 (N_1417,In_1104,N_467);
nand U1418 (N_1418,In_245,N_339);
and U1419 (N_1419,N_1085,In_345);
and U1420 (N_1420,In_170,In_1689);
nand U1421 (N_1421,In_1905,N_1167);
xnor U1422 (N_1422,In_2421,N_1068);
xor U1423 (N_1423,N_1269,N_1217);
nor U1424 (N_1424,In_390,In_1245);
nor U1425 (N_1425,N_808,N_389);
and U1426 (N_1426,N_614,In_2609);
and U1427 (N_1427,N_548,N_296);
xnor U1428 (N_1428,In_1538,In_1111);
nand U1429 (N_1429,N_1263,In_112);
nand U1430 (N_1430,N_1228,N_1338);
nor U1431 (N_1431,N_892,N_531);
xor U1432 (N_1432,In_2438,In_1371);
nand U1433 (N_1433,In_523,N_1313);
nand U1434 (N_1434,In_1228,N_1327);
xnor U1435 (N_1435,N_78,N_971);
nor U1436 (N_1436,In_1600,N_1267);
nor U1437 (N_1437,In_1723,N_1205);
xor U1438 (N_1438,N_967,N_1046);
xnor U1439 (N_1439,N_1254,In_2774);
xor U1440 (N_1440,N_846,N_1303);
nand U1441 (N_1441,In_794,N_1344);
nand U1442 (N_1442,In_1753,In_315);
xnor U1443 (N_1443,N_1146,N_571);
xnor U1444 (N_1444,In_2645,N_787);
nand U1445 (N_1445,In_2779,N_977);
or U1446 (N_1446,In_1540,In_2881);
nor U1447 (N_1447,In_702,In_1534);
xor U1448 (N_1448,In_1471,In_2362);
and U1449 (N_1449,N_1342,N_1275);
nor U1450 (N_1450,N_894,In_2750);
nor U1451 (N_1451,In_1895,In_1770);
nor U1452 (N_1452,N_371,N_68);
nand U1453 (N_1453,N_862,In_1431);
xnor U1454 (N_1454,N_415,N_1224);
or U1455 (N_1455,N_1226,In_1660);
and U1456 (N_1456,N_769,N_1109);
nor U1457 (N_1457,N_719,N_839);
xor U1458 (N_1458,N_1385,N_1154);
and U1459 (N_1459,N_1055,N_437);
nor U1460 (N_1460,In_1943,In_1197);
nand U1461 (N_1461,N_1316,In_82);
nand U1462 (N_1462,In_2449,In_2403);
nand U1463 (N_1463,In_989,In_155);
xor U1464 (N_1464,In_1260,N_1251);
nand U1465 (N_1465,N_564,In_2661);
or U1466 (N_1466,In_1615,In_344);
xor U1467 (N_1467,In_1030,N_1178);
nor U1468 (N_1468,In_2476,In_1402);
nand U1469 (N_1469,N_194,In_2058);
xnor U1470 (N_1470,In_2875,N_1340);
and U1471 (N_1471,N_1025,In_1021);
nand U1472 (N_1472,In_2497,N_1105);
nand U1473 (N_1473,N_1089,In_1589);
xor U1474 (N_1474,In_2967,In_2123);
nand U1475 (N_1475,N_800,N_316);
xor U1476 (N_1476,In_1446,In_2014);
or U1477 (N_1477,N_1330,In_462);
or U1478 (N_1478,N_1354,In_2654);
and U1479 (N_1479,In_2261,In_1238);
nand U1480 (N_1480,N_731,N_1079);
nand U1481 (N_1481,N_71,In_498);
or U1482 (N_1482,In_516,In_219);
xor U1483 (N_1483,In_1851,N_284);
nor U1484 (N_1484,In_623,In_2849);
xnor U1485 (N_1485,N_934,N_933);
and U1486 (N_1486,N_764,N_969);
or U1487 (N_1487,N_509,N_1200);
or U1488 (N_1488,In_763,N_1098);
and U1489 (N_1489,N_785,N_197);
xnor U1490 (N_1490,N_1011,In_1915);
xor U1491 (N_1491,In_954,N_1333);
or U1492 (N_1492,In_880,N_875);
nor U1493 (N_1493,In_787,N_937);
and U1494 (N_1494,In_848,In_1525);
nor U1495 (N_1495,N_493,N_1122);
nor U1496 (N_1496,In_1103,N_1063);
xor U1497 (N_1497,N_469,N_1090);
and U1498 (N_1498,N_1300,N_588);
xor U1499 (N_1499,In_1991,N_665);
and U1500 (N_1500,In_260,N_948);
xor U1501 (N_1501,N_1075,In_2030);
xnor U1502 (N_1502,In_1037,N_546);
nor U1503 (N_1503,N_1336,In_1951);
nor U1504 (N_1504,In_1169,N_1111);
and U1505 (N_1505,In_1349,N_1023);
and U1506 (N_1506,In_2619,In_947);
nor U1507 (N_1507,In_2195,N_1119);
or U1508 (N_1508,N_1188,N_234);
nand U1509 (N_1509,N_1266,N_88);
nor U1510 (N_1510,In_31,N_1234);
and U1511 (N_1511,In_1931,N_1140);
nor U1512 (N_1512,In_1300,N_1243);
or U1513 (N_1513,In_1500,N_919);
xor U1514 (N_1514,N_1381,N_480);
nor U1515 (N_1515,In_25,In_507);
nor U1516 (N_1516,N_991,N_814);
nor U1517 (N_1517,In_1673,In_1924);
or U1518 (N_1518,N_385,In_2304);
xnor U1519 (N_1519,N_1260,N_1049);
and U1520 (N_1520,N_1304,N_1306);
or U1521 (N_1521,In_1440,N_1157);
nand U1522 (N_1522,N_1194,In_341);
nor U1523 (N_1523,N_900,In_928);
xor U1524 (N_1524,In_104,N_1233);
nor U1525 (N_1525,N_1211,In_258);
and U1526 (N_1526,In_1921,In_187);
nand U1527 (N_1527,N_1239,In_2889);
and U1528 (N_1528,N_957,In_2838);
nor U1529 (N_1529,In_1092,In_1436);
nand U1530 (N_1530,N_1163,In_1011);
and U1531 (N_1531,In_116,N_481);
or U1532 (N_1532,In_1334,In_1233);
or U1533 (N_1533,In_1470,N_108);
nor U1534 (N_1534,In_335,N_1286);
xnor U1535 (N_1535,N_1076,N_1322);
or U1536 (N_1536,N_910,In_1222);
xnor U1537 (N_1537,In_21,In_1125);
and U1538 (N_1538,In_803,N_586);
xor U1539 (N_1539,In_1545,In_2210);
xor U1540 (N_1540,In_1962,N_1253);
and U1541 (N_1541,In_635,In_456);
nand U1542 (N_1542,In_1972,In_2314);
nor U1543 (N_1543,In_2822,In_2942);
nor U1544 (N_1544,In_1860,In_2474);
or U1545 (N_1545,In_1801,In_735);
and U1546 (N_1546,In_1448,In_2220);
and U1547 (N_1547,N_1345,In_1986);
xnor U1548 (N_1548,N_902,N_1183);
or U1549 (N_1549,N_1291,N_1201);
and U1550 (N_1550,In_1073,N_1114);
xnor U1551 (N_1551,In_2306,In_1048);
and U1552 (N_1552,In_2718,In_1940);
or U1553 (N_1553,In_1551,N_725);
nand U1554 (N_1554,N_1043,In_4);
nand U1555 (N_1555,N_166,In_823);
or U1556 (N_1556,N_1207,N_1360);
or U1557 (N_1557,In_843,In_1528);
and U1558 (N_1558,In_2397,N_1019);
xnor U1559 (N_1559,N_1190,N_1144);
and U1560 (N_1560,In_641,N_653);
xor U1561 (N_1561,In_897,In_883);
or U1562 (N_1562,N_1281,In_2064);
nor U1563 (N_1563,In_2020,N_1231);
nand U1564 (N_1564,In_1664,N_754);
and U1565 (N_1565,N_597,N_423);
and U1566 (N_1566,N_1092,N_533);
xnor U1567 (N_1567,In_12,In_460);
or U1568 (N_1568,N_488,N_393);
nand U1569 (N_1569,In_2324,N_425);
nand U1570 (N_1570,In_2239,In_950);
nor U1571 (N_1571,In_2757,N_866);
and U1572 (N_1572,In_1836,In_328);
or U1573 (N_1573,In_83,In_1351);
xor U1574 (N_1574,N_1007,N_1351);
nand U1575 (N_1575,N_1379,N_121);
or U1576 (N_1576,N_344,N_660);
or U1577 (N_1577,N_351,N_75);
nand U1578 (N_1578,N_365,N_1160);
xnor U1579 (N_1579,In_1678,N_1245);
or U1580 (N_1580,N_1397,In_41);
xnor U1581 (N_1581,In_264,N_482);
or U1582 (N_1582,In_1419,In_216);
or U1583 (N_1583,In_2702,In_1939);
or U1584 (N_1584,N_1034,In_2986);
nor U1585 (N_1585,In_317,N_1334);
nand U1586 (N_1586,In_748,In_1118);
xor U1587 (N_1587,N_618,In_2308);
nand U1588 (N_1588,N_874,N_523);
or U1589 (N_1589,In_2944,N_254);
nor U1590 (N_1590,In_2511,N_55);
nand U1591 (N_1591,In_440,In_1176);
nor U1592 (N_1592,In_911,N_1380);
xor U1593 (N_1593,In_821,N_984);
xnor U1594 (N_1594,In_2105,N_1358);
nor U1595 (N_1595,N_1315,N_694);
or U1596 (N_1596,In_1057,N_388);
xnor U1597 (N_1597,N_1366,In_815);
and U1598 (N_1598,In_2012,N_92);
nor U1599 (N_1599,N_885,N_1040);
nor U1600 (N_1600,In_1789,N_1257);
or U1601 (N_1601,N_698,In_629);
nor U1602 (N_1602,In_1160,N_1343);
and U1603 (N_1603,N_684,N_1537);
and U1604 (N_1604,N_490,In_2787);
xor U1605 (N_1605,N_1426,In_1868);
nor U1606 (N_1606,In_1748,In_694);
xor U1607 (N_1607,N_849,N_1446);
nor U1608 (N_1608,In_68,In_493);
nand U1609 (N_1609,N_861,In_1560);
nand U1610 (N_1610,N_988,In_2550);
nor U1611 (N_1611,In_1954,N_1541);
or U1612 (N_1612,N_1348,N_832);
or U1613 (N_1613,In_2596,N_627);
xor U1614 (N_1614,In_177,In_597);
xnor U1615 (N_1615,In_2146,In_2372);
nand U1616 (N_1616,In_525,N_577);
and U1617 (N_1617,N_1248,N_346);
nor U1618 (N_1618,In_2138,N_241);
nand U1619 (N_1619,N_833,N_1432);
nand U1620 (N_1620,N_1573,In_1263);
or U1621 (N_1621,N_1355,In_2361);
and U1622 (N_1622,In_1529,N_179);
or U1623 (N_1623,N_979,In_1463);
and U1624 (N_1624,In_2339,N_943);
nor U1625 (N_1625,In_1784,N_1593);
and U1626 (N_1626,N_391,In_1138);
or U1627 (N_1627,N_925,In_2735);
and U1628 (N_1628,N_836,In_1232);
or U1629 (N_1629,N_705,In_1821);
xor U1630 (N_1630,N_1522,N_706);
and U1631 (N_1631,In_543,In_2766);
or U1632 (N_1632,N_1270,In_2639);
or U1633 (N_1633,N_1284,In_547);
nor U1634 (N_1634,N_405,N_1074);
or U1635 (N_1635,N_1529,In_1170);
or U1636 (N_1636,N_1301,In_1717);
and U1637 (N_1637,N_1508,N_1186);
xnor U1638 (N_1638,N_1215,N_863);
and U1639 (N_1639,N_293,N_913);
nor U1640 (N_1640,N_1472,In_1981);
xnor U1641 (N_1641,In_142,In_1557);
nor U1642 (N_1642,N_1264,In_2428);
and U1643 (N_1643,N_983,In_476);
and U1644 (N_1644,N_717,N_1179);
or U1645 (N_1645,N_1371,N_1383);
and U1646 (N_1646,N_266,N_1265);
nand U1647 (N_1647,In_2729,N_534);
xnor U1648 (N_1648,In_1758,In_2906);
xnor U1649 (N_1649,In_2029,N_1525);
or U1650 (N_1650,In_1662,N_635);
nand U1651 (N_1651,In_2913,In_1364);
nor U1652 (N_1652,N_384,N_95);
nor U1653 (N_1653,N_1010,In_204);
nor U1654 (N_1654,N_1374,N_1137);
nand U1655 (N_1655,N_120,In_1547);
xor U1656 (N_1656,N_1174,N_345);
and U1657 (N_1657,N_1051,In_2369);
nand U1658 (N_1658,In_795,In_373);
xnor U1659 (N_1659,In_1818,N_1428);
or U1660 (N_1660,N_941,In_212);
and U1661 (N_1661,In_1609,In_1705);
and U1662 (N_1662,N_746,N_1212);
nor U1663 (N_1663,In_503,N_1297);
xnor U1664 (N_1664,In_1350,In_1880);
nand U1665 (N_1665,In_119,N_1060);
nand U1666 (N_1666,N_775,N_1324);
xor U1667 (N_1667,In_1028,In_874);
nand U1668 (N_1668,N_670,N_1073);
or U1669 (N_1669,N_1524,N_131);
and U1670 (N_1670,In_533,In_1076);
nor U1671 (N_1671,In_2524,In_720);
and U1672 (N_1672,N_576,In_2204);
and U1673 (N_1673,In_2443,In_188);
xor U1674 (N_1674,N_1285,N_1455);
xor U1675 (N_1675,N_827,In_885);
and U1676 (N_1676,In_2823,In_938);
xor U1677 (N_1677,In_1958,N_1363);
nor U1678 (N_1678,N_647,In_2329);
nor U1679 (N_1679,In_2614,N_1347);
xor U1680 (N_1680,In_1287,N_1252);
or U1681 (N_1681,N_1312,N_1480);
nor U1682 (N_1682,In_889,N_1328);
or U1683 (N_1683,N_987,In_810);
xor U1684 (N_1684,N_549,In_1227);
and U1685 (N_1685,N_85,In_1157);
or U1686 (N_1686,In_870,In_2861);
nor U1687 (N_1687,N_1590,In_557);
nor U1688 (N_1688,In_161,In_902);
nand U1689 (N_1689,In_318,N_1405);
nor U1690 (N_1690,N_953,In_2592);
xnor U1691 (N_1691,In_1283,N_674);
xor U1692 (N_1692,N_1588,In_2049);
and U1693 (N_1693,In_1458,In_1521);
and U1694 (N_1694,In_2241,N_1516);
xor U1695 (N_1695,N_1484,In_2425);
and U1696 (N_1696,N_1589,N_930);
or U1697 (N_1697,N_246,N_938);
xor U1698 (N_1698,N_1511,N_646);
nor U1699 (N_1699,In_775,In_2500);
and U1700 (N_1700,In_973,N_524);
xnor U1701 (N_1701,N_31,N_829);
nand U1702 (N_1702,N_1554,N_1298);
or U1703 (N_1703,N_1372,In_652);
nand U1704 (N_1704,In_458,In_1383);
nor U1705 (N_1705,In_1347,N_1483);
xnor U1706 (N_1706,N_544,N_1392);
or U1707 (N_1707,In_692,N_1527);
or U1708 (N_1708,N_695,N_450);
and U1709 (N_1709,N_1457,N_1);
nand U1710 (N_1710,In_1327,N_1552);
nand U1711 (N_1711,In_2043,N_1434);
and U1712 (N_1712,In_454,In_1391);
xor U1713 (N_1713,N_87,In_208);
nand U1714 (N_1714,In_2610,In_1054);
nor U1715 (N_1715,N_12,In_1095);
nand U1716 (N_1716,In_797,In_1520);
nand U1717 (N_1717,In_1478,In_92);
nor U1718 (N_1718,N_1546,In_1318);
or U1719 (N_1719,N_1341,N_1436);
or U1720 (N_1720,N_1500,In_1303);
nor U1721 (N_1721,In_486,N_1171);
nor U1722 (N_1722,N_1420,In_878);
nor U1723 (N_1723,N_1377,N_868);
nand U1724 (N_1724,N_1408,In_1671);
xnor U1725 (N_1725,N_1125,N_1216);
or U1726 (N_1726,In_2177,In_1906);
nor U1727 (N_1727,N_1172,In_1837);
xor U1728 (N_1728,N_1557,N_1504);
nand U1729 (N_1729,In_2199,In_430);
xor U1730 (N_1730,N_1445,In_2710);
xor U1731 (N_1731,N_1501,In_2703);
or U1732 (N_1732,N_1112,In_899);
nor U1733 (N_1733,In_2475,N_1476);
nor U1734 (N_1734,In_257,In_2953);
nor U1735 (N_1735,N_1028,N_1214);
nand U1736 (N_1736,In_263,N_1280);
or U1737 (N_1737,In_1719,N_602);
xor U1738 (N_1738,N_1394,In_2256);
or U1739 (N_1739,In_2542,N_504);
xor U1740 (N_1740,N_759,N_1481);
nor U1741 (N_1741,In_2966,In_411);
and U1742 (N_1742,N_893,In_340);
and U1743 (N_1743,In_1523,N_782);
or U1744 (N_1744,N_1352,N_654);
or U1745 (N_1745,N_1531,N_1387);
xor U1746 (N_1746,N_20,In_1061);
nand U1747 (N_1747,In_2284,N_1502);
xnor U1748 (N_1748,In_1059,N_630);
and U1749 (N_1749,In_1042,N_831);
xnor U1750 (N_1750,In_2890,N_1162);
and U1751 (N_1751,N_1473,In_819);
or U1752 (N_1752,N_905,N_1350);
xor U1753 (N_1753,N_587,In_2359);
nand U1754 (N_1754,N_1056,N_1130);
nor U1755 (N_1755,N_1451,N_1042);
nor U1756 (N_1756,N_362,N_1542);
and U1757 (N_1757,N_1321,In_2168);
xnor U1758 (N_1758,In_1348,In_2505);
and U1759 (N_1759,N_462,N_1030);
xor U1760 (N_1760,In_1670,In_541);
nand U1761 (N_1761,N_1026,N_1449);
xnor U1762 (N_1762,N_1412,In_2282);
nand U1763 (N_1763,N_1307,In_2395);
and U1764 (N_1764,N_1505,N_1404);
nand U1765 (N_1765,N_1124,N_1104);
nand U1766 (N_1766,N_1169,In_968);
nand U1767 (N_1767,N_1274,In_1741);
nor U1768 (N_1768,In_2523,N_547);
xnor U1769 (N_1769,N_1575,N_1429);
or U1770 (N_1770,In_2877,N_214);
xor U1771 (N_1771,N_15,In_2089);
and U1772 (N_1772,N_1533,In_877);
nand U1773 (N_1773,In_986,N_1293);
nor U1774 (N_1774,N_1339,N_118);
nand U1775 (N_1775,N_1571,N_400);
nand U1776 (N_1776,In_2066,N_687);
or U1777 (N_1777,In_1274,N_1320);
xnor U1778 (N_1778,N_176,In_2069);
xor U1779 (N_1779,N_1282,In_401);
nor U1780 (N_1780,In_42,In_2327);
nand U1781 (N_1781,N_774,In_354);
nand U1782 (N_1782,In_1425,In_463);
or U1783 (N_1783,In_2170,In_841);
and U1784 (N_1784,In_1252,N_851);
nor U1785 (N_1785,In_1044,In_1110);
and U1786 (N_1786,N_143,N_1453);
nor U1787 (N_1787,N_397,N_477);
or U1788 (N_1788,N_927,N_168);
nor U1789 (N_1789,N_752,In_211);
or U1790 (N_1790,N_1465,In_1809);
xnor U1791 (N_1791,N_203,N_1273);
nor U1792 (N_1792,N_1288,In_1385);
or U1793 (N_1793,In_852,In_1862);
xnor U1794 (N_1794,In_1834,N_1583);
or U1795 (N_1795,N_1219,In_996);
xor U1796 (N_1796,N_1255,N_1033);
nand U1797 (N_1797,In_1039,N_1337);
xnor U1798 (N_1798,N_1568,In_1816);
and U1799 (N_1799,In_1994,N_1402);
nor U1800 (N_1800,N_838,In_1619);
and U1801 (N_1801,N_1602,N_1494);
xor U1802 (N_1802,In_347,In_1393);
nand U1803 (N_1803,In_2883,In_2251);
xnor U1804 (N_1804,In_2394,N_939);
nor U1805 (N_1805,In_1345,N_1548);
nor U1806 (N_1806,In_2818,N_1638);
nand U1807 (N_1807,N_1401,In_1432);
nand U1808 (N_1808,N_353,In_964);
nand U1809 (N_1809,N_1711,N_738);
and U1810 (N_1810,In_1113,N_952);
xor U1811 (N_1811,In_45,In_1386);
nor U1812 (N_1812,N_1678,N_1003);
and U1813 (N_1813,In_2865,N_395);
and U1814 (N_1814,In_955,In_2553);
or U1815 (N_1815,In_2496,In_1083);
and U1816 (N_1816,N_1784,N_1764);
and U1817 (N_1817,N_1462,In_1542);
nand U1818 (N_1818,In_2600,In_1293);
xor U1819 (N_1819,In_686,N_1213);
and U1820 (N_1820,In_867,N_1368);
nor U1821 (N_1821,N_1607,N_1564);
nor U1822 (N_1822,N_1549,N_302);
and U1823 (N_1823,In_2455,N_1742);
xnor U1824 (N_1824,In_2391,In_99);
or U1825 (N_1825,N_1706,N_1702);
and U1826 (N_1826,In_95,In_2432);
nand U1827 (N_1827,In_1856,N_1599);
xnor U1828 (N_1828,N_1772,In_561);
or U1829 (N_1829,N_703,In_2909);
or U1830 (N_1830,In_1257,In_1970);
or U1831 (N_1831,N_1353,In_1435);
nand U1832 (N_1832,In_2860,N_1425);
xnor U1833 (N_1833,In_736,N_883);
or U1834 (N_1834,In_1840,N_593);
or U1835 (N_1835,In_1932,N_946);
nor U1836 (N_1836,N_1096,N_1734);
xnor U1837 (N_1837,N_1606,N_1609);
nor U1838 (N_1838,In_1569,In_0);
nor U1839 (N_1839,N_1470,N_1400);
nor U1840 (N_1840,N_1153,In_1737);
or U1841 (N_1841,N_1622,N_1660);
xor U1842 (N_1842,N_1675,In_617);
nand U1843 (N_1843,N_1367,N_1047);
nor U1844 (N_1844,In_1850,N_1570);
or U1845 (N_1845,In_958,In_707);
or U1846 (N_1846,N_1536,In_461);
xnor U1847 (N_1847,In_1941,In_859);
nor U1848 (N_1848,In_2382,N_1331);
or U1849 (N_1849,In_2529,N_1038);
xor U1850 (N_1850,In_1275,In_2559);
or U1851 (N_1851,N_1302,In_627);
xor U1852 (N_1852,N_1621,N_1238);
nand U1853 (N_1853,N_1625,In_1599);
or U1854 (N_1854,In_2586,In_1004);
or U1855 (N_1855,N_323,In_2618);
nor U1856 (N_1856,In_26,In_215);
or U1857 (N_1857,In_1031,N_243);
or U1858 (N_1858,In_2481,N_1329);
nand U1859 (N_1859,In_574,N_1519);
and U1860 (N_1860,In_2291,N_1095);
nor U1861 (N_1861,In_2590,N_842);
and U1862 (N_1862,In_2024,N_1559);
xnor U1863 (N_1863,N_1659,In_266);
xnor U1864 (N_1864,In_554,N_1478);
xor U1865 (N_1865,N_1142,In_387);
or U1866 (N_1866,N_1540,N_792);
nand U1867 (N_1867,N_949,N_1725);
nor U1868 (N_1868,N_881,N_1662);
nor U1869 (N_1869,In_711,N_1521);
or U1870 (N_1870,N_1650,N_1770);
or U1871 (N_1871,In_1646,N_1720);
and U1872 (N_1872,N_445,N_1152);
nor U1873 (N_1873,N_1474,N_553);
xor U1874 (N_1874,N_1618,In_1246);
nor U1875 (N_1875,N_1057,In_2911);
xnor U1876 (N_1876,N_797,N_1459);
and U1877 (N_1877,N_465,N_303);
xnor U1878 (N_1878,In_976,In_576);
xnor U1879 (N_1879,In_85,In_2330);
xor U1880 (N_1880,In_995,N_783);
xor U1881 (N_1881,In_1687,N_1229);
xor U1882 (N_1882,N_1580,In_2479);
xnor U1883 (N_1883,N_1701,In_289);
nand U1884 (N_1884,N_1308,N_1673);
nand U1885 (N_1885,In_1617,N_1723);
and U1886 (N_1886,N_1417,N_1416);
nor U1887 (N_1887,In_2267,In_81);
nor U1888 (N_1888,In_2519,In_957);
xor U1889 (N_1889,N_1563,N_834);
nand U1890 (N_1890,N_1515,In_2044);
xor U1891 (N_1891,N_1492,N_1278);
nand U1892 (N_1892,N_1684,N_1319);
nor U1893 (N_1893,N_151,In_232);
xor U1894 (N_1894,N_1765,N_372);
nor U1895 (N_1895,N_1247,N_1558);
and U1896 (N_1896,N_857,In_1607);
or U1897 (N_1897,N_1705,N_882);
nor U1898 (N_1898,In_1080,N_1672);
or U1899 (N_1899,N_521,N_715);
and U1900 (N_1900,N_708,N_60);
xnor U1901 (N_1901,N_1464,In_338);
xnor U1902 (N_1902,In_1240,N_483);
xnor U1903 (N_1903,In_1372,In_2217);
or U1904 (N_1904,N_1458,In_2332);
xor U1905 (N_1905,In_1734,N_807);
or U1906 (N_1906,N_1235,N_1509);
and U1907 (N_1907,N_1290,In_2656);
nand U1908 (N_1908,N_1628,N_1463);
and U1909 (N_1909,In_1661,N_1619);
nor U1910 (N_1910,In_2311,N_433);
xnor U1911 (N_1911,N_865,N_343);
xor U1912 (N_1912,N_876,In_101);
and U1913 (N_1913,N_700,In_1632);
nand U1914 (N_1914,In_922,N_1745);
nor U1915 (N_1915,In_1332,N_890);
or U1916 (N_1916,N_1689,N_1682);
nand U1917 (N_1917,N_1017,N_222);
xor U1918 (N_1918,N_922,N_1761);
nor U1919 (N_1919,N_1454,N_1732);
xor U1920 (N_1920,In_108,N_825);
or U1921 (N_1921,N_1012,In_2867);
nor U1922 (N_1922,N_156,N_487);
xor U1923 (N_1923,N_1712,In_2225);
and U1924 (N_1924,N_1587,In_1333);
or U1925 (N_1925,N_1595,N_1221);
xor U1926 (N_1926,N_1389,In_6);
and U1927 (N_1927,N_1657,N_1714);
or U1928 (N_1928,N_411,N_1578);
nand U1929 (N_1929,N_555,N_1626);
xnor U1930 (N_1930,N_1168,N_52);
nor U1931 (N_1931,In_27,N_1107);
nand U1932 (N_1932,In_587,In_431);
or U1933 (N_1933,N_742,In_246);
and U1934 (N_1934,In_729,N_607);
nand U1935 (N_1935,N_1724,N_1582);
nor U1936 (N_1936,N_1735,N_750);
nand U1937 (N_1937,N_1574,N_1674);
nor U1938 (N_1938,N_1738,N_1579);
nor U1939 (N_1939,N_608,In_1688);
and U1940 (N_1940,In_1976,N_506);
nor U1941 (N_1941,In_1069,N_1147);
xor U1942 (N_1942,N_1192,N_1733);
or U1943 (N_1943,N_164,N_1370);
xor U1944 (N_1944,N_1210,In_1624);
and U1945 (N_1945,N_989,N_1671);
or U1946 (N_1946,N_1677,N_1526);
and U1947 (N_1947,In_2091,N_1780);
nor U1948 (N_1948,N_1757,N_599);
nand U1949 (N_1949,In_1716,N_1693);
xnor U1950 (N_1950,N_1781,N_1614);
or U1951 (N_1951,N_820,N_878);
nor U1952 (N_1952,N_557,N_1612);
nor U1953 (N_1953,N_1259,N_1409);
nand U1954 (N_1954,N_718,N_909);
nand U1955 (N_1955,N_707,In_2928);
and U1956 (N_1956,In_1649,N_1700);
xnor U1957 (N_1957,In_129,N_1667);
nor U1958 (N_1958,N_854,N_1692);
xnor U1959 (N_1959,In_1313,N_566);
nor U1960 (N_1960,N_439,N_1295);
or U1961 (N_1961,N_1127,In_2765);
and U1962 (N_1962,In_110,N_583);
and U1963 (N_1963,N_1369,In_2400);
nor U1964 (N_1964,N_872,In_2490);
or U1965 (N_1965,In_1026,N_1386);
or U1966 (N_1966,N_244,N_455);
nor U1967 (N_1967,In_2978,In_106);
or U1968 (N_1968,In_2269,In_1702);
xnor U1969 (N_1969,In_800,N_1795);
xnor U1970 (N_1970,N_497,N_788);
and U1971 (N_1971,N_1256,N_976);
nor U1972 (N_1972,In_2346,N_1410);
or U1973 (N_1973,N_1769,N_870);
or U1974 (N_1974,In_1653,N_1448);
xnor U1975 (N_1975,N_1680,In_2111);
and U1976 (N_1976,N_204,In_1116);
nor U1977 (N_1977,N_525,In_659);
and U1978 (N_1978,N_540,N_1161);
or U1979 (N_1979,N_1204,N_966);
nor U1980 (N_1980,In_2776,In_2632);
xor U1981 (N_1981,N_1039,N_1080);
xor U1982 (N_1982,N_1332,N_1283);
nor U1983 (N_1983,In_649,N_794);
nand U1984 (N_1984,N_110,In_2994);
nand U1985 (N_1985,N_307,In_696);
and U1986 (N_1986,N_747,N_1517);
xnor U1987 (N_1987,In_1797,In_2354);
nand U1988 (N_1988,N_1777,In_912);
nand U1989 (N_1989,N_1384,N_844);
or U1990 (N_1990,In_1946,In_1107);
xnor U1991 (N_1991,N_206,N_373);
and U1992 (N_1992,N_1035,In_1411);
or U1993 (N_1993,N_392,N_1503);
and U1994 (N_1994,N_1414,N_1276);
nand U1995 (N_1995,N_239,N_858);
nor U1996 (N_1996,N_982,N_1748);
nor U1997 (N_1997,N_1513,In_1893);
or U1998 (N_1998,N_142,N_529);
or U1999 (N_1999,N_478,In_23);
xor U2000 (N_2000,In_647,In_1942);
and U2001 (N_2001,In_1833,In_1559);
or U2002 (N_2002,In_2377,In_1456);
nor U2003 (N_2003,N_1666,N_1982);
and U2004 (N_2004,N_1937,N_1690);
and U2005 (N_2005,N_1953,N_1150);
nor U2006 (N_2006,In_1532,N_1987);
or U2007 (N_2007,In_1641,N_1683);
nor U2008 (N_2008,N_1317,N_28);
nor U2009 (N_2009,N_1923,N_102);
nand U2010 (N_2010,N_1903,In_926);
xor U2011 (N_2011,N_1899,In_1150);
or U2012 (N_2012,N_1305,N_1685);
nor U2013 (N_2013,N_1670,N_1886);
xor U2014 (N_2014,N_1403,N_1016);
nor U2015 (N_2015,N_818,N_167);
nand U2016 (N_2016,N_1747,N_1876);
nand U2017 (N_2017,In_1866,In_838);
nor U2018 (N_2018,N_1827,N_1783);
xor U2019 (N_2019,N_1822,N_1794);
and U2020 (N_2020,In_1882,In_569);
and U2021 (N_2021,N_1950,N_1835);
nor U2022 (N_2022,N_208,N_335);
xor U2023 (N_2023,N_1045,In_2634);
nand U2024 (N_2024,In_1518,N_1156);
nor U2025 (N_2025,N_1857,In_2738);
and U2026 (N_2026,N_1195,N_1900);
and U2027 (N_2027,In_2441,N_321);
or U2028 (N_2028,N_1957,N_907);
nand U2029 (N_2029,N_1837,N_619);
nor U2030 (N_2030,N_1362,N_682);
or U2031 (N_2031,N_629,N_1013);
and U2032 (N_2032,In_362,N_474);
nor U2033 (N_2033,N_1357,N_1811);
nand U2034 (N_2034,In_261,N_1629);
nor U2035 (N_2035,In_2689,N_1036);
nor U2036 (N_2036,N_1785,N_1647);
nand U2037 (N_2037,N_960,N_1261);
and U2038 (N_2038,N_1489,N_1361);
nor U2039 (N_2039,N_1037,N_1158);
nor U2040 (N_2040,In_1360,In_397);
nor U2041 (N_2041,N_1945,N_122);
nor U2042 (N_2042,N_961,N_1246);
xor U2043 (N_2043,N_1995,N_1727);
or U2044 (N_2044,N_1450,N_1911);
nand U2045 (N_2045,In_1978,N_512);
xor U2046 (N_2046,In_73,N_1704);
nor U2047 (N_2047,N_377,N_1709);
xor U2048 (N_2048,In_2963,N_1933);
nand U2049 (N_2049,In_1144,N_1289);
or U2050 (N_2050,N_1861,N_1750);
and U2051 (N_2051,In_2184,N_1165);
nand U2052 (N_2052,N_1956,N_1032);
or U2053 (N_2053,N_1433,N_895);
and U2054 (N_2054,N_1209,N_579);
nand U2055 (N_2055,In_689,In_2289);
and U2056 (N_2056,N_1817,N_1108);
nand U2057 (N_2057,N_1912,N_1843);
nor U2058 (N_2058,N_1376,N_1232);
nand U2059 (N_2059,N_1439,N_1065);
or U2060 (N_2060,In_75,In_863);
and U2061 (N_2061,N_1002,N_1695);
xor U2062 (N_2062,N_406,N_1335);
xor U2063 (N_2063,N_1115,In_2134);
xor U2064 (N_2064,N_1506,N_962);
or U2065 (N_2065,N_1479,N_1006);
nor U2066 (N_2066,In_1132,In_2769);
or U2067 (N_2067,N_1960,N_451);
or U2068 (N_2068,N_508,In_1992);
xor U2069 (N_2069,N_1773,N_1499);
xnor U2070 (N_2070,N_1896,N_1807);
or U2071 (N_2071,N_663,N_1177);
nand U2072 (N_2072,In_1331,N_856);
nand U2073 (N_2073,N_912,N_1828);
and U2074 (N_2074,In_1068,In_2588);
nor U2075 (N_2075,N_572,N_340);
or U2076 (N_2076,N_42,N_1431);
or U2077 (N_2077,N_624,N_1863);
nand U2078 (N_2078,N_1983,N_1721);
and U2079 (N_2079,N_1959,In_1601);
or U2080 (N_2080,N_1430,N_1222);
and U2081 (N_2081,N_1642,In_1762);
xor U2082 (N_2082,In_2910,N_926);
or U2083 (N_2083,In_1344,N_1810);
or U2084 (N_2084,N_1867,N_1419);
xnor U2085 (N_2085,In_1121,N_1838);
or U2086 (N_2086,In_2898,In_2228);
nor U2087 (N_2087,In_1676,N_1963);
or U2088 (N_2088,In_1401,N_1885);
nand U2089 (N_2089,In_1714,N_1914);
and U2090 (N_2090,In_858,N_1523);
or U2091 (N_2091,N_1787,N_1832);
nor U2092 (N_2092,In_2675,In_2520);
or U2093 (N_2093,In_2360,N_1884);
nand U2094 (N_2094,In_2683,In_566);
xnor U2095 (N_2095,In_1325,In_564);
xor U2096 (N_2096,N_1873,N_1927);
or U2097 (N_2097,N_1825,In_320);
nor U2098 (N_2098,N_855,In_1495);
xnor U2099 (N_2099,N_1964,N_1545);
or U2100 (N_2100,N_1613,N_1935);
or U2101 (N_2101,N_1155,N_1688);
nor U2102 (N_2102,N_1925,In_172);
or U2103 (N_2103,N_1736,N_1364);
nand U2104 (N_2104,N_1907,In_342);
or U2105 (N_2105,N_1475,N_1974);
nor U2106 (N_2106,In_1041,In_275);
xor U2107 (N_2107,In_2539,N_809);
nor U2108 (N_2108,N_1815,N_914);
nand U2109 (N_2109,N_1924,N_1880);
nor U2110 (N_2110,In_2674,N_1743);
and U2111 (N_2111,N_1965,N_1497);
and U2112 (N_2112,N_1296,N_1901);
nand U2113 (N_2113,N_1968,In_2997);
nand U2114 (N_2114,N_917,N_1346);
nand U2115 (N_2115,N_1632,N_1992);
nand U2116 (N_2116,In_1728,N_410);
or U2117 (N_2117,In_545,N_1084);
xor U2118 (N_2118,N_1145,In_2992);
and U2119 (N_2119,N_625,In_2074);
or U2120 (N_2120,N_1889,N_1648);
or U2121 (N_2121,In_438,N_1093);
xor U2122 (N_2122,In_1749,In_1575);
nor U2123 (N_2123,N_1759,N_1739);
xor U2124 (N_2124,N_1636,N_1971);
and U2125 (N_2125,N_802,N_1443);
nand U2126 (N_2126,N_1020,In_2567);
or U2127 (N_2127,N_1868,In_292);
xnor U2128 (N_2128,N_1771,In_2120);
nand U2129 (N_2129,N_1751,N_997);
or U2130 (N_2130,N_668,N_1616);
and U2131 (N_2131,N_446,In_2383);
xor U2132 (N_2132,N_1543,N_1600);
and U2133 (N_2133,N_1468,N_1803);
or U2134 (N_2134,N_1722,N_743);
nand U2135 (N_2135,N_1314,N_1586);
and U2136 (N_2136,In_981,N_1833);
nor U2137 (N_2137,In_2671,In_2402);
xor U2138 (N_2138,N_304,N_1653);
xor U2139 (N_2139,N_1801,N_1973);
nor U2140 (N_2140,N_1800,N_336);
nand U2141 (N_2141,N_1908,N_396);
xnor U2142 (N_2142,N_1947,In_2631);
and U2143 (N_2143,In_682,N_1493);
xor U2144 (N_2144,N_1697,N_1962);
or U2145 (N_2145,N_801,In_348);
or U2146 (N_2146,In_599,N_1486);
and U2147 (N_2147,N_1550,N_1792);
xnor U2148 (N_2148,N_1881,N_767);
nand U2149 (N_2149,N_1191,N_1934);
nor U2150 (N_2150,N_262,N_1994);
or U2151 (N_2151,In_2122,N_1719);
xnor U2152 (N_2152,N_1102,N_768);
or U2153 (N_2153,N_1651,N_1623);
nor U2154 (N_2154,In_668,In_2378);
or U2155 (N_2155,N_1708,N_1768);
or U2156 (N_2156,N_649,N_1001);
xor U2157 (N_2157,N_1729,In_147);
nand U2158 (N_2158,N_1904,N_1840);
nor U2159 (N_2159,In_656,N_1116);
and U2160 (N_2160,N_1422,N_1310);
xor U2161 (N_2161,In_2246,N_1681);
nand U2162 (N_2162,In_1200,N_1620);
and U2163 (N_2163,N_1311,In_1473);
or U2164 (N_2164,In_1810,N_1922);
and U2165 (N_2165,N_248,N_1991);
xor U2166 (N_2166,N_1611,N_1617);
or U2167 (N_2167,N_144,N_1665);
xor U2168 (N_2168,N_1566,N_1944);
nand U2169 (N_2169,N_1788,N_191);
or U2170 (N_2170,N_1936,N_1854);
or U2171 (N_2171,N_1749,In_2799);
nand U2172 (N_2172,N_1654,N_1831);
and U2173 (N_2173,In_1474,N_1902);
nand U2174 (N_2174,N_1180,In_1550);
xnor U2175 (N_2175,N_219,N_1746);
and U2176 (N_2176,N_1005,In_396);
xnor U2177 (N_2177,N_65,N_1244);
or U2178 (N_2178,N_1603,In_58);
and U2179 (N_2179,In_967,N_1948);
xnor U2180 (N_2180,In_2355,N_264);
xor U2181 (N_2181,In_2940,N_1591);
or U2182 (N_2182,N_1940,N_1052);
nor U2183 (N_2183,In_316,N_1989);
and U2184 (N_2184,N_1853,N_1892);
nand U2185 (N_2185,N_1604,N_1883);
xnor U2186 (N_2186,N_1668,N_1421);
and U2187 (N_2187,N_1477,N_963);
and U2188 (N_2188,N_1758,N_1029);
nor U2189 (N_2189,N_628,N_1044);
and U2190 (N_2190,N_1447,N_1652);
nand U2191 (N_2191,N_1637,N_1645);
nor U2192 (N_2192,In_2578,In_2746);
nand U2193 (N_2193,N_1133,In_423);
nand U2194 (N_2194,In_2347,In_2888);
nand U2195 (N_2195,In_1281,N_1299);
or U2196 (N_2196,In_2802,N_1818);
xor U2197 (N_2197,In_138,N_1894);
nand U2198 (N_2198,N_702,N_1805);
and U2199 (N_2199,In_1023,N_1814);
nand U2200 (N_2200,N_2107,N_1841);
or U2201 (N_2201,N_1507,N_1388);
or U2202 (N_2202,N_2137,N_1560);
and U2203 (N_2203,N_1895,N_1495);
and U2204 (N_2204,In_1315,N_2086);
and U2205 (N_2205,N_1997,N_2051);
nor U2206 (N_2206,N_1970,N_2191);
or U2207 (N_2207,N_2007,N_2064);
or U2208 (N_2208,In_1201,In_2856);
or U2209 (N_2209,N_2176,In_2174);
nor U2210 (N_2210,In_2960,N_2126);
xnor U2211 (N_2211,N_2183,N_1528);
nor U2212 (N_2212,N_2106,In_751);
nand U2213 (N_2213,In_2016,In_93);
and U2214 (N_2214,N_1148,N_1236);
or U2215 (N_2215,N_2123,In_965);
nand U2216 (N_2216,N_399,N_2174);
and U2217 (N_2217,N_1691,In_1278);
xnor U2218 (N_2218,In_179,N_2150);
nand U2219 (N_2219,N_1471,N_2092);
nor U2220 (N_2220,N_1159,N_1919);
and U2221 (N_2221,In_2544,N_848);
and U2222 (N_2222,N_2160,N_2057);
or U2223 (N_2223,In_287,In_770);
or U2224 (N_2224,N_2154,In_799);
or U2225 (N_2225,In_2057,N_1891);
xor U2226 (N_2226,N_1272,N_1487);
and U2227 (N_2227,In_2234,N_1535);
or U2228 (N_2228,N_1829,N_2021);
nor U2229 (N_2229,N_2136,N_1534);
xor U2230 (N_2230,N_1225,N_1812);
nand U2231 (N_2231,N_2010,N_2149);
and U2232 (N_2232,In_2522,N_2077);
nand U2233 (N_2233,N_2144,N_1461);
nor U2234 (N_2234,N_1893,In_2157);
xor U2235 (N_2235,N_1663,N_422);
nand U2236 (N_2236,N_1086,N_1981);
nor U2237 (N_2237,N_2190,N_2169);
nor U2238 (N_2238,N_349,N_1848);
xor U2239 (N_2239,In_2466,N_1318);
nor U2240 (N_2240,N_1698,N_2193);
or U2241 (N_2241,N_2002,In_2836);
nand U2242 (N_2242,N_1796,In_306);
or U2243 (N_2243,N_2097,N_1808);
or U2244 (N_2244,N_1565,N_1577);
or U2245 (N_2245,N_2058,N_1091);
nor U2246 (N_2246,N_1556,In_2620);
and U2247 (N_2247,N_819,N_1496);
or U2248 (N_2248,In_603,In_1739);
nor U2249 (N_2249,N_1067,N_955);
or U2250 (N_2250,N_1279,N_1999);
xor U2251 (N_2251,N_2196,N_1469);
nor U2252 (N_2252,N_2096,In_2281);
and U2253 (N_2253,In_367,N_2050);
nand U2254 (N_2254,N_2017,N_1791);
nand U2255 (N_2255,N_1726,N_1988);
and U2256 (N_2256,N_1605,N_1898);
xor U2257 (N_2257,N_1954,N_2068);
nor U2258 (N_2258,N_1866,In_2743);
xor U2259 (N_2259,N_2109,N_519);
nand U2260 (N_2260,N_1520,N_226);
nor U2261 (N_2261,In_2921,N_2094);
nor U2262 (N_2262,In_727,N_1860);
nor U2263 (N_2263,N_2161,N_1939);
xor U2264 (N_2264,In_779,N_1943);
xor U2265 (N_2265,N_1227,N_1782);
nand U2266 (N_2266,N_319,N_906);
xnor U2267 (N_2267,N_1752,N_1058);
and U2268 (N_2268,N_2105,N_290);
nand U2269 (N_2269,N_291,In_141);
nor U2270 (N_2270,N_973,N_2053);
nand U2271 (N_2271,N_1393,N_357);
nand U2272 (N_2272,N_1512,N_1839);
nand U2273 (N_2273,N_1661,N_1237);
or U2274 (N_2274,N_1041,N_2192);
xor U2275 (N_2275,In_1692,N_2155);
nor U2276 (N_2276,N_1268,N_1643);
nand U2277 (N_2277,N_1427,N_1594);
xor U2278 (N_2278,In_753,N_1395);
and U2279 (N_2279,N_2061,N_526);
nor U2280 (N_2280,N_62,In_979);
nand U2281 (N_2281,N_2110,N_2166);
xor U2282 (N_2282,In_2676,N_1717);
xnor U2283 (N_2283,In_2121,N_1767);
or U2284 (N_2284,N_1713,In_2027);
xnor U2285 (N_2285,N_1703,In_937);
nand U2286 (N_2286,N_2066,N_1952);
or U2287 (N_2287,N_1597,N_1113);
or U2288 (N_2288,N_920,N_1715);
and U2289 (N_2289,N_2114,In_448);
and U2290 (N_2290,N_2025,N_485);
xor U2291 (N_2291,N_134,N_1882);
nand U2292 (N_2292,N_954,N_904);
nand U2293 (N_2293,N_552,N_1646);
or U2294 (N_2294,N_1864,N_929);
xor U2295 (N_2295,In_2892,N_366);
xnor U2296 (N_2296,N_1031,In_2869);
or U2297 (N_2297,N_2165,N_1027);
or U2298 (N_2298,N_2128,N_896);
and U2299 (N_2299,N_2152,N_2005);
and U2300 (N_2300,N_447,N_471);
nor U2301 (N_2301,N_2060,N_1826);
xor U2302 (N_2302,N_1967,N_1631);
and U2303 (N_2303,N_2001,N_1398);
nor U2304 (N_2304,N_2019,N_1920);
nand U2305 (N_2305,In_1380,N_1581);
nand U2306 (N_2306,N_1932,In_451);
nor U2307 (N_2307,N_2036,In_2839);
and U2308 (N_2308,N_2013,N_1862);
and U2309 (N_2309,N_847,N_1852);
xor U2310 (N_2310,In_2739,N_1262);
nand U2311 (N_2311,N_2093,N_2198);
nor U2312 (N_2312,N_1555,N_1890);
nor U2313 (N_2313,N_1993,In_1494);
xnor U2314 (N_2314,N_2041,N_2099);
or U2315 (N_2315,N_975,N_1686);
or U2316 (N_2316,N_2142,N_1887);
nor U2317 (N_2317,N_2091,N_1220);
or U2318 (N_2318,N_2177,N_2186);
nand U2319 (N_2319,In_2627,N_1879);
and U2320 (N_2320,N_916,N_2029);
and U2321 (N_2321,N_1553,N_978);
nor U2322 (N_2322,In_2764,N_1941);
and U2323 (N_2323,N_1598,N_1202);
nor U2324 (N_2324,N_1406,N_1187);
or U2325 (N_2325,N_2129,N_1921);
xor U2326 (N_2326,N_1802,N_1949);
nor U2327 (N_2327,In_1109,N_2087);
and U2328 (N_2328,N_637,N_1173);
or U2329 (N_2329,N_603,N_645);
xnor U2330 (N_2330,N_1601,In_1210);
nand U2331 (N_2331,N_1407,In_2515);
xor U2332 (N_2332,N_489,N_1572);
and U2333 (N_2333,N_1123,N_2184);
xor U2334 (N_2334,N_1655,N_2069);
nand U2335 (N_2335,N_2127,N_1799);
xnor U2336 (N_2336,N_1567,In_46);
or U2337 (N_2337,In_1056,N_1488);
or U2338 (N_2338,N_1467,N_1778);
and U2339 (N_2339,N_2103,N_1004);
nand U2340 (N_2340,N_2048,N_1189);
and U2341 (N_2341,N_1888,N_2164);
or U2342 (N_2342,N_2181,N_620);
nand U2343 (N_2343,N_1744,N_1326);
xnor U2344 (N_2344,In_1585,N_2101);
xor U2345 (N_2345,N_2117,N_2065);
nor U2346 (N_2346,N_1624,N_1518);
nor U2347 (N_2347,N_2052,N_1585);
xor U2348 (N_2348,N_1930,N_1596);
or U2349 (N_2349,N_2056,N_1918);
xor U2350 (N_2350,N_1530,N_1009);
or U2351 (N_2351,N_2098,In_183);
nand U2352 (N_2352,N_1849,N_1287);
xor U2353 (N_2353,N_1865,N_2046);
nand U2354 (N_2354,N_2024,In_2273);
nor U2355 (N_2355,N_1875,N_1608);
nor U2356 (N_2356,N_1766,N_1390);
and U2357 (N_2357,N_417,N_2082);
nor U2358 (N_2358,N_1961,N_1415);
or U2359 (N_2359,N_1977,N_1905);
nor U2360 (N_2360,N_84,N_1203);
and U2361 (N_2361,N_1615,N_273);
nor U2362 (N_2362,N_2032,N_2023);
and U2363 (N_2363,In_1863,In_1743);
and U2364 (N_2364,N_1798,N_1756);
and U2365 (N_2365,N_2195,N_1699);
or U2366 (N_2366,N_1878,In_1406);
or U2367 (N_2367,N_2074,In_48);
xor U2368 (N_2368,In_1766,N_1855);
and U2369 (N_2369,N_1975,N_1561);
or U2370 (N_2370,N_1951,N_1022);
xor U2371 (N_2371,N_1929,N_942);
xor U2372 (N_2372,N_1966,N_1490);
nand U2373 (N_2373,N_2100,N_908);
xor U2374 (N_2374,N_1423,N_2009);
and U2375 (N_2375,N_867,N_1544);
nand U2376 (N_2376,N_2042,N_1066);
nand U2377 (N_2377,N_341,N_594);
or U2378 (N_2378,N_1634,In_1507);
or U2379 (N_2379,N_2015,N_1185);
nand U2380 (N_2380,N_2075,N_2139);
or U2381 (N_2381,N_232,N_2134);
or U2382 (N_2382,N_992,N_1980);
and U2383 (N_2383,N_1452,N_1972);
nor U2384 (N_2384,N_1669,N_633);
and U2385 (N_2385,N_2153,N_330);
nand U2386 (N_2386,N_2076,N_1538);
nor U2387 (N_2387,In_312,N_1872);
xnor U2388 (N_2388,N_1592,N_753);
nor U2389 (N_2389,N_1437,In_2453);
xor U2390 (N_2390,N_1928,N_2033);
nand U2391 (N_2391,In_1870,N_1793);
and U2392 (N_2392,In_38,N_688);
xnor U2393 (N_2393,N_1610,In_1146);
and U2394 (N_2394,N_1819,N_2004);
xnor U2395 (N_2395,N_897,N_1779);
nor U2396 (N_2396,In_1130,N_1438);
nand U2397 (N_2397,N_859,N_428);
and U2398 (N_2398,N_2138,N_1774);
nand U2399 (N_2399,In_2952,N_2147);
nand U2400 (N_2400,N_1737,N_2280);
nand U2401 (N_2401,N_1349,N_2267);
nand U2402 (N_2402,N_590,In_1504);
and U2403 (N_2403,N_2067,N_1365);
nor U2404 (N_2404,N_1375,N_2210);
xor U2405 (N_2405,N_1869,N_1456);
or U2406 (N_2406,N_13,N_1906);
or U2407 (N_2407,N_2335,N_72);
and U2408 (N_2408,N_1760,N_1208);
and U2409 (N_2409,N_835,N_1249);
xnor U2410 (N_2410,N_2390,N_2336);
nand U2411 (N_2411,N_2258,N_1836);
and U2412 (N_2412,N_1969,N_1218);
xor U2413 (N_2413,In_2508,N_2008);
nand U2414 (N_2414,N_2080,N_2263);
nor U2415 (N_2415,N_2292,N_799);
xor U2416 (N_2416,N_2018,N_2132);
and U2417 (N_2417,In_551,N_1441);
or U2418 (N_2418,In_755,In_921);
and U2419 (N_2419,N_1182,N_1562);
or U2420 (N_2420,In_1623,N_2217);
and U2421 (N_2421,N_2320,N_2313);
nor U2422 (N_2422,N_1753,N_667);
nand U2423 (N_2423,N_1442,N_1391);
or U2424 (N_2424,N_2385,In_2385);
nand U2425 (N_2425,N_2016,N_2115);
and U2426 (N_2426,N_2391,N_1644);
nor U2427 (N_2427,N_2311,N_2167);
nand U2428 (N_2428,In_1052,In_2215);
and U2429 (N_2429,N_2000,N_1938);
xnor U2430 (N_2430,N_2379,N_1931);
nand U2431 (N_2431,In_1539,In_1341);
or U2432 (N_2432,In_598,N_2244);
xor U2433 (N_2433,In_2464,N_2316);
nor U2434 (N_2434,N_2281,N_1440);
nor U2435 (N_2435,N_1411,N_2072);
and U2436 (N_2436,In_450,N_709);
or U2437 (N_2437,N_1070,In_669);
and U2438 (N_2438,N_2189,N_683);
or U2439 (N_2439,N_2314,N_1740);
or U2440 (N_2440,N_64,N_202);
or U2441 (N_2441,N_2156,N_541);
or U2442 (N_2442,N_2070,N_1184);
xor U2443 (N_2443,N_2141,N_2230);
nand U2444 (N_2444,N_2211,In_1255);
nor U2445 (N_2445,In_2629,N_1664);
and U2446 (N_2446,N_2326,N_2324);
nand U2447 (N_2447,N_1271,N_2118);
nand U2448 (N_2448,N_1754,N_1728);
and U2449 (N_2449,N_2371,N_2011);
nor U2450 (N_2450,N_2393,N_2089);
nand U2451 (N_2451,N_1763,N_2112);
xor U2452 (N_2452,N_1913,N_1910);
nand U2453 (N_2453,N_2084,N_1584);
and U2454 (N_2454,N_2397,In_1475);
nand U2455 (N_2455,N_2333,N_1081);
nor U2456 (N_2456,N_1460,In_931);
or U2457 (N_2457,N_2245,N_69);
nand U2458 (N_2458,N_2073,N_1676);
or U2459 (N_2459,N_2376,N_1915);
xnor U2460 (N_2460,N_2220,N_2090);
nand U2461 (N_2461,N_318,N_1206);
nor U2462 (N_2462,N_2378,N_2315);
and U2463 (N_2463,N_1117,In_2741);
nand U2464 (N_2464,N_1120,In_1796);
or U2465 (N_2465,In_674,In_1177);
nor U2466 (N_2466,N_2305,N_2205);
nand U2467 (N_2467,N_1696,N_2380);
nand U2468 (N_2468,N_2124,N_1859);
and U2469 (N_2469,N_2387,N_2221);
or U2470 (N_2470,In_1267,N_837);
or U2471 (N_2471,N_1687,N_2043);
and U2472 (N_2472,N_958,N_672);
and U2473 (N_2473,In_2863,N_2374);
and U2474 (N_2474,N_2182,N_2256);
xor U2475 (N_2475,N_2257,N_2291);
xnor U2476 (N_2476,N_1958,N_2085);
and U2477 (N_2477,N_2355,N_598);
xor U2478 (N_2478,N_1850,N_2269);
nor U2479 (N_2479,N_1823,N_1359);
or U2480 (N_2480,N_2347,N_2047);
or U2481 (N_2481,N_2297,N_816);
or U2482 (N_2482,N_2243,N_1170);
xor U2483 (N_2483,N_1824,N_1718);
nand U2484 (N_2484,N_1741,N_2253);
and U2485 (N_2485,N_616,N_1323);
nor U2486 (N_2486,In_856,N_2308);
or U2487 (N_2487,N_864,N_2236);
or U2488 (N_2488,In_80,N_2022);
and U2489 (N_2489,N_2224,N_2353);
xnor U2490 (N_2490,N_2396,N_1979);
nand U2491 (N_2491,N_2163,N_2342);
nand U2492 (N_2492,N_2222,N_2235);
nor U2493 (N_2493,N_2383,N_1955);
and U2494 (N_2494,N_691,N_2354);
or U2495 (N_2495,N_1539,N_811);
nor U2496 (N_2496,N_921,In_243);
and U2497 (N_2497,N_1630,N_2202);
or U2498 (N_2498,N_2040,N_1166);
and U2499 (N_2499,N_2290,N_518);
and U2500 (N_2500,N_2071,N_2225);
xnor U2501 (N_2501,N_1978,N_1196);
or U2502 (N_2502,N_2330,N_2063);
nor U2503 (N_2503,N_2295,N_1806);
xnor U2504 (N_2504,N_2304,N_2208);
xor U2505 (N_2505,N_879,N_2337);
nor U2506 (N_2506,N_2020,N_2254);
and U2507 (N_2507,N_463,N_1277);
and U2508 (N_2508,N_2125,N_2301);
nor U2509 (N_2509,In_747,N_1984);
nand U2510 (N_2510,In_443,N_1996);
and U2511 (N_2511,N_2259,N_884);
xor U2512 (N_2512,N_1141,N_2345);
or U2513 (N_2513,N_2356,N_1656);
xor U2514 (N_2514,N_2157,N_2034);
nand U2515 (N_2515,N_2204,N_1199);
and U2516 (N_2516,N_681,N_2327);
or U2517 (N_2517,N_2031,N_1858);
xor U2518 (N_2518,N_2095,N_1786);
and U2519 (N_2519,N_2054,N_2006);
nand U2520 (N_2520,In_1919,In_37);
nand U2521 (N_2521,N_180,In_1582);
nor U2522 (N_2522,N_2045,N_2216);
nand U2523 (N_2523,N_2158,N_2215);
nor U2524 (N_2524,N_1466,N_2014);
xor U2525 (N_2525,N_2207,In_2302);
xor U2526 (N_2526,N_2240,N_2146);
nand U2527 (N_2527,N_2030,N_2234);
xor U2528 (N_2528,N_2352,N_2261);
and U2529 (N_2529,In_1184,N_2395);
and U2530 (N_2530,N_2296,N_2332);
nor U2531 (N_2531,N_2120,N_2367);
nor U2532 (N_2532,N_1809,N_1990);
xnor U2533 (N_2533,N_2386,N_2351);
or U2534 (N_2534,N_2275,N_514);
and U2535 (N_2535,N_454,N_1551);
nor U2536 (N_2536,N_1240,N_1053);
xor U2537 (N_2537,N_2283,N_1821);
nand U2538 (N_2538,N_2398,N_1424);
xor U2539 (N_2539,N_2178,N_2302);
nor U2540 (N_2540,N_1106,N_2108);
nand U2541 (N_2541,N_2370,N_1874);
or U2542 (N_2542,N_2218,N_2349);
nand U2543 (N_2543,N_2248,N_1730);
nand U2544 (N_2544,N_2277,N_911);
xnor U2545 (N_2545,N_2180,N_2055);
nand U2546 (N_2546,N_2242,N_1498);
nor U2547 (N_2547,N_2012,In_607);
nor U2548 (N_2548,N_2122,N_2368);
xor U2549 (N_2549,N_1510,In_2658);
xnor U2550 (N_2550,N_2294,N_2188);
or U2551 (N_2551,N_2306,N_403);
and U2552 (N_2552,N_1649,N_1762);
nor U2553 (N_2553,In_2734,In_384);
nand U2554 (N_2554,N_261,N_83);
nor U2555 (N_2555,N_520,N_2049);
xor U2556 (N_2556,N_2237,N_1844);
nor U2557 (N_2557,N_209,N_2365);
nor U2558 (N_2558,N_2119,N_1435);
nand U2559 (N_2559,N_96,N_974);
xnor U2560 (N_2560,N_1064,In_197);
nand U2561 (N_2561,N_1842,N_815);
and U2562 (N_2562,N_1926,N_2239);
and U2563 (N_2563,N_1088,N_2173);
nor U2564 (N_2564,N_2362,N_2175);
nand U2565 (N_2565,N_2272,In_2151);
nand U2566 (N_2566,N_2081,N_2131);
nor U2567 (N_2567,N_1871,N_1640);
and U2568 (N_2568,N_2317,N_659);
xor U2569 (N_2569,N_2249,In_1555);
nor U2570 (N_2570,N_1635,N_1514);
and U2571 (N_2571,N_1797,N_2044);
and U2572 (N_2572,N_1309,N_2231);
nand U2573 (N_2573,N_1942,N_1128);
xnor U2574 (N_2574,N_1250,N_2185);
nand U2575 (N_2575,N_636,In_2167);
nand U2576 (N_2576,N_2318,N_1707);
nor U2577 (N_2577,N_2285,N_2251);
nand U2578 (N_2578,N_2026,N_2260);
nor U2579 (N_2579,In_2469,N_2348);
nand U2580 (N_2580,In_2584,N_1008);
xor U2581 (N_2581,N_124,N_2179);
nand U2582 (N_2582,In_1420,In_1995);
or U2583 (N_2583,N_632,N_2121);
nand U2584 (N_2584,N_1813,N_1087);
nor U2585 (N_2585,N_2162,In_124);
nor U2586 (N_2586,N_2219,N_1138);
and U2587 (N_2587,N_796,N_2287);
nor U2588 (N_2588,N_1804,N_1633);
nand U2589 (N_2589,N_1694,N_2323);
xnor U2590 (N_2590,N_730,N_1679);
nor U2591 (N_2591,N_2037,N_207);
nor U2592 (N_2592,N_1356,N_2268);
nor U2593 (N_2593,In_193,N_2270);
nand U2594 (N_2594,N_2187,N_2375);
xnor U2595 (N_2595,N_2307,N_1877);
xor U2596 (N_2596,N_2145,N_2135);
nand U2597 (N_2597,N_2238,N_2338);
nand U2598 (N_2598,N_2194,N_2170);
or U2599 (N_2599,N_1856,N_1325);
nor U2600 (N_2600,N_2223,In_2820);
nor U2601 (N_2601,N_2171,N_2469);
nor U2602 (N_2602,N_2418,N_2405);
and U2603 (N_2603,N_1847,In_632);
xnor U2604 (N_2604,N_2116,N_2214);
xor U2605 (N_2605,N_2430,N_2399);
nand U2606 (N_2606,N_2282,N_2421);
nor U2607 (N_2607,In_615,N_2276);
or U2608 (N_2608,N_2572,N_1176);
or U2609 (N_2609,N_2595,N_2366);
and U2610 (N_2610,N_2556,N_2384);
xor U2611 (N_2611,N_2457,N_2485);
nand U2612 (N_2612,N_2599,N_2598);
nand U2613 (N_2613,N_2419,N_604);
or U2614 (N_2614,N_2228,N_2159);
xor U2615 (N_2615,N_1230,N_736);
nand U2616 (N_2616,N_432,N_2558);
nand U2617 (N_2617,N_2413,N_2414);
nand U2618 (N_2618,N_1851,N_2441);
xnor U2619 (N_2619,N_2534,N_2437);
xnor U2620 (N_2620,N_2489,N_2459);
nor U2621 (N_2621,N_2113,N_2501);
and U2622 (N_2622,N_1755,N_1845);
or U2623 (N_2623,N_2543,N_2201);
xor U2624 (N_2624,In_1038,N_2583);
and U2625 (N_2625,N_99,N_2596);
or U2626 (N_2626,N_2328,N_2452);
xor U2627 (N_2627,N_2447,N_2229);
nand U2628 (N_2628,N_2442,N_2580);
xnor U2629 (N_2629,N_1294,N_2403);
nor U2630 (N_2630,N_1834,N_2467);
nor U2631 (N_2631,N_2364,N_2530);
or U2632 (N_2632,In_824,N_2392);
nand U2633 (N_2633,In_2010,N_1820);
nor U2634 (N_2634,N_2523,N_2592);
xor U2635 (N_2635,N_2451,N_1482);
nor U2636 (N_2636,N_2533,N_216);
or U2637 (N_2637,N_2565,N_2148);
nand U2638 (N_2638,N_2591,N_2411);
nand U2639 (N_2639,N_2197,N_2232);
and U2640 (N_2640,In_509,N_2466);
and U2641 (N_2641,N_2241,N_1658);
and U2642 (N_2642,N_2408,N_1396);
xnor U2643 (N_2643,N_2431,N_2284);
xnor U2644 (N_2644,N_2593,N_2472);
xor U2645 (N_2645,N_2444,N_2438);
nor U2646 (N_2646,N_1976,N_2478);
xor U2647 (N_2647,N_2456,N_2344);
nand U2648 (N_2648,N_2246,In_404);
nor U2649 (N_2649,N_2588,N_1639);
nand U2650 (N_2650,N_2547,N_2529);
nor U2651 (N_2651,In_1450,N_2586);
nor U2652 (N_2652,N_2548,N_2559);
and U2653 (N_2653,N_2331,N_2300);
xnor U2654 (N_2654,N_2203,N_2515);
nor U2655 (N_2655,N_2079,N_196);
nand U2656 (N_2656,N_2476,N_2400);
and U2657 (N_2657,N_2422,N_2039);
nand U2658 (N_2658,N_2209,N_2566);
xnor U2659 (N_2659,N_2303,In_1900);
nor U2660 (N_2660,N_2477,N_2484);
nand U2661 (N_2661,N_1444,N_2443);
or U2662 (N_2662,N_2493,In_494);
and U2663 (N_2663,N_2540,N_2521);
and U2664 (N_2664,N_2455,N_2410);
and U2665 (N_2665,N_1292,N_2445);
nor U2666 (N_2666,N_1641,N_2581);
nor U2667 (N_2667,N_2461,N_2357);
or U2668 (N_2668,N_1710,N_2589);
nand U2669 (N_2669,N_2550,N_2401);
or U2670 (N_2670,N_2462,N_2264);
and U2671 (N_2671,N_2504,N_2412);
nor U2672 (N_2672,N_2541,N_2289);
nand U2673 (N_2673,N_2088,N_2130);
xor U2674 (N_2674,N_1198,N_2499);
xor U2675 (N_2675,N_2526,N_2511);
nand U2676 (N_2676,N_2377,N_2382);
xnor U2677 (N_2677,N_2587,N_2524);
nand U2678 (N_2678,In_1512,N_1413);
or U2679 (N_2679,N_2293,N_2552);
nor U2680 (N_2680,N_2463,N_1998);
nor U2681 (N_2681,N_2537,N_2279);
xor U2682 (N_2682,N_2481,N_2329);
or U2683 (N_2683,N_2563,N_2200);
nand U2684 (N_2684,N_2473,N_2434);
and U2685 (N_2685,N_2582,N_2078);
nand U2686 (N_2686,N_2503,N_2460);
or U2687 (N_2687,N_2579,N_2532);
xor U2688 (N_2688,N_2363,N_2340);
nor U2689 (N_2689,N_2574,N_1916);
or U2690 (N_2690,N_2226,N_2502);
xnor U2691 (N_2691,N_2555,N_2527);
or U2692 (N_2692,N_2250,N_2359);
and U2693 (N_2693,N_2500,N_2465);
and U2694 (N_2694,N_2564,N_2325);
nor U2695 (N_2695,N_2520,N_1917);
nand U2696 (N_2696,N_172,N_2199);
or U2697 (N_2697,N_2546,N_2266);
and U2698 (N_2698,N_2104,N_2567);
xnor U2699 (N_2699,N_1716,N_1491);
xor U2700 (N_2700,N_2360,N_724);
nand U2701 (N_2701,N_2420,N_2426);
and U2702 (N_2702,N_2495,N_2322);
xor U2703 (N_2703,N_2545,N_2450);
or U2704 (N_2704,N_2425,N_2577);
nor U2705 (N_2705,N_2498,N_2373);
or U2706 (N_2706,N_2439,N_2212);
and U2707 (N_2707,N_2433,N_2339);
nand U2708 (N_2708,N_2027,N_2518);
nor U2709 (N_2709,N_2561,N_2538);
and U2710 (N_2710,N_2102,N_2406);
or U2711 (N_2711,N_1373,N_2389);
xnor U2712 (N_2712,N_2369,N_2341);
or U2713 (N_2713,In_2760,N_1846);
xnor U2714 (N_2714,N_2570,N_1547);
and U2715 (N_2715,N_2436,N_2312);
xor U2716 (N_2716,N_2562,N_2554);
or U2717 (N_2717,N_2151,N_1816);
nor U2718 (N_2718,N_2482,In_1552);
xor U2719 (N_2719,N_1985,N_2551);
or U2720 (N_2720,N_2585,N_2539);
and U2721 (N_2721,N_2525,N_2449);
and U2722 (N_2722,N_1830,N_2213);
xor U2723 (N_2723,N_2038,N_1897);
nand U2724 (N_2724,N_2062,N_2133);
or U2725 (N_2725,N_2505,N_2343);
nand U2726 (N_2726,N_2429,N_2458);
nand U2727 (N_2727,In_5,N_2571);
or U2728 (N_2728,N_2227,In_144);
and U2729 (N_2729,N_2544,N_2233);
xnor U2730 (N_2730,N_2483,N_2517);
nand U2731 (N_2731,N_947,N_2278);
nand U2732 (N_2732,N_2409,N_2492);
nand U2733 (N_2733,N_2454,N_2475);
nand U2734 (N_2734,N_1485,N_2361);
and U2735 (N_2735,N_1870,N_2404);
xor U2736 (N_2736,N_2255,N_2553);
nor U2737 (N_2737,N_2486,N_2578);
xnor U2738 (N_2738,N_2083,N_2479);
and U2739 (N_2739,N_2516,N_2407);
or U2740 (N_2740,N_2428,N_1789);
or U2741 (N_2741,In_70,N_2573);
nor U2742 (N_2742,N_2568,N_2415);
or U2743 (N_2743,N_2346,N_2334);
nand U2744 (N_2744,In_2357,N_2273);
or U2745 (N_2745,N_2509,N_1775);
xnor U2746 (N_2746,N_2470,N_2597);
nor U2747 (N_2747,N_2519,N_2496);
xor U2748 (N_2748,N_2059,N_2549);
or U2749 (N_2749,N_2480,N_2416);
nand U2750 (N_2750,N_1569,N_2522);
xnor U2751 (N_2751,N_9,N_1223);
nor U2752 (N_2752,N_2262,N_2265);
and U2753 (N_2753,N_1418,N_1790);
and U2754 (N_2754,N_2494,In_646);
nor U2755 (N_2755,N_2286,N_2172);
nand U2756 (N_2756,In_1586,N_2453);
nor U2757 (N_2757,N_2319,N_2247);
and U2758 (N_2758,N_2372,In_2957);
or U2759 (N_2759,N_2423,N_2448);
and U2760 (N_2760,N_2388,In_195);
or U2761 (N_2761,N_2402,N_539);
and U2762 (N_2762,N_2508,N_1776);
nor U2763 (N_2763,N_1909,N_2474);
nand U2764 (N_2764,N_1731,N_1986);
or U2765 (N_2765,N_1627,N_2497);
and U2766 (N_2766,N_2490,N_2514);
or U2767 (N_2767,In_2095,In_63);
xnor U2768 (N_2768,N_2298,N_2394);
or U2769 (N_2769,N_2531,N_2536);
and U2770 (N_2770,N_1242,N_2003);
nor U2771 (N_2771,N_2569,N_2274);
nand U2772 (N_2772,N_2542,N_2506);
nand U2773 (N_2773,N_2309,N_2590);
nor U2774 (N_2774,N_2468,N_2427);
or U2775 (N_2775,N_2424,N_501);
nor U2776 (N_2776,N_2035,N_2321);
nand U2777 (N_2777,N_2487,N_2381);
nand U2778 (N_2778,N_2575,N_2350);
xor U2779 (N_2779,N_2576,N_2417);
xnor U2780 (N_2780,N_2594,In_820);
or U2781 (N_2781,N_2491,N_2143);
and U2782 (N_2782,N_2584,N_2140);
and U2783 (N_2783,N_1946,N_1532);
xor U2784 (N_2784,N_2535,N_2168);
or U2785 (N_2785,N_2557,N_2488);
xnor U2786 (N_2786,N_2507,N_2464);
xnor U2787 (N_2787,N_2435,N_532);
and U2788 (N_2788,N_2560,N_2471);
nor U2789 (N_2789,In_1537,N_2206);
and U2790 (N_2790,N_2252,N_2358);
or U2791 (N_2791,N_558,N_2446);
and U2792 (N_2792,N_2528,N_2288);
xnor U2793 (N_2793,N_2271,N_2111);
and U2794 (N_2794,N_2432,N_2513);
xnor U2795 (N_2795,N_2440,N_2512);
nand U2796 (N_2796,N_1576,N_2510);
or U2797 (N_2797,N_299,N_2028);
nor U2798 (N_2798,N_898,N_2299);
and U2799 (N_2799,N_1118,N_2310);
or U2800 (N_2800,N_2756,N_2632);
nor U2801 (N_2801,N_2721,N_2604);
nor U2802 (N_2802,N_2694,N_2787);
and U2803 (N_2803,N_2736,N_2691);
nand U2804 (N_2804,N_2754,N_2657);
nor U2805 (N_2805,N_2779,N_2705);
and U2806 (N_2806,N_2626,N_2681);
nand U2807 (N_2807,N_2726,N_2675);
xor U2808 (N_2808,N_2695,N_2624);
xor U2809 (N_2809,N_2615,N_2739);
or U2810 (N_2810,N_2761,N_2621);
and U2811 (N_2811,N_2767,N_2640);
and U2812 (N_2812,N_2798,N_2744);
and U2813 (N_2813,N_2762,N_2777);
or U2814 (N_2814,N_2707,N_2783);
nor U2815 (N_2815,N_2785,N_2697);
nand U2816 (N_2816,N_2636,N_2651);
nor U2817 (N_2817,N_2745,N_2631);
nor U2818 (N_2818,N_2720,N_2608);
xnor U2819 (N_2819,N_2637,N_2740);
nor U2820 (N_2820,N_2679,N_2693);
or U2821 (N_2821,N_2627,N_2618);
xor U2822 (N_2822,N_2771,N_2670);
nor U2823 (N_2823,N_2778,N_2698);
and U2824 (N_2824,N_2799,N_2750);
xnor U2825 (N_2825,N_2704,N_2642);
xor U2826 (N_2826,N_2710,N_2663);
and U2827 (N_2827,N_2752,N_2669);
xor U2828 (N_2828,N_2641,N_2743);
nor U2829 (N_2829,N_2727,N_2732);
nor U2830 (N_2830,N_2639,N_2620);
and U2831 (N_2831,N_2729,N_2759);
xnor U2832 (N_2832,N_2780,N_2737);
nor U2833 (N_2833,N_2605,N_2746);
nand U2834 (N_2834,N_2687,N_2645);
or U2835 (N_2835,N_2765,N_2775);
xnor U2836 (N_2836,N_2725,N_2661);
nand U2837 (N_2837,N_2797,N_2635);
or U2838 (N_2838,N_2706,N_2610);
nand U2839 (N_2839,N_2749,N_2611);
nand U2840 (N_2840,N_2617,N_2760);
nand U2841 (N_2841,N_2680,N_2728);
or U2842 (N_2842,N_2703,N_2602);
nand U2843 (N_2843,N_2688,N_2763);
nor U2844 (N_2844,N_2731,N_2716);
nor U2845 (N_2845,N_2646,N_2796);
xnor U2846 (N_2846,N_2733,N_2794);
xor U2847 (N_2847,N_2724,N_2690);
nor U2848 (N_2848,N_2723,N_2711);
xnor U2849 (N_2849,N_2676,N_2689);
nand U2850 (N_2850,N_2672,N_2658);
and U2851 (N_2851,N_2623,N_2748);
and U2852 (N_2852,N_2792,N_2769);
nor U2853 (N_2853,N_2768,N_2677);
nand U2854 (N_2854,N_2648,N_2644);
nor U2855 (N_2855,N_2758,N_2664);
xnor U2856 (N_2856,N_2666,N_2629);
and U2857 (N_2857,N_2738,N_2685);
xor U2858 (N_2858,N_2766,N_2678);
nand U2859 (N_2859,N_2730,N_2702);
nand U2860 (N_2860,N_2751,N_2671);
or U2861 (N_2861,N_2795,N_2628);
nor U2862 (N_2862,N_2742,N_2782);
nor U2863 (N_2863,N_2786,N_2665);
nand U2864 (N_2864,N_2790,N_2655);
nor U2865 (N_2865,N_2619,N_2789);
nor U2866 (N_2866,N_2699,N_2653);
and U2867 (N_2867,N_2791,N_2638);
or U2868 (N_2868,N_2757,N_2607);
nor U2869 (N_2869,N_2741,N_2659);
and U2870 (N_2870,N_2696,N_2734);
nor U2871 (N_2871,N_2643,N_2715);
or U2872 (N_2872,N_2634,N_2674);
or U2873 (N_2873,N_2770,N_2708);
nand U2874 (N_2874,N_2719,N_2709);
nor U2875 (N_2875,N_2753,N_2601);
and U2876 (N_2876,N_2660,N_2647);
nor U2877 (N_2877,N_2625,N_2701);
and U2878 (N_2878,N_2683,N_2686);
nand U2879 (N_2879,N_2772,N_2735);
nor U2880 (N_2880,N_2612,N_2793);
nand U2881 (N_2881,N_2722,N_2684);
and U2882 (N_2882,N_2656,N_2654);
and U2883 (N_2883,N_2667,N_2630);
xor U2884 (N_2884,N_2781,N_2717);
and U2885 (N_2885,N_2614,N_2700);
nand U2886 (N_2886,N_2668,N_2633);
xnor U2887 (N_2887,N_2788,N_2692);
nor U2888 (N_2888,N_2600,N_2603);
xnor U2889 (N_2889,N_2682,N_2609);
nand U2890 (N_2890,N_2774,N_2649);
or U2891 (N_2891,N_2652,N_2606);
xor U2892 (N_2892,N_2713,N_2764);
xnor U2893 (N_2893,N_2784,N_2673);
nor U2894 (N_2894,N_2613,N_2662);
nand U2895 (N_2895,N_2755,N_2718);
xnor U2896 (N_2896,N_2773,N_2622);
and U2897 (N_2897,N_2776,N_2616);
nor U2898 (N_2898,N_2712,N_2650);
or U2899 (N_2899,N_2714,N_2747);
and U2900 (N_2900,N_2704,N_2764);
or U2901 (N_2901,N_2686,N_2768);
or U2902 (N_2902,N_2707,N_2646);
nand U2903 (N_2903,N_2686,N_2777);
and U2904 (N_2904,N_2631,N_2656);
or U2905 (N_2905,N_2786,N_2653);
and U2906 (N_2906,N_2721,N_2633);
nor U2907 (N_2907,N_2656,N_2700);
and U2908 (N_2908,N_2684,N_2765);
nor U2909 (N_2909,N_2671,N_2635);
nand U2910 (N_2910,N_2681,N_2766);
nor U2911 (N_2911,N_2646,N_2630);
nand U2912 (N_2912,N_2667,N_2730);
or U2913 (N_2913,N_2779,N_2706);
or U2914 (N_2914,N_2779,N_2624);
and U2915 (N_2915,N_2618,N_2720);
and U2916 (N_2916,N_2627,N_2694);
nor U2917 (N_2917,N_2724,N_2732);
nand U2918 (N_2918,N_2631,N_2728);
nand U2919 (N_2919,N_2719,N_2769);
and U2920 (N_2920,N_2660,N_2661);
and U2921 (N_2921,N_2688,N_2614);
nand U2922 (N_2922,N_2647,N_2671);
xnor U2923 (N_2923,N_2640,N_2666);
nor U2924 (N_2924,N_2659,N_2740);
or U2925 (N_2925,N_2724,N_2682);
or U2926 (N_2926,N_2782,N_2659);
and U2927 (N_2927,N_2771,N_2607);
xnor U2928 (N_2928,N_2603,N_2796);
xnor U2929 (N_2929,N_2759,N_2772);
nor U2930 (N_2930,N_2687,N_2718);
and U2931 (N_2931,N_2735,N_2629);
nor U2932 (N_2932,N_2626,N_2643);
and U2933 (N_2933,N_2695,N_2765);
xor U2934 (N_2934,N_2700,N_2650);
or U2935 (N_2935,N_2648,N_2756);
nor U2936 (N_2936,N_2719,N_2767);
xor U2937 (N_2937,N_2700,N_2721);
nor U2938 (N_2938,N_2723,N_2632);
or U2939 (N_2939,N_2784,N_2787);
or U2940 (N_2940,N_2665,N_2663);
and U2941 (N_2941,N_2648,N_2629);
or U2942 (N_2942,N_2658,N_2724);
nor U2943 (N_2943,N_2735,N_2720);
xnor U2944 (N_2944,N_2672,N_2730);
nand U2945 (N_2945,N_2713,N_2729);
nor U2946 (N_2946,N_2751,N_2784);
nor U2947 (N_2947,N_2712,N_2688);
xor U2948 (N_2948,N_2654,N_2614);
or U2949 (N_2949,N_2775,N_2779);
or U2950 (N_2950,N_2646,N_2768);
and U2951 (N_2951,N_2792,N_2658);
or U2952 (N_2952,N_2606,N_2641);
xor U2953 (N_2953,N_2658,N_2638);
xor U2954 (N_2954,N_2628,N_2742);
xor U2955 (N_2955,N_2647,N_2763);
and U2956 (N_2956,N_2609,N_2683);
and U2957 (N_2957,N_2716,N_2677);
and U2958 (N_2958,N_2778,N_2799);
or U2959 (N_2959,N_2637,N_2708);
xor U2960 (N_2960,N_2655,N_2640);
xor U2961 (N_2961,N_2742,N_2744);
nor U2962 (N_2962,N_2757,N_2721);
xnor U2963 (N_2963,N_2769,N_2677);
xnor U2964 (N_2964,N_2791,N_2645);
xnor U2965 (N_2965,N_2776,N_2603);
xnor U2966 (N_2966,N_2608,N_2743);
or U2967 (N_2967,N_2653,N_2798);
and U2968 (N_2968,N_2641,N_2731);
nor U2969 (N_2969,N_2765,N_2631);
or U2970 (N_2970,N_2652,N_2646);
xor U2971 (N_2971,N_2626,N_2637);
and U2972 (N_2972,N_2659,N_2649);
nor U2973 (N_2973,N_2764,N_2743);
nand U2974 (N_2974,N_2791,N_2624);
or U2975 (N_2975,N_2613,N_2640);
nand U2976 (N_2976,N_2626,N_2684);
and U2977 (N_2977,N_2799,N_2786);
nor U2978 (N_2978,N_2621,N_2643);
and U2979 (N_2979,N_2772,N_2763);
xor U2980 (N_2980,N_2729,N_2620);
nor U2981 (N_2981,N_2710,N_2725);
nor U2982 (N_2982,N_2692,N_2605);
nor U2983 (N_2983,N_2792,N_2683);
or U2984 (N_2984,N_2602,N_2693);
nand U2985 (N_2985,N_2627,N_2647);
nor U2986 (N_2986,N_2711,N_2604);
and U2987 (N_2987,N_2704,N_2724);
and U2988 (N_2988,N_2730,N_2775);
and U2989 (N_2989,N_2721,N_2703);
and U2990 (N_2990,N_2758,N_2739);
xor U2991 (N_2991,N_2634,N_2790);
nand U2992 (N_2992,N_2604,N_2627);
nand U2993 (N_2993,N_2682,N_2634);
xnor U2994 (N_2994,N_2728,N_2727);
nand U2995 (N_2995,N_2745,N_2705);
and U2996 (N_2996,N_2642,N_2762);
nor U2997 (N_2997,N_2754,N_2600);
and U2998 (N_2998,N_2784,N_2642);
nand U2999 (N_2999,N_2657,N_2649);
and U3000 (N_3000,N_2930,N_2844);
nor U3001 (N_3001,N_2883,N_2869);
nor U3002 (N_3002,N_2903,N_2982);
nand U3003 (N_3003,N_2898,N_2858);
xor U3004 (N_3004,N_2966,N_2814);
nor U3005 (N_3005,N_2948,N_2839);
and U3006 (N_3006,N_2905,N_2983);
nor U3007 (N_3007,N_2841,N_2893);
xnor U3008 (N_3008,N_2807,N_2840);
and U3009 (N_3009,N_2846,N_2963);
and U3010 (N_3010,N_2877,N_2917);
xnor U3011 (N_3011,N_2927,N_2842);
nand U3012 (N_3012,N_2936,N_2934);
xnor U3013 (N_3013,N_2899,N_2811);
nor U3014 (N_3014,N_2831,N_2856);
and U3015 (N_3015,N_2889,N_2955);
and U3016 (N_3016,N_2808,N_2829);
xnor U3017 (N_3017,N_2981,N_2988);
nand U3018 (N_3018,N_2824,N_2896);
or U3019 (N_3019,N_2962,N_2822);
and U3020 (N_3020,N_2993,N_2880);
and U3021 (N_3021,N_2901,N_2876);
xnor U3022 (N_3022,N_2892,N_2951);
and U3023 (N_3023,N_2915,N_2870);
nor U3024 (N_3024,N_2868,N_2851);
or U3025 (N_3025,N_2830,N_2859);
nand U3026 (N_3026,N_2912,N_2849);
and U3027 (N_3027,N_2825,N_2800);
or U3028 (N_3028,N_2989,N_2873);
nand U3029 (N_3029,N_2996,N_2897);
nor U3030 (N_3030,N_2823,N_2909);
nor U3031 (N_3031,N_2965,N_2960);
nor U3032 (N_3032,N_2956,N_2910);
and U3033 (N_3033,N_2837,N_2947);
xnor U3034 (N_3034,N_2959,N_2997);
and U3035 (N_3035,N_2806,N_2994);
nor U3036 (N_3036,N_2933,N_2843);
nand U3037 (N_3037,N_2815,N_2872);
and U3038 (N_3038,N_2967,N_2838);
nor U3039 (N_3039,N_2961,N_2921);
xnor U3040 (N_3040,N_2946,N_2802);
or U3041 (N_3041,N_2976,N_2950);
or U3042 (N_3042,N_2939,N_2801);
nor U3043 (N_3043,N_2971,N_2879);
nand U3044 (N_3044,N_2954,N_2958);
nand U3045 (N_3045,N_2866,N_2826);
and U3046 (N_3046,N_2977,N_2985);
xnor U3047 (N_3047,N_2827,N_2875);
and U3048 (N_3048,N_2862,N_2820);
or U3049 (N_3049,N_2845,N_2940);
nor U3050 (N_3050,N_2992,N_2925);
nand U3051 (N_3051,N_2902,N_2894);
nor U3052 (N_3052,N_2860,N_2972);
nand U3053 (N_3053,N_2973,N_2855);
or U3054 (N_3054,N_2987,N_2979);
nand U3055 (N_3055,N_2864,N_2881);
or U3056 (N_3056,N_2920,N_2874);
nand U3057 (N_3057,N_2968,N_2949);
or U3058 (N_3058,N_2813,N_2978);
nor U3059 (N_3059,N_2836,N_2803);
nand U3060 (N_3060,N_2945,N_2888);
and U3061 (N_3061,N_2919,N_2891);
xnor U3062 (N_3062,N_2964,N_2931);
xor U3063 (N_3063,N_2904,N_2911);
xnor U3064 (N_3064,N_2857,N_2913);
xnor U3065 (N_3065,N_2929,N_2926);
nor U3066 (N_3066,N_2928,N_2995);
and U3067 (N_3067,N_2944,N_2907);
nand U3068 (N_3068,N_2882,N_2974);
nor U3069 (N_3069,N_2908,N_2835);
xor U3070 (N_3070,N_2834,N_2812);
or U3071 (N_3071,N_2818,N_2980);
nand U3072 (N_3072,N_2938,N_2942);
xnor U3073 (N_3073,N_2885,N_2999);
xor U3074 (N_3074,N_2865,N_2819);
nand U3075 (N_3075,N_2867,N_2853);
nor U3076 (N_3076,N_2918,N_2854);
and U3077 (N_3077,N_2887,N_2817);
nand U3078 (N_3078,N_2991,N_2861);
nor U3079 (N_3079,N_2914,N_2937);
and U3080 (N_3080,N_2922,N_2941);
xnor U3081 (N_3081,N_2906,N_2804);
nor U3082 (N_3082,N_2969,N_2828);
nor U3083 (N_3083,N_2863,N_2809);
nand U3084 (N_3084,N_2986,N_2953);
nand U3085 (N_3085,N_2900,N_2878);
and U3086 (N_3086,N_2821,N_2833);
or U3087 (N_3087,N_2847,N_2805);
xnor U3088 (N_3088,N_2890,N_2810);
nand U3089 (N_3089,N_2884,N_2970);
and U3090 (N_3090,N_2871,N_2975);
nand U3091 (N_3091,N_2832,N_2957);
and U3092 (N_3092,N_2916,N_2852);
nand U3093 (N_3093,N_2935,N_2943);
nor U3094 (N_3094,N_2984,N_2848);
xnor U3095 (N_3095,N_2990,N_2850);
xor U3096 (N_3096,N_2886,N_2952);
and U3097 (N_3097,N_2816,N_2998);
or U3098 (N_3098,N_2924,N_2923);
nor U3099 (N_3099,N_2895,N_2932);
xor U3100 (N_3100,N_2897,N_2920);
or U3101 (N_3101,N_2874,N_2993);
and U3102 (N_3102,N_2993,N_2914);
nor U3103 (N_3103,N_2911,N_2810);
and U3104 (N_3104,N_2856,N_2868);
or U3105 (N_3105,N_2905,N_2881);
nand U3106 (N_3106,N_2870,N_2970);
nand U3107 (N_3107,N_2821,N_2988);
nor U3108 (N_3108,N_2965,N_2961);
xnor U3109 (N_3109,N_2822,N_2955);
nor U3110 (N_3110,N_2927,N_2925);
or U3111 (N_3111,N_2938,N_2812);
or U3112 (N_3112,N_2928,N_2921);
nand U3113 (N_3113,N_2808,N_2893);
or U3114 (N_3114,N_2871,N_2935);
and U3115 (N_3115,N_2949,N_2848);
nor U3116 (N_3116,N_2924,N_2952);
or U3117 (N_3117,N_2870,N_2909);
nand U3118 (N_3118,N_2842,N_2934);
nor U3119 (N_3119,N_2954,N_2872);
nand U3120 (N_3120,N_2815,N_2933);
xor U3121 (N_3121,N_2943,N_2897);
nand U3122 (N_3122,N_2898,N_2933);
and U3123 (N_3123,N_2994,N_2960);
or U3124 (N_3124,N_2938,N_2993);
xnor U3125 (N_3125,N_2901,N_2938);
nand U3126 (N_3126,N_2976,N_2991);
and U3127 (N_3127,N_2881,N_2821);
or U3128 (N_3128,N_2815,N_2972);
nand U3129 (N_3129,N_2964,N_2999);
or U3130 (N_3130,N_2809,N_2910);
nand U3131 (N_3131,N_2824,N_2840);
xnor U3132 (N_3132,N_2911,N_2840);
and U3133 (N_3133,N_2843,N_2807);
nand U3134 (N_3134,N_2805,N_2818);
xor U3135 (N_3135,N_2949,N_2831);
xnor U3136 (N_3136,N_2896,N_2909);
xor U3137 (N_3137,N_2972,N_2914);
nand U3138 (N_3138,N_2864,N_2875);
xnor U3139 (N_3139,N_2859,N_2939);
and U3140 (N_3140,N_2960,N_2997);
or U3141 (N_3141,N_2970,N_2929);
and U3142 (N_3142,N_2990,N_2816);
xor U3143 (N_3143,N_2880,N_2803);
nand U3144 (N_3144,N_2879,N_2937);
and U3145 (N_3145,N_2923,N_2845);
nand U3146 (N_3146,N_2913,N_2802);
and U3147 (N_3147,N_2898,N_2937);
and U3148 (N_3148,N_2882,N_2833);
nand U3149 (N_3149,N_2888,N_2803);
xor U3150 (N_3150,N_2843,N_2828);
and U3151 (N_3151,N_2993,N_2896);
nor U3152 (N_3152,N_2945,N_2956);
and U3153 (N_3153,N_2962,N_2865);
nor U3154 (N_3154,N_2931,N_2884);
xnor U3155 (N_3155,N_2855,N_2845);
or U3156 (N_3156,N_2834,N_2883);
xor U3157 (N_3157,N_2842,N_2886);
xor U3158 (N_3158,N_2863,N_2938);
xnor U3159 (N_3159,N_2848,N_2989);
or U3160 (N_3160,N_2908,N_2824);
xor U3161 (N_3161,N_2829,N_2896);
nor U3162 (N_3162,N_2825,N_2940);
nand U3163 (N_3163,N_2990,N_2910);
xnor U3164 (N_3164,N_2889,N_2956);
and U3165 (N_3165,N_2813,N_2833);
nand U3166 (N_3166,N_2947,N_2962);
nor U3167 (N_3167,N_2905,N_2997);
nor U3168 (N_3168,N_2944,N_2823);
nor U3169 (N_3169,N_2948,N_2942);
or U3170 (N_3170,N_2956,N_2978);
and U3171 (N_3171,N_2986,N_2971);
or U3172 (N_3172,N_2945,N_2964);
nor U3173 (N_3173,N_2953,N_2941);
nand U3174 (N_3174,N_2828,N_2861);
or U3175 (N_3175,N_2992,N_2922);
xnor U3176 (N_3176,N_2965,N_2852);
nand U3177 (N_3177,N_2860,N_2941);
or U3178 (N_3178,N_2848,N_2922);
nand U3179 (N_3179,N_2996,N_2966);
nand U3180 (N_3180,N_2860,N_2908);
nand U3181 (N_3181,N_2947,N_2896);
or U3182 (N_3182,N_2837,N_2821);
nor U3183 (N_3183,N_2890,N_2881);
xnor U3184 (N_3184,N_2946,N_2902);
nand U3185 (N_3185,N_2827,N_2908);
or U3186 (N_3186,N_2863,N_2835);
or U3187 (N_3187,N_2939,N_2995);
nand U3188 (N_3188,N_2970,N_2811);
or U3189 (N_3189,N_2865,N_2898);
nor U3190 (N_3190,N_2973,N_2870);
nand U3191 (N_3191,N_2867,N_2886);
nand U3192 (N_3192,N_2803,N_2846);
nand U3193 (N_3193,N_2859,N_2990);
nand U3194 (N_3194,N_2890,N_2827);
and U3195 (N_3195,N_2893,N_2889);
nand U3196 (N_3196,N_2816,N_2870);
and U3197 (N_3197,N_2973,N_2838);
xnor U3198 (N_3198,N_2922,N_2967);
nand U3199 (N_3199,N_2811,N_2873);
nor U3200 (N_3200,N_3113,N_3140);
xnor U3201 (N_3201,N_3179,N_3102);
nand U3202 (N_3202,N_3144,N_3164);
nor U3203 (N_3203,N_3111,N_3183);
nand U3204 (N_3204,N_3075,N_3105);
or U3205 (N_3205,N_3193,N_3044);
nor U3206 (N_3206,N_3172,N_3199);
nand U3207 (N_3207,N_3117,N_3191);
and U3208 (N_3208,N_3133,N_3024);
or U3209 (N_3209,N_3167,N_3054);
and U3210 (N_3210,N_3171,N_3166);
nand U3211 (N_3211,N_3168,N_3196);
nand U3212 (N_3212,N_3066,N_3156);
nor U3213 (N_3213,N_3148,N_3058);
nor U3214 (N_3214,N_3143,N_3136);
nand U3215 (N_3215,N_3047,N_3122);
nand U3216 (N_3216,N_3000,N_3025);
nand U3217 (N_3217,N_3173,N_3026);
and U3218 (N_3218,N_3006,N_3003);
nor U3219 (N_3219,N_3197,N_3083);
or U3220 (N_3220,N_3021,N_3126);
nand U3221 (N_3221,N_3190,N_3112);
xnor U3222 (N_3222,N_3028,N_3005);
nor U3223 (N_3223,N_3062,N_3125);
nand U3224 (N_3224,N_3115,N_3162);
nand U3225 (N_3225,N_3084,N_3081);
nand U3226 (N_3226,N_3157,N_3029);
xor U3227 (N_3227,N_3187,N_3192);
nand U3228 (N_3228,N_3034,N_3063);
nor U3229 (N_3229,N_3068,N_3139);
or U3230 (N_3230,N_3001,N_3060);
nand U3231 (N_3231,N_3134,N_3077);
nand U3232 (N_3232,N_3169,N_3056);
nor U3233 (N_3233,N_3076,N_3118);
nand U3234 (N_3234,N_3040,N_3067);
nand U3235 (N_3235,N_3004,N_3074);
nor U3236 (N_3236,N_3051,N_3178);
nand U3237 (N_3237,N_3095,N_3163);
and U3238 (N_3238,N_3131,N_3093);
nor U3239 (N_3239,N_3107,N_3079);
xnor U3240 (N_3240,N_3036,N_3155);
and U3241 (N_3241,N_3033,N_3100);
or U3242 (N_3242,N_3008,N_3186);
nor U3243 (N_3243,N_3045,N_3127);
or U3244 (N_3244,N_3038,N_3061);
or U3245 (N_3245,N_3072,N_3154);
xor U3246 (N_3246,N_3142,N_3039);
and U3247 (N_3247,N_3007,N_3094);
nand U3248 (N_3248,N_3009,N_3129);
nor U3249 (N_3249,N_3035,N_3141);
nor U3250 (N_3250,N_3106,N_3046);
or U3251 (N_3251,N_3052,N_3069);
nand U3252 (N_3252,N_3032,N_3120);
and U3253 (N_3253,N_3091,N_3119);
and U3254 (N_3254,N_3145,N_3014);
or U3255 (N_3255,N_3099,N_3110);
xnor U3256 (N_3256,N_3124,N_3177);
and U3257 (N_3257,N_3088,N_3059);
nand U3258 (N_3258,N_3086,N_3188);
nand U3259 (N_3259,N_3055,N_3104);
xor U3260 (N_3260,N_3185,N_3082);
xnor U3261 (N_3261,N_3050,N_3108);
xnor U3262 (N_3262,N_3037,N_3116);
or U3263 (N_3263,N_3031,N_3096);
nand U3264 (N_3264,N_3138,N_3174);
nand U3265 (N_3265,N_3073,N_3194);
or U3266 (N_3266,N_3152,N_3195);
or U3267 (N_3267,N_3130,N_3098);
and U3268 (N_3268,N_3153,N_3176);
or U3269 (N_3269,N_3146,N_3182);
xor U3270 (N_3270,N_3023,N_3048);
xor U3271 (N_3271,N_3010,N_3070);
nor U3272 (N_3272,N_3103,N_3041);
and U3273 (N_3273,N_3128,N_3158);
nor U3274 (N_3274,N_3097,N_3198);
or U3275 (N_3275,N_3042,N_3180);
or U3276 (N_3276,N_3022,N_3150);
nand U3277 (N_3277,N_3064,N_3019);
or U3278 (N_3278,N_3012,N_3085);
nor U3279 (N_3279,N_3017,N_3175);
nor U3280 (N_3280,N_3149,N_3101);
nand U3281 (N_3281,N_3087,N_3132);
nand U3282 (N_3282,N_3049,N_3137);
xor U3283 (N_3283,N_3057,N_3165);
and U3284 (N_3284,N_3011,N_3123);
or U3285 (N_3285,N_3147,N_3020);
xor U3286 (N_3286,N_3109,N_3159);
nor U3287 (N_3287,N_3015,N_3018);
nand U3288 (N_3288,N_3065,N_3053);
and U3289 (N_3289,N_3151,N_3092);
or U3290 (N_3290,N_3089,N_3016);
xor U3291 (N_3291,N_3080,N_3135);
and U3292 (N_3292,N_3181,N_3170);
xnor U3293 (N_3293,N_3114,N_3160);
xnor U3294 (N_3294,N_3090,N_3161);
nand U3295 (N_3295,N_3189,N_3013);
and U3296 (N_3296,N_3184,N_3027);
nand U3297 (N_3297,N_3030,N_3078);
nor U3298 (N_3298,N_3002,N_3121);
nand U3299 (N_3299,N_3043,N_3071);
nor U3300 (N_3300,N_3117,N_3062);
xnor U3301 (N_3301,N_3074,N_3062);
nor U3302 (N_3302,N_3178,N_3126);
nand U3303 (N_3303,N_3068,N_3129);
nor U3304 (N_3304,N_3068,N_3001);
nor U3305 (N_3305,N_3171,N_3037);
xor U3306 (N_3306,N_3008,N_3019);
nor U3307 (N_3307,N_3079,N_3012);
nor U3308 (N_3308,N_3008,N_3172);
nand U3309 (N_3309,N_3179,N_3096);
xor U3310 (N_3310,N_3076,N_3173);
or U3311 (N_3311,N_3171,N_3001);
and U3312 (N_3312,N_3189,N_3068);
nand U3313 (N_3313,N_3125,N_3132);
or U3314 (N_3314,N_3078,N_3151);
nor U3315 (N_3315,N_3115,N_3188);
xor U3316 (N_3316,N_3107,N_3005);
nand U3317 (N_3317,N_3025,N_3178);
nor U3318 (N_3318,N_3047,N_3017);
nand U3319 (N_3319,N_3067,N_3110);
nor U3320 (N_3320,N_3106,N_3034);
nand U3321 (N_3321,N_3172,N_3056);
nor U3322 (N_3322,N_3031,N_3170);
and U3323 (N_3323,N_3169,N_3004);
or U3324 (N_3324,N_3076,N_3132);
xnor U3325 (N_3325,N_3118,N_3064);
nand U3326 (N_3326,N_3001,N_3092);
nor U3327 (N_3327,N_3164,N_3170);
nand U3328 (N_3328,N_3052,N_3006);
nor U3329 (N_3329,N_3069,N_3102);
nor U3330 (N_3330,N_3093,N_3194);
or U3331 (N_3331,N_3080,N_3050);
nor U3332 (N_3332,N_3036,N_3083);
and U3333 (N_3333,N_3004,N_3192);
xnor U3334 (N_3334,N_3010,N_3191);
nor U3335 (N_3335,N_3064,N_3094);
or U3336 (N_3336,N_3186,N_3173);
nand U3337 (N_3337,N_3135,N_3140);
or U3338 (N_3338,N_3049,N_3031);
nand U3339 (N_3339,N_3122,N_3196);
or U3340 (N_3340,N_3035,N_3016);
or U3341 (N_3341,N_3163,N_3151);
nand U3342 (N_3342,N_3089,N_3131);
nand U3343 (N_3343,N_3141,N_3188);
nand U3344 (N_3344,N_3077,N_3102);
nor U3345 (N_3345,N_3027,N_3126);
nor U3346 (N_3346,N_3062,N_3186);
xnor U3347 (N_3347,N_3146,N_3054);
and U3348 (N_3348,N_3028,N_3187);
and U3349 (N_3349,N_3172,N_3193);
nand U3350 (N_3350,N_3057,N_3027);
xor U3351 (N_3351,N_3062,N_3105);
or U3352 (N_3352,N_3178,N_3133);
or U3353 (N_3353,N_3182,N_3079);
nand U3354 (N_3354,N_3150,N_3186);
and U3355 (N_3355,N_3159,N_3040);
xnor U3356 (N_3356,N_3138,N_3132);
or U3357 (N_3357,N_3184,N_3041);
xor U3358 (N_3358,N_3099,N_3137);
or U3359 (N_3359,N_3113,N_3015);
or U3360 (N_3360,N_3177,N_3100);
xor U3361 (N_3361,N_3173,N_3016);
nor U3362 (N_3362,N_3147,N_3151);
xnor U3363 (N_3363,N_3033,N_3157);
or U3364 (N_3364,N_3198,N_3117);
nor U3365 (N_3365,N_3120,N_3074);
nor U3366 (N_3366,N_3124,N_3160);
nor U3367 (N_3367,N_3116,N_3199);
nand U3368 (N_3368,N_3103,N_3099);
nand U3369 (N_3369,N_3086,N_3055);
xnor U3370 (N_3370,N_3132,N_3082);
nand U3371 (N_3371,N_3121,N_3198);
xor U3372 (N_3372,N_3057,N_3189);
nor U3373 (N_3373,N_3063,N_3004);
xnor U3374 (N_3374,N_3133,N_3164);
nand U3375 (N_3375,N_3178,N_3067);
and U3376 (N_3376,N_3091,N_3083);
and U3377 (N_3377,N_3005,N_3185);
xnor U3378 (N_3378,N_3046,N_3176);
or U3379 (N_3379,N_3122,N_3128);
nor U3380 (N_3380,N_3119,N_3170);
nor U3381 (N_3381,N_3041,N_3053);
or U3382 (N_3382,N_3014,N_3067);
nand U3383 (N_3383,N_3068,N_3178);
xor U3384 (N_3384,N_3104,N_3125);
or U3385 (N_3385,N_3044,N_3136);
xnor U3386 (N_3386,N_3187,N_3132);
and U3387 (N_3387,N_3138,N_3126);
or U3388 (N_3388,N_3000,N_3162);
nand U3389 (N_3389,N_3088,N_3122);
nor U3390 (N_3390,N_3126,N_3166);
and U3391 (N_3391,N_3085,N_3122);
and U3392 (N_3392,N_3179,N_3160);
or U3393 (N_3393,N_3045,N_3019);
and U3394 (N_3394,N_3197,N_3114);
nand U3395 (N_3395,N_3083,N_3193);
and U3396 (N_3396,N_3112,N_3098);
and U3397 (N_3397,N_3068,N_3006);
or U3398 (N_3398,N_3180,N_3034);
nor U3399 (N_3399,N_3057,N_3192);
nand U3400 (N_3400,N_3318,N_3371);
nand U3401 (N_3401,N_3352,N_3280);
nand U3402 (N_3402,N_3309,N_3209);
xnor U3403 (N_3403,N_3340,N_3338);
xor U3404 (N_3404,N_3238,N_3216);
nor U3405 (N_3405,N_3291,N_3233);
and U3406 (N_3406,N_3239,N_3248);
nand U3407 (N_3407,N_3220,N_3255);
xor U3408 (N_3408,N_3213,N_3336);
nor U3409 (N_3409,N_3296,N_3237);
xor U3410 (N_3410,N_3397,N_3387);
and U3411 (N_3411,N_3288,N_3279);
or U3412 (N_3412,N_3268,N_3315);
and U3413 (N_3413,N_3393,N_3210);
xnor U3414 (N_3414,N_3326,N_3354);
nand U3415 (N_3415,N_3365,N_3205);
or U3416 (N_3416,N_3339,N_3258);
or U3417 (N_3417,N_3359,N_3245);
xnor U3418 (N_3418,N_3289,N_3388);
and U3419 (N_3419,N_3277,N_3232);
nand U3420 (N_3420,N_3287,N_3240);
or U3421 (N_3421,N_3379,N_3310);
xnor U3422 (N_3422,N_3269,N_3367);
nor U3423 (N_3423,N_3314,N_3254);
xnor U3424 (N_3424,N_3283,N_3218);
nand U3425 (N_3425,N_3284,N_3293);
xor U3426 (N_3426,N_3350,N_3368);
and U3427 (N_3427,N_3380,N_3271);
and U3428 (N_3428,N_3300,N_3235);
and U3429 (N_3429,N_3321,N_3249);
or U3430 (N_3430,N_3372,N_3250);
xor U3431 (N_3431,N_3259,N_3217);
nor U3432 (N_3432,N_3341,N_3215);
or U3433 (N_3433,N_3301,N_3317);
xnor U3434 (N_3434,N_3332,N_3224);
nand U3435 (N_3435,N_3292,N_3234);
xnor U3436 (N_3436,N_3261,N_3211);
and U3437 (N_3437,N_3323,N_3312);
and U3438 (N_3438,N_3353,N_3394);
nand U3439 (N_3439,N_3230,N_3247);
nand U3440 (N_3440,N_3319,N_3242);
and U3441 (N_3441,N_3222,N_3355);
or U3442 (N_3442,N_3256,N_3363);
nor U3443 (N_3443,N_3270,N_3334);
nand U3444 (N_3444,N_3398,N_3327);
xnor U3445 (N_3445,N_3274,N_3275);
or U3446 (N_3446,N_3236,N_3399);
nor U3447 (N_3447,N_3223,N_3252);
nor U3448 (N_3448,N_3200,N_3281);
nor U3449 (N_3449,N_3297,N_3201);
and U3450 (N_3450,N_3349,N_3335);
nor U3451 (N_3451,N_3361,N_3266);
or U3452 (N_3452,N_3212,N_3263);
xor U3453 (N_3453,N_3386,N_3313);
xor U3454 (N_3454,N_3303,N_3290);
and U3455 (N_3455,N_3364,N_3298);
nand U3456 (N_3456,N_3294,N_3357);
xor U3457 (N_3457,N_3251,N_3241);
and U3458 (N_3458,N_3366,N_3356);
and U3459 (N_3459,N_3342,N_3381);
and U3460 (N_3460,N_3203,N_3304);
nor U3461 (N_3461,N_3362,N_3351);
nor U3462 (N_3462,N_3331,N_3337);
nand U3463 (N_3463,N_3378,N_3396);
or U3464 (N_3464,N_3390,N_3295);
and U3465 (N_3465,N_3308,N_3276);
nor U3466 (N_3466,N_3302,N_3243);
nand U3467 (N_3467,N_3273,N_3330);
xor U3468 (N_3468,N_3391,N_3329);
nor U3469 (N_3469,N_3262,N_3225);
or U3470 (N_3470,N_3376,N_3265);
nor U3471 (N_3471,N_3369,N_3320);
nor U3472 (N_3472,N_3374,N_3253);
and U3473 (N_3473,N_3347,N_3227);
xor U3474 (N_3474,N_3219,N_3395);
or U3475 (N_3475,N_3316,N_3324);
nor U3476 (N_3476,N_3373,N_3383);
xnor U3477 (N_3477,N_3392,N_3343);
or U3478 (N_3478,N_3344,N_3267);
nor U3479 (N_3479,N_3272,N_3382);
nand U3480 (N_3480,N_3285,N_3231);
nor U3481 (N_3481,N_3360,N_3286);
or U3482 (N_3482,N_3260,N_3264);
nor U3483 (N_3483,N_3375,N_3299);
and U3484 (N_3484,N_3389,N_3206);
nor U3485 (N_3485,N_3370,N_3328);
nand U3486 (N_3486,N_3384,N_3377);
nand U3487 (N_3487,N_3348,N_3226);
nor U3488 (N_3488,N_3306,N_3257);
nor U3489 (N_3489,N_3346,N_3307);
nand U3490 (N_3490,N_3214,N_3246);
or U3491 (N_3491,N_3202,N_3311);
or U3492 (N_3492,N_3229,N_3204);
nor U3493 (N_3493,N_3228,N_3385);
nand U3494 (N_3494,N_3325,N_3278);
xor U3495 (N_3495,N_3282,N_3244);
or U3496 (N_3496,N_3305,N_3208);
nor U3497 (N_3497,N_3322,N_3358);
and U3498 (N_3498,N_3207,N_3333);
nor U3499 (N_3499,N_3345,N_3221);
xnor U3500 (N_3500,N_3324,N_3217);
or U3501 (N_3501,N_3336,N_3221);
or U3502 (N_3502,N_3285,N_3298);
or U3503 (N_3503,N_3224,N_3370);
xnor U3504 (N_3504,N_3287,N_3301);
nor U3505 (N_3505,N_3243,N_3203);
and U3506 (N_3506,N_3206,N_3224);
or U3507 (N_3507,N_3234,N_3286);
and U3508 (N_3508,N_3290,N_3250);
nand U3509 (N_3509,N_3330,N_3309);
nor U3510 (N_3510,N_3384,N_3335);
nand U3511 (N_3511,N_3239,N_3330);
nand U3512 (N_3512,N_3366,N_3203);
and U3513 (N_3513,N_3262,N_3219);
xnor U3514 (N_3514,N_3299,N_3270);
nand U3515 (N_3515,N_3375,N_3352);
xnor U3516 (N_3516,N_3378,N_3368);
and U3517 (N_3517,N_3368,N_3334);
xor U3518 (N_3518,N_3335,N_3333);
nor U3519 (N_3519,N_3335,N_3216);
nor U3520 (N_3520,N_3333,N_3247);
or U3521 (N_3521,N_3322,N_3382);
or U3522 (N_3522,N_3207,N_3254);
nor U3523 (N_3523,N_3372,N_3307);
and U3524 (N_3524,N_3264,N_3351);
nand U3525 (N_3525,N_3271,N_3322);
xnor U3526 (N_3526,N_3330,N_3265);
and U3527 (N_3527,N_3287,N_3385);
or U3528 (N_3528,N_3260,N_3297);
or U3529 (N_3529,N_3250,N_3255);
xor U3530 (N_3530,N_3350,N_3205);
xor U3531 (N_3531,N_3220,N_3346);
nand U3532 (N_3532,N_3221,N_3378);
xor U3533 (N_3533,N_3202,N_3398);
nor U3534 (N_3534,N_3325,N_3255);
and U3535 (N_3535,N_3312,N_3314);
nand U3536 (N_3536,N_3208,N_3219);
and U3537 (N_3537,N_3398,N_3219);
or U3538 (N_3538,N_3255,N_3245);
nand U3539 (N_3539,N_3250,N_3218);
nand U3540 (N_3540,N_3227,N_3233);
nand U3541 (N_3541,N_3215,N_3335);
xnor U3542 (N_3542,N_3269,N_3253);
and U3543 (N_3543,N_3256,N_3362);
nor U3544 (N_3544,N_3369,N_3223);
nand U3545 (N_3545,N_3280,N_3301);
or U3546 (N_3546,N_3335,N_3259);
nor U3547 (N_3547,N_3287,N_3200);
nor U3548 (N_3548,N_3276,N_3213);
or U3549 (N_3549,N_3375,N_3226);
nor U3550 (N_3550,N_3221,N_3322);
or U3551 (N_3551,N_3342,N_3273);
nand U3552 (N_3552,N_3396,N_3256);
nand U3553 (N_3553,N_3209,N_3395);
nor U3554 (N_3554,N_3210,N_3222);
nor U3555 (N_3555,N_3240,N_3378);
and U3556 (N_3556,N_3213,N_3374);
xor U3557 (N_3557,N_3284,N_3374);
and U3558 (N_3558,N_3301,N_3385);
and U3559 (N_3559,N_3233,N_3389);
nand U3560 (N_3560,N_3251,N_3395);
nand U3561 (N_3561,N_3264,N_3263);
nor U3562 (N_3562,N_3228,N_3281);
xor U3563 (N_3563,N_3389,N_3332);
or U3564 (N_3564,N_3374,N_3351);
or U3565 (N_3565,N_3244,N_3348);
or U3566 (N_3566,N_3379,N_3378);
and U3567 (N_3567,N_3294,N_3386);
nor U3568 (N_3568,N_3398,N_3320);
or U3569 (N_3569,N_3353,N_3325);
and U3570 (N_3570,N_3396,N_3205);
and U3571 (N_3571,N_3232,N_3285);
nand U3572 (N_3572,N_3386,N_3332);
and U3573 (N_3573,N_3353,N_3288);
and U3574 (N_3574,N_3325,N_3366);
xor U3575 (N_3575,N_3202,N_3285);
nand U3576 (N_3576,N_3263,N_3335);
or U3577 (N_3577,N_3351,N_3271);
nand U3578 (N_3578,N_3262,N_3358);
nand U3579 (N_3579,N_3293,N_3332);
or U3580 (N_3580,N_3273,N_3395);
and U3581 (N_3581,N_3230,N_3276);
nor U3582 (N_3582,N_3353,N_3214);
nor U3583 (N_3583,N_3244,N_3219);
and U3584 (N_3584,N_3222,N_3214);
xnor U3585 (N_3585,N_3340,N_3394);
nor U3586 (N_3586,N_3398,N_3282);
nand U3587 (N_3587,N_3310,N_3204);
or U3588 (N_3588,N_3251,N_3268);
and U3589 (N_3589,N_3361,N_3230);
and U3590 (N_3590,N_3349,N_3375);
nor U3591 (N_3591,N_3235,N_3290);
nor U3592 (N_3592,N_3297,N_3316);
nand U3593 (N_3593,N_3252,N_3294);
xor U3594 (N_3594,N_3265,N_3299);
xor U3595 (N_3595,N_3394,N_3223);
and U3596 (N_3596,N_3244,N_3232);
or U3597 (N_3597,N_3207,N_3311);
nor U3598 (N_3598,N_3375,N_3247);
nor U3599 (N_3599,N_3277,N_3286);
and U3600 (N_3600,N_3527,N_3481);
and U3601 (N_3601,N_3496,N_3442);
or U3602 (N_3602,N_3456,N_3466);
xnor U3603 (N_3603,N_3507,N_3416);
or U3604 (N_3604,N_3433,N_3404);
and U3605 (N_3605,N_3434,N_3516);
xnor U3606 (N_3606,N_3440,N_3444);
and U3607 (N_3607,N_3423,N_3502);
xor U3608 (N_3608,N_3537,N_3427);
nor U3609 (N_3609,N_3504,N_3483);
and U3610 (N_3610,N_3556,N_3555);
xor U3611 (N_3611,N_3493,N_3551);
nor U3612 (N_3612,N_3531,N_3468);
nand U3613 (N_3613,N_3492,N_3574);
nand U3614 (N_3614,N_3413,N_3569);
or U3615 (N_3615,N_3443,N_3584);
xor U3616 (N_3616,N_3534,N_3491);
xor U3617 (N_3617,N_3418,N_3535);
xor U3618 (N_3618,N_3591,N_3463);
nor U3619 (N_3619,N_3566,N_3559);
nor U3620 (N_3620,N_3594,N_3562);
and U3621 (N_3621,N_3596,N_3577);
nand U3622 (N_3622,N_3564,N_3500);
nor U3623 (N_3623,N_3477,N_3479);
xnor U3624 (N_3624,N_3494,N_3408);
nand U3625 (N_3625,N_3454,N_3573);
and U3626 (N_3626,N_3542,N_3445);
xor U3627 (N_3627,N_3498,N_3478);
or U3628 (N_3628,N_3536,N_3576);
and U3629 (N_3629,N_3464,N_3452);
xnor U3630 (N_3630,N_3490,N_3460);
or U3631 (N_3631,N_3593,N_3592);
and U3632 (N_3632,N_3582,N_3595);
nand U3633 (N_3633,N_3450,N_3458);
nand U3634 (N_3634,N_3470,N_3550);
xor U3635 (N_3635,N_3401,N_3517);
or U3636 (N_3636,N_3518,N_3563);
or U3637 (N_3637,N_3532,N_3539);
xor U3638 (N_3638,N_3515,N_3422);
nand U3639 (N_3639,N_3484,N_3472);
or U3640 (N_3640,N_3462,N_3590);
and U3641 (N_3641,N_3522,N_3560);
xnor U3642 (N_3642,N_3431,N_3469);
and U3643 (N_3643,N_3449,N_3414);
nor U3644 (N_3644,N_3541,N_3540);
nor U3645 (N_3645,N_3587,N_3424);
or U3646 (N_3646,N_3457,N_3580);
nor U3647 (N_3647,N_3571,N_3448);
xor U3648 (N_3648,N_3529,N_3432);
nand U3649 (N_3649,N_3525,N_3475);
nor U3650 (N_3650,N_3497,N_3524);
xor U3651 (N_3651,N_3411,N_3552);
nor U3652 (N_3652,N_3501,N_3575);
and U3653 (N_3653,N_3488,N_3538);
nand U3654 (N_3654,N_3553,N_3461);
and U3655 (N_3655,N_3505,N_3425);
xnor U3656 (N_3656,N_3568,N_3561);
or U3657 (N_3657,N_3459,N_3447);
nand U3658 (N_3658,N_3597,N_3400);
nand U3659 (N_3659,N_3503,N_3549);
or U3660 (N_3660,N_3495,N_3511);
nor U3661 (N_3661,N_3436,N_3428);
nand U3662 (N_3662,N_3499,N_3429);
xnor U3663 (N_3663,N_3512,N_3545);
xnor U3664 (N_3664,N_3579,N_3514);
and U3665 (N_3665,N_3557,N_3417);
and U3666 (N_3666,N_3485,N_3521);
nand U3667 (N_3667,N_3509,N_3430);
xor U3668 (N_3668,N_3403,N_3510);
nand U3669 (N_3669,N_3438,N_3420);
nand U3670 (N_3670,N_3405,N_3589);
xor U3671 (N_3671,N_3506,N_3528);
nand U3672 (N_3672,N_3544,N_3439);
and U3673 (N_3673,N_3415,N_3547);
nor U3674 (N_3674,N_3426,N_3513);
or U3675 (N_3675,N_3530,N_3533);
or U3676 (N_3676,N_3523,N_3409);
nor U3677 (N_3677,N_3586,N_3419);
nand U3678 (N_3678,N_3519,N_3471);
nand U3679 (N_3679,N_3548,N_3410);
nand U3680 (N_3680,N_3480,N_3402);
nand U3681 (N_3681,N_3543,N_3467);
xor U3682 (N_3682,N_3482,N_3565);
xor U3683 (N_3683,N_3486,N_3583);
xnor U3684 (N_3684,N_3599,N_3508);
xor U3685 (N_3685,N_3406,N_3455);
nand U3686 (N_3686,N_3546,N_3489);
nand U3687 (N_3687,N_3446,N_3451);
nand U3688 (N_3688,N_3585,N_3558);
nand U3689 (N_3689,N_3578,N_3407);
and U3690 (N_3690,N_3476,N_3412);
nor U3691 (N_3691,N_3581,N_3526);
xnor U3692 (N_3692,N_3567,N_3520);
nor U3693 (N_3693,N_3598,N_3453);
or U3694 (N_3694,N_3487,N_3441);
nand U3695 (N_3695,N_3465,N_3474);
nor U3696 (N_3696,N_3572,N_3437);
nand U3697 (N_3697,N_3588,N_3473);
and U3698 (N_3698,N_3554,N_3421);
or U3699 (N_3699,N_3570,N_3435);
or U3700 (N_3700,N_3573,N_3572);
xor U3701 (N_3701,N_3570,N_3477);
or U3702 (N_3702,N_3485,N_3573);
or U3703 (N_3703,N_3586,N_3420);
xnor U3704 (N_3704,N_3596,N_3517);
nand U3705 (N_3705,N_3537,N_3466);
nand U3706 (N_3706,N_3410,N_3415);
xnor U3707 (N_3707,N_3425,N_3460);
nand U3708 (N_3708,N_3481,N_3520);
xnor U3709 (N_3709,N_3523,N_3478);
or U3710 (N_3710,N_3514,N_3478);
nand U3711 (N_3711,N_3458,N_3440);
nor U3712 (N_3712,N_3485,N_3411);
nand U3713 (N_3713,N_3439,N_3599);
nor U3714 (N_3714,N_3539,N_3565);
nor U3715 (N_3715,N_3453,N_3568);
nand U3716 (N_3716,N_3568,N_3571);
or U3717 (N_3717,N_3587,N_3591);
nor U3718 (N_3718,N_3413,N_3587);
or U3719 (N_3719,N_3580,N_3489);
and U3720 (N_3720,N_3457,N_3472);
xor U3721 (N_3721,N_3518,N_3526);
xor U3722 (N_3722,N_3462,N_3416);
and U3723 (N_3723,N_3450,N_3477);
nand U3724 (N_3724,N_3551,N_3403);
xor U3725 (N_3725,N_3478,N_3407);
nand U3726 (N_3726,N_3599,N_3565);
or U3727 (N_3727,N_3549,N_3406);
xor U3728 (N_3728,N_3443,N_3515);
xnor U3729 (N_3729,N_3457,N_3404);
or U3730 (N_3730,N_3569,N_3598);
xor U3731 (N_3731,N_3495,N_3468);
or U3732 (N_3732,N_3425,N_3484);
or U3733 (N_3733,N_3493,N_3420);
or U3734 (N_3734,N_3416,N_3497);
xnor U3735 (N_3735,N_3424,N_3462);
xor U3736 (N_3736,N_3535,N_3598);
and U3737 (N_3737,N_3499,N_3562);
and U3738 (N_3738,N_3409,N_3599);
and U3739 (N_3739,N_3411,N_3570);
or U3740 (N_3740,N_3578,N_3405);
or U3741 (N_3741,N_3412,N_3582);
xnor U3742 (N_3742,N_3490,N_3548);
xnor U3743 (N_3743,N_3462,N_3478);
or U3744 (N_3744,N_3501,N_3531);
nand U3745 (N_3745,N_3432,N_3475);
nor U3746 (N_3746,N_3453,N_3406);
nor U3747 (N_3747,N_3470,N_3497);
or U3748 (N_3748,N_3438,N_3433);
and U3749 (N_3749,N_3566,N_3470);
or U3750 (N_3750,N_3417,N_3530);
xnor U3751 (N_3751,N_3574,N_3446);
or U3752 (N_3752,N_3424,N_3571);
or U3753 (N_3753,N_3474,N_3418);
or U3754 (N_3754,N_3595,N_3461);
and U3755 (N_3755,N_3560,N_3466);
nor U3756 (N_3756,N_3587,N_3464);
or U3757 (N_3757,N_3519,N_3555);
and U3758 (N_3758,N_3467,N_3548);
xnor U3759 (N_3759,N_3507,N_3536);
nand U3760 (N_3760,N_3420,N_3578);
or U3761 (N_3761,N_3488,N_3506);
nand U3762 (N_3762,N_3486,N_3522);
nand U3763 (N_3763,N_3415,N_3455);
and U3764 (N_3764,N_3416,N_3505);
or U3765 (N_3765,N_3555,N_3509);
or U3766 (N_3766,N_3535,N_3568);
or U3767 (N_3767,N_3449,N_3497);
nand U3768 (N_3768,N_3408,N_3597);
xnor U3769 (N_3769,N_3478,N_3559);
nand U3770 (N_3770,N_3586,N_3580);
nand U3771 (N_3771,N_3591,N_3540);
nand U3772 (N_3772,N_3431,N_3502);
and U3773 (N_3773,N_3527,N_3580);
and U3774 (N_3774,N_3464,N_3541);
nor U3775 (N_3775,N_3480,N_3440);
and U3776 (N_3776,N_3407,N_3539);
and U3777 (N_3777,N_3447,N_3427);
nor U3778 (N_3778,N_3578,N_3468);
or U3779 (N_3779,N_3410,N_3509);
and U3780 (N_3780,N_3458,N_3513);
xnor U3781 (N_3781,N_3584,N_3421);
xnor U3782 (N_3782,N_3407,N_3401);
xnor U3783 (N_3783,N_3464,N_3479);
or U3784 (N_3784,N_3460,N_3427);
nand U3785 (N_3785,N_3464,N_3429);
or U3786 (N_3786,N_3418,N_3597);
xor U3787 (N_3787,N_3572,N_3485);
nand U3788 (N_3788,N_3568,N_3410);
or U3789 (N_3789,N_3470,N_3448);
xnor U3790 (N_3790,N_3440,N_3408);
or U3791 (N_3791,N_3419,N_3559);
xor U3792 (N_3792,N_3555,N_3508);
xnor U3793 (N_3793,N_3539,N_3537);
xor U3794 (N_3794,N_3586,N_3593);
xor U3795 (N_3795,N_3419,N_3551);
and U3796 (N_3796,N_3567,N_3422);
or U3797 (N_3797,N_3486,N_3410);
nor U3798 (N_3798,N_3417,N_3501);
or U3799 (N_3799,N_3491,N_3500);
nor U3800 (N_3800,N_3624,N_3648);
or U3801 (N_3801,N_3726,N_3760);
or U3802 (N_3802,N_3784,N_3757);
nand U3803 (N_3803,N_3708,N_3636);
or U3804 (N_3804,N_3650,N_3663);
nand U3805 (N_3805,N_3627,N_3783);
nor U3806 (N_3806,N_3697,N_3681);
or U3807 (N_3807,N_3647,N_3785);
nand U3808 (N_3808,N_3696,N_3670);
xnor U3809 (N_3809,N_3637,N_3664);
or U3810 (N_3810,N_3680,N_3679);
nand U3811 (N_3811,N_3691,N_3619);
xnor U3812 (N_3812,N_3676,N_3613);
nand U3813 (N_3813,N_3787,N_3751);
or U3814 (N_3814,N_3622,N_3793);
xor U3815 (N_3815,N_3626,N_3700);
nor U3816 (N_3816,N_3705,N_3629);
or U3817 (N_3817,N_3771,N_3738);
and U3818 (N_3818,N_3749,N_3702);
nand U3819 (N_3819,N_3639,N_3645);
or U3820 (N_3820,N_3661,N_3605);
nand U3821 (N_3821,N_3699,N_3657);
xor U3822 (N_3822,N_3735,N_3740);
nand U3823 (N_3823,N_3786,N_3745);
xor U3824 (N_3824,N_3668,N_3736);
nand U3825 (N_3825,N_3776,N_3611);
nand U3826 (N_3826,N_3712,N_3658);
and U3827 (N_3827,N_3640,N_3798);
nand U3828 (N_3828,N_3788,N_3651);
nand U3829 (N_3829,N_3685,N_3616);
nor U3830 (N_3830,N_3672,N_3765);
nand U3831 (N_3831,N_3683,N_3659);
xnor U3832 (N_3832,N_3630,N_3728);
nor U3833 (N_3833,N_3775,N_3709);
and U3834 (N_3834,N_3742,N_3752);
nand U3835 (N_3835,N_3673,N_3772);
nor U3836 (N_3836,N_3759,N_3649);
xor U3837 (N_3837,N_3719,N_3695);
nand U3838 (N_3838,N_3612,N_3628);
xnor U3839 (N_3839,N_3754,N_3755);
and U3840 (N_3840,N_3758,N_3790);
and U3841 (N_3841,N_3753,N_3703);
nor U3842 (N_3842,N_3782,N_3618);
and U3843 (N_3843,N_3766,N_3701);
nor U3844 (N_3844,N_3761,N_3731);
xor U3845 (N_3845,N_3644,N_3737);
nor U3846 (N_3846,N_3791,N_3666);
or U3847 (N_3847,N_3780,N_3756);
or U3848 (N_3848,N_3656,N_3667);
xnor U3849 (N_3849,N_3698,N_3723);
and U3850 (N_3850,N_3646,N_3714);
nor U3851 (N_3851,N_3643,N_3686);
or U3852 (N_3852,N_3795,N_3693);
nor U3853 (N_3853,N_3721,N_3704);
xnor U3854 (N_3854,N_3778,N_3621);
or U3855 (N_3855,N_3732,N_3678);
and U3856 (N_3856,N_3733,N_3660);
nor U3857 (N_3857,N_3654,N_3614);
or U3858 (N_3858,N_3777,N_3770);
nor U3859 (N_3859,N_3750,N_3720);
or U3860 (N_3860,N_3655,N_3781);
nand U3861 (N_3861,N_3615,N_3779);
xor U3862 (N_3862,N_3747,N_3674);
xor U3863 (N_3863,N_3716,N_3687);
xor U3864 (N_3864,N_3609,N_3707);
or U3865 (N_3865,N_3604,N_3665);
xnor U3866 (N_3866,N_3690,N_3662);
nand U3867 (N_3867,N_3796,N_3689);
xor U3868 (N_3868,N_3789,N_3715);
or U3869 (N_3869,N_3684,N_3635);
xor U3870 (N_3870,N_3692,N_3764);
or U3871 (N_3871,N_3724,N_3631);
xor U3872 (N_3872,N_3722,N_3768);
nand U3873 (N_3873,N_3743,N_3706);
nor U3874 (N_3874,N_3677,N_3682);
xnor U3875 (N_3875,N_3797,N_3769);
xor U3876 (N_3876,N_3711,N_3671);
xor U3877 (N_3877,N_3741,N_3610);
nor U3878 (N_3878,N_3675,N_3620);
nor U3879 (N_3879,N_3652,N_3794);
nand U3880 (N_3880,N_3617,N_3792);
xor U3881 (N_3881,N_3727,N_3606);
nor U3882 (N_3882,N_3748,N_3600);
or U3883 (N_3883,N_3762,N_3634);
xor U3884 (N_3884,N_3729,N_3730);
xor U3885 (N_3885,N_3774,N_3718);
nor U3886 (N_3886,N_3746,N_3744);
nor U3887 (N_3887,N_3799,N_3734);
nand U3888 (N_3888,N_3669,N_3763);
and U3889 (N_3889,N_3625,N_3739);
and U3890 (N_3890,N_3688,N_3694);
or U3891 (N_3891,N_3713,N_3633);
or U3892 (N_3892,N_3632,N_3623);
nand U3893 (N_3893,N_3717,N_3642);
nor U3894 (N_3894,N_3607,N_3725);
nand U3895 (N_3895,N_3773,N_3641);
and U3896 (N_3896,N_3653,N_3603);
or U3897 (N_3897,N_3602,N_3767);
or U3898 (N_3898,N_3638,N_3710);
nor U3899 (N_3899,N_3601,N_3608);
xnor U3900 (N_3900,N_3750,N_3712);
xor U3901 (N_3901,N_3716,N_3711);
xnor U3902 (N_3902,N_3760,N_3722);
or U3903 (N_3903,N_3661,N_3639);
nor U3904 (N_3904,N_3744,N_3741);
nand U3905 (N_3905,N_3703,N_3621);
xnor U3906 (N_3906,N_3691,N_3700);
nand U3907 (N_3907,N_3759,N_3674);
nand U3908 (N_3908,N_3681,N_3665);
nor U3909 (N_3909,N_3634,N_3700);
nor U3910 (N_3910,N_3731,N_3716);
nor U3911 (N_3911,N_3667,N_3699);
nand U3912 (N_3912,N_3759,N_3680);
or U3913 (N_3913,N_3753,N_3623);
xor U3914 (N_3914,N_3769,N_3664);
nand U3915 (N_3915,N_3651,N_3758);
nand U3916 (N_3916,N_3727,N_3761);
or U3917 (N_3917,N_3756,N_3647);
nand U3918 (N_3918,N_3609,N_3694);
nand U3919 (N_3919,N_3608,N_3602);
and U3920 (N_3920,N_3651,N_3786);
xnor U3921 (N_3921,N_3714,N_3689);
or U3922 (N_3922,N_3764,N_3702);
xor U3923 (N_3923,N_3767,N_3665);
nand U3924 (N_3924,N_3749,N_3616);
nand U3925 (N_3925,N_3748,N_3632);
xnor U3926 (N_3926,N_3630,N_3645);
nand U3927 (N_3927,N_3774,N_3690);
and U3928 (N_3928,N_3610,N_3759);
nand U3929 (N_3929,N_3717,N_3627);
nand U3930 (N_3930,N_3654,N_3730);
nor U3931 (N_3931,N_3663,N_3617);
and U3932 (N_3932,N_3766,N_3744);
or U3933 (N_3933,N_3709,N_3611);
xnor U3934 (N_3934,N_3794,N_3619);
and U3935 (N_3935,N_3679,N_3601);
and U3936 (N_3936,N_3785,N_3727);
and U3937 (N_3937,N_3701,N_3726);
or U3938 (N_3938,N_3763,N_3799);
or U3939 (N_3939,N_3788,N_3748);
xnor U3940 (N_3940,N_3779,N_3771);
nand U3941 (N_3941,N_3692,N_3695);
nor U3942 (N_3942,N_3789,N_3658);
nand U3943 (N_3943,N_3696,N_3761);
nor U3944 (N_3944,N_3618,N_3781);
or U3945 (N_3945,N_3630,N_3654);
nor U3946 (N_3946,N_3695,N_3746);
nor U3947 (N_3947,N_3768,N_3744);
or U3948 (N_3948,N_3780,N_3750);
and U3949 (N_3949,N_3628,N_3620);
and U3950 (N_3950,N_3757,N_3781);
or U3951 (N_3951,N_3644,N_3659);
nor U3952 (N_3952,N_3625,N_3659);
xor U3953 (N_3953,N_3697,N_3638);
nor U3954 (N_3954,N_3681,N_3656);
nand U3955 (N_3955,N_3672,N_3710);
xor U3956 (N_3956,N_3641,N_3697);
and U3957 (N_3957,N_3719,N_3623);
nor U3958 (N_3958,N_3686,N_3655);
and U3959 (N_3959,N_3602,N_3675);
nor U3960 (N_3960,N_3793,N_3630);
and U3961 (N_3961,N_3667,N_3706);
or U3962 (N_3962,N_3659,N_3664);
xor U3963 (N_3963,N_3672,N_3616);
and U3964 (N_3964,N_3757,N_3674);
nor U3965 (N_3965,N_3620,N_3692);
nor U3966 (N_3966,N_3772,N_3788);
and U3967 (N_3967,N_3630,N_3705);
and U3968 (N_3968,N_3602,N_3770);
xor U3969 (N_3969,N_3693,N_3672);
xnor U3970 (N_3970,N_3784,N_3622);
xor U3971 (N_3971,N_3795,N_3785);
nand U3972 (N_3972,N_3685,N_3702);
xor U3973 (N_3973,N_3646,N_3738);
nand U3974 (N_3974,N_3636,N_3613);
xnor U3975 (N_3975,N_3712,N_3752);
xor U3976 (N_3976,N_3619,N_3604);
nand U3977 (N_3977,N_3680,N_3640);
nor U3978 (N_3978,N_3790,N_3626);
nand U3979 (N_3979,N_3663,N_3735);
and U3980 (N_3980,N_3768,N_3618);
nor U3981 (N_3981,N_3716,N_3697);
and U3982 (N_3982,N_3779,N_3616);
nor U3983 (N_3983,N_3698,N_3732);
nor U3984 (N_3984,N_3715,N_3744);
nor U3985 (N_3985,N_3660,N_3617);
nor U3986 (N_3986,N_3651,N_3682);
xnor U3987 (N_3987,N_3728,N_3611);
nor U3988 (N_3988,N_3664,N_3728);
and U3989 (N_3989,N_3741,N_3679);
or U3990 (N_3990,N_3688,N_3683);
and U3991 (N_3991,N_3767,N_3738);
xor U3992 (N_3992,N_3698,N_3615);
xor U3993 (N_3993,N_3645,N_3773);
and U3994 (N_3994,N_3725,N_3629);
or U3995 (N_3995,N_3757,N_3742);
nor U3996 (N_3996,N_3615,N_3659);
or U3997 (N_3997,N_3689,N_3669);
and U3998 (N_3998,N_3635,N_3794);
xnor U3999 (N_3999,N_3711,N_3793);
and U4000 (N_4000,N_3866,N_3997);
nand U4001 (N_4001,N_3990,N_3966);
nand U4002 (N_4002,N_3905,N_3899);
nand U4003 (N_4003,N_3960,N_3986);
xnor U4004 (N_4004,N_3902,N_3929);
nor U4005 (N_4005,N_3946,N_3947);
xnor U4006 (N_4006,N_3857,N_3871);
xnor U4007 (N_4007,N_3994,N_3979);
nor U4008 (N_4008,N_3992,N_3900);
nor U4009 (N_4009,N_3989,N_3827);
xnor U4010 (N_4010,N_3837,N_3848);
nor U4011 (N_4011,N_3872,N_3865);
xor U4012 (N_4012,N_3800,N_3885);
nor U4013 (N_4013,N_3803,N_3910);
nor U4014 (N_4014,N_3977,N_3843);
or U4015 (N_4015,N_3876,N_3835);
nand U4016 (N_4016,N_3841,N_3808);
and U4017 (N_4017,N_3907,N_3906);
xnor U4018 (N_4018,N_3809,N_3927);
and U4019 (N_4019,N_3955,N_3895);
nand U4020 (N_4020,N_3833,N_3894);
nand U4021 (N_4021,N_3883,N_3951);
and U4022 (N_4022,N_3874,N_3959);
nand U4023 (N_4023,N_3911,N_3957);
xor U4024 (N_4024,N_3903,N_3846);
xor U4025 (N_4025,N_3854,N_3931);
or U4026 (N_4026,N_3944,N_3880);
nand U4027 (N_4027,N_3998,N_3971);
and U4028 (N_4028,N_3982,N_3969);
xor U4029 (N_4029,N_3812,N_3888);
nor U4030 (N_4030,N_3858,N_3856);
xnor U4031 (N_4031,N_3853,N_3873);
nor U4032 (N_4032,N_3805,N_3818);
nor U4033 (N_4033,N_3904,N_3840);
nor U4034 (N_4034,N_3893,N_3834);
xor U4035 (N_4035,N_3807,N_3915);
xor U4036 (N_4036,N_3839,N_3983);
and U4037 (N_4037,N_3922,N_3867);
or U4038 (N_4038,N_3925,N_3822);
xor U4039 (N_4039,N_3829,N_3847);
or U4040 (N_4040,N_3875,N_3806);
xnor U4041 (N_4041,N_3914,N_3917);
and U4042 (N_4042,N_3996,N_3934);
nor U4043 (N_4043,N_3830,N_3926);
nor U4044 (N_4044,N_3889,N_3984);
or U4045 (N_4045,N_3993,N_3988);
xor U4046 (N_4046,N_3862,N_3801);
nand U4047 (N_4047,N_3878,N_3991);
nand U4048 (N_4048,N_3891,N_3956);
and U4049 (N_4049,N_3975,N_3849);
or U4050 (N_4050,N_3826,N_3901);
and U4051 (N_4051,N_3949,N_3831);
nor U4052 (N_4052,N_3981,N_3896);
and U4053 (N_4053,N_3816,N_3933);
xor U4054 (N_4054,N_3963,N_3919);
nor U4055 (N_4055,N_3819,N_3886);
nor U4056 (N_4056,N_3802,N_3921);
nand U4057 (N_4057,N_3924,N_3953);
or U4058 (N_4058,N_3937,N_3908);
nor U4059 (N_4059,N_3887,N_3964);
xnor U4060 (N_4060,N_3870,N_3940);
or U4061 (N_4061,N_3820,N_3973);
nor U4062 (N_4062,N_3823,N_3976);
xnor U4063 (N_4063,N_3980,N_3836);
nor U4064 (N_4064,N_3968,N_3970);
nand U4065 (N_4065,N_3954,N_3923);
xnor U4066 (N_4066,N_3860,N_3952);
nand U4067 (N_4067,N_3811,N_3828);
nor U4068 (N_4068,N_3824,N_3851);
nand U4069 (N_4069,N_3897,N_3882);
and U4070 (N_4070,N_3999,N_3821);
nor U4071 (N_4071,N_3939,N_3909);
xnor U4072 (N_4072,N_3916,N_3961);
nand U4073 (N_4073,N_3863,N_3850);
nand U4074 (N_4074,N_3913,N_3935);
and U4075 (N_4075,N_3918,N_3974);
xor U4076 (N_4076,N_3928,N_3864);
nand U4077 (N_4077,N_3932,N_3879);
nand U4078 (N_4078,N_3890,N_3950);
nor U4079 (N_4079,N_3884,N_3813);
nor U4080 (N_4080,N_3814,N_3972);
or U4081 (N_4081,N_3958,N_3965);
xnor U4082 (N_4082,N_3938,N_3962);
nand U4083 (N_4083,N_3810,N_3985);
nor U4084 (N_4084,N_3898,N_3942);
xor U4085 (N_4085,N_3877,N_3892);
or U4086 (N_4086,N_3804,N_3995);
xnor U4087 (N_4087,N_3869,N_3855);
and U4088 (N_4088,N_3936,N_3912);
or U4089 (N_4089,N_3943,N_3948);
or U4090 (N_4090,N_3817,N_3978);
nor U4091 (N_4091,N_3844,N_3941);
xor U4092 (N_4092,N_3945,N_3842);
nor U4093 (N_4093,N_3881,N_3825);
nor U4094 (N_4094,N_3861,N_3920);
nor U4095 (N_4095,N_3838,N_3832);
nor U4096 (N_4096,N_3930,N_3845);
and U4097 (N_4097,N_3987,N_3868);
nand U4098 (N_4098,N_3852,N_3859);
nand U4099 (N_4099,N_3815,N_3967);
or U4100 (N_4100,N_3879,N_3929);
nor U4101 (N_4101,N_3916,N_3822);
and U4102 (N_4102,N_3994,N_3893);
and U4103 (N_4103,N_3840,N_3896);
or U4104 (N_4104,N_3836,N_3989);
and U4105 (N_4105,N_3847,N_3975);
and U4106 (N_4106,N_3821,N_3939);
or U4107 (N_4107,N_3816,N_3907);
and U4108 (N_4108,N_3849,N_3982);
nor U4109 (N_4109,N_3988,N_3836);
nor U4110 (N_4110,N_3832,N_3822);
nor U4111 (N_4111,N_3947,N_3930);
nand U4112 (N_4112,N_3950,N_3923);
and U4113 (N_4113,N_3980,N_3947);
nor U4114 (N_4114,N_3844,N_3812);
nand U4115 (N_4115,N_3838,N_3851);
xnor U4116 (N_4116,N_3864,N_3909);
xor U4117 (N_4117,N_3998,N_3896);
xnor U4118 (N_4118,N_3932,N_3933);
and U4119 (N_4119,N_3855,N_3992);
and U4120 (N_4120,N_3975,N_3923);
or U4121 (N_4121,N_3873,N_3919);
xnor U4122 (N_4122,N_3875,N_3934);
nand U4123 (N_4123,N_3863,N_3818);
nand U4124 (N_4124,N_3877,N_3986);
and U4125 (N_4125,N_3889,N_3811);
or U4126 (N_4126,N_3946,N_3802);
nand U4127 (N_4127,N_3953,N_3895);
nor U4128 (N_4128,N_3940,N_3960);
nor U4129 (N_4129,N_3931,N_3960);
xnor U4130 (N_4130,N_3912,N_3922);
and U4131 (N_4131,N_3953,N_3862);
nor U4132 (N_4132,N_3854,N_3974);
and U4133 (N_4133,N_3830,N_3879);
and U4134 (N_4134,N_3978,N_3929);
or U4135 (N_4135,N_3819,N_3921);
nand U4136 (N_4136,N_3885,N_3955);
nor U4137 (N_4137,N_3819,N_3956);
and U4138 (N_4138,N_3877,N_3838);
nor U4139 (N_4139,N_3941,N_3981);
and U4140 (N_4140,N_3894,N_3913);
nand U4141 (N_4141,N_3968,N_3967);
nand U4142 (N_4142,N_3820,N_3906);
xnor U4143 (N_4143,N_3956,N_3837);
or U4144 (N_4144,N_3859,N_3911);
and U4145 (N_4145,N_3869,N_3868);
and U4146 (N_4146,N_3832,N_3804);
xnor U4147 (N_4147,N_3961,N_3922);
xnor U4148 (N_4148,N_3954,N_3902);
nand U4149 (N_4149,N_3877,N_3850);
nand U4150 (N_4150,N_3884,N_3851);
or U4151 (N_4151,N_3946,N_3924);
or U4152 (N_4152,N_3949,N_3975);
nor U4153 (N_4153,N_3940,N_3830);
nor U4154 (N_4154,N_3949,N_3920);
and U4155 (N_4155,N_3806,N_3993);
or U4156 (N_4156,N_3950,N_3818);
and U4157 (N_4157,N_3954,N_3977);
nand U4158 (N_4158,N_3824,N_3813);
and U4159 (N_4159,N_3886,N_3983);
and U4160 (N_4160,N_3834,N_3885);
xor U4161 (N_4161,N_3952,N_3825);
or U4162 (N_4162,N_3873,N_3916);
nand U4163 (N_4163,N_3992,N_3831);
xor U4164 (N_4164,N_3958,N_3974);
nand U4165 (N_4165,N_3970,N_3932);
xor U4166 (N_4166,N_3982,N_3872);
nand U4167 (N_4167,N_3876,N_3900);
and U4168 (N_4168,N_3843,N_3936);
nor U4169 (N_4169,N_3954,N_3909);
nand U4170 (N_4170,N_3879,N_3873);
or U4171 (N_4171,N_3992,N_3986);
nand U4172 (N_4172,N_3898,N_3873);
xor U4173 (N_4173,N_3948,N_3814);
xor U4174 (N_4174,N_3998,N_3807);
or U4175 (N_4175,N_3989,N_3998);
nand U4176 (N_4176,N_3945,N_3983);
xnor U4177 (N_4177,N_3986,N_3844);
nand U4178 (N_4178,N_3964,N_3998);
nand U4179 (N_4179,N_3910,N_3811);
or U4180 (N_4180,N_3848,N_3875);
nand U4181 (N_4181,N_3814,N_3838);
nor U4182 (N_4182,N_3915,N_3991);
or U4183 (N_4183,N_3825,N_3842);
or U4184 (N_4184,N_3997,N_3899);
and U4185 (N_4185,N_3930,N_3943);
nand U4186 (N_4186,N_3941,N_3970);
and U4187 (N_4187,N_3905,N_3963);
or U4188 (N_4188,N_3811,N_3805);
nand U4189 (N_4189,N_3805,N_3814);
nand U4190 (N_4190,N_3857,N_3858);
xnor U4191 (N_4191,N_3822,N_3906);
and U4192 (N_4192,N_3800,N_3872);
xor U4193 (N_4193,N_3954,N_3816);
nand U4194 (N_4194,N_3992,N_3803);
and U4195 (N_4195,N_3921,N_3971);
xor U4196 (N_4196,N_3916,N_3867);
xnor U4197 (N_4197,N_3900,N_3890);
nor U4198 (N_4198,N_3847,N_3805);
xor U4199 (N_4199,N_3975,N_3971);
xnor U4200 (N_4200,N_4114,N_4000);
xor U4201 (N_4201,N_4048,N_4068);
and U4202 (N_4202,N_4035,N_4125);
and U4203 (N_4203,N_4132,N_4038);
nand U4204 (N_4204,N_4163,N_4039);
or U4205 (N_4205,N_4115,N_4161);
and U4206 (N_4206,N_4138,N_4084);
or U4207 (N_4207,N_4196,N_4172);
nor U4208 (N_4208,N_4086,N_4144);
xnor U4209 (N_4209,N_4185,N_4102);
xor U4210 (N_4210,N_4120,N_4079);
or U4211 (N_4211,N_4093,N_4131);
and U4212 (N_4212,N_4013,N_4190);
or U4213 (N_4213,N_4165,N_4029);
or U4214 (N_4214,N_4097,N_4117);
or U4215 (N_4215,N_4073,N_4152);
and U4216 (N_4216,N_4014,N_4025);
or U4217 (N_4217,N_4149,N_4123);
nand U4218 (N_4218,N_4150,N_4191);
and U4219 (N_4219,N_4175,N_4006);
nand U4220 (N_4220,N_4101,N_4176);
nand U4221 (N_4221,N_4072,N_4042);
xnor U4222 (N_4222,N_4027,N_4067);
nand U4223 (N_4223,N_4178,N_4021);
and U4224 (N_4224,N_4112,N_4151);
xor U4225 (N_4225,N_4063,N_4140);
nor U4226 (N_4226,N_4045,N_4023);
and U4227 (N_4227,N_4137,N_4103);
and U4228 (N_4228,N_4077,N_4107);
nor U4229 (N_4229,N_4085,N_4181);
or U4230 (N_4230,N_4145,N_4057);
and U4231 (N_4231,N_4080,N_4022);
and U4232 (N_4232,N_4075,N_4130);
nand U4233 (N_4233,N_4094,N_4100);
and U4234 (N_4234,N_4003,N_4174);
or U4235 (N_4235,N_4009,N_4139);
and U4236 (N_4236,N_4011,N_4189);
and U4237 (N_4237,N_4054,N_4106);
nand U4238 (N_4238,N_4058,N_4168);
and U4239 (N_4239,N_4089,N_4095);
nand U4240 (N_4240,N_4083,N_4171);
nor U4241 (N_4241,N_4160,N_4078);
and U4242 (N_4242,N_4017,N_4076);
nor U4243 (N_4243,N_4064,N_4096);
nand U4244 (N_4244,N_4199,N_4026);
and U4245 (N_4245,N_4030,N_4002);
or U4246 (N_4246,N_4135,N_4183);
and U4247 (N_4247,N_4142,N_4055);
or U4248 (N_4248,N_4105,N_4173);
or U4249 (N_4249,N_4194,N_4056);
nor U4250 (N_4250,N_4012,N_4060);
xor U4251 (N_4251,N_4001,N_4005);
xor U4252 (N_4252,N_4179,N_4157);
nand U4253 (N_4253,N_4069,N_4071);
xnor U4254 (N_4254,N_4113,N_4154);
nand U4255 (N_4255,N_4156,N_4052);
nand U4256 (N_4256,N_4197,N_4153);
and U4257 (N_4257,N_4122,N_4040);
or U4258 (N_4258,N_4164,N_4099);
xor U4259 (N_4259,N_4195,N_4050);
xnor U4260 (N_4260,N_4193,N_4186);
or U4261 (N_4261,N_4159,N_4169);
nand U4262 (N_4262,N_4010,N_4028);
xnor U4263 (N_4263,N_4133,N_4020);
and U4264 (N_4264,N_4110,N_4129);
nor U4265 (N_4265,N_4004,N_4118);
xnor U4266 (N_4266,N_4043,N_4108);
xor U4267 (N_4267,N_4128,N_4031);
nand U4268 (N_4268,N_4015,N_4034);
and U4269 (N_4269,N_4111,N_4182);
and U4270 (N_4270,N_4074,N_4170);
or U4271 (N_4271,N_4007,N_4016);
or U4272 (N_4272,N_4167,N_4090);
nor U4273 (N_4273,N_4036,N_4098);
and U4274 (N_4274,N_4059,N_4126);
nand U4275 (N_4275,N_4092,N_4033);
xor U4276 (N_4276,N_4124,N_4192);
xor U4277 (N_4277,N_4177,N_4008);
or U4278 (N_4278,N_4070,N_4061);
nor U4279 (N_4279,N_4116,N_4155);
and U4280 (N_4280,N_4032,N_4104);
nor U4281 (N_4281,N_4162,N_4081);
nand U4282 (N_4282,N_4018,N_4082);
nor U4283 (N_4283,N_4134,N_4166);
and U4284 (N_4284,N_4180,N_4119);
and U4285 (N_4285,N_4066,N_4062);
xnor U4286 (N_4286,N_4148,N_4091);
xor U4287 (N_4287,N_4147,N_4127);
nand U4288 (N_4288,N_4141,N_4047);
or U4289 (N_4289,N_4146,N_4051);
nor U4290 (N_4290,N_4136,N_4053);
xor U4291 (N_4291,N_4019,N_4121);
xnor U4292 (N_4292,N_4087,N_4158);
nand U4293 (N_4293,N_4109,N_4188);
xor U4294 (N_4294,N_4143,N_4198);
and U4295 (N_4295,N_4024,N_4049);
nor U4296 (N_4296,N_4065,N_4187);
xnor U4297 (N_4297,N_4184,N_4088);
xor U4298 (N_4298,N_4044,N_4037);
and U4299 (N_4299,N_4041,N_4046);
and U4300 (N_4300,N_4010,N_4125);
nor U4301 (N_4301,N_4000,N_4029);
nor U4302 (N_4302,N_4184,N_4141);
or U4303 (N_4303,N_4140,N_4159);
xnor U4304 (N_4304,N_4193,N_4189);
or U4305 (N_4305,N_4149,N_4155);
nor U4306 (N_4306,N_4090,N_4061);
xor U4307 (N_4307,N_4081,N_4123);
nor U4308 (N_4308,N_4074,N_4175);
xor U4309 (N_4309,N_4068,N_4020);
and U4310 (N_4310,N_4070,N_4091);
and U4311 (N_4311,N_4197,N_4170);
and U4312 (N_4312,N_4165,N_4080);
nand U4313 (N_4313,N_4059,N_4027);
or U4314 (N_4314,N_4136,N_4062);
xor U4315 (N_4315,N_4196,N_4056);
or U4316 (N_4316,N_4097,N_4066);
nor U4317 (N_4317,N_4195,N_4175);
nand U4318 (N_4318,N_4106,N_4176);
nor U4319 (N_4319,N_4198,N_4197);
and U4320 (N_4320,N_4145,N_4193);
nor U4321 (N_4321,N_4073,N_4008);
and U4322 (N_4322,N_4074,N_4094);
and U4323 (N_4323,N_4185,N_4030);
and U4324 (N_4324,N_4111,N_4079);
xnor U4325 (N_4325,N_4127,N_4135);
xor U4326 (N_4326,N_4133,N_4119);
nor U4327 (N_4327,N_4142,N_4180);
and U4328 (N_4328,N_4003,N_4112);
nor U4329 (N_4329,N_4170,N_4019);
nand U4330 (N_4330,N_4122,N_4070);
and U4331 (N_4331,N_4133,N_4141);
xor U4332 (N_4332,N_4067,N_4018);
nor U4333 (N_4333,N_4073,N_4103);
nand U4334 (N_4334,N_4142,N_4050);
or U4335 (N_4335,N_4156,N_4151);
nor U4336 (N_4336,N_4007,N_4147);
nor U4337 (N_4337,N_4056,N_4052);
xnor U4338 (N_4338,N_4075,N_4000);
nor U4339 (N_4339,N_4065,N_4001);
or U4340 (N_4340,N_4058,N_4143);
nand U4341 (N_4341,N_4181,N_4099);
nand U4342 (N_4342,N_4090,N_4139);
nor U4343 (N_4343,N_4017,N_4022);
or U4344 (N_4344,N_4141,N_4050);
xor U4345 (N_4345,N_4041,N_4035);
or U4346 (N_4346,N_4115,N_4031);
nand U4347 (N_4347,N_4103,N_4163);
or U4348 (N_4348,N_4147,N_4119);
or U4349 (N_4349,N_4164,N_4187);
or U4350 (N_4350,N_4185,N_4004);
or U4351 (N_4351,N_4106,N_4047);
and U4352 (N_4352,N_4021,N_4074);
xor U4353 (N_4353,N_4175,N_4120);
nand U4354 (N_4354,N_4198,N_4005);
nor U4355 (N_4355,N_4058,N_4173);
or U4356 (N_4356,N_4010,N_4181);
and U4357 (N_4357,N_4136,N_4095);
nand U4358 (N_4358,N_4196,N_4087);
nand U4359 (N_4359,N_4065,N_4064);
nand U4360 (N_4360,N_4150,N_4115);
xor U4361 (N_4361,N_4113,N_4079);
xor U4362 (N_4362,N_4009,N_4140);
xnor U4363 (N_4363,N_4179,N_4025);
and U4364 (N_4364,N_4020,N_4042);
nand U4365 (N_4365,N_4010,N_4087);
nor U4366 (N_4366,N_4079,N_4075);
and U4367 (N_4367,N_4067,N_4076);
and U4368 (N_4368,N_4154,N_4083);
xor U4369 (N_4369,N_4017,N_4161);
xor U4370 (N_4370,N_4196,N_4052);
and U4371 (N_4371,N_4062,N_4003);
nor U4372 (N_4372,N_4091,N_4087);
nand U4373 (N_4373,N_4093,N_4195);
xor U4374 (N_4374,N_4182,N_4029);
or U4375 (N_4375,N_4057,N_4149);
or U4376 (N_4376,N_4129,N_4199);
nor U4377 (N_4377,N_4130,N_4154);
xnor U4378 (N_4378,N_4150,N_4185);
nand U4379 (N_4379,N_4100,N_4190);
and U4380 (N_4380,N_4146,N_4088);
or U4381 (N_4381,N_4186,N_4056);
nand U4382 (N_4382,N_4012,N_4049);
xnor U4383 (N_4383,N_4128,N_4071);
and U4384 (N_4384,N_4036,N_4011);
xnor U4385 (N_4385,N_4005,N_4098);
xnor U4386 (N_4386,N_4193,N_4039);
nor U4387 (N_4387,N_4185,N_4083);
nor U4388 (N_4388,N_4189,N_4034);
or U4389 (N_4389,N_4070,N_4198);
nand U4390 (N_4390,N_4008,N_4087);
nor U4391 (N_4391,N_4188,N_4091);
and U4392 (N_4392,N_4046,N_4195);
or U4393 (N_4393,N_4175,N_4078);
and U4394 (N_4394,N_4048,N_4096);
nor U4395 (N_4395,N_4156,N_4006);
xor U4396 (N_4396,N_4134,N_4154);
or U4397 (N_4397,N_4139,N_4010);
xnor U4398 (N_4398,N_4112,N_4143);
xor U4399 (N_4399,N_4144,N_4083);
nor U4400 (N_4400,N_4361,N_4296);
and U4401 (N_4401,N_4297,N_4219);
nand U4402 (N_4402,N_4278,N_4250);
and U4403 (N_4403,N_4254,N_4249);
nand U4404 (N_4404,N_4318,N_4258);
or U4405 (N_4405,N_4367,N_4263);
and U4406 (N_4406,N_4330,N_4344);
nand U4407 (N_4407,N_4291,N_4280);
and U4408 (N_4408,N_4224,N_4244);
nor U4409 (N_4409,N_4369,N_4204);
or U4410 (N_4410,N_4373,N_4309);
nand U4411 (N_4411,N_4307,N_4283);
nor U4412 (N_4412,N_4279,N_4349);
xnor U4413 (N_4413,N_4354,N_4394);
xnor U4414 (N_4414,N_4228,N_4285);
nor U4415 (N_4415,N_4341,N_4362);
or U4416 (N_4416,N_4357,N_4339);
nor U4417 (N_4417,N_4332,N_4333);
nand U4418 (N_4418,N_4397,N_4276);
xor U4419 (N_4419,N_4268,N_4260);
and U4420 (N_4420,N_4399,N_4310);
nor U4421 (N_4421,N_4311,N_4377);
nand U4422 (N_4422,N_4363,N_4313);
nor U4423 (N_4423,N_4372,N_4221);
and U4424 (N_4424,N_4201,N_4286);
nor U4425 (N_4425,N_4380,N_4240);
nand U4426 (N_4426,N_4247,N_4387);
nand U4427 (N_4427,N_4382,N_4203);
and U4428 (N_4428,N_4323,N_4265);
and U4429 (N_4429,N_4355,N_4384);
or U4430 (N_4430,N_4237,N_4319);
xor U4431 (N_4431,N_4386,N_4337);
nand U4432 (N_4432,N_4383,N_4293);
and U4433 (N_4433,N_4206,N_4329);
nand U4434 (N_4434,N_4395,N_4359);
and U4435 (N_4435,N_4266,N_4336);
nor U4436 (N_4436,N_4366,N_4284);
or U4437 (N_4437,N_4277,N_4379);
xnor U4438 (N_4438,N_4234,N_4300);
and U4439 (N_4439,N_4375,N_4390);
xnor U4440 (N_4440,N_4396,N_4312);
or U4441 (N_4441,N_4338,N_4346);
and U4442 (N_4442,N_4232,N_4289);
and U4443 (N_4443,N_4374,N_4231);
xnor U4444 (N_4444,N_4290,N_4342);
or U4445 (N_4445,N_4385,N_4371);
nand U4446 (N_4446,N_4202,N_4281);
nand U4447 (N_4447,N_4398,N_4327);
nor U4448 (N_4448,N_4245,N_4236);
or U4449 (N_4449,N_4350,N_4218);
and U4450 (N_4450,N_4261,N_4340);
nor U4451 (N_4451,N_4320,N_4217);
nor U4452 (N_4452,N_4360,N_4251);
nand U4453 (N_4453,N_4226,N_4264);
nor U4454 (N_4454,N_4392,N_4267);
or U4455 (N_4455,N_4239,N_4322);
or U4456 (N_4456,N_4314,N_4317);
xor U4457 (N_4457,N_4220,N_4316);
or U4458 (N_4458,N_4256,N_4364);
and U4459 (N_4459,N_4345,N_4315);
xor U4460 (N_4460,N_4262,N_4306);
or U4461 (N_4461,N_4325,N_4351);
nor U4462 (N_4462,N_4370,N_4225);
xnor U4463 (N_4463,N_4272,N_4208);
nand U4464 (N_4464,N_4230,N_4227);
and U4465 (N_4465,N_4275,N_4348);
or U4466 (N_4466,N_4302,N_4381);
nand U4467 (N_4467,N_4305,N_4303);
or U4468 (N_4468,N_4246,N_4238);
or U4469 (N_4469,N_4207,N_4271);
or U4470 (N_4470,N_4298,N_4353);
nor U4471 (N_4471,N_4388,N_4255);
and U4472 (N_4472,N_4343,N_4335);
or U4473 (N_4473,N_4292,N_4321);
nor U4474 (N_4474,N_4269,N_4331);
xor U4475 (N_4475,N_4200,N_4212);
and U4476 (N_4476,N_4259,N_4214);
nand U4477 (N_4477,N_4326,N_4299);
and U4478 (N_4478,N_4213,N_4308);
or U4479 (N_4479,N_4241,N_4274);
nand U4480 (N_4480,N_4282,N_4235);
nor U4481 (N_4481,N_4242,N_4270);
xor U4482 (N_4482,N_4301,N_4287);
xnor U4483 (N_4483,N_4347,N_4295);
or U4484 (N_4484,N_4273,N_4328);
xor U4485 (N_4485,N_4222,N_4365);
nand U4486 (N_4486,N_4378,N_4352);
and U4487 (N_4487,N_4210,N_4376);
xnor U4488 (N_4488,N_4243,N_4393);
nor U4489 (N_4489,N_4334,N_4391);
nor U4490 (N_4490,N_4288,N_4253);
or U4491 (N_4491,N_4233,N_4205);
nand U4492 (N_4492,N_4389,N_4229);
and U4493 (N_4493,N_4223,N_4211);
or U4494 (N_4494,N_4216,N_4257);
nand U4495 (N_4495,N_4294,N_4358);
nand U4496 (N_4496,N_4368,N_4209);
nor U4497 (N_4497,N_4356,N_4304);
nand U4498 (N_4498,N_4324,N_4252);
or U4499 (N_4499,N_4215,N_4248);
and U4500 (N_4500,N_4215,N_4242);
or U4501 (N_4501,N_4298,N_4337);
nand U4502 (N_4502,N_4305,N_4357);
xnor U4503 (N_4503,N_4241,N_4212);
and U4504 (N_4504,N_4312,N_4210);
xor U4505 (N_4505,N_4215,N_4237);
nor U4506 (N_4506,N_4353,N_4280);
and U4507 (N_4507,N_4278,N_4217);
xnor U4508 (N_4508,N_4204,N_4257);
xnor U4509 (N_4509,N_4206,N_4294);
and U4510 (N_4510,N_4363,N_4272);
or U4511 (N_4511,N_4247,N_4226);
or U4512 (N_4512,N_4221,N_4362);
and U4513 (N_4513,N_4321,N_4226);
nand U4514 (N_4514,N_4349,N_4381);
or U4515 (N_4515,N_4288,N_4313);
nand U4516 (N_4516,N_4288,N_4334);
nand U4517 (N_4517,N_4200,N_4249);
nor U4518 (N_4518,N_4329,N_4211);
and U4519 (N_4519,N_4300,N_4243);
nand U4520 (N_4520,N_4227,N_4317);
and U4521 (N_4521,N_4200,N_4396);
nand U4522 (N_4522,N_4300,N_4399);
and U4523 (N_4523,N_4306,N_4360);
or U4524 (N_4524,N_4326,N_4215);
xnor U4525 (N_4525,N_4277,N_4278);
and U4526 (N_4526,N_4205,N_4317);
and U4527 (N_4527,N_4286,N_4326);
nor U4528 (N_4528,N_4368,N_4363);
and U4529 (N_4529,N_4207,N_4203);
or U4530 (N_4530,N_4379,N_4398);
xnor U4531 (N_4531,N_4246,N_4208);
nor U4532 (N_4532,N_4371,N_4342);
nand U4533 (N_4533,N_4364,N_4245);
and U4534 (N_4534,N_4300,N_4332);
and U4535 (N_4535,N_4268,N_4290);
nor U4536 (N_4536,N_4267,N_4286);
and U4537 (N_4537,N_4299,N_4353);
and U4538 (N_4538,N_4302,N_4249);
nand U4539 (N_4539,N_4237,N_4228);
nor U4540 (N_4540,N_4261,N_4251);
xor U4541 (N_4541,N_4277,N_4355);
or U4542 (N_4542,N_4225,N_4319);
xnor U4543 (N_4543,N_4302,N_4312);
or U4544 (N_4544,N_4336,N_4215);
or U4545 (N_4545,N_4316,N_4273);
nor U4546 (N_4546,N_4238,N_4213);
and U4547 (N_4547,N_4208,N_4264);
nor U4548 (N_4548,N_4220,N_4378);
xor U4549 (N_4549,N_4374,N_4358);
and U4550 (N_4550,N_4287,N_4205);
or U4551 (N_4551,N_4270,N_4258);
or U4552 (N_4552,N_4287,N_4213);
and U4553 (N_4553,N_4318,N_4207);
or U4554 (N_4554,N_4272,N_4224);
and U4555 (N_4555,N_4375,N_4269);
nand U4556 (N_4556,N_4374,N_4344);
xnor U4557 (N_4557,N_4287,N_4268);
or U4558 (N_4558,N_4385,N_4208);
nand U4559 (N_4559,N_4266,N_4244);
and U4560 (N_4560,N_4381,N_4282);
nand U4561 (N_4561,N_4284,N_4381);
nor U4562 (N_4562,N_4319,N_4299);
nand U4563 (N_4563,N_4261,N_4364);
nand U4564 (N_4564,N_4263,N_4349);
nand U4565 (N_4565,N_4323,N_4340);
nand U4566 (N_4566,N_4209,N_4272);
or U4567 (N_4567,N_4326,N_4272);
nand U4568 (N_4568,N_4225,N_4261);
and U4569 (N_4569,N_4301,N_4364);
and U4570 (N_4570,N_4315,N_4330);
nand U4571 (N_4571,N_4203,N_4230);
or U4572 (N_4572,N_4321,N_4274);
nor U4573 (N_4573,N_4344,N_4296);
and U4574 (N_4574,N_4267,N_4272);
nor U4575 (N_4575,N_4297,N_4298);
and U4576 (N_4576,N_4200,N_4219);
or U4577 (N_4577,N_4393,N_4328);
and U4578 (N_4578,N_4389,N_4320);
nor U4579 (N_4579,N_4303,N_4233);
nor U4580 (N_4580,N_4286,N_4310);
or U4581 (N_4581,N_4273,N_4310);
nand U4582 (N_4582,N_4394,N_4265);
xnor U4583 (N_4583,N_4308,N_4325);
and U4584 (N_4584,N_4279,N_4295);
nor U4585 (N_4585,N_4254,N_4360);
nor U4586 (N_4586,N_4210,N_4320);
and U4587 (N_4587,N_4353,N_4227);
or U4588 (N_4588,N_4358,N_4300);
nand U4589 (N_4589,N_4300,N_4395);
xor U4590 (N_4590,N_4334,N_4370);
or U4591 (N_4591,N_4276,N_4234);
xnor U4592 (N_4592,N_4301,N_4213);
nor U4593 (N_4593,N_4228,N_4267);
nor U4594 (N_4594,N_4261,N_4350);
xnor U4595 (N_4595,N_4269,N_4381);
nand U4596 (N_4596,N_4220,N_4286);
and U4597 (N_4597,N_4297,N_4289);
xnor U4598 (N_4598,N_4395,N_4354);
xor U4599 (N_4599,N_4242,N_4208);
xnor U4600 (N_4600,N_4488,N_4523);
or U4601 (N_4601,N_4493,N_4466);
and U4602 (N_4602,N_4515,N_4450);
and U4603 (N_4603,N_4563,N_4579);
or U4604 (N_4604,N_4569,N_4418);
nor U4605 (N_4605,N_4492,N_4494);
or U4606 (N_4606,N_4528,N_4419);
xor U4607 (N_4607,N_4541,N_4598);
or U4608 (N_4608,N_4470,N_4473);
xor U4609 (N_4609,N_4547,N_4434);
nand U4610 (N_4610,N_4461,N_4489);
or U4611 (N_4611,N_4420,N_4445);
and U4612 (N_4612,N_4559,N_4487);
and U4613 (N_4613,N_4520,N_4503);
nor U4614 (N_4614,N_4463,N_4527);
xnor U4615 (N_4615,N_4453,N_4562);
and U4616 (N_4616,N_4584,N_4435);
nor U4617 (N_4617,N_4480,N_4412);
nor U4618 (N_4618,N_4431,N_4406);
or U4619 (N_4619,N_4537,N_4501);
nand U4620 (N_4620,N_4572,N_4530);
or U4621 (N_4621,N_4560,N_4575);
or U4622 (N_4622,N_4585,N_4400);
nor U4623 (N_4623,N_4554,N_4482);
or U4624 (N_4624,N_4401,N_4405);
nor U4625 (N_4625,N_4533,N_4427);
xor U4626 (N_4626,N_4573,N_4452);
nand U4627 (N_4627,N_4446,N_4404);
nand U4628 (N_4628,N_4467,N_4556);
or U4629 (N_4629,N_4459,N_4447);
or U4630 (N_4630,N_4415,N_4521);
xnor U4631 (N_4631,N_4490,N_4464);
xor U4632 (N_4632,N_4544,N_4444);
nand U4633 (N_4633,N_4529,N_4505);
nor U4634 (N_4634,N_4589,N_4430);
nor U4635 (N_4635,N_4451,N_4506);
nand U4636 (N_4636,N_4582,N_4524);
nor U4637 (N_4637,N_4586,N_4549);
or U4638 (N_4638,N_4477,N_4468);
xnor U4639 (N_4639,N_4491,N_4518);
nor U4640 (N_4640,N_4571,N_4496);
nand U4641 (N_4641,N_4593,N_4597);
nand U4642 (N_4642,N_4499,N_4535);
xor U4643 (N_4643,N_4546,N_4476);
or U4644 (N_4644,N_4539,N_4436);
nor U4645 (N_4645,N_4587,N_4526);
nor U4646 (N_4646,N_4484,N_4510);
and U4647 (N_4647,N_4507,N_4411);
or U4648 (N_4648,N_4532,N_4580);
xor U4649 (N_4649,N_4407,N_4522);
xor U4650 (N_4650,N_4458,N_4566);
and U4651 (N_4651,N_4410,N_4551);
nand U4652 (N_4652,N_4429,N_4567);
or U4653 (N_4653,N_4416,N_4591);
xnor U4654 (N_4654,N_4497,N_4481);
and U4655 (N_4655,N_4495,N_4565);
xor U4656 (N_4656,N_4592,N_4465);
nand U4657 (N_4657,N_4456,N_4574);
nor U4658 (N_4658,N_4460,N_4514);
and U4659 (N_4659,N_4536,N_4543);
or U4660 (N_4660,N_4564,N_4432);
and U4661 (N_4661,N_4408,N_4561);
and U4662 (N_4662,N_4545,N_4448);
xnor U4663 (N_4663,N_4454,N_4421);
or U4664 (N_4664,N_4553,N_4511);
and U4665 (N_4665,N_4439,N_4517);
or U4666 (N_4666,N_4462,N_4540);
xnor U4667 (N_4667,N_4504,N_4590);
nor U4668 (N_4668,N_4525,N_4440);
nand U4669 (N_4669,N_4512,N_4438);
xnor U4670 (N_4670,N_4548,N_4478);
xor U4671 (N_4671,N_4469,N_4449);
and U4672 (N_4672,N_4509,N_4542);
xor U4673 (N_4673,N_4581,N_4403);
nand U4674 (N_4674,N_4513,N_4576);
nand U4675 (N_4675,N_4486,N_4538);
nor U4676 (N_4676,N_4516,N_4502);
xor U4677 (N_4677,N_4425,N_4588);
xnor U4678 (N_4678,N_4485,N_4474);
or U4679 (N_4679,N_4578,N_4471);
and U4680 (N_4680,N_4409,N_4552);
nand U4681 (N_4681,N_4500,N_4426);
nand U4682 (N_4682,N_4433,N_4422);
xor U4683 (N_4683,N_4595,N_4417);
nor U4684 (N_4684,N_4596,N_4402);
or U4685 (N_4685,N_4443,N_4498);
or U4686 (N_4686,N_4568,N_4531);
or U4687 (N_4687,N_4442,N_4413);
or U4688 (N_4688,N_4558,N_4550);
and U4689 (N_4689,N_4441,N_4534);
nor U4690 (N_4690,N_4594,N_4423);
xnor U4691 (N_4691,N_4555,N_4414);
nand U4692 (N_4692,N_4519,N_4424);
or U4693 (N_4693,N_4508,N_4457);
nor U4694 (N_4694,N_4570,N_4483);
or U4695 (N_4695,N_4479,N_4472);
or U4696 (N_4696,N_4557,N_4455);
nand U4697 (N_4697,N_4437,N_4583);
and U4698 (N_4698,N_4428,N_4475);
nor U4699 (N_4699,N_4577,N_4599);
and U4700 (N_4700,N_4457,N_4521);
nor U4701 (N_4701,N_4522,N_4519);
nand U4702 (N_4702,N_4504,N_4521);
and U4703 (N_4703,N_4538,N_4520);
xnor U4704 (N_4704,N_4447,N_4497);
nor U4705 (N_4705,N_4586,N_4587);
xor U4706 (N_4706,N_4597,N_4415);
and U4707 (N_4707,N_4543,N_4508);
nand U4708 (N_4708,N_4582,N_4409);
nor U4709 (N_4709,N_4518,N_4576);
and U4710 (N_4710,N_4553,N_4441);
xnor U4711 (N_4711,N_4594,N_4509);
or U4712 (N_4712,N_4571,N_4514);
and U4713 (N_4713,N_4508,N_4548);
and U4714 (N_4714,N_4596,N_4560);
xor U4715 (N_4715,N_4475,N_4599);
nand U4716 (N_4716,N_4511,N_4598);
xnor U4717 (N_4717,N_4534,N_4580);
nand U4718 (N_4718,N_4420,N_4504);
and U4719 (N_4719,N_4415,N_4430);
or U4720 (N_4720,N_4450,N_4500);
or U4721 (N_4721,N_4577,N_4444);
and U4722 (N_4722,N_4441,N_4455);
and U4723 (N_4723,N_4475,N_4477);
nand U4724 (N_4724,N_4503,N_4458);
or U4725 (N_4725,N_4596,N_4493);
nor U4726 (N_4726,N_4560,N_4402);
nor U4727 (N_4727,N_4509,N_4520);
xor U4728 (N_4728,N_4479,N_4561);
nand U4729 (N_4729,N_4419,N_4405);
and U4730 (N_4730,N_4579,N_4445);
or U4731 (N_4731,N_4586,N_4439);
nand U4732 (N_4732,N_4444,N_4471);
and U4733 (N_4733,N_4427,N_4412);
and U4734 (N_4734,N_4441,N_4540);
nand U4735 (N_4735,N_4402,N_4540);
or U4736 (N_4736,N_4469,N_4490);
nor U4737 (N_4737,N_4423,N_4448);
or U4738 (N_4738,N_4482,N_4425);
nor U4739 (N_4739,N_4510,N_4553);
nor U4740 (N_4740,N_4497,N_4598);
xnor U4741 (N_4741,N_4423,N_4408);
xor U4742 (N_4742,N_4403,N_4543);
nand U4743 (N_4743,N_4465,N_4558);
xor U4744 (N_4744,N_4431,N_4502);
or U4745 (N_4745,N_4532,N_4414);
nand U4746 (N_4746,N_4563,N_4524);
xor U4747 (N_4747,N_4524,N_4445);
nand U4748 (N_4748,N_4458,N_4516);
xor U4749 (N_4749,N_4597,N_4499);
and U4750 (N_4750,N_4487,N_4446);
nor U4751 (N_4751,N_4418,N_4562);
nor U4752 (N_4752,N_4468,N_4546);
or U4753 (N_4753,N_4511,N_4452);
and U4754 (N_4754,N_4540,N_4452);
or U4755 (N_4755,N_4591,N_4493);
and U4756 (N_4756,N_4586,N_4501);
nand U4757 (N_4757,N_4437,N_4489);
or U4758 (N_4758,N_4586,N_4418);
xnor U4759 (N_4759,N_4535,N_4409);
or U4760 (N_4760,N_4459,N_4418);
and U4761 (N_4761,N_4436,N_4459);
xnor U4762 (N_4762,N_4405,N_4517);
nor U4763 (N_4763,N_4459,N_4452);
or U4764 (N_4764,N_4540,N_4585);
or U4765 (N_4765,N_4592,N_4443);
and U4766 (N_4766,N_4478,N_4583);
xnor U4767 (N_4767,N_4551,N_4453);
and U4768 (N_4768,N_4401,N_4459);
and U4769 (N_4769,N_4508,N_4581);
or U4770 (N_4770,N_4525,N_4596);
nand U4771 (N_4771,N_4446,N_4407);
xor U4772 (N_4772,N_4549,N_4486);
nor U4773 (N_4773,N_4499,N_4527);
and U4774 (N_4774,N_4501,N_4536);
or U4775 (N_4775,N_4429,N_4496);
xor U4776 (N_4776,N_4518,N_4461);
nor U4777 (N_4777,N_4527,N_4421);
or U4778 (N_4778,N_4525,N_4447);
and U4779 (N_4779,N_4471,N_4599);
or U4780 (N_4780,N_4509,N_4598);
nand U4781 (N_4781,N_4403,N_4551);
nor U4782 (N_4782,N_4576,N_4430);
nand U4783 (N_4783,N_4525,N_4471);
and U4784 (N_4784,N_4513,N_4471);
and U4785 (N_4785,N_4557,N_4516);
nor U4786 (N_4786,N_4448,N_4501);
nand U4787 (N_4787,N_4413,N_4578);
xor U4788 (N_4788,N_4568,N_4578);
xor U4789 (N_4789,N_4564,N_4402);
xnor U4790 (N_4790,N_4552,N_4587);
xor U4791 (N_4791,N_4502,N_4520);
or U4792 (N_4792,N_4592,N_4588);
nor U4793 (N_4793,N_4548,N_4420);
or U4794 (N_4794,N_4449,N_4424);
and U4795 (N_4795,N_4420,N_4556);
or U4796 (N_4796,N_4538,N_4523);
and U4797 (N_4797,N_4496,N_4468);
nor U4798 (N_4798,N_4437,N_4473);
and U4799 (N_4799,N_4408,N_4440);
or U4800 (N_4800,N_4649,N_4635);
xnor U4801 (N_4801,N_4758,N_4754);
and U4802 (N_4802,N_4699,N_4652);
xor U4803 (N_4803,N_4792,N_4664);
or U4804 (N_4804,N_4711,N_4604);
and U4805 (N_4805,N_4796,N_4615);
or U4806 (N_4806,N_4782,N_4606);
and U4807 (N_4807,N_4746,N_4666);
nand U4808 (N_4808,N_4614,N_4707);
xnor U4809 (N_4809,N_4704,N_4736);
and U4810 (N_4810,N_4709,N_4793);
or U4811 (N_4811,N_4623,N_4610);
nor U4812 (N_4812,N_4621,N_4759);
and U4813 (N_4813,N_4742,N_4688);
nor U4814 (N_4814,N_4633,N_4745);
nor U4815 (N_4815,N_4647,N_4689);
nand U4816 (N_4816,N_4613,N_4786);
xor U4817 (N_4817,N_4720,N_4772);
nor U4818 (N_4818,N_4708,N_4719);
xor U4819 (N_4819,N_4629,N_4655);
or U4820 (N_4820,N_4676,N_4732);
nand U4821 (N_4821,N_4631,N_4739);
nor U4822 (N_4822,N_4799,N_4744);
or U4823 (N_4823,N_4729,N_4774);
or U4824 (N_4824,N_4737,N_4616);
xnor U4825 (N_4825,N_4685,N_4797);
and U4826 (N_4826,N_4663,N_4778);
nand U4827 (N_4827,N_4728,N_4602);
nand U4828 (N_4828,N_4740,N_4632);
nand U4829 (N_4829,N_4640,N_4617);
nand U4830 (N_4830,N_4757,N_4651);
nor U4831 (N_4831,N_4641,N_4748);
and U4832 (N_4832,N_4715,N_4787);
or U4833 (N_4833,N_4625,N_4696);
nand U4834 (N_4834,N_4675,N_4779);
and U4835 (N_4835,N_4700,N_4743);
or U4836 (N_4836,N_4752,N_4670);
xnor U4837 (N_4837,N_4622,N_4682);
xor U4838 (N_4838,N_4644,N_4601);
xor U4839 (N_4839,N_4712,N_4726);
xor U4840 (N_4840,N_4607,N_4738);
nand U4841 (N_4841,N_4668,N_4727);
nor U4842 (N_4842,N_4687,N_4656);
or U4843 (N_4843,N_4769,N_4612);
nand U4844 (N_4844,N_4791,N_4630);
nor U4845 (N_4845,N_4654,N_4624);
or U4846 (N_4846,N_4751,N_4705);
and U4847 (N_4847,N_4662,N_4628);
and U4848 (N_4848,N_4777,N_4694);
xor U4849 (N_4849,N_4725,N_4721);
nor U4850 (N_4850,N_4788,N_4773);
nor U4851 (N_4851,N_4653,N_4648);
and U4852 (N_4852,N_4780,N_4673);
and U4853 (N_4853,N_4620,N_4749);
xnor U4854 (N_4854,N_4784,N_4771);
xor U4855 (N_4855,N_4781,N_4611);
or U4856 (N_4856,N_4710,N_4645);
nand U4857 (N_4857,N_4717,N_4686);
and U4858 (N_4858,N_4723,N_4761);
nor U4859 (N_4859,N_4683,N_4697);
nand U4860 (N_4860,N_4733,N_4693);
and U4861 (N_4861,N_4659,N_4747);
xnor U4862 (N_4862,N_4701,N_4605);
xor U4863 (N_4863,N_4785,N_4718);
nor U4864 (N_4864,N_4724,N_4608);
nor U4865 (N_4865,N_4627,N_4619);
and U4866 (N_4866,N_4661,N_4763);
xor U4867 (N_4867,N_4716,N_4756);
nor U4868 (N_4868,N_4750,N_4677);
and U4869 (N_4869,N_4684,N_4678);
xnor U4870 (N_4870,N_4681,N_4714);
nand U4871 (N_4871,N_4762,N_4760);
or U4872 (N_4872,N_4735,N_4671);
nor U4873 (N_4873,N_4703,N_4789);
xnor U4874 (N_4874,N_4639,N_4665);
nand U4875 (N_4875,N_4667,N_4646);
and U4876 (N_4876,N_4775,N_4698);
xnor U4877 (N_4877,N_4638,N_4672);
xnor U4878 (N_4878,N_4706,N_4755);
nor U4879 (N_4879,N_4734,N_4764);
nand U4880 (N_4880,N_4669,N_4753);
xor U4881 (N_4881,N_4722,N_4626);
xor U4882 (N_4882,N_4795,N_4770);
xor U4883 (N_4883,N_4643,N_4776);
nand U4884 (N_4884,N_4766,N_4600);
nor U4885 (N_4885,N_4692,N_4790);
nor U4886 (N_4886,N_4657,N_4741);
or U4887 (N_4887,N_4765,N_4702);
nand U4888 (N_4888,N_4783,N_4636);
and U4889 (N_4889,N_4695,N_4730);
nand U4890 (N_4890,N_4679,N_4618);
or U4891 (N_4891,N_4603,N_4660);
and U4892 (N_4892,N_4731,N_4658);
or U4893 (N_4893,N_4674,N_4680);
nor U4894 (N_4894,N_4767,N_4642);
nor U4895 (N_4895,N_4794,N_4691);
nor U4896 (N_4896,N_4650,N_4713);
and U4897 (N_4897,N_4768,N_4798);
xnor U4898 (N_4898,N_4637,N_4609);
xnor U4899 (N_4899,N_4634,N_4690);
or U4900 (N_4900,N_4648,N_4758);
nor U4901 (N_4901,N_4739,N_4772);
or U4902 (N_4902,N_4706,N_4771);
xor U4903 (N_4903,N_4615,N_4676);
nand U4904 (N_4904,N_4626,N_4631);
xnor U4905 (N_4905,N_4786,N_4632);
and U4906 (N_4906,N_4789,N_4750);
nor U4907 (N_4907,N_4780,N_4719);
nor U4908 (N_4908,N_4691,N_4670);
xnor U4909 (N_4909,N_4730,N_4779);
nand U4910 (N_4910,N_4672,N_4792);
nor U4911 (N_4911,N_4707,N_4694);
or U4912 (N_4912,N_4607,N_4742);
xor U4913 (N_4913,N_4796,N_4757);
and U4914 (N_4914,N_4650,N_4692);
nor U4915 (N_4915,N_4658,N_4606);
nor U4916 (N_4916,N_4658,N_4759);
nor U4917 (N_4917,N_4764,N_4796);
xor U4918 (N_4918,N_4694,N_4673);
nand U4919 (N_4919,N_4630,N_4756);
xor U4920 (N_4920,N_4608,N_4702);
nand U4921 (N_4921,N_4724,N_4751);
nand U4922 (N_4922,N_4706,N_4722);
or U4923 (N_4923,N_4762,N_4799);
xor U4924 (N_4924,N_4628,N_4695);
and U4925 (N_4925,N_4672,N_4605);
or U4926 (N_4926,N_4631,N_4794);
nor U4927 (N_4927,N_4725,N_4674);
xor U4928 (N_4928,N_4643,N_4737);
nor U4929 (N_4929,N_4685,N_4604);
nand U4930 (N_4930,N_4745,N_4637);
nand U4931 (N_4931,N_4714,N_4754);
or U4932 (N_4932,N_4600,N_4742);
and U4933 (N_4933,N_4660,N_4794);
and U4934 (N_4934,N_4759,N_4777);
and U4935 (N_4935,N_4613,N_4658);
nand U4936 (N_4936,N_4766,N_4736);
or U4937 (N_4937,N_4708,N_4691);
xnor U4938 (N_4938,N_4748,N_4654);
or U4939 (N_4939,N_4676,N_4779);
nand U4940 (N_4940,N_4600,N_4621);
or U4941 (N_4941,N_4738,N_4604);
nor U4942 (N_4942,N_4642,N_4719);
or U4943 (N_4943,N_4795,N_4799);
nand U4944 (N_4944,N_4718,N_4675);
and U4945 (N_4945,N_4716,N_4610);
nand U4946 (N_4946,N_4675,N_4613);
or U4947 (N_4947,N_4610,N_4738);
xnor U4948 (N_4948,N_4781,N_4707);
and U4949 (N_4949,N_4735,N_4698);
nor U4950 (N_4950,N_4647,N_4648);
or U4951 (N_4951,N_4705,N_4604);
xnor U4952 (N_4952,N_4752,N_4661);
and U4953 (N_4953,N_4672,N_4705);
xor U4954 (N_4954,N_4731,N_4754);
or U4955 (N_4955,N_4698,N_4653);
xor U4956 (N_4956,N_4658,N_4689);
xor U4957 (N_4957,N_4638,N_4646);
xnor U4958 (N_4958,N_4694,N_4624);
nor U4959 (N_4959,N_4755,N_4605);
nand U4960 (N_4960,N_4667,N_4616);
and U4961 (N_4961,N_4730,N_4692);
xnor U4962 (N_4962,N_4630,N_4652);
and U4963 (N_4963,N_4632,N_4747);
xor U4964 (N_4964,N_4741,N_4679);
or U4965 (N_4965,N_4628,N_4610);
nor U4966 (N_4966,N_4752,N_4716);
and U4967 (N_4967,N_4766,N_4618);
or U4968 (N_4968,N_4735,N_4721);
xor U4969 (N_4969,N_4664,N_4666);
nor U4970 (N_4970,N_4716,N_4768);
xnor U4971 (N_4971,N_4670,N_4722);
xor U4972 (N_4972,N_4756,N_4763);
or U4973 (N_4973,N_4798,N_4762);
or U4974 (N_4974,N_4638,N_4793);
nand U4975 (N_4975,N_4652,N_4659);
xnor U4976 (N_4976,N_4626,N_4693);
nand U4977 (N_4977,N_4665,N_4602);
nor U4978 (N_4978,N_4706,N_4660);
nor U4979 (N_4979,N_4683,N_4766);
xnor U4980 (N_4980,N_4795,N_4758);
or U4981 (N_4981,N_4784,N_4774);
xnor U4982 (N_4982,N_4755,N_4602);
or U4983 (N_4983,N_4685,N_4701);
or U4984 (N_4984,N_4608,N_4655);
xnor U4985 (N_4985,N_4612,N_4771);
or U4986 (N_4986,N_4788,N_4690);
and U4987 (N_4987,N_4789,N_4721);
nand U4988 (N_4988,N_4651,N_4705);
nand U4989 (N_4989,N_4611,N_4740);
nand U4990 (N_4990,N_4631,N_4695);
xor U4991 (N_4991,N_4792,N_4704);
or U4992 (N_4992,N_4716,N_4661);
or U4993 (N_4993,N_4708,N_4695);
xnor U4994 (N_4994,N_4722,N_4614);
or U4995 (N_4995,N_4632,N_4722);
and U4996 (N_4996,N_4766,N_4641);
xnor U4997 (N_4997,N_4794,N_4601);
nor U4998 (N_4998,N_4725,N_4693);
and U4999 (N_4999,N_4694,N_4690);
xnor U5000 (N_5000,N_4912,N_4962);
nand U5001 (N_5001,N_4980,N_4909);
nor U5002 (N_5002,N_4932,N_4856);
xor U5003 (N_5003,N_4851,N_4849);
and U5004 (N_5004,N_4908,N_4954);
nand U5005 (N_5005,N_4844,N_4850);
or U5006 (N_5006,N_4821,N_4956);
or U5007 (N_5007,N_4842,N_4863);
nor U5008 (N_5008,N_4910,N_4959);
xor U5009 (N_5009,N_4978,N_4883);
nor U5010 (N_5010,N_4893,N_4835);
xor U5011 (N_5011,N_4871,N_4867);
and U5012 (N_5012,N_4934,N_4963);
xnor U5013 (N_5013,N_4936,N_4941);
nor U5014 (N_5014,N_4981,N_4872);
nor U5015 (N_5015,N_4896,N_4999);
and U5016 (N_5016,N_4989,N_4824);
and U5017 (N_5017,N_4974,N_4917);
nand U5018 (N_5018,N_4820,N_4929);
xnor U5019 (N_5019,N_4894,N_4803);
xnor U5020 (N_5020,N_4923,N_4855);
nor U5021 (N_5021,N_4916,N_4944);
and U5022 (N_5022,N_4887,N_4951);
xor U5023 (N_5023,N_4837,N_4841);
and U5024 (N_5024,N_4906,N_4848);
or U5025 (N_5025,N_4890,N_4976);
nor U5026 (N_5026,N_4957,N_4858);
xor U5027 (N_5027,N_4965,N_4995);
xnor U5028 (N_5028,N_4886,N_4878);
xnor U5029 (N_5029,N_4831,N_4950);
or U5030 (N_5030,N_4809,N_4960);
or U5031 (N_5031,N_4970,N_4975);
and U5032 (N_5032,N_4961,N_4972);
nor U5033 (N_5033,N_4977,N_4829);
nand U5034 (N_5034,N_4808,N_4928);
or U5035 (N_5035,N_4805,N_4876);
or U5036 (N_5036,N_4862,N_4922);
and U5037 (N_5037,N_4816,N_4845);
nor U5038 (N_5038,N_4983,N_4881);
nand U5039 (N_5039,N_4826,N_4869);
xnor U5040 (N_5040,N_4888,N_4992);
nor U5041 (N_5041,N_4882,N_4939);
xor U5042 (N_5042,N_4840,N_4924);
nor U5043 (N_5043,N_4815,N_4830);
or U5044 (N_5044,N_4846,N_4880);
nand U5045 (N_5045,N_4938,N_4898);
and U5046 (N_5046,N_4897,N_4994);
xor U5047 (N_5047,N_4966,N_4813);
nor U5048 (N_5048,N_4919,N_4901);
xor U5049 (N_5049,N_4879,N_4873);
nor U5050 (N_5050,N_4877,N_4996);
or U5051 (N_5051,N_4953,N_4931);
or U5052 (N_5052,N_4902,N_4834);
or U5053 (N_5053,N_4870,N_4860);
nor U5054 (N_5054,N_4895,N_4986);
or U5055 (N_5055,N_4971,N_4920);
nand U5056 (N_5056,N_4905,N_4955);
and U5057 (N_5057,N_4921,N_4811);
nor U5058 (N_5058,N_4952,N_4943);
nor U5059 (N_5059,N_4817,N_4822);
nor U5060 (N_5060,N_4868,N_4969);
and U5061 (N_5061,N_4949,N_4812);
nand U5062 (N_5062,N_4991,N_4839);
or U5063 (N_5063,N_4899,N_4925);
nor U5064 (N_5064,N_4979,N_4987);
or U5065 (N_5065,N_4804,N_4827);
nor U5066 (N_5066,N_4942,N_4935);
nand U5067 (N_5067,N_4884,N_4800);
xnor U5068 (N_5068,N_4927,N_4801);
or U5069 (N_5069,N_4865,N_4930);
nor U5070 (N_5070,N_4967,N_4903);
nand U5071 (N_5071,N_4875,N_4854);
or U5072 (N_5072,N_4926,N_4940);
nor U5073 (N_5073,N_4914,N_4833);
or U5074 (N_5074,N_4892,N_4885);
nand U5075 (N_5075,N_4904,N_4866);
nand U5076 (N_5076,N_4984,N_4832);
xnor U5077 (N_5077,N_4861,N_4982);
or U5078 (N_5078,N_4937,N_4946);
or U5079 (N_5079,N_4857,N_4948);
xnor U5080 (N_5080,N_4990,N_4945);
and U5081 (N_5081,N_4973,N_4889);
and U5082 (N_5082,N_4859,N_4819);
nand U5083 (N_5083,N_4853,N_4998);
nand U5084 (N_5084,N_4907,N_4818);
and U5085 (N_5085,N_4874,N_4985);
nand U5086 (N_5086,N_4852,N_4847);
nand U5087 (N_5087,N_4993,N_4988);
or U5088 (N_5088,N_4828,N_4933);
nor U5089 (N_5089,N_4838,N_4968);
xnor U5090 (N_5090,N_4843,N_4814);
nand U5091 (N_5091,N_4997,N_4900);
nor U5092 (N_5092,N_4810,N_4947);
nor U5093 (N_5093,N_4802,N_4806);
nor U5094 (N_5094,N_4823,N_4918);
nand U5095 (N_5095,N_4964,N_4807);
xor U5096 (N_5096,N_4891,N_4864);
nor U5097 (N_5097,N_4836,N_4913);
nor U5098 (N_5098,N_4915,N_4911);
xnor U5099 (N_5099,N_4958,N_4825);
xnor U5100 (N_5100,N_4956,N_4932);
and U5101 (N_5101,N_4911,N_4821);
and U5102 (N_5102,N_4840,N_4944);
nor U5103 (N_5103,N_4955,N_4866);
or U5104 (N_5104,N_4952,N_4859);
or U5105 (N_5105,N_4871,N_4843);
nand U5106 (N_5106,N_4951,N_4984);
and U5107 (N_5107,N_4903,N_4802);
or U5108 (N_5108,N_4885,N_4900);
xnor U5109 (N_5109,N_4816,N_4817);
xnor U5110 (N_5110,N_4814,N_4900);
or U5111 (N_5111,N_4843,N_4986);
or U5112 (N_5112,N_4973,N_4958);
nand U5113 (N_5113,N_4914,N_4981);
nand U5114 (N_5114,N_4965,N_4829);
nor U5115 (N_5115,N_4884,N_4984);
or U5116 (N_5116,N_4952,N_4981);
and U5117 (N_5117,N_4802,N_4891);
xor U5118 (N_5118,N_4951,N_4885);
or U5119 (N_5119,N_4820,N_4956);
or U5120 (N_5120,N_4940,N_4943);
xor U5121 (N_5121,N_4828,N_4895);
or U5122 (N_5122,N_4998,N_4988);
xor U5123 (N_5123,N_4817,N_4932);
nand U5124 (N_5124,N_4818,N_4800);
nor U5125 (N_5125,N_4872,N_4921);
nor U5126 (N_5126,N_4807,N_4847);
and U5127 (N_5127,N_4948,N_4894);
or U5128 (N_5128,N_4897,N_4965);
nand U5129 (N_5129,N_4951,N_4940);
nor U5130 (N_5130,N_4886,N_4806);
and U5131 (N_5131,N_4828,N_4923);
and U5132 (N_5132,N_4884,N_4819);
xnor U5133 (N_5133,N_4852,N_4973);
or U5134 (N_5134,N_4815,N_4997);
nor U5135 (N_5135,N_4975,N_4878);
and U5136 (N_5136,N_4983,N_4951);
nor U5137 (N_5137,N_4891,N_4882);
nand U5138 (N_5138,N_4988,N_4965);
nor U5139 (N_5139,N_4880,N_4935);
or U5140 (N_5140,N_4891,N_4975);
or U5141 (N_5141,N_4981,N_4852);
nand U5142 (N_5142,N_4980,N_4911);
nor U5143 (N_5143,N_4892,N_4932);
nand U5144 (N_5144,N_4863,N_4819);
or U5145 (N_5145,N_4983,N_4981);
nor U5146 (N_5146,N_4935,N_4907);
or U5147 (N_5147,N_4809,N_4880);
and U5148 (N_5148,N_4808,N_4875);
nand U5149 (N_5149,N_4978,N_4987);
nor U5150 (N_5150,N_4880,N_4953);
or U5151 (N_5151,N_4907,N_4993);
xnor U5152 (N_5152,N_4892,N_4896);
and U5153 (N_5153,N_4930,N_4996);
and U5154 (N_5154,N_4878,N_4923);
and U5155 (N_5155,N_4820,N_4810);
nor U5156 (N_5156,N_4885,N_4801);
xnor U5157 (N_5157,N_4903,N_4951);
or U5158 (N_5158,N_4865,N_4878);
and U5159 (N_5159,N_4902,N_4891);
nor U5160 (N_5160,N_4865,N_4992);
nor U5161 (N_5161,N_4923,N_4873);
nor U5162 (N_5162,N_4973,N_4966);
nand U5163 (N_5163,N_4857,N_4820);
or U5164 (N_5164,N_4981,N_4957);
nand U5165 (N_5165,N_4822,N_4998);
or U5166 (N_5166,N_4967,N_4976);
nand U5167 (N_5167,N_4960,N_4976);
nand U5168 (N_5168,N_4846,N_4866);
nor U5169 (N_5169,N_4806,N_4835);
nor U5170 (N_5170,N_4935,N_4908);
and U5171 (N_5171,N_4886,N_4914);
nor U5172 (N_5172,N_4924,N_4954);
nor U5173 (N_5173,N_4939,N_4926);
nand U5174 (N_5174,N_4878,N_4843);
and U5175 (N_5175,N_4867,N_4849);
xor U5176 (N_5176,N_4991,N_4985);
nand U5177 (N_5177,N_4861,N_4893);
nor U5178 (N_5178,N_4883,N_4859);
nor U5179 (N_5179,N_4818,N_4887);
or U5180 (N_5180,N_4909,N_4984);
xnor U5181 (N_5181,N_4828,N_4824);
or U5182 (N_5182,N_4841,N_4996);
and U5183 (N_5183,N_4963,N_4883);
or U5184 (N_5184,N_4930,N_4848);
nand U5185 (N_5185,N_4943,N_4944);
nand U5186 (N_5186,N_4858,N_4908);
and U5187 (N_5187,N_4961,N_4816);
nor U5188 (N_5188,N_4914,N_4980);
and U5189 (N_5189,N_4889,N_4999);
xor U5190 (N_5190,N_4826,N_4902);
xnor U5191 (N_5191,N_4984,N_4899);
nand U5192 (N_5192,N_4926,N_4973);
nand U5193 (N_5193,N_4834,N_4850);
nand U5194 (N_5194,N_4822,N_4834);
and U5195 (N_5195,N_4802,N_4912);
nor U5196 (N_5196,N_4916,N_4836);
and U5197 (N_5197,N_4985,N_4993);
nor U5198 (N_5198,N_4805,N_4940);
and U5199 (N_5199,N_4909,N_4973);
nand U5200 (N_5200,N_5076,N_5069);
xor U5201 (N_5201,N_5043,N_5017);
and U5202 (N_5202,N_5002,N_5150);
or U5203 (N_5203,N_5044,N_5041);
nor U5204 (N_5204,N_5158,N_5174);
or U5205 (N_5205,N_5062,N_5065);
and U5206 (N_5206,N_5194,N_5055);
xor U5207 (N_5207,N_5006,N_5135);
or U5208 (N_5208,N_5033,N_5164);
and U5209 (N_5209,N_5104,N_5068);
and U5210 (N_5210,N_5145,N_5079);
or U5211 (N_5211,N_5110,N_5122);
nand U5212 (N_5212,N_5107,N_5120);
nand U5213 (N_5213,N_5163,N_5175);
or U5214 (N_5214,N_5151,N_5116);
or U5215 (N_5215,N_5003,N_5167);
nand U5216 (N_5216,N_5064,N_5028);
xnor U5217 (N_5217,N_5013,N_5102);
xor U5218 (N_5218,N_5086,N_5010);
and U5219 (N_5219,N_5057,N_5052);
or U5220 (N_5220,N_5058,N_5075);
nor U5221 (N_5221,N_5106,N_5072);
nor U5222 (N_5222,N_5063,N_5087);
xor U5223 (N_5223,N_5112,N_5166);
nor U5224 (N_5224,N_5004,N_5051);
xor U5225 (N_5225,N_5040,N_5146);
xor U5226 (N_5226,N_5142,N_5084);
or U5227 (N_5227,N_5162,N_5159);
or U5228 (N_5228,N_5067,N_5071);
nand U5229 (N_5229,N_5114,N_5094);
nor U5230 (N_5230,N_5190,N_5161);
nand U5231 (N_5231,N_5054,N_5129);
or U5232 (N_5232,N_5137,N_5053);
xnor U5233 (N_5233,N_5191,N_5083);
nand U5234 (N_5234,N_5088,N_5005);
nand U5235 (N_5235,N_5093,N_5082);
nor U5236 (N_5236,N_5188,N_5173);
nand U5237 (N_5237,N_5049,N_5179);
or U5238 (N_5238,N_5035,N_5187);
xnor U5239 (N_5239,N_5061,N_5123);
nand U5240 (N_5240,N_5019,N_5000);
or U5241 (N_5241,N_5176,N_5144);
or U5242 (N_5242,N_5073,N_5039);
xnor U5243 (N_5243,N_5130,N_5012);
and U5244 (N_5244,N_5070,N_5155);
and U5245 (N_5245,N_5115,N_5074);
nor U5246 (N_5246,N_5133,N_5143);
nor U5247 (N_5247,N_5147,N_5030);
and U5248 (N_5248,N_5031,N_5118);
xor U5249 (N_5249,N_5056,N_5016);
nand U5250 (N_5250,N_5152,N_5050);
nor U5251 (N_5251,N_5127,N_5092);
nand U5252 (N_5252,N_5117,N_5189);
nor U5253 (N_5253,N_5091,N_5183);
nor U5254 (N_5254,N_5136,N_5078);
nand U5255 (N_5255,N_5193,N_5108);
nor U5256 (N_5256,N_5148,N_5021);
nor U5257 (N_5257,N_5022,N_5170);
nand U5258 (N_5258,N_5103,N_5128);
or U5259 (N_5259,N_5037,N_5184);
nand U5260 (N_5260,N_5066,N_5134);
xor U5261 (N_5261,N_5197,N_5077);
nor U5262 (N_5262,N_5192,N_5060);
nor U5263 (N_5263,N_5090,N_5149);
or U5264 (N_5264,N_5080,N_5015);
nor U5265 (N_5265,N_5042,N_5124);
xnor U5266 (N_5266,N_5113,N_5096);
nor U5267 (N_5267,N_5100,N_5157);
xnor U5268 (N_5268,N_5001,N_5026);
nor U5269 (N_5269,N_5105,N_5154);
and U5270 (N_5270,N_5139,N_5126);
nand U5271 (N_5271,N_5089,N_5132);
xnor U5272 (N_5272,N_5023,N_5195);
and U5273 (N_5273,N_5007,N_5009);
and U5274 (N_5274,N_5098,N_5185);
and U5275 (N_5275,N_5034,N_5181);
or U5276 (N_5276,N_5109,N_5140);
nor U5277 (N_5277,N_5171,N_5048);
nor U5278 (N_5278,N_5198,N_5111);
and U5279 (N_5279,N_5008,N_5165);
and U5280 (N_5280,N_5172,N_5036);
nand U5281 (N_5281,N_5099,N_5029);
or U5282 (N_5282,N_5046,N_5101);
nor U5283 (N_5283,N_5097,N_5119);
nor U5284 (N_5284,N_5047,N_5059);
and U5285 (N_5285,N_5025,N_5027);
nand U5286 (N_5286,N_5196,N_5182);
nand U5287 (N_5287,N_5032,N_5186);
nand U5288 (N_5288,N_5014,N_5169);
xor U5289 (N_5289,N_5199,N_5138);
nand U5290 (N_5290,N_5018,N_5125);
xnor U5291 (N_5291,N_5085,N_5131);
nor U5292 (N_5292,N_5038,N_5177);
and U5293 (N_5293,N_5011,N_5160);
and U5294 (N_5294,N_5121,N_5081);
nor U5295 (N_5295,N_5024,N_5141);
or U5296 (N_5296,N_5178,N_5020);
nor U5297 (N_5297,N_5095,N_5168);
and U5298 (N_5298,N_5180,N_5156);
and U5299 (N_5299,N_5045,N_5153);
nor U5300 (N_5300,N_5074,N_5089);
and U5301 (N_5301,N_5093,N_5161);
xnor U5302 (N_5302,N_5044,N_5126);
and U5303 (N_5303,N_5175,N_5196);
nor U5304 (N_5304,N_5031,N_5192);
xor U5305 (N_5305,N_5157,N_5104);
xor U5306 (N_5306,N_5086,N_5157);
xor U5307 (N_5307,N_5064,N_5037);
xor U5308 (N_5308,N_5148,N_5177);
and U5309 (N_5309,N_5147,N_5072);
and U5310 (N_5310,N_5090,N_5180);
or U5311 (N_5311,N_5184,N_5146);
xnor U5312 (N_5312,N_5004,N_5113);
or U5313 (N_5313,N_5139,N_5157);
nand U5314 (N_5314,N_5082,N_5065);
nor U5315 (N_5315,N_5018,N_5029);
and U5316 (N_5316,N_5152,N_5008);
nor U5317 (N_5317,N_5118,N_5046);
or U5318 (N_5318,N_5101,N_5000);
and U5319 (N_5319,N_5030,N_5150);
nor U5320 (N_5320,N_5011,N_5108);
and U5321 (N_5321,N_5164,N_5091);
nor U5322 (N_5322,N_5183,N_5115);
and U5323 (N_5323,N_5191,N_5048);
nor U5324 (N_5324,N_5005,N_5063);
or U5325 (N_5325,N_5102,N_5156);
nor U5326 (N_5326,N_5058,N_5090);
nor U5327 (N_5327,N_5098,N_5186);
nand U5328 (N_5328,N_5047,N_5124);
nand U5329 (N_5329,N_5199,N_5118);
nor U5330 (N_5330,N_5197,N_5099);
xnor U5331 (N_5331,N_5145,N_5058);
or U5332 (N_5332,N_5153,N_5162);
or U5333 (N_5333,N_5155,N_5103);
xor U5334 (N_5334,N_5024,N_5096);
nor U5335 (N_5335,N_5096,N_5029);
and U5336 (N_5336,N_5161,N_5092);
xor U5337 (N_5337,N_5130,N_5165);
xnor U5338 (N_5338,N_5157,N_5030);
nor U5339 (N_5339,N_5037,N_5137);
nand U5340 (N_5340,N_5071,N_5191);
or U5341 (N_5341,N_5157,N_5060);
xnor U5342 (N_5342,N_5084,N_5196);
nor U5343 (N_5343,N_5179,N_5133);
nor U5344 (N_5344,N_5084,N_5038);
xnor U5345 (N_5345,N_5006,N_5023);
xor U5346 (N_5346,N_5088,N_5174);
nand U5347 (N_5347,N_5088,N_5139);
xor U5348 (N_5348,N_5060,N_5069);
nor U5349 (N_5349,N_5006,N_5067);
xnor U5350 (N_5350,N_5003,N_5099);
nand U5351 (N_5351,N_5015,N_5128);
nor U5352 (N_5352,N_5103,N_5134);
or U5353 (N_5353,N_5162,N_5010);
xnor U5354 (N_5354,N_5127,N_5015);
or U5355 (N_5355,N_5105,N_5143);
nor U5356 (N_5356,N_5023,N_5059);
nor U5357 (N_5357,N_5171,N_5159);
and U5358 (N_5358,N_5119,N_5037);
xor U5359 (N_5359,N_5104,N_5180);
or U5360 (N_5360,N_5162,N_5185);
and U5361 (N_5361,N_5031,N_5074);
xnor U5362 (N_5362,N_5029,N_5124);
and U5363 (N_5363,N_5006,N_5163);
nand U5364 (N_5364,N_5078,N_5140);
or U5365 (N_5365,N_5127,N_5131);
nand U5366 (N_5366,N_5121,N_5199);
or U5367 (N_5367,N_5066,N_5049);
or U5368 (N_5368,N_5191,N_5045);
nor U5369 (N_5369,N_5174,N_5039);
xor U5370 (N_5370,N_5141,N_5057);
xnor U5371 (N_5371,N_5055,N_5060);
xnor U5372 (N_5372,N_5076,N_5179);
nor U5373 (N_5373,N_5137,N_5091);
or U5374 (N_5374,N_5166,N_5047);
xnor U5375 (N_5375,N_5194,N_5187);
xor U5376 (N_5376,N_5075,N_5176);
and U5377 (N_5377,N_5148,N_5114);
nor U5378 (N_5378,N_5107,N_5166);
xnor U5379 (N_5379,N_5061,N_5070);
or U5380 (N_5380,N_5081,N_5060);
xnor U5381 (N_5381,N_5013,N_5175);
nand U5382 (N_5382,N_5101,N_5131);
xnor U5383 (N_5383,N_5018,N_5175);
xor U5384 (N_5384,N_5012,N_5147);
and U5385 (N_5385,N_5057,N_5026);
nor U5386 (N_5386,N_5036,N_5144);
and U5387 (N_5387,N_5066,N_5190);
nand U5388 (N_5388,N_5184,N_5062);
and U5389 (N_5389,N_5051,N_5022);
nor U5390 (N_5390,N_5028,N_5069);
nand U5391 (N_5391,N_5018,N_5017);
or U5392 (N_5392,N_5026,N_5133);
xnor U5393 (N_5393,N_5080,N_5027);
nor U5394 (N_5394,N_5080,N_5070);
nor U5395 (N_5395,N_5087,N_5180);
or U5396 (N_5396,N_5172,N_5170);
or U5397 (N_5397,N_5194,N_5037);
xnor U5398 (N_5398,N_5015,N_5025);
nand U5399 (N_5399,N_5187,N_5121);
or U5400 (N_5400,N_5284,N_5322);
nor U5401 (N_5401,N_5226,N_5266);
or U5402 (N_5402,N_5363,N_5259);
and U5403 (N_5403,N_5305,N_5232);
nand U5404 (N_5404,N_5308,N_5248);
xnor U5405 (N_5405,N_5332,N_5272);
xnor U5406 (N_5406,N_5224,N_5207);
xnor U5407 (N_5407,N_5345,N_5391);
nand U5408 (N_5408,N_5228,N_5374);
nand U5409 (N_5409,N_5244,N_5213);
and U5410 (N_5410,N_5376,N_5261);
and U5411 (N_5411,N_5202,N_5393);
xor U5412 (N_5412,N_5307,N_5375);
nor U5413 (N_5413,N_5209,N_5344);
xnor U5414 (N_5414,N_5392,N_5329);
and U5415 (N_5415,N_5319,N_5301);
nor U5416 (N_5416,N_5324,N_5201);
nand U5417 (N_5417,N_5204,N_5221);
nand U5418 (N_5418,N_5241,N_5263);
nand U5419 (N_5419,N_5220,N_5208);
nand U5420 (N_5420,N_5382,N_5317);
nor U5421 (N_5421,N_5397,N_5291);
or U5422 (N_5422,N_5326,N_5269);
or U5423 (N_5423,N_5369,N_5318);
and U5424 (N_5424,N_5249,N_5271);
nor U5425 (N_5425,N_5388,N_5304);
and U5426 (N_5426,N_5359,N_5377);
or U5427 (N_5427,N_5298,N_5235);
xor U5428 (N_5428,N_5245,N_5358);
and U5429 (N_5429,N_5306,N_5311);
nand U5430 (N_5430,N_5355,N_5340);
nand U5431 (N_5431,N_5357,N_5383);
and U5432 (N_5432,N_5323,N_5227);
and U5433 (N_5433,N_5243,N_5257);
nor U5434 (N_5434,N_5297,N_5264);
nand U5435 (N_5435,N_5315,N_5282);
and U5436 (N_5436,N_5293,N_5370);
or U5437 (N_5437,N_5260,N_5362);
or U5438 (N_5438,N_5251,N_5217);
nand U5439 (N_5439,N_5210,N_5237);
xnor U5440 (N_5440,N_5250,N_5247);
and U5441 (N_5441,N_5278,N_5330);
nor U5442 (N_5442,N_5342,N_5381);
and U5443 (N_5443,N_5236,N_5270);
and U5444 (N_5444,N_5312,N_5333);
xnor U5445 (N_5445,N_5273,N_5335);
nand U5446 (N_5446,N_5200,N_5368);
and U5447 (N_5447,N_5215,N_5339);
nand U5448 (N_5448,N_5379,N_5222);
and U5449 (N_5449,N_5255,N_5239);
xor U5450 (N_5450,N_5341,N_5299);
or U5451 (N_5451,N_5292,N_5240);
nand U5452 (N_5452,N_5225,N_5294);
xnor U5453 (N_5453,N_5296,N_5238);
nand U5454 (N_5454,N_5218,N_5366);
xor U5455 (N_5455,N_5351,N_5219);
nor U5456 (N_5456,N_5206,N_5394);
and U5457 (N_5457,N_5398,N_5229);
or U5458 (N_5458,N_5203,N_5328);
xnor U5459 (N_5459,N_5290,N_5399);
or U5460 (N_5460,N_5371,N_5216);
nor U5461 (N_5461,N_5295,N_5354);
and U5462 (N_5462,N_5364,N_5380);
and U5463 (N_5463,N_5276,N_5242);
nor U5464 (N_5464,N_5390,N_5395);
and U5465 (N_5465,N_5253,N_5265);
or U5466 (N_5466,N_5230,N_5288);
nand U5467 (N_5467,N_5205,N_5289);
or U5468 (N_5468,N_5321,N_5385);
nor U5469 (N_5469,N_5246,N_5350);
xor U5470 (N_5470,N_5331,N_5372);
or U5471 (N_5471,N_5353,N_5274);
and U5472 (N_5472,N_5389,N_5268);
or U5473 (N_5473,N_5384,N_5283);
nand U5474 (N_5474,N_5347,N_5254);
xor U5475 (N_5475,N_5378,N_5336);
nand U5476 (N_5476,N_5310,N_5386);
nor U5477 (N_5477,N_5300,N_5281);
nand U5478 (N_5478,N_5313,N_5258);
xnor U5479 (N_5479,N_5231,N_5275);
nand U5480 (N_5480,N_5356,N_5334);
xor U5481 (N_5481,N_5302,N_5352);
nor U5482 (N_5482,N_5277,N_5214);
nor U5483 (N_5483,N_5367,N_5387);
and U5484 (N_5484,N_5349,N_5223);
nand U5485 (N_5485,N_5338,N_5396);
nor U5486 (N_5486,N_5262,N_5346);
and U5487 (N_5487,N_5373,N_5211);
xor U5488 (N_5488,N_5287,N_5337);
and U5489 (N_5489,N_5314,N_5233);
xnor U5490 (N_5490,N_5285,N_5361);
nor U5491 (N_5491,N_5267,N_5303);
nor U5492 (N_5492,N_5286,N_5325);
nor U5493 (N_5493,N_5360,N_5309);
or U5494 (N_5494,N_5365,N_5234);
xor U5495 (N_5495,N_5320,N_5348);
and U5496 (N_5496,N_5316,N_5256);
or U5497 (N_5497,N_5327,N_5279);
nand U5498 (N_5498,N_5343,N_5212);
nand U5499 (N_5499,N_5252,N_5280);
or U5500 (N_5500,N_5249,N_5351);
or U5501 (N_5501,N_5338,N_5204);
or U5502 (N_5502,N_5253,N_5225);
or U5503 (N_5503,N_5249,N_5320);
and U5504 (N_5504,N_5269,N_5289);
nand U5505 (N_5505,N_5241,N_5351);
or U5506 (N_5506,N_5369,N_5215);
nand U5507 (N_5507,N_5373,N_5213);
xnor U5508 (N_5508,N_5249,N_5268);
xor U5509 (N_5509,N_5229,N_5273);
xnor U5510 (N_5510,N_5350,N_5393);
xnor U5511 (N_5511,N_5359,N_5226);
xor U5512 (N_5512,N_5370,N_5272);
xor U5513 (N_5513,N_5311,N_5227);
nand U5514 (N_5514,N_5339,N_5279);
xnor U5515 (N_5515,N_5280,N_5303);
nor U5516 (N_5516,N_5242,N_5370);
nand U5517 (N_5517,N_5256,N_5350);
xnor U5518 (N_5518,N_5335,N_5201);
xnor U5519 (N_5519,N_5331,N_5300);
or U5520 (N_5520,N_5391,N_5318);
or U5521 (N_5521,N_5258,N_5232);
nand U5522 (N_5522,N_5242,N_5332);
nor U5523 (N_5523,N_5339,N_5367);
or U5524 (N_5524,N_5374,N_5225);
nor U5525 (N_5525,N_5333,N_5264);
and U5526 (N_5526,N_5315,N_5222);
nand U5527 (N_5527,N_5231,N_5393);
xor U5528 (N_5528,N_5328,N_5327);
nor U5529 (N_5529,N_5352,N_5369);
and U5530 (N_5530,N_5235,N_5251);
or U5531 (N_5531,N_5226,N_5323);
or U5532 (N_5532,N_5254,N_5302);
or U5533 (N_5533,N_5285,N_5326);
and U5534 (N_5534,N_5237,N_5371);
and U5535 (N_5535,N_5332,N_5346);
nand U5536 (N_5536,N_5232,N_5348);
nor U5537 (N_5537,N_5244,N_5291);
xor U5538 (N_5538,N_5215,N_5243);
nand U5539 (N_5539,N_5323,N_5349);
nand U5540 (N_5540,N_5276,N_5326);
nand U5541 (N_5541,N_5366,N_5208);
nand U5542 (N_5542,N_5326,N_5394);
or U5543 (N_5543,N_5377,N_5225);
nor U5544 (N_5544,N_5367,N_5218);
xor U5545 (N_5545,N_5386,N_5225);
or U5546 (N_5546,N_5377,N_5358);
nand U5547 (N_5547,N_5384,N_5389);
nor U5548 (N_5548,N_5328,N_5362);
or U5549 (N_5549,N_5239,N_5396);
nand U5550 (N_5550,N_5214,N_5350);
xnor U5551 (N_5551,N_5251,N_5269);
nor U5552 (N_5552,N_5317,N_5320);
xor U5553 (N_5553,N_5376,N_5266);
nand U5554 (N_5554,N_5257,N_5357);
or U5555 (N_5555,N_5260,N_5349);
and U5556 (N_5556,N_5374,N_5312);
and U5557 (N_5557,N_5209,N_5329);
xor U5558 (N_5558,N_5319,N_5372);
and U5559 (N_5559,N_5358,N_5202);
xnor U5560 (N_5560,N_5370,N_5358);
and U5561 (N_5561,N_5262,N_5363);
and U5562 (N_5562,N_5387,N_5246);
nor U5563 (N_5563,N_5267,N_5314);
and U5564 (N_5564,N_5237,N_5289);
nand U5565 (N_5565,N_5208,N_5260);
xor U5566 (N_5566,N_5290,N_5279);
and U5567 (N_5567,N_5281,N_5298);
nand U5568 (N_5568,N_5218,N_5217);
nand U5569 (N_5569,N_5368,N_5215);
nor U5570 (N_5570,N_5380,N_5279);
xnor U5571 (N_5571,N_5317,N_5221);
xor U5572 (N_5572,N_5235,N_5314);
and U5573 (N_5573,N_5251,N_5282);
and U5574 (N_5574,N_5382,N_5298);
xor U5575 (N_5575,N_5243,N_5383);
xnor U5576 (N_5576,N_5251,N_5359);
xor U5577 (N_5577,N_5288,N_5339);
xor U5578 (N_5578,N_5339,N_5226);
or U5579 (N_5579,N_5225,N_5209);
or U5580 (N_5580,N_5234,N_5277);
nor U5581 (N_5581,N_5277,N_5388);
nor U5582 (N_5582,N_5365,N_5251);
and U5583 (N_5583,N_5204,N_5392);
and U5584 (N_5584,N_5385,N_5230);
or U5585 (N_5585,N_5253,N_5382);
xor U5586 (N_5586,N_5292,N_5303);
or U5587 (N_5587,N_5299,N_5252);
nand U5588 (N_5588,N_5312,N_5305);
or U5589 (N_5589,N_5388,N_5350);
xnor U5590 (N_5590,N_5259,N_5299);
or U5591 (N_5591,N_5277,N_5370);
and U5592 (N_5592,N_5357,N_5372);
xor U5593 (N_5593,N_5314,N_5393);
nor U5594 (N_5594,N_5299,N_5248);
nor U5595 (N_5595,N_5370,N_5220);
nor U5596 (N_5596,N_5333,N_5306);
xnor U5597 (N_5597,N_5211,N_5225);
and U5598 (N_5598,N_5286,N_5206);
and U5599 (N_5599,N_5224,N_5388);
and U5600 (N_5600,N_5414,N_5454);
nor U5601 (N_5601,N_5494,N_5583);
xnor U5602 (N_5602,N_5443,N_5462);
nor U5603 (N_5603,N_5472,N_5545);
xor U5604 (N_5604,N_5516,N_5572);
nand U5605 (N_5605,N_5445,N_5406);
or U5606 (N_5606,N_5528,N_5456);
xor U5607 (N_5607,N_5448,N_5519);
nor U5608 (N_5608,N_5424,N_5587);
or U5609 (N_5609,N_5559,N_5418);
and U5610 (N_5610,N_5506,N_5490);
nor U5611 (N_5611,N_5586,N_5492);
nor U5612 (N_5612,N_5577,N_5440);
or U5613 (N_5613,N_5473,N_5495);
xor U5614 (N_5614,N_5573,N_5557);
nor U5615 (N_5615,N_5449,N_5599);
nor U5616 (N_5616,N_5501,N_5520);
or U5617 (N_5617,N_5512,N_5493);
nor U5618 (N_5618,N_5482,N_5489);
nor U5619 (N_5619,N_5487,N_5517);
and U5620 (N_5620,N_5581,N_5483);
or U5621 (N_5621,N_5560,N_5530);
nor U5622 (N_5622,N_5485,N_5568);
nor U5623 (N_5623,N_5410,N_5542);
nor U5624 (N_5624,N_5514,N_5533);
nand U5625 (N_5625,N_5550,N_5475);
or U5626 (N_5626,N_5423,N_5480);
xor U5627 (N_5627,N_5417,N_5419);
and U5628 (N_5628,N_5434,N_5467);
and U5629 (N_5629,N_5416,N_5428);
and U5630 (N_5630,N_5561,N_5515);
or U5631 (N_5631,N_5579,N_5479);
or U5632 (N_5632,N_5526,N_5567);
xor U5633 (N_5633,N_5458,N_5543);
and U5634 (N_5634,N_5455,N_5405);
nand U5635 (N_5635,N_5409,N_5584);
or U5636 (N_5636,N_5465,N_5529);
nand U5637 (N_5637,N_5548,N_5461);
xnor U5638 (N_5638,N_5429,N_5447);
xor U5639 (N_5639,N_5558,N_5594);
nand U5640 (N_5640,N_5499,N_5498);
xor U5641 (N_5641,N_5537,N_5438);
or U5642 (N_5642,N_5502,N_5566);
nand U5643 (N_5643,N_5415,N_5401);
nor U5644 (N_5644,N_5470,N_5436);
nor U5645 (N_5645,N_5522,N_5532);
or U5646 (N_5646,N_5574,N_5556);
or U5647 (N_5647,N_5582,N_5547);
and U5648 (N_5648,N_5507,N_5544);
xnor U5649 (N_5649,N_5432,N_5598);
or U5650 (N_5650,N_5408,N_5481);
nor U5651 (N_5651,N_5508,N_5403);
xor U5652 (N_5652,N_5518,N_5565);
or U5653 (N_5653,N_5437,N_5576);
nor U5654 (N_5654,N_5484,N_5442);
nand U5655 (N_5655,N_5477,N_5476);
nand U5656 (N_5656,N_5471,N_5412);
and U5657 (N_5657,N_5555,N_5446);
and U5658 (N_5658,N_5564,N_5578);
nor U5659 (N_5659,N_5597,N_5588);
and U5660 (N_5660,N_5504,N_5531);
xor U5661 (N_5661,N_5400,N_5411);
or U5662 (N_5662,N_5500,N_5538);
nand U5663 (N_5663,N_5523,N_5413);
and U5664 (N_5664,N_5402,N_5503);
xor U5665 (N_5665,N_5505,N_5425);
nor U5666 (N_5666,N_5497,N_5536);
nor U5667 (N_5667,N_5596,N_5552);
nor U5668 (N_5668,N_5585,N_5421);
nor U5669 (N_5669,N_5591,N_5422);
xnor U5670 (N_5670,N_5427,N_5433);
xor U5671 (N_5671,N_5541,N_5453);
xnor U5672 (N_5672,N_5589,N_5486);
nor U5673 (N_5673,N_5444,N_5580);
nor U5674 (N_5674,N_5513,N_5464);
or U5675 (N_5675,N_5459,N_5469);
nand U5676 (N_5676,N_5549,N_5540);
xor U5677 (N_5677,N_5491,N_5592);
nor U5678 (N_5678,N_5407,N_5450);
or U5679 (N_5679,N_5539,N_5524);
nor U5680 (N_5680,N_5570,N_5595);
and U5681 (N_5681,N_5474,N_5451);
or U5682 (N_5682,N_5511,N_5457);
nand U5683 (N_5683,N_5554,N_5510);
and U5684 (N_5684,N_5546,N_5466);
nor U5685 (N_5685,N_5509,N_5468);
nand U5686 (N_5686,N_5535,N_5478);
or U5687 (N_5687,N_5553,N_5551);
and U5688 (N_5688,N_5430,N_5431);
xnor U5689 (N_5689,N_5527,N_5404);
xnor U5690 (N_5690,N_5562,N_5441);
or U5691 (N_5691,N_5525,N_5452);
and U5692 (N_5692,N_5420,N_5426);
nor U5693 (N_5693,N_5534,N_5439);
xor U5694 (N_5694,N_5460,N_5496);
nand U5695 (N_5695,N_5435,N_5521);
and U5696 (N_5696,N_5488,N_5563);
nand U5697 (N_5697,N_5571,N_5569);
or U5698 (N_5698,N_5593,N_5463);
or U5699 (N_5699,N_5575,N_5590);
nand U5700 (N_5700,N_5595,N_5448);
or U5701 (N_5701,N_5438,N_5406);
nand U5702 (N_5702,N_5540,N_5467);
and U5703 (N_5703,N_5417,N_5501);
and U5704 (N_5704,N_5498,N_5460);
or U5705 (N_5705,N_5454,N_5474);
and U5706 (N_5706,N_5526,N_5457);
xor U5707 (N_5707,N_5541,N_5428);
and U5708 (N_5708,N_5486,N_5454);
nand U5709 (N_5709,N_5584,N_5504);
or U5710 (N_5710,N_5405,N_5480);
nor U5711 (N_5711,N_5516,N_5450);
nor U5712 (N_5712,N_5558,N_5583);
nand U5713 (N_5713,N_5543,N_5545);
xor U5714 (N_5714,N_5533,N_5537);
nand U5715 (N_5715,N_5422,N_5524);
xor U5716 (N_5716,N_5461,N_5573);
and U5717 (N_5717,N_5416,N_5508);
nand U5718 (N_5718,N_5492,N_5464);
nor U5719 (N_5719,N_5494,N_5507);
nor U5720 (N_5720,N_5479,N_5471);
or U5721 (N_5721,N_5429,N_5478);
xor U5722 (N_5722,N_5507,N_5522);
or U5723 (N_5723,N_5422,N_5435);
or U5724 (N_5724,N_5521,N_5469);
or U5725 (N_5725,N_5568,N_5477);
or U5726 (N_5726,N_5445,N_5572);
nand U5727 (N_5727,N_5547,N_5409);
nor U5728 (N_5728,N_5515,N_5494);
nand U5729 (N_5729,N_5555,N_5586);
and U5730 (N_5730,N_5595,N_5477);
nor U5731 (N_5731,N_5537,N_5597);
and U5732 (N_5732,N_5447,N_5591);
or U5733 (N_5733,N_5473,N_5591);
or U5734 (N_5734,N_5538,N_5512);
and U5735 (N_5735,N_5414,N_5544);
nor U5736 (N_5736,N_5518,N_5526);
and U5737 (N_5737,N_5473,N_5463);
and U5738 (N_5738,N_5530,N_5541);
nor U5739 (N_5739,N_5416,N_5482);
xor U5740 (N_5740,N_5537,N_5433);
or U5741 (N_5741,N_5535,N_5429);
or U5742 (N_5742,N_5466,N_5461);
nor U5743 (N_5743,N_5473,N_5588);
xnor U5744 (N_5744,N_5530,N_5563);
and U5745 (N_5745,N_5580,N_5541);
xnor U5746 (N_5746,N_5578,N_5415);
nand U5747 (N_5747,N_5504,N_5407);
and U5748 (N_5748,N_5593,N_5465);
or U5749 (N_5749,N_5556,N_5533);
or U5750 (N_5750,N_5404,N_5505);
nand U5751 (N_5751,N_5558,N_5587);
and U5752 (N_5752,N_5587,N_5472);
nor U5753 (N_5753,N_5404,N_5461);
or U5754 (N_5754,N_5490,N_5587);
xnor U5755 (N_5755,N_5573,N_5402);
nand U5756 (N_5756,N_5522,N_5418);
and U5757 (N_5757,N_5549,N_5571);
xnor U5758 (N_5758,N_5469,N_5518);
or U5759 (N_5759,N_5523,N_5457);
xor U5760 (N_5760,N_5553,N_5476);
nor U5761 (N_5761,N_5419,N_5544);
or U5762 (N_5762,N_5574,N_5498);
nor U5763 (N_5763,N_5598,N_5596);
or U5764 (N_5764,N_5416,N_5540);
and U5765 (N_5765,N_5573,N_5423);
nand U5766 (N_5766,N_5415,N_5591);
xnor U5767 (N_5767,N_5519,N_5464);
xor U5768 (N_5768,N_5409,N_5493);
nor U5769 (N_5769,N_5479,N_5430);
nor U5770 (N_5770,N_5437,N_5400);
nor U5771 (N_5771,N_5554,N_5405);
nor U5772 (N_5772,N_5455,N_5509);
xor U5773 (N_5773,N_5556,N_5576);
nand U5774 (N_5774,N_5445,N_5463);
nor U5775 (N_5775,N_5531,N_5543);
xnor U5776 (N_5776,N_5515,N_5549);
or U5777 (N_5777,N_5500,N_5543);
or U5778 (N_5778,N_5541,N_5508);
and U5779 (N_5779,N_5500,N_5484);
xnor U5780 (N_5780,N_5437,N_5484);
xnor U5781 (N_5781,N_5555,N_5565);
or U5782 (N_5782,N_5482,N_5408);
nor U5783 (N_5783,N_5573,N_5536);
and U5784 (N_5784,N_5447,N_5522);
or U5785 (N_5785,N_5482,N_5529);
xnor U5786 (N_5786,N_5508,N_5423);
nand U5787 (N_5787,N_5505,N_5533);
and U5788 (N_5788,N_5463,N_5542);
nor U5789 (N_5789,N_5442,N_5448);
xnor U5790 (N_5790,N_5513,N_5488);
and U5791 (N_5791,N_5427,N_5594);
nand U5792 (N_5792,N_5473,N_5449);
nand U5793 (N_5793,N_5525,N_5421);
or U5794 (N_5794,N_5408,N_5458);
and U5795 (N_5795,N_5495,N_5445);
xnor U5796 (N_5796,N_5527,N_5414);
nor U5797 (N_5797,N_5558,N_5512);
and U5798 (N_5798,N_5562,N_5554);
nand U5799 (N_5799,N_5549,N_5403);
xor U5800 (N_5800,N_5686,N_5661);
xor U5801 (N_5801,N_5743,N_5723);
and U5802 (N_5802,N_5621,N_5649);
nand U5803 (N_5803,N_5745,N_5768);
nand U5804 (N_5804,N_5642,N_5648);
nor U5805 (N_5805,N_5662,N_5641);
nor U5806 (N_5806,N_5714,N_5780);
nand U5807 (N_5807,N_5630,N_5611);
or U5808 (N_5808,N_5706,N_5719);
or U5809 (N_5809,N_5756,N_5668);
nand U5810 (N_5810,N_5628,N_5610);
and U5811 (N_5811,N_5680,N_5626);
nand U5812 (N_5812,N_5620,N_5650);
or U5813 (N_5813,N_5637,N_5689);
nand U5814 (N_5814,N_5785,N_5761);
nor U5815 (N_5815,N_5713,N_5767);
nand U5816 (N_5816,N_5683,N_5773);
or U5817 (N_5817,N_5770,N_5658);
xnor U5818 (N_5818,N_5652,N_5685);
and U5819 (N_5819,N_5734,N_5754);
nor U5820 (N_5820,N_5678,N_5697);
or U5821 (N_5821,N_5640,N_5715);
nor U5822 (N_5822,N_5669,N_5794);
and U5823 (N_5823,N_5736,N_5717);
nand U5824 (N_5824,N_5732,N_5791);
nand U5825 (N_5825,N_5744,N_5741);
and U5826 (N_5826,N_5607,N_5722);
nor U5827 (N_5827,N_5625,N_5639);
nand U5828 (N_5828,N_5646,N_5727);
or U5829 (N_5829,N_5696,N_5692);
nand U5830 (N_5830,N_5733,N_5600);
nand U5831 (N_5831,N_5796,N_5687);
nor U5832 (N_5832,N_5726,N_5693);
xor U5833 (N_5833,N_5790,N_5647);
and U5834 (N_5834,N_5704,N_5694);
nor U5835 (N_5835,N_5615,N_5627);
nor U5836 (N_5836,N_5663,N_5731);
nor U5837 (N_5837,N_5645,N_5720);
xor U5838 (N_5838,N_5673,N_5749);
xor U5839 (N_5839,N_5711,N_5608);
xnor U5840 (N_5840,N_5624,N_5769);
nor U5841 (N_5841,N_5721,N_5710);
nand U5842 (N_5842,N_5609,N_5783);
xnor U5843 (N_5843,N_5701,N_5671);
nor U5844 (N_5844,N_5777,N_5602);
nand U5845 (N_5845,N_5651,N_5670);
nor U5846 (N_5846,N_5656,N_5739);
and U5847 (N_5847,N_5665,N_5632);
nor U5848 (N_5848,N_5601,N_5771);
nor U5849 (N_5849,N_5753,N_5677);
and U5850 (N_5850,N_5666,N_5638);
or U5851 (N_5851,N_5606,N_5622);
nand U5852 (N_5852,N_5654,N_5707);
xor U5853 (N_5853,N_5763,N_5792);
nor U5854 (N_5854,N_5629,N_5682);
xor U5855 (N_5855,N_5784,N_5764);
or U5856 (N_5856,N_5644,N_5667);
nand U5857 (N_5857,N_5603,N_5725);
xor U5858 (N_5858,N_5766,N_5737);
xor U5859 (N_5859,N_5798,N_5674);
or U5860 (N_5860,N_5708,N_5765);
xnor U5861 (N_5861,N_5635,N_5659);
nor U5862 (N_5862,N_5728,N_5762);
nand U5863 (N_5863,N_5688,N_5613);
and U5864 (N_5864,N_5679,N_5695);
and U5865 (N_5865,N_5786,N_5752);
nand U5866 (N_5866,N_5740,N_5779);
xor U5867 (N_5867,N_5758,N_5718);
or U5868 (N_5868,N_5748,N_5604);
xor U5869 (N_5869,N_5699,N_5657);
and U5870 (N_5870,N_5788,N_5757);
nor U5871 (N_5871,N_5774,N_5623);
and U5872 (N_5872,N_5747,N_5681);
and U5873 (N_5873,N_5690,N_5729);
and U5874 (N_5874,N_5751,N_5705);
nand U5875 (N_5875,N_5775,N_5614);
or U5876 (N_5876,N_5776,N_5793);
or U5877 (N_5877,N_5612,N_5698);
nor U5878 (N_5878,N_5619,N_5660);
and U5879 (N_5879,N_5738,N_5617);
nand U5880 (N_5880,N_5760,N_5746);
or U5881 (N_5881,N_5634,N_5799);
and U5882 (N_5882,N_5709,N_5675);
xnor U5883 (N_5883,N_5605,N_5618);
nor U5884 (N_5884,N_5789,N_5724);
and U5885 (N_5885,N_5702,N_5742);
nand U5886 (N_5886,N_5655,N_5664);
nor U5887 (N_5887,N_5616,N_5703);
or U5888 (N_5888,N_5750,N_5672);
nor U5889 (N_5889,N_5730,N_5631);
xor U5890 (N_5890,N_5782,N_5781);
xnor U5891 (N_5891,N_5778,N_5735);
nor U5892 (N_5892,N_5712,N_5636);
and U5893 (N_5893,N_5797,N_5691);
xnor U5894 (N_5894,N_5676,N_5759);
xnor U5895 (N_5895,N_5787,N_5795);
or U5896 (N_5896,N_5755,N_5643);
and U5897 (N_5897,N_5700,N_5684);
or U5898 (N_5898,N_5772,N_5716);
and U5899 (N_5899,N_5633,N_5653);
and U5900 (N_5900,N_5691,N_5739);
and U5901 (N_5901,N_5717,N_5648);
nand U5902 (N_5902,N_5727,N_5653);
nor U5903 (N_5903,N_5630,N_5704);
nor U5904 (N_5904,N_5787,N_5663);
or U5905 (N_5905,N_5727,N_5713);
nand U5906 (N_5906,N_5737,N_5775);
nor U5907 (N_5907,N_5653,N_5664);
or U5908 (N_5908,N_5644,N_5614);
nor U5909 (N_5909,N_5620,N_5677);
nand U5910 (N_5910,N_5616,N_5630);
or U5911 (N_5911,N_5764,N_5620);
xor U5912 (N_5912,N_5774,N_5601);
and U5913 (N_5913,N_5675,N_5714);
or U5914 (N_5914,N_5627,N_5606);
or U5915 (N_5915,N_5723,N_5670);
nand U5916 (N_5916,N_5683,N_5664);
or U5917 (N_5917,N_5728,N_5611);
xor U5918 (N_5918,N_5743,N_5786);
xor U5919 (N_5919,N_5634,N_5603);
nand U5920 (N_5920,N_5671,N_5727);
nand U5921 (N_5921,N_5665,N_5790);
xnor U5922 (N_5922,N_5680,N_5682);
nand U5923 (N_5923,N_5778,N_5793);
and U5924 (N_5924,N_5652,N_5720);
nor U5925 (N_5925,N_5771,N_5759);
nor U5926 (N_5926,N_5698,N_5610);
nor U5927 (N_5927,N_5627,N_5766);
xor U5928 (N_5928,N_5782,N_5723);
nor U5929 (N_5929,N_5768,N_5644);
nor U5930 (N_5930,N_5722,N_5785);
nor U5931 (N_5931,N_5642,N_5733);
nor U5932 (N_5932,N_5728,N_5610);
and U5933 (N_5933,N_5675,N_5755);
nand U5934 (N_5934,N_5636,N_5615);
nor U5935 (N_5935,N_5704,N_5635);
and U5936 (N_5936,N_5740,N_5795);
and U5937 (N_5937,N_5640,N_5788);
and U5938 (N_5938,N_5657,N_5719);
or U5939 (N_5939,N_5619,N_5764);
nand U5940 (N_5940,N_5647,N_5769);
nor U5941 (N_5941,N_5620,N_5664);
xor U5942 (N_5942,N_5719,N_5603);
nor U5943 (N_5943,N_5745,N_5788);
nor U5944 (N_5944,N_5700,N_5656);
and U5945 (N_5945,N_5687,N_5717);
nand U5946 (N_5946,N_5667,N_5688);
or U5947 (N_5947,N_5638,N_5793);
or U5948 (N_5948,N_5615,N_5754);
or U5949 (N_5949,N_5675,N_5797);
or U5950 (N_5950,N_5616,N_5695);
xor U5951 (N_5951,N_5620,N_5767);
xor U5952 (N_5952,N_5626,N_5729);
nand U5953 (N_5953,N_5757,N_5684);
and U5954 (N_5954,N_5759,N_5711);
nor U5955 (N_5955,N_5719,N_5628);
and U5956 (N_5956,N_5795,N_5603);
and U5957 (N_5957,N_5634,N_5702);
xnor U5958 (N_5958,N_5738,N_5780);
nor U5959 (N_5959,N_5702,N_5632);
nor U5960 (N_5960,N_5638,N_5655);
nand U5961 (N_5961,N_5657,N_5728);
xnor U5962 (N_5962,N_5744,N_5798);
or U5963 (N_5963,N_5787,N_5707);
xnor U5964 (N_5964,N_5764,N_5660);
nand U5965 (N_5965,N_5796,N_5740);
and U5966 (N_5966,N_5689,N_5639);
xnor U5967 (N_5967,N_5792,N_5614);
xor U5968 (N_5968,N_5705,N_5770);
nand U5969 (N_5969,N_5637,N_5711);
nand U5970 (N_5970,N_5667,N_5640);
nor U5971 (N_5971,N_5600,N_5666);
and U5972 (N_5972,N_5632,N_5794);
or U5973 (N_5973,N_5707,N_5788);
and U5974 (N_5974,N_5648,N_5702);
or U5975 (N_5975,N_5735,N_5737);
and U5976 (N_5976,N_5603,N_5665);
or U5977 (N_5977,N_5642,N_5600);
xnor U5978 (N_5978,N_5659,N_5728);
nand U5979 (N_5979,N_5754,N_5787);
xnor U5980 (N_5980,N_5720,N_5713);
nor U5981 (N_5981,N_5611,N_5696);
and U5982 (N_5982,N_5669,N_5673);
or U5983 (N_5983,N_5701,N_5774);
nor U5984 (N_5984,N_5610,N_5629);
nand U5985 (N_5985,N_5746,N_5664);
or U5986 (N_5986,N_5680,N_5764);
xnor U5987 (N_5987,N_5650,N_5623);
xor U5988 (N_5988,N_5756,N_5798);
xnor U5989 (N_5989,N_5793,N_5633);
and U5990 (N_5990,N_5707,N_5715);
nand U5991 (N_5991,N_5672,N_5653);
or U5992 (N_5992,N_5673,N_5722);
nand U5993 (N_5993,N_5688,N_5676);
nand U5994 (N_5994,N_5709,N_5652);
nor U5995 (N_5995,N_5746,N_5786);
nand U5996 (N_5996,N_5643,N_5765);
nor U5997 (N_5997,N_5715,N_5782);
xor U5998 (N_5998,N_5659,N_5796);
xor U5999 (N_5999,N_5713,N_5635);
or U6000 (N_6000,N_5965,N_5899);
nor U6001 (N_6001,N_5919,N_5912);
or U6002 (N_6002,N_5944,N_5857);
or U6003 (N_6003,N_5847,N_5973);
xor U6004 (N_6004,N_5822,N_5892);
or U6005 (N_6005,N_5909,N_5924);
and U6006 (N_6006,N_5981,N_5947);
nand U6007 (N_6007,N_5861,N_5957);
nand U6008 (N_6008,N_5879,N_5978);
nor U6009 (N_6009,N_5935,N_5870);
nor U6010 (N_6010,N_5926,N_5827);
nor U6011 (N_6011,N_5936,N_5998);
and U6012 (N_6012,N_5910,N_5969);
xor U6013 (N_6013,N_5887,N_5888);
xnor U6014 (N_6014,N_5992,N_5880);
or U6015 (N_6015,N_5933,N_5873);
or U6016 (N_6016,N_5840,N_5946);
nand U6017 (N_6017,N_5803,N_5804);
or U6018 (N_6018,N_5882,N_5913);
and U6019 (N_6019,N_5982,N_5930);
and U6020 (N_6020,N_5956,N_5963);
or U6021 (N_6021,N_5989,N_5846);
and U6022 (N_6022,N_5921,N_5825);
xor U6023 (N_6023,N_5897,N_5810);
or U6024 (N_6024,N_5995,N_5948);
and U6025 (N_6025,N_5971,N_5937);
nor U6026 (N_6026,N_5865,N_5968);
xor U6027 (N_6027,N_5871,N_5869);
xnor U6028 (N_6028,N_5943,N_5829);
or U6029 (N_6029,N_5811,N_5920);
and U6030 (N_6030,N_5986,N_5934);
or U6031 (N_6031,N_5806,N_5862);
nor U6032 (N_6032,N_5818,N_5979);
nand U6033 (N_6033,N_5851,N_5849);
xor U6034 (N_6034,N_5884,N_5848);
or U6035 (N_6035,N_5940,N_5839);
nand U6036 (N_6036,N_5842,N_5864);
nor U6037 (N_6037,N_5801,N_5898);
or U6038 (N_6038,N_5994,N_5895);
and U6039 (N_6039,N_5923,N_5860);
nor U6040 (N_6040,N_5931,N_5925);
and U6041 (N_6041,N_5932,N_5966);
nor U6042 (N_6042,N_5807,N_5900);
xnor U6043 (N_6043,N_5875,N_5872);
or U6044 (N_6044,N_5881,N_5830);
nand U6045 (N_6045,N_5955,N_5843);
and U6046 (N_6046,N_5904,N_5855);
xnor U6047 (N_6047,N_5821,N_5903);
nor U6048 (N_6048,N_5951,N_5988);
xor U6049 (N_6049,N_5826,N_5853);
and U6050 (N_6050,N_5908,N_5834);
or U6051 (N_6051,N_5812,N_5967);
or U6052 (N_6052,N_5852,N_5841);
nand U6053 (N_6053,N_5914,N_5954);
and U6054 (N_6054,N_5885,N_5958);
nor U6055 (N_6055,N_5858,N_5942);
or U6056 (N_6056,N_5817,N_5962);
xnor U6057 (N_6057,N_5809,N_5927);
xnor U6058 (N_6058,N_5859,N_5990);
nor U6059 (N_6059,N_5844,N_5867);
and U6060 (N_6060,N_5953,N_5876);
and U6061 (N_6061,N_5993,N_5974);
or U6062 (N_6062,N_5964,N_5906);
nor U6063 (N_6063,N_5959,N_5883);
or U6064 (N_6064,N_5877,N_5890);
nor U6065 (N_6065,N_5894,N_5970);
nand U6066 (N_6066,N_5836,N_5939);
xor U6067 (N_6067,N_5866,N_5854);
nand U6068 (N_6068,N_5991,N_5893);
or U6069 (N_6069,N_5863,N_5975);
xnor U6070 (N_6070,N_5949,N_5985);
xor U6071 (N_6071,N_5952,N_5916);
and U6072 (N_6072,N_5878,N_5902);
or U6073 (N_6073,N_5838,N_5960);
xnor U6074 (N_6074,N_5856,N_5805);
xor U6075 (N_6075,N_5996,N_5845);
xor U6076 (N_6076,N_5983,N_5980);
and U6077 (N_6077,N_5833,N_5972);
and U6078 (N_6078,N_5929,N_5945);
and U6079 (N_6079,N_5907,N_5961);
nand U6080 (N_6080,N_5901,N_5891);
or U6081 (N_6081,N_5874,N_5823);
and U6082 (N_6082,N_5820,N_5828);
nand U6083 (N_6083,N_5889,N_5950);
or U6084 (N_6084,N_5819,N_5886);
and U6085 (N_6085,N_5915,N_5917);
xor U6086 (N_6086,N_5832,N_5850);
and U6087 (N_6087,N_5835,N_5918);
and U6088 (N_6088,N_5922,N_5941);
or U6089 (N_6089,N_5977,N_5808);
nor U6090 (N_6090,N_5905,N_5976);
or U6091 (N_6091,N_5816,N_5802);
nand U6092 (N_6092,N_5831,N_5999);
or U6093 (N_6093,N_5813,N_5987);
nor U6094 (N_6094,N_5911,N_5824);
xor U6095 (N_6095,N_5928,N_5868);
nor U6096 (N_6096,N_5997,N_5938);
and U6097 (N_6097,N_5837,N_5896);
xor U6098 (N_6098,N_5800,N_5984);
nand U6099 (N_6099,N_5814,N_5815);
and U6100 (N_6100,N_5972,N_5872);
nor U6101 (N_6101,N_5947,N_5931);
or U6102 (N_6102,N_5837,N_5827);
and U6103 (N_6103,N_5954,N_5904);
nor U6104 (N_6104,N_5857,N_5886);
nor U6105 (N_6105,N_5804,N_5881);
nand U6106 (N_6106,N_5822,N_5856);
and U6107 (N_6107,N_5950,N_5958);
and U6108 (N_6108,N_5832,N_5882);
nor U6109 (N_6109,N_5875,N_5881);
nor U6110 (N_6110,N_5886,N_5885);
nor U6111 (N_6111,N_5936,N_5907);
and U6112 (N_6112,N_5865,N_5992);
xor U6113 (N_6113,N_5890,N_5809);
and U6114 (N_6114,N_5825,N_5838);
xor U6115 (N_6115,N_5888,N_5850);
xnor U6116 (N_6116,N_5829,N_5854);
or U6117 (N_6117,N_5929,N_5965);
nand U6118 (N_6118,N_5953,N_5864);
or U6119 (N_6119,N_5973,N_5855);
or U6120 (N_6120,N_5979,N_5895);
xor U6121 (N_6121,N_5862,N_5947);
or U6122 (N_6122,N_5819,N_5851);
xnor U6123 (N_6123,N_5937,N_5840);
nor U6124 (N_6124,N_5958,N_5938);
or U6125 (N_6125,N_5885,N_5976);
nor U6126 (N_6126,N_5853,N_5805);
or U6127 (N_6127,N_5921,N_5850);
nor U6128 (N_6128,N_5896,N_5855);
xnor U6129 (N_6129,N_5932,N_5885);
and U6130 (N_6130,N_5966,N_5934);
nand U6131 (N_6131,N_5955,N_5911);
xor U6132 (N_6132,N_5825,N_5947);
xnor U6133 (N_6133,N_5981,N_5942);
nor U6134 (N_6134,N_5812,N_5938);
and U6135 (N_6135,N_5883,N_5963);
or U6136 (N_6136,N_5930,N_5968);
nand U6137 (N_6137,N_5821,N_5863);
nor U6138 (N_6138,N_5876,N_5911);
or U6139 (N_6139,N_5942,N_5967);
nand U6140 (N_6140,N_5951,N_5925);
and U6141 (N_6141,N_5953,N_5841);
or U6142 (N_6142,N_5999,N_5818);
xnor U6143 (N_6143,N_5882,N_5928);
xnor U6144 (N_6144,N_5899,N_5902);
nor U6145 (N_6145,N_5915,N_5908);
nor U6146 (N_6146,N_5898,N_5873);
nand U6147 (N_6147,N_5832,N_5955);
or U6148 (N_6148,N_5916,N_5875);
xor U6149 (N_6149,N_5898,N_5945);
nor U6150 (N_6150,N_5845,N_5863);
nor U6151 (N_6151,N_5896,N_5922);
xnor U6152 (N_6152,N_5934,N_5809);
xor U6153 (N_6153,N_5817,N_5882);
nand U6154 (N_6154,N_5986,N_5831);
nand U6155 (N_6155,N_5901,N_5949);
or U6156 (N_6156,N_5994,N_5837);
nand U6157 (N_6157,N_5901,N_5945);
nor U6158 (N_6158,N_5932,N_5880);
nor U6159 (N_6159,N_5837,N_5976);
nand U6160 (N_6160,N_5933,N_5805);
nand U6161 (N_6161,N_5890,N_5938);
and U6162 (N_6162,N_5974,N_5856);
or U6163 (N_6163,N_5859,N_5962);
nor U6164 (N_6164,N_5871,N_5986);
xor U6165 (N_6165,N_5872,N_5870);
nand U6166 (N_6166,N_5818,N_5953);
nand U6167 (N_6167,N_5812,N_5979);
or U6168 (N_6168,N_5957,N_5982);
or U6169 (N_6169,N_5805,N_5904);
or U6170 (N_6170,N_5932,N_5857);
and U6171 (N_6171,N_5804,N_5897);
or U6172 (N_6172,N_5976,N_5981);
or U6173 (N_6173,N_5865,N_5985);
xnor U6174 (N_6174,N_5837,N_5901);
xor U6175 (N_6175,N_5949,N_5988);
or U6176 (N_6176,N_5867,N_5802);
and U6177 (N_6177,N_5917,N_5828);
or U6178 (N_6178,N_5848,N_5894);
and U6179 (N_6179,N_5982,N_5873);
xor U6180 (N_6180,N_5941,N_5850);
or U6181 (N_6181,N_5827,N_5953);
and U6182 (N_6182,N_5890,N_5947);
or U6183 (N_6183,N_5801,N_5844);
and U6184 (N_6184,N_5864,N_5936);
nand U6185 (N_6185,N_5811,N_5861);
nand U6186 (N_6186,N_5967,N_5869);
xnor U6187 (N_6187,N_5966,N_5892);
or U6188 (N_6188,N_5932,N_5817);
nand U6189 (N_6189,N_5915,N_5965);
nor U6190 (N_6190,N_5947,N_5823);
and U6191 (N_6191,N_5812,N_5874);
or U6192 (N_6192,N_5809,N_5824);
or U6193 (N_6193,N_5859,N_5898);
xnor U6194 (N_6194,N_5907,N_5849);
or U6195 (N_6195,N_5807,N_5929);
xor U6196 (N_6196,N_5999,N_5867);
and U6197 (N_6197,N_5884,N_5814);
or U6198 (N_6198,N_5917,N_5895);
and U6199 (N_6199,N_5823,N_5828);
and U6200 (N_6200,N_6040,N_6032);
nand U6201 (N_6201,N_6077,N_6172);
or U6202 (N_6202,N_6076,N_6117);
nor U6203 (N_6203,N_6183,N_6021);
or U6204 (N_6204,N_6069,N_6163);
xor U6205 (N_6205,N_6093,N_6050);
or U6206 (N_6206,N_6031,N_6166);
xor U6207 (N_6207,N_6131,N_6136);
or U6208 (N_6208,N_6177,N_6044);
nor U6209 (N_6209,N_6068,N_6070);
and U6210 (N_6210,N_6173,N_6062);
nand U6211 (N_6211,N_6162,N_6009);
nor U6212 (N_6212,N_6164,N_6098);
or U6213 (N_6213,N_6128,N_6022);
and U6214 (N_6214,N_6147,N_6013);
nor U6215 (N_6215,N_6006,N_6111);
nand U6216 (N_6216,N_6081,N_6198);
nand U6217 (N_6217,N_6135,N_6138);
nand U6218 (N_6218,N_6058,N_6012);
and U6219 (N_6219,N_6127,N_6185);
xor U6220 (N_6220,N_6046,N_6097);
and U6221 (N_6221,N_6010,N_6179);
or U6222 (N_6222,N_6158,N_6026);
xor U6223 (N_6223,N_6197,N_6051);
or U6224 (N_6224,N_6186,N_6004);
nor U6225 (N_6225,N_6096,N_6000);
xor U6226 (N_6226,N_6168,N_6153);
and U6227 (N_6227,N_6084,N_6104);
xnor U6228 (N_6228,N_6071,N_6122);
nand U6229 (N_6229,N_6079,N_6165);
nor U6230 (N_6230,N_6073,N_6120);
nand U6231 (N_6231,N_6118,N_6132);
or U6232 (N_6232,N_6015,N_6041);
or U6233 (N_6233,N_6149,N_6099);
nand U6234 (N_6234,N_6140,N_6161);
and U6235 (N_6235,N_6049,N_6123);
nor U6236 (N_6236,N_6059,N_6055);
xor U6237 (N_6237,N_6142,N_6089);
or U6238 (N_6238,N_6083,N_6060);
xor U6239 (N_6239,N_6126,N_6189);
nor U6240 (N_6240,N_6190,N_6087);
or U6241 (N_6241,N_6152,N_6029);
nand U6242 (N_6242,N_6092,N_6106);
xor U6243 (N_6243,N_6066,N_6052);
or U6244 (N_6244,N_6074,N_6056);
or U6245 (N_6245,N_6160,N_6078);
xor U6246 (N_6246,N_6105,N_6180);
nand U6247 (N_6247,N_6003,N_6144);
and U6248 (N_6248,N_6024,N_6016);
nand U6249 (N_6249,N_6054,N_6080);
and U6250 (N_6250,N_6005,N_6178);
nor U6251 (N_6251,N_6108,N_6171);
or U6252 (N_6252,N_6036,N_6038);
nor U6253 (N_6253,N_6184,N_6167);
and U6254 (N_6254,N_6170,N_6039);
or U6255 (N_6255,N_6008,N_6125);
or U6256 (N_6256,N_6001,N_6192);
and U6257 (N_6257,N_6134,N_6042);
and U6258 (N_6258,N_6035,N_6034);
nand U6259 (N_6259,N_6033,N_6103);
xnor U6260 (N_6260,N_6176,N_6191);
and U6261 (N_6261,N_6182,N_6061);
nand U6262 (N_6262,N_6095,N_6114);
nand U6263 (N_6263,N_6159,N_6150);
or U6264 (N_6264,N_6057,N_6094);
xnor U6265 (N_6265,N_6143,N_6157);
and U6266 (N_6266,N_6011,N_6017);
and U6267 (N_6267,N_6133,N_6027);
nand U6268 (N_6268,N_6072,N_6102);
nand U6269 (N_6269,N_6018,N_6063);
and U6270 (N_6270,N_6043,N_6065);
nand U6271 (N_6271,N_6116,N_6047);
nand U6272 (N_6272,N_6086,N_6124);
nand U6273 (N_6273,N_6045,N_6019);
xnor U6274 (N_6274,N_6002,N_6188);
or U6275 (N_6275,N_6181,N_6129);
and U6276 (N_6276,N_6139,N_6107);
xor U6277 (N_6277,N_6053,N_6175);
xnor U6278 (N_6278,N_6085,N_6151);
xnor U6279 (N_6279,N_6014,N_6148);
nand U6280 (N_6280,N_6156,N_6028);
xor U6281 (N_6281,N_6193,N_6025);
nor U6282 (N_6282,N_6199,N_6115);
and U6283 (N_6283,N_6090,N_6048);
or U6284 (N_6284,N_6110,N_6169);
or U6285 (N_6285,N_6091,N_6088);
xnor U6286 (N_6286,N_6112,N_6100);
xor U6287 (N_6287,N_6155,N_6082);
or U6288 (N_6288,N_6067,N_6037);
or U6289 (N_6289,N_6145,N_6030);
and U6290 (N_6290,N_6121,N_6075);
nor U6291 (N_6291,N_6023,N_6113);
nand U6292 (N_6292,N_6154,N_6146);
nor U6293 (N_6293,N_6109,N_6141);
nor U6294 (N_6294,N_6020,N_6119);
or U6295 (N_6295,N_6101,N_6174);
xnor U6296 (N_6296,N_6137,N_6194);
and U6297 (N_6297,N_6007,N_6196);
and U6298 (N_6298,N_6064,N_6187);
nor U6299 (N_6299,N_6130,N_6195);
or U6300 (N_6300,N_6103,N_6156);
or U6301 (N_6301,N_6024,N_6094);
and U6302 (N_6302,N_6177,N_6066);
or U6303 (N_6303,N_6153,N_6066);
or U6304 (N_6304,N_6139,N_6136);
nand U6305 (N_6305,N_6076,N_6099);
or U6306 (N_6306,N_6137,N_6044);
nor U6307 (N_6307,N_6070,N_6134);
and U6308 (N_6308,N_6108,N_6169);
nand U6309 (N_6309,N_6007,N_6025);
nand U6310 (N_6310,N_6157,N_6102);
nor U6311 (N_6311,N_6145,N_6029);
xnor U6312 (N_6312,N_6030,N_6017);
nand U6313 (N_6313,N_6113,N_6021);
or U6314 (N_6314,N_6098,N_6199);
xnor U6315 (N_6315,N_6061,N_6090);
and U6316 (N_6316,N_6082,N_6190);
xor U6317 (N_6317,N_6038,N_6195);
xor U6318 (N_6318,N_6101,N_6091);
nor U6319 (N_6319,N_6062,N_6013);
nand U6320 (N_6320,N_6029,N_6086);
nand U6321 (N_6321,N_6157,N_6035);
nor U6322 (N_6322,N_6129,N_6029);
and U6323 (N_6323,N_6041,N_6191);
nor U6324 (N_6324,N_6071,N_6037);
xnor U6325 (N_6325,N_6113,N_6135);
and U6326 (N_6326,N_6110,N_6148);
xnor U6327 (N_6327,N_6109,N_6179);
and U6328 (N_6328,N_6140,N_6019);
xnor U6329 (N_6329,N_6154,N_6047);
nand U6330 (N_6330,N_6137,N_6066);
nor U6331 (N_6331,N_6175,N_6184);
nand U6332 (N_6332,N_6095,N_6002);
or U6333 (N_6333,N_6173,N_6070);
and U6334 (N_6334,N_6058,N_6074);
nand U6335 (N_6335,N_6133,N_6110);
nand U6336 (N_6336,N_6104,N_6158);
xnor U6337 (N_6337,N_6134,N_6114);
or U6338 (N_6338,N_6056,N_6053);
and U6339 (N_6339,N_6020,N_6133);
and U6340 (N_6340,N_6136,N_6151);
and U6341 (N_6341,N_6089,N_6155);
nand U6342 (N_6342,N_6000,N_6035);
nor U6343 (N_6343,N_6124,N_6181);
xnor U6344 (N_6344,N_6016,N_6015);
nor U6345 (N_6345,N_6071,N_6115);
nor U6346 (N_6346,N_6024,N_6082);
and U6347 (N_6347,N_6186,N_6129);
nor U6348 (N_6348,N_6170,N_6087);
or U6349 (N_6349,N_6134,N_6181);
or U6350 (N_6350,N_6199,N_6134);
nor U6351 (N_6351,N_6013,N_6150);
nor U6352 (N_6352,N_6199,N_6192);
and U6353 (N_6353,N_6077,N_6127);
nand U6354 (N_6354,N_6159,N_6118);
xor U6355 (N_6355,N_6171,N_6098);
nand U6356 (N_6356,N_6104,N_6188);
and U6357 (N_6357,N_6125,N_6070);
nor U6358 (N_6358,N_6044,N_6168);
or U6359 (N_6359,N_6198,N_6129);
xor U6360 (N_6360,N_6130,N_6156);
and U6361 (N_6361,N_6032,N_6039);
xnor U6362 (N_6362,N_6006,N_6177);
or U6363 (N_6363,N_6025,N_6113);
nand U6364 (N_6364,N_6033,N_6080);
xor U6365 (N_6365,N_6085,N_6090);
nor U6366 (N_6366,N_6193,N_6185);
xor U6367 (N_6367,N_6168,N_6183);
and U6368 (N_6368,N_6171,N_6009);
nand U6369 (N_6369,N_6158,N_6144);
nand U6370 (N_6370,N_6122,N_6194);
xor U6371 (N_6371,N_6024,N_6112);
nand U6372 (N_6372,N_6198,N_6122);
or U6373 (N_6373,N_6159,N_6035);
nor U6374 (N_6374,N_6187,N_6000);
or U6375 (N_6375,N_6063,N_6108);
nor U6376 (N_6376,N_6180,N_6133);
xnor U6377 (N_6377,N_6106,N_6143);
or U6378 (N_6378,N_6041,N_6164);
xor U6379 (N_6379,N_6136,N_6197);
and U6380 (N_6380,N_6004,N_6074);
nand U6381 (N_6381,N_6152,N_6190);
nand U6382 (N_6382,N_6020,N_6123);
nand U6383 (N_6383,N_6050,N_6060);
or U6384 (N_6384,N_6162,N_6093);
and U6385 (N_6385,N_6097,N_6064);
nor U6386 (N_6386,N_6082,N_6021);
nand U6387 (N_6387,N_6160,N_6196);
or U6388 (N_6388,N_6124,N_6083);
or U6389 (N_6389,N_6060,N_6195);
and U6390 (N_6390,N_6168,N_6029);
or U6391 (N_6391,N_6043,N_6057);
and U6392 (N_6392,N_6023,N_6160);
or U6393 (N_6393,N_6165,N_6029);
nor U6394 (N_6394,N_6071,N_6055);
and U6395 (N_6395,N_6198,N_6152);
nand U6396 (N_6396,N_6101,N_6181);
and U6397 (N_6397,N_6149,N_6137);
xor U6398 (N_6398,N_6043,N_6108);
and U6399 (N_6399,N_6100,N_6095);
or U6400 (N_6400,N_6257,N_6280);
and U6401 (N_6401,N_6259,N_6308);
nand U6402 (N_6402,N_6311,N_6231);
and U6403 (N_6403,N_6247,N_6254);
nand U6404 (N_6404,N_6300,N_6301);
and U6405 (N_6405,N_6314,N_6356);
nor U6406 (N_6406,N_6232,N_6249);
or U6407 (N_6407,N_6267,N_6317);
nor U6408 (N_6408,N_6378,N_6335);
nand U6409 (N_6409,N_6395,N_6226);
or U6410 (N_6410,N_6384,N_6228);
or U6411 (N_6411,N_6273,N_6253);
xor U6412 (N_6412,N_6270,N_6292);
xnor U6413 (N_6413,N_6385,N_6203);
xnor U6414 (N_6414,N_6318,N_6245);
nand U6415 (N_6415,N_6398,N_6397);
xor U6416 (N_6416,N_6305,N_6279);
nor U6417 (N_6417,N_6227,N_6334);
xor U6418 (N_6418,N_6342,N_6368);
nand U6419 (N_6419,N_6216,N_6269);
and U6420 (N_6420,N_6331,N_6348);
and U6421 (N_6421,N_6307,N_6213);
or U6422 (N_6422,N_6241,N_6258);
xnor U6423 (N_6423,N_6202,N_6392);
xnor U6424 (N_6424,N_6353,N_6322);
nor U6425 (N_6425,N_6239,N_6256);
nand U6426 (N_6426,N_6349,N_6380);
xnor U6427 (N_6427,N_6347,N_6362);
and U6428 (N_6428,N_6338,N_6373);
xnor U6429 (N_6429,N_6360,N_6211);
nand U6430 (N_6430,N_6350,N_6387);
and U6431 (N_6431,N_6248,N_6365);
or U6432 (N_6432,N_6371,N_6265);
or U6433 (N_6433,N_6215,N_6312);
nand U6434 (N_6434,N_6277,N_6382);
nand U6435 (N_6435,N_6286,N_6386);
or U6436 (N_6436,N_6251,N_6323);
and U6437 (N_6437,N_6377,N_6274);
or U6438 (N_6438,N_6275,N_6313);
xor U6439 (N_6439,N_6246,N_6341);
xor U6440 (N_6440,N_6363,N_6324);
nor U6441 (N_6441,N_6304,N_6271);
xor U6442 (N_6442,N_6302,N_6396);
xor U6443 (N_6443,N_6326,N_6372);
nand U6444 (N_6444,N_6358,N_6221);
xor U6445 (N_6445,N_6238,N_6242);
xnor U6446 (N_6446,N_6381,N_6220);
nor U6447 (N_6447,N_6264,N_6357);
and U6448 (N_6448,N_6268,N_6388);
nor U6449 (N_6449,N_6339,N_6272);
nand U6450 (N_6450,N_6329,N_6336);
and U6451 (N_6451,N_6320,N_6235);
or U6452 (N_6452,N_6315,N_6252);
or U6453 (N_6453,N_6306,N_6205);
or U6454 (N_6454,N_6343,N_6370);
and U6455 (N_6455,N_6303,N_6207);
or U6456 (N_6456,N_6288,N_6218);
xnor U6457 (N_6457,N_6376,N_6325);
xor U6458 (N_6458,N_6204,N_6255);
and U6459 (N_6459,N_6262,N_6355);
and U6460 (N_6460,N_6332,N_6345);
nand U6461 (N_6461,N_6276,N_6217);
nand U6462 (N_6462,N_6285,N_6240);
nand U6463 (N_6463,N_6293,N_6209);
and U6464 (N_6464,N_6354,N_6224);
nand U6465 (N_6465,N_6310,N_6237);
xor U6466 (N_6466,N_6399,N_6290);
nor U6467 (N_6467,N_6321,N_6250);
or U6468 (N_6468,N_6340,N_6201);
nor U6469 (N_6469,N_6236,N_6208);
and U6470 (N_6470,N_6351,N_6243);
xor U6471 (N_6471,N_6244,N_6346);
or U6472 (N_6472,N_6281,N_6219);
and U6473 (N_6473,N_6291,N_6352);
nor U6474 (N_6474,N_6327,N_6223);
xor U6475 (N_6475,N_6263,N_6284);
nand U6476 (N_6476,N_6210,N_6366);
or U6477 (N_6477,N_6309,N_6283);
xnor U6478 (N_6478,N_6282,N_6330);
or U6479 (N_6479,N_6333,N_6374);
or U6480 (N_6480,N_6229,N_6225);
nand U6481 (N_6481,N_6266,N_6369);
and U6482 (N_6482,N_6289,N_6379);
xor U6483 (N_6483,N_6296,N_6212);
nand U6484 (N_6484,N_6200,N_6337);
and U6485 (N_6485,N_6230,N_6297);
xnor U6486 (N_6486,N_6389,N_6393);
or U6487 (N_6487,N_6214,N_6278);
or U6488 (N_6488,N_6316,N_6234);
or U6489 (N_6489,N_6364,N_6222);
xor U6490 (N_6490,N_6295,N_6367);
nand U6491 (N_6491,N_6260,N_6391);
nand U6492 (N_6492,N_6359,N_6394);
or U6493 (N_6493,N_6361,N_6319);
nor U6494 (N_6494,N_6328,N_6261);
or U6495 (N_6495,N_6344,N_6383);
xnor U6496 (N_6496,N_6233,N_6390);
nor U6497 (N_6497,N_6294,N_6206);
or U6498 (N_6498,N_6299,N_6298);
xnor U6499 (N_6499,N_6287,N_6375);
xor U6500 (N_6500,N_6265,N_6275);
or U6501 (N_6501,N_6388,N_6320);
and U6502 (N_6502,N_6327,N_6346);
xnor U6503 (N_6503,N_6279,N_6254);
xor U6504 (N_6504,N_6327,N_6260);
nand U6505 (N_6505,N_6293,N_6268);
nor U6506 (N_6506,N_6379,N_6354);
or U6507 (N_6507,N_6334,N_6235);
nor U6508 (N_6508,N_6212,N_6215);
and U6509 (N_6509,N_6309,N_6364);
xnor U6510 (N_6510,N_6343,N_6288);
xor U6511 (N_6511,N_6272,N_6261);
xor U6512 (N_6512,N_6244,N_6230);
nor U6513 (N_6513,N_6398,N_6294);
and U6514 (N_6514,N_6356,N_6206);
and U6515 (N_6515,N_6374,N_6245);
xnor U6516 (N_6516,N_6398,N_6235);
or U6517 (N_6517,N_6231,N_6247);
and U6518 (N_6518,N_6287,N_6257);
nor U6519 (N_6519,N_6329,N_6338);
nand U6520 (N_6520,N_6207,N_6205);
or U6521 (N_6521,N_6216,N_6295);
xor U6522 (N_6522,N_6298,N_6318);
or U6523 (N_6523,N_6214,N_6304);
or U6524 (N_6524,N_6294,N_6227);
or U6525 (N_6525,N_6320,N_6211);
xnor U6526 (N_6526,N_6325,N_6337);
nand U6527 (N_6527,N_6313,N_6227);
xor U6528 (N_6528,N_6373,N_6249);
nor U6529 (N_6529,N_6306,N_6278);
or U6530 (N_6530,N_6201,N_6207);
nand U6531 (N_6531,N_6378,N_6205);
xnor U6532 (N_6532,N_6374,N_6218);
and U6533 (N_6533,N_6356,N_6359);
nand U6534 (N_6534,N_6228,N_6329);
xnor U6535 (N_6535,N_6248,N_6244);
and U6536 (N_6536,N_6288,N_6242);
nor U6537 (N_6537,N_6305,N_6351);
nor U6538 (N_6538,N_6292,N_6291);
nor U6539 (N_6539,N_6223,N_6381);
nor U6540 (N_6540,N_6294,N_6314);
or U6541 (N_6541,N_6397,N_6249);
nand U6542 (N_6542,N_6292,N_6248);
nand U6543 (N_6543,N_6223,N_6279);
nand U6544 (N_6544,N_6222,N_6235);
and U6545 (N_6545,N_6253,N_6285);
or U6546 (N_6546,N_6303,N_6353);
nand U6547 (N_6547,N_6278,N_6274);
xor U6548 (N_6548,N_6205,N_6297);
and U6549 (N_6549,N_6399,N_6224);
nor U6550 (N_6550,N_6256,N_6204);
or U6551 (N_6551,N_6293,N_6201);
and U6552 (N_6552,N_6260,N_6230);
or U6553 (N_6553,N_6386,N_6253);
nor U6554 (N_6554,N_6202,N_6304);
nor U6555 (N_6555,N_6303,N_6358);
nor U6556 (N_6556,N_6253,N_6340);
xnor U6557 (N_6557,N_6216,N_6359);
nor U6558 (N_6558,N_6271,N_6251);
xnor U6559 (N_6559,N_6290,N_6323);
and U6560 (N_6560,N_6207,N_6329);
nor U6561 (N_6561,N_6268,N_6385);
xor U6562 (N_6562,N_6305,N_6274);
nand U6563 (N_6563,N_6339,N_6295);
and U6564 (N_6564,N_6303,N_6333);
and U6565 (N_6565,N_6300,N_6270);
nand U6566 (N_6566,N_6265,N_6377);
and U6567 (N_6567,N_6281,N_6371);
or U6568 (N_6568,N_6331,N_6350);
xnor U6569 (N_6569,N_6205,N_6287);
xor U6570 (N_6570,N_6364,N_6297);
or U6571 (N_6571,N_6327,N_6323);
and U6572 (N_6572,N_6249,N_6318);
xnor U6573 (N_6573,N_6255,N_6294);
or U6574 (N_6574,N_6235,N_6230);
and U6575 (N_6575,N_6395,N_6232);
nand U6576 (N_6576,N_6279,N_6241);
nand U6577 (N_6577,N_6233,N_6308);
and U6578 (N_6578,N_6374,N_6352);
or U6579 (N_6579,N_6209,N_6206);
nor U6580 (N_6580,N_6384,N_6226);
nor U6581 (N_6581,N_6253,N_6249);
and U6582 (N_6582,N_6370,N_6382);
xor U6583 (N_6583,N_6313,N_6345);
nand U6584 (N_6584,N_6306,N_6217);
or U6585 (N_6585,N_6388,N_6333);
nand U6586 (N_6586,N_6371,N_6339);
and U6587 (N_6587,N_6276,N_6393);
and U6588 (N_6588,N_6378,N_6329);
nand U6589 (N_6589,N_6206,N_6381);
xor U6590 (N_6590,N_6328,N_6395);
nor U6591 (N_6591,N_6270,N_6391);
or U6592 (N_6592,N_6239,N_6327);
and U6593 (N_6593,N_6209,N_6291);
xor U6594 (N_6594,N_6218,N_6231);
nand U6595 (N_6595,N_6376,N_6316);
and U6596 (N_6596,N_6247,N_6238);
and U6597 (N_6597,N_6245,N_6212);
nor U6598 (N_6598,N_6225,N_6264);
or U6599 (N_6599,N_6280,N_6284);
and U6600 (N_6600,N_6419,N_6469);
and U6601 (N_6601,N_6545,N_6479);
and U6602 (N_6602,N_6564,N_6482);
or U6603 (N_6603,N_6474,N_6503);
or U6604 (N_6604,N_6560,N_6446);
or U6605 (N_6605,N_6417,N_6444);
nor U6606 (N_6606,N_6527,N_6486);
nor U6607 (N_6607,N_6595,N_6478);
or U6608 (N_6608,N_6483,N_6459);
nand U6609 (N_6609,N_6568,N_6462);
or U6610 (N_6610,N_6430,N_6575);
nor U6611 (N_6611,N_6422,N_6463);
and U6612 (N_6612,N_6596,N_6535);
and U6613 (N_6613,N_6520,N_6497);
nand U6614 (N_6614,N_6490,N_6500);
nor U6615 (N_6615,N_6401,N_6461);
nor U6616 (N_6616,N_6528,N_6404);
xor U6617 (N_6617,N_6484,N_6412);
xnor U6618 (N_6618,N_6519,N_6517);
and U6619 (N_6619,N_6439,N_6584);
xor U6620 (N_6620,N_6526,N_6505);
and U6621 (N_6621,N_6578,N_6453);
nor U6622 (N_6622,N_6570,N_6576);
nand U6623 (N_6623,N_6567,N_6443);
or U6624 (N_6624,N_6590,N_6423);
and U6625 (N_6625,N_6433,N_6544);
or U6626 (N_6626,N_6425,N_6427);
nand U6627 (N_6627,N_6554,N_6559);
nor U6628 (N_6628,N_6466,N_6518);
and U6629 (N_6629,N_6496,N_6543);
nand U6630 (N_6630,N_6408,N_6438);
nor U6631 (N_6631,N_6541,N_6524);
xor U6632 (N_6632,N_6485,N_6562);
or U6633 (N_6633,N_6566,N_6441);
nand U6634 (N_6634,N_6548,N_6592);
and U6635 (N_6635,N_6514,N_6416);
and U6636 (N_6636,N_6458,N_6599);
nor U6637 (N_6637,N_6569,N_6550);
xnor U6638 (N_6638,N_6581,N_6471);
nand U6639 (N_6639,N_6480,N_6525);
or U6640 (N_6640,N_6556,N_6579);
xor U6641 (N_6641,N_6561,N_6472);
nand U6642 (N_6642,N_6494,N_6598);
nand U6643 (N_6643,N_6491,N_6418);
or U6644 (N_6644,N_6531,N_6421);
nand U6645 (N_6645,N_6555,N_6492);
and U6646 (N_6646,N_6530,N_6467);
xnor U6647 (N_6647,N_6452,N_6504);
nor U6648 (N_6648,N_6552,N_6539);
xnor U6649 (N_6649,N_6434,N_6426);
and U6650 (N_6650,N_6481,N_6523);
or U6651 (N_6651,N_6499,N_6410);
nand U6652 (N_6652,N_6583,N_6487);
xnor U6653 (N_6653,N_6411,N_6587);
and U6654 (N_6654,N_6400,N_6515);
or U6655 (N_6655,N_6432,N_6589);
nand U6656 (N_6656,N_6551,N_6502);
nor U6657 (N_6657,N_6546,N_6455);
xnor U6658 (N_6658,N_6457,N_6488);
nor U6659 (N_6659,N_6473,N_6431);
xnor U6660 (N_6660,N_6477,N_6521);
and U6661 (N_6661,N_6495,N_6597);
xnor U6662 (N_6662,N_6435,N_6538);
and U6663 (N_6663,N_6407,N_6454);
nand U6664 (N_6664,N_6507,N_6413);
nand U6665 (N_6665,N_6537,N_6445);
and U6666 (N_6666,N_6571,N_6456);
or U6667 (N_6667,N_6415,N_6588);
xor U6668 (N_6668,N_6428,N_6509);
and U6669 (N_6669,N_6489,N_6448);
and U6670 (N_6670,N_6573,N_6508);
nor U6671 (N_6671,N_6549,N_6510);
nand U6672 (N_6672,N_6437,N_6475);
nand U6673 (N_6673,N_6464,N_6512);
nor U6674 (N_6674,N_6536,N_6501);
or U6675 (N_6675,N_6436,N_6513);
xnor U6676 (N_6676,N_6440,N_6547);
or U6677 (N_6677,N_6470,N_6468);
nand U6678 (N_6678,N_6558,N_6593);
and U6679 (N_6679,N_6580,N_6534);
or U6680 (N_6680,N_6451,N_6409);
xnor U6681 (N_6681,N_6406,N_6585);
xnor U6682 (N_6682,N_6540,N_6405);
xnor U6683 (N_6683,N_6506,N_6572);
nor U6684 (N_6684,N_6529,N_6460);
nand U6685 (N_6685,N_6429,N_6577);
and U6686 (N_6686,N_6557,N_6522);
or U6687 (N_6687,N_6402,N_6449);
nor U6688 (N_6688,N_6424,N_6465);
or U6689 (N_6689,N_6594,N_6420);
or U6690 (N_6690,N_6565,N_6586);
or U6691 (N_6691,N_6533,N_6574);
xnor U6692 (N_6692,N_6450,N_6542);
xor U6693 (N_6693,N_6591,N_6403);
nand U6694 (N_6694,N_6553,N_6563);
xor U6695 (N_6695,N_6532,N_6493);
and U6696 (N_6696,N_6476,N_6442);
nor U6697 (N_6697,N_6498,N_6582);
and U6698 (N_6698,N_6511,N_6414);
and U6699 (N_6699,N_6447,N_6516);
or U6700 (N_6700,N_6482,N_6468);
nor U6701 (N_6701,N_6479,N_6547);
nand U6702 (N_6702,N_6518,N_6505);
nor U6703 (N_6703,N_6548,N_6414);
nand U6704 (N_6704,N_6478,N_6561);
or U6705 (N_6705,N_6452,N_6598);
xor U6706 (N_6706,N_6531,N_6469);
and U6707 (N_6707,N_6591,N_6554);
nor U6708 (N_6708,N_6530,N_6546);
xnor U6709 (N_6709,N_6470,N_6485);
xor U6710 (N_6710,N_6469,N_6564);
xnor U6711 (N_6711,N_6581,N_6483);
xnor U6712 (N_6712,N_6400,N_6506);
nor U6713 (N_6713,N_6544,N_6508);
nor U6714 (N_6714,N_6579,N_6559);
and U6715 (N_6715,N_6586,N_6476);
xor U6716 (N_6716,N_6535,N_6494);
or U6717 (N_6717,N_6519,N_6587);
or U6718 (N_6718,N_6545,N_6451);
nand U6719 (N_6719,N_6445,N_6402);
nand U6720 (N_6720,N_6502,N_6576);
and U6721 (N_6721,N_6462,N_6496);
and U6722 (N_6722,N_6549,N_6423);
nand U6723 (N_6723,N_6566,N_6459);
or U6724 (N_6724,N_6436,N_6549);
nand U6725 (N_6725,N_6544,N_6566);
nand U6726 (N_6726,N_6422,N_6527);
nand U6727 (N_6727,N_6502,N_6577);
and U6728 (N_6728,N_6560,N_6585);
or U6729 (N_6729,N_6556,N_6441);
or U6730 (N_6730,N_6589,N_6422);
or U6731 (N_6731,N_6459,N_6402);
nor U6732 (N_6732,N_6556,N_6580);
and U6733 (N_6733,N_6457,N_6563);
or U6734 (N_6734,N_6563,N_6424);
or U6735 (N_6735,N_6538,N_6492);
nand U6736 (N_6736,N_6429,N_6580);
nand U6737 (N_6737,N_6408,N_6495);
xor U6738 (N_6738,N_6578,N_6509);
or U6739 (N_6739,N_6530,N_6452);
nor U6740 (N_6740,N_6401,N_6536);
nand U6741 (N_6741,N_6538,N_6599);
xnor U6742 (N_6742,N_6496,N_6571);
nand U6743 (N_6743,N_6509,N_6528);
xnor U6744 (N_6744,N_6418,N_6558);
xor U6745 (N_6745,N_6405,N_6518);
and U6746 (N_6746,N_6411,N_6530);
and U6747 (N_6747,N_6528,N_6582);
nor U6748 (N_6748,N_6554,N_6431);
nor U6749 (N_6749,N_6567,N_6414);
xnor U6750 (N_6750,N_6578,N_6499);
and U6751 (N_6751,N_6570,N_6475);
nand U6752 (N_6752,N_6403,N_6546);
xor U6753 (N_6753,N_6472,N_6519);
or U6754 (N_6754,N_6534,N_6508);
xor U6755 (N_6755,N_6560,N_6575);
nor U6756 (N_6756,N_6532,N_6514);
or U6757 (N_6757,N_6479,N_6548);
xor U6758 (N_6758,N_6576,N_6532);
and U6759 (N_6759,N_6445,N_6508);
nor U6760 (N_6760,N_6407,N_6420);
nor U6761 (N_6761,N_6481,N_6559);
and U6762 (N_6762,N_6544,N_6502);
nand U6763 (N_6763,N_6587,N_6569);
and U6764 (N_6764,N_6571,N_6547);
and U6765 (N_6765,N_6460,N_6532);
and U6766 (N_6766,N_6451,N_6415);
and U6767 (N_6767,N_6477,N_6401);
or U6768 (N_6768,N_6579,N_6401);
nor U6769 (N_6769,N_6430,N_6422);
and U6770 (N_6770,N_6542,N_6595);
and U6771 (N_6771,N_6439,N_6410);
nand U6772 (N_6772,N_6519,N_6442);
nor U6773 (N_6773,N_6467,N_6512);
xnor U6774 (N_6774,N_6417,N_6528);
nand U6775 (N_6775,N_6488,N_6400);
and U6776 (N_6776,N_6455,N_6483);
nor U6777 (N_6777,N_6567,N_6465);
nand U6778 (N_6778,N_6428,N_6577);
nor U6779 (N_6779,N_6508,N_6564);
xnor U6780 (N_6780,N_6543,N_6508);
xnor U6781 (N_6781,N_6587,N_6486);
nor U6782 (N_6782,N_6429,N_6442);
nand U6783 (N_6783,N_6477,N_6454);
and U6784 (N_6784,N_6454,N_6473);
xor U6785 (N_6785,N_6511,N_6496);
or U6786 (N_6786,N_6476,N_6592);
or U6787 (N_6787,N_6412,N_6560);
nor U6788 (N_6788,N_6505,N_6448);
nand U6789 (N_6789,N_6409,N_6594);
and U6790 (N_6790,N_6532,N_6547);
nor U6791 (N_6791,N_6495,N_6544);
nand U6792 (N_6792,N_6426,N_6406);
nand U6793 (N_6793,N_6590,N_6503);
and U6794 (N_6794,N_6498,N_6499);
and U6795 (N_6795,N_6491,N_6557);
xnor U6796 (N_6796,N_6527,N_6469);
nor U6797 (N_6797,N_6413,N_6449);
and U6798 (N_6798,N_6452,N_6589);
or U6799 (N_6799,N_6565,N_6437);
or U6800 (N_6800,N_6682,N_6685);
and U6801 (N_6801,N_6790,N_6651);
and U6802 (N_6802,N_6735,N_6636);
or U6803 (N_6803,N_6742,N_6763);
and U6804 (N_6804,N_6678,N_6628);
and U6805 (N_6805,N_6662,N_6773);
nand U6806 (N_6806,N_6644,N_6686);
nor U6807 (N_6807,N_6648,N_6778);
and U6808 (N_6808,N_6769,N_6788);
and U6809 (N_6809,N_6745,N_6676);
or U6810 (N_6810,N_6620,N_6670);
xor U6811 (N_6811,N_6689,N_6796);
or U6812 (N_6812,N_6654,N_6627);
xnor U6813 (N_6813,N_6797,N_6663);
and U6814 (N_6814,N_6657,N_6690);
nand U6815 (N_6815,N_6658,N_6641);
or U6816 (N_6816,N_6780,N_6711);
and U6817 (N_6817,N_6738,N_6737);
xor U6818 (N_6818,N_6691,N_6710);
nand U6819 (N_6819,N_6615,N_6709);
and U6820 (N_6820,N_6656,N_6762);
nor U6821 (N_6821,N_6713,N_6772);
or U6822 (N_6822,N_6633,N_6617);
or U6823 (N_6823,N_6770,N_6698);
nor U6824 (N_6824,N_6688,N_6647);
or U6825 (N_6825,N_6766,N_6792);
and U6826 (N_6826,N_6704,N_6640);
nor U6827 (N_6827,N_6666,N_6629);
nor U6828 (N_6828,N_6734,N_6605);
nand U6829 (N_6829,N_6652,N_6746);
xor U6830 (N_6830,N_6736,N_6750);
or U6831 (N_6831,N_6779,N_6692);
nor U6832 (N_6832,N_6785,N_6791);
or U6833 (N_6833,N_6731,N_6621);
and U6834 (N_6834,N_6696,N_6661);
and U6835 (N_6835,N_6799,N_6673);
and U6836 (N_6836,N_6700,N_6624);
xor U6837 (N_6837,N_6757,N_6755);
nor U6838 (N_6838,N_6600,N_6608);
xnor U6839 (N_6839,N_6715,N_6753);
and U6840 (N_6840,N_6758,N_6752);
xor U6841 (N_6841,N_6606,N_6639);
nor U6842 (N_6842,N_6725,N_6722);
xnor U6843 (N_6843,N_6703,N_6717);
xnor U6844 (N_6844,N_6756,N_6759);
xor U6845 (N_6845,N_6705,N_6635);
and U6846 (N_6846,N_6783,N_6614);
and U6847 (N_6847,N_6706,N_6789);
nor U6848 (N_6848,N_6681,N_6687);
nand U6849 (N_6849,N_6665,N_6623);
or U6850 (N_6850,N_6795,N_6695);
and U6851 (N_6851,N_6760,N_6694);
or U6852 (N_6852,N_6649,N_6754);
nor U6853 (N_6853,N_6630,N_6727);
and U6854 (N_6854,N_6743,N_6776);
or U6855 (N_6855,N_6612,N_6764);
and U6856 (N_6856,N_6642,N_6765);
or U6857 (N_6857,N_6718,N_6677);
xor U6858 (N_6858,N_6619,N_6626);
xnor U6859 (N_6859,N_6781,N_6748);
nand U6860 (N_6860,N_6723,N_6714);
xnor U6861 (N_6861,N_6740,N_6786);
or U6862 (N_6862,N_6611,N_6732);
nor U6863 (N_6863,N_6645,N_6733);
and U6864 (N_6864,N_6664,N_6684);
and U6865 (N_6865,N_6650,N_6716);
nor U6866 (N_6866,N_6749,N_6609);
nor U6867 (N_6867,N_6712,N_6613);
or U6868 (N_6868,N_6634,N_6798);
and U6869 (N_6869,N_6697,N_6653);
or U6870 (N_6870,N_6669,N_6768);
and U6871 (N_6871,N_6637,N_6702);
or U6872 (N_6872,N_6674,N_6777);
xor U6873 (N_6873,N_6782,N_6784);
nand U6874 (N_6874,N_6604,N_6679);
xor U6875 (N_6875,N_6631,N_6659);
nand U6876 (N_6876,N_6701,N_6601);
nor U6877 (N_6877,N_6618,N_6767);
and U6878 (N_6878,N_6729,N_6668);
nor U6879 (N_6879,N_6708,N_6720);
nor U6880 (N_6880,N_6793,N_6646);
or U6881 (N_6881,N_6775,N_6787);
xnor U6882 (N_6882,N_6707,N_6622);
xor U6883 (N_6883,N_6728,N_6751);
and U6884 (N_6884,N_6616,N_6602);
xnor U6885 (N_6885,N_6747,N_6726);
xor U6886 (N_6886,N_6680,N_6660);
nor U6887 (N_6887,N_6603,N_6724);
nand U6888 (N_6888,N_6632,N_6643);
and U6889 (N_6889,N_6761,N_6774);
nand U6890 (N_6890,N_6655,N_6744);
xnor U6891 (N_6891,N_6699,N_6719);
nand U6892 (N_6892,N_6607,N_6683);
or U6893 (N_6893,N_6625,N_6730);
xor U6894 (N_6894,N_6794,N_6693);
xnor U6895 (N_6895,N_6741,N_6675);
nand U6896 (N_6896,N_6610,N_6721);
xor U6897 (N_6897,N_6671,N_6667);
nor U6898 (N_6898,N_6638,N_6672);
xor U6899 (N_6899,N_6739,N_6771);
or U6900 (N_6900,N_6654,N_6768);
or U6901 (N_6901,N_6672,N_6795);
xor U6902 (N_6902,N_6624,N_6780);
nand U6903 (N_6903,N_6799,N_6761);
nand U6904 (N_6904,N_6743,N_6734);
and U6905 (N_6905,N_6688,N_6783);
xor U6906 (N_6906,N_6764,N_6713);
nand U6907 (N_6907,N_6708,N_6665);
nand U6908 (N_6908,N_6756,N_6797);
nand U6909 (N_6909,N_6765,N_6648);
xnor U6910 (N_6910,N_6608,N_6756);
nand U6911 (N_6911,N_6698,N_6697);
and U6912 (N_6912,N_6757,N_6662);
nor U6913 (N_6913,N_6712,N_6698);
xnor U6914 (N_6914,N_6664,N_6631);
or U6915 (N_6915,N_6747,N_6746);
or U6916 (N_6916,N_6698,N_6686);
and U6917 (N_6917,N_6763,N_6792);
nand U6918 (N_6918,N_6706,N_6602);
nand U6919 (N_6919,N_6772,N_6793);
and U6920 (N_6920,N_6740,N_6727);
xor U6921 (N_6921,N_6640,N_6786);
xnor U6922 (N_6922,N_6786,N_6779);
or U6923 (N_6923,N_6770,N_6645);
nor U6924 (N_6924,N_6787,N_6780);
xnor U6925 (N_6925,N_6625,N_6742);
nor U6926 (N_6926,N_6776,N_6768);
nand U6927 (N_6927,N_6724,N_6742);
xor U6928 (N_6928,N_6621,N_6730);
and U6929 (N_6929,N_6741,N_6637);
nor U6930 (N_6930,N_6717,N_6770);
and U6931 (N_6931,N_6635,N_6774);
or U6932 (N_6932,N_6601,N_6732);
xor U6933 (N_6933,N_6681,N_6691);
or U6934 (N_6934,N_6701,N_6740);
xor U6935 (N_6935,N_6766,N_6711);
and U6936 (N_6936,N_6740,N_6764);
or U6937 (N_6937,N_6735,N_6610);
xnor U6938 (N_6938,N_6778,N_6754);
and U6939 (N_6939,N_6711,N_6637);
nand U6940 (N_6940,N_6791,N_6780);
or U6941 (N_6941,N_6638,N_6739);
nand U6942 (N_6942,N_6669,N_6729);
nor U6943 (N_6943,N_6752,N_6777);
or U6944 (N_6944,N_6720,N_6662);
nand U6945 (N_6945,N_6780,N_6726);
and U6946 (N_6946,N_6783,N_6765);
and U6947 (N_6947,N_6654,N_6699);
nand U6948 (N_6948,N_6651,N_6770);
or U6949 (N_6949,N_6630,N_6711);
xnor U6950 (N_6950,N_6752,N_6697);
nor U6951 (N_6951,N_6759,N_6785);
nor U6952 (N_6952,N_6666,N_6797);
nand U6953 (N_6953,N_6713,N_6747);
and U6954 (N_6954,N_6744,N_6792);
xnor U6955 (N_6955,N_6627,N_6643);
nand U6956 (N_6956,N_6752,N_6696);
and U6957 (N_6957,N_6687,N_6787);
xnor U6958 (N_6958,N_6707,N_6682);
or U6959 (N_6959,N_6698,N_6606);
nor U6960 (N_6960,N_6708,N_6600);
xnor U6961 (N_6961,N_6600,N_6747);
nand U6962 (N_6962,N_6763,N_6774);
xnor U6963 (N_6963,N_6727,N_6658);
or U6964 (N_6964,N_6750,N_6674);
xor U6965 (N_6965,N_6621,N_6619);
xnor U6966 (N_6966,N_6785,N_6795);
nand U6967 (N_6967,N_6718,N_6692);
and U6968 (N_6968,N_6784,N_6620);
nand U6969 (N_6969,N_6626,N_6603);
nor U6970 (N_6970,N_6709,N_6676);
and U6971 (N_6971,N_6738,N_6679);
nor U6972 (N_6972,N_6620,N_6741);
nand U6973 (N_6973,N_6671,N_6680);
nand U6974 (N_6974,N_6666,N_6746);
xnor U6975 (N_6975,N_6784,N_6755);
nor U6976 (N_6976,N_6695,N_6685);
nand U6977 (N_6977,N_6791,N_6712);
nand U6978 (N_6978,N_6761,N_6760);
and U6979 (N_6979,N_6793,N_6602);
xor U6980 (N_6980,N_6628,N_6641);
nor U6981 (N_6981,N_6784,N_6739);
nand U6982 (N_6982,N_6703,N_6755);
nand U6983 (N_6983,N_6695,N_6760);
nand U6984 (N_6984,N_6609,N_6719);
or U6985 (N_6985,N_6690,N_6601);
xor U6986 (N_6986,N_6791,N_6639);
or U6987 (N_6987,N_6632,N_6723);
or U6988 (N_6988,N_6753,N_6713);
xor U6989 (N_6989,N_6731,N_6716);
nand U6990 (N_6990,N_6786,N_6790);
and U6991 (N_6991,N_6708,N_6690);
nor U6992 (N_6992,N_6671,N_6787);
nor U6993 (N_6993,N_6618,N_6768);
nor U6994 (N_6994,N_6629,N_6704);
nand U6995 (N_6995,N_6664,N_6648);
nand U6996 (N_6996,N_6695,N_6636);
nand U6997 (N_6997,N_6621,N_6661);
nor U6998 (N_6998,N_6754,N_6715);
nor U6999 (N_6999,N_6661,N_6625);
or U7000 (N_7000,N_6810,N_6952);
xor U7001 (N_7001,N_6857,N_6907);
xor U7002 (N_7002,N_6839,N_6830);
nor U7003 (N_7003,N_6884,N_6987);
nor U7004 (N_7004,N_6920,N_6828);
or U7005 (N_7005,N_6937,N_6893);
xor U7006 (N_7006,N_6914,N_6980);
or U7007 (N_7007,N_6860,N_6995);
and U7008 (N_7008,N_6803,N_6879);
and U7009 (N_7009,N_6872,N_6912);
nand U7010 (N_7010,N_6918,N_6926);
nand U7011 (N_7011,N_6925,N_6855);
nor U7012 (N_7012,N_6984,N_6886);
and U7013 (N_7013,N_6852,N_6845);
or U7014 (N_7014,N_6835,N_6801);
nor U7015 (N_7015,N_6858,N_6955);
nor U7016 (N_7016,N_6924,N_6969);
or U7017 (N_7017,N_6878,N_6881);
and U7018 (N_7018,N_6967,N_6862);
and U7019 (N_7019,N_6934,N_6947);
xor U7020 (N_7020,N_6919,N_6948);
nor U7021 (N_7021,N_6829,N_6856);
or U7022 (N_7022,N_6994,N_6951);
nor U7023 (N_7023,N_6929,N_6885);
nor U7024 (N_7024,N_6811,N_6807);
nor U7025 (N_7025,N_6815,N_6910);
and U7026 (N_7026,N_6968,N_6804);
nand U7027 (N_7027,N_6996,N_6961);
xnor U7028 (N_7028,N_6818,N_6978);
xnor U7029 (N_7029,N_6981,N_6876);
nor U7030 (N_7030,N_6888,N_6826);
nand U7031 (N_7031,N_6932,N_6941);
nand U7032 (N_7032,N_6846,N_6911);
xor U7033 (N_7033,N_6843,N_6887);
or U7034 (N_7034,N_6960,N_6901);
or U7035 (N_7035,N_6859,N_6966);
xor U7036 (N_7036,N_6809,N_6800);
or U7037 (N_7037,N_6896,N_6870);
and U7038 (N_7038,N_6903,N_6900);
nand U7039 (N_7039,N_6850,N_6827);
or U7040 (N_7040,N_6864,N_6849);
or U7041 (N_7041,N_6805,N_6820);
or U7042 (N_7042,N_6953,N_6848);
nand U7043 (N_7043,N_6923,N_6821);
xor U7044 (N_7044,N_6871,N_6808);
nor U7045 (N_7045,N_6959,N_6970);
and U7046 (N_7046,N_6935,N_6931);
xnor U7047 (N_7047,N_6847,N_6812);
or U7048 (N_7048,N_6939,N_6913);
or U7049 (N_7049,N_6868,N_6892);
xor U7050 (N_7050,N_6963,N_6989);
xnor U7051 (N_7051,N_6999,N_6840);
nor U7052 (N_7052,N_6854,N_6942);
nor U7053 (N_7053,N_6957,N_6950);
and U7054 (N_7054,N_6956,N_6902);
nor U7055 (N_7055,N_6825,N_6930);
or U7056 (N_7056,N_6917,N_6979);
or U7057 (N_7057,N_6928,N_6927);
nor U7058 (N_7058,N_6844,N_6891);
or U7059 (N_7059,N_6832,N_6822);
nand U7060 (N_7060,N_6975,N_6972);
and U7061 (N_7061,N_6904,N_6816);
xnor U7062 (N_7062,N_6863,N_6874);
nor U7063 (N_7063,N_6938,N_6806);
nor U7064 (N_7064,N_6992,N_6986);
or U7065 (N_7065,N_6853,N_6958);
nand U7066 (N_7066,N_6976,N_6851);
and U7067 (N_7067,N_6819,N_6915);
and U7068 (N_7068,N_6817,N_6833);
and U7069 (N_7069,N_6869,N_6988);
or U7070 (N_7070,N_6883,N_6895);
nor U7071 (N_7071,N_6965,N_6875);
nand U7072 (N_7072,N_6991,N_6880);
nor U7073 (N_7073,N_6873,N_6823);
nand U7074 (N_7074,N_6985,N_6824);
and U7075 (N_7075,N_6894,N_6866);
nor U7076 (N_7076,N_6921,N_6905);
nor U7077 (N_7077,N_6922,N_6946);
xor U7078 (N_7078,N_6813,N_6841);
or U7079 (N_7079,N_6971,N_6802);
and U7080 (N_7080,N_6834,N_6974);
nand U7081 (N_7081,N_6936,N_6977);
nor U7082 (N_7082,N_6916,N_6889);
xnor U7083 (N_7083,N_6964,N_6983);
or U7084 (N_7084,N_6982,N_6890);
nand U7085 (N_7085,N_6877,N_6962);
and U7086 (N_7086,N_6973,N_6997);
xor U7087 (N_7087,N_6831,N_6906);
or U7088 (N_7088,N_6998,N_6908);
xnor U7089 (N_7089,N_6909,N_6949);
or U7090 (N_7090,N_6940,N_6943);
nor U7091 (N_7091,N_6944,N_6945);
nor U7092 (N_7092,N_6842,N_6993);
and U7093 (N_7093,N_6838,N_6867);
xor U7094 (N_7094,N_6882,N_6990);
xor U7095 (N_7095,N_6898,N_6899);
xor U7096 (N_7096,N_6837,N_6897);
nor U7097 (N_7097,N_6861,N_6836);
and U7098 (N_7098,N_6933,N_6954);
and U7099 (N_7099,N_6865,N_6814);
nor U7100 (N_7100,N_6918,N_6903);
and U7101 (N_7101,N_6809,N_6904);
nor U7102 (N_7102,N_6962,N_6925);
nand U7103 (N_7103,N_6827,N_6831);
xor U7104 (N_7104,N_6940,N_6945);
nand U7105 (N_7105,N_6847,N_6895);
nor U7106 (N_7106,N_6817,N_6897);
and U7107 (N_7107,N_6944,N_6826);
xnor U7108 (N_7108,N_6977,N_6953);
nand U7109 (N_7109,N_6939,N_6847);
nand U7110 (N_7110,N_6915,N_6904);
or U7111 (N_7111,N_6802,N_6929);
nand U7112 (N_7112,N_6820,N_6929);
nor U7113 (N_7113,N_6899,N_6833);
nor U7114 (N_7114,N_6904,N_6801);
or U7115 (N_7115,N_6857,N_6896);
xnor U7116 (N_7116,N_6880,N_6833);
or U7117 (N_7117,N_6953,N_6956);
and U7118 (N_7118,N_6910,N_6955);
xnor U7119 (N_7119,N_6902,N_6995);
nand U7120 (N_7120,N_6822,N_6868);
xor U7121 (N_7121,N_6822,N_6846);
or U7122 (N_7122,N_6886,N_6942);
xor U7123 (N_7123,N_6825,N_6879);
nand U7124 (N_7124,N_6999,N_6828);
nor U7125 (N_7125,N_6958,N_6991);
and U7126 (N_7126,N_6932,N_6804);
nor U7127 (N_7127,N_6928,N_6972);
nor U7128 (N_7128,N_6984,N_6982);
or U7129 (N_7129,N_6888,N_6874);
nand U7130 (N_7130,N_6945,N_6949);
or U7131 (N_7131,N_6988,N_6893);
or U7132 (N_7132,N_6955,N_6871);
nand U7133 (N_7133,N_6965,N_6979);
xnor U7134 (N_7134,N_6846,N_6805);
xor U7135 (N_7135,N_6943,N_6838);
xor U7136 (N_7136,N_6866,N_6833);
or U7137 (N_7137,N_6808,N_6885);
xnor U7138 (N_7138,N_6942,N_6882);
and U7139 (N_7139,N_6928,N_6975);
nand U7140 (N_7140,N_6929,N_6873);
or U7141 (N_7141,N_6951,N_6946);
nor U7142 (N_7142,N_6838,N_6825);
or U7143 (N_7143,N_6819,N_6958);
and U7144 (N_7144,N_6864,N_6826);
or U7145 (N_7145,N_6907,N_6855);
nand U7146 (N_7146,N_6935,N_6970);
or U7147 (N_7147,N_6803,N_6998);
xor U7148 (N_7148,N_6904,N_6832);
nor U7149 (N_7149,N_6858,N_6864);
nand U7150 (N_7150,N_6967,N_6935);
and U7151 (N_7151,N_6967,N_6835);
or U7152 (N_7152,N_6975,N_6935);
and U7153 (N_7153,N_6999,N_6849);
nand U7154 (N_7154,N_6901,N_6986);
or U7155 (N_7155,N_6949,N_6996);
and U7156 (N_7156,N_6860,N_6922);
nor U7157 (N_7157,N_6984,N_6989);
and U7158 (N_7158,N_6823,N_6966);
or U7159 (N_7159,N_6956,N_6938);
nand U7160 (N_7160,N_6907,N_6843);
or U7161 (N_7161,N_6993,N_6853);
and U7162 (N_7162,N_6947,N_6951);
and U7163 (N_7163,N_6831,N_6869);
nand U7164 (N_7164,N_6889,N_6884);
nor U7165 (N_7165,N_6967,N_6879);
nor U7166 (N_7166,N_6865,N_6910);
xnor U7167 (N_7167,N_6804,N_6930);
and U7168 (N_7168,N_6862,N_6868);
nand U7169 (N_7169,N_6980,N_6900);
xor U7170 (N_7170,N_6889,N_6836);
or U7171 (N_7171,N_6904,N_6858);
xor U7172 (N_7172,N_6837,N_6836);
or U7173 (N_7173,N_6805,N_6891);
or U7174 (N_7174,N_6818,N_6981);
and U7175 (N_7175,N_6807,N_6871);
xnor U7176 (N_7176,N_6816,N_6886);
xor U7177 (N_7177,N_6870,N_6998);
or U7178 (N_7178,N_6980,N_6898);
xnor U7179 (N_7179,N_6970,N_6898);
nand U7180 (N_7180,N_6805,N_6849);
or U7181 (N_7181,N_6831,N_6962);
or U7182 (N_7182,N_6836,N_6873);
xor U7183 (N_7183,N_6819,N_6969);
nor U7184 (N_7184,N_6875,N_6917);
nor U7185 (N_7185,N_6865,N_6984);
nor U7186 (N_7186,N_6916,N_6876);
and U7187 (N_7187,N_6858,N_6820);
and U7188 (N_7188,N_6923,N_6808);
and U7189 (N_7189,N_6955,N_6815);
nor U7190 (N_7190,N_6935,N_6854);
nand U7191 (N_7191,N_6945,N_6818);
xor U7192 (N_7192,N_6869,N_6911);
or U7193 (N_7193,N_6949,N_6811);
nand U7194 (N_7194,N_6862,N_6993);
nand U7195 (N_7195,N_6873,N_6944);
xor U7196 (N_7196,N_6951,N_6932);
or U7197 (N_7197,N_6957,N_6951);
or U7198 (N_7198,N_6875,N_6823);
nor U7199 (N_7199,N_6940,N_6972);
nand U7200 (N_7200,N_7072,N_7091);
nand U7201 (N_7201,N_7136,N_7045);
or U7202 (N_7202,N_7040,N_7095);
xnor U7203 (N_7203,N_7033,N_7148);
nand U7204 (N_7204,N_7104,N_7153);
nor U7205 (N_7205,N_7079,N_7083);
nand U7206 (N_7206,N_7180,N_7143);
nand U7207 (N_7207,N_7028,N_7071);
nor U7208 (N_7208,N_7019,N_7139);
nor U7209 (N_7209,N_7081,N_7087);
nor U7210 (N_7210,N_7069,N_7176);
or U7211 (N_7211,N_7170,N_7077);
nor U7212 (N_7212,N_7166,N_7149);
or U7213 (N_7213,N_7175,N_7154);
or U7214 (N_7214,N_7052,N_7080);
nor U7215 (N_7215,N_7043,N_7085);
and U7216 (N_7216,N_7044,N_7185);
nor U7217 (N_7217,N_7165,N_7084);
xor U7218 (N_7218,N_7075,N_7106);
xnor U7219 (N_7219,N_7012,N_7022);
and U7220 (N_7220,N_7112,N_7066);
or U7221 (N_7221,N_7169,N_7163);
nand U7222 (N_7222,N_7096,N_7189);
xnor U7223 (N_7223,N_7046,N_7062);
nor U7224 (N_7224,N_7060,N_7086);
nand U7225 (N_7225,N_7042,N_7172);
xnor U7226 (N_7226,N_7182,N_7032);
or U7227 (N_7227,N_7034,N_7184);
xor U7228 (N_7228,N_7105,N_7097);
xnor U7229 (N_7229,N_7151,N_7199);
nor U7230 (N_7230,N_7132,N_7197);
or U7231 (N_7231,N_7137,N_7050);
and U7232 (N_7232,N_7061,N_7140);
or U7233 (N_7233,N_7101,N_7076);
and U7234 (N_7234,N_7146,N_7002);
or U7235 (N_7235,N_7121,N_7004);
nor U7236 (N_7236,N_7051,N_7018);
nand U7237 (N_7237,N_7026,N_7057);
nand U7238 (N_7238,N_7001,N_7119);
or U7239 (N_7239,N_7025,N_7194);
xor U7240 (N_7240,N_7115,N_7094);
nor U7241 (N_7241,N_7187,N_7054);
or U7242 (N_7242,N_7122,N_7017);
and U7243 (N_7243,N_7183,N_7009);
nand U7244 (N_7244,N_7107,N_7109);
nor U7245 (N_7245,N_7056,N_7053);
nand U7246 (N_7246,N_7098,N_7073);
xor U7247 (N_7247,N_7141,N_7055);
and U7248 (N_7248,N_7015,N_7021);
nand U7249 (N_7249,N_7114,N_7117);
and U7250 (N_7250,N_7047,N_7116);
nand U7251 (N_7251,N_7067,N_7088);
or U7252 (N_7252,N_7171,N_7031);
nor U7253 (N_7253,N_7063,N_7014);
and U7254 (N_7254,N_7005,N_7145);
nand U7255 (N_7255,N_7158,N_7124);
or U7256 (N_7256,N_7036,N_7190);
and U7257 (N_7257,N_7135,N_7192);
and U7258 (N_7258,N_7039,N_7168);
nand U7259 (N_7259,N_7010,N_7173);
xor U7260 (N_7260,N_7130,N_7029);
nand U7261 (N_7261,N_7038,N_7120);
or U7262 (N_7262,N_7089,N_7155);
and U7263 (N_7263,N_7152,N_7160);
and U7264 (N_7264,N_7150,N_7157);
xor U7265 (N_7265,N_7048,N_7131);
or U7266 (N_7266,N_7142,N_7164);
nor U7267 (N_7267,N_7195,N_7006);
xnor U7268 (N_7268,N_7024,N_7161);
nor U7269 (N_7269,N_7147,N_7070);
or U7270 (N_7270,N_7159,N_7059);
xnor U7271 (N_7271,N_7099,N_7126);
nor U7272 (N_7272,N_7196,N_7123);
nand U7273 (N_7273,N_7007,N_7138);
or U7274 (N_7274,N_7092,N_7008);
and U7275 (N_7275,N_7016,N_7003);
nor U7276 (N_7276,N_7167,N_7078);
and U7277 (N_7277,N_7118,N_7134);
nand U7278 (N_7278,N_7041,N_7074);
nor U7279 (N_7279,N_7108,N_7020);
nand U7280 (N_7280,N_7193,N_7191);
xnor U7281 (N_7281,N_7198,N_7188);
xor U7282 (N_7282,N_7000,N_7093);
and U7283 (N_7283,N_7133,N_7162);
and U7284 (N_7284,N_7179,N_7058);
xnor U7285 (N_7285,N_7100,N_7049);
and U7286 (N_7286,N_7068,N_7102);
and U7287 (N_7287,N_7064,N_7037);
nor U7288 (N_7288,N_7065,N_7127);
xnor U7289 (N_7289,N_7129,N_7181);
and U7290 (N_7290,N_7178,N_7013);
nand U7291 (N_7291,N_7113,N_7090);
and U7292 (N_7292,N_7174,N_7177);
nand U7293 (N_7293,N_7030,N_7156);
xor U7294 (N_7294,N_7110,N_7027);
or U7295 (N_7295,N_7144,N_7011);
xnor U7296 (N_7296,N_7023,N_7111);
or U7297 (N_7297,N_7103,N_7186);
nor U7298 (N_7298,N_7035,N_7125);
or U7299 (N_7299,N_7128,N_7082);
and U7300 (N_7300,N_7124,N_7117);
or U7301 (N_7301,N_7147,N_7049);
and U7302 (N_7302,N_7119,N_7151);
xor U7303 (N_7303,N_7017,N_7110);
or U7304 (N_7304,N_7015,N_7165);
or U7305 (N_7305,N_7171,N_7097);
xnor U7306 (N_7306,N_7130,N_7165);
or U7307 (N_7307,N_7180,N_7186);
nor U7308 (N_7308,N_7042,N_7065);
or U7309 (N_7309,N_7084,N_7102);
and U7310 (N_7310,N_7167,N_7014);
nand U7311 (N_7311,N_7057,N_7105);
nor U7312 (N_7312,N_7008,N_7023);
or U7313 (N_7313,N_7058,N_7115);
nor U7314 (N_7314,N_7034,N_7131);
and U7315 (N_7315,N_7057,N_7120);
or U7316 (N_7316,N_7067,N_7111);
xor U7317 (N_7317,N_7009,N_7116);
nor U7318 (N_7318,N_7105,N_7145);
nor U7319 (N_7319,N_7073,N_7145);
or U7320 (N_7320,N_7096,N_7087);
xnor U7321 (N_7321,N_7108,N_7162);
or U7322 (N_7322,N_7147,N_7000);
or U7323 (N_7323,N_7008,N_7075);
xnor U7324 (N_7324,N_7197,N_7035);
xnor U7325 (N_7325,N_7006,N_7129);
xnor U7326 (N_7326,N_7175,N_7076);
nor U7327 (N_7327,N_7074,N_7129);
or U7328 (N_7328,N_7019,N_7073);
nand U7329 (N_7329,N_7014,N_7147);
and U7330 (N_7330,N_7131,N_7122);
nand U7331 (N_7331,N_7008,N_7162);
nand U7332 (N_7332,N_7145,N_7079);
nand U7333 (N_7333,N_7143,N_7134);
xor U7334 (N_7334,N_7073,N_7030);
nand U7335 (N_7335,N_7123,N_7188);
or U7336 (N_7336,N_7060,N_7112);
and U7337 (N_7337,N_7008,N_7067);
xnor U7338 (N_7338,N_7159,N_7132);
or U7339 (N_7339,N_7103,N_7049);
and U7340 (N_7340,N_7097,N_7133);
xnor U7341 (N_7341,N_7133,N_7074);
and U7342 (N_7342,N_7068,N_7024);
and U7343 (N_7343,N_7146,N_7023);
nor U7344 (N_7344,N_7036,N_7161);
nor U7345 (N_7345,N_7087,N_7084);
xor U7346 (N_7346,N_7082,N_7139);
or U7347 (N_7347,N_7029,N_7067);
nand U7348 (N_7348,N_7146,N_7089);
xnor U7349 (N_7349,N_7164,N_7078);
or U7350 (N_7350,N_7062,N_7063);
or U7351 (N_7351,N_7085,N_7184);
xnor U7352 (N_7352,N_7195,N_7111);
nand U7353 (N_7353,N_7096,N_7120);
and U7354 (N_7354,N_7008,N_7177);
xnor U7355 (N_7355,N_7105,N_7051);
nor U7356 (N_7356,N_7053,N_7023);
nor U7357 (N_7357,N_7065,N_7059);
or U7358 (N_7358,N_7194,N_7195);
nand U7359 (N_7359,N_7052,N_7032);
or U7360 (N_7360,N_7044,N_7037);
nor U7361 (N_7361,N_7171,N_7167);
or U7362 (N_7362,N_7071,N_7002);
nor U7363 (N_7363,N_7091,N_7112);
and U7364 (N_7364,N_7114,N_7137);
nor U7365 (N_7365,N_7082,N_7161);
xnor U7366 (N_7366,N_7014,N_7068);
and U7367 (N_7367,N_7163,N_7024);
xnor U7368 (N_7368,N_7052,N_7127);
nand U7369 (N_7369,N_7116,N_7101);
nand U7370 (N_7370,N_7167,N_7187);
nor U7371 (N_7371,N_7024,N_7009);
and U7372 (N_7372,N_7063,N_7188);
xor U7373 (N_7373,N_7083,N_7100);
or U7374 (N_7374,N_7114,N_7154);
nor U7375 (N_7375,N_7025,N_7111);
nor U7376 (N_7376,N_7017,N_7182);
nand U7377 (N_7377,N_7029,N_7160);
or U7378 (N_7378,N_7002,N_7097);
xnor U7379 (N_7379,N_7018,N_7041);
and U7380 (N_7380,N_7110,N_7021);
or U7381 (N_7381,N_7156,N_7199);
nor U7382 (N_7382,N_7186,N_7081);
and U7383 (N_7383,N_7102,N_7195);
nor U7384 (N_7384,N_7148,N_7175);
nor U7385 (N_7385,N_7052,N_7089);
or U7386 (N_7386,N_7104,N_7013);
xnor U7387 (N_7387,N_7180,N_7025);
nor U7388 (N_7388,N_7178,N_7177);
and U7389 (N_7389,N_7025,N_7129);
xor U7390 (N_7390,N_7123,N_7096);
nor U7391 (N_7391,N_7141,N_7129);
xnor U7392 (N_7392,N_7197,N_7008);
nor U7393 (N_7393,N_7022,N_7115);
nor U7394 (N_7394,N_7189,N_7026);
and U7395 (N_7395,N_7116,N_7177);
xor U7396 (N_7396,N_7156,N_7082);
and U7397 (N_7397,N_7070,N_7120);
or U7398 (N_7398,N_7184,N_7078);
or U7399 (N_7399,N_7026,N_7121);
nand U7400 (N_7400,N_7240,N_7353);
xor U7401 (N_7401,N_7289,N_7330);
xor U7402 (N_7402,N_7380,N_7385);
or U7403 (N_7403,N_7360,N_7344);
nand U7404 (N_7404,N_7216,N_7267);
xor U7405 (N_7405,N_7284,N_7341);
nor U7406 (N_7406,N_7224,N_7366);
or U7407 (N_7407,N_7391,N_7227);
nor U7408 (N_7408,N_7221,N_7223);
or U7409 (N_7409,N_7218,N_7246);
xor U7410 (N_7410,N_7364,N_7318);
xnor U7411 (N_7411,N_7258,N_7348);
and U7412 (N_7412,N_7354,N_7269);
nand U7413 (N_7413,N_7243,N_7356);
xor U7414 (N_7414,N_7302,N_7307);
nor U7415 (N_7415,N_7395,N_7247);
nor U7416 (N_7416,N_7324,N_7310);
xnor U7417 (N_7417,N_7248,N_7379);
or U7418 (N_7418,N_7278,N_7288);
and U7419 (N_7419,N_7249,N_7371);
nor U7420 (N_7420,N_7349,N_7304);
nor U7421 (N_7421,N_7333,N_7235);
xor U7422 (N_7422,N_7206,N_7337);
or U7423 (N_7423,N_7219,N_7378);
and U7424 (N_7424,N_7351,N_7338);
xor U7425 (N_7425,N_7311,N_7208);
nor U7426 (N_7426,N_7272,N_7386);
and U7427 (N_7427,N_7398,N_7301);
or U7428 (N_7428,N_7239,N_7376);
nand U7429 (N_7429,N_7295,N_7325);
nor U7430 (N_7430,N_7211,N_7375);
xnor U7431 (N_7431,N_7233,N_7222);
nor U7432 (N_7432,N_7260,N_7266);
xor U7433 (N_7433,N_7271,N_7322);
or U7434 (N_7434,N_7382,N_7389);
and U7435 (N_7435,N_7357,N_7290);
nor U7436 (N_7436,N_7207,N_7231);
xor U7437 (N_7437,N_7228,N_7299);
nand U7438 (N_7438,N_7241,N_7226);
xnor U7439 (N_7439,N_7273,N_7372);
nor U7440 (N_7440,N_7369,N_7399);
or U7441 (N_7441,N_7286,N_7257);
or U7442 (N_7442,N_7362,N_7253);
and U7443 (N_7443,N_7204,N_7281);
xnor U7444 (N_7444,N_7323,N_7319);
nand U7445 (N_7445,N_7292,N_7336);
and U7446 (N_7446,N_7205,N_7358);
and U7447 (N_7447,N_7368,N_7268);
nand U7448 (N_7448,N_7236,N_7392);
or U7449 (N_7449,N_7201,N_7237);
and U7450 (N_7450,N_7220,N_7270);
and U7451 (N_7451,N_7328,N_7320);
nor U7452 (N_7452,N_7332,N_7282);
or U7453 (N_7453,N_7234,N_7213);
xor U7454 (N_7454,N_7256,N_7346);
xnor U7455 (N_7455,N_7232,N_7339);
or U7456 (N_7456,N_7264,N_7342);
nand U7457 (N_7457,N_7308,N_7255);
or U7458 (N_7458,N_7277,N_7276);
nor U7459 (N_7459,N_7209,N_7285);
nand U7460 (N_7460,N_7203,N_7335);
nor U7461 (N_7461,N_7293,N_7244);
and U7462 (N_7462,N_7365,N_7200);
nor U7463 (N_7463,N_7230,N_7212);
or U7464 (N_7464,N_7381,N_7396);
or U7465 (N_7465,N_7298,N_7377);
xor U7466 (N_7466,N_7261,N_7259);
xnor U7467 (N_7467,N_7355,N_7210);
nand U7468 (N_7468,N_7397,N_7202);
nor U7469 (N_7469,N_7363,N_7225);
and U7470 (N_7470,N_7314,N_7294);
or U7471 (N_7471,N_7297,N_7312);
and U7472 (N_7472,N_7343,N_7352);
nand U7473 (N_7473,N_7340,N_7217);
xor U7474 (N_7474,N_7242,N_7251);
nand U7475 (N_7475,N_7296,N_7279);
xor U7476 (N_7476,N_7331,N_7374);
nand U7477 (N_7477,N_7274,N_7287);
or U7478 (N_7478,N_7306,N_7316);
nand U7479 (N_7479,N_7327,N_7263);
nor U7480 (N_7480,N_7347,N_7326);
or U7481 (N_7481,N_7214,N_7291);
or U7482 (N_7482,N_7275,N_7252);
or U7483 (N_7483,N_7305,N_7254);
xnor U7484 (N_7484,N_7309,N_7384);
nor U7485 (N_7485,N_7393,N_7370);
or U7486 (N_7486,N_7313,N_7245);
nand U7487 (N_7487,N_7388,N_7373);
xor U7488 (N_7488,N_7321,N_7303);
nand U7489 (N_7489,N_7315,N_7238);
or U7490 (N_7490,N_7280,N_7387);
or U7491 (N_7491,N_7262,N_7229);
and U7492 (N_7492,N_7215,N_7394);
xor U7493 (N_7493,N_7300,N_7283);
nand U7494 (N_7494,N_7367,N_7390);
nor U7495 (N_7495,N_7383,N_7334);
nor U7496 (N_7496,N_7361,N_7350);
or U7497 (N_7497,N_7345,N_7359);
nor U7498 (N_7498,N_7329,N_7265);
nor U7499 (N_7499,N_7317,N_7250);
or U7500 (N_7500,N_7241,N_7382);
or U7501 (N_7501,N_7350,N_7218);
nand U7502 (N_7502,N_7214,N_7213);
nand U7503 (N_7503,N_7222,N_7338);
xor U7504 (N_7504,N_7344,N_7261);
xnor U7505 (N_7505,N_7271,N_7335);
or U7506 (N_7506,N_7231,N_7312);
and U7507 (N_7507,N_7286,N_7303);
xor U7508 (N_7508,N_7305,N_7319);
nand U7509 (N_7509,N_7379,N_7382);
nand U7510 (N_7510,N_7336,N_7274);
nor U7511 (N_7511,N_7222,N_7368);
or U7512 (N_7512,N_7367,N_7259);
xor U7513 (N_7513,N_7379,N_7387);
and U7514 (N_7514,N_7275,N_7261);
or U7515 (N_7515,N_7381,N_7329);
and U7516 (N_7516,N_7299,N_7223);
or U7517 (N_7517,N_7379,N_7314);
nand U7518 (N_7518,N_7387,N_7357);
and U7519 (N_7519,N_7272,N_7321);
xor U7520 (N_7520,N_7259,N_7394);
nand U7521 (N_7521,N_7297,N_7386);
and U7522 (N_7522,N_7344,N_7297);
xor U7523 (N_7523,N_7225,N_7311);
or U7524 (N_7524,N_7255,N_7322);
xnor U7525 (N_7525,N_7248,N_7398);
and U7526 (N_7526,N_7286,N_7332);
xnor U7527 (N_7527,N_7232,N_7266);
nand U7528 (N_7528,N_7358,N_7395);
or U7529 (N_7529,N_7307,N_7246);
xor U7530 (N_7530,N_7234,N_7231);
and U7531 (N_7531,N_7334,N_7306);
xor U7532 (N_7532,N_7325,N_7228);
and U7533 (N_7533,N_7319,N_7308);
or U7534 (N_7534,N_7302,N_7309);
nand U7535 (N_7535,N_7289,N_7224);
or U7536 (N_7536,N_7246,N_7297);
or U7537 (N_7537,N_7215,N_7288);
xor U7538 (N_7538,N_7250,N_7268);
nand U7539 (N_7539,N_7206,N_7324);
and U7540 (N_7540,N_7350,N_7206);
nor U7541 (N_7541,N_7393,N_7279);
or U7542 (N_7542,N_7219,N_7321);
xnor U7543 (N_7543,N_7314,N_7289);
or U7544 (N_7544,N_7222,N_7321);
xnor U7545 (N_7545,N_7277,N_7203);
nand U7546 (N_7546,N_7280,N_7313);
nand U7547 (N_7547,N_7393,N_7291);
nor U7548 (N_7548,N_7230,N_7222);
or U7549 (N_7549,N_7377,N_7203);
xor U7550 (N_7550,N_7301,N_7323);
or U7551 (N_7551,N_7348,N_7280);
nand U7552 (N_7552,N_7393,N_7352);
nand U7553 (N_7553,N_7218,N_7278);
nand U7554 (N_7554,N_7240,N_7290);
nor U7555 (N_7555,N_7248,N_7395);
or U7556 (N_7556,N_7348,N_7207);
nor U7557 (N_7557,N_7205,N_7230);
nand U7558 (N_7558,N_7305,N_7253);
nor U7559 (N_7559,N_7252,N_7256);
xor U7560 (N_7560,N_7305,N_7287);
nor U7561 (N_7561,N_7255,N_7246);
or U7562 (N_7562,N_7396,N_7345);
nor U7563 (N_7563,N_7282,N_7226);
or U7564 (N_7564,N_7268,N_7205);
nand U7565 (N_7565,N_7205,N_7312);
nand U7566 (N_7566,N_7331,N_7275);
nor U7567 (N_7567,N_7305,N_7271);
and U7568 (N_7568,N_7354,N_7247);
and U7569 (N_7569,N_7301,N_7262);
nor U7570 (N_7570,N_7352,N_7222);
nand U7571 (N_7571,N_7273,N_7260);
xor U7572 (N_7572,N_7211,N_7338);
and U7573 (N_7573,N_7286,N_7234);
or U7574 (N_7574,N_7250,N_7292);
nand U7575 (N_7575,N_7238,N_7324);
xor U7576 (N_7576,N_7280,N_7223);
nor U7577 (N_7577,N_7320,N_7204);
nor U7578 (N_7578,N_7326,N_7246);
nand U7579 (N_7579,N_7396,N_7346);
and U7580 (N_7580,N_7303,N_7272);
nand U7581 (N_7581,N_7378,N_7276);
or U7582 (N_7582,N_7397,N_7373);
nand U7583 (N_7583,N_7242,N_7359);
xor U7584 (N_7584,N_7390,N_7203);
or U7585 (N_7585,N_7289,N_7382);
nor U7586 (N_7586,N_7278,N_7225);
and U7587 (N_7587,N_7349,N_7339);
or U7588 (N_7588,N_7395,N_7296);
or U7589 (N_7589,N_7207,N_7324);
and U7590 (N_7590,N_7388,N_7240);
or U7591 (N_7591,N_7369,N_7233);
xor U7592 (N_7592,N_7287,N_7326);
nand U7593 (N_7593,N_7308,N_7369);
nor U7594 (N_7594,N_7304,N_7388);
and U7595 (N_7595,N_7270,N_7238);
xor U7596 (N_7596,N_7383,N_7374);
nor U7597 (N_7597,N_7241,N_7383);
or U7598 (N_7598,N_7369,N_7327);
nand U7599 (N_7599,N_7361,N_7365);
and U7600 (N_7600,N_7405,N_7487);
and U7601 (N_7601,N_7479,N_7582);
nor U7602 (N_7602,N_7588,N_7411);
xor U7603 (N_7603,N_7587,N_7508);
or U7604 (N_7604,N_7501,N_7570);
and U7605 (N_7605,N_7591,N_7447);
or U7606 (N_7606,N_7518,N_7435);
and U7607 (N_7607,N_7482,N_7412);
xor U7608 (N_7608,N_7503,N_7516);
or U7609 (N_7609,N_7598,N_7509);
or U7610 (N_7610,N_7415,N_7549);
nor U7611 (N_7611,N_7421,N_7504);
xnor U7612 (N_7612,N_7586,N_7440);
nor U7613 (N_7613,N_7523,N_7420);
xor U7614 (N_7614,N_7510,N_7595);
or U7615 (N_7615,N_7417,N_7481);
nor U7616 (N_7616,N_7414,N_7454);
nand U7617 (N_7617,N_7490,N_7455);
and U7618 (N_7618,N_7429,N_7497);
and U7619 (N_7619,N_7558,N_7538);
and U7620 (N_7620,N_7521,N_7584);
nor U7621 (N_7621,N_7541,N_7571);
nand U7622 (N_7622,N_7577,N_7542);
nand U7623 (N_7623,N_7581,N_7484);
xnor U7624 (N_7624,N_7574,N_7453);
nor U7625 (N_7625,N_7513,N_7562);
and U7626 (N_7626,N_7597,N_7400);
and U7627 (N_7627,N_7404,N_7526);
or U7628 (N_7628,N_7529,N_7568);
and U7629 (N_7629,N_7443,N_7572);
or U7630 (N_7630,N_7536,N_7528);
or U7631 (N_7631,N_7451,N_7520);
nand U7632 (N_7632,N_7459,N_7486);
and U7633 (N_7633,N_7410,N_7456);
or U7634 (N_7634,N_7553,N_7580);
xnor U7635 (N_7635,N_7458,N_7550);
or U7636 (N_7636,N_7496,N_7579);
or U7637 (N_7637,N_7533,N_7556);
nor U7638 (N_7638,N_7439,N_7507);
and U7639 (N_7639,N_7476,N_7555);
and U7640 (N_7640,N_7431,N_7422);
xnor U7641 (N_7641,N_7480,N_7448);
or U7642 (N_7642,N_7511,N_7475);
xnor U7643 (N_7643,N_7530,N_7428);
nor U7644 (N_7644,N_7467,N_7423);
xor U7645 (N_7645,N_7464,N_7534);
and U7646 (N_7646,N_7444,N_7547);
and U7647 (N_7647,N_7540,N_7418);
nor U7648 (N_7648,N_7543,N_7514);
and U7649 (N_7649,N_7519,N_7596);
and U7650 (N_7650,N_7485,N_7407);
and U7651 (N_7651,N_7499,N_7567);
or U7652 (N_7652,N_7537,N_7468);
xnor U7653 (N_7653,N_7470,N_7413);
nor U7654 (N_7654,N_7594,N_7452);
xor U7655 (N_7655,N_7546,N_7491);
nand U7656 (N_7656,N_7446,N_7522);
and U7657 (N_7657,N_7564,N_7563);
xnor U7658 (N_7658,N_7460,N_7576);
nand U7659 (N_7659,N_7474,N_7436);
nor U7660 (N_7660,N_7472,N_7416);
nand U7661 (N_7661,N_7461,N_7599);
nand U7662 (N_7662,N_7560,N_7495);
nor U7663 (N_7663,N_7544,N_7593);
and U7664 (N_7664,N_7442,N_7573);
and U7665 (N_7665,N_7438,N_7477);
nor U7666 (N_7666,N_7424,N_7465);
or U7667 (N_7667,N_7515,N_7483);
nand U7668 (N_7668,N_7441,N_7432);
xor U7669 (N_7669,N_7589,N_7489);
xnor U7670 (N_7670,N_7450,N_7434);
nand U7671 (N_7671,N_7531,N_7437);
nor U7672 (N_7672,N_7505,N_7539);
or U7673 (N_7673,N_7426,N_7561);
or U7674 (N_7674,N_7527,N_7578);
nand U7675 (N_7675,N_7506,N_7552);
xnor U7676 (N_7676,N_7466,N_7535);
nor U7677 (N_7677,N_7569,N_7524);
xnor U7678 (N_7678,N_7427,N_7502);
and U7679 (N_7679,N_7430,N_7402);
or U7680 (N_7680,N_7449,N_7512);
and U7681 (N_7681,N_7492,N_7532);
nor U7682 (N_7682,N_7565,N_7463);
or U7683 (N_7683,N_7575,N_7548);
nand U7684 (N_7684,N_7557,N_7592);
nand U7685 (N_7685,N_7457,N_7583);
and U7686 (N_7686,N_7471,N_7488);
and U7687 (N_7687,N_7478,N_7559);
nand U7688 (N_7688,N_7498,N_7462);
and U7689 (N_7689,N_7419,N_7473);
and U7690 (N_7690,N_7408,N_7517);
and U7691 (N_7691,N_7433,N_7525);
nor U7692 (N_7692,N_7494,N_7585);
and U7693 (N_7693,N_7409,N_7469);
and U7694 (N_7694,N_7551,N_7566);
nand U7695 (N_7695,N_7401,N_7445);
xor U7696 (N_7696,N_7554,N_7500);
nand U7697 (N_7697,N_7590,N_7403);
nand U7698 (N_7698,N_7425,N_7493);
or U7699 (N_7699,N_7406,N_7545);
nor U7700 (N_7700,N_7481,N_7495);
xor U7701 (N_7701,N_7466,N_7503);
or U7702 (N_7702,N_7591,N_7501);
nand U7703 (N_7703,N_7556,N_7532);
nand U7704 (N_7704,N_7551,N_7446);
nor U7705 (N_7705,N_7411,N_7415);
xor U7706 (N_7706,N_7417,N_7525);
nand U7707 (N_7707,N_7549,N_7590);
nor U7708 (N_7708,N_7456,N_7406);
xor U7709 (N_7709,N_7442,N_7585);
nand U7710 (N_7710,N_7402,N_7491);
nand U7711 (N_7711,N_7446,N_7539);
xor U7712 (N_7712,N_7590,N_7436);
nor U7713 (N_7713,N_7472,N_7535);
xnor U7714 (N_7714,N_7459,N_7481);
nor U7715 (N_7715,N_7440,N_7505);
xor U7716 (N_7716,N_7562,N_7525);
nor U7717 (N_7717,N_7584,N_7520);
xnor U7718 (N_7718,N_7453,N_7520);
nor U7719 (N_7719,N_7428,N_7417);
nor U7720 (N_7720,N_7521,N_7530);
nor U7721 (N_7721,N_7539,N_7589);
xnor U7722 (N_7722,N_7465,N_7520);
and U7723 (N_7723,N_7583,N_7571);
xnor U7724 (N_7724,N_7511,N_7411);
nand U7725 (N_7725,N_7562,N_7568);
or U7726 (N_7726,N_7402,N_7463);
xor U7727 (N_7727,N_7436,N_7475);
nor U7728 (N_7728,N_7440,N_7409);
and U7729 (N_7729,N_7523,N_7444);
or U7730 (N_7730,N_7591,N_7445);
nand U7731 (N_7731,N_7436,N_7518);
nor U7732 (N_7732,N_7482,N_7508);
or U7733 (N_7733,N_7464,N_7537);
or U7734 (N_7734,N_7508,N_7544);
nand U7735 (N_7735,N_7429,N_7528);
xor U7736 (N_7736,N_7473,N_7474);
nand U7737 (N_7737,N_7456,N_7422);
nand U7738 (N_7738,N_7418,N_7427);
or U7739 (N_7739,N_7585,N_7518);
xnor U7740 (N_7740,N_7417,N_7465);
nor U7741 (N_7741,N_7466,N_7509);
nand U7742 (N_7742,N_7504,N_7430);
and U7743 (N_7743,N_7594,N_7413);
or U7744 (N_7744,N_7595,N_7598);
or U7745 (N_7745,N_7500,N_7580);
xnor U7746 (N_7746,N_7494,N_7506);
nor U7747 (N_7747,N_7463,N_7429);
nand U7748 (N_7748,N_7511,N_7504);
nor U7749 (N_7749,N_7410,N_7467);
nand U7750 (N_7750,N_7486,N_7597);
xor U7751 (N_7751,N_7401,N_7485);
and U7752 (N_7752,N_7532,N_7592);
nand U7753 (N_7753,N_7565,N_7428);
or U7754 (N_7754,N_7438,N_7406);
nor U7755 (N_7755,N_7504,N_7571);
nor U7756 (N_7756,N_7435,N_7450);
xnor U7757 (N_7757,N_7583,N_7415);
xor U7758 (N_7758,N_7572,N_7403);
or U7759 (N_7759,N_7474,N_7457);
nor U7760 (N_7760,N_7594,N_7543);
nor U7761 (N_7761,N_7407,N_7471);
nor U7762 (N_7762,N_7578,N_7407);
and U7763 (N_7763,N_7560,N_7593);
nor U7764 (N_7764,N_7580,N_7443);
or U7765 (N_7765,N_7453,N_7567);
xnor U7766 (N_7766,N_7582,N_7552);
xor U7767 (N_7767,N_7540,N_7484);
and U7768 (N_7768,N_7400,N_7515);
or U7769 (N_7769,N_7509,N_7445);
nand U7770 (N_7770,N_7434,N_7465);
nor U7771 (N_7771,N_7451,N_7556);
nand U7772 (N_7772,N_7503,N_7424);
nand U7773 (N_7773,N_7563,N_7432);
and U7774 (N_7774,N_7404,N_7426);
or U7775 (N_7775,N_7426,N_7498);
nand U7776 (N_7776,N_7448,N_7552);
nand U7777 (N_7777,N_7495,N_7556);
nand U7778 (N_7778,N_7507,N_7579);
or U7779 (N_7779,N_7565,N_7519);
and U7780 (N_7780,N_7503,N_7443);
nand U7781 (N_7781,N_7411,N_7510);
and U7782 (N_7782,N_7501,N_7505);
xnor U7783 (N_7783,N_7462,N_7426);
and U7784 (N_7784,N_7427,N_7430);
xor U7785 (N_7785,N_7476,N_7443);
and U7786 (N_7786,N_7584,N_7452);
xnor U7787 (N_7787,N_7476,N_7523);
or U7788 (N_7788,N_7504,N_7598);
or U7789 (N_7789,N_7405,N_7478);
or U7790 (N_7790,N_7443,N_7567);
or U7791 (N_7791,N_7563,N_7570);
and U7792 (N_7792,N_7595,N_7532);
nand U7793 (N_7793,N_7474,N_7595);
and U7794 (N_7794,N_7560,N_7409);
nor U7795 (N_7795,N_7581,N_7478);
nand U7796 (N_7796,N_7580,N_7400);
nand U7797 (N_7797,N_7443,N_7422);
xnor U7798 (N_7798,N_7540,N_7514);
xor U7799 (N_7799,N_7541,N_7468);
and U7800 (N_7800,N_7760,N_7771);
and U7801 (N_7801,N_7696,N_7708);
or U7802 (N_7802,N_7799,N_7782);
nor U7803 (N_7803,N_7648,N_7661);
nand U7804 (N_7804,N_7740,N_7616);
nor U7805 (N_7805,N_7718,N_7775);
or U7806 (N_7806,N_7652,N_7713);
and U7807 (N_7807,N_7629,N_7654);
xnor U7808 (N_7808,N_7737,N_7780);
and U7809 (N_7809,N_7767,N_7716);
xor U7810 (N_7810,N_7604,N_7777);
and U7811 (N_7811,N_7602,N_7662);
nor U7812 (N_7812,N_7744,N_7660);
or U7813 (N_7813,N_7726,N_7689);
or U7814 (N_7814,N_7626,N_7765);
nand U7815 (N_7815,N_7632,N_7722);
and U7816 (N_7816,N_7634,N_7641);
or U7817 (N_7817,N_7728,N_7768);
nor U7818 (N_7818,N_7693,N_7645);
and U7819 (N_7819,N_7734,N_7720);
and U7820 (N_7820,N_7736,N_7723);
nand U7821 (N_7821,N_7789,N_7677);
and U7822 (N_7822,N_7676,N_7717);
nor U7823 (N_7823,N_7701,N_7738);
or U7824 (N_7824,N_7699,N_7757);
nand U7825 (N_7825,N_7609,N_7621);
nor U7826 (N_7826,N_7637,N_7747);
nor U7827 (N_7827,N_7613,N_7732);
and U7828 (N_7828,N_7715,N_7761);
and U7829 (N_7829,N_7651,N_7608);
or U7830 (N_7830,N_7684,N_7628);
xnor U7831 (N_7831,N_7706,N_7688);
or U7832 (N_7832,N_7749,N_7748);
or U7833 (N_7833,N_7646,N_7638);
or U7834 (N_7834,N_7786,N_7630);
nor U7835 (N_7835,N_7709,N_7611);
xor U7836 (N_7836,N_7750,N_7697);
xor U7837 (N_7837,N_7668,N_7745);
nor U7838 (N_7838,N_7614,N_7791);
and U7839 (N_7839,N_7776,N_7623);
and U7840 (N_7840,N_7653,N_7746);
xor U7841 (N_7841,N_7659,N_7759);
or U7842 (N_7842,N_7779,N_7766);
nor U7843 (N_7843,N_7773,N_7640);
and U7844 (N_7844,N_7612,N_7650);
nand U7845 (N_7845,N_7601,N_7633);
or U7846 (N_7846,N_7698,N_7694);
nand U7847 (N_7847,N_7669,N_7783);
nand U7848 (N_7848,N_7731,N_7673);
nand U7849 (N_7849,N_7670,N_7798);
and U7850 (N_7850,N_7667,N_7664);
nand U7851 (N_7851,N_7756,N_7624);
xor U7852 (N_7852,N_7655,N_7691);
xor U7853 (N_7853,N_7674,N_7785);
nor U7854 (N_7854,N_7649,N_7686);
nor U7855 (N_7855,N_7772,N_7781);
xnor U7856 (N_7856,N_7647,N_7685);
and U7857 (N_7857,N_7663,N_7679);
nor U7858 (N_7858,N_7687,N_7743);
xnor U7859 (N_7859,N_7622,N_7741);
and U7860 (N_7860,N_7603,N_7695);
and U7861 (N_7861,N_7600,N_7636);
nor U7862 (N_7862,N_7755,N_7733);
and U7863 (N_7863,N_7666,N_7619);
or U7864 (N_7864,N_7797,N_7702);
and U7865 (N_7865,N_7784,N_7703);
xor U7866 (N_7866,N_7778,N_7627);
or U7867 (N_7867,N_7704,N_7625);
nand U7868 (N_7868,N_7700,N_7770);
or U7869 (N_7869,N_7721,N_7714);
nand U7870 (N_7870,N_7739,N_7707);
nand U7871 (N_7871,N_7751,N_7793);
or U7872 (N_7872,N_7665,N_7610);
xor U7873 (N_7873,N_7692,N_7711);
or U7874 (N_7874,N_7735,N_7725);
and U7875 (N_7875,N_7795,N_7729);
or U7876 (N_7876,N_7657,N_7787);
and U7877 (N_7877,N_7658,N_7605);
or U7878 (N_7878,N_7792,N_7682);
or U7879 (N_7879,N_7752,N_7671);
nor U7880 (N_7880,N_7642,N_7754);
xor U7881 (N_7881,N_7790,N_7678);
xor U7882 (N_7882,N_7690,N_7617);
xnor U7883 (N_7883,N_7615,N_7675);
and U7884 (N_7884,N_7719,N_7764);
nand U7885 (N_7885,N_7769,N_7794);
and U7886 (N_7886,N_7730,N_7796);
nor U7887 (N_7887,N_7727,N_7680);
nand U7888 (N_7888,N_7774,N_7672);
nand U7889 (N_7889,N_7724,N_7742);
and U7890 (N_7890,N_7753,N_7788);
or U7891 (N_7891,N_7683,N_7618);
nand U7892 (N_7892,N_7644,N_7643);
and U7893 (N_7893,N_7762,N_7639);
xor U7894 (N_7894,N_7712,N_7606);
nor U7895 (N_7895,N_7635,N_7705);
nor U7896 (N_7896,N_7758,N_7656);
and U7897 (N_7897,N_7631,N_7763);
or U7898 (N_7898,N_7681,N_7620);
xnor U7899 (N_7899,N_7710,N_7607);
or U7900 (N_7900,N_7605,N_7634);
xor U7901 (N_7901,N_7774,N_7730);
xnor U7902 (N_7902,N_7695,N_7624);
and U7903 (N_7903,N_7652,N_7667);
or U7904 (N_7904,N_7609,N_7732);
nand U7905 (N_7905,N_7729,N_7761);
nor U7906 (N_7906,N_7722,N_7644);
nor U7907 (N_7907,N_7793,N_7664);
or U7908 (N_7908,N_7680,N_7784);
xor U7909 (N_7909,N_7680,N_7653);
nor U7910 (N_7910,N_7721,N_7780);
nand U7911 (N_7911,N_7644,N_7676);
and U7912 (N_7912,N_7619,N_7679);
and U7913 (N_7913,N_7712,N_7760);
or U7914 (N_7914,N_7726,N_7704);
xnor U7915 (N_7915,N_7699,N_7771);
nor U7916 (N_7916,N_7612,N_7713);
and U7917 (N_7917,N_7769,N_7719);
nand U7918 (N_7918,N_7794,N_7600);
and U7919 (N_7919,N_7608,N_7753);
or U7920 (N_7920,N_7606,N_7764);
xor U7921 (N_7921,N_7622,N_7639);
or U7922 (N_7922,N_7779,N_7778);
xnor U7923 (N_7923,N_7796,N_7631);
and U7924 (N_7924,N_7604,N_7797);
and U7925 (N_7925,N_7748,N_7798);
xnor U7926 (N_7926,N_7685,N_7619);
xor U7927 (N_7927,N_7785,N_7617);
or U7928 (N_7928,N_7770,N_7784);
or U7929 (N_7929,N_7621,N_7702);
nor U7930 (N_7930,N_7730,N_7751);
or U7931 (N_7931,N_7601,N_7659);
nand U7932 (N_7932,N_7702,N_7649);
nor U7933 (N_7933,N_7782,N_7609);
and U7934 (N_7934,N_7729,N_7619);
nor U7935 (N_7935,N_7777,N_7776);
nor U7936 (N_7936,N_7694,N_7610);
nand U7937 (N_7937,N_7759,N_7648);
nor U7938 (N_7938,N_7682,N_7635);
or U7939 (N_7939,N_7647,N_7663);
xor U7940 (N_7940,N_7742,N_7735);
nand U7941 (N_7941,N_7780,N_7631);
and U7942 (N_7942,N_7697,N_7726);
nand U7943 (N_7943,N_7601,N_7694);
nand U7944 (N_7944,N_7660,N_7737);
nor U7945 (N_7945,N_7785,N_7762);
or U7946 (N_7946,N_7663,N_7643);
nand U7947 (N_7947,N_7686,N_7681);
and U7948 (N_7948,N_7735,N_7680);
or U7949 (N_7949,N_7672,N_7681);
nand U7950 (N_7950,N_7740,N_7609);
xnor U7951 (N_7951,N_7684,N_7685);
and U7952 (N_7952,N_7644,N_7762);
nand U7953 (N_7953,N_7640,N_7734);
nand U7954 (N_7954,N_7739,N_7772);
nor U7955 (N_7955,N_7699,N_7659);
xor U7956 (N_7956,N_7618,N_7777);
nand U7957 (N_7957,N_7694,N_7737);
nor U7958 (N_7958,N_7659,N_7744);
xor U7959 (N_7959,N_7616,N_7780);
nor U7960 (N_7960,N_7695,N_7683);
xnor U7961 (N_7961,N_7784,N_7763);
xor U7962 (N_7962,N_7658,N_7688);
xnor U7963 (N_7963,N_7628,N_7735);
nand U7964 (N_7964,N_7607,N_7637);
or U7965 (N_7965,N_7611,N_7688);
nand U7966 (N_7966,N_7665,N_7716);
and U7967 (N_7967,N_7798,N_7733);
nand U7968 (N_7968,N_7761,N_7666);
nand U7969 (N_7969,N_7610,N_7766);
nand U7970 (N_7970,N_7608,N_7741);
or U7971 (N_7971,N_7662,N_7785);
and U7972 (N_7972,N_7722,N_7743);
xor U7973 (N_7973,N_7792,N_7787);
nand U7974 (N_7974,N_7634,N_7612);
or U7975 (N_7975,N_7710,N_7718);
xnor U7976 (N_7976,N_7676,N_7747);
nor U7977 (N_7977,N_7623,N_7768);
xor U7978 (N_7978,N_7765,N_7706);
or U7979 (N_7979,N_7717,N_7651);
and U7980 (N_7980,N_7683,N_7691);
nand U7981 (N_7981,N_7777,N_7786);
nor U7982 (N_7982,N_7615,N_7791);
xnor U7983 (N_7983,N_7770,N_7664);
nor U7984 (N_7984,N_7675,N_7692);
and U7985 (N_7985,N_7786,N_7637);
xor U7986 (N_7986,N_7657,N_7604);
or U7987 (N_7987,N_7733,N_7665);
xnor U7988 (N_7988,N_7793,N_7622);
nand U7989 (N_7989,N_7730,N_7658);
nand U7990 (N_7990,N_7706,N_7692);
xor U7991 (N_7991,N_7764,N_7720);
nand U7992 (N_7992,N_7697,N_7713);
and U7993 (N_7993,N_7685,N_7771);
nand U7994 (N_7994,N_7798,N_7768);
nand U7995 (N_7995,N_7762,N_7635);
xor U7996 (N_7996,N_7693,N_7747);
xnor U7997 (N_7997,N_7721,N_7653);
and U7998 (N_7998,N_7763,N_7762);
and U7999 (N_7999,N_7693,N_7699);
xor U8000 (N_8000,N_7874,N_7977);
nand U8001 (N_8001,N_7959,N_7800);
nand U8002 (N_8002,N_7892,N_7824);
nor U8003 (N_8003,N_7889,N_7913);
or U8004 (N_8004,N_7944,N_7838);
or U8005 (N_8005,N_7962,N_7866);
and U8006 (N_8006,N_7813,N_7832);
xor U8007 (N_8007,N_7958,N_7907);
and U8008 (N_8008,N_7952,N_7965);
nor U8009 (N_8009,N_7950,N_7922);
or U8010 (N_8010,N_7928,N_7815);
and U8011 (N_8011,N_7975,N_7938);
and U8012 (N_8012,N_7893,N_7820);
nor U8013 (N_8013,N_7908,N_7853);
nor U8014 (N_8014,N_7829,N_7859);
nand U8015 (N_8015,N_7926,N_7896);
xnor U8016 (N_8016,N_7803,N_7851);
or U8017 (N_8017,N_7823,N_7826);
xnor U8018 (N_8018,N_7996,N_7894);
xnor U8019 (N_8019,N_7912,N_7854);
nor U8020 (N_8020,N_7917,N_7817);
nor U8021 (N_8021,N_7867,N_7870);
or U8022 (N_8022,N_7953,N_7946);
nand U8023 (N_8023,N_7964,N_7997);
nor U8024 (N_8024,N_7916,N_7970);
nand U8025 (N_8025,N_7807,N_7849);
or U8026 (N_8026,N_7981,N_7985);
nor U8027 (N_8027,N_7895,N_7860);
and U8028 (N_8028,N_7809,N_7973);
xor U8029 (N_8029,N_7819,N_7903);
or U8030 (N_8030,N_7844,N_7841);
nand U8031 (N_8031,N_7871,N_7967);
xor U8032 (N_8032,N_7939,N_7891);
xor U8033 (N_8033,N_7899,N_7877);
xnor U8034 (N_8034,N_7805,N_7811);
and U8035 (N_8035,N_7808,N_7888);
nand U8036 (N_8036,N_7974,N_7995);
nand U8037 (N_8037,N_7992,N_7937);
and U8038 (N_8038,N_7818,N_7918);
xnor U8039 (N_8039,N_7898,N_7986);
or U8040 (N_8040,N_7998,N_7837);
xnor U8041 (N_8041,N_7846,N_7949);
xnor U8042 (N_8042,N_7857,N_7845);
nand U8043 (N_8043,N_7833,N_7827);
and U8044 (N_8044,N_7927,N_7885);
nand U8045 (N_8045,N_7925,N_7910);
and U8046 (N_8046,N_7872,N_7930);
and U8047 (N_8047,N_7887,N_7881);
and U8048 (N_8048,N_7835,N_7929);
or U8049 (N_8049,N_7839,N_7993);
and U8050 (N_8050,N_7951,N_7816);
or U8051 (N_8051,N_7957,N_7904);
nor U8052 (N_8052,N_7842,N_7906);
xnor U8053 (N_8053,N_7982,N_7848);
xor U8054 (N_8054,N_7968,N_7836);
xnor U8055 (N_8055,N_7999,N_7802);
nand U8056 (N_8056,N_7931,N_7932);
xor U8057 (N_8057,N_7915,N_7933);
nand U8058 (N_8058,N_7861,N_7810);
or U8059 (N_8059,N_7976,N_7831);
nand U8060 (N_8060,N_7942,N_7980);
xor U8061 (N_8061,N_7814,N_7840);
and U8062 (N_8062,N_7869,N_7943);
xnor U8063 (N_8063,N_7941,N_7882);
nor U8064 (N_8064,N_7897,N_7905);
xor U8065 (N_8065,N_7945,N_7878);
xor U8066 (N_8066,N_7911,N_7972);
or U8067 (N_8067,N_7960,N_7954);
xor U8068 (N_8068,N_7863,N_7924);
xnor U8069 (N_8069,N_7936,N_7821);
or U8070 (N_8070,N_7804,N_7847);
or U8071 (N_8071,N_7822,N_7855);
and U8072 (N_8072,N_7858,N_7961);
nand U8073 (N_8073,N_7879,N_7948);
xnor U8074 (N_8074,N_7890,N_7990);
xor U8075 (N_8075,N_7963,N_7801);
nand U8076 (N_8076,N_7979,N_7934);
nand U8077 (N_8077,N_7984,N_7884);
and U8078 (N_8078,N_7856,N_7806);
nor U8079 (N_8079,N_7828,N_7880);
xnor U8080 (N_8080,N_7983,N_7988);
and U8081 (N_8081,N_7978,N_7921);
nor U8082 (N_8082,N_7909,N_7902);
nand U8083 (N_8083,N_7843,N_7868);
xor U8084 (N_8084,N_7852,N_7994);
and U8085 (N_8085,N_7830,N_7812);
xnor U8086 (N_8086,N_7923,N_7875);
or U8087 (N_8087,N_7876,N_7991);
or U8088 (N_8088,N_7886,N_7971);
xnor U8089 (N_8089,N_7864,N_7834);
nor U8090 (N_8090,N_7883,N_7862);
nor U8091 (N_8091,N_7873,N_7901);
and U8092 (N_8092,N_7969,N_7914);
or U8093 (N_8093,N_7987,N_7935);
and U8094 (N_8094,N_7865,N_7955);
nor U8095 (N_8095,N_7825,N_7956);
xnor U8096 (N_8096,N_7920,N_7900);
nor U8097 (N_8097,N_7989,N_7947);
xor U8098 (N_8098,N_7940,N_7966);
and U8099 (N_8099,N_7850,N_7919);
nand U8100 (N_8100,N_7951,N_7825);
and U8101 (N_8101,N_7810,N_7868);
or U8102 (N_8102,N_7902,N_7893);
nor U8103 (N_8103,N_7813,N_7917);
or U8104 (N_8104,N_7978,N_7872);
or U8105 (N_8105,N_7861,N_7813);
or U8106 (N_8106,N_7827,N_7893);
xor U8107 (N_8107,N_7922,N_7824);
and U8108 (N_8108,N_7806,N_7847);
nor U8109 (N_8109,N_7900,N_7839);
and U8110 (N_8110,N_7912,N_7887);
nand U8111 (N_8111,N_7860,N_7969);
or U8112 (N_8112,N_7960,N_7856);
xor U8113 (N_8113,N_7961,N_7918);
or U8114 (N_8114,N_7992,N_7832);
nor U8115 (N_8115,N_7953,N_7859);
and U8116 (N_8116,N_7992,N_7855);
xor U8117 (N_8117,N_7905,N_7800);
xor U8118 (N_8118,N_7917,N_7840);
and U8119 (N_8119,N_7941,N_7920);
and U8120 (N_8120,N_7819,N_7927);
or U8121 (N_8121,N_7943,N_7801);
nand U8122 (N_8122,N_7997,N_7854);
nor U8123 (N_8123,N_7958,N_7978);
nand U8124 (N_8124,N_7860,N_7980);
xor U8125 (N_8125,N_7873,N_7853);
and U8126 (N_8126,N_7958,N_7953);
or U8127 (N_8127,N_7838,N_7996);
or U8128 (N_8128,N_7908,N_7805);
nor U8129 (N_8129,N_7819,N_7937);
nor U8130 (N_8130,N_7944,N_7904);
or U8131 (N_8131,N_7920,N_7914);
or U8132 (N_8132,N_7927,N_7860);
nand U8133 (N_8133,N_7892,N_7995);
or U8134 (N_8134,N_7922,N_7802);
xor U8135 (N_8135,N_7972,N_7915);
or U8136 (N_8136,N_7807,N_7891);
xor U8137 (N_8137,N_7807,N_7887);
nor U8138 (N_8138,N_7987,N_7850);
nand U8139 (N_8139,N_7959,N_7932);
and U8140 (N_8140,N_7870,N_7923);
and U8141 (N_8141,N_7818,N_7983);
nand U8142 (N_8142,N_7941,N_7847);
or U8143 (N_8143,N_7977,N_7968);
and U8144 (N_8144,N_7923,N_7825);
or U8145 (N_8145,N_7910,N_7924);
and U8146 (N_8146,N_7878,N_7827);
xor U8147 (N_8147,N_7911,N_7942);
and U8148 (N_8148,N_7950,N_7867);
xor U8149 (N_8149,N_7923,N_7819);
or U8150 (N_8150,N_7902,N_7854);
nand U8151 (N_8151,N_7833,N_7950);
nor U8152 (N_8152,N_7823,N_7877);
nor U8153 (N_8153,N_7974,N_7866);
nor U8154 (N_8154,N_7916,N_7989);
nand U8155 (N_8155,N_7996,N_7910);
or U8156 (N_8156,N_7889,N_7991);
nand U8157 (N_8157,N_7899,N_7855);
xor U8158 (N_8158,N_7919,N_7991);
nor U8159 (N_8159,N_7992,N_7800);
or U8160 (N_8160,N_7986,N_7985);
xor U8161 (N_8161,N_7958,N_7834);
or U8162 (N_8162,N_7995,N_7878);
nor U8163 (N_8163,N_7802,N_7843);
and U8164 (N_8164,N_7877,N_7858);
or U8165 (N_8165,N_7963,N_7824);
nor U8166 (N_8166,N_7846,N_7952);
or U8167 (N_8167,N_7872,N_7818);
xnor U8168 (N_8168,N_7931,N_7940);
and U8169 (N_8169,N_7804,N_7848);
nand U8170 (N_8170,N_7868,N_7884);
nand U8171 (N_8171,N_7895,N_7973);
nor U8172 (N_8172,N_7962,N_7848);
and U8173 (N_8173,N_7894,N_7832);
nand U8174 (N_8174,N_7974,N_7999);
nand U8175 (N_8175,N_7861,N_7926);
and U8176 (N_8176,N_7909,N_7836);
or U8177 (N_8177,N_7816,N_7856);
xnor U8178 (N_8178,N_7870,N_7916);
nor U8179 (N_8179,N_7901,N_7833);
nand U8180 (N_8180,N_7823,N_7929);
or U8181 (N_8181,N_7969,N_7867);
nor U8182 (N_8182,N_7953,N_7954);
and U8183 (N_8183,N_7977,N_7974);
nor U8184 (N_8184,N_7918,N_7820);
nor U8185 (N_8185,N_7854,N_7800);
and U8186 (N_8186,N_7985,N_7864);
or U8187 (N_8187,N_7865,N_7963);
or U8188 (N_8188,N_7816,N_7940);
and U8189 (N_8189,N_7980,N_7842);
nor U8190 (N_8190,N_7939,N_7830);
and U8191 (N_8191,N_7942,N_7826);
nand U8192 (N_8192,N_7912,N_7885);
nor U8193 (N_8193,N_7811,N_7818);
xnor U8194 (N_8194,N_7921,N_7992);
or U8195 (N_8195,N_7956,N_7968);
nor U8196 (N_8196,N_7837,N_7841);
xor U8197 (N_8197,N_7869,N_7981);
or U8198 (N_8198,N_7856,N_7844);
or U8199 (N_8199,N_7924,N_7854);
xnor U8200 (N_8200,N_8116,N_8172);
and U8201 (N_8201,N_8196,N_8126);
xnor U8202 (N_8202,N_8000,N_8088);
and U8203 (N_8203,N_8007,N_8125);
and U8204 (N_8204,N_8193,N_8189);
and U8205 (N_8205,N_8072,N_8122);
nor U8206 (N_8206,N_8142,N_8145);
or U8207 (N_8207,N_8129,N_8131);
xor U8208 (N_8208,N_8030,N_8031);
xor U8209 (N_8209,N_8109,N_8104);
or U8210 (N_8210,N_8026,N_8112);
and U8211 (N_8211,N_8044,N_8182);
or U8212 (N_8212,N_8074,N_8139);
nand U8213 (N_8213,N_8056,N_8093);
or U8214 (N_8214,N_8035,N_8002);
and U8215 (N_8215,N_8071,N_8147);
and U8216 (N_8216,N_8134,N_8014);
nand U8217 (N_8217,N_8005,N_8114);
xor U8218 (N_8218,N_8113,N_8043);
or U8219 (N_8219,N_8190,N_8177);
nand U8220 (N_8220,N_8017,N_8127);
xnor U8221 (N_8221,N_8187,N_8089);
nor U8222 (N_8222,N_8064,N_8060);
or U8223 (N_8223,N_8135,N_8040);
or U8224 (N_8224,N_8012,N_8146);
xor U8225 (N_8225,N_8055,N_8160);
or U8226 (N_8226,N_8132,N_8083);
and U8227 (N_8227,N_8124,N_8161);
nand U8228 (N_8228,N_8198,N_8025);
and U8229 (N_8229,N_8108,N_8174);
or U8230 (N_8230,N_8156,N_8168);
or U8231 (N_8231,N_8118,N_8171);
or U8232 (N_8232,N_8154,N_8021);
nor U8233 (N_8233,N_8049,N_8105);
and U8234 (N_8234,N_8119,N_8117);
or U8235 (N_8235,N_8130,N_8042);
xor U8236 (N_8236,N_8143,N_8167);
or U8237 (N_8237,N_8090,N_8022);
xnor U8238 (N_8238,N_8149,N_8063);
nor U8239 (N_8239,N_8050,N_8151);
nor U8240 (N_8240,N_8033,N_8004);
or U8241 (N_8241,N_8194,N_8184);
and U8242 (N_8242,N_8029,N_8098);
nand U8243 (N_8243,N_8091,N_8065);
nand U8244 (N_8244,N_8183,N_8008);
xor U8245 (N_8245,N_8138,N_8195);
and U8246 (N_8246,N_8045,N_8057);
xor U8247 (N_8247,N_8169,N_8192);
and U8248 (N_8248,N_8013,N_8095);
or U8249 (N_8249,N_8121,N_8164);
and U8250 (N_8250,N_8039,N_8162);
xor U8251 (N_8251,N_8053,N_8062);
xor U8252 (N_8252,N_8067,N_8069);
and U8253 (N_8253,N_8082,N_8123);
or U8254 (N_8254,N_8024,N_8155);
or U8255 (N_8255,N_8041,N_8085);
nand U8256 (N_8256,N_8015,N_8163);
xnor U8257 (N_8257,N_8032,N_8068);
nor U8258 (N_8258,N_8179,N_8188);
and U8259 (N_8259,N_8077,N_8028);
nor U8260 (N_8260,N_8199,N_8128);
xnor U8261 (N_8261,N_8115,N_8166);
xnor U8262 (N_8262,N_8175,N_8019);
and U8263 (N_8263,N_8106,N_8170);
nand U8264 (N_8264,N_8011,N_8101);
or U8265 (N_8265,N_8086,N_8052);
xnor U8266 (N_8266,N_8111,N_8152);
nor U8267 (N_8267,N_8080,N_8159);
nor U8268 (N_8268,N_8165,N_8046);
nand U8269 (N_8269,N_8075,N_8178);
or U8270 (N_8270,N_8191,N_8059);
nor U8271 (N_8271,N_8003,N_8079);
nor U8272 (N_8272,N_8100,N_8150);
or U8273 (N_8273,N_8010,N_8070);
nand U8274 (N_8274,N_8006,N_8137);
nand U8275 (N_8275,N_8001,N_8103);
nand U8276 (N_8276,N_8173,N_8141);
xor U8277 (N_8277,N_8061,N_8096);
nand U8278 (N_8278,N_8054,N_8157);
nor U8279 (N_8279,N_8066,N_8099);
nand U8280 (N_8280,N_8087,N_8153);
xor U8281 (N_8281,N_8009,N_8120);
and U8282 (N_8282,N_8107,N_8027);
or U8283 (N_8283,N_8036,N_8140);
and U8284 (N_8284,N_8076,N_8158);
xor U8285 (N_8285,N_8048,N_8051);
nand U8286 (N_8286,N_8110,N_8037);
or U8287 (N_8287,N_8081,N_8136);
or U8288 (N_8288,N_8018,N_8197);
and U8289 (N_8289,N_8181,N_8176);
nor U8290 (N_8290,N_8047,N_8084);
xor U8291 (N_8291,N_8185,N_8102);
nand U8292 (N_8292,N_8186,N_8034);
or U8293 (N_8293,N_8144,N_8133);
nor U8294 (N_8294,N_8078,N_8058);
nor U8295 (N_8295,N_8020,N_8016);
nor U8296 (N_8296,N_8092,N_8097);
or U8297 (N_8297,N_8094,N_8038);
nand U8298 (N_8298,N_8148,N_8180);
nor U8299 (N_8299,N_8073,N_8023);
nor U8300 (N_8300,N_8109,N_8100);
or U8301 (N_8301,N_8168,N_8100);
nor U8302 (N_8302,N_8047,N_8064);
or U8303 (N_8303,N_8193,N_8014);
nor U8304 (N_8304,N_8027,N_8035);
or U8305 (N_8305,N_8113,N_8198);
or U8306 (N_8306,N_8164,N_8103);
or U8307 (N_8307,N_8154,N_8051);
xor U8308 (N_8308,N_8011,N_8055);
nand U8309 (N_8309,N_8072,N_8098);
nor U8310 (N_8310,N_8159,N_8135);
nand U8311 (N_8311,N_8029,N_8134);
nor U8312 (N_8312,N_8185,N_8110);
xor U8313 (N_8313,N_8073,N_8132);
xor U8314 (N_8314,N_8177,N_8078);
nor U8315 (N_8315,N_8107,N_8161);
or U8316 (N_8316,N_8197,N_8147);
nor U8317 (N_8317,N_8059,N_8069);
or U8318 (N_8318,N_8127,N_8134);
or U8319 (N_8319,N_8118,N_8115);
nor U8320 (N_8320,N_8193,N_8090);
nor U8321 (N_8321,N_8095,N_8118);
and U8322 (N_8322,N_8184,N_8186);
nor U8323 (N_8323,N_8142,N_8127);
nand U8324 (N_8324,N_8183,N_8070);
xnor U8325 (N_8325,N_8052,N_8079);
and U8326 (N_8326,N_8123,N_8163);
nor U8327 (N_8327,N_8090,N_8107);
nand U8328 (N_8328,N_8087,N_8164);
or U8329 (N_8329,N_8025,N_8146);
or U8330 (N_8330,N_8129,N_8080);
nand U8331 (N_8331,N_8003,N_8107);
xnor U8332 (N_8332,N_8192,N_8198);
nand U8333 (N_8333,N_8033,N_8175);
or U8334 (N_8334,N_8110,N_8054);
xor U8335 (N_8335,N_8036,N_8088);
or U8336 (N_8336,N_8170,N_8041);
nor U8337 (N_8337,N_8199,N_8179);
xor U8338 (N_8338,N_8143,N_8157);
and U8339 (N_8339,N_8040,N_8064);
or U8340 (N_8340,N_8079,N_8053);
or U8341 (N_8341,N_8176,N_8099);
xnor U8342 (N_8342,N_8009,N_8157);
and U8343 (N_8343,N_8064,N_8132);
nand U8344 (N_8344,N_8173,N_8043);
nor U8345 (N_8345,N_8122,N_8070);
xnor U8346 (N_8346,N_8160,N_8146);
nor U8347 (N_8347,N_8084,N_8062);
and U8348 (N_8348,N_8167,N_8007);
nand U8349 (N_8349,N_8014,N_8099);
or U8350 (N_8350,N_8041,N_8020);
or U8351 (N_8351,N_8197,N_8162);
nor U8352 (N_8352,N_8027,N_8032);
nor U8353 (N_8353,N_8113,N_8179);
xnor U8354 (N_8354,N_8094,N_8035);
nand U8355 (N_8355,N_8153,N_8094);
or U8356 (N_8356,N_8086,N_8051);
nor U8357 (N_8357,N_8168,N_8127);
xnor U8358 (N_8358,N_8091,N_8115);
nor U8359 (N_8359,N_8174,N_8107);
nor U8360 (N_8360,N_8136,N_8066);
and U8361 (N_8361,N_8187,N_8175);
and U8362 (N_8362,N_8097,N_8060);
or U8363 (N_8363,N_8033,N_8015);
nor U8364 (N_8364,N_8131,N_8119);
xor U8365 (N_8365,N_8011,N_8195);
nand U8366 (N_8366,N_8014,N_8131);
or U8367 (N_8367,N_8185,N_8135);
nand U8368 (N_8368,N_8002,N_8075);
or U8369 (N_8369,N_8061,N_8095);
nand U8370 (N_8370,N_8024,N_8106);
nand U8371 (N_8371,N_8068,N_8072);
xnor U8372 (N_8372,N_8124,N_8189);
and U8373 (N_8373,N_8169,N_8195);
or U8374 (N_8374,N_8140,N_8189);
and U8375 (N_8375,N_8195,N_8153);
xor U8376 (N_8376,N_8098,N_8096);
nand U8377 (N_8377,N_8116,N_8170);
or U8378 (N_8378,N_8195,N_8119);
nor U8379 (N_8379,N_8155,N_8164);
nand U8380 (N_8380,N_8172,N_8095);
xor U8381 (N_8381,N_8041,N_8169);
nand U8382 (N_8382,N_8109,N_8070);
nand U8383 (N_8383,N_8144,N_8029);
nor U8384 (N_8384,N_8009,N_8181);
and U8385 (N_8385,N_8054,N_8005);
nor U8386 (N_8386,N_8134,N_8033);
nand U8387 (N_8387,N_8072,N_8149);
and U8388 (N_8388,N_8040,N_8140);
xor U8389 (N_8389,N_8107,N_8187);
nand U8390 (N_8390,N_8196,N_8165);
nand U8391 (N_8391,N_8013,N_8073);
and U8392 (N_8392,N_8108,N_8042);
and U8393 (N_8393,N_8057,N_8180);
and U8394 (N_8394,N_8003,N_8191);
nand U8395 (N_8395,N_8074,N_8134);
nor U8396 (N_8396,N_8078,N_8044);
nand U8397 (N_8397,N_8054,N_8169);
or U8398 (N_8398,N_8089,N_8007);
or U8399 (N_8399,N_8125,N_8086);
nor U8400 (N_8400,N_8328,N_8237);
nor U8401 (N_8401,N_8316,N_8334);
or U8402 (N_8402,N_8214,N_8205);
or U8403 (N_8403,N_8294,N_8275);
or U8404 (N_8404,N_8279,N_8301);
nor U8405 (N_8405,N_8319,N_8272);
nor U8406 (N_8406,N_8253,N_8386);
and U8407 (N_8407,N_8399,N_8336);
and U8408 (N_8408,N_8332,N_8363);
nor U8409 (N_8409,N_8208,N_8267);
nor U8410 (N_8410,N_8255,N_8276);
or U8411 (N_8411,N_8280,N_8360);
xor U8412 (N_8412,N_8317,N_8300);
nor U8413 (N_8413,N_8254,N_8362);
nand U8414 (N_8414,N_8233,N_8221);
xor U8415 (N_8415,N_8384,N_8344);
xor U8416 (N_8416,N_8232,N_8358);
nor U8417 (N_8417,N_8248,N_8296);
or U8418 (N_8418,N_8282,N_8258);
nand U8419 (N_8419,N_8203,N_8241);
nand U8420 (N_8420,N_8343,N_8377);
or U8421 (N_8421,N_8318,N_8326);
and U8422 (N_8422,N_8378,N_8393);
and U8423 (N_8423,N_8329,N_8310);
nor U8424 (N_8424,N_8234,N_8207);
or U8425 (N_8425,N_8307,N_8368);
nand U8426 (N_8426,N_8213,N_8201);
nor U8427 (N_8427,N_8212,N_8298);
nand U8428 (N_8428,N_8284,N_8251);
nand U8429 (N_8429,N_8222,N_8339);
nand U8430 (N_8430,N_8244,N_8229);
and U8431 (N_8431,N_8322,N_8398);
or U8432 (N_8432,N_8261,N_8337);
nor U8433 (N_8433,N_8293,N_8364);
and U8434 (N_8434,N_8256,N_8288);
xnor U8435 (N_8435,N_8395,N_8309);
nor U8436 (N_8436,N_8359,N_8306);
xor U8437 (N_8437,N_8291,N_8320);
or U8438 (N_8438,N_8346,N_8223);
and U8439 (N_8439,N_8313,N_8262);
nand U8440 (N_8440,N_8374,N_8312);
and U8441 (N_8441,N_8246,N_8397);
nand U8442 (N_8442,N_8369,N_8314);
nor U8443 (N_8443,N_8274,N_8373);
nand U8444 (N_8444,N_8392,N_8264);
nand U8445 (N_8445,N_8218,N_8361);
or U8446 (N_8446,N_8224,N_8219);
xnor U8447 (N_8447,N_8270,N_8210);
and U8448 (N_8448,N_8265,N_8348);
nor U8449 (N_8449,N_8257,N_8209);
nand U8450 (N_8450,N_8323,N_8349);
xor U8451 (N_8451,N_8220,N_8236);
xnor U8452 (N_8452,N_8228,N_8305);
or U8453 (N_8453,N_8338,N_8299);
nand U8454 (N_8454,N_8350,N_8394);
nand U8455 (N_8455,N_8324,N_8303);
and U8456 (N_8456,N_8331,N_8297);
or U8457 (N_8457,N_8315,N_8259);
nand U8458 (N_8458,N_8200,N_8281);
xnor U8459 (N_8459,N_8375,N_8240);
nand U8460 (N_8460,N_8330,N_8295);
xor U8461 (N_8461,N_8268,N_8277);
nor U8462 (N_8462,N_8372,N_8242);
or U8463 (N_8463,N_8341,N_8273);
xnor U8464 (N_8464,N_8391,N_8290);
or U8465 (N_8465,N_8204,N_8227);
and U8466 (N_8466,N_8249,N_8216);
and U8467 (N_8467,N_8333,N_8217);
xnor U8468 (N_8468,N_8225,N_8390);
nor U8469 (N_8469,N_8283,N_8380);
nor U8470 (N_8470,N_8206,N_8271);
xor U8471 (N_8471,N_8367,N_8347);
nand U8472 (N_8472,N_8231,N_8289);
and U8473 (N_8473,N_8247,N_8335);
or U8474 (N_8474,N_8355,N_8260);
or U8475 (N_8475,N_8340,N_8357);
or U8476 (N_8476,N_8286,N_8245);
and U8477 (N_8477,N_8252,N_8376);
and U8478 (N_8478,N_8356,N_8387);
nand U8479 (N_8479,N_8287,N_8266);
and U8480 (N_8480,N_8215,N_8389);
and U8481 (N_8481,N_8311,N_8381);
nor U8482 (N_8482,N_8292,N_8285);
or U8483 (N_8483,N_8354,N_8321);
and U8484 (N_8484,N_8243,N_8351);
and U8485 (N_8485,N_8345,N_8352);
nand U8486 (N_8486,N_8383,N_8211);
xor U8487 (N_8487,N_8327,N_8370);
or U8488 (N_8488,N_8278,N_8366);
nand U8489 (N_8489,N_8302,N_8269);
or U8490 (N_8490,N_8385,N_8365);
nor U8491 (N_8491,N_8353,N_8239);
nor U8492 (N_8492,N_8202,N_8263);
nand U8493 (N_8493,N_8379,N_8308);
or U8494 (N_8494,N_8396,N_8382);
nand U8495 (N_8495,N_8250,N_8304);
or U8496 (N_8496,N_8226,N_8230);
nor U8497 (N_8497,N_8235,N_8342);
nand U8498 (N_8498,N_8371,N_8238);
and U8499 (N_8499,N_8388,N_8325);
or U8500 (N_8500,N_8273,N_8382);
and U8501 (N_8501,N_8228,N_8313);
or U8502 (N_8502,N_8367,N_8239);
nor U8503 (N_8503,N_8210,N_8293);
or U8504 (N_8504,N_8366,N_8358);
xor U8505 (N_8505,N_8247,N_8392);
nor U8506 (N_8506,N_8326,N_8301);
nor U8507 (N_8507,N_8201,N_8392);
nor U8508 (N_8508,N_8356,N_8268);
xnor U8509 (N_8509,N_8290,N_8274);
or U8510 (N_8510,N_8324,N_8287);
nand U8511 (N_8511,N_8222,N_8395);
or U8512 (N_8512,N_8205,N_8201);
or U8513 (N_8513,N_8249,N_8228);
or U8514 (N_8514,N_8292,N_8312);
xnor U8515 (N_8515,N_8396,N_8330);
and U8516 (N_8516,N_8295,N_8246);
xor U8517 (N_8517,N_8369,N_8327);
nand U8518 (N_8518,N_8242,N_8362);
nor U8519 (N_8519,N_8375,N_8380);
nand U8520 (N_8520,N_8316,N_8281);
nand U8521 (N_8521,N_8310,N_8242);
nor U8522 (N_8522,N_8328,N_8225);
and U8523 (N_8523,N_8396,N_8315);
and U8524 (N_8524,N_8207,N_8299);
xor U8525 (N_8525,N_8371,N_8274);
nor U8526 (N_8526,N_8299,N_8241);
xor U8527 (N_8527,N_8326,N_8222);
xnor U8528 (N_8528,N_8359,N_8373);
xnor U8529 (N_8529,N_8257,N_8366);
nand U8530 (N_8530,N_8318,N_8377);
nand U8531 (N_8531,N_8309,N_8374);
and U8532 (N_8532,N_8301,N_8374);
xor U8533 (N_8533,N_8265,N_8330);
nand U8534 (N_8534,N_8259,N_8307);
and U8535 (N_8535,N_8339,N_8275);
nand U8536 (N_8536,N_8244,N_8335);
nor U8537 (N_8537,N_8263,N_8302);
and U8538 (N_8538,N_8339,N_8366);
nand U8539 (N_8539,N_8338,N_8357);
nand U8540 (N_8540,N_8241,N_8234);
and U8541 (N_8541,N_8312,N_8207);
xor U8542 (N_8542,N_8296,N_8234);
and U8543 (N_8543,N_8360,N_8295);
or U8544 (N_8544,N_8289,N_8224);
nor U8545 (N_8545,N_8277,N_8221);
xnor U8546 (N_8546,N_8303,N_8342);
or U8547 (N_8547,N_8262,N_8236);
xnor U8548 (N_8548,N_8285,N_8210);
and U8549 (N_8549,N_8314,N_8229);
or U8550 (N_8550,N_8234,N_8311);
or U8551 (N_8551,N_8355,N_8230);
xnor U8552 (N_8552,N_8266,N_8282);
or U8553 (N_8553,N_8261,N_8379);
or U8554 (N_8554,N_8278,N_8383);
nand U8555 (N_8555,N_8240,N_8215);
or U8556 (N_8556,N_8343,N_8203);
and U8557 (N_8557,N_8330,N_8337);
nand U8558 (N_8558,N_8311,N_8269);
or U8559 (N_8559,N_8213,N_8364);
and U8560 (N_8560,N_8209,N_8386);
or U8561 (N_8561,N_8315,N_8201);
xnor U8562 (N_8562,N_8396,N_8227);
nor U8563 (N_8563,N_8365,N_8369);
or U8564 (N_8564,N_8209,N_8283);
or U8565 (N_8565,N_8281,N_8251);
nor U8566 (N_8566,N_8341,N_8388);
xor U8567 (N_8567,N_8372,N_8360);
nand U8568 (N_8568,N_8218,N_8291);
and U8569 (N_8569,N_8231,N_8293);
xor U8570 (N_8570,N_8238,N_8257);
nand U8571 (N_8571,N_8387,N_8273);
xor U8572 (N_8572,N_8242,N_8334);
and U8573 (N_8573,N_8324,N_8222);
nand U8574 (N_8574,N_8311,N_8270);
or U8575 (N_8575,N_8238,N_8309);
nand U8576 (N_8576,N_8264,N_8386);
or U8577 (N_8577,N_8252,N_8298);
nand U8578 (N_8578,N_8320,N_8321);
or U8579 (N_8579,N_8344,N_8359);
and U8580 (N_8580,N_8398,N_8252);
nor U8581 (N_8581,N_8319,N_8318);
nand U8582 (N_8582,N_8329,N_8221);
and U8583 (N_8583,N_8261,N_8274);
xnor U8584 (N_8584,N_8328,N_8205);
nand U8585 (N_8585,N_8352,N_8205);
and U8586 (N_8586,N_8299,N_8305);
nand U8587 (N_8587,N_8306,N_8346);
nor U8588 (N_8588,N_8219,N_8393);
nor U8589 (N_8589,N_8206,N_8371);
nor U8590 (N_8590,N_8273,N_8364);
nand U8591 (N_8591,N_8216,N_8316);
nor U8592 (N_8592,N_8281,N_8226);
and U8593 (N_8593,N_8368,N_8240);
nand U8594 (N_8594,N_8275,N_8245);
nor U8595 (N_8595,N_8222,N_8374);
or U8596 (N_8596,N_8388,N_8369);
nand U8597 (N_8597,N_8346,N_8299);
nor U8598 (N_8598,N_8330,N_8359);
xnor U8599 (N_8599,N_8293,N_8268);
nor U8600 (N_8600,N_8464,N_8444);
or U8601 (N_8601,N_8410,N_8581);
or U8602 (N_8602,N_8407,N_8448);
nor U8603 (N_8603,N_8512,N_8494);
nor U8604 (N_8604,N_8588,N_8405);
nand U8605 (N_8605,N_8576,N_8457);
nor U8606 (N_8606,N_8451,N_8491);
nand U8607 (N_8607,N_8490,N_8557);
xor U8608 (N_8608,N_8470,N_8569);
nor U8609 (N_8609,N_8486,N_8406);
or U8610 (N_8610,N_8511,N_8566);
or U8611 (N_8611,N_8515,N_8475);
and U8612 (N_8612,N_8446,N_8432);
xor U8613 (N_8613,N_8440,N_8596);
or U8614 (N_8614,N_8426,N_8453);
and U8615 (N_8615,N_8528,N_8431);
nand U8616 (N_8616,N_8597,N_8594);
or U8617 (N_8617,N_8516,N_8501);
nand U8618 (N_8618,N_8423,N_8577);
or U8619 (N_8619,N_8415,N_8555);
nor U8620 (N_8620,N_8598,N_8493);
and U8621 (N_8621,N_8531,N_8584);
nand U8622 (N_8622,N_8578,N_8402);
xnor U8623 (N_8623,N_8445,N_8541);
or U8624 (N_8624,N_8537,N_8414);
and U8625 (N_8625,N_8585,N_8489);
nor U8626 (N_8626,N_8590,N_8484);
and U8627 (N_8627,N_8538,N_8458);
xor U8628 (N_8628,N_8556,N_8495);
xor U8629 (N_8629,N_8480,N_8473);
nor U8630 (N_8630,N_8565,N_8403);
nand U8631 (N_8631,N_8504,N_8465);
and U8632 (N_8632,N_8409,N_8467);
nor U8633 (N_8633,N_8466,N_8529);
nor U8634 (N_8634,N_8450,N_8530);
nand U8635 (N_8635,N_8573,N_8424);
xor U8636 (N_8636,N_8505,N_8455);
nor U8637 (N_8637,N_8499,N_8476);
and U8638 (N_8638,N_8582,N_8502);
nand U8639 (N_8639,N_8564,N_8449);
and U8640 (N_8640,N_8519,N_8419);
nor U8641 (N_8641,N_8420,N_8485);
nand U8642 (N_8642,N_8474,N_8553);
xor U8643 (N_8643,N_8593,N_8483);
or U8644 (N_8644,N_8547,N_8524);
and U8645 (N_8645,N_8418,N_8487);
or U8646 (N_8646,N_8412,N_8523);
nand U8647 (N_8647,N_8526,N_8521);
or U8648 (N_8648,N_8401,N_8518);
and U8649 (N_8649,N_8463,N_8514);
xor U8650 (N_8650,N_8575,N_8425);
or U8651 (N_8651,N_8472,N_8429);
nor U8652 (N_8652,N_8545,N_8452);
or U8653 (N_8653,N_8550,N_8535);
xor U8654 (N_8654,N_8548,N_8468);
nor U8655 (N_8655,N_8442,N_8513);
xnor U8656 (N_8656,N_8471,N_8498);
nand U8657 (N_8657,N_8503,N_8542);
nand U8658 (N_8658,N_8427,N_8579);
nand U8659 (N_8659,N_8533,N_8430);
nor U8660 (N_8660,N_8536,N_8544);
nand U8661 (N_8661,N_8534,N_8438);
and U8662 (N_8662,N_8477,N_8560);
and U8663 (N_8663,N_8562,N_8478);
nor U8664 (N_8664,N_8539,N_8587);
and U8665 (N_8665,N_8496,N_8592);
and U8666 (N_8666,N_8558,N_8488);
xor U8667 (N_8667,N_8492,N_8416);
or U8668 (N_8668,N_8561,N_8517);
or U8669 (N_8669,N_8580,N_8589);
xnor U8670 (N_8670,N_8408,N_8479);
nand U8671 (N_8671,N_8583,N_8482);
or U8672 (N_8672,N_8509,N_8552);
and U8673 (N_8673,N_8434,N_8571);
or U8674 (N_8674,N_8568,N_8574);
nor U8675 (N_8675,N_8439,N_8462);
or U8676 (N_8676,N_8549,N_8447);
xnor U8677 (N_8677,N_8563,N_8481);
nor U8678 (N_8678,N_8508,N_8532);
xnor U8679 (N_8679,N_8520,N_8599);
or U8680 (N_8680,N_8400,N_8497);
nand U8681 (N_8681,N_8460,N_8417);
or U8682 (N_8682,N_8404,N_8554);
and U8683 (N_8683,N_8469,N_8522);
and U8684 (N_8684,N_8570,N_8421);
and U8685 (N_8685,N_8436,N_8567);
nor U8686 (N_8686,N_8413,N_8456);
xor U8687 (N_8687,N_8510,N_8437);
xor U8688 (N_8688,N_8595,N_8422);
nor U8689 (N_8689,N_8527,N_8461);
nand U8690 (N_8690,N_8411,N_8428);
nand U8691 (N_8691,N_8500,N_8433);
or U8692 (N_8692,N_8435,N_8559);
and U8693 (N_8693,N_8540,N_8506);
nor U8694 (N_8694,N_8459,N_8525);
nor U8695 (N_8695,N_8546,N_8586);
xnor U8696 (N_8696,N_8454,N_8507);
and U8697 (N_8697,N_8441,N_8551);
nor U8698 (N_8698,N_8543,N_8443);
nor U8699 (N_8699,N_8572,N_8591);
or U8700 (N_8700,N_8514,N_8555);
or U8701 (N_8701,N_8476,N_8587);
and U8702 (N_8702,N_8596,N_8405);
and U8703 (N_8703,N_8503,N_8582);
nand U8704 (N_8704,N_8520,N_8526);
xnor U8705 (N_8705,N_8510,N_8478);
nor U8706 (N_8706,N_8425,N_8424);
and U8707 (N_8707,N_8557,N_8563);
xnor U8708 (N_8708,N_8412,N_8564);
nor U8709 (N_8709,N_8493,N_8535);
nand U8710 (N_8710,N_8564,N_8554);
xor U8711 (N_8711,N_8517,N_8473);
nor U8712 (N_8712,N_8566,N_8494);
and U8713 (N_8713,N_8538,N_8494);
nor U8714 (N_8714,N_8551,N_8429);
or U8715 (N_8715,N_8426,N_8508);
and U8716 (N_8716,N_8522,N_8510);
and U8717 (N_8717,N_8515,N_8473);
xnor U8718 (N_8718,N_8490,N_8454);
xor U8719 (N_8719,N_8505,N_8588);
or U8720 (N_8720,N_8469,N_8563);
nor U8721 (N_8721,N_8508,N_8511);
nand U8722 (N_8722,N_8464,N_8492);
xor U8723 (N_8723,N_8518,N_8427);
nand U8724 (N_8724,N_8556,N_8493);
nand U8725 (N_8725,N_8405,N_8466);
and U8726 (N_8726,N_8571,N_8455);
nor U8727 (N_8727,N_8482,N_8592);
xor U8728 (N_8728,N_8486,N_8484);
or U8729 (N_8729,N_8563,N_8402);
or U8730 (N_8730,N_8433,N_8459);
and U8731 (N_8731,N_8583,N_8413);
xor U8732 (N_8732,N_8521,N_8439);
or U8733 (N_8733,N_8495,N_8428);
or U8734 (N_8734,N_8476,N_8413);
xor U8735 (N_8735,N_8426,N_8504);
nand U8736 (N_8736,N_8557,N_8502);
xnor U8737 (N_8737,N_8453,N_8420);
and U8738 (N_8738,N_8565,N_8504);
nand U8739 (N_8739,N_8414,N_8556);
xnor U8740 (N_8740,N_8588,N_8449);
nand U8741 (N_8741,N_8526,N_8495);
and U8742 (N_8742,N_8480,N_8426);
nand U8743 (N_8743,N_8502,N_8563);
xor U8744 (N_8744,N_8473,N_8463);
and U8745 (N_8745,N_8472,N_8591);
xnor U8746 (N_8746,N_8548,N_8582);
nor U8747 (N_8747,N_8596,N_8532);
nand U8748 (N_8748,N_8549,N_8506);
or U8749 (N_8749,N_8500,N_8587);
and U8750 (N_8750,N_8596,N_8491);
nor U8751 (N_8751,N_8474,N_8560);
xnor U8752 (N_8752,N_8502,N_8535);
xnor U8753 (N_8753,N_8524,N_8404);
nor U8754 (N_8754,N_8469,N_8585);
nor U8755 (N_8755,N_8599,N_8418);
xnor U8756 (N_8756,N_8515,N_8461);
nand U8757 (N_8757,N_8452,N_8470);
and U8758 (N_8758,N_8456,N_8536);
nand U8759 (N_8759,N_8595,N_8532);
nor U8760 (N_8760,N_8405,N_8552);
and U8761 (N_8761,N_8496,N_8492);
nor U8762 (N_8762,N_8502,N_8435);
or U8763 (N_8763,N_8508,N_8568);
xor U8764 (N_8764,N_8540,N_8516);
nand U8765 (N_8765,N_8432,N_8441);
nor U8766 (N_8766,N_8482,N_8401);
and U8767 (N_8767,N_8415,N_8423);
and U8768 (N_8768,N_8591,N_8521);
or U8769 (N_8769,N_8402,N_8531);
xor U8770 (N_8770,N_8485,N_8402);
xnor U8771 (N_8771,N_8426,N_8461);
nor U8772 (N_8772,N_8572,N_8545);
nand U8773 (N_8773,N_8517,N_8433);
xnor U8774 (N_8774,N_8543,N_8569);
or U8775 (N_8775,N_8526,N_8483);
or U8776 (N_8776,N_8522,N_8441);
nand U8777 (N_8777,N_8421,N_8544);
nor U8778 (N_8778,N_8514,N_8570);
xnor U8779 (N_8779,N_8508,N_8557);
xnor U8780 (N_8780,N_8507,N_8595);
xor U8781 (N_8781,N_8525,N_8418);
nand U8782 (N_8782,N_8414,N_8409);
or U8783 (N_8783,N_8543,N_8567);
nand U8784 (N_8784,N_8438,N_8599);
or U8785 (N_8785,N_8563,N_8457);
nand U8786 (N_8786,N_8539,N_8426);
nor U8787 (N_8787,N_8449,N_8418);
and U8788 (N_8788,N_8560,N_8462);
xor U8789 (N_8789,N_8478,N_8447);
and U8790 (N_8790,N_8520,N_8408);
and U8791 (N_8791,N_8567,N_8401);
nand U8792 (N_8792,N_8449,N_8453);
and U8793 (N_8793,N_8426,N_8593);
nand U8794 (N_8794,N_8413,N_8506);
xnor U8795 (N_8795,N_8447,N_8513);
or U8796 (N_8796,N_8437,N_8542);
and U8797 (N_8797,N_8449,N_8556);
nand U8798 (N_8798,N_8463,N_8578);
xor U8799 (N_8799,N_8489,N_8510);
xor U8800 (N_8800,N_8661,N_8621);
nor U8801 (N_8801,N_8715,N_8696);
xnor U8802 (N_8802,N_8607,N_8615);
xor U8803 (N_8803,N_8639,N_8718);
nand U8804 (N_8804,N_8669,N_8641);
xnor U8805 (N_8805,N_8699,N_8774);
xnor U8806 (N_8806,N_8731,N_8740);
nand U8807 (N_8807,N_8690,N_8671);
or U8808 (N_8808,N_8741,N_8609);
nor U8809 (N_8809,N_8706,N_8784);
nor U8810 (N_8810,N_8640,N_8781);
nand U8811 (N_8811,N_8733,N_8724);
and U8812 (N_8812,N_8680,N_8780);
and U8813 (N_8813,N_8771,N_8611);
or U8814 (N_8814,N_8748,N_8701);
nor U8815 (N_8815,N_8704,N_8678);
nor U8816 (N_8816,N_8664,N_8745);
nor U8817 (N_8817,N_8764,N_8676);
nand U8818 (N_8818,N_8684,N_8682);
nor U8819 (N_8819,N_8642,N_8707);
nor U8820 (N_8820,N_8633,N_8666);
xor U8821 (N_8821,N_8747,N_8790);
and U8822 (N_8822,N_8742,N_8672);
and U8823 (N_8823,N_8732,N_8605);
xor U8824 (N_8824,N_8687,N_8758);
nand U8825 (N_8825,N_8726,N_8799);
nor U8826 (N_8826,N_8667,N_8759);
or U8827 (N_8827,N_8779,N_8662);
xor U8828 (N_8828,N_8694,N_8749);
nand U8829 (N_8829,N_8643,N_8651);
or U8830 (N_8830,N_8761,N_8627);
and U8831 (N_8831,N_8735,N_8760);
nand U8832 (N_8832,N_8645,N_8789);
nor U8833 (N_8833,N_8729,N_8616);
and U8834 (N_8834,N_8685,N_8739);
nand U8835 (N_8835,N_8637,N_8751);
nand U8836 (N_8836,N_8711,N_8623);
and U8837 (N_8837,N_8619,N_8673);
or U8838 (N_8838,N_8765,N_8603);
nand U8839 (N_8839,N_8730,N_8757);
nor U8840 (N_8840,N_8743,N_8721);
or U8841 (N_8841,N_8768,N_8670);
nor U8842 (N_8842,N_8752,N_8791);
nor U8843 (N_8843,N_8775,N_8697);
and U8844 (N_8844,N_8700,N_8776);
xnor U8845 (N_8845,N_8796,N_8773);
or U8846 (N_8846,N_8653,N_8798);
xnor U8847 (N_8847,N_8649,N_8770);
nor U8848 (N_8848,N_8652,N_8636);
nor U8849 (N_8849,N_8663,N_8622);
and U8850 (N_8850,N_8675,N_8736);
and U8851 (N_8851,N_8665,N_8785);
or U8852 (N_8852,N_8793,N_8668);
xnor U8853 (N_8853,N_8788,N_8612);
and U8854 (N_8854,N_8755,N_8646);
and U8855 (N_8855,N_8746,N_8604);
xnor U8856 (N_8856,N_8703,N_8769);
xor U8857 (N_8857,N_8650,N_8762);
xor U8858 (N_8858,N_8722,N_8647);
or U8859 (N_8859,N_8705,N_8691);
nand U8860 (N_8860,N_8632,N_8783);
xor U8861 (N_8861,N_8716,N_8602);
nand U8862 (N_8862,N_8689,N_8708);
and U8863 (N_8863,N_8683,N_8756);
nor U8864 (N_8864,N_8608,N_8644);
nand U8865 (N_8865,N_8763,N_8618);
nor U8866 (N_8866,N_8654,N_8631);
and U8867 (N_8867,N_8695,N_8795);
and U8868 (N_8868,N_8766,N_8772);
and U8869 (N_8869,N_8734,N_8629);
xor U8870 (N_8870,N_8625,N_8606);
nor U8871 (N_8871,N_8738,N_8717);
nand U8872 (N_8872,N_8600,N_8648);
nor U8873 (N_8873,N_8767,N_8712);
nand U8874 (N_8874,N_8725,N_8709);
nand U8875 (N_8875,N_8728,N_8679);
nor U8876 (N_8876,N_8744,N_8681);
or U8877 (N_8877,N_8713,N_8754);
xor U8878 (N_8878,N_8659,N_8794);
nor U8879 (N_8879,N_8660,N_8624);
nand U8880 (N_8880,N_8714,N_8720);
or U8881 (N_8881,N_8686,N_8656);
nor U8882 (N_8882,N_8628,N_8655);
or U8883 (N_8883,N_8727,N_8710);
xor U8884 (N_8884,N_8635,N_8634);
nand U8885 (N_8885,N_8601,N_8626);
xor U8886 (N_8886,N_8778,N_8630);
nor U8887 (N_8887,N_8613,N_8688);
nor U8888 (N_8888,N_8617,N_8750);
nor U8889 (N_8889,N_8797,N_8614);
and U8890 (N_8890,N_8777,N_8658);
nand U8891 (N_8891,N_8638,N_8723);
xor U8892 (N_8892,N_8702,N_8792);
xnor U8893 (N_8893,N_8610,N_8620);
nor U8894 (N_8894,N_8674,N_8698);
nand U8895 (N_8895,N_8657,N_8677);
nand U8896 (N_8896,N_8782,N_8692);
xor U8897 (N_8897,N_8693,N_8737);
and U8898 (N_8898,N_8787,N_8786);
xor U8899 (N_8899,N_8719,N_8753);
nand U8900 (N_8900,N_8613,N_8746);
and U8901 (N_8901,N_8793,N_8789);
and U8902 (N_8902,N_8727,N_8632);
xor U8903 (N_8903,N_8661,N_8715);
or U8904 (N_8904,N_8713,N_8601);
or U8905 (N_8905,N_8683,N_8670);
or U8906 (N_8906,N_8682,N_8600);
nand U8907 (N_8907,N_8743,N_8784);
or U8908 (N_8908,N_8672,N_8700);
or U8909 (N_8909,N_8799,N_8665);
nand U8910 (N_8910,N_8623,N_8726);
and U8911 (N_8911,N_8625,N_8714);
nor U8912 (N_8912,N_8746,N_8630);
xor U8913 (N_8913,N_8684,N_8608);
xor U8914 (N_8914,N_8785,N_8715);
or U8915 (N_8915,N_8663,N_8789);
nor U8916 (N_8916,N_8782,N_8682);
or U8917 (N_8917,N_8795,N_8615);
nor U8918 (N_8918,N_8760,N_8666);
xor U8919 (N_8919,N_8646,N_8643);
nor U8920 (N_8920,N_8640,N_8677);
nor U8921 (N_8921,N_8780,N_8745);
xnor U8922 (N_8922,N_8749,N_8724);
or U8923 (N_8923,N_8688,N_8685);
nand U8924 (N_8924,N_8701,N_8642);
and U8925 (N_8925,N_8787,N_8628);
nor U8926 (N_8926,N_8672,N_8638);
or U8927 (N_8927,N_8697,N_8611);
and U8928 (N_8928,N_8697,N_8619);
or U8929 (N_8929,N_8719,N_8718);
nand U8930 (N_8930,N_8782,N_8648);
nor U8931 (N_8931,N_8683,N_8639);
nor U8932 (N_8932,N_8716,N_8635);
nand U8933 (N_8933,N_8712,N_8689);
xor U8934 (N_8934,N_8690,N_8719);
nor U8935 (N_8935,N_8771,N_8722);
nor U8936 (N_8936,N_8678,N_8762);
nand U8937 (N_8937,N_8605,N_8705);
nor U8938 (N_8938,N_8650,N_8792);
or U8939 (N_8939,N_8702,N_8688);
or U8940 (N_8940,N_8663,N_8696);
xnor U8941 (N_8941,N_8785,N_8673);
xor U8942 (N_8942,N_8705,N_8644);
nor U8943 (N_8943,N_8621,N_8671);
nor U8944 (N_8944,N_8627,N_8640);
nor U8945 (N_8945,N_8666,N_8609);
and U8946 (N_8946,N_8731,N_8720);
and U8947 (N_8947,N_8658,N_8770);
and U8948 (N_8948,N_8784,N_8697);
xnor U8949 (N_8949,N_8606,N_8785);
nor U8950 (N_8950,N_8616,N_8711);
and U8951 (N_8951,N_8674,N_8609);
nand U8952 (N_8952,N_8799,N_8737);
xor U8953 (N_8953,N_8708,N_8643);
and U8954 (N_8954,N_8609,N_8685);
and U8955 (N_8955,N_8707,N_8688);
nor U8956 (N_8956,N_8646,N_8625);
xor U8957 (N_8957,N_8751,N_8710);
nand U8958 (N_8958,N_8753,N_8791);
or U8959 (N_8959,N_8651,N_8646);
or U8960 (N_8960,N_8679,N_8664);
xor U8961 (N_8961,N_8733,N_8691);
nand U8962 (N_8962,N_8692,N_8792);
nand U8963 (N_8963,N_8632,N_8620);
nor U8964 (N_8964,N_8624,N_8618);
or U8965 (N_8965,N_8673,N_8777);
nor U8966 (N_8966,N_8652,N_8795);
xor U8967 (N_8967,N_8628,N_8693);
or U8968 (N_8968,N_8708,N_8665);
nand U8969 (N_8969,N_8797,N_8753);
xnor U8970 (N_8970,N_8737,N_8796);
xnor U8971 (N_8971,N_8635,N_8720);
nand U8972 (N_8972,N_8611,N_8689);
xnor U8973 (N_8973,N_8653,N_8689);
nor U8974 (N_8974,N_8600,N_8705);
xor U8975 (N_8975,N_8787,N_8690);
nor U8976 (N_8976,N_8677,N_8703);
and U8977 (N_8977,N_8776,N_8762);
nor U8978 (N_8978,N_8776,N_8610);
nor U8979 (N_8979,N_8702,N_8765);
nand U8980 (N_8980,N_8731,N_8612);
or U8981 (N_8981,N_8618,N_8787);
and U8982 (N_8982,N_8617,N_8702);
nand U8983 (N_8983,N_8658,N_8668);
nor U8984 (N_8984,N_8782,N_8641);
nor U8985 (N_8985,N_8754,N_8661);
xnor U8986 (N_8986,N_8715,N_8716);
and U8987 (N_8987,N_8744,N_8755);
nand U8988 (N_8988,N_8753,N_8609);
and U8989 (N_8989,N_8612,N_8626);
and U8990 (N_8990,N_8639,N_8728);
nor U8991 (N_8991,N_8666,N_8701);
and U8992 (N_8992,N_8730,N_8610);
nand U8993 (N_8993,N_8699,N_8608);
and U8994 (N_8994,N_8659,N_8650);
and U8995 (N_8995,N_8789,N_8662);
nor U8996 (N_8996,N_8739,N_8693);
xor U8997 (N_8997,N_8740,N_8786);
nor U8998 (N_8998,N_8787,N_8781);
nand U8999 (N_8999,N_8689,N_8789);
or U9000 (N_9000,N_8854,N_8992);
nand U9001 (N_9001,N_8893,N_8882);
and U9002 (N_9002,N_8869,N_8819);
and U9003 (N_9003,N_8946,N_8955);
nor U9004 (N_9004,N_8921,N_8866);
or U9005 (N_9005,N_8836,N_8934);
or U9006 (N_9006,N_8917,N_8896);
xor U9007 (N_9007,N_8802,N_8830);
xor U9008 (N_9008,N_8833,N_8909);
or U9009 (N_9009,N_8990,N_8883);
nor U9010 (N_9010,N_8911,N_8860);
and U9011 (N_9011,N_8863,N_8959);
xnor U9012 (N_9012,N_8899,N_8935);
nor U9013 (N_9013,N_8978,N_8815);
nand U9014 (N_9014,N_8816,N_8903);
and U9015 (N_9015,N_8821,N_8898);
xor U9016 (N_9016,N_8850,N_8969);
nand U9017 (N_9017,N_8993,N_8801);
nor U9018 (N_9018,N_8902,N_8931);
xnor U9019 (N_9019,N_8956,N_8864);
nand U9020 (N_9020,N_8865,N_8929);
xnor U9021 (N_9021,N_8840,N_8939);
nor U9022 (N_9022,N_8800,N_8976);
xor U9023 (N_9023,N_8950,N_8867);
or U9024 (N_9024,N_8835,N_8878);
or U9025 (N_9025,N_8817,N_8940);
xnor U9026 (N_9026,N_8908,N_8843);
nor U9027 (N_9027,N_8960,N_8897);
or U9028 (N_9028,N_8853,N_8822);
and U9029 (N_9029,N_8937,N_8857);
nor U9030 (N_9030,N_8973,N_8888);
xor U9031 (N_9031,N_8998,N_8811);
nand U9032 (N_9032,N_8928,N_8904);
or U9033 (N_9033,N_8871,N_8873);
nor U9034 (N_9034,N_8832,N_8982);
xnor U9035 (N_9035,N_8927,N_8858);
nor U9036 (N_9036,N_8812,N_8831);
and U9037 (N_9037,N_8827,N_8887);
or U9038 (N_9038,N_8846,N_8914);
and U9039 (N_9039,N_8844,N_8979);
xor U9040 (N_9040,N_8974,N_8838);
nand U9041 (N_9041,N_8967,N_8825);
nand U9042 (N_9042,N_8972,N_8834);
and U9043 (N_9043,N_8987,N_8975);
or U9044 (N_9044,N_8926,N_8932);
nor U9045 (N_9045,N_8818,N_8900);
xor U9046 (N_9046,N_8839,N_8848);
or U9047 (N_9047,N_8901,N_8841);
nand U9048 (N_9048,N_8852,N_8813);
or U9049 (N_9049,N_8999,N_8949);
nor U9050 (N_9050,N_8962,N_8954);
xor U9051 (N_9051,N_8820,N_8997);
nor U9052 (N_9052,N_8837,N_8905);
nor U9053 (N_9053,N_8930,N_8913);
nand U9054 (N_9054,N_8925,N_8884);
xor U9055 (N_9055,N_8983,N_8994);
or U9056 (N_9056,N_8910,N_8907);
and U9057 (N_9057,N_8996,N_8951);
and U9058 (N_9058,N_8991,N_8922);
and U9059 (N_9059,N_8906,N_8923);
xor U9060 (N_9060,N_8938,N_8891);
or U9061 (N_9061,N_8958,N_8824);
xnor U9062 (N_9062,N_8814,N_8989);
or U9063 (N_9063,N_8880,N_8804);
nand U9064 (N_9064,N_8879,N_8872);
and U9065 (N_9065,N_8957,N_8868);
nor U9066 (N_9066,N_8933,N_8952);
nor U9067 (N_9067,N_8803,N_8948);
nand U9068 (N_9068,N_8876,N_8826);
xor U9069 (N_9069,N_8963,N_8915);
and U9070 (N_9070,N_8870,N_8851);
or U9071 (N_9071,N_8890,N_8980);
nand U9072 (N_9072,N_8920,N_8855);
nor U9073 (N_9073,N_8845,N_8895);
and U9074 (N_9074,N_8995,N_8968);
or U9075 (N_9075,N_8981,N_8966);
nor U9076 (N_9076,N_8965,N_8861);
nand U9077 (N_9077,N_8808,N_8964);
nand U9078 (N_9078,N_8859,N_8977);
nor U9079 (N_9079,N_8889,N_8807);
or U9080 (N_9080,N_8936,N_8862);
xnor U9081 (N_9081,N_8856,N_8953);
xnor U9082 (N_9082,N_8886,N_8810);
nor U9083 (N_9083,N_8971,N_8942);
xnor U9084 (N_9084,N_8809,N_8894);
and U9085 (N_9085,N_8892,N_8874);
xnor U9086 (N_9086,N_8947,N_8945);
and U9087 (N_9087,N_8877,N_8988);
nand U9088 (N_9088,N_8823,N_8806);
xor U9089 (N_9089,N_8829,N_8943);
and U9090 (N_9090,N_8885,N_8805);
nand U9091 (N_9091,N_8924,N_8912);
nor U9092 (N_9092,N_8875,N_8916);
xnor U9093 (N_9093,N_8985,N_8944);
or U9094 (N_9094,N_8918,N_8847);
xnor U9095 (N_9095,N_8941,N_8842);
xor U9096 (N_9096,N_8984,N_8970);
nand U9097 (N_9097,N_8881,N_8961);
xnor U9098 (N_9098,N_8986,N_8919);
or U9099 (N_9099,N_8849,N_8828);
xnor U9100 (N_9100,N_8846,N_8866);
xor U9101 (N_9101,N_8843,N_8898);
or U9102 (N_9102,N_8953,N_8951);
and U9103 (N_9103,N_8981,N_8961);
or U9104 (N_9104,N_8921,N_8953);
nor U9105 (N_9105,N_8867,N_8879);
nand U9106 (N_9106,N_8913,N_8985);
and U9107 (N_9107,N_8809,N_8945);
or U9108 (N_9108,N_8879,N_8817);
or U9109 (N_9109,N_8873,N_8953);
nor U9110 (N_9110,N_8821,N_8969);
nor U9111 (N_9111,N_8860,N_8882);
xnor U9112 (N_9112,N_8816,N_8813);
xnor U9113 (N_9113,N_8981,N_8852);
xnor U9114 (N_9114,N_8991,N_8973);
nor U9115 (N_9115,N_8947,N_8873);
xnor U9116 (N_9116,N_8964,N_8967);
or U9117 (N_9117,N_8902,N_8963);
nor U9118 (N_9118,N_8825,N_8998);
or U9119 (N_9119,N_8964,N_8897);
nand U9120 (N_9120,N_8817,N_8841);
nor U9121 (N_9121,N_8848,N_8878);
nor U9122 (N_9122,N_8855,N_8935);
nor U9123 (N_9123,N_8901,N_8862);
nand U9124 (N_9124,N_8820,N_8980);
nand U9125 (N_9125,N_8805,N_8972);
xor U9126 (N_9126,N_8883,N_8942);
xor U9127 (N_9127,N_8835,N_8814);
nor U9128 (N_9128,N_8856,N_8977);
or U9129 (N_9129,N_8849,N_8810);
xnor U9130 (N_9130,N_8995,N_8841);
and U9131 (N_9131,N_8948,N_8997);
and U9132 (N_9132,N_8832,N_8830);
and U9133 (N_9133,N_8888,N_8971);
and U9134 (N_9134,N_8827,N_8915);
xnor U9135 (N_9135,N_8869,N_8912);
and U9136 (N_9136,N_8895,N_8864);
nand U9137 (N_9137,N_8845,N_8962);
or U9138 (N_9138,N_8860,N_8909);
and U9139 (N_9139,N_8898,N_8858);
and U9140 (N_9140,N_8988,N_8802);
nand U9141 (N_9141,N_8826,N_8969);
nor U9142 (N_9142,N_8986,N_8806);
xor U9143 (N_9143,N_8811,N_8977);
nor U9144 (N_9144,N_8899,N_8872);
and U9145 (N_9145,N_8903,N_8802);
and U9146 (N_9146,N_8841,N_8883);
xor U9147 (N_9147,N_8805,N_8806);
or U9148 (N_9148,N_8848,N_8828);
xor U9149 (N_9149,N_8923,N_8952);
nand U9150 (N_9150,N_8874,N_8979);
nand U9151 (N_9151,N_8912,N_8824);
nand U9152 (N_9152,N_8931,N_8894);
or U9153 (N_9153,N_8885,N_8974);
nand U9154 (N_9154,N_8979,N_8830);
xnor U9155 (N_9155,N_8964,N_8814);
or U9156 (N_9156,N_8960,N_8909);
nand U9157 (N_9157,N_8924,N_8886);
and U9158 (N_9158,N_8911,N_8938);
or U9159 (N_9159,N_8965,N_8828);
nor U9160 (N_9160,N_8939,N_8865);
or U9161 (N_9161,N_8810,N_8825);
nand U9162 (N_9162,N_8983,N_8908);
xor U9163 (N_9163,N_8806,N_8993);
nand U9164 (N_9164,N_8981,N_8959);
nor U9165 (N_9165,N_8869,N_8928);
nor U9166 (N_9166,N_8844,N_8828);
nand U9167 (N_9167,N_8845,N_8876);
and U9168 (N_9168,N_8978,N_8958);
xnor U9169 (N_9169,N_8954,N_8896);
and U9170 (N_9170,N_8919,N_8960);
and U9171 (N_9171,N_8803,N_8846);
and U9172 (N_9172,N_8942,N_8862);
nand U9173 (N_9173,N_8920,N_8816);
nand U9174 (N_9174,N_8979,N_8930);
nand U9175 (N_9175,N_8927,N_8844);
or U9176 (N_9176,N_8879,N_8942);
xnor U9177 (N_9177,N_8882,N_8846);
or U9178 (N_9178,N_8893,N_8885);
nor U9179 (N_9179,N_8992,N_8843);
xnor U9180 (N_9180,N_8951,N_8974);
xor U9181 (N_9181,N_8945,N_8964);
and U9182 (N_9182,N_8818,N_8927);
or U9183 (N_9183,N_8833,N_8966);
or U9184 (N_9184,N_8825,N_8917);
nand U9185 (N_9185,N_8874,N_8818);
or U9186 (N_9186,N_8891,N_8858);
xnor U9187 (N_9187,N_8848,N_8940);
or U9188 (N_9188,N_8995,N_8922);
nand U9189 (N_9189,N_8838,N_8901);
or U9190 (N_9190,N_8970,N_8944);
or U9191 (N_9191,N_8817,N_8908);
nand U9192 (N_9192,N_8993,N_8956);
xnor U9193 (N_9193,N_8821,N_8932);
xnor U9194 (N_9194,N_8828,N_8898);
and U9195 (N_9195,N_8914,N_8815);
nand U9196 (N_9196,N_8902,N_8997);
nand U9197 (N_9197,N_8870,N_8918);
xnor U9198 (N_9198,N_8851,N_8942);
xor U9199 (N_9199,N_8850,N_8809);
xnor U9200 (N_9200,N_9131,N_9001);
xnor U9201 (N_9201,N_9090,N_9165);
or U9202 (N_9202,N_9034,N_9028);
nand U9203 (N_9203,N_9190,N_9006);
nor U9204 (N_9204,N_9104,N_9149);
and U9205 (N_9205,N_9000,N_9067);
nand U9206 (N_9206,N_9144,N_9089);
and U9207 (N_9207,N_9013,N_9194);
nor U9208 (N_9208,N_9055,N_9022);
and U9209 (N_9209,N_9062,N_9118);
or U9210 (N_9210,N_9075,N_9069);
or U9211 (N_9211,N_9113,N_9170);
xor U9212 (N_9212,N_9093,N_9136);
nand U9213 (N_9213,N_9198,N_9079);
nand U9214 (N_9214,N_9116,N_9180);
nand U9215 (N_9215,N_9066,N_9120);
nor U9216 (N_9216,N_9082,N_9160);
nand U9217 (N_9217,N_9094,N_9157);
nand U9218 (N_9218,N_9138,N_9121);
nor U9219 (N_9219,N_9193,N_9056);
xnor U9220 (N_9220,N_9133,N_9026);
xnor U9221 (N_9221,N_9130,N_9168);
nor U9222 (N_9222,N_9073,N_9112);
xor U9223 (N_9223,N_9105,N_9040);
nor U9224 (N_9224,N_9103,N_9027);
nand U9225 (N_9225,N_9122,N_9123);
nor U9226 (N_9226,N_9057,N_9024);
and U9227 (N_9227,N_9096,N_9020);
and U9228 (N_9228,N_9145,N_9197);
or U9229 (N_9229,N_9183,N_9085);
nor U9230 (N_9230,N_9182,N_9014);
and U9231 (N_9231,N_9010,N_9095);
nand U9232 (N_9232,N_9166,N_9156);
and U9233 (N_9233,N_9011,N_9009);
nand U9234 (N_9234,N_9171,N_9106);
nand U9235 (N_9235,N_9107,N_9036);
nor U9236 (N_9236,N_9155,N_9035);
nor U9237 (N_9237,N_9008,N_9119);
or U9238 (N_9238,N_9100,N_9007);
nor U9239 (N_9239,N_9045,N_9037);
nand U9240 (N_9240,N_9021,N_9049);
nor U9241 (N_9241,N_9172,N_9162);
or U9242 (N_9242,N_9175,N_9101);
or U9243 (N_9243,N_9151,N_9061);
xor U9244 (N_9244,N_9032,N_9152);
xor U9245 (N_9245,N_9132,N_9043);
xnor U9246 (N_9246,N_9063,N_9184);
nor U9247 (N_9247,N_9199,N_9033);
and U9248 (N_9248,N_9059,N_9052);
or U9249 (N_9249,N_9051,N_9046);
nor U9250 (N_9250,N_9139,N_9081);
nand U9251 (N_9251,N_9054,N_9004);
or U9252 (N_9252,N_9091,N_9044);
nand U9253 (N_9253,N_9195,N_9060);
nor U9254 (N_9254,N_9177,N_9047);
and U9255 (N_9255,N_9039,N_9005);
nor U9256 (N_9256,N_9117,N_9186);
nor U9257 (N_9257,N_9111,N_9153);
or U9258 (N_9258,N_9187,N_9072);
nand U9259 (N_9259,N_9108,N_9154);
nor U9260 (N_9260,N_9088,N_9159);
nor U9261 (N_9261,N_9185,N_9053);
nor U9262 (N_9262,N_9140,N_9179);
nand U9263 (N_9263,N_9142,N_9128);
nor U9264 (N_9264,N_9178,N_9109);
nor U9265 (N_9265,N_9124,N_9003);
and U9266 (N_9266,N_9110,N_9023);
or U9267 (N_9267,N_9174,N_9097);
or U9268 (N_9268,N_9076,N_9070);
nor U9269 (N_9269,N_9176,N_9192);
and U9270 (N_9270,N_9012,N_9098);
nand U9271 (N_9271,N_9084,N_9071);
and U9272 (N_9272,N_9181,N_9102);
or U9273 (N_9273,N_9031,N_9016);
and U9274 (N_9274,N_9163,N_9041);
nand U9275 (N_9275,N_9064,N_9025);
and U9276 (N_9276,N_9125,N_9150);
xnor U9277 (N_9277,N_9114,N_9078);
nand U9278 (N_9278,N_9146,N_9188);
and U9279 (N_9279,N_9191,N_9137);
nand U9280 (N_9280,N_9148,N_9029);
nand U9281 (N_9281,N_9196,N_9083);
xnor U9282 (N_9282,N_9092,N_9164);
and U9283 (N_9283,N_9135,N_9080);
nor U9284 (N_9284,N_9169,N_9141);
and U9285 (N_9285,N_9167,N_9030);
and U9286 (N_9286,N_9065,N_9189);
xnor U9287 (N_9287,N_9017,N_9126);
or U9288 (N_9288,N_9086,N_9129);
or U9289 (N_9289,N_9018,N_9127);
nor U9290 (N_9290,N_9158,N_9058);
xor U9291 (N_9291,N_9087,N_9115);
and U9292 (N_9292,N_9015,N_9143);
and U9293 (N_9293,N_9147,N_9099);
xor U9294 (N_9294,N_9134,N_9173);
nor U9295 (N_9295,N_9042,N_9050);
nor U9296 (N_9296,N_9002,N_9074);
nand U9297 (N_9297,N_9019,N_9077);
or U9298 (N_9298,N_9068,N_9048);
or U9299 (N_9299,N_9161,N_9038);
nand U9300 (N_9300,N_9080,N_9078);
nor U9301 (N_9301,N_9129,N_9032);
or U9302 (N_9302,N_9142,N_9037);
or U9303 (N_9303,N_9172,N_9155);
nor U9304 (N_9304,N_9007,N_9118);
nand U9305 (N_9305,N_9166,N_9130);
xnor U9306 (N_9306,N_9046,N_9035);
nand U9307 (N_9307,N_9042,N_9015);
nor U9308 (N_9308,N_9072,N_9068);
or U9309 (N_9309,N_9030,N_9113);
or U9310 (N_9310,N_9063,N_9044);
nand U9311 (N_9311,N_9164,N_9030);
xor U9312 (N_9312,N_9027,N_9052);
nand U9313 (N_9313,N_9094,N_9055);
xnor U9314 (N_9314,N_9119,N_9028);
nand U9315 (N_9315,N_9000,N_9174);
and U9316 (N_9316,N_9092,N_9049);
and U9317 (N_9317,N_9068,N_9190);
and U9318 (N_9318,N_9195,N_9196);
nor U9319 (N_9319,N_9018,N_9173);
nor U9320 (N_9320,N_9026,N_9058);
xor U9321 (N_9321,N_9078,N_9066);
xnor U9322 (N_9322,N_9075,N_9124);
nor U9323 (N_9323,N_9113,N_9020);
nand U9324 (N_9324,N_9040,N_9041);
xor U9325 (N_9325,N_9189,N_9028);
nor U9326 (N_9326,N_9143,N_9037);
nor U9327 (N_9327,N_9105,N_9007);
nor U9328 (N_9328,N_9012,N_9182);
and U9329 (N_9329,N_9137,N_9004);
nand U9330 (N_9330,N_9090,N_9016);
xor U9331 (N_9331,N_9113,N_9166);
nor U9332 (N_9332,N_9137,N_9105);
xor U9333 (N_9333,N_9074,N_9150);
and U9334 (N_9334,N_9088,N_9160);
nand U9335 (N_9335,N_9167,N_9040);
nand U9336 (N_9336,N_9024,N_9144);
nor U9337 (N_9337,N_9178,N_9157);
or U9338 (N_9338,N_9104,N_9003);
or U9339 (N_9339,N_9152,N_9101);
nand U9340 (N_9340,N_9032,N_9115);
nor U9341 (N_9341,N_9140,N_9184);
xnor U9342 (N_9342,N_9139,N_9181);
or U9343 (N_9343,N_9058,N_9040);
xnor U9344 (N_9344,N_9058,N_9138);
or U9345 (N_9345,N_9148,N_9119);
nand U9346 (N_9346,N_9050,N_9018);
or U9347 (N_9347,N_9105,N_9143);
or U9348 (N_9348,N_9102,N_9057);
nor U9349 (N_9349,N_9112,N_9134);
xor U9350 (N_9350,N_9068,N_9199);
or U9351 (N_9351,N_9096,N_9082);
xor U9352 (N_9352,N_9003,N_9145);
nand U9353 (N_9353,N_9028,N_9153);
nand U9354 (N_9354,N_9009,N_9054);
nand U9355 (N_9355,N_9195,N_9062);
nand U9356 (N_9356,N_9054,N_9063);
nor U9357 (N_9357,N_9026,N_9089);
or U9358 (N_9358,N_9157,N_9016);
nand U9359 (N_9359,N_9186,N_9111);
xor U9360 (N_9360,N_9087,N_9038);
or U9361 (N_9361,N_9196,N_9108);
nor U9362 (N_9362,N_9051,N_9121);
or U9363 (N_9363,N_9112,N_9116);
and U9364 (N_9364,N_9076,N_9180);
nand U9365 (N_9365,N_9130,N_9030);
and U9366 (N_9366,N_9161,N_9042);
nand U9367 (N_9367,N_9080,N_9102);
or U9368 (N_9368,N_9127,N_9004);
nand U9369 (N_9369,N_9111,N_9052);
or U9370 (N_9370,N_9176,N_9020);
or U9371 (N_9371,N_9196,N_9166);
or U9372 (N_9372,N_9198,N_9152);
nand U9373 (N_9373,N_9007,N_9155);
or U9374 (N_9374,N_9069,N_9137);
xor U9375 (N_9375,N_9103,N_9186);
or U9376 (N_9376,N_9147,N_9137);
nand U9377 (N_9377,N_9164,N_9178);
nor U9378 (N_9378,N_9130,N_9091);
or U9379 (N_9379,N_9127,N_9168);
xor U9380 (N_9380,N_9126,N_9038);
and U9381 (N_9381,N_9135,N_9120);
or U9382 (N_9382,N_9165,N_9092);
nand U9383 (N_9383,N_9175,N_9086);
or U9384 (N_9384,N_9021,N_9155);
nand U9385 (N_9385,N_9077,N_9120);
or U9386 (N_9386,N_9065,N_9191);
nor U9387 (N_9387,N_9054,N_9192);
nand U9388 (N_9388,N_9082,N_9014);
nor U9389 (N_9389,N_9105,N_9199);
xor U9390 (N_9390,N_9028,N_9151);
nand U9391 (N_9391,N_9005,N_9122);
xnor U9392 (N_9392,N_9036,N_9190);
nand U9393 (N_9393,N_9049,N_9056);
or U9394 (N_9394,N_9085,N_9180);
xnor U9395 (N_9395,N_9026,N_9197);
nand U9396 (N_9396,N_9094,N_9024);
xnor U9397 (N_9397,N_9170,N_9034);
or U9398 (N_9398,N_9131,N_9186);
and U9399 (N_9399,N_9029,N_9066);
xor U9400 (N_9400,N_9308,N_9384);
nand U9401 (N_9401,N_9385,N_9216);
xnor U9402 (N_9402,N_9206,N_9322);
nor U9403 (N_9403,N_9347,N_9200);
nor U9404 (N_9404,N_9369,N_9379);
xnor U9405 (N_9405,N_9215,N_9260);
nand U9406 (N_9406,N_9246,N_9343);
xnor U9407 (N_9407,N_9247,N_9381);
nand U9408 (N_9408,N_9305,N_9386);
nand U9409 (N_9409,N_9396,N_9209);
nor U9410 (N_9410,N_9229,N_9250);
xor U9411 (N_9411,N_9211,N_9208);
or U9412 (N_9412,N_9276,N_9254);
nor U9413 (N_9413,N_9320,N_9226);
and U9414 (N_9414,N_9382,N_9251);
nor U9415 (N_9415,N_9271,N_9397);
nor U9416 (N_9416,N_9335,N_9368);
nand U9417 (N_9417,N_9205,N_9249);
xnor U9418 (N_9418,N_9367,N_9302);
or U9419 (N_9419,N_9275,N_9267);
and U9420 (N_9420,N_9348,N_9314);
xor U9421 (N_9421,N_9277,N_9274);
nand U9422 (N_9422,N_9395,N_9283);
or U9423 (N_9423,N_9350,N_9270);
nand U9424 (N_9424,N_9364,N_9339);
or U9425 (N_9425,N_9374,N_9378);
and U9426 (N_9426,N_9311,N_9312);
xnor U9427 (N_9427,N_9228,N_9316);
or U9428 (N_9428,N_9235,N_9213);
nor U9429 (N_9429,N_9224,N_9220);
or U9430 (N_9430,N_9262,N_9307);
or U9431 (N_9431,N_9344,N_9280);
nor U9432 (N_9432,N_9324,N_9287);
nor U9433 (N_9433,N_9256,N_9393);
nor U9434 (N_9434,N_9399,N_9243);
xor U9435 (N_9435,N_9398,N_9273);
nor U9436 (N_9436,N_9295,N_9303);
or U9437 (N_9437,N_9331,N_9357);
nor U9438 (N_9438,N_9266,N_9351);
xnor U9439 (N_9439,N_9263,N_9244);
nand U9440 (N_9440,N_9334,N_9362);
nor U9441 (N_9441,N_9240,N_9372);
xor U9442 (N_9442,N_9293,N_9317);
or U9443 (N_9443,N_9282,N_9291);
nor U9444 (N_9444,N_9242,N_9297);
and U9445 (N_9445,N_9376,N_9222);
xnor U9446 (N_9446,N_9201,N_9259);
nor U9447 (N_9447,N_9204,N_9325);
xor U9448 (N_9448,N_9341,N_9354);
xnor U9449 (N_9449,N_9365,N_9371);
nor U9450 (N_9450,N_9239,N_9258);
xnor U9451 (N_9451,N_9261,N_9203);
xnor U9452 (N_9452,N_9337,N_9252);
and U9453 (N_9453,N_9284,N_9333);
or U9454 (N_9454,N_9234,N_9321);
and U9455 (N_9455,N_9202,N_9310);
xnor U9456 (N_9456,N_9309,N_9387);
and U9457 (N_9457,N_9377,N_9285);
and U9458 (N_9458,N_9232,N_9214);
nand U9459 (N_9459,N_9373,N_9225);
xnor U9460 (N_9460,N_9352,N_9210);
xor U9461 (N_9461,N_9326,N_9299);
xnor U9462 (N_9462,N_9353,N_9292);
nor U9463 (N_9463,N_9338,N_9319);
and U9464 (N_9464,N_9355,N_9360);
nor U9465 (N_9465,N_9233,N_9392);
and U9466 (N_9466,N_9272,N_9238);
nor U9467 (N_9467,N_9207,N_9346);
and U9468 (N_9468,N_9342,N_9301);
or U9469 (N_9469,N_9332,N_9217);
or U9470 (N_9470,N_9264,N_9300);
xnor U9471 (N_9471,N_9218,N_9230);
nand U9472 (N_9472,N_9288,N_9231);
and U9473 (N_9473,N_9219,N_9340);
nor U9474 (N_9474,N_9390,N_9313);
and U9475 (N_9475,N_9370,N_9236);
nor U9476 (N_9476,N_9294,N_9358);
xnor U9477 (N_9477,N_9265,N_9363);
xor U9478 (N_9478,N_9329,N_9361);
or U9479 (N_9479,N_9327,N_9290);
and U9480 (N_9480,N_9296,N_9279);
nor U9481 (N_9481,N_9253,N_9356);
nand U9482 (N_9482,N_9255,N_9269);
xor U9483 (N_9483,N_9241,N_9389);
or U9484 (N_9484,N_9281,N_9278);
xnor U9485 (N_9485,N_9268,N_9304);
nand U9486 (N_9486,N_9359,N_9328);
and U9487 (N_9487,N_9257,N_9306);
or U9488 (N_9488,N_9227,N_9221);
and U9489 (N_9489,N_9388,N_9212);
and U9490 (N_9490,N_9298,N_9286);
xnor U9491 (N_9491,N_9366,N_9248);
or U9492 (N_9492,N_9336,N_9349);
or U9493 (N_9493,N_9323,N_9237);
nand U9494 (N_9494,N_9245,N_9383);
and U9495 (N_9495,N_9315,N_9318);
nor U9496 (N_9496,N_9345,N_9330);
nor U9497 (N_9497,N_9223,N_9289);
nor U9498 (N_9498,N_9380,N_9391);
nand U9499 (N_9499,N_9375,N_9394);
nor U9500 (N_9500,N_9360,N_9206);
and U9501 (N_9501,N_9327,N_9338);
nand U9502 (N_9502,N_9307,N_9302);
nor U9503 (N_9503,N_9223,N_9320);
or U9504 (N_9504,N_9329,N_9385);
nand U9505 (N_9505,N_9371,N_9222);
and U9506 (N_9506,N_9379,N_9229);
nand U9507 (N_9507,N_9247,N_9220);
or U9508 (N_9508,N_9306,N_9360);
and U9509 (N_9509,N_9278,N_9241);
xnor U9510 (N_9510,N_9365,N_9349);
xnor U9511 (N_9511,N_9367,N_9357);
or U9512 (N_9512,N_9375,N_9288);
and U9513 (N_9513,N_9293,N_9389);
or U9514 (N_9514,N_9226,N_9344);
or U9515 (N_9515,N_9341,N_9309);
or U9516 (N_9516,N_9258,N_9335);
or U9517 (N_9517,N_9341,N_9380);
and U9518 (N_9518,N_9389,N_9315);
xor U9519 (N_9519,N_9240,N_9232);
and U9520 (N_9520,N_9204,N_9251);
or U9521 (N_9521,N_9369,N_9321);
nand U9522 (N_9522,N_9372,N_9253);
xnor U9523 (N_9523,N_9243,N_9248);
xnor U9524 (N_9524,N_9343,N_9250);
and U9525 (N_9525,N_9261,N_9227);
nand U9526 (N_9526,N_9324,N_9303);
and U9527 (N_9527,N_9260,N_9396);
or U9528 (N_9528,N_9359,N_9342);
xor U9529 (N_9529,N_9326,N_9363);
and U9530 (N_9530,N_9375,N_9264);
nand U9531 (N_9531,N_9254,N_9267);
and U9532 (N_9532,N_9216,N_9272);
or U9533 (N_9533,N_9215,N_9360);
and U9534 (N_9534,N_9202,N_9356);
nor U9535 (N_9535,N_9391,N_9265);
xor U9536 (N_9536,N_9255,N_9251);
xor U9537 (N_9537,N_9251,N_9211);
or U9538 (N_9538,N_9383,N_9233);
nor U9539 (N_9539,N_9314,N_9346);
nor U9540 (N_9540,N_9324,N_9356);
nand U9541 (N_9541,N_9246,N_9391);
and U9542 (N_9542,N_9331,N_9399);
and U9543 (N_9543,N_9363,N_9222);
xnor U9544 (N_9544,N_9305,N_9316);
or U9545 (N_9545,N_9399,N_9340);
or U9546 (N_9546,N_9202,N_9230);
nor U9547 (N_9547,N_9278,N_9223);
or U9548 (N_9548,N_9295,N_9280);
or U9549 (N_9549,N_9285,N_9309);
and U9550 (N_9550,N_9325,N_9255);
and U9551 (N_9551,N_9307,N_9373);
or U9552 (N_9552,N_9209,N_9270);
nand U9553 (N_9553,N_9297,N_9395);
or U9554 (N_9554,N_9246,N_9225);
and U9555 (N_9555,N_9266,N_9393);
xor U9556 (N_9556,N_9224,N_9354);
and U9557 (N_9557,N_9356,N_9365);
and U9558 (N_9558,N_9275,N_9232);
nand U9559 (N_9559,N_9206,N_9236);
and U9560 (N_9560,N_9242,N_9355);
and U9561 (N_9561,N_9270,N_9283);
xnor U9562 (N_9562,N_9254,N_9256);
and U9563 (N_9563,N_9367,N_9248);
xor U9564 (N_9564,N_9362,N_9306);
and U9565 (N_9565,N_9393,N_9304);
xnor U9566 (N_9566,N_9360,N_9343);
nand U9567 (N_9567,N_9256,N_9201);
nand U9568 (N_9568,N_9380,N_9265);
nand U9569 (N_9569,N_9267,N_9302);
nand U9570 (N_9570,N_9234,N_9357);
nand U9571 (N_9571,N_9348,N_9399);
and U9572 (N_9572,N_9295,N_9221);
and U9573 (N_9573,N_9275,N_9260);
xor U9574 (N_9574,N_9320,N_9241);
or U9575 (N_9575,N_9325,N_9214);
or U9576 (N_9576,N_9219,N_9373);
xnor U9577 (N_9577,N_9371,N_9211);
xnor U9578 (N_9578,N_9337,N_9277);
and U9579 (N_9579,N_9265,N_9240);
nor U9580 (N_9580,N_9344,N_9274);
and U9581 (N_9581,N_9228,N_9265);
nand U9582 (N_9582,N_9288,N_9264);
or U9583 (N_9583,N_9237,N_9336);
xnor U9584 (N_9584,N_9232,N_9369);
and U9585 (N_9585,N_9280,N_9352);
xor U9586 (N_9586,N_9347,N_9259);
xor U9587 (N_9587,N_9335,N_9206);
nand U9588 (N_9588,N_9335,N_9246);
xnor U9589 (N_9589,N_9210,N_9229);
and U9590 (N_9590,N_9350,N_9313);
xnor U9591 (N_9591,N_9399,N_9382);
and U9592 (N_9592,N_9332,N_9395);
and U9593 (N_9593,N_9242,N_9289);
xnor U9594 (N_9594,N_9340,N_9330);
xor U9595 (N_9595,N_9363,N_9384);
or U9596 (N_9596,N_9244,N_9217);
nand U9597 (N_9597,N_9288,N_9305);
or U9598 (N_9598,N_9256,N_9220);
nor U9599 (N_9599,N_9366,N_9289);
or U9600 (N_9600,N_9421,N_9528);
nand U9601 (N_9601,N_9448,N_9461);
nor U9602 (N_9602,N_9542,N_9581);
xnor U9603 (N_9603,N_9447,N_9456);
and U9604 (N_9604,N_9597,N_9533);
nor U9605 (N_9605,N_9577,N_9426);
and U9606 (N_9606,N_9526,N_9455);
or U9607 (N_9607,N_9407,N_9502);
nand U9608 (N_9608,N_9419,N_9536);
nand U9609 (N_9609,N_9403,N_9532);
nand U9610 (N_9610,N_9452,N_9439);
xor U9611 (N_9611,N_9466,N_9510);
nand U9612 (N_9612,N_9445,N_9595);
nand U9613 (N_9613,N_9563,N_9568);
or U9614 (N_9614,N_9593,N_9443);
nor U9615 (N_9615,N_9404,N_9575);
or U9616 (N_9616,N_9571,N_9566);
nand U9617 (N_9617,N_9497,N_9414);
xnor U9618 (N_9618,N_9406,N_9435);
nor U9619 (N_9619,N_9525,N_9498);
xor U9620 (N_9620,N_9531,N_9440);
xor U9621 (N_9621,N_9586,N_9470);
or U9622 (N_9622,N_9411,N_9583);
or U9623 (N_9623,N_9534,N_9431);
nor U9624 (N_9624,N_9549,N_9505);
xor U9625 (N_9625,N_9541,N_9416);
xnor U9626 (N_9626,N_9500,N_9599);
xor U9627 (N_9627,N_9491,N_9418);
nand U9628 (N_9628,N_9481,N_9441);
nand U9629 (N_9629,N_9468,N_9496);
or U9630 (N_9630,N_9574,N_9430);
nor U9631 (N_9631,N_9592,N_9584);
nand U9632 (N_9632,N_9442,N_9587);
nor U9633 (N_9633,N_9543,N_9567);
xor U9634 (N_9634,N_9508,N_9538);
nor U9635 (N_9635,N_9569,N_9400);
nand U9636 (N_9636,N_9504,N_9450);
or U9637 (N_9637,N_9509,N_9513);
xnor U9638 (N_9638,N_9487,N_9476);
or U9639 (N_9639,N_9486,N_9520);
or U9640 (N_9640,N_9417,N_9515);
or U9641 (N_9641,N_9425,N_9507);
and U9642 (N_9642,N_9449,N_9553);
xor U9643 (N_9643,N_9463,N_9578);
and U9644 (N_9644,N_9588,N_9555);
nand U9645 (N_9645,N_9492,N_9514);
xor U9646 (N_9646,N_9573,N_9557);
or U9647 (N_9647,N_9444,N_9524);
or U9648 (N_9648,N_9482,N_9545);
nand U9649 (N_9649,N_9493,N_9453);
and U9650 (N_9650,N_9576,N_9495);
and U9651 (N_9651,N_9535,N_9519);
nor U9652 (N_9652,N_9518,N_9454);
nor U9653 (N_9653,N_9548,N_9427);
nor U9654 (N_9654,N_9589,N_9562);
and U9655 (N_9655,N_9479,N_9530);
xor U9656 (N_9656,N_9590,N_9483);
and U9657 (N_9657,N_9410,N_9544);
and U9658 (N_9658,N_9517,N_9598);
and U9659 (N_9659,N_9477,N_9499);
nand U9660 (N_9660,N_9484,N_9462);
nor U9661 (N_9661,N_9446,N_9547);
xor U9662 (N_9662,N_9506,N_9488);
xnor U9663 (N_9663,N_9432,N_9436);
nor U9664 (N_9664,N_9550,N_9591);
xor U9665 (N_9665,N_9434,N_9424);
nand U9666 (N_9666,N_9537,N_9478);
and U9667 (N_9667,N_9523,N_9580);
nand U9668 (N_9668,N_9596,N_9511);
nor U9669 (N_9669,N_9554,N_9458);
or U9670 (N_9670,N_9539,N_9420);
nand U9671 (N_9671,N_9494,N_9579);
nand U9672 (N_9672,N_9469,N_9451);
or U9673 (N_9673,N_9570,N_9480);
nor U9674 (N_9674,N_9474,N_9459);
nor U9675 (N_9675,N_9512,N_9422);
nor U9676 (N_9676,N_9561,N_9594);
or U9677 (N_9677,N_9503,N_9582);
or U9678 (N_9678,N_9401,N_9433);
nand U9679 (N_9679,N_9413,N_9428);
nor U9680 (N_9680,N_9529,N_9501);
xnor U9681 (N_9681,N_9437,N_9565);
xor U9682 (N_9682,N_9467,N_9429);
and U9683 (N_9683,N_9521,N_9415);
nor U9684 (N_9684,N_9408,N_9473);
and U9685 (N_9685,N_9490,N_9402);
or U9686 (N_9686,N_9409,N_9559);
xnor U9687 (N_9687,N_9540,N_9438);
nor U9688 (N_9688,N_9558,N_9423);
nor U9689 (N_9689,N_9546,N_9522);
and U9690 (N_9690,N_9516,N_9405);
nor U9691 (N_9691,N_9412,N_9572);
and U9692 (N_9692,N_9564,N_9465);
and U9693 (N_9693,N_9471,N_9585);
and U9694 (N_9694,N_9457,N_9464);
nor U9695 (N_9695,N_9560,N_9472);
nor U9696 (N_9696,N_9460,N_9527);
and U9697 (N_9697,N_9475,N_9552);
nor U9698 (N_9698,N_9551,N_9556);
nor U9699 (N_9699,N_9485,N_9489);
or U9700 (N_9700,N_9551,N_9596);
nor U9701 (N_9701,N_9455,N_9459);
or U9702 (N_9702,N_9513,N_9562);
xor U9703 (N_9703,N_9406,N_9488);
or U9704 (N_9704,N_9590,N_9424);
or U9705 (N_9705,N_9596,N_9413);
xor U9706 (N_9706,N_9571,N_9454);
or U9707 (N_9707,N_9496,N_9566);
nand U9708 (N_9708,N_9542,N_9586);
or U9709 (N_9709,N_9577,N_9405);
and U9710 (N_9710,N_9533,N_9556);
nand U9711 (N_9711,N_9512,N_9510);
and U9712 (N_9712,N_9415,N_9559);
and U9713 (N_9713,N_9581,N_9492);
and U9714 (N_9714,N_9481,N_9456);
nor U9715 (N_9715,N_9422,N_9511);
and U9716 (N_9716,N_9494,N_9581);
xor U9717 (N_9717,N_9515,N_9542);
and U9718 (N_9718,N_9456,N_9582);
or U9719 (N_9719,N_9440,N_9431);
or U9720 (N_9720,N_9499,N_9528);
xor U9721 (N_9721,N_9585,N_9417);
and U9722 (N_9722,N_9534,N_9423);
or U9723 (N_9723,N_9544,N_9574);
xor U9724 (N_9724,N_9458,N_9504);
nand U9725 (N_9725,N_9468,N_9508);
nor U9726 (N_9726,N_9586,N_9599);
nand U9727 (N_9727,N_9484,N_9550);
nor U9728 (N_9728,N_9426,N_9464);
nor U9729 (N_9729,N_9534,N_9577);
nor U9730 (N_9730,N_9530,N_9598);
and U9731 (N_9731,N_9530,N_9415);
and U9732 (N_9732,N_9520,N_9586);
xnor U9733 (N_9733,N_9572,N_9461);
nand U9734 (N_9734,N_9598,N_9415);
nand U9735 (N_9735,N_9431,N_9583);
and U9736 (N_9736,N_9437,N_9408);
nand U9737 (N_9737,N_9440,N_9525);
xnor U9738 (N_9738,N_9589,N_9523);
xnor U9739 (N_9739,N_9431,N_9477);
nor U9740 (N_9740,N_9430,N_9439);
and U9741 (N_9741,N_9483,N_9499);
nor U9742 (N_9742,N_9515,N_9540);
or U9743 (N_9743,N_9448,N_9574);
nor U9744 (N_9744,N_9522,N_9500);
xnor U9745 (N_9745,N_9438,N_9580);
or U9746 (N_9746,N_9543,N_9497);
or U9747 (N_9747,N_9457,N_9437);
or U9748 (N_9748,N_9475,N_9460);
or U9749 (N_9749,N_9457,N_9403);
nand U9750 (N_9750,N_9434,N_9413);
nor U9751 (N_9751,N_9534,N_9476);
and U9752 (N_9752,N_9504,N_9574);
or U9753 (N_9753,N_9476,N_9590);
and U9754 (N_9754,N_9479,N_9457);
nor U9755 (N_9755,N_9446,N_9590);
or U9756 (N_9756,N_9478,N_9534);
nor U9757 (N_9757,N_9508,N_9560);
xnor U9758 (N_9758,N_9551,N_9540);
xor U9759 (N_9759,N_9424,N_9432);
nand U9760 (N_9760,N_9557,N_9592);
nand U9761 (N_9761,N_9547,N_9556);
nand U9762 (N_9762,N_9542,N_9557);
or U9763 (N_9763,N_9554,N_9429);
nor U9764 (N_9764,N_9482,N_9515);
or U9765 (N_9765,N_9448,N_9519);
xnor U9766 (N_9766,N_9437,N_9548);
xnor U9767 (N_9767,N_9402,N_9565);
nor U9768 (N_9768,N_9456,N_9483);
nor U9769 (N_9769,N_9548,N_9506);
nand U9770 (N_9770,N_9553,N_9533);
xnor U9771 (N_9771,N_9477,N_9457);
and U9772 (N_9772,N_9531,N_9421);
nor U9773 (N_9773,N_9510,N_9446);
and U9774 (N_9774,N_9577,N_9436);
nor U9775 (N_9775,N_9538,N_9406);
xor U9776 (N_9776,N_9576,N_9533);
and U9777 (N_9777,N_9480,N_9593);
and U9778 (N_9778,N_9599,N_9468);
xnor U9779 (N_9779,N_9492,N_9419);
or U9780 (N_9780,N_9517,N_9531);
and U9781 (N_9781,N_9514,N_9500);
xnor U9782 (N_9782,N_9426,N_9581);
and U9783 (N_9783,N_9413,N_9488);
xnor U9784 (N_9784,N_9430,N_9567);
or U9785 (N_9785,N_9431,N_9509);
nand U9786 (N_9786,N_9523,N_9525);
nor U9787 (N_9787,N_9472,N_9554);
nand U9788 (N_9788,N_9403,N_9494);
xnor U9789 (N_9789,N_9471,N_9518);
xor U9790 (N_9790,N_9435,N_9559);
nor U9791 (N_9791,N_9567,N_9579);
and U9792 (N_9792,N_9477,N_9448);
nand U9793 (N_9793,N_9483,N_9485);
xor U9794 (N_9794,N_9452,N_9570);
and U9795 (N_9795,N_9526,N_9598);
xor U9796 (N_9796,N_9505,N_9441);
nor U9797 (N_9797,N_9555,N_9481);
and U9798 (N_9798,N_9467,N_9475);
or U9799 (N_9799,N_9548,N_9564);
nor U9800 (N_9800,N_9627,N_9745);
or U9801 (N_9801,N_9684,N_9666);
nand U9802 (N_9802,N_9714,N_9604);
or U9803 (N_9803,N_9648,N_9734);
xnor U9804 (N_9804,N_9699,N_9629);
and U9805 (N_9805,N_9744,N_9774);
or U9806 (N_9806,N_9635,N_9611);
xor U9807 (N_9807,N_9702,N_9689);
nand U9808 (N_9808,N_9783,N_9773);
and U9809 (N_9809,N_9756,N_9697);
or U9810 (N_9810,N_9610,N_9690);
xnor U9811 (N_9811,N_9735,N_9712);
and U9812 (N_9812,N_9638,N_9766);
nor U9813 (N_9813,N_9623,N_9716);
nor U9814 (N_9814,N_9726,N_9797);
xor U9815 (N_9815,N_9780,N_9655);
and U9816 (N_9816,N_9755,N_9705);
xor U9817 (N_9817,N_9752,N_9609);
or U9818 (N_9818,N_9758,N_9622);
nand U9819 (N_9819,N_9748,N_9625);
or U9820 (N_9820,N_9747,N_9796);
nand U9821 (N_9821,N_9672,N_9686);
nor U9822 (N_9822,N_9736,N_9757);
nor U9823 (N_9823,N_9695,N_9651);
nor U9824 (N_9824,N_9637,N_9709);
nand U9825 (N_9825,N_9665,N_9767);
or U9826 (N_9826,N_9606,N_9759);
nand U9827 (N_9827,N_9602,N_9667);
nand U9828 (N_9828,N_9680,N_9663);
and U9829 (N_9829,N_9794,N_9652);
or U9830 (N_9830,N_9704,N_9701);
xnor U9831 (N_9831,N_9643,N_9720);
and U9832 (N_9832,N_9644,N_9742);
nand U9833 (N_9833,N_9787,N_9642);
and U9834 (N_9834,N_9628,N_9673);
nand U9835 (N_9835,N_9683,N_9791);
or U9836 (N_9836,N_9784,N_9750);
xor U9837 (N_9837,N_9723,N_9654);
and U9838 (N_9838,N_9775,N_9799);
or U9839 (N_9839,N_9708,N_9694);
or U9840 (N_9840,N_9614,N_9624);
nand U9841 (N_9841,N_9790,N_9616);
xor U9842 (N_9842,N_9727,N_9731);
or U9843 (N_9843,N_9728,N_9741);
nand U9844 (N_9844,N_9688,N_9786);
or U9845 (N_9845,N_9707,N_9687);
and U9846 (N_9846,N_9678,N_9724);
nand U9847 (N_9847,N_9743,N_9711);
or U9848 (N_9848,N_9658,N_9732);
nand U9849 (N_9849,N_9691,N_9615);
or U9850 (N_9850,N_9785,N_9721);
or U9851 (N_9851,N_9769,N_9782);
nor U9852 (N_9852,N_9659,N_9605);
nand U9853 (N_9853,N_9753,N_9778);
or U9854 (N_9854,N_9675,N_9698);
xnor U9855 (N_9855,N_9657,N_9779);
nor U9856 (N_9856,N_9607,N_9633);
and U9857 (N_9857,N_9647,N_9718);
xnor U9858 (N_9858,N_9660,N_9679);
and U9859 (N_9859,N_9739,N_9781);
and U9860 (N_9860,N_9662,N_9761);
or U9861 (N_9861,N_9612,N_9763);
or U9862 (N_9862,N_9746,N_9608);
nor U9863 (N_9863,N_9600,N_9613);
and U9864 (N_9864,N_9646,N_9703);
or U9865 (N_9865,N_9789,N_9645);
nand U9866 (N_9866,N_9618,N_9661);
and U9867 (N_9867,N_9649,N_9765);
and U9868 (N_9868,N_9674,N_9700);
and U9869 (N_9869,N_9603,N_9715);
nor U9870 (N_9870,N_9617,N_9792);
nor U9871 (N_9871,N_9696,N_9740);
xor U9872 (N_9872,N_9621,N_9771);
and U9873 (N_9873,N_9636,N_9631);
xnor U9874 (N_9874,N_9664,N_9764);
and U9875 (N_9875,N_9762,N_9776);
xor U9876 (N_9876,N_9671,N_9669);
and U9877 (N_9877,N_9733,N_9768);
xnor U9878 (N_9878,N_9737,N_9730);
or U9879 (N_9879,N_9738,N_9706);
xnor U9880 (N_9880,N_9630,N_9681);
nor U9881 (N_9881,N_9793,N_9620);
nand U9882 (N_9882,N_9626,N_9717);
or U9883 (N_9883,N_9754,N_9713);
nand U9884 (N_9884,N_9719,N_9722);
and U9885 (N_9885,N_9685,N_9653);
and U9886 (N_9886,N_9751,N_9772);
and U9887 (N_9887,N_9601,N_9639);
or U9888 (N_9888,N_9668,N_9760);
or U9889 (N_9889,N_9788,N_9641);
and U9890 (N_9890,N_9692,N_9795);
xnor U9891 (N_9891,N_9777,N_9798);
nand U9892 (N_9892,N_9677,N_9729);
nand U9893 (N_9893,N_9632,N_9682);
nor U9894 (N_9894,N_9656,N_9634);
or U9895 (N_9895,N_9710,N_9749);
or U9896 (N_9896,N_9676,N_9770);
nand U9897 (N_9897,N_9619,N_9725);
and U9898 (N_9898,N_9650,N_9693);
xor U9899 (N_9899,N_9670,N_9640);
or U9900 (N_9900,N_9680,N_9679);
and U9901 (N_9901,N_9797,N_9663);
or U9902 (N_9902,N_9655,N_9723);
and U9903 (N_9903,N_9764,N_9635);
or U9904 (N_9904,N_9725,N_9686);
nand U9905 (N_9905,N_9700,N_9652);
xor U9906 (N_9906,N_9666,N_9660);
and U9907 (N_9907,N_9677,N_9689);
or U9908 (N_9908,N_9626,N_9735);
nand U9909 (N_9909,N_9714,N_9728);
nand U9910 (N_9910,N_9708,N_9625);
xor U9911 (N_9911,N_9735,N_9659);
xor U9912 (N_9912,N_9643,N_9695);
nor U9913 (N_9913,N_9676,N_9720);
and U9914 (N_9914,N_9764,N_9756);
or U9915 (N_9915,N_9759,N_9611);
nor U9916 (N_9916,N_9689,N_9645);
nor U9917 (N_9917,N_9646,N_9727);
xor U9918 (N_9918,N_9790,N_9711);
nor U9919 (N_9919,N_9655,N_9732);
nand U9920 (N_9920,N_9607,N_9666);
or U9921 (N_9921,N_9639,N_9673);
nand U9922 (N_9922,N_9704,N_9722);
and U9923 (N_9923,N_9789,N_9736);
and U9924 (N_9924,N_9649,N_9623);
and U9925 (N_9925,N_9632,N_9671);
and U9926 (N_9926,N_9788,N_9655);
nor U9927 (N_9927,N_9654,N_9725);
nand U9928 (N_9928,N_9707,N_9626);
xnor U9929 (N_9929,N_9673,N_9615);
and U9930 (N_9930,N_9756,N_9651);
nand U9931 (N_9931,N_9657,N_9712);
nand U9932 (N_9932,N_9608,N_9775);
xnor U9933 (N_9933,N_9797,N_9635);
or U9934 (N_9934,N_9738,N_9665);
xnor U9935 (N_9935,N_9789,N_9799);
nand U9936 (N_9936,N_9631,N_9766);
or U9937 (N_9937,N_9645,N_9738);
or U9938 (N_9938,N_9644,N_9698);
nand U9939 (N_9939,N_9642,N_9790);
or U9940 (N_9940,N_9672,N_9773);
xnor U9941 (N_9941,N_9785,N_9641);
nand U9942 (N_9942,N_9746,N_9668);
xor U9943 (N_9943,N_9784,N_9743);
nor U9944 (N_9944,N_9792,N_9799);
or U9945 (N_9945,N_9671,N_9691);
nand U9946 (N_9946,N_9728,N_9717);
xor U9947 (N_9947,N_9643,N_9706);
or U9948 (N_9948,N_9779,N_9617);
nand U9949 (N_9949,N_9633,N_9704);
and U9950 (N_9950,N_9761,N_9770);
xor U9951 (N_9951,N_9765,N_9797);
xor U9952 (N_9952,N_9760,N_9610);
nand U9953 (N_9953,N_9718,N_9649);
nor U9954 (N_9954,N_9606,N_9719);
and U9955 (N_9955,N_9719,N_9658);
nand U9956 (N_9956,N_9715,N_9773);
or U9957 (N_9957,N_9662,N_9634);
xnor U9958 (N_9958,N_9608,N_9704);
xnor U9959 (N_9959,N_9750,N_9653);
nand U9960 (N_9960,N_9792,N_9722);
nand U9961 (N_9961,N_9705,N_9643);
or U9962 (N_9962,N_9640,N_9786);
and U9963 (N_9963,N_9773,N_9633);
or U9964 (N_9964,N_9770,N_9793);
nor U9965 (N_9965,N_9743,N_9628);
and U9966 (N_9966,N_9787,N_9672);
or U9967 (N_9967,N_9634,N_9716);
or U9968 (N_9968,N_9799,N_9701);
xor U9969 (N_9969,N_9672,N_9763);
or U9970 (N_9970,N_9798,N_9700);
or U9971 (N_9971,N_9766,N_9686);
xor U9972 (N_9972,N_9705,N_9760);
xnor U9973 (N_9973,N_9793,N_9772);
or U9974 (N_9974,N_9723,N_9766);
and U9975 (N_9975,N_9618,N_9791);
nor U9976 (N_9976,N_9751,N_9660);
nor U9977 (N_9977,N_9642,N_9722);
or U9978 (N_9978,N_9785,N_9768);
or U9979 (N_9979,N_9668,N_9602);
xnor U9980 (N_9980,N_9616,N_9676);
and U9981 (N_9981,N_9625,N_9718);
xor U9982 (N_9982,N_9703,N_9710);
and U9983 (N_9983,N_9698,N_9646);
nand U9984 (N_9984,N_9651,N_9601);
xor U9985 (N_9985,N_9634,N_9746);
nand U9986 (N_9986,N_9636,N_9757);
and U9987 (N_9987,N_9725,N_9798);
nor U9988 (N_9988,N_9679,N_9655);
xor U9989 (N_9989,N_9718,N_9637);
and U9990 (N_9990,N_9758,N_9750);
nand U9991 (N_9991,N_9618,N_9629);
xor U9992 (N_9992,N_9637,N_9756);
and U9993 (N_9993,N_9659,N_9797);
or U9994 (N_9994,N_9688,N_9778);
and U9995 (N_9995,N_9791,N_9610);
nand U9996 (N_9996,N_9790,N_9738);
or U9997 (N_9997,N_9651,N_9638);
and U9998 (N_9998,N_9729,N_9628);
and U9999 (N_9999,N_9749,N_9788);
nand U10000 (N_10000,N_9982,N_9888);
and U10001 (N_10001,N_9912,N_9955);
and U10002 (N_10002,N_9943,N_9842);
or U10003 (N_10003,N_9853,N_9939);
xor U10004 (N_10004,N_9926,N_9855);
and U10005 (N_10005,N_9812,N_9821);
nor U10006 (N_10006,N_9937,N_9995);
nand U10007 (N_10007,N_9971,N_9984);
xor U10008 (N_10008,N_9934,N_9819);
and U10009 (N_10009,N_9991,N_9829);
and U10010 (N_10010,N_9870,N_9845);
nor U10011 (N_10011,N_9807,N_9980);
or U10012 (N_10012,N_9826,N_9999);
or U10013 (N_10013,N_9915,N_9820);
nand U10014 (N_10014,N_9840,N_9814);
nand U10015 (N_10015,N_9871,N_9837);
xnor U10016 (N_10016,N_9886,N_9931);
nand U10017 (N_10017,N_9959,N_9881);
or U10018 (N_10018,N_9909,N_9911);
or U10019 (N_10019,N_9897,N_9811);
and U10020 (N_10020,N_9866,N_9921);
or U10021 (N_10021,N_9856,N_9913);
or U10022 (N_10022,N_9867,N_9816);
nor U10023 (N_10023,N_9832,N_9850);
and U10024 (N_10024,N_9815,N_9876);
or U10025 (N_10025,N_9925,N_9875);
xnor U10026 (N_10026,N_9975,N_9804);
nor U10027 (N_10027,N_9834,N_9877);
xor U10028 (N_10028,N_9802,N_9967);
and U10029 (N_10029,N_9960,N_9849);
or U10030 (N_10030,N_9930,N_9946);
nor U10031 (N_10031,N_9818,N_9803);
or U10032 (N_10032,N_9938,N_9974);
and U10033 (N_10033,N_9806,N_9836);
nor U10034 (N_10034,N_9903,N_9863);
nand U10035 (N_10035,N_9827,N_9882);
nor U10036 (N_10036,N_9981,N_9824);
and U10037 (N_10037,N_9851,N_9823);
or U10038 (N_10038,N_9973,N_9989);
xnor U10039 (N_10039,N_9940,N_9892);
nand U10040 (N_10040,N_9963,N_9987);
nor U10041 (N_10041,N_9904,N_9800);
xor U10042 (N_10042,N_9988,N_9872);
nor U10043 (N_10043,N_9838,N_9906);
and U10044 (N_10044,N_9962,N_9965);
nor U10045 (N_10045,N_9861,N_9890);
nor U10046 (N_10046,N_9922,N_9828);
nor U10047 (N_10047,N_9864,N_9935);
and U10048 (N_10048,N_9964,N_9932);
nand U10049 (N_10049,N_9933,N_9918);
nand U10050 (N_10050,N_9953,N_9862);
and U10051 (N_10051,N_9908,N_9810);
xnor U10052 (N_10052,N_9944,N_9843);
xor U10053 (N_10053,N_9894,N_9978);
or U10054 (N_10054,N_9961,N_9927);
and U10055 (N_10055,N_9868,N_9902);
xnor U10056 (N_10056,N_9801,N_9948);
or U10057 (N_10057,N_9919,N_9994);
xor U10058 (N_10058,N_9972,N_9899);
xor U10059 (N_10059,N_9859,N_9901);
or U10060 (N_10060,N_9969,N_9883);
and U10061 (N_10061,N_9949,N_9896);
nor U10062 (N_10062,N_9952,N_9822);
xor U10063 (N_10063,N_9900,N_9880);
nand U10064 (N_10064,N_9945,N_9905);
xnor U10065 (N_10065,N_9841,N_9986);
and U10066 (N_10066,N_9839,N_9993);
nor U10067 (N_10067,N_9966,N_9929);
or U10068 (N_10068,N_9907,N_9893);
and U10069 (N_10069,N_9898,N_9983);
or U10070 (N_10070,N_9977,N_9809);
nor U10071 (N_10071,N_9885,N_9916);
nand U10072 (N_10072,N_9990,N_9817);
xor U10073 (N_10073,N_9844,N_9954);
nand U10074 (N_10074,N_9928,N_9830);
nor U10075 (N_10075,N_9854,N_9825);
or U10076 (N_10076,N_9847,N_9852);
or U10077 (N_10077,N_9956,N_9968);
nand U10078 (N_10078,N_9805,N_9910);
and U10079 (N_10079,N_9941,N_9958);
or U10080 (N_10080,N_9985,N_9917);
or U10081 (N_10081,N_9950,N_9857);
xor U10082 (N_10082,N_9874,N_9992);
and U10083 (N_10083,N_9808,N_9848);
xnor U10084 (N_10084,N_9884,N_9895);
nor U10085 (N_10085,N_9887,N_9835);
nand U10086 (N_10086,N_9942,N_9979);
nor U10087 (N_10087,N_9951,N_9957);
nor U10088 (N_10088,N_9858,N_9914);
and U10089 (N_10089,N_9879,N_9860);
and U10090 (N_10090,N_9936,N_9833);
and U10091 (N_10091,N_9831,N_9970);
or U10092 (N_10092,N_9998,N_9865);
xor U10093 (N_10093,N_9846,N_9997);
and U10094 (N_10094,N_9924,N_9813);
and U10095 (N_10095,N_9869,N_9873);
xor U10096 (N_10096,N_9891,N_9878);
and U10097 (N_10097,N_9920,N_9947);
and U10098 (N_10098,N_9976,N_9923);
nor U10099 (N_10099,N_9889,N_9996);
nor U10100 (N_10100,N_9971,N_9972);
and U10101 (N_10101,N_9885,N_9959);
and U10102 (N_10102,N_9840,N_9880);
nand U10103 (N_10103,N_9963,N_9980);
nand U10104 (N_10104,N_9854,N_9852);
nor U10105 (N_10105,N_9898,N_9846);
xnor U10106 (N_10106,N_9910,N_9945);
xnor U10107 (N_10107,N_9984,N_9864);
xnor U10108 (N_10108,N_9918,N_9938);
nand U10109 (N_10109,N_9818,N_9837);
nor U10110 (N_10110,N_9903,N_9959);
nand U10111 (N_10111,N_9948,N_9972);
or U10112 (N_10112,N_9846,N_9832);
nand U10113 (N_10113,N_9902,N_9928);
nand U10114 (N_10114,N_9812,N_9926);
or U10115 (N_10115,N_9890,N_9880);
nor U10116 (N_10116,N_9848,N_9990);
xnor U10117 (N_10117,N_9986,N_9921);
xor U10118 (N_10118,N_9914,N_9919);
or U10119 (N_10119,N_9881,N_9913);
and U10120 (N_10120,N_9940,N_9842);
nor U10121 (N_10121,N_9817,N_9888);
and U10122 (N_10122,N_9815,N_9920);
or U10123 (N_10123,N_9822,N_9963);
nor U10124 (N_10124,N_9884,N_9963);
xor U10125 (N_10125,N_9919,N_9987);
and U10126 (N_10126,N_9958,N_9995);
or U10127 (N_10127,N_9855,N_9971);
nor U10128 (N_10128,N_9978,N_9887);
and U10129 (N_10129,N_9854,N_9809);
nor U10130 (N_10130,N_9963,N_9826);
xor U10131 (N_10131,N_9845,N_9884);
and U10132 (N_10132,N_9820,N_9888);
nor U10133 (N_10133,N_9802,N_9921);
xnor U10134 (N_10134,N_9986,N_9997);
or U10135 (N_10135,N_9883,N_9882);
and U10136 (N_10136,N_9826,N_9948);
or U10137 (N_10137,N_9886,N_9841);
or U10138 (N_10138,N_9814,N_9821);
nand U10139 (N_10139,N_9898,N_9989);
nor U10140 (N_10140,N_9802,N_9962);
and U10141 (N_10141,N_9859,N_9898);
xor U10142 (N_10142,N_9921,N_9832);
nand U10143 (N_10143,N_9813,N_9878);
and U10144 (N_10144,N_9881,N_9808);
and U10145 (N_10145,N_9807,N_9916);
and U10146 (N_10146,N_9859,N_9888);
nor U10147 (N_10147,N_9960,N_9956);
nand U10148 (N_10148,N_9857,N_9802);
nor U10149 (N_10149,N_9882,N_9855);
nor U10150 (N_10150,N_9901,N_9854);
and U10151 (N_10151,N_9832,N_9829);
or U10152 (N_10152,N_9805,N_9920);
or U10153 (N_10153,N_9978,N_9973);
or U10154 (N_10154,N_9948,N_9844);
and U10155 (N_10155,N_9847,N_9891);
or U10156 (N_10156,N_9825,N_9929);
and U10157 (N_10157,N_9870,N_9893);
and U10158 (N_10158,N_9934,N_9824);
nor U10159 (N_10159,N_9930,N_9818);
xor U10160 (N_10160,N_9888,N_9913);
and U10161 (N_10161,N_9920,N_9999);
nand U10162 (N_10162,N_9854,N_9985);
or U10163 (N_10163,N_9995,N_9855);
and U10164 (N_10164,N_9878,N_9826);
or U10165 (N_10165,N_9980,N_9934);
xor U10166 (N_10166,N_9909,N_9853);
xnor U10167 (N_10167,N_9802,N_9994);
xnor U10168 (N_10168,N_9909,N_9848);
and U10169 (N_10169,N_9866,N_9938);
nor U10170 (N_10170,N_9879,N_9974);
or U10171 (N_10171,N_9846,N_9964);
or U10172 (N_10172,N_9941,N_9995);
and U10173 (N_10173,N_9887,N_9879);
and U10174 (N_10174,N_9920,N_9829);
xor U10175 (N_10175,N_9943,N_9867);
xor U10176 (N_10176,N_9877,N_9923);
nor U10177 (N_10177,N_9891,N_9848);
nand U10178 (N_10178,N_9963,N_9986);
and U10179 (N_10179,N_9870,N_9912);
nand U10180 (N_10180,N_9880,N_9882);
nand U10181 (N_10181,N_9867,N_9959);
and U10182 (N_10182,N_9829,N_9818);
and U10183 (N_10183,N_9893,N_9895);
nor U10184 (N_10184,N_9828,N_9908);
xnor U10185 (N_10185,N_9851,N_9887);
or U10186 (N_10186,N_9961,N_9928);
or U10187 (N_10187,N_9945,N_9800);
nor U10188 (N_10188,N_9984,N_9884);
nor U10189 (N_10189,N_9863,N_9896);
or U10190 (N_10190,N_9907,N_9957);
nand U10191 (N_10191,N_9849,N_9975);
xnor U10192 (N_10192,N_9819,N_9867);
nor U10193 (N_10193,N_9950,N_9853);
nand U10194 (N_10194,N_9886,N_9910);
or U10195 (N_10195,N_9866,N_9956);
xor U10196 (N_10196,N_9962,N_9975);
and U10197 (N_10197,N_9858,N_9943);
xor U10198 (N_10198,N_9993,N_9982);
nor U10199 (N_10199,N_9939,N_9921);
and U10200 (N_10200,N_10148,N_10146);
or U10201 (N_10201,N_10044,N_10152);
or U10202 (N_10202,N_10119,N_10021);
and U10203 (N_10203,N_10185,N_10117);
and U10204 (N_10204,N_10032,N_10093);
and U10205 (N_10205,N_10058,N_10045);
nand U10206 (N_10206,N_10094,N_10090);
or U10207 (N_10207,N_10017,N_10001);
or U10208 (N_10208,N_10006,N_10123);
nand U10209 (N_10209,N_10091,N_10081);
xor U10210 (N_10210,N_10173,N_10019);
and U10211 (N_10211,N_10193,N_10057);
or U10212 (N_10212,N_10089,N_10102);
nor U10213 (N_10213,N_10160,N_10086);
nor U10214 (N_10214,N_10142,N_10171);
nand U10215 (N_10215,N_10186,N_10197);
or U10216 (N_10216,N_10129,N_10015);
or U10217 (N_10217,N_10043,N_10083);
and U10218 (N_10218,N_10188,N_10155);
and U10219 (N_10219,N_10048,N_10029);
and U10220 (N_10220,N_10149,N_10095);
nand U10221 (N_10221,N_10069,N_10114);
nand U10222 (N_10222,N_10011,N_10087);
or U10223 (N_10223,N_10031,N_10050);
nand U10224 (N_10224,N_10002,N_10139);
nand U10225 (N_10225,N_10157,N_10153);
and U10226 (N_10226,N_10070,N_10012);
xor U10227 (N_10227,N_10159,N_10108);
nand U10228 (N_10228,N_10099,N_10107);
or U10229 (N_10229,N_10135,N_10097);
nand U10230 (N_10230,N_10198,N_10144);
xor U10231 (N_10231,N_10079,N_10130);
xor U10232 (N_10232,N_10164,N_10049);
or U10233 (N_10233,N_10065,N_10098);
and U10234 (N_10234,N_10053,N_10059);
nand U10235 (N_10235,N_10109,N_10167);
nor U10236 (N_10236,N_10163,N_10178);
xnor U10237 (N_10237,N_10132,N_10055);
nand U10238 (N_10238,N_10092,N_10022);
xor U10239 (N_10239,N_10143,N_10066);
nand U10240 (N_10240,N_10072,N_10115);
or U10241 (N_10241,N_10191,N_10003);
or U10242 (N_10242,N_10187,N_10008);
xor U10243 (N_10243,N_10141,N_10116);
nor U10244 (N_10244,N_10088,N_10184);
nand U10245 (N_10245,N_10131,N_10041);
and U10246 (N_10246,N_10038,N_10101);
and U10247 (N_10247,N_10013,N_10016);
or U10248 (N_10248,N_10025,N_10118);
xor U10249 (N_10249,N_10111,N_10181);
or U10250 (N_10250,N_10126,N_10156);
xor U10251 (N_10251,N_10174,N_10120);
and U10252 (N_10252,N_10165,N_10009);
xor U10253 (N_10253,N_10145,N_10176);
nor U10254 (N_10254,N_10140,N_10122);
nor U10255 (N_10255,N_10068,N_10096);
nor U10256 (N_10256,N_10084,N_10138);
nand U10257 (N_10257,N_10196,N_10128);
or U10258 (N_10258,N_10195,N_10158);
nor U10259 (N_10259,N_10104,N_10051);
xnor U10260 (N_10260,N_10054,N_10082);
and U10261 (N_10261,N_10047,N_10035);
or U10262 (N_10262,N_10067,N_10113);
or U10263 (N_10263,N_10162,N_10037);
nand U10264 (N_10264,N_10034,N_10033);
nor U10265 (N_10265,N_10103,N_10080);
nand U10266 (N_10266,N_10075,N_10180);
or U10267 (N_10267,N_10136,N_10040);
xnor U10268 (N_10268,N_10150,N_10077);
nor U10269 (N_10269,N_10039,N_10170);
nand U10270 (N_10270,N_10060,N_10175);
xor U10271 (N_10271,N_10154,N_10190);
or U10272 (N_10272,N_10023,N_10183);
nor U10273 (N_10273,N_10161,N_10036);
and U10274 (N_10274,N_10172,N_10074);
nor U10275 (N_10275,N_10056,N_10134);
nor U10276 (N_10276,N_10133,N_10100);
nand U10277 (N_10277,N_10169,N_10042);
nand U10278 (N_10278,N_10137,N_10199);
xor U10279 (N_10279,N_10147,N_10078);
nand U10280 (N_10280,N_10192,N_10177);
nor U10281 (N_10281,N_10020,N_10125);
nor U10282 (N_10282,N_10046,N_10194);
and U10283 (N_10283,N_10018,N_10182);
and U10284 (N_10284,N_10179,N_10024);
nand U10285 (N_10285,N_10007,N_10105);
xor U10286 (N_10286,N_10028,N_10064);
xor U10287 (N_10287,N_10005,N_10076);
and U10288 (N_10288,N_10014,N_10052);
and U10289 (N_10289,N_10189,N_10071);
or U10290 (N_10290,N_10112,N_10026);
nor U10291 (N_10291,N_10010,N_10061);
nand U10292 (N_10292,N_10106,N_10166);
xor U10293 (N_10293,N_10124,N_10063);
and U10294 (N_10294,N_10030,N_10073);
xnor U10295 (N_10295,N_10085,N_10168);
nand U10296 (N_10296,N_10000,N_10004);
and U10297 (N_10297,N_10110,N_10121);
or U10298 (N_10298,N_10062,N_10027);
xor U10299 (N_10299,N_10151,N_10127);
or U10300 (N_10300,N_10032,N_10173);
nor U10301 (N_10301,N_10111,N_10083);
nor U10302 (N_10302,N_10139,N_10167);
xor U10303 (N_10303,N_10048,N_10189);
nor U10304 (N_10304,N_10009,N_10001);
xnor U10305 (N_10305,N_10055,N_10051);
or U10306 (N_10306,N_10004,N_10063);
xnor U10307 (N_10307,N_10042,N_10087);
nand U10308 (N_10308,N_10146,N_10154);
nor U10309 (N_10309,N_10108,N_10186);
xor U10310 (N_10310,N_10125,N_10084);
or U10311 (N_10311,N_10055,N_10084);
or U10312 (N_10312,N_10000,N_10171);
and U10313 (N_10313,N_10021,N_10027);
and U10314 (N_10314,N_10043,N_10024);
nand U10315 (N_10315,N_10161,N_10042);
or U10316 (N_10316,N_10180,N_10126);
nand U10317 (N_10317,N_10086,N_10151);
or U10318 (N_10318,N_10103,N_10104);
nor U10319 (N_10319,N_10111,N_10023);
or U10320 (N_10320,N_10116,N_10187);
xnor U10321 (N_10321,N_10173,N_10104);
or U10322 (N_10322,N_10124,N_10045);
nand U10323 (N_10323,N_10137,N_10061);
nor U10324 (N_10324,N_10177,N_10038);
nor U10325 (N_10325,N_10004,N_10025);
xor U10326 (N_10326,N_10158,N_10180);
and U10327 (N_10327,N_10166,N_10109);
xnor U10328 (N_10328,N_10161,N_10106);
and U10329 (N_10329,N_10030,N_10063);
nor U10330 (N_10330,N_10107,N_10105);
xor U10331 (N_10331,N_10038,N_10168);
and U10332 (N_10332,N_10158,N_10153);
xor U10333 (N_10333,N_10166,N_10090);
or U10334 (N_10334,N_10032,N_10127);
nand U10335 (N_10335,N_10113,N_10068);
or U10336 (N_10336,N_10013,N_10073);
and U10337 (N_10337,N_10027,N_10061);
or U10338 (N_10338,N_10011,N_10154);
nand U10339 (N_10339,N_10050,N_10108);
nor U10340 (N_10340,N_10166,N_10182);
nand U10341 (N_10341,N_10075,N_10190);
and U10342 (N_10342,N_10078,N_10154);
xnor U10343 (N_10343,N_10026,N_10193);
nand U10344 (N_10344,N_10190,N_10170);
nor U10345 (N_10345,N_10169,N_10065);
nand U10346 (N_10346,N_10078,N_10059);
nand U10347 (N_10347,N_10117,N_10079);
nand U10348 (N_10348,N_10029,N_10198);
or U10349 (N_10349,N_10067,N_10115);
and U10350 (N_10350,N_10007,N_10070);
nor U10351 (N_10351,N_10167,N_10009);
and U10352 (N_10352,N_10110,N_10011);
xnor U10353 (N_10353,N_10181,N_10026);
nand U10354 (N_10354,N_10176,N_10162);
or U10355 (N_10355,N_10175,N_10024);
nand U10356 (N_10356,N_10062,N_10146);
nor U10357 (N_10357,N_10151,N_10101);
and U10358 (N_10358,N_10022,N_10037);
nor U10359 (N_10359,N_10094,N_10178);
or U10360 (N_10360,N_10155,N_10112);
xor U10361 (N_10361,N_10089,N_10084);
and U10362 (N_10362,N_10116,N_10179);
nor U10363 (N_10363,N_10033,N_10069);
or U10364 (N_10364,N_10051,N_10190);
xor U10365 (N_10365,N_10078,N_10063);
xor U10366 (N_10366,N_10190,N_10123);
nand U10367 (N_10367,N_10058,N_10155);
or U10368 (N_10368,N_10158,N_10166);
xnor U10369 (N_10369,N_10115,N_10175);
nor U10370 (N_10370,N_10138,N_10009);
nor U10371 (N_10371,N_10122,N_10068);
and U10372 (N_10372,N_10138,N_10143);
nand U10373 (N_10373,N_10000,N_10135);
nor U10374 (N_10374,N_10066,N_10003);
or U10375 (N_10375,N_10066,N_10081);
or U10376 (N_10376,N_10002,N_10044);
and U10377 (N_10377,N_10034,N_10004);
and U10378 (N_10378,N_10191,N_10043);
or U10379 (N_10379,N_10015,N_10189);
xor U10380 (N_10380,N_10055,N_10048);
xnor U10381 (N_10381,N_10127,N_10136);
xor U10382 (N_10382,N_10090,N_10109);
or U10383 (N_10383,N_10051,N_10006);
nor U10384 (N_10384,N_10143,N_10067);
xor U10385 (N_10385,N_10105,N_10137);
nand U10386 (N_10386,N_10073,N_10152);
xnor U10387 (N_10387,N_10089,N_10132);
xnor U10388 (N_10388,N_10155,N_10192);
and U10389 (N_10389,N_10177,N_10150);
xor U10390 (N_10390,N_10138,N_10073);
or U10391 (N_10391,N_10010,N_10116);
nand U10392 (N_10392,N_10023,N_10070);
or U10393 (N_10393,N_10173,N_10035);
nand U10394 (N_10394,N_10173,N_10195);
and U10395 (N_10395,N_10152,N_10097);
nor U10396 (N_10396,N_10027,N_10145);
and U10397 (N_10397,N_10088,N_10083);
nand U10398 (N_10398,N_10177,N_10106);
or U10399 (N_10399,N_10025,N_10146);
nor U10400 (N_10400,N_10236,N_10388);
or U10401 (N_10401,N_10283,N_10262);
xor U10402 (N_10402,N_10218,N_10281);
and U10403 (N_10403,N_10264,N_10325);
nor U10404 (N_10404,N_10329,N_10304);
xor U10405 (N_10405,N_10291,N_10373);
nor U10406 (N_10406,N_10247,N_10275);
xnor U10407 (N_10407,N_10386,N_10313);
and U10408 (N_10408,N_10284,N_10278);
or U10409 (N_10409,N_10277,N_10255);
and U10410 (N_10410,N_10316,N_10273);
nor U10411 (N_10411,N_10308,N_10225);
xnor U10412 (N_10412,N_10384,N_10245);
xor U10413 (N_10413,N_10372,N_10323);
xnor U10414 (N_10414,N_10259,N_10357);
and U10415 (N_10415,N_10363,N_10379);
nand U10416 (N_10416,N_10294,N_10345);
or U10417 (N_10417,N_10209,N_10341);
and U10418 (N_10418,N_10370,N_10267);
nor U10419 (N_10419,N_10269,N_10237);
xor U10420 (N_10420,N_10383,N_10358);
nand U10421 (N_10421,N_10274,N_10367);
nand U10422 (N_10422,N_10314,N_10227);
nor U10423 (N_10423,N_10265,N_10380);
nor U10424 (N_10424,N_10261,N_10207);
or U10425 (N_10425,N_10289,N_10331);
nand U10426 (N_10426,N_10397,N_10365);
nand U10427 (N_10427,N_10217,N_10344);
and U10428 (N_10428,N_10266,N_10303);
xnor U10429 (N_10429,N_10223,N_10296);
nand U10430 (N_10430,N_10307,N_10254);
and U10431 (N_10431,N_10276,N_10216);
nand U10432 (N_10432,N_10221,N_10208);
or U10433 (N_10433,N_10375,N_10203);
nor U10434 (N_10434,N_10298,N_10324);
nand U10435 (N_10435,N_10250,N_10224);
or U10436 (N_10436,N_10239,N_10387);
and U10437 (N_10437,N_10231,N_10299);
nand U10438 (N_10438,N_10311,N_10263);
xor U10439 (N_10439,N_10390,N_10200);
nor U10440 (N_10440,N_10315,N_10286);
nor U10441 (N_10441,N_10288,N_10394);
and U10442 (N_10442,N_10335,N_10346);
xnor U10443 (N_10443,N_10252,N_10310);
nand U10444 (N_10444,N_10292,N_10336);
nor U10445 (N_10445,N_10321,N_10234);
and U10446 (N_10446,N_10347,N_10360);
xor U10447 (N_10447,N_10282,N_10333);
xor U10448 (N_10448,N_10251,N_10319);
and U10449 (N_10449,N_10215,N_10359);
xor U10450 (N_10450,N_10272,N_10369);
or U10451 (N_10451,N_10328,N_10280);
nor U10452 (N_10452,N_10240,N_10248);
xor U10453 (N_10453,N_10212,N_10257);
xor U10454 (N_10454,N_10312,N_10391);
xnor U10455 (N_10455,N_10342,N_10256);
nand U10456 (N_10456,N_10242,N_10230);
nor U10457 (N_10457,N_10356,N_10253);
nand U10458 (N_10458,N_10349,N_10305);
or U10459 (N_10459,N_10233,N_10340);
and U10460 (N_10460,N_10332,N_10211);
nor U10461 (N_10461,N_10213,N_10300);
and U10462 (N_10462,N_10297,N_10279);
nand U10463 (N_10463,N_10355,N_10326);
and U10464 (N_10464,N_10205,N_10399);
and U10465 (N_10465,N_10318,N_10398);
nand U10466 (N_10466,N_10210,N_10320);
and U10467 (N_10467,N_10374,N_10334);
nand U10468 (N_10468,N_10389,N_10220);
xnor U10469 (N_10469,N_10382,N_10222);
or U10470 (N_10470,N_10235,N_10371);
xnor U10471 (N_10471,N_10317,N_10271);
or U10472 (N_10472,N_10244,N_10241);
and U10473 (N_10473,N_10396,N_10229);
nor U10474 (N_10474,N_10302,N_10362);
or U10475 (N_10475,N_10260,N_10226);
or U10476 (N_10476,N_10381,N_10364);
nor U10477 (N_10477,N_10366,N_10219);
nand U10478 (N_10478,N_10368,N_10202);
nor U10479 (N_10479,N_10393,N_10339);
xor U10480 (N_10480,N_10301,N_10353);
xor U10481 (N_10481,N_10258,N_10204);
xnor U10482 (N_10482,N_10232,N_10361);
nand U10483 (N_10483,N_10376,N_10354);
nor U10484 (N_10484,N_10228,N_10270);
or U10485 (N_10485,N_10293,N_10322);
nand U10486 (N_10486,N_10343,N_10348);
nor U10487 (N_10487,N_10238,N_10352);
xnor U10488 (N_10488,N_10285,N_10268);
or U10489 (N_10489,N_10350,N_10330);
or U10490 (N_10490,N_10214,N_10246);
or U10491 (N_10491,N_10327,N_10306);
nand U10492 (N_10492,N_10338,N_10337);
xor U10493 (N_10493,N_10206,N_10287);
and U10494 (N_10494,N_10392,N_10377);
nand U10495 (N_10495,N_10395,N_10290);
xor U10496 (N_10496,N_10385,N_10249);
nand U10497 (N_10497,N_10201,N_10295);
nor U10498 (N_10498,N_10378,N_10309);
and U10499 (N_10499,N_10351,N_10243);
nand U10500 (N_10500,N_10212,N_10351);
and U10501 (N_10501,N_10344,N_10272);
or U10502 (N_10502,N_10307,N_10242);
or U10503 (N_10503,N_10263,N_10315);
xor U10504 (N_10504,N_10340,N_10388);
and U10505 (N_10505,N_10319,N_10258);
nor U10506 (N_10506,N_10390,N_10283);
and U10507 (N_10507,N_10292,N_10332);
and U10508 (N_10508,N_10308,N_10213);
nand U10509 (N_10509,N_10350,N_10261);
and U10510 (N_10510,N_10323,N_10268);
nor U10511 (N_10511,N_10384,N_10293);
xor U10512 (N_10512,N_10281,N_10361);
xnor U10513 (N_10513,N_10341,N_10225);
nor U10514 (N_10514,N_10215,N_10268);
xnor U10515 (N_10515,N_10287,N_10370);
xnor U10516 (N_10516,N_10266,N_10224);
nand U10517 (N_10517,N_10361,N_10328);
xor U10518 (N_10518,N_10238,N_10219);
nor U10519 (N_10519,N_10280,N_10321);
or U10520 (N_10520,N_10269,N_10336);
or U10521 (N_10521,N_10384,N_10287);
nor U10522 (N_10522,N_10231,N_10243);
nand U10523 (N_10523,N_10398,N_10395);
or U10524 (N_10524,N_10250,N_10303);
nand U10525 (N_10525,N_10386,N_10392);
xor U10526 (N_10526,N_10377,N_10282);
or U10527 (N_10527,N_10228,N_10359);
nor U10528 (N_10528,N_10252,N_10373);
or U10529 (N_10529,N_10212,N_10325);
and U10530 (N_10530,N_10375,N_10200);
nor U10531 (N_10531,N_10315,N_10363);
nand U10532 (N_10532,N_10269,N_10266);
and U10533 (N_10533,N_10237,N_10334);
and U10534 (N_10534,N_10371,N_10290);
nand U10535 (N_10535,N_10246,N_10320);
nor U10536 (N_10536,N_10224,N_10310);
xnor U10537 (N_10537,N_10268,N_10328);
or U10538 (N_10538,N_10219,N_10310);
or U10539 (N_10539,N_10370,N_10315);
xor U10540 (N_10540,N_10206,N_10365);
xnor U10541 (N_10541,N_10232,N_10216);
nor U10542 (N_10542,N_10332,N_10239);
and U10543 (N_10543,N_10257,N_10268);
and U10544 (N_10544,N_10314,N_10210);
nor U10545 (N_10545,N_10320,N_10357);
and U10546 (N_10546,N_10238,N_10215);
or U10547 (N_10547,N_10279,N_10289);
or U10548 (N_10548,N_10291,N_10278);
nand U10549 (N_10549,N_10309,N_10204);
nand U10550 (N_10550,N_10356,N_10261);
and U10551 (N_10551,N_10357,N_10299);
or U10552 (N_10552,N_10294,N_10315);
or U10553 (N_10553,N_10370,N_10385);
or U10554 (N_10554,N_10263,N_10314);
or U10555 (N_10555,N_10230,N_10277);
nor U10556 (N_10556,N_10289,N_10262);
xor U10557 (N_10557,N_10231,N_10314);
nand U10558 (N_10558,N_10253,N_10327);
xnor U10559 (N_10559,N_10360,N_10303);
xnor U10560 (N_10560,N_10344,N_10323);
or U10561 (N_10561,N_10229,N_10246);
nor U10562 (N_10562,N_10385,N_10272);
nand U10563 (N_10563,N_10390,N_10208);
or U10564 (N_10564,N_10389,N_10236);
and U10565 (N_10565,N_10365,N_10348);
nand U10566 (N_10566,N_10357,N_10344);
nand U10567 (N_10567,N_10266,N_10380);
nor U10568 (N_10568,N_10243,N_10251);
or U10569 (N_10569,N_10368,N_10287);
nand U10570 (N_10570,N_10332,N_10313);
and U10571 (N_10571,N_10314,N_10214);
and U10572 (N_10572,N_10300,N_10349);
or U10573 (N_10573,N_10345,N_10348);
and U10574 (N_10574,N_10227,N_10385);
and U10575 (N_10575,N_10352,N_10310);
and U10576 (N_10576,N_10307,N_10374);
or U10577 (N_10577,N_10201,N_10219);
or U10578 (N_10578,N_10341,N_10230);
and U10579 (N_10579,N_10358,N_10397);
nor U10580 (N_10580,N_10237,N_10207);
nor U10581 (N_10581,N_10277,N_10273);
nor U10582 (N_10582,N_10241,N_10257);
xnor U10583 (N_10583,N_10245,N_10224);
nand U10584 (N_10584,N_10258,N_10369);
or U10585 (N_10585,N_10245,N_10297);
nand U10586 (N_10586,N_10248,N_10396);
xor U10587 (N_10587,N_10298,N_10334);
and U10588 (N_10588,N_10278,N_10295);
nand U10589 (N_10589,N_10236,N_10359);
or U10590 (N_10590,N_10349,N_10357);
nor U10591 (N_10591,N_10325,N_10333);
and U10592 (N_10592,N_10313,N_10252);
xnor U10593 (N_10593,N_10363,N_10290);
and U10594 (N_10594,N_10390,N_10296);
nor U10595 (N_10595,N_10350,N_10226);
nor U10596 (N_10596,N_10224,N_10359);
and U10597 (N_10597,N_10328,N_10318);
nand U10598 (N_10598,N_10339,N_10303);
or U10599 (N_10599,N_10216,N_10236);
nand U10600 (N_10600,N_10470,N_10401);
nand U10601 (N_10601,N_10554,N_10512);
or U10602 (N_10602,N_10580,N_10471);
and U10603 (N_10603,N_10566,N_10567);
or U10604 (N_10604,N_10559,N_10496);
xnor U10605 (N_10605,N_10436,N_10492);
nor U10606 (N_10606,N_10596,N_10411);
and U10607 (N_10607,N_10502,N_10485);
or U10608 (N_10608,N_10523,N_10557);
and U10609 (N_10609,N_10572,N_10460);
nand U10610 (N_10610,N_10534,N_10467);
and U10611 (N_10611,N_10585,N_10521);
and U10612 (N_10612,N_10586,N_10597);
and U10613 (N_10613,N_10561,N_10420);
nand U10614 (N_10614,N_10447,N_10574);
nand U10615 (N_10615,N_10484,N_10402);
nor U10616 (N_10616,N_10590,N_10422);
and U10617 (N_10617,N_10466,N_10419);
nor U10618 (N_10618,N_10594,N_10493);
xnor U10619 (N_10619,N_10469,N_10475);
nand U10620 (N_10620,N_10591,N_10431);
nor U10621 (N_10621,N_10463,N_10457);
xnor U10622 (N_10622,N_10491,N_10576);
nor U10623 (N_10623,N_10589,N_10588);
nand U10624 (N_10624,N_10548,N_10499);
or U10625 (N_10625,N_10480,N_10515);
nand U10626 (N_10626,N_10509,N_10456);
and U10627 (N_10627,N_10505,N_10525);
and U10628 (N_10628,N_10595,N_10528);
nand U10629 (N_10629,N_10508,N_10448);
or U10630 (N_10630,N_10568,N_10433);
or U10631 (N_10631,N_10516,N_10524);
nand U10632 (N_10632,N_10430,N_10405);
and U10633 (N_10633,N_10479,N_10550);
nand U10634 (N_10634,N_10562,N_10497);
and U10635 (N_10635,N_10472,N_10584);
nor U10636 (N_10636,N_10409,N_10582);
xnor U10637 (N_10637,N_10407,N_10477);
nand U10638 (N_10638,N_10426,N_10579);
nor U10639 (N_10639,N_10565,N_10536);
and U10640 (N_10640,N_10545,N_10526);
and U10641 (N_10641,N_10531,N_10518);
or U10642 (N_10642,N_10424,N_10533);
nor U10643 (N_10643,N_10483,N_10450);
and U10644 (N_10644,N_10446,N_10489);
and U10645 (N_10645,N_10519,N_10546);
nand U10646 (N_10646,N_10558,N_10439);
nor U10647 (N_10647,N_10541,N_10547);
and U10648 (N_10648,N_10520,N_10569);
xnor U10649 (N_10649,N_10474,N_10503);
and U10650 (N_10650,N_10454,N_10410);
nand U10651 (N_10651,N_10458,N_10560);
nand U10652 (N_10652,N_10425,N_10434);
nor U10653 (N_10653,N_10486,N_10412);
nand U10654 (N_10654,N_10476,N_10532);
nand U10655 (N_10655,N_10473,N_10564);
or U10656 (N_10656,N_10495,N_10598);
xnor U10657 (N_10657,N_10538,N_10452);
nand U10658 (N_10658,N_10513,N_10573);
xnor U10659 (N_10659,N_10592,N_10432);
xor U10660 (N_10660,N_10529,N_10465);
nor U10661 (N_10661,N_10552,N_10498);
nor U10662 (N_10662,N_10404,N_10488);
nor U10663 (N_10663,N_10549,N_10514);
xnor U10664 (N_10664,N_10577,N_10535);
nor U10665 (N_10665,N_10442,N_10464);
nor U10666 (N_10666,N_10500,N_10429);
and U10667 (N_10667,N_10435,N_10408);
xor U10668 (N_10668,N_10438,N_10428);
or U10669 (N_10669,N_10555,N_10414);
xor U10670 (N_10670,N_10423,N_10571);
xor U10671 (N_10671,N_10462,N_10482);
nand U10672 (N_10672,N_10583,N_10453);
and U10673 (N_10673,N_10530,N_10490);
and U10674 (N_10674,N_10504,N_10406);
nor U10675 (N_10675,N_10413,N_10444);
and U10676 (N_10676,N_10421,N_10587);
or U10677 (N_10677,N_10468,N_10522);
xnor U10678 (N_10678,N_10581,N_10501);
or U10679 (N_10679,N_10517,N_10494);
and U10680 (N_10680,N_10563,N_10461);
nand U10681 (N_10681,N_10455,N_10539);
nor U10682 (N_10682,N_10556,N_10506);
and U10683 (N_10683,N_10544,N_10570);
xor U10684 (N_10684,N_10478,N_10449);
nor U10685 (N_10685,N_10481,N_10511);
or U10686 (N_10686,N_10400,N_10540);
xnor U10687 (N_10687,N_10510,N_10527);
nor U10688 (N_10688,N_10443,N_10451);
and U10689 (N_10689,N_10578,N_10440);
and U10690 (N_10690,N_10441,N_10593);
and U10691 (N_10691,N_10543,N_10459);
or U10692 (N_10692,N_10417,N_10415);
nand U10693 (N_10693,N_10599,N_10418);
nor U10694 (N_10694,N_10553,N_10487);
nand U10695 (N_10695,N_10416,N_10427);
nor U10696 (N_10696,N_10542,N_10507);
xor U10697 (N_10697,N_10403,N_10537);
nand U10698 (N_10698,N_10575,N_10437);
xor U10699 (N_10699,N_10445,N_10551);
or U10700 (N_10700,N_10429,N_10444);
xnor U10701 (N_10701,N_10493,N_10464);
nor U10702 (N_10702,N_10589,N_10488);
nor U10703 (N_10703,N_10533,N_10509);
nand U10704 (N_10704,N_10545,N_10410);
nand U10705 (N_10705,N_10500,N_10597);
and U10706 (N_10706,N_10568,N_10402);
nor U10707 (N_10707,N_10542,N_10413);
and U10708 (N_10708,N_10444,N_10405);
nand U10709 (N_10709,N_10562,N_10459);
or U10710 (N_10710,N_10564,N_10511);
or U10711 (N_10711,N_10468,N_10525);
or U10712 (N_10712,N_10475,N_10437);
xnor U10713 (N_10713,N_10523,N_10586);
and U10714 (N_10714,N_10479,N_10530);
and U10715 (N_10715,N_10451,N_10579);
nor U10716 (N_10716,N_10417,N_10487);
or U10717 (N_10717,N_10450,N_10464);
nand U10718 (N_10718,N_10405,N_10532);
xor U10719 (N_10719,N_10425,N_10546);
or U10720 (N_10720,N_10574,N_10439);
and U10721 (N_10721,N_10469,N_10520);
or U10722 (N_10722,N_10496,N_10595);
xor U10723 (N_10723,N_10578,N_10593);
nor U10724 (N_10724,N_10415,N_10453);
and U10725 (N_10725,N_10543,N_10529);
nor U10726 (N_10726,N_10485,N_10552);
nand U10727 (N_10727,N_10404,N_10461);
nor U10728 (N_10728,N_10522,N_10561);
and U10729 (N_10729,N_10451,N_10472);
nand U10730 (N_10730,N_10465,N_10598);
or U10731 (N_10731,N_10432,N_10502);
xor U10732 (N_10732,N_10545,N_10491);
nand U10733 (N_10733,N_10540,N_10554);
or U10734 (N_10734,N_10464,N_10514);
nand U10735 (N_10735,N_10454,N_10407);
nor U10736 (N_10736,N_10488,N_10557);
xnor U10737 (N_10737,N_10570,N_10574);
xnor U10738 (N_10738,N_10461,N_10440);
xor U10739 (N_10739,N_10473,N_10527);
nand U10740 (N_10740,N_10543,N_10436);
nor U10741 (N_10741,N_10467,N_10413);
nand U10742 (N_10742,N_10478,N_10477);
and U10743 (N_10743,N_10559,N_10422);
and U10744 (N_10744,N_10453,N_10465);
xnor U10745 (N_10745,N_10568,N_10422);
nor U10746 (N_10746,N_10534,N_10463);
or U10747 (N_10747,N_10438,N_10585);
nand U10748 (N_10748,N_10424,N_10566);
and U10749 (N_10749,N_10467,N_10515);
or U10750 (N_10750,N_10421,N_10477);
and U10751 (N_10751,N_10596,N_10584);
xnor U10752 (N_10752,N_10560,N_10433);
nand U10753 (N_10753,N_10475,N_10480);
nor U10754 (N_10754,N_10524,N_10459);
nand U10755 (N_10755,N_10405,N_10517);
xor U10756 (N_10756,N_10442,N_10519);
or U10757 (N_10757,N_10590,N_10440);
or U10758 (N_10758,N_10520,N_10568);
or U10759 (N_10759,N_10424,N_10461);
nor U10760 (N_10760,N_10530,N_10410);
or U10761 (N_10761,N_10489,N_10539);
nor U10762 (N_10762,N_10578,N_10561);
xnor U10763 (N_10763,N_10409,N_10515);
nand U10764 (N_10764,N_10492,N_10487);
xnor U10765 (N_10765,N_10580,N_10485);
nor U10766 (N_10766,N_10544,N_10400);
xor U10767 (N_10767,N_10498,N_10411);
xor U10768 (N_10768,N_10526,N_10575);
xor U10769 (N_10769,N_10416,N_10469);
xor U10770 (N_10770,N_10531,N_10459);
xor U10771 (N_10771,N_10426,N_10572);
xor U10772 (N_10772,N_10429,N_10595);
xnor U10773 (N_10773,N_10531,N_10461);
nand U10774 (N_10774,N_10514,N_10558);
and U10775 (N_10775,N_10575,N_10554);
xor U10776 (N_10776,N_10419,N_10552);
nor U10777 (N_10777,N_10535,N_10485);
nand U10778 (N_10778,N_10587,N_10429);
and U10779 (N_10779,N_10541,N_10489);
nand U10780 (N_10780,N_10539,N_10591);
xor U10781 (N_10781,N_10541,N_10538);
or U10782 (N_10782,N_10432,N_10550);
or U10783 (N_10783,N_10485,N_10413);
and U10784 (N_10784,N_10591,N_10433);
and U10785 (N_10785,N_10578,N_10403);
xnor U10786 (N_10786,N_10556,N_10403);
or U10787 (N_10787,N_10531,N_10529);
and U10788 (N_10788,N_10536,N_10527);
nor U10789 (N_10789,N_10509,N_10500);
nand U10790 (N_10790,N_10430,N_10452);
or U10791 (N_10791,N_10497,N_10450);
xor U10792 (N_10792,N_10422,N_10563);
xnor U10793 (N_10793,N_10544,N_10403);
nand U10794 (N_10794,N_10556,N_10543);
xnor U10795 (N_10795,N_10413,N_10436);
nand U10796 (N_10796,N_10477,N_10506);
and U10797 (N_10797,N_10431,N_10401);
or U10798 (N_10798,N_10416,N_10596);
and U10799 (N_10799,N_10438,N_10422);
and U10800 (N_10800,N_10722,N_10603);
and U10801 (N_10801,N_10763,N_10700);
nor U10802 (N_10802,N_10629,N_10671);
or U10803 (N_10803,N_10652,N_10684);
and U10804 (N_10804,N_10719,N_10689);
or U10805 (N_10805,N_10678,N_10787);
nand U10806 (N_10806,N_10724,N_10609);
xor U10807 (N_10807,N_10674,N_10693);
or U10808 (N_10808,N_10707,N_10645);
xnor U10809 (N_10809,N_10610,N_10696);
or U10810 (N_10810,N_10628,N_10737);
nor U10811 (N_10811,N_10682,N_10602);
or U10812 (N_10812,N_10607,N_10711);
xnor U10813 (N_10813,N_10751,N_10714);
nand U10814 (N_10814,N_10611,N_10782);
xor U10815 (N_10815,N_10762,N_10744);
xor U10816 (N_10816,N_10663,N_10771);
or U10817 (N_10817,N_10661,N_10765);
nand U10818 (N_10818,N_10735,N_10646);
and U10819 (N_10819,N_10699,N_10760);
nor U10820 (N_10820,N_10638,N_10709);
xor U10821 (N_10821,N_10620,N_10656);
and U10822 (N_10822,N_10701,N_10746);
and U10823 (N_10823,N_10758,N_10604);
and U10824 (N_10824,N_10742,N_10727);
or U10825 (N_10825,N_10740,N_10739);
nand U10826 (N_10826,N_10770,N_10605);
nand U10827 (N_10827,N_10778,N_10692);
nor U10828 (N_10828,N_10676,N_10748);
or U10829 (N_10829,N_10710,N_10725);
xor U10830 (N_10830,N_10755,N_10649);
nor U10831 (N_10831,N_10720,N_10768);
and U10832 (N_10832,N_10776,N_10639);
nand U10833 (N_10833,N_10614,N_10792);
nand U10834 (N_10834,N_10713,N_10706);
or U10835 (N_10835,N_10750,N_10736);
nor U10836 (N_10836,N_10774,N_10679);
or U10837 (N_10837,N_10631,N_10759);
and U10838 (N_10838,N_10741,N_10647);
and U10839 (N_10839,N_10769,N_10749);
and U10840 (N_10840,N_10657,N_10718);
or U10841 (N_10841,N_10613,N_10636);
and U10842 (N_10842,N_10665,N_10777);
and U10843 (N_10843,N_10716,N_10723);
nand U10844 (N_10844,N_10756,N_10772);
nand U10845 (N_10845,N_10686,N_10643);
nor U10846 (N_10846,N_10673,N_10797);
xnor U10847 (N_10847,N_10670,N_10781);
and U10848 (N_10848,N_10695,N_10767);
nor U10849 (N_10849,N_10773,N_10654);
and U10850 (N_10850,N_10627,N_10785);
or U10851 (N_10851,N_10738,N_10675);
nand U10852 (N_10852,N_10618,N_10705);
or U10853 (N_10853,N_10612,N_10795);
xnor U10854 (N_10854,N_10685,N_10616);
or U10855 (N_10855,N_10664,N_10621);
and U10856 (N_10856,N_10789,N_10623);
and U10857 (N_10857,N_10615,N_10653);
nor U10858 (N_10858,N_10690,N_10786);
or U10859 (N_10859,N_10667,N_10731);
xnor U10860 (N_10860,N_10668,N_10747);
nand U10861 (N_10861,N_10681,N_10677);
xor U10862 (N_10862,N_10753,N_10788);
nand U10863 (N_10863,N_10680,N_10633);
or U10864 (N_10864,N_10761,N_10625);
and U10865 (N_10865,N_10703,N_10644);
xor U10866 (N_10866,N_10712,N_10779);
nor U10867 (N_10867,N_10624,N_10691);
or U10868 (N_10868,N_10622,N_10650);
nand U10869 (N_10869,N_10728,N_10617);
xor U10870 (N_10870,N_10632,N_10635);
xor U10871 (N_10871,N_10702,N_10626);
xnor U10872 (N_10872,N_10642,N_10743);
nand U10873 (N_10873,N_10648,N_10662);
nand U10874 (N_10874,N_10775,N_10660);
nor U10875 (N_10875,N_10688,N_10784);
nand U10876 (N_10876,N_10694,N_10697);
or U10877 (N_10877,N_10793,N_10732);
and U10878 (N_10878,N_10754,N_10658);
xor U10879 (N_10879,N_10726,N_10794);
nand U10880 (N_10880,N_10637,N_10619);
nand U10881 (N_10881,N_10730,N_10606);
nor U10882 (N_10882,N_10683,N_10634);
nor U10883 (N_10883,N_10752,N_10640);
nand U10884 (N_10884,N_10698,N_10757);
nor U10885 (N_10885,N_10601,N_10608);
nor U10886 (N_10886,N_10745,N_10790);
and U10887 (N_10887,N_10687,N_10659);
nor U10888 (N_10888,N_10780,N_10799);
and U10889 (N_10889,N_10669,N_10783);
nand U10890 (N_10890,N_10766,N_10717);
and U10891 (N_10891,N_10721,N_10666);
nand U10892 (N_10892,N_10798,N_10672);
nor U10893 (N_10893,N_10641,N_10630);
or U10894 (N_10894,N_10791,N_10708);
or U10895 (N_10895,N_10796,N_10733);
nor U10896 (N_10896,N_10734,N_10729);
or U10897 (N_10897,N_10600,N_10704);
and U10898 (N_10898,N_10651,N_10715);
or U10899 (N_10899,N_10764,N_10655);
xnor U10900 (N_10900,N_10690,N_10799);
nand U10901 (N_10901,N_10699,N_10733);
xor U10902 (N_10902,N_10741,N_10663);
nand U10903 (N_10903,N_10776,N_10708);
or U10904 (N_10904,N_10646,N_10755);
xor U10905 (N_10905,N_10654,N_10640);
nand U10906 (N_10906,N_10735,N_10759);
and U10907 (N_10907,N_10642,N_10779);
nor U10908 (N_10908,N_10619,N_10731);
and U10909 (N_10909,N_10647,N_10761);
or U10910 (N_10910,N_10734,N_10693);
or U10911 (N_10911,N_10635,N_10627);
or U10912 (N_10912,N_10660,N_10786);
xnor U10913 (N_10913,N_10637,N_10770);
or U10914 (N_10914,N_10627,N_10753);
nand U10915 (N_10915,N_10694,N_10791);
nor U10916 (N_10916,N_10659,N_10752);
nor U10917 (N_10917,N_10731,N_10610);
or U10918 (N_10918,N_10675,N_10618);
and U10919 (N_10919,N_10610,N_10737);
xor U10920 (N_10920,N_10606,N_10781);
xor U10921 (N_10921,N_10794,N_10757);
or U10922 (N_10922,N_10648,N_10716);
xor U10923 (N_10923,N_10695,N_10746);
nand U10924 (N_10924,N_10793,N_10718);
nor U10925 (N_10925,N_10643,N_10721);
and U10926 (N_10926,N_10692,N_10631);
and U10927 (N_10927,N_10620,N_10789);
or U10928 (N_10928,N_10744,N_10678);
and U10929 (N_10929,N_10693,N_10680);
nand U10930 (N_10930,N_10787,N_10726);
nor U10931 (N_10931,N_10605,N_10746);
and U10932 (N_10932,N_10649,N_10635);
or U10933 (N_10933,N_10644,N_10712);
and U10934 (N_10934,N_10663,N_10747);
nor U10935 (N_10935,N_10693,N_10710);
or U10936 (N_10936,N_10744,N_10671);
nor U10937 (N_10937,N_10614,N_10632);
nand U10938 (N_10938,N_10636,N_10660);
nor U10939 (N_10939,N_10615,N_10759);
and U10940 (N_10940,N_10767,N_10749);
nand U10941 (N_10941,N_10646,N_10602);
nand U10942 (N_10942,N_10733,N_10743);
xnor U10943 (N_10943,N_10675,N_10794);
and U10944 (N_10944,N_10660,N_10622);
nor U10945 (N_10945,N_10758,N_10649);
and U10946 (N_10946,N_10717,N_10659);
and U10947 (N_10947,N_10715,N_10686);
xnor U10948 (N_10948,N_10719,N_10755);
or U10949 (N_10949,N_10659,N_10608);
or U10950 (N_10950,N_10755,N_10691);
nand U10951 (N_10951,N_10687,N_10601);
xnor U10952 (N_10952,N_10755,N_10791);
nor U10953 (N_10953,N_10643,N_10626);
xor U10954 (N_10954,N_10712,N_10671);
nor U10955 (N_10955,N_10652,N_10780);
xor U10956 (N_10956,N_10615,N_10701);
nor U10957 (N_10957,N_10706,N_10701);
and U10958 (N_10958,N_10732,N_10657);
or U10959 (N_10959,N_10635,N_10797);
and U10960 (N_10960,N_10619,N_10720);
and U10961 (N_10961,N_10799,N_10669);
nor U10962 (N_10962,N_10604,N_10686);
or U10963 (N_10963,N_10720,N_10765);
or U10964 (N_10964,N_10640,N_10703);
xnor U10965 (N_10965,N_10637,N_10776);
or U10966 (N_10966,N_10740,N_10760);
or U10967 (N_10967,N_10607,N_10610);
or U10968 (N_10968,N_10710,N_10787);
xor U10969 (N_10969,N_10695,N_10758);
or U10970 (N_10970,N_10623,N_10680);
xor U10971 (N_10971,N_10725,N_10653);
nor U10972 (N_10972,N_10621,N_10628);
nor U10973 (N_10973,N_10749,N_10794);
nand U10974 (N_10974,N_10787,N_10606);
and U10975 (N_10975,N_10635,N_10685);
nand U10976 (N_10976,N_10659,N_10697);
xnor U10977 (N_10977,N_10725,N_10734);
and U10978 (N_10978,N_10707,N_10749);
xnor U10979 (N_10979,N_10639,N_10748);
and U10980 (N_10980,N_10756,N_10780);
nor U10981 (N_10981,N_10621,N_10615);
nor U10982 (N_10982,N_10703,N_10781);
nand U10983 (N_10983,N_10783,N_10702);
nand U10984 (N_10984,N_10717,N_10617);
xor U10985 (N_10985,N_10685,N_10607);
nand U10986 (N_10986,N_10618,N_10665);
nand U10987 (N_10987,N_10741,N_10772);
xnor U10988 (N_10988,N_10647,N_10768);
or U10989 (N_10989,N_10775,N_10639);
or U10990 (N_10990,N_10646,N_10748);
xor U10991 (N_10991,N_10611,N_10726);
or U10992 (N_10992,N_10642,N_10732);
and U10993 (N_10993,N_10611,N_10689);
or U10994 (N_10994,N_10646,N_10667);
nand U10995 (N_10995,N_10675,N_10764);
or U10996 (N_10996,N_10643,N_10735);
nor U10997 (N_10997,N_10626,N_10745);
nand U10998 (N_10998,N_10755,N_10798);
or U10999 (N_10999,N_10717,N_10699);
or U11000 (N_11000,N_10920,N_10951);
xnor U11001 (N_11001,N_10832,N_10834);
nor U11002 (N_11002,N_10986,N_10935);
nor U11003 (N_11003,N_10806,N_10898);
xor U11004 (N_11004,N_10840,N_10896);
xnor U11005 (N_11005,N_10821,N_10836);
nor U11006 (N_11006,N_10918,N_10838);
nand U11007 (N_11007,N_10844,N_10944);
and U11008 (N_11008,N_10833,N_10987);
and U11009 (N_11009,N_10881,N_10810);
nor U11010 (N_11010,N_10938,N_10850);
and U11011 (N_11011,N_10890,N_10965);
nor U11012 (N_11012,N_10801,N_10887);
nor U11013 (N_11013,N_10997,N_10961);
xor U11014 (N_11014,N_10830,N_10870);
and U11015 (N_11015,N_10979,N_10908);
and U11016 (N_11016,N_10919,N_10975);
nand U11017 (N_11017,N_10876,N_10846);
or U11018 (N_11018,N_10991,N_10839);
xor U11019 (N_11019,N_10863,N_10968);
nor U11020 (N_11020,N_10814,N_10827);
or U11021 (N_11021,N_10936,N_10861);
or U11022 (N_11022,N_10989,N_10928);
nand U11023 (N_11023,N_10958,N_10809);
or U11024 (N_11024,N_10963,N_10828);
nor U11025 (N_11025,N_10995,N_10868);
or U11026 (N_11026,N_10813,N_10990);
nand U11027 (N_11027,N_10962,N_10946);
nor U11028 (N_11028,N_10816,N_10931);
xor U11029 (N_11029,N_10800,N_10969);
xor U11030 (N_11030,N_10978,N_10815);
nor U11031 (N_11031,N_10903,N_10802);
nand U11032 (N_11032,N_10970,N_10880);
nor U11033 (N_11033,N_10947,N_10817);
nor U11034 (N_11034,N_10885,N_10912);
nand U11035 (N_11035,N_10929,N_10874);
nand U11036 (N_11036,N_10998,N_10917);
xnor U11037 (N_11037,N_10875,N_10824);
nor U11038 (N_11038,N_10825,N_10845);
nor U11039 (N_11039,N_10954,N_10945);
and U11040 (N_11040,N_10866,N_10909);
nand U11041 (N_11041,N_10983,N_10900);
and U11042 (N_11042,N_10973,N_10930);
and U11043 (N_11043,N_10932,N_10923);
and U11044 (N_11044,N_10822,N_10939);
nand U11045 (N_11045,N_10924,N_10872);
xnor U11046 (N_11046,N_10808,N_10843);
nor U11047 (N_11047,N_10882,N_10977);
nand U11048 (N_11048,N_10959,N_10829);
xor U11049 (N_11049,N_10867,N_10835);
nand U11050 (N_11050,N_10858,N_10904);
or U11051 (N_11051,N_10901,N_10811);
and U11052 (N_11052,N_10907,N_10883);
nor U11053 (N_11053,N_10807,N_10894);
or U11054 (N_11054,N_10860,N_10952);
nor U11055 (N_11055,N_10855,N_10878);
nor U11056 (N_11056,N_10902,N_10915);
and U11057 (N_11057,N_10950,N_10967);
nand U11058 (N_11058,N_10826,N_10842);
and U11059 (N_11059,N_10984,N_10857);
or U11060 (N_11060,N_10974,N_10999);
and U11061 (N_11061,N_10921,N_10862);
or U11062 (N_11062,N_10916,N_10992);
nand U11063 (N_11063,N_10893,N_10812);
and U11064 (N_11064,N_10966,N_10927);
nor U11065 (N_11065,N_10994,N_10864);
nand U11066 (N_11066,N_10888,N_10895);
or U11067 (N_11067,N_10933,N_10853);
and U11068 (N_11068,N_10926,N_10837);
and U11069 (N_11069,N_10976,N_10852);
nand U11070 (N_11070,N_10922,N_10911);
nor U11071 (N_11071,N_10892,N_10906);
nor U11072 (N_11072,N_10993,N_10971);
and U11073 (N_11073,N_10803,N_10905);
or U11074 (N_11074,N_10960,N_10982);
xor U11075 (N_11075,N_10856,N_10914);
nand U11076 (N_11076,N_10873,N_10879);
and U11077 (N_11077,N_10877,N_10957);
nor U11078 (N_11078,N_10831,N_10884);
nand U11079 (N_11079,N_10985,N_10942);
or U11080 (N_11080,N_10848,N_10820);
and U11081 (N_11081,N_10871,N_10988);
xor U11082 (N_11082,N_10851,N_10913);
nor U11083 (N_11083,N_10805,N_10948);
or U11084 (N_11084,N_10981,N_10891);
and U11085 (N_11085,N_10949,N_10934);
or U11086 (N_11086,N_10953,N_10943);
nand U11087 (N_11087,N_10940,N_10823);
nor U11088 (N_11088,N_10899,N_10937);
and U11089 (N_11089,N_10804,N_10964);
and U11090 (N_11090,N_10910,N_10847);
or U11091 (N_11091,N_10897,N_10849);
nand U11092 (N_11092,N_10941,N_10886);
or U11093 (N_11093,N_10818,N_10819);
or U11094 (N_11094,N_10972,N_10865);
xor U11095 (N_11095,N_10859,N_10925);
or U11096 (N_11096,N_10996,N_10869);
nor U11097 (N_11097,N_10980,N_10955);
nand U11098 (N_11098,N_10841,N_10854);
and U11099 (N_11099,N_10889,N_10956);
and U11100 (N_11100,N_10835,N_10895);
or U11101 (N_11101,N_10981,N_10922);
nor U11102 (N_11102,N_10900,N_10972);
or U11103 (N_11103,N_10865,N_10890);
xnor U11104 (N_11104,N_10813,N_10986);
or U11105 (N_11105,N_10895,N_10840);
nor U11106 (N_11106,N_10890,N_10802);
xor U11107 (N_11107,N_10870,N_10932);
nand U11108 (N_11108,N_10856,N_10821);
nor U11109 (N_11109,N_10849,N_10829);
nor U11110 (N_11110,N_10953,N_10889);
xor U11111 (N_11111,N_10842,N_10824);
or U11112 (N_11112,N_10994,N_10837);
nor U11113 (N_11113,N_10853,N_10953);
xor U11114 (N_11114,N_10862,N_10940);
xnor U11115 (N_11115,N_10801,N_10998);
or U11116 (N_11116,N_10900,N_10842);
and U11117 (N_11117,N_10823,N_10979);
nand U11118 (N_11118,N_10949,N_10870);
nand U11119 (N_11119,N_10991,N_10809);
nand U11120 (N_11120,N_10970,N_10873);
nor U11121 (N_11121,N_10832,N_10937);
or U11122 (N_11122,N_10881,N_10963);
and U11123 (N_11123,N_10934,N_10972);
xnor U11124 (N_11124,N_10807,N_10913);
or U11125 (N_11125,N_10931,N_10996);
nor U11126 (N_11126,N_10980,N_10933);
or U11127 (N_11127,N_10927,N_10931);
nor U11128 (N_11128,N_10853,N_10912);
or U11129 (N_11129,N_10833,N_10918);
or U11130 (N_11130,N_10887,N_10886);
nor U11131 (N_11131,N_10851,N_10985);
nor U11132 (N_11132,N_10809,N_10818);
xor U11133 (N_11133,N_10934,N_10832);
xnor U11134 (N_11134,N_10948,N_10802);
and U11135 (N_11135,N_10956,N_10989);
and U11136 (N_11136,N_10937,N_10822);
nand U11137 (N_11137,N_10849,N_10823);
nor U11138 (N_11138,N_10905,N_10973);
nand U11139 (N_11139,N_10842,N_10976);
and U11140 (N_11140,N_10822,N_10815);
nor U11141 (N_11141,N_10832,N_10825);
nor U11142 (N_11142,N_10909,N_10826);
and U11143 (N_11143,N_10842,N_10851);
nor U11144 (N_11144,N_10991,N_10831);
nor U11145 (N_11145,N_10930,N_10983);
nand U11146 (N_11146,N_10895,N_10811);
and U11147 (N_11147,N_10909,N_10837);
nand U11148 (N_11148,N_10912,N_10988);
xnor U11149 (N_11149,N_10931,N_10807);
nor U11150 (N_11150,N_10819,N_10892);
or U11151 (N_11151,N_10880,N_10889);
nor U11152 (N_11152,N_10910,N_10845);
nand U11153 (N_11153,N_10879,N_10840);
xor U11154 (N_11154,N_10957,N_10836);
or U11155 (N_11155,N_10817,N_10860);
xnor U11156 (N_11156,N_10992,N_10895);
and U11157 (N_11157,N_10825,N_10997);
and U11158 (N_11158,N_10951,N_10923);
nand U11159 (N_11159,N_10958,N_10995);
or U11160 (N_11160,N_10814,N_10965);
xor U11161 (N_11161,N_10828,N_10833);
and U11162 (N_11162,N_10991,N_10802);
nand U11163 (N_11163,N_10947,N_10992);
nand U11164 (N_11164,N_10933,N_10849);
nor U11165 (N_11165,N_10942,N_10884);
xnor U11166 (N_11166,N_10845,N_10859);
and U11167 (N_11167,N_10820,N_10903);
nor U11168 (N_11168,N_10946,N_10984);
or U11169 (N_11169,N_10818,N_10899);
or U11170 (N_11170,N_10966,N_10970);
nand U11171 (N_11171,N_10968,N_10827);
or U11172 (N_11172,N_10875,N_10800);
nand U11173 (N_11173,N_10969,N_10862);
nand U11174 (N_11174,N_10931,N_10838);
and U11175 (N_11175,N_10935,N_10906);
nor U11176 (N_11176,N_10962,N_10840);
and U11177 (N_11177,N_10901,N_10972);
and U11178 (N_11178,N_10992,N_10984);
xor U11179 (N_11179,N_10996,N_10876);
nor U11180 (N_11180,N_10829,N_10952);
xor U11181 (N_11181,N_10891,N_10895);
xor U11182 (N_11182,N_10814,N_10857);
and U11183 (N_11183,N_10999,N_10973);
xor U11184 (N_11184,N_10840,N_10845);
nor U11185 (N_11185,N_10875,N_10897);
and U11186 (N_11186,N_10879,N_10812);
xor U11187 (N_11187,N_10811,N_10886);
or U11188 (N_11188,N_10879,N_10903);
nand U11189 (N_11189,N_10825,N_10850);
or U11190 (N_11190,N_10988,N_10806);
xor U11191 (N_11191,N_10945,N_10932);
nor U11192 (N_11192,N_10968,N_10956);
xor U11193 (N_11193,N_10983,N_10856);
and U11194 (N_11194,N_10928,N_10867);
xnor U11195 (N_11195,N_10955,N_10925);
xnor U11196 (N_11196,N_10804,N_10888);
nor U11197 (N_11197,N_10925,N_10969);
nor U11198 (N_11198,N_10868,N_10863);
or U11199 (N_11199,N_10914,N_10984);
nor U11200 (N_11200,N_11195,N_11052);
and U11201 (N_11201,N_11046,N_11030);
or U11202 (N_11202,N_11071,N_11019);
nor U11203 (N_11203,N_11044,N_11074);
nor U11204 (N_11204,N_11197,N_11017);
and U11205 (N_11205,N_11142,N_11167);
and U11206 (N_11206,N_11118,N_11025);
and U11207 (N_11207,N_11063,N_11012);
nand U11208 (N_11208,N_11054,N_11156);
or U11209 (N_11209,N_11053,N_11005);
or U11210 (N_11210,N_11159,N_11043);
or U11211 (N_11211,N_11033,N_11069);
and U11212 (N_11212,N_11088,N_11080);
xnor U11213 (N_11213,N_11151,N_11163);
and U11214 (N_11214,N_11193,N_11048);
nand U11215 (N_11215,N_11014,N_11127);
and U11216 (N_11216,N_11113,N_11067);
nor U11217 (N_11217,N_11087,N_11196);
and U11218 (N_11218,N_11172,N_11082);
nand U11219 (N_11219,N_11031,N_11162);
nand U11220 (N_11220,N_11115,N_11021);
or U11221 (N_11221,N_11068,N_11157);
nand U11222 (N_11222,N_11002,N_11184);
and U11223 (N_11223,N_11171,N_11011);
nor U11224 (N_11224,N_11094,N_11060);
and U11225 (N_11225,N_11182,N_11050);
xor U11226 (N_11226,N_11018,N_11160);
or U11227 (N_11227,N_11190,N_11147);
and U11228 (N_11228,N_11004,N_11168);
nor U11229 (N_11229,N_11098,N_11103);
and U11230 (N_11230,N_11199,N_11089);
nor U11231 (N_11231,N_11008,N_11007);
or U11232 (N_11232,N_11149,N_11108);
nand U11233 (N_11233,N_11055,N_11116);
nor U11234 (N_11234,N_11148,N_11145);
nand U11235 (N_11235,N_11085,N_11102);
nand U11236 (N_11236,N_11020,N_11059);
or U11237 (N_11237,N_11003,N_11169);
nor U11238 (N_11238,N_11176,N_11039);
nor U11239 (N_11239,N_11180,N_11078);
nor U11240 (N_11240,N_11122,N_11064);
xnor U11241 (N_11241,N_11035,N_11049);
or U11242 (N_11242,N_11024,N_11126);
nand U11243 (N_11243,N_11010,N_11066);
nor U11244 (N_11244,N_11022,N_11016);
xor U11245 (N_11245,N_11164,N_11183);
xor U11246 (N_11246,N_11042,N_11161);
or U11247 (N_11247,N_11015,N_11106);
nand U11248 (N_11248,N_11137,N_11131);
nand U11249 (N_11249,N_11186,N_11029);
xnor U11250 (N_11250,N_11191,N_11105);
nor U11251 (N_11251,N_11194,N_11081);
or U11252 (N_11252,N_11075,N_11083);
nor U11253 (N_11253,N_11177,N_11136);
or U11254 (N_11254,N_11129,N_11170);
nand U11255 (N_11255,N_11144,N_11150);
and U11256 (N_11256,N_11155,N_11013);
and U11257 (N_11257,N_11092,N_11065);
or U11258 (N_11258,N_11109,N_11135);
nor U11259 (N_11259,N_11188,N_11198);
and U11260 (N_11260,N_11152,N_11045);
xor U11261 (N_11261,N_11100,N_11175);
or U11262 (N_11262,N_11097,N_11073);
or U11263 (N_11263,N_11036,N_11076);
and U11264 (N_11264,N_11166,N_11143);
nand U11265 (N_11265,N_11140,N_11112);
nor U11266 (N_11266,N_11146,N_11124);
nand U11267 (N_11267,N_11111,N_11099);
xor U11268 (N_11268,N_11090,N_11040);
and U11269 (N_11269,N_11041,N_11062);
or U11270 (N_11270,N_11077,N_11086);
and U11271 (N_11271,N_11091,N_11070);
nand U11272 (N_11272,N_11051,N_11173);
or U11273 (N_11273,N_11117,N_11178);
or U11274 (N_11274,N_11079,N_11189);
or U11275 (N_11275,N_11123,N_11138);
xor U11276 (N_11276,N_11139,N_11000);
xor U11277 (N_11277,N_11101,N_11125);
xnor U11278 (N_11278,N_11134,N_11027);
nor U11279 (N_11279,N_11130,N_11179);
and U11280 (N_11280,N_11120,N_11174);
xnor U11281 (N_11281,N_11093,N_11181);
and U11282 (N_11282,N_11121,N_11119);
nand U11283 (N_11283,N_11056,N_11132);
nand U11284 (N_11284,N_11128,N_11023);
nand U11285 (N_11285,N_11158,N_11107);
and U11286 (N_11286,N_11026,N_11009);
nand U11287 (N_11287,N_11028,N_11096);
xor U11288 (N_11288,N_11187,N_11006);
nor U11289 (N_11289,N_11047,N_11095);
nor U11290 (N_11290,N_11037,N_11034);
nand U11291 (N_11291,N_11061,N_11154);
xor U11292 (N_11292,N_11057,N_11038);
and U11293 (N_11293,N_11133,N_11072);
or U11294 (N_11294,N_11141,N_11058);
nand U11295 (N_11295,N_11114,N_11185);
or U11296 (N_11296,N_11153,N_11110);
nor U11297 (N_11297,N_11192,N_11165);
or U11298 (N_11298,N_11104,N_11001);
nor U11299 (N_11299,N_11084,N_11032);
or U11300 (N_11300,N_11026,N_11016);
and U11301 (N_11301,N_11131,N_11086);
xnor U11302 (N_11302,N_11090,N_11184);
nor U11303 (N_11303,N_11145,N_11042);
and U11304 (N_11304,N_11134,N_11057);
or U11305 (N_11305,N_11081,N_11006);
nor U11306 (N_11306,N_11095,N_11098);
nor U11307 (N_11307,N_11161,N_11084);
xor U11308 (N_11308,N_11176,N_11043);
xor U11309 (N_11309,N_11144,N_11035);
or U11310 (N_11310,N_11013,N_11148);
nand U11311 (N_11311,N_11177,N_11175);
and U11312 (N_11312,N_11009,N_11078);
and U11313 (N_11313,N_11143,N_11003);
nor U11314 (N_11314,N_11107,N_11119);
nand U11315 (N_11315,N_11150,N_11185);
and U11316 (N_11316,N_11023,N_11031);
or U11317 (N_11317,N_11154,N_11116);
or U11318 (N_11318,N_11165,N_11167);
xnor U11319 (N_11319,N_11158,N_11090);
and U11320 (N_11320,N_11158,N_11152);
xnor U11321 (N_11321,N_11170,N_11179);
nor U11322 (N_11322,N_11056,N_11157);
nand U11323 (N_11323,N_11080,N_11065);
xor U11324 (N_11324,N_11199,N_11042);
nand U11325 (N_11325,N_11198,N_11016);
and U11326 (N_11326,N_11147,N_11079);
or U11327 (N_11327,N_11196,N_11179);
or U11328 (N_11328,N_11159,N_11079);
or U11329 (N_11329,N_11116,N_11076);
and U11330 (N_11330,N_11010,N_11038);
and U11331 (N_11331,N_11195,N_11127);
xnor U11332 (N_11332,N_11178,N_11040);
and U11333 (N_11333,N_11168,N_11073);
nand U11334 (N_11334,N_11153,N_11172);
or U11335 (N_11335,N_11140,N_11176);
xnor U11336 (N_11336,N_11095,N_11139);
and U11337 (N_11337,N_11123,N_11112);
nor U11338 (N_11338,N_11113,N_11035);
or U11339 (N_11339,N_11124,N_11084);
xor U11340 (N_11340,N_11175,N_11185);
or U11341 (N_11341,N_11046,N_11156);
or U11342 (N_11342,N_11022,N_11065);
nand U11343 (N_11343,N_11074,N_11167);
nor U11344 (N_11344,N_11055,N_11133);
nand U11345 (N_11345,N_11180,N_11006);
nand U11346 (N_11346,N_11105,N_11090);
nand U11347 (N_11347,N_11146,N_11096);
nor U11348 (N_11348,N_11197,N_11035);
and U11349 (N_11349,N_11048,N_11009);
xor U11350 (N_11350,N_11145,N_11116);
and U11351 (N_11351,N_11025,N_11076);
and U11352 (N_11352,N_11163,N_11066);
and U11353 (N_11353,N_11102,N_11172);
and U11354 (N_11354,N_11191,N_11064);
or U11355 (N_11355,N_11030,N_11092);
xnor U11356 (N_11356,N_11185,N_11074);
nand U11357 (N_11357,N_11144,N_11028);
nand U11358 (N_11358,N_11096,N_11186);
and U11359 (N_11359,N_11045,N_11170);
nor U11360 (N_11360,N_11170,N_11159);
nor U11361 (N_11361,N_11087,N_11048);
nand U11362 (N_11362,N_11019,N_11013);
xor U11363 (N_11363,N_11131,N_11193);
xor U11364 (N_11364,N_11063,N_11120);
nor U11365 (N_11365,N_11090,N_11009);
nor U11366 (N_11366,N_11109,N_11102);
nand U11367 (N_11367,N_11145,N_11129);
nand U11368 (N_11368,N_11013,N_11152);
xor U11369 (N_11369,N_11048,N_11139);
and U11370 (N_11370,N_11031,N_11010);
xnor U11371 (N_11371,N_11165,N_11128);
nor U11372 (N_11372,N_11195,N_11076);
and U11373 (N_11373,N_11129,N_11001);
or U11374 (N_11374,N_11075,N_11085);
nor U11375 (N_11375,N_11115,N_11104);
nand U11376 (N_11376,N_11134,N_11126);
nand U11377 (N_11377,N_11057,N_11028);
xnor U11378 (N_11378,N_11006,N_11194);
xnor U11379 (N_11379,N_11079,N_11033);
or U11380 (N_11380,N_11085,N_11082);
nor U11381 (N_11381,N_11072,N_11118);
nand U11382 (N_11382,N_11122,N_11190);
or U11383 (N_11383,N_11048,N_11196);
xnor U11384 (N_11384,N_11042,N_11039);
xor U11385 (N_11385,N_11116,N_11135);
or U11386 (N_11386,N_11090,N_11066);
nand U11387 (N_11387,N_11087,N_11003);
or U11388 (N_11388,N_11074,N_11090);
or U11389 (N_11389,N_11045,N_11059);
or U11390 (N_11390,N_11054,N_11095);
or U11391 (N_11391,N_11155,N_11118);
nor U11392 (N_11392,N_11033,N_11162);
xor U11393 (N_11393,N_11119,N_11023);
or U11394 (N_11394,N_11111,N_11049);
xor U11395 (N_11395,N_11161,N_11086);
nor U11396 (N_11396,N_11023,N_11091);
xnor U11397 (N_11397,N_11083,N_11092);
nand U11398 (N_11398,N_11017,N_11098);
nand U11399 (N_11399,N_11162,N_11161);
xor U11400 (N_11400,N_11327,N_11348);
and U11401 (N_11401,N_11370,N_11258);
nor U11402 (N_11402,N_11344,N_11218);
and U11403 (N_11403,N_11378,N_11393);
nand U11404 (N_11404,N_11245,N_11354);
and U11405 (N_11405,N_11294,N_11306);
or U11406 (N_11406,N_11203,N_11215);
and U11407 (N_11407,N_11238,N_11376);
nand U11408 (N_11408,N_11338,N_11261);
nor U11409 (N_11409,N_11364,N_11275);
xor U11410 (N_11410,N_11267,N_11304);
or U11411 (N_11411,N_11228,N_11325);
and U11412 (N_11412,N_11207,N_11384);
nand U11413 (N_11413,N_11232,N_11334);
xor U11414 (N_11414,N_11230,N_11315);
xor U11415 (N_11415,N_11291,N_11358);
xnor U11416 (N_11416,N_11367,N_11309);
nand U11417 (N_11417,N_11337,N_11310);
xor U11418 (N_11418,N_11229,N_11254);
nor U11419 (N_11419,N_11336,N_11270);
xor U11420 (N_11420,N_11278,N_11302);
nor U11421 (N_11421,N_11339,N_11242);
nand U11422 (N_11422,N_11368,N_11298);
nand U11423 (N_11423,N_11365,N_11382);
and U11424 (N_11424,N_11255,N_11269);
or U11425 (N_11425,N_11293,N_11347);
nor U11426 (N_11426,N_11305,N_11287);
nor U11427 (N_11427,N_11226,N_11231);
nand U11428 (N_11428,N_11394,N_11271);
nand U11429 (N_11429,N_11353,N_11324);
and U11430 (N_11430,N_11395,N_11379);
or U11431 (N_11431,N_11239,N_11280);
and U11432 (N_11432,N_11221,N_11352);
nor U11433 (N_11433,N_11371,N_11385);
xnor U11434 (N_11434,N_11276,N_11251);
xor U11435 (N_11435,N_11388,N_11316);
nand U11436 (N_11436,N_11292,N_11274);
nor U11437 (N_11437,N_11329,N_11330);
and U11438 (N_11438,N_11248,N_11256);
nand U11439 (N_11439,N_11277,N_11219);
nor U11440 (N_11440,N_11204,N_11297);
or U11441 (N_11441,N_11345,N_11321);
and U11442 (N_11442,N_11260,N_11244);
nand U11443 (N_11443,N_11361,N_11213);
and U11444 (N_11444,N_11381,N_11268);
xnor U11445 (N_11445,N_11296,N_11363);
nor U11446 (N_11446,N_11224,N_11286);
nor U11447 (N_11447,N_11257,N_11240);
nand U11448 (N_11448,N_11216,N_11279);
or U11449 (N_11449,N_11366,N_11225);
nand U11450 (N_11450,N_11283,N_11234);
nor U11451 (N_11451,N_11317,N_11308);
xor U11452 (N_11452,N_11399,N_11300);
and U11453 (N_11453,N_11375,N_11272);
nand U11454 (N_11454,N_11243,N_11335);
and U11455 (N_11455,N_11266,N_11202);
or U11456 (N_11456,N_11214,N_11200);
and U11457 (N_11457,N_11397,N_11343);
and U11458 (N_11458,N_11212,N_11252);
xnor U11459 (N_11459,N_11360,N_11357);
or U11460 (N_11460,N_11217,N_11398);
or U11461 (N_11461,N_11295,N_11211);
xor U11462 (N_11462,N_11355,N_11246);
and U11463 (N_11463,N_11391,N_11359);
or U11464 (N_11464,N_11265,N_11220);
nor U11465 (N_11465,N_11311,N_11326);
nor U11466 (N_11466,N_11333,N_11284);
or U11467 (N_11467,N_11386,N_11303);
and U11468 (N_11468,N_11247,N_11262);
nand U11469 (N_11469,N_11320,N_11223);
and U11470 (N_11470,N_11342,N_11289);
and U11471 (N_11471,N_11235,N_11383);
xor U11472 (N_11472,N_11377,N_11322);
and U11473 (N_11473,N_11374,N_11273);
xnor U11474 (N_11474,N_11372,N_11233);
and U11475 (N_11475,N_11288,N_11341);
nor U11476 (N_11476,N_11249,N_11206);
xor U11477 (N_11477,N_11222,N_11227);
and U11478 (N_11478,N_11328,N_11373);
nand U11479 (N_11479,N_11318,N_11362);
or U11480 (N_11480,N_11253,N_11299);
xor U11481 (N_11481,N_11346,N_11369);
nand U11482 (N_11482,N_11281,N_11392);
nor U11483 (N_11483,N_11209,N_11210);
xnor U11484 (N_11484,N_11351,N_11350);
nand U11485 (N_11485,N_11340,N_11241);
and U11486 (N_11486,N_11319,N_11250);
nor U11487 (N_11487,N_11263,N_11331);
and U11488 (N_11488,N_11390,N_11282);
or U11489 (N_11489,N_11356,N_11205);
nand U11490 (N_11490,N_11236,N_11389);
nor U11491 (N_11491,N_11314,N_11208);
nor U11492 (N_11492,N_11332,N_11290);
nand U11493 (N_11493,N_11264,N_11285);
nor U11494 (N_11494,N_11396,N_11301);
and U11495 (N_11495,N_11349,N_11201);
or U11496 (N_11496,N_11237,N_11380);
xor U11497 (N_11497,N_11307,N_11312);
or U11498 (N_11498,N_11387,N_11313);
or U11499 (N_11499,N_11259,N_11323);
and U11500 (N_11500,N_11207,N_11301);
or U11501 (N_11501,N_11309,N_11248);
xor U11502 (N_11502,N_11360,N_11392);
or U11503 (N_11503,N_11345,N_11287);
and U11504 (N_11504,N_11216,N_11277);
xor U11505 (N_11505,N_11343,N_11308);
or U11506 (N_11506,N_11319,N_11207);
xnor U11507 (N_11507,N_11372,N_11258);
or U11508 (N_11508,N_11264,N_11376);
or U11509 (N_11509,N_11387,N_11382);
nor U11510 (N_11510,N_11279,N_11211);
or U11511 (N_11511,N_11399,N_11298);
or U11512 (N_11512,N_11273,N_11267);
nor U11513 (N_11513,N_11265,N_11348);
nor U11514 (N_11514,N_11313,N_11255);
nand U11515 (N_11515,N_11243,N_11368);
and U11516 (N_11516,N_11207,N_11388);
xnor U11517 (N_11517,N_11279,N_11275);
nor U11518 (N_11518,N_11371,N_11290);
and U11519 (N_11519,N_11239,N_11211);
nand U11520 (N_11520,N_11211,N_11361);
xor U11521 (N_11521,N_11265,N_11367);
and U11522 (N_11522,N_11273,N_11247);
nor U11523 (N_11523,N_11344,N_11338);
or U11524 (N_11524,N_11268,N_11316);
or U11525 (N_11525,N_11228,N_11305);
and U11526 (N_11526,N_11262,N_11290);
and U11527 (N_11527,N_11257,N_11293);
xor U11528 (N_11528,N_11261,N_11226);
and U11529 (N_11529,N_11204,N_11353);
nor U11530 (N_11530,N_11222,N_11215);
or U11531 (N_11531,N_11226,N_11257);
or U11532 (N_11532,N_11219,N_11303);
or U11533 (N_11533,N_11344,N_11222);
or U11534 (N_11534,N_11392,N_11208);
or U11535 (N_11535,N_11398,N_11379);
and U11536 (N_11536,N_11277,N_11314);
nand U11537 (N_11537,N_11381,N_11339);
nor U11538 (N_11538,N_11211,N_11212);
or U11539 (N_11539,N_11216,N_11252);
nand U11540 (N_11540,N_11360,N_11331);
nor U11541 (N_11541,N_11208,N_11232);
and U11542 (N_11542,N_11383,N_11280);
nor U11543 (N_11543,N_11282,N_11374);
nand U11544 (N_11544,N_11316,N_11225);
and U11545 (N_11545,N_11202,N_11200);
nand U11546 (N_11546,N_11392,N_11275);
and U11547 (N_11547,N_11290,N_11291);
nor U11548 (N_11548,N_11318,N_11298);
or U11549 (N_11549,N_11239,N_11261);
nor U11550 (N_11550,N_11388,N_11329);
nor U11551 (N_11551,N_11264,N_11288);
or U11552 (N_11552,N_11242,N_11308);
nor U11553 (N_11553,N_11249,N_11377);
xnor U11554 (N_11554,N_11210,N_11273);
nand U11555 (N_11555,N_11249,N_11327);
nor U11556 (N_11556,N_11299,N_11294);
nor U11557 (N_11557,N_11318,N_11345);
and U11558 (N_11558,N_11227,N_11220);
or U11559 (N_11559,N_11307,N_11273);
or U11560 (N_11560,N_11253,N_11380);
and U11561 (N_11561,N_11395,N_11255);
and U11562 (N_11562,N_11322,N_11372);
nand U11563 (N_11563,N_11335,N_11340);
nand U11564 (N_11564,N_11280,N_11271);
nand U11565 (N_11565,N_11332,N_11239);
and U11566 (N_11566,N_11257,N_11242);
nor U11567 (N_11567,N_11335,N_11363);
or U11568 (N_11568,N_11324,N_11334);
nor U11569 (N_11569,N_11222,N_11207);
xor U11570 (N_11570,N_11375,N_11227);
xor U11571 (N_11571,N_11317,N_11208);
nand U11572 (N_11572,N_11337,N_11309);
xor U11573 (N_11573,N_11230,N_11347);
nor U11574 (N_11574,N_11251,N_11266);
or U11575 (N_11575,N_11259,N_11308);
xnor U11576 (N_11576,N_11235,N_11309);
and U11577 (N_11577,N_11254,N_11241);
and U11578 (N_11578,N_11217,N_11213);
nand U11579 (N_11579,N_11213,N_11249);
and U11580 (N_11580,N_11311,N_11212);
xor U11581 (N_11581,N_11340,N_11350);
xor U11582 (N_11582,N_11240,N_11380);
xnor U11583 (N_11583,N_11300,N_11342);
nand U11584 (N_11584,N_11253,N_11338);
or U11585 (N_11585,N_11337,N_11383);
or U11586 (N_11586,N_11359,N_11311);
or U11587 (N_11587,N_11222,N_11276);
xnor U11588 (N_11588,N_11272,N_11355);
and U11589 (N_11589,N_11376,N_11314);
nand U11590 (N_11590,N_11345,N_11202);
nand U11591 (N_11591,N_11267,N_11213);
xnor U11592 (N_11592,N_11290,N_11308);
nand U11593 (N_11593,N_11228,N_11389);
or U11594 (N_11594,N_11264,N_11250);
xnor U11595 (N_11595,N_11219,N_11335);
xnor U11596 (N_11596,N_11215,N_11252);
or U11597 (N_11597,N_11392,N_11302);
xnor U11598 (N_11598,N_11377,N_11269);
nor U11599 (N_11599,N_11242,N_11226);
nand U11600 (N_11600,N_11499,N_11522);
and U11601 (N_11601,N_11508,N_11476);
or U11602 (N_11602,N_11430,N_11560);
nand U11603 (N_11603,N_11518,N_11491);
nor U11604 (N_11604,N_11484,N_11489);
xor U11605 (N_11605,N_11497,N_11597);
nand U11606 (N_11606,N_11524,N_11593);
nand U11607 (N_11607,N_11485,N_11556);
nand U11608 (N_11608,N_11490,N_11561);
nand U11609 (N_11609,N_11441,N_11423);
nand U11610 (N_11610,N_11465,N_11553);
nor U11611 (N_11611,N_11510,N_11534);
and U11612 (N_11612,N_11535,N_11589);
or U11613 (N_11613,N_11580,N_11543);
xnor U11614 (N_11614,N_11462,N_11448);
or U11615 (N_11615,N_11449,N_11502);
or U11616 (N_11616,N_11509,N_11526);
and U11617 (N_11617,N_11411,N_11408);
nand U11618 (N_11618,N_11487,N_11416);
and U11619 (N_11619,N_11488,N_11467);
or U11620 (N_11620,N_11514,N_11594);
or U11621 (N_11621,N_11463,N_11520);
nand U11622 (N_11622,N_11532,N_11472);
and U11623 (N_11623,N_11421,N_11453);
and U11624 (N_11624,N_11460,N_11440);
nand U11625 (N_11625,N_11422,N_11405);
nand U11626 (N_11626,N_11574,N_11576);
or U11627 (N_11627,N_11447,N_11595);
or U11628 (N_11628,N_11400,N_11505);
and U11629 (N_11629,N_11470,N_11598);
nand U11630 (N_11630,N_11541,N_11578);
nand U11631 (N_11631,N_11434,N_11538);
xor U11632 (N_11632,N_11419,N_11555);
nand U11633 (N_11633,N_11410,N_11503);
xnor U11634 (N_11634,N_11468,N_11500);
nor U11635 (N_11635,N_11572,N_11481);
xnor U11636 (N_11636,N_11455,N_11540);
nand U11637 (N_11637,N_11542,N_11401);
nand U11638 (N_11638,N_11436,N_11480);
or U11639 (N_11639,N_11588,N_11512);
xor U11640 (N_11640,N_11424,N_11412);
xnor U11641 (N_11641,N_11471,N_11523);
nor U11642 (N_11642,N_11404,N_11426);
xor U11643 (N_11643,N_11511,N_11494);
or U11644 (N_11644,N_11516,N_11566);
xor U11645 (N_11645,N_11452,N_11482);
or U11646 (N_11646,N_11483,N_11564);
xnor U11647 (N_11647,N_11461,N_11429);
or U11648 (N_11648,N_11547,N_11517);
nand U11649 (N_11649,N_11591,N_11415);
nor U11650 (N_11650,N_11439,N_11562);
nand U11651 (N_11651,N_11456,N_11443);
nand U11652 (N_11652,N_11486,N_11528);
and U11653 (N_11653,N_11457,N_11446);
or U11654 (N_11654,N_11464,N_11582);
nand U11655 (N_11655,N_11552,N_11466);
and U11656 (N_11656,N_11563,N_11417);
and U11657 (N_11657,N_11406,N_11513);
nand U11658 (N_11658,N_11496,N_11533);
xor U11659 (N_11659,N_11557,N_11437);
nand U11660 (N_11660,N_11568,N_11495);
xor U11661 (N_11661,N_11550,N_11565);
or U11662 (N_11662,N_11587,N_11573);
xor U11663 (N_11663,N_11402,N_11435);
or U11664 (N_11664,N_11530,N_11432);
or U11665 (N_11665,N_11519,N_11585);
nor U11666 (N_11666,N_11409,N_11442);
nor U11667 (N_11667,N_11549,N_11586);
xnor U11668 (N_11668,N_11407,N_11403);
and U11669 (N_11669,N_11444,N_11438);
or U11670 (N_11670,N_11569,N_11433);
xor U11671 (N_11671,N_11599,N_11531);
or U11672 (N_11672,N_11473,N_11420);
nor U11673 (N_11673,N_11567,N_11474);
and U11674 (N_11674,N_11575,N_11581);
nand U11675 (N_11675,N_11479,N_11537);
nand U11676 (N_11676,N_11525,N_11504);
nand U11677 (N_11677,N_11584,N_11529);
and U11678 (N_11678,N_11425,N_11431);
and U11679 (N_11679,N_11558,N_11451);
nor U11680 (N_11680,N_11428,N_11527);
xor U11681 (N_11681,N_11413,N_11507);
and U11682 (N_11682,N_11459,N_11536);
or U11683 (N_11683,N_11427,N_11515);
or U11684 (N_11684,N_11478,N_11521);
xnor U11685 (N_11685,N_11498,N_11551);
and U11686 (N_11686,N_11596,N_11570);
and U11687 (N_11687,N_11544,N_11546);
or U11688 (N_11688,N_11592,N_11454);
and U11689 (N_11689,N_11545,N_11590);
xnor U11690 (N_11690,N_11577,N_11559);
nand U11691 (N_11691,N_11469,N_11571);
xnor U11692 (N_11692,N_11450,N_11418);
or U11693 (N_11693,N_11539,N_11414);
nand U11694 (N_11694,N_11506,N_11493);
xnor U11695 (N_11695,N_11492,N_11583);
and U11696 (N_11696,N_11548,N_11458);
nor U11697 (N_11697,N_11501,N_11554);
nand U11698 (N_11698,N_11579,N_11475);
nor U11699 (N_11699,N_11477,N_11445);
and U11700 (N_11700,N_11467,N_11518);
nand U11701 (N_11701,N_11457,N_11406);
xor U11702 (N_11702,N_11472,N_11572);
nor U11703 (N_11703,N_11535,N_11471);
and U11704 (N_11704,N_11571,N_11477);
and U11705 (N_11705,N_11488,N_11443);
nor U11706 (N_11706,N_11484,N_11542);
or U11707 (N_11707,N_11483,N_11571);
xnor U11708 (N_11708,N_11483,N_11461);
and U11709 (N_11709,N_11439,N_11519);
nor U11710 (N_11710,N_11540,N_11490);
nand U11711 (N_11711,N_11514,N_11566);
or U11712 (N_11712,N_11441,N_11476);
nor U11713 (N_11713,N_11555,N_11552);
or U11714 (N_11714,N_11534,N_11493);
nor U11715 (N_11715,N_11405,N_11534);
and U11716 (N_11716,N_11486,N_11492);
xnor U11717 (N_11717,N_11451,N_11457);
xor U11718 (N_11718,N_11511,N_11468);
nor U11719 (N_11719,N_11585,N_11419);
nand U11720 (N_11720,N_11570,N_11512);
nor U11721 (N_11721,N_11533,N_11545);
xor U11722 (N_11722,N_11449,N_11435);
or U11723 (N_11723,N_11481,N_11474);
xor U11724 (N_11724,N_11547,N_11413);
xnor U11725 (N_11725,N_11559,N_11545);
xor U11726 (N_11726,N_11401,N_11482);
nand U11727 (N_11727,N_11543,N_11468);
xor U11728 (N_11728,N_11457,N_11578);
and U11729 (N_11729,N_11538,N_11405);
nor U11730 (N_11730,N_11462,N_11542);
or U11731 (N_11731,N_11434,N_11593);
nor U11732 (N_11732,N_11422,N_11587);
or U11733 (N_11733,N_11455,N_11553);
and U11734 (N_11734,N_11588,N_11480);
nand U11735 (N_11735,N_11505,N_11513);
or U11736 (N_11736,N_11506,N_11545);
nor U11737 (N_11737,N_11593,N_11532);
or U11738 (N_11738,N_11449,N_11478);
nor U11739 (N_11739,N_11520,N_11536);
and U11740 (N_11740,N_11447,N_11414);
xnor U11741 (N_11741,N_11566,N_11577);
nand U11742 (N_11742,N_11440,N_11550);
and U11743 (N_11743,N_11436,N_11583);
nor U11744 (N_11744,N_11577,N_11598);
xnor U11745 (N_11745,N_11562,N_11529);
and U11746 (N_11746,N_11567,N_11530);
or U11747 (N_11747,N_11448,N_11567);
nand U11748 (N_11748,N_11491,N_11542);
nand U11749 (N_11749,N_11411,N_11535);
xor U11750 (N_11750,N_11521,N_11542);
or U11751 (N_11751,N_11441,N_11413);
nand U11752 (N_11752,N_11518,N_11488);
nand U11753 (N_11753,N_11462,N_11449);
or U11754 (N_11754,N_11498,N_11599);
and U11755 (N_11755,N_11465,N_11437);
nor U11756 (N_11756,N_11443,N_11492);
or U11757 (N_11757,N_11549,N_11459);
or U11758 (N_11758,N_11414,N_11598);
nand U11759 (N_11759,N_11464,N_11481);
nand U11760 (N_11760,N_11466,N_11553);
xnor U11761 (N_11761,N_11488,N_11406);
nor U11762 (N_11762,N_11441,N_11494);
xnor U11763 (N_11763,N_11586,N_11512);
or U11764 (N_11764,N_11459,N_11496);
nand U11765 (N_11765,N_11421,N_11540);
or U11766 (N_11766,N_11453,N_11403);
or U11767 (N_11767,N_11422,N_11493);
nand U11768 (N_11768,N_11525,N_11519);
and U11769 (N_11769,N_11470,N_11487);
nand U11770 (N_11770,N_11461,N_11553);
nand U11771 (N_11771,N_11400,N_11549);
nor U11772 (N_11772,N_11584,N_11512);
xnor U11773 (N_11773,N_11557,N_11566);
or U11774 (N_11774,N_11593,N_11572);
xor U11775 (N_11775,N_11467,N_11572);
or U11776 (N_11776,N_11420,N_11466);
nor U11777 (N_11777,N_11439,N_11498);
or U11778 (N_11778,N_11586,N_11452);
and U11779 (N_11779,N_11473,N_11443);
xnor U11780 (N_11780,N_11483,N_11438);
xor U11781 (N_11781,N_11412,N_11536);
xor U11782 (N_11782,N_11592,N_11562);
nor U11783 (N_11783,N_11579,N_11542);
nor U11784 (N_11784,N_11409,N_11468);
xor U11785 (N_11785,N_11474,N_11495);
xor U11786 (N_11786,N_11445,N_11594);
xor U11787 (N_11787,N_11534,N_11598);
nand U11788 (N_11788,N_11423,N_11479);
or U11789 (N_11789,N_11579,N_11431);
nand U11790 (N_11790,N_11521,N_11594);
nand U11791 (N_11791,N_11572,N_11599);
or U11792 (N_11792,N_11585,N_11550);
nor U11793 (N_11793,N_11407,N_11562);
nand U11794 (N_11794,N_11551,N_11550);
xor U11795 (N_11795,N_11415,N_11515);
or U11796 (N_11796,N_11455,N_11551);
and U11797 (N_11797,N_11414,N_11566);
xor U11798 (N_11798,N_11535,N_11432);
and U11799 (N_11799,N_11400,N_11552);
or U11800 (N_11800,N_11760,N_11659);
xnor U11801 (N_11801,N_11726,N_11662);
xor U11802 (N_11802,N_11787,N_11754);
xor U11803 (N_11803,N_11668,N_11703);
nand U11804 (N_11804,N_11674,N_11764);
xnor U11805 (N_11805,N_11691,N_11628);
xnor U11806 (N_11806,N_11742,N_11644);
nand U11807 (N_11807,N_11684,N_11686);
nor U11808 (N_11808,N_11707,N_11601);
xnor U11809 (N_11809,N_11763,N_11692);
nor U11810 (N_11810,N_11779,N_11716);
nand U11811 (N_11811,N_11788,N_11685);
nand U11812 (N_11812,N_11743,N_11609);
nand U11813 (N_11813,N_11734,N_11654);
and U11814 (N_11814,N_11617,N_11664);
nand U11815 (N_11815,N_11634,N_11652);
nand U11816 (N_11816,N_11629,N_11759);
and U11817 (N_11817,N_11665,N_11649);
and U11818 (N_11818,N_11778,N_11728);
or U11819 (N_11819,N_11783,N_11675);
nor U11820 (N_11820,N_11711,N_11637);
or U11821 (N_11821,N_11614,N_11635);
xnor U11822 (N_11822,N_11640,N_11616);
nand U11823 (N_11823,N_11768,N_11706);
xnor U11824 (N_11824,N_11749,N_11639);
nand U11825 (N_11825,N_11653,N_11702);
xor U11826 (N_11826,N_11750,N_11736);
and U11827 (N_11827,N_11758,N_11751);
nand U11828 (N_11828,N_11713,N_11618);
and U11829 (N_11829,N_11735,N_11648);
and U11830 (N_11830,N_11766,N_11689);
and U11831 (N_11831,N_11602,N_11714);
nand U11832 (N_11832,N_11770,N_11796);
xor U11833 (N_11833,N_11789,N_11776);
or U11834 (N_11834,N_11670,N_11730);
xnor U11835 (N_11835,N_11645,N_11781);
and U11836 (N_11836,N_11688,N_11721);
and U11837 (N_11837,N_11641,N_11625);
or U11838 (N_11838,N_11679,N_11697);
xor U11839 (N_11839,N_11704,N_11615);
and U11840 (N_11840,N_11606,N_11693);
nor U11841 (N_11841,N_11677,N_11744);
nand U11842 (N_11842,N_11636,N_11699);
nor U11843 (N_11843,N_11701,N_11723);
and U11844 (N_11844,N_11633,N_11785);
nor U11845 (N_11845,N_11666,N_11769);
or U11846 (N_11846,N_11620,N_11612);
or U11847 (N_11847,N_11738,N_11604);
or U11848 (N_11848,N_11798,N_11746);
and U11849 (N_11849,N_11650,N_11772);
and U11850 (N_11850,N_11727,N_11718);
nand U11851 (N_11851,N_11739,N_11792);
or U11852 (N_11852,N_11700,N_11761);
xnor U11853 (N_11853,N_11762,N_11627);
nand U11854 (N_11854,N_11780,N_11740);
nand U11855 (N_11855,N_11729,N_11756);
and U11856 (N_11856,N_11773,N_11724);
xnor U11857 (N_11857,N_11791,N_11624);
nor U11858 (N_11858,N_11682,N_11782);
or U11859 (N_11859,N_11709,N_11630);
nor U11860 (N_11860,N_11611,N_11632);
and U11861 (N_11861,N_11671,N_11622);
or U11862 (N_11862,N_11715,N_11698);
xnor U11863 (N_11863,N_11748,N_11631);
and U11864 (N_11864,N_11676,N_11708);
and U11865 (N_11865,N_11799,N_11667);
xnor U11866 (N_11866,N_11673,N_11603);
nand U11867 (N_11867,N_11794,N_11757);
or U11868 (N_11868,N_11720,N_11681);
xor U11869 (N_11869,N_11605,N_11643);
xnor U11870 (N_11870,N_11680,N_11790);
xor U11871 (N_11871,N_11663,N_11745);
nor U11872 (N_11872,N_11646,N_11719);
nor U11873 (N_11873,N_11775,N_11705);
and U11874 (N_11874,N_11657,N_11747);
xor U11875 (N_11875,N_11610,N_11786);
nand U11876 (N_11876,N_11755,N_11784);
xnor U11877 (N_11877,N_11765,N_11690);
or U11878 (N_11878,N_11658,N_11793);
xor U11879 (N_11879,N_11607,N_11725);
nand U11880 (N_11880,N_11717,N_11600);
xor U11881 (N_11881,N_11638,N_11733);
nor U11882 (N_11882,N_11647,N_11613);
xnor U11883 (N_11883,N_11777,N_11623);
nor U11884 (N_11884,N_11737,N_11687);
nand U11885 (N_11885,N_11678,N_11621);
xor U11886 (N_11886,N_11722,N_11672);
nand U11887 (N_11887,N_11642,N_11669);
and U11888 (N_11888,N_11797,N_11767);
xor U11889 (N_11889,N_11753,N_11741);
or U11890 (N_11890,N_11661,N_11774);
nand U11891 (N_11891,N_11694,N_11683);
and U11892 (N_11892,N_11655,N_11608);
xnor U11893 (N_11893,N_11752,N_11710);
xor U11894 (N_11894,N_11656,N_11732);
xnor U11895 (N_11895,N_11626,N_11731);
or U11896 (N_11896,N_11712,N_11696);
nor U11897 (N_11897,N_11771,N_11660);
and U11898 (N_11898,N_11651,N_11795);
nand U11899 (N_11899,N_11695,N_11619);
nand U11900 (N_11900,N_11687,N_11660);
xnor U11901 (N_11901,N_11761,N_11725);
nor U11902 (N_11902,N_11766,N_11613);
nor U11903 (N_11903,N_11699,N_11772);
or U11904 (N_11904,N_11668,N_11644);
nand U11905 (N_11905,N_11656,N_11739);
or U11906 (N_11906,N_11608,N_11694);
nand U11907 (N_11907,N_11779,N_11767);
xor U11908 (N_11908,N_11661,N_11687);
or U11909 (N_11909,N_11682,N_11720);
nor U11910 (N_11910,N_11738,N_11705);
and U11911 (N_11911,N_11645,N_11741);
or U11912 (N_11912,N_11798,N_11617);
nor U11913 (N_11913,N_11702,N_11724);
nor U11914 (N_11914,N_11753,N_11779);
or U11915 (N_11915,N_11757,N_11623);
and U11916 (N_11916,N_11755,N_11608);
or U11917 (N_11917,N_11703,N_11601);
xnor U11918 (N_11918,N_11655,N_11702);
nand U11919 (N_11919,N_11697,N_11765);
or U11920 (N_11920,N_11601,N_11610);
nor U11921 (N_11921,N_11696,N_11695);
and U11922 (N_11922,N_11607,N_11648);
xnor U11923 (N_11923,N_11644,N_11737);
xnor U11924 (N_11924,N_11614,N_11607);
nor U11925 (N_11925,N_11797,N_11779);
nor U11926 (N_11926,N_11725,N_11605);
or U11927 (N_11927,N_11686,N_11624);
xor U11928 (N_11928,N_11613,N_11717);
xor U11929 (N_11929,N_11712,N_11610);
xor U11930 (N_11930,N_11765,N_11602);
xor U11931 (N_11931,N_11786,N_11721);
nand U11932 (N_11932,N_11719,N_11750);
or U11933 (N_11933,N_11638,N_11780);
and U11934 (N_11934,N_11729,N_11733);
xor U11935 (N_11935,N_11603,N_11707);
and U11936 (N_11936,N_11785,N_11763);
and U11937 (N_11937,N_11668,N_11675);
or U11938 (N_11938,N_11702,N_11730);
nand U11939 (N_11939,N_11797,N_11785);
nor U11940 (N_11940,N_11601,N_11698);
and U11941 (N_11941,N_11741,N_11752);
nand U11942 (N_11942,N_11766,N_11639);
nand U11943 (N_11943,N_11625,N_11686);
nand U11944 (N_11944,N_11652,N_11651);
or U11945 (N_11945,N_11736,N_11623);
and U11946 (N_11946,N_11623,N_11629);
nand U11947 (N_11947,N_11750,N_11746);
nand U11948 (N_11948,N_11702,N_11779);
nor U11949 (N_11949,N_11621,N_11764);
and U11950 (N_11950,N_11682,N_11745);
or U11951 (N_11951,N_11783,N_11695);
and U11952 (N_11952,N_11619,N_11640);
and U11953 (N_11953,N_11714,N_11716);
nand U11954 (N_11954,N_11608,N_11609);
nand U11955 (N_11955,N_11636,N_11732);
and U11956 (N_11956,N_11713,N_11756);
nor U11957 (N_11957,N_11767,N_11621);
and U11958 (N_11958,N_11659,N_11720);
or U11959 (N_11959,N_11689,N_11672);
nand U11960 (N_11960,N_11738,N_11786);
and U11961 (N_11961,N_11632,N_11720);
nand U11962 (N_11962,N_11751,N_11637);
xor U11963 (N_11963,N_11798,N_11607);
or U11964 (N_11964,N_11676,N_11642);
and U11965 (N_11965,N_11631,N_11644);
nand U11966 (N_11966,N_11733,N_11682);
and U11967 (N_11967,N_11646,N_11625);
xnor U11968 (N_11968,N_11752,N_11626);
nand U11969 (N_11969,N_11792,N_11709);
nor U11970 (N_11970,N_11759,N_11712);
or U11971 (N_11971,N_11666,N_11692);
nor U11972 (N_11972,N_11603,N_11754);
nor U11973 (N_11973,N_11609,N_11666);
or U11974 (N_11974,N_11785,N_11687);
or U11975 (N_11975,N_11689,N_11683);
nor U11976 (N_11976,N_11638,N_11771);
nor U11977 (N_11977,N_11656,N_11652);
or U11978 (N_11978,N_11777,N_11683);
nor U11979 (N_11979,N_11793,N_11761);
nor U11980 (N_11980,N_11622,N_11652);
xnor U11981 (N_11981,N_11637,N_11695);
and U11982 (N_11982,N_11627,N_11743);
or U11983 (N_11983,N_11637,N_11775);
and U11984 (N_11984,N_11760,N_11723);
nor U11985 (N_11985,N_11680,N_11635);
nor U11986 (N_11986,N_11728,N_11784);
nand U11987 (N_11987,N_11751,N_11683);
and U11988 (N_11988,N_11739,N_11729);
and U11989 (N_11989,N_11762,N_11713);
xnor U11990 (N_11990,N_11722,N_11678);
or U11991 (N_11991,N_11792,N_11751);
or U11992 (N_11992,N_11799,N_11791);
xnor U11993 (N_11993,N_11607,N_11698);
nand U11994 (N_11994,N_11717,N_11615);
or U11995 (N_11995,N_11742,N_11758);
xnor U11996 (N_11996,N_11721,N_11702);
xor U11997 (N_11997,N_11746,N_11730);
xnor U11998 (N_11998,N_11765,N_11745);
and U11999 (N_11999,N_11772,N_11745);
nand U12000 (N_12000,N_11926,N_11979);
and U12001 (N_12001,N_11889,N_11930);
xnor U12002 (N_12002,N_11876,N_11984);
and U12003 (N_12003,N_11936,N_11809);
nor U12004 (N_12004,N_11818,N_11929);
or U12005 (N_12005,N_11968,N_11865);
and U12006 (N_12006,N_11967,N_11831);
xnor U12007 (N_12007,N_11909,N_11855);
or U12008 (N_12008,N_11966,N_11942);
nand U12009 (N_12009,N_11888,N_11923);
nor U12010 (N_12010,N_11849,N_11802);
or U12011 (N_12011,N_11801,N_11952);
and U12012 (N_12012,N_11907,N_11971);
xor U12013 (N_12013,N_11974,N_11875);
or U12014 (N_12014,N_11981,N_11994);
nand U12015 (N_12015,N_11864,N_11985);
nand U12016 (N_12016,N_11975,N_11805);
nor U12017 (N_12017,N_11877,N_11867);
nor U12018 (N_12018,N_11949,N_11870);
nand U12019 (N_12019,N_11814,N_11822);
nor U12020 (N_12020,N_11950,N_11919);
and U12021 (N_12021,N_11914,N_11808);
or U12022 (N_12022,N_11963,N_11838);
or U12023 (N_12023,N_11921,N_11991);
nor U12024 (N_12024,N_11955,N_11862);
or U12025 (N_12025,N_11938,N_11941);
nand U12026 (N_12026,N_11885,N_11839);
or U12027 (N_12027,N_11937,N_11866);
or U12028 (N_12028,N_11816,N_11881);
xor U12029 (N_12029,N_11863,N_11844);
or U12030 (N_12030,N_11846,N_11810);
xor U12031 (N_12031,N_11961,N_11990);
and U12032 (N_12032,N_11946,N_11807);
nor U12033 (N_12033,N_11986,N_11860);
nand U12034 (N_12034,N_11964,N_11958);
nor U12035 (N_12035,N_11900,N_11912);
nand U12036 (N_12036,N_11983,N_11918);
or U12037 (N_12037,N_11886,N_11944);
xor U12038 (N_12038,N_11819,N_11848);
xnor U12039 (N_12039,N_11934,N_11882);
nand U12040 (N_12040,N_11834,N_11940);
nor U12041 (N_12041,N_11891,N_11970);
nor U12042 (N_12042,N_11957,N_11911);
and U12043 (N_12043,N_11962,N_11917);
nand U12044 (N_12044,N_11976,N_11995);
nand U12045 (N_12045,N_11851,N_11933);
or U12046 (N_12046,N_11993,N_11910);
xor U12047 (N_12047,N_11916,N_11813);
xnor U12048 (N_12048,N_11825,N_11803);
nand U12049 (N_12049,N_11965,N_11823);
nand U12050 (N_12050,N_11943,N_11956);
xnor U12051 (N_12051,N_11817,N_11811);
or U12052 (N_12052,N_11883,N_11879);
nand U12053 (N_12053,N_11806,N_11827);
or U12054 (N_12054,N_11924,N_11913);
or U12055 (N_12055,N_11977,N_11939);
xor U12056 (N_12056,N_11898,N_11932);
nor U12057 (N_12057,N_11892,N_11953);
nor U12058 (N_12058,N_11880,N_11947);
nor U12059 (N_12059,N_11821,N_11854);
xnor U12060 (N_12060,N_11904,N_11843);
nand U12061 (N_12061,N_11987,N_11897);
or U12062 (N_12062,N_11928,N_11873);
and U12063 (N_12063,N_11894,N_11812);
xor U12064 (N_12064,N_11905,N_11842);
xor U12065 (N_12065,N_11973,N_11887);
nand U12066 (N_12066,N_11997,N_11954);
xnor U12067 (N_12067,N_11982,N_11832);
and U12068 (N_12068,N_11858,N_11830);
nand U12069 (N_12069,N_11815,N_11895);
or U12070 (N_12070,N_11925,N_11906);
and U12071 (N_12071,N_11980,N_11874);
xor U12072 (N_12072,N_11972,N_11902);
xnor U12073 (N_12073,N_11996,N_11890);
nor U12074 (N_12074,N_11804,N_11969);
nor U12075 (N_12075,N_11989,N_11959);
or U12076 (N_12076,N_11853,N_11857);
nand U12077 (N_12077,N_11869,N_11960);
or U12078 (N_12078,N_11931,N_11868);
and U12079 (N_12079,N_11903,N_11836);
nor U12080 (N_12080,N_11820,N_11847);
xnor U12081 (N_12081,N_11837,N_11840);
xor U12082 (N_12082,N_11978,N_11872);
and U12083 (N_12083,N_11999,N_11861);
or U12084 (N_12084,N_11951,N_11878);
nor U12085 (N_12085,N_11988,N_11845);
nor U12086 (N_12086,N_11920,N_11992);
nand U12087 (N_12087,N_11859,N_11901);
nand U12088 (N_12088,N_11948,N_11998);
and U12089 (N_12089,N_11829,N_11871);
or U12090 (N_12090,N_11908,N_11893);
and U12091 (N_12091,N_11824,N_11896);
nand U12092 (N_12092,N_11850,N_11835);
nand U12093 (N_12093,N_11935,N_11841);
and U12094 (N_12094,N_11828,N_11884);
and U12095 (N_12095,N_11927,N_11852);
or U12096 (N_12096,N_11833,N_11915);
nand U12097 (N_12097,N_11826,N_11899);
nor U12098 (N_12098,N_11945,N_11922);
xnor U12099 (N_12099,N_11856,N_11800);
nand U12100 (N_12100,N_11951,N_11880);
and U12101 (N_12101,N_11865,N_11848);
xnor U12102 (N_12102,N_11832,N_11941);
or U12103 (N_12103,N_11898,N_11849);
or U12104 (N_12104,N_11949,N_11821);
nor U12105 (N_12105,N_11821,N_11974);
or U12106 (N_12106,N_11922,N_11965);
or U12107 (N_12107,N_11963,N_11821);
xnor U12108 (N_12108,N_11816,N_11927);
nor U12109 (N_12109,N_11984,N_11987);
nand U12110 (N_12110,N_11884,N_11981);
or U12111 (N_12111,N_11866,N_11978);
nand U12112 (N_12112,N_11819,N_11956);
nor U12113 (N_12113,N_11972,N_11818);
and U12114 (N_12114,N_11905,N_11801);
and U12115 (N_12115,N_11989,N_11913);
xnor U12116 (N_12116,N_11936,N_11912);
nand U12117 (N_12117,N_11998,N_11876);
xor U12118 (N_12118,N_11890,N_11886);
nor U12119 (N_12119,N_11877,N_11946);
xor U12120 (N_12120,N_11820,N_11887);
or U12121 (N_12121,N_11885,N_11989);
nand U12122 (N_12122,N_11829,N_11855);
and U12123 (N_12123,N_11981,N_11870);
and U12124 (N_12124,N_11848,N_11890);
or U12125 (N_12125,N_11875,N_11962);
nand U12126 (N_12126,N_11873,N_11896);
and U12127 (N_12127,N_11935,N_11863);
nand U12128 (N_12128,N_11911,N_11841);
and U12129 (N_12129,N_11819,N_11840);
or U12130 (N_12130,N_11977,N_11841);
nor U12131 (N_12131,N_11869,N_11827);
nand U12132 (N_12132,N_11870,N_11886);
nand U12133 (N_12133,N_11835,N_11918);
xor U12134 (N_12134,N_11969,N_11930);
nor U12135 (N_12135,N_11919,N_11967);
xor U12136 (N_12136,N_11985,N_11807);
nor U12137 (N_12137,N_11874,N_11942);
nand U12138 (N_12138,N_11991,N_11904);
nor U12139 (N_12139,N_11845,N_11869);
or U12140 (N_12140,N_11945,N_11999);
and U12141 (N_12141,N_11924,N_11849);
xnor U12142 (N_12142,N_11878,N_11836);
or U12143 (N_12143,N_11871,N_11821);
and U12144 (N_12144,N_11898,N_11949);
or U12145 (N_12145,N_11847,N_11947);
and U12146 (N_12146,N_11975,N_11832);
or U12147 (N_12147,N_11964,N_11913);
or U12148 (N_12148,N_11977,N_11830);
or U12149 (N_12149,N_11813,N_11902);
or U12150 (N_12150,N_11940,N_11946);
nor U12151 (N_12151,N_11973,N_11997);
nand U12152 (N_12152,N_11831,N_11901);
or U12153 (N_12153,N_11966,N_11912);
or U12154 (N_12154,N_11864,N_11861);
xor U12155 (N_12155,N_11999,N_11900);
and U12156 (N_12156,N_11875,N_11816);
xnor U12157 (N_12157,N_11908,N_11995);
or U12158 (N_12158,N_11966,N_11834);
or U12159 (N_12159,N_11987,N_11845);
or U12160 (N_12160,N_11931,N_11844);
nand U12161 (N_12161,N_11822,N_11940);
nand U12162 (N_12162,N_11953,N_11861);
nor U12163 (N_12163,N_11858,N_11940);
xnor U12164 (N_12164,N_11840,N_11846);
xnor U12165 (N_12165,N_11958,N_11849);
xnor U12166 (N_12166,N_11827,N_11993);
or U12167 (N_12167,N_11956,N_11816);
nor U12168 (N_12168,N_11971,N_11801);
xor U12169 (N_12169,N_11920,N_11824);
nor U12170 (N_12170,N_11940,N_11964);
and U12171 (N_12171,N_11974,N_11814);
nand U12172 (N_12172,N_11887,N_11846);
nand U12173 (N_12173,N_11854,N_11863);
and U12174 (N_12174,N_11899,N_11845);
nand U12175 (N_12175,N_11883,N_11913);
xnor U12176 (N_12176,N_11990,N_11932);
nand U12177 (N_12177,N_11805,N_11827);
nand U12178 (N_12178,N_11967,N_11911);
and U12179 (N_12179,N_11869,N_11882);
and U12180 (N_12180,N_11973,N_11920);
nand U12181 (N_12181,N_11882,N_11881);
nand U12182 (N_12182,N_11821,N_11828);
and U12183 (N_12183,N_11891,N_11903);
nor U12184 (N_12184,N_11909,N_11979);
or U12185 (N_12185,N_11834,N_11898);
or U12186 (N_12186,N_11819,N_11876);
or U12187 (N_12187,N_11802,N_11818);
and U12188 (N_12188,N_11854,N_11910);
or U12189 (N_12189,N_11933,N_11807);
and U12190 (N_12190,N_11872,N_11982);
nand U12191 (N_12191,N_11994,N_11982);
or U12192 (N_12192,N_11840,N_11862);
nor U12193 (N_12193,N_11838,N_11893);
nand U12194 (N_12194,N_11861,N_11977);
nand U12195 (N_12195,N_11961,N_11943);
and U12196 (N_12196,N_11910,N_11876);
xnor U12197 (N_12197,N_11890,N_11831);
xnor U12198 (N_12198,N_11882,N_11933);
or U12199 (N_12199,N_11936,N_11907);
and U12200 (N_12200,N_12111,N_12090);
nor U12201 (N_12201,N_12129,N_12061);
xnor U12202 (N_12202,N_12065,N_12126);
nor U12203 (N_12203,N_12094,N_12143);
xnor U12204 (N_12204,N_12142,N_12085);
xor U12205 (N_12205,N_12165,N_12071);
xor U12206 (N_12206,N_12150,N_12058);
xor U12207 (N_12207,N_12175,N_12192);
xnor U12208 (N_12208,N_12104,N_12154);
or U12209 (N_12209,N_12123,N_12169);
nor U12210 (N_12210,N_12188,N_12108);
and U12211 (N_12211,N_12029,N_12190);
and U12212 (N_12212,N_12109,N_12124);
and U12213 (N_12213,N_12055,N_12146);
and U12214 (N_12214,N_12189,N_12044);
and U12215 (N_12215,N_12046,N_12014);
or U12216 (N_12216,N_12196,N_12103);
and U12217 (N_12217,N_12005,N_12186);
nand U12218 (N_12218,N_12114,N_12092);
xor U12219 (N_12219,N_12102,N_12031);
and U12220 (N_12220,N_12032,N_12183);
and U12221 (N_12221,N_12054,N_12132);
or U12222 (N_12222,N_12130,N_12067);
or U12223 (N_12223,N_12101,N_12088);
nand U12224 (N_12224,N_12069,N_12135);
nor U12225 (N_12225,N_12082,N_12195);
xor U12226 (N_12226,N_12068,N_12034);
xnor U12227 (N_12227,N_12181,N_12073);
and U12228 (N_12228,N_12157,N_12095);
and U12229 (N_12229,N_12149,N_12078);
nand U12230 (N_12230,N_12030,N_12180);
and U12231 (N_12231,N_12053,N_12127);
nand U12232 (N_12232,N_12076,N_12019);
and U12233 (N_12233,N_12139,N_12152);
or U12234 (N_12234,N_12096,N_12170);
and U12235 (N_12235,N_12084,N_12017);
nor U12236 (N_12236,N_12159,N_12059);
and U12237 (N_12237,N_12194,N_12125);
or U12238 (N_12238,N_12107,N_12145);
xnor U12239 (N_12239,N_12039,N_12110);
or U12240 (N_12240,N_12026,N_12003);
or U12241 (N_12241,N_12037,N_12010);
xor U12242 (N_12242,N_12160,N_12177);
nor U12243 (N_12243,N_12122,N_12072);
xor U12244 (N_12244,N_12155,N_12070);
xnor U12245 (N_12245,N_12040,N_12021);
or U12246 (N_12246,N_12156,N_12052);
or U12247 (N_12247,N_12178,N_12057);
nor U12248 (N_12248,N_12041,N_12133);
xor U12249 (N_12249,N_12042,N_12027);
and U12250 (N_12250,N_12171,N_12063);
or U12251 (N_12251,N_12161,N_12011);
nor U12252 (N_12252,N_12187,N_12064);
and U12253 (N_12253,N_12038,N_12047);
nand U12254 (N_12254,N_12147,N_12164);
and U12255 (N_12255,N_12079,N_12174);
nand U12256 (N_12256,N_12080,N_12148);
and U12257 (N_12257,N_12086,N_12167);
or U12258 (N_12258,N_12006,N_12136);
and U12259 (N_12259,N_12120,N_12004);
xor U12260 (N_12260,N_12013,N_12001);
nor U12261 (N_12261,N_12134,N_12153);
nor U12262 (N_12262,N_12117,N_12179);
nor U12263 (N_12263,N_12199,N_12028);
and U12264 (N_12264,N_12131,N_12191);
and U12265 (N_12265,N_12115,N_12007);
xnor U12266 (N_12266,N_12158,N_12024);
nand U12267 (N_12267,N_12193,N_12043);
and U12268 (N_12268,N_12118,N_12062);
nand U12269 (N_12269,N_12151,N_12106);
xor U12270 (N_12270,N_12018,N_12050);
and U12271 (N_12271,N_12012,N_12002);
nand U12272 (N_12272,N_12098,N_12128);
xnor U12273 (N_12273,N_12141,N_12066);
nand U12274 (N_12274,N_12144,N_12009);
nand U12275 (N_12275,N_12087,N_12045);
or U12276 (N_12276,N_12051,N_12198);
nand U12277 (N_12277,N_12099,N_12138);
and U12278 (N_12278,N_12035,N_12137);
nand U12279 (N_12279,N_12182,N_12000);
nand U12280 (N_12280,N_12091,N_12056);
xnor U12281 (N_12281,N_12168,N_12116);
xor U12282 (N_12282,N_12162,N_12081);
xnor U12283 (N_12283,N_12197,N_12166);
or U12284 (N_12284,N_12016,N_12060);
nor U12285 (N_12285,N_12172,N_12048);
nand U12286 (N_12286,N_12176,N_12097);
nand U12287 (N_12287,N_12077,N_12020);
or U12288 (N_12288,N_12075,N_12074);
and U12289 (N_12289,N_12173,N_12036);
or U12290 (N_12290,N_12184,N_12015);
nand U12291 (N_12291,N_12083,N_12025);
xnor U12292 (N_12292,N_12185,N_12121);
nor U12293 (N_12293,N_12105,N_12023);
nand U12294 (N_12294,N_12119,N_12089);
xnor U12295 (N_12295,N_12049,N_12008);
xnor U12296 (N_12296,N_12113,N_12100);
nor U12297 (N_12297,N_12163,N_12022);
nor U12298 (N_12298,N_12112,N_12140);
and U12299 (N_12299,N_12033,N_12093);
nand U12300 (N_12300,N_12061,N_12103);
nand U12301 (N_12301,N_12142,N_12051);
and U12302 (N_12302,N_12118,N_12153);
and U12303 (N_12303,N_12145,N_12198);
and U12304 (N_12304,N_12147,N_12165);
nor U12305 (N_12305,N_12145,N_12014);
nand U12306 (N_12306,N_12081,N_12138);
xnor U12307 (N_12307,N_12184,N_12035);
or U12308 (N_12308,N_12046,N_12176);
nand U12309 (N_12309,N_12049,N_12138);
nor U12310 (N_12310,N_12073,N_12098);
nand U12311 (N_12311,N_12118,N_12015);
nor U12312 (N_12312,N_12065,N_12149);
xnor U12313 (N_12313,N_12168,N_12043);
xnor U12314 (N_12314,N_12098,N_12052);
or U12315 (N_12315,N_12088,N_12023);
and U12316 (N_12316,N_12147,N_12086);
nor U12317 (N_12317,N_12104,N_12155);
and U12318 (N_12318,N_12035,N_12043);
xor U12319 (N_12319,N_12126,N_12070);
and U12320 (N_12320,N_12021,N_12156);
or U12321 (N_12321,N_12081,N_12008);
nand U12322 (N_12322,N_12181,N_12001);
xnor U12323 (N_12323,N_12127,N_12078);
nand U12324 (N_12324,N_12109,N_12176);
or U12325 (N_12325,N_12049,N_12080);
xnor U12326 (N_12326,N_12013,N_12105);
xor U12327 (N_12327,N_12176,N_12126);
and U12328 (N_12328,N_12035,N_12028);
and U12329 (N_12329,N_12134,N_12013);
nor U12330 (N_12330,N_12151,N_12005);
nor U12331 (N_12331,N_12190,N_12053);
nor U12332 (N_12332,N_12047,N_12177);
and U12333 (N_12333,N_12185,N_12017);
nor U12334 (N_12334,N_12186,N_12068);
nand U12335 (N_12335,N_12076,N_12185);
xnor U12336 (N_12336,N_12168,N_12046);
xnor U12337 (N_12337,N_12020,N_12004);
and U12338 (N_12338,N_12188,N_12132);
nand U12339 (N_12339,N_12008,N_12123);
xor U12340 (N_12340,N_12092,N_12174);
xnor U12341 (N_12341,N_12022,N_12013);
nand U12342 (N_12342,N_12068,N_12120);
and U12343 (N_12343,N_12183,N_12035);
and U12344 (N_12344,N_12158,N_12100);
nor U12345 (N_12345,N_12013,N_12029);
and U12346 (N_12346,N_12013,N_12040);
nor U12347 (N_12347,N_12011,N_12059);
nand U12348 (N_12348,N_12118,N_12192);
nand U12349 (N_12349,N_12081,N_12113);
xor U12350 (N_12350,N_12030,N_12110);
nor U12351 (N_12351,N_12118,N_12132);
and U12352 (N_12352,N_12035,N_12078);
xor U12353 (N_12353,N_12190,N_12195);
nor U12354 (N_12354,N_12079,N_12120);
nor U12355 (N_12355,N_12125,N_12028);
nor U12356 (N_12356,N_12003,N_12070);
and U12357 (N_12357,N_12081,N_12137);
xor U12358 (N_12358,N_12104,N_12015);
nor U12359 (N_12359,N_12193,N_12024);
xor U12360 (N_12360,N_12157,N_12161);
nand U12361 (N_12361,N_12025,N_12052);
nor U12362 (N_12362,N_12127,N_12030);
or U12363 (N_12363,N_12131,N_12067);
nor U12364 (N_12364,N_12072,N_12180);
nand U12365 (N_12365,N_12175,N_12086);
and U12366 (N_12366,N_12133,N_12050);
or U12367 (N_12367,N_12116,N_12187);
or U12368 (N_12368,N_12164,N_12171);
xor U12369 (N_12369,N_12137,N_12020);
or U12370 (N_12370,N_12008,N_12078);
nand U12371 (N_12371,N_12043,N_12147);
xor U12372 (N_12372,N_12025,N_12054);
and U12373 (N_12373,N_12018,N_12195);
nand U12374 (N_12374,N_12120,N_12196);
and U12375 (N_12375,N_12130,N_12199);
and U12376 (N_12376,N_12101,N_12184);
nand U12377 (N_12377,N_12179,N_12142);
xor U12378 (N_12378,N_12047,N_12041);
and U12379 (N_12379,N_12199,N_12069);
nand U12380 (N_12380,N_12175,N_12107);
nor U12381 (N_12381,N_12031,N_12161);
nor U12382 (N_12382,N_12152,N_12024);
or U12383 (N_12383,N_12191,N_12132);
xor U12384 (N_12384,N_12108,N_12065);
or U12385 (N_12385,N_12044,N_12013);
and U12386 (N_12386,N_12027,N_12153);
nand U12387 (N_12387,N_12016,N_12032);
nor U12388 (N_12388,N_12182,N_12120);
or U12389 (N_12389,N_12122,N_12081);
or U12390 (N_12390,N_12059,N_12187);
nand U12391 (N_12391,N_12178,N_12152);
and U12392 (N_12392,N_12169,N_12083);
or U12393 (N_12393,N_12040,N_12167);
nand U12394 (N_12394,N_12029,N_12119);
and U12395 (N_12395,N_12085,N_12175);
nor U12396 (N_12396,N_12054,N_12019);
nor U12397 (N_12397,N_12157,N_12111);
or U12398 (N_12398,N_12058,N_12105);
nand U12399 (N_12399,N_12152,N_12186);
or U12400 (N_12400,N_12312,N_12349);
or U12401 (N_12401,N_12395,N_12339);
nand U12402 (N_12402,N_12207,N_12314);
nor U12403 (N_12403,N_12383,N_12391);
xor U12404 (N_12404,N_12264,N_12374);
xor U12405 (N_12405,N_12239,N_12318);
or U12406 (N_12406,N_12371,N_12352);
and U12407 (N_12407,N_12233,N_12222);
and U12408 (N_12408,N_12386,N_12321);
and U12409 (N_12409,N_12240,N_12385);
nand U12410 (N_12410,N_12364,N_12235);
and U12411 (N_12411,N_12320,N_12229);
or U12412 (N_12412,N_12389,N_12242);
or U12413 (N_12413,N_12357,N_12367);
nand U12414 (N_12414,N_12319,N_12382);
nor U12415 (N_12415,N_12204,N_12377);
nor U12416 (N_12416,N_12288,N_12201);
and U12417 (N_12417,N_12297,N_12211);
xnor U12418 (N_12418,N_12337,N_12263);
nor U12419 (N_12419,N_12252,N_12330);
or U12420 (N_12420,N_12244,N_12203);
and U12421 (N_12421,N_12311,N_12202);
and U12422 (N_12422,N_12296,N_12209);
or U12423 (N_12423,N_12380,N_12375);
and U12424 (N_12424,N_12336,N_12206);
xor U12425 (N_12425,N_12226,N_12373);
or U12426 (N_12426,N_12213,N_12208);
nand U12427 (N_12427,N_12258,N_12309);
nor U12428 (N_12428,N_12248,N_12228);
xnor U12429 (N_12429,N_12295,N_12398);
nor U12430 (N_12430,N_12259,N_12266);
and U12431 (N_12431,N_12344,N_12232);
xor U12432 (N_12432,N_12351,N_12269);
and U12433 (N_12433,N_12348,N_12246);
nand U12434 (N_12434,N_12200,N_12326);
xor U12435 (N_12435,N_12260,N_12363);
or U12436 (N_12436,N_12335,N_12315);
and U12437 (N_12437,N_12217,N_12331);
or U12438 (N_12438,N_12298,N_12212);
xnor U12439 (N_12439,N_12234,N_12343);
xor U12440 (N_12440,N_12238,N_12341);
nor U12441 (N_12441,N_12275,N_12270);
nor U12442 (N_12442,N_12265,N_12280);
and U12443 (N_12443,N_12334,N_12274);
xnor U12444 (N_12444,N_12362,N_12291);
nor U12445 (N_12445,N_12305,N_12237);
nor U12446 (N_12446,N_12210,N_12300);
or U12447 (N_12447,N_12254,N_12243);
xnor U12448 (N_12448,N_12227,N_12359);
nand U12449 (N_12449,N_12340,N_12354);
xnor U12450 (N_12450,N_12327,N_12215);
xor U12451 (N_12451,N_12366,N_12281);
and U12452 (N_12452,N_12332,N_12286);
nor U12453 (N_12453,N_12325,N_12308);
nor U12454 (N_12454,N_12249,N_12282);
nor U12455 (N_12455,N_12292,N_12310);
nor U12456 (N_12456,N_12294,N_12276);
nand U12457 (N_12457,N_12333,N_12283);
nand U12458 (N_12458,N_12221,N_12390);
nand U12459 (N_12459,N_12342,N_12353);
nor U12460 (N_12460,N_12247,N_12220);
nor U12461 (N_12461,N_12316,N_12378);
nor U12462 (N_12462,N_12345,N_12278);
and U12463 (N_12463,N_12306,N_12271);
or U12464 (N_12464,N_12223,N_12301);
nand U12465 (N_12465,N_12329,N_12360);
xnor U12466 (N_12466,N_12272,N_12290);
or U12467 (N_12467,N_12392,N_12324);
xnor U12468 (N_12468,N_12225,N_12284);
or U12469 (N_12469,N_12356,N_12287);
or U12470 (N_12470,N_12273,N_12379);
nand U12471 (N_12471,N_12350,N_12257);
nand U12472 (N_12472,N_12256,N_12313);
nand U12473 (N_12473,N_12396,N_12381);
xor U12474 (N_12474,N_12255,N_12224);
nor U12475 (N_12475,N_12304,N_12368);
or U12476 (N_12476,N_12338,N_12230);
xnor U12477 (N_12477,N_12393,N_12236);
xnor U12478 (N_12478,N_12279,N_12268);
and U12479 (N_12479,N_12388,N_12251);
nor U12480 (N_12480,N_12369,N_12376);
nor U12481 (N_12481,N_12372,N_12328);
nor U12482 (N_12482,N_12358,N_12262);
or U12483 (N_12483,N_12384,N_12250);
xnor U12484 (N_12484,N_12245,N_12293);
xnor U12485 (N_12485,N_12231,N_12299);
nand U12486 (N_12486,N_12355,N_12399);
xnor U12487 (N_12487,N_12277,N_12397);
nor U12488 (N_12488,N_12394,N_12307);
and U12489 (N_12489,N_12214,N_12289);
and U12490 (N_12490,N_12285,N_12205);
xor U12491 (N_12491,N_12365,N_12323);
or U12492 (N_12492,N_12261,N_12322);
or U12493 (N_12493,N_12387,N_12347);
xor U12494 (N_12494,N_12267,N_12253);
and U12495 (N_12495,N_12219,N_12218);
xnor U12496 (N_12496,N_12346,N_12370);
xnor U12497 (N_12497,N_12241,N_12317);
nor U12498 (N_12498,N_12216,N_12361);
nor U12499 (N_12499,N_12303,N_12302);
or U12500 (N_12500,N_12225,N_12302);
nor U12501 (N_12501,N_12307,N_12233);
nand U12502 (N_12502,N_12350,N_12248);
xor U12503 (N_12503,N_12395,N_12255);
xor U12504 (N_12504,N_12293,N_12226);
nor U12505 (N_12505,N_12279,N_12372);
nor U12506 (N_12506,N_12381,N_12259);
or U12507 (N_12507,N_12287,N_12274);
nand U12508 (N_12508,N_12355,N_12262);
and U12509 (N_12509,N_12331,N_12324);
nand U12510 (N_12510,N_12306,N_12210);
xor U12511 (N_12511,N_12354,N_12360);
or U12512 (N_12512,N_12275,N_12328);
or U12513 (N_12513,N_12205,N_12341);
xor U12514 (N_12514,N_12352,N_12303);
and U12515 (N_12515,N_12380,N_12348);
nand U12516 (N_12516,N_12261,N_12367);
nor U12517 (N_12517,N_12226,N_12362);
nor U12518 (N_12518,N_12270,N_12380);
and U12519 (N_12519,N_12319,N_12260);
and U12520 (N_12520,N_12358,N_12274);
or U12521 (N_12521,N_12293,N_12316);
or U12522 (N_12522,N_12357,N_12261);
nor U12523 (N_12523,N_12335,N_12329);
or U12524 (N_12524,N_12300,N_12325);
and U12525 (N_12525,N_12215,N_12250);
or U12526 (N_12526,N_12398,N_12216);
nor U12527 (N_12527,N_12270,N_12269);
and U12528 (N_12528,N_12280,N_12262);
and U12529 (N_12529,N_12217,N_12399);
or U12530 (N_12530,N_12323,N_12344);
and U12531 (N_12531,N_12324,N_12242);
nand U12532 (N_12532,N_12319,N_12315);
xnor U12533 (N_12533,N_12388,N_12309);
nor U12534 (N_12534,N_12200,N_12224);
nand U12535 (N_12535,N_12290,N_12327);
and U12536 (N_12536,N_12314,N_12245);
xor U12537 (N_12537,N_12362,N_12391);
xor U12538 (N_12538,N_12246,N_12398);
nor U12539 (N_12539,N_12296,N_12213);
or U12540 (N_12540,N_12344,N_12251);
and U12541 (N_12541,N_12205,N_12224);
nand U12542 (N_12542,N_12310,N_12257);
nand U12543 (N_12543,N_12208,N_12276);
xnor U12544 (N_12544,N_12335,N_12233);
and U12545 (N_12545,N_12241,N_12247);
and U12546 (N_12546,N_12378,N_12237);
nand U12547 (N_12547,N_12317,N_12356);
nand U12548 (N_12548,N_12212,N_12277);
and U12549 (N_12549,N_12394,N_12240);
and U12550 (N_12550,N_12273,N_12390);
or U12551 (N_12551,N_12380,N_12343);
nor U12552 (N_12552,N_12304,N_12257);
or U12553 (N_12553,N_12215,N_12289);
xor U12554 (N_12554,N_12322,N_12271);
xor U12555 (N_12555,N_12299,N_12343);
xor U12556 (N_12556,N_12369,N_12210);
and U12557 (N_12557,N_12244,N_12369);
or U12558 (N_12558,N_12257,N_12318);
nor U12559 (N_12559,N_12245,N_12279);
nor U12560 (N_12560,N_12297,N_12236);
nand U12561 (N_12561,N_12222,N_12280);
nor U12562 (N_12562,N_12201,N_12251);
nand U12563 (N_12563,N_12381,N_12308);
nor U12564 (N_12564,N_12390,N_12367);
and U12565 (N_12565,N_12217,N_12253);
nand U12566 (N_12566,N_12222,N_12242);
and U12567 (N_12567,N_12367,N_12311);
nand U12568 (N_12568,N_12261,N_12392);
and U12569 (N_12569,N_12399,N_12224);
nand U12570 (N_12570,N_12251,N_12339);
nor U12571 (N_12571,N_12245,N_12261);
nand U12572 (N_12572,N_12381,N_12235);
nand U12573 (N_12573,N_12377,N_12328);
or U12574 (N_12574,N_12260,N_12271);
nand U12575 (N_12575,N_12385,N_12380);
or U12576 (N_12576,N_12398,N_12262);
and U12577 (N_12577,N_12227,N_12371);
or U12578 (N_12578,N_12282,N_12293);
and U12579 (N_12579,N_12394,N_12285);
or U12580 (N_12580,N_12347,N_12300);
and U12581 (N_12581,N_12209,N_12388);
or U12582 (N_12582,N_12388,N_12213);
and U12583 (N_12583,N_12223,N_12215);
or U12584 (N_12584,N_12377,N_12289);
nor U12585 (N_12585,N_12245,N_12322);
and U12586 (N_12586,N_12220,N_12273);
nor U12587 (N_12587,N_12281,N_12291);
nor U12588 (N_12588,N_12206,N_12322);
or U12589 (N_12589,N_12365,N_12201);
and U12590 (N_12590,N_12255,N_12334);
nor U12591 (N_12591,N_12223,N_12267);
or U12592 (N_12592,N_12326,N_12238);
xnor U12593 (N_12593,N_12285,N_12261);
nand U12594 (N_12594,N_12371,N_12395);
xor U12595 (N_12595,N_12383,N_12249);
xnor U12596 (N_12596,N_12241,N_12229);
and U12597 (N_12597,N_12243,N_12371);
xnor U12598 (N_12598,N_12307,N_12243);
and U12599 (N_12599,N_12310,N_12354);
xnor U12600 (N_12600,N_12468,N_12453);
nand U12601 (N_12601,N_12461,N_12558);
xnor U12602 (N_12602,N_12596,N_12538);
nand U12603 (N_12603,N_12526,N_12430);
or U12604 (N_12604,N_12496,N_12583);
or U12605 (N_12605,N_12597,N_12432);
nor U12606 (N_12606,N_12582,N_12549);
and U12607 (N_12607,N_12515,N_12463);
or U12608 (N_12608,N_12564,N_12545);
nand U12609 (N_12609,N_12493,N_12537);
nor U12610 (N_12610,N_12444,N_12551);
or U12611 (N_12611,N_12404,N_12428);
and U12612 (N_12612,N_12403,N_12501);
nor U12613 (N_12613,N_12525,N_12556);
and U12614 (N_12614,N_12504,N_12502);
nor U12615 (N_12615,N_12443,N_12530);
nand U12616 (N_12616,N_12512,N_12497);
and U12617 (N_12617,N_12466,N_12449);
nand U12618 (N_12618,N_12535,N_12481);
xor U12619 (N_12619,N_12578,N_12547);
or U12620 (N_12620,N_12407,N_12567);
nor U12621 (N_12621,N_12450,N_12479);
nand U12622 (N_12622,N_12555,N_12541);
or U12623 (N_12623,N_12577,N_12536);
or U12624 (N_12624,N_12492,N_12474);
xnor U12625 (N_12625,N_12565,N_12445);
xnor U12626 (N_12626,N_12495,N_12516);
or U12627 (N_12627,N_12417,N_12506);
or U12628 (N_12628,N_12408,N_12429);
nor U12629 (N_12629,N_12451,N_12457);
xor U12630 (N_12630,N_12410,N_12472);
nand U12631 (N_12631,N_12452,N_12476);
nand U12632 (N_12632,N_12589,N_12586);
and U12633 (N_12633,N_12469,N_12503);
xnor U12634 (N_12634,N_12458,N_12478);
nand U12635 (N_12635,N_12522,N_12459);
xnor U12636 (N_12636,N_12579,N_12509);
nand U12637 (N_12637,N_12462,N_12592);
nor U12638 (N_12638,N_12447,N_12553);
nand U12639 (N_12639,N_12508,N_12507);
xor U12640 (N_12640,N_12548,N_12499);
nand U12641 (N_12641,N_12409,N_12500);
xnor U12642 (N_12642,N_12483,N_12464);
nand U12643 (N_12643,N_12573,N_12411);
and U12644 (N_12644,N_12414,N_12405);
xor U12645 (N_12645,N_12470,N_12568);
and U12646 (N_12646,N_12595,N_12560);
and U12647 (N_12647,N_12524,N_12446);
nor U12648 (N_12648,N_12570,N_12510);
xnor U12649 (N_12649,N_12585,N_12511);
xor U12650 (N_12650,N_12591,N_12415);
and U12651 (N_12651,N_12563,N_12491);
xnor U12652 (N_12652,N_12482,N_12521);
xor U12653 (N_12653,N_12598,N_12437);
nand U12654 (N_12654,N_12566,N_12574);
and U12655 (N_12655,N_12486,N_12471);
and U12656 (N_12656,N_12599,N_12529);
xnor U12657 (N_12657,N_12534,N_12473);
xor U12658 (N_12658,N_12532,N_12520);
or U12659 (N_12659,N_12571,N_12422);
or U12660 (N_12660,N_12434,N_12456);
xor U12661 (N_12661,N_12413,N_12581);
nand U12662 (N_12662,N_12528,N_12518);
xor U12663 (N_12663,N_12490,N_12523);
or U12664 (N_12664,N_12552,N_12401);
or U12665 (N_12665,N_12477,N_12416);
and U12666 (N_12666,N_12489,N_12440);
nor U12667 (N_12667,N_12484,N_12554);
nor U12668 (N_12668,N_12433,N_12519);
nor U12669 (N_12669,N_12546,N_12587);
nand U12670 (N_12670,N_12527,N_12562);
nor U12671 (N_12671,N_12543,N_12455);
or U12672 (N_12672,N_12427,N_12424);
or U12673 (N_12673,N_12423,N_12425);
or U12674 (N_12674,N_12533,N_12494);
xnor U12675 (N_12675,N_12419,N_12561);
nand U12676 (N_12676,N_12448,N_12465);
nor U12677 (N_12677,N_12406,N_12505);
or U12678 (N_12678,N_12435,N_12485);
nand U12679 (N_12679,N_12498,N_12487);
and U12680 (N_12680,N_12420,N_12531);
or U12681 (N_12681,N_12580,N_12569);
or U12682 (N_12682,N_12439,N_12593);
or U12683 (N_12683,N_12576,N_12544);
or U12684 (N_12684,N_12426,N_12514);
or U12685 (N_12685,N_12418,N_12588);
nor U12686 (N_12686,N_12488,N_12557);
and U12687 (N_12687,N_12542,N_12480);
nor U12688 (N_12688,N_12559,N_12475);
and U12689 (N_12689,N_12402,N_12421);
and U12690 (N_12690,N_12400,N_12441);
nor U12691 (N_12691,N_12572,N_12436);
or U12692 (N_12692,N_12539,N_12517);
nor U12693 (N_12693,N_12594,N_12513);
or U12694 (N_12694,N_12584,N_12412);
or U12695 (N_12695,N_12550,N_12460);
and U12696 (N_12696,N_12467,N_12438);
xnor U12697 (N_12697,N_12590,N_12575);
xnor U12698 (N_12698,N_12540,N_12431);
nor U12699 (N_12699,N_12454,N_12442);
and U12700 (N_12700,N_12494,N_12532);
nor U12701 (N_12701,N_12478,N_12454);
nand U12702 (N_12702,N_12566,N_12485);
xor U12703 (N_12703,N_12499,N_12549);
nand U12704 (N_12704,N_12445,N_12465);
xor U12705 (N_12705,N_12503,N_12506);
nor U12706 (N_12706,N_12443,N_12420);
and U12707 (N_12707,N_12539,N_12478);
and U12708 (N_12708,N_12433,N_12498);
nor U12709 (N_12709,N_12483,N_12541);
and U12710 (N_12710,N_12449,N_12432);
xnor U12711 (N_12711,N_12448,N_12470);
xor U12712 (N_12712,N_12525,N_12581);
xnor U12713 (N_12713,N_12565,N_12430);
or U12714 (N_12714,N_12578,N_12590);
nand U12715 (N_12715,N_12589,N_12504);
and U12716 (N_12716,N_12545,N_12412);
nor U12717 (N_12717,N_12521,N_12513);
and U12718 (N_12718,N_12482,N_12552);
and U12719 (N_12719,N_12475,N_12440);
xnor U12720 (N_12720,N_12419,N_12569);
nor U12721 (N_12721,N_12549,N_12459);
xnor U12722 (N_12722,N_12557,N_12505);
nand U12723 (N_12723,N_12530,N_12418);
or U12724 (N_12724,N_12443,N_12497);
and U12725 (N_12725,N_12458,N_12509);
and U12726 (N_12726,N_12474,N_12513);
xnor U12727 (N_12727,N_12508,N_12425);
and U12728 (N_12728,N_12497,N_12475);
xnor U12729 (N_12729,N_12419,N_12542);
nor U12730 (N_12730,N_12575,N_12466);
and U12731 (N_12731,N_12417,N_12412);
nand U12732 (N_12732,N_12496,N_12406);
nand U12733 (N_12733,N_12558,N_12487);
or U12734 (N_12734,N_12595,N_12523);
and U12735 (N_12735,N_12405,N_12579);
or U12736 (N_12736,N_12420,N_12542);
or U12737 (N_12737,N_12567,N_12467);
nor U12738 (N_12738,N_12415,N_12501);
nand U12739 (N_12739,N_12561,N_12580);
and U12740 (N_12740,N_12445,N_12492);
and U12741 (N_12741,N_12556,N_12540);
xnor U12742 (N_12742,N_12586,N_12595);
xnor U12743 (N_12743,N_12492,N_12461);
or U12744 (N_12744,N_12438,N_12472);
and U12745 (N_12745,N_12503,N_12579);
nand U12746 (N_12746,N_12482,N_12484);
xor U12747 (N_12747,N_12528,N_12555);
xnor U12748 (N_12748,N_12559,N_12513);
nand U12749 (N_12749,N_12442,N_12465);
and U12750 (N_12750,N_12564,N_12551);
nand U12751 (N_12751,N_12431,N_12415);
and U12752 (N_12752,N_12582,N_12407);
xnor U12753 (N_12753,N_12542,N_12535);
nor U12754 (N_12754,N_12464,N_12540);
and U12755 (N_12755,N_12474,N_12452);
nor U12756 (N_12756,N_12479,N_12437);
and U12757 (N_12757,N_12581,N_12418);
nor U12758 (N_12758,N_12499,N_12518);
or U12759 (N_12759,N_12592,N_12428);
xnor U12760 (N_12760,N_12400,N_12531);
nand U12761 (N_12761,N_12459,N_12463);
or U12762 (N_12762,N_12470,N_12579);
and U12763 (N_12763,N_12442,N_12500);
and U12764 (N_12764,N_12590,N_12496);
or U12765 (N_12765,N_12478,N_12532);
nor U12766 (N_12766,N_12510,N_12509);
xor U12767 (N_12767,N_12483,N_12517);
or U12768 (N_12768,N_12404,N_12505);
nand U12769 (N_12769,N_12493,N_12428);
xor U12770 (N_12770,N_12550,N_12400);
and U12771 (N_12771,N_12448,N_12509);
xor U12772 (N_12772,N_12536,N_12504);
nand U12773 (N_12773,N_12499,N_12473);
xnor U12774 (N_12774,N_12499,N_12412);
or U12775 (N_12775,N_12405,N_12527);
nand U12776 (N_12776,N_12470,N_12578);
and U12777 (N_12777,N_12514,N_12533);
and U12778 (N_12778,N_12577,N_12496);
or U12779 (N_12779,N_12586,N_12501);
xnor U12780 (N_12780,N_12461,N_12596);
nand U12781 (N_12781,N_12568,N_12594);
and U12782 (N_12782,N_12598,N_12583);
or U12783 (N_12783,N_12509,N_12524);
or U12784 (N_12784,N_12488,N_12562);
xnor U12785 (N_12785,N_12589,N_12447);
xor U12786 (N_12786,N_12418,N_12438);
nor U12787 (N_12787,N_12560,N_12588);
and U12788 (N_12788,N_12562,N_12478);
or U12789 (N_12789,N_12521,N_12504);
xnor U12790 (N_12790,N_12412,N_12420);
nor U12791 (N_12791,N_12590,N_12523);
nand U12792 (N_12792,N_12575,N_12465);
xor U12793 (N_12793,N_12464,N_12446);
and U12794 (N_12794,N_12568,N_12496);
xnor U12795 (N_12795,N_12539,N_12491);
or U12796 (N_12796,N_12573,N_12574);
nor U12797 (N_12797,N_12552,N_12551);
and U12798 (N_12798,N_12466,N_12558);
or U12799 (N_12799,N_12453,N_12560);
nor U12800 (N_12800,N_12680,N_12642);
xor U12801 (N_12801,N_12673,N_12745);
nor U12802 (N_12802,N_12782,N_12754);
and U12803 (N_12803,N_12726,N_12601);
or U12804 (N_12804,N_12794,N_12689);
or U12805 (N_12805,N_12693,N_12767);
nor U12806 (N_12806,N_12663,N_12780);
or U12807 (N_12807,N_12790,N_12609);
xnor U12808 (N_12808,N_12773,N_12694);
nor U12809 (N_12809,N_12686,N_12799);
nand U12810 (N_12810,N_12775,N_12644);
nand U12811 (N_12811,N_12727,N_12721);
nor U12812 (N_12812,N_12662,N_12690);
xor U12813 (N_12813,N_12743,N_12651);
nor U12814 (N_12814,N_12655,N_12765);
nor U12815 (N_12815,N_12738,N_12714);
nor U12816 (N_12816,N_12712,N_12633);
and U12817 (N_12817,N_12755,N_12634);
or U12818 (N_12818,N_12747,N_12795);
xnor U12819 (N_12819,N_12730,N_12623);
or U12820 (N_12820,N_12778,N_12719);
xnor U12821 (N_12821,N_12716,N_12798);
xor U12822 (N_12822,N_12613,N_12620);
or U12823 (N_12823,N_12762,N_12626);
nand U12824 (N_12824,N_12611,N_12704);
nand U12825 (N_12825,N_12783,N_12621);
xnor U12826 (N_12826,N_12768,N_12698);
xnor U12827 (N_12827,N_12707,N_12641);
or U12828 (N_12828,N_12682,N_12701);
and U12829 (N_12829,N_12606,N_12696);
nand U12830 (N_12830,N_12630,N_12725);
nor U12831 (N_12831,N_12756,N_12757);
xnor U12832 (N_12832,N_12687,N_12793);
nor U12833 (N_12833,N_12771,N_12784);
nand U12834 (N_12834,N_12739,N_12785);
nand U12835 (N_12835,N_12781,N_12617);
and U12836 (N_12836,N_12792,N_12615);
nand U12837 (N_12837,N_12670,N_12728);
and U12838 (N_12838,N_12618,N_12643);
nor U12839 (N_12839,N_12700,N_12763);
nor U12840 (N_12840,N_12632,N_12607);
nand U12841 (N_12841,N_12668,N_12647);
and U12842 (N_12842,N_12779,N_12628);
or U12843 (N_12843,N_12675,N_12759);
nand U12844 (N_12844,N_12665,N_12603);
xnor U12845 (N_12845,N_12761,N_12608);
or U12846 (N_12846,N_12602,N_12629);
nor U12847 (N_12847,N_12695,N_12681);
and U12848 (N_12848,N_12614,N_12666);
or U12849 (N_12849,N_12637,N_12791);
or U12850 (N_12850,N_12660,N_12731);
and U12851 (N_12851,N_12657,N_12656);
xor U12852 (N_12852,N_12669,N_12764);
and U12853 (N_12853,N_12649,N_12683);
and U12854 (N_12854,N_12729,N_12766);
and U12855 (N_12855,N_12679,N_12604);
xor U12856 (N_12856,N_12708,N_12751);
or U12857 (N_12857,N_12646,N_12658);
xor U12858 (N_12858,N_12744,N_12688);
nor U12859 (N_12859,N_12749,N_12638);
nor U12860 (N_12860,N_12684,N_12760);
nor U12861 (N_12861,N_12741,N_12624);
or U12862 (N_12862,N_12640,N_12667);
and U12863 (N_12863,N_12713,N_12718);
xor U12864 (N_12864,N_12625,N_12769);
nand U12865 (N_12865,N_12652,N_12786);
nor U12866 (N_12866,N_12742,N_12612);
and U12867 (N_12867,N_12692,N_12664);
or U12868 (N_12868,N_12674,N_12705);
nand U12869 (N_12869,N_12723,N_12672);
or U12870 (N_12870,N_12702,N_12631);
xor U12871 (N_12871,N_12699,N_12736);
xor U12872 (N_12872,N_12671,N_12619);
nor U12873 (N_12873,N_12788,N_12645);
and U12874 (N_12874,N_12709,N_12627);
and U12875 (N_12875,N_12737,N_12648);
nand U12876 (N_12876,N_12770,N_12636);
nor U12877 (N_12877,N_12616,N_12722);
xnor U12878 (N_12878,N_12772,N_12639);
and U12879 (N_12879,N_12750,N_12740);
nand U12880 (N_12880,N_12691,N_12676);
and U12881 (N_12881,N_12789,N_12605);
or U12882 (N_12882,N_12635,N_12610);
xor U12883 (N_12883,N_12720,N_12733);
nand U12884 (N_12884,N_12703,N_12734);
or U12885 (N_12885,N_12732,N_12774);
nand U12886 (N_12886,N_12653,N_12661);
nor U12887 (N_12887,N_12735,N_12753);
xnor U12888 (N_12888,N_12717,N_12710);
or U12889 (N_12889,N_12697,N_12711);
nor U12890 (N_12890,N_12650,N_12622);
or U12891 (N_12891,N_12776,N_12715);
and U12892 (N_12892,N_12654,N_12787);
xor U12893 (N_12893,N_12659,N_12678);
and U12894 (N_12894,N_12748,N_12797);
xor U12895 (N_12895,N_12746,N_12758);
or U12896 (N_12896,N_12685,N_12777);
nor U12897 (N_12897,N_12796,N_12724);
or U12898 (N_12898,N_12677,N_12706);
xnor U12899 (N_12899,N_12752,N_12600);
xnor U12900 (N_12900,N_12608,N_12783);
nand U12901 (N_12901,N_12683,N_12645);
nand U12902 (N_12902,N_12717,N_12769);
and U12903 (N_12903,N_12706,N_12671);
nor U12904 (N_12904,N_12651,N_12791);
or U12905 (N_12905,N_12609,N_12793);
nor U12906 (N_12906,N_12639,N_12775);
xor U12907 (N_12907,N_12766,N_12705);
or U12908 (N_12908,N_12754,N_12720);
or U12909 (N_12909,N_12608,N_12726);
nor U12910 (N_12910,N_12684,N_12731);
nand U12911 (N_12911,N_12749,N_12697);
nand U12912 (N_12912,N_12694,N_12607);
nand U12913 (N_12913,N_12662,N_12615);
and U12914 (N_12914,N_12693,N_12702);
and U12915 (N_12915,N_12677,N_12756);
and U12916 (N_12916,N_12732,N_12747);
nand U12917 (N_12917,N_12637,N_12670);
or U12918 (N_12918,N_12659,N_12799);
xnor U12919 (N_12919,N_12661,N_12649);
nand U12920 (N_12920,N_12733,N_12782);
and U12921 (N_12921,N_12787,N_12658);
nand U12922 (N_12922,N_12609,N_12717);
and U12923 (N_12923,N_12738,N_12637);
xor U12924 (N_12924,N_12668,N_12672);
xnor U12925 (N_12925,N_12642,N_12666);
nor U12926 (N_12926,N_12706,N_12661);
and U12927 (N_12927,N_12745,N_12773);
and U12928 (N_12928,N_12677,N_12763);
nand U12929 (N_12929,N_12661,N_12681);
or U12930 (N_12930,N_12797,N_12745);
or U12931 (N_12931,N_12725,N_12723);
or U12932 (N_12932,N_12735,N_12769);
nand U12933 (N_12933,N_12799,N_12721);
or U12934 (N_12934,N_12641,N_12797);
nor U12935 (N_12935,N_12714,N_12730);
or U12936 (N_12936,N_12687,N_12702);
and U12937 (N_12937,N_12742,N_12672);
nand U12938 (N_12938,N_12748,N_12738);
and U12939 (N_12939,N_12765,N_12790);
nand U12940 (N_12940,N_12724,N_12641);
xor U12941 (N_12941,N_12601,N_12710);
xnor U12942 (N_12942,N_12762,N_12761);
nor U12943 (N_12943,N_12736,N_12660);
nor U12944 (N_12944,N_12774,N_12636);
xor U12945 (N_12945,N_12610,N_12676);
xor U12946 (N_12946,N_12657,N_12742);
nor U12947 (N_12947,N_12769,N_12796);
nand U12948 (N_12948,N_12657,N_12606);
xor U12949 (N_12949,N_12769,N_12606);
and U12950 (N_12950,N_12622,N_12797);
nor U12951 (N_12951,N_12688,N_12726);
nand U12952 (N_12952,N_12663,N_12729);
nor U12953 (N_12953,N_12782,N_12659);
nand U12954 (N_12954,N_12786,N_12746);
xnor U12955 (N_12955,N_12616,N_12602);
or U12956 (N_12956,N_12620,N_12732);
xnor U12957 (N_12957,N_12681,N_12685);
nand U12958 (N_12958,N_12649,N_12762);
xor U12959 (N_12959,N_12689,N_12617);
nor U12960 (N_12960,N_12617,N_12676);
nand U12961 (N_12961,N_12782,N_12661);
nor U12962 (N_12962,N_12733,N_12763);
and U12963 (N_12963,N_12649,N_12687);
and U12964 (N_12964,N_12756,N_12682);
or U12965 (N_12965,N_12683,N_12616);
nor U12966 (N_12966,N_12738,N_12745);
or U12967 (N_12967,N_12700,N_12676);
or U12968 (N_12968,N_12722,N_12665);
or U12969 (N_12969,N_12794,N_12706);
and U12970 (N_12970,N_12674,N_12665);
nor U12971 (N_12971,N_12766,N_12776);
xor U12972 (N_12972,N_12781,N_12620);
nand U12973 (N_12973,N_12626,N_12708);
nand U12974 (N_12974,N_12723,N_12757);
or U12975 (N_12975,N_12748,N_12641);
or U12976 (N_12976,N_12699,N_12693);
and U12977 (N_12977,N_12649,N_12711);
nor U12978 (N_12978,N_12600,N_12734);
nor U12979 (N_12979,N_12657,N_12766);
and U12980 (N_12980,N_12712,N_12693);
and U12981 (N_12981,N_12768,N_12630);
or U12982 (N_12982,N_12764,N_12729);
and U12983 (N_12983,N_12644,N_12625);
xor U12984 (N_12984,N_12695,N_12757);
or U12985 (N_12985,N_12646,N_12744);
xnor U12986 (N_12986,N_12746,N_12662);
or U12987 (N_12987,N_12620,N_12698);
xor U12988 (N_12988,N_12690,N_12790);
xor U12989 (N_12989,N_12765,N_12696);
xor U12990 (N_12990,N_12663,N_12615);
nor U12991 (N_12991,N_12734,N_12791);
nand U12992 (N_12992,N_12639,N_12793);
or U12993 (N_12993,N_12784,N_12711);
xnor U12994 (N_12994,N_12676,N_12694);
and U12995 (N_12995,N_12737,N_12644);
or U12996 (N_12996,N_12789,N_12689);
nor U12997 (N_12997,N_12700,N_12654);
xor U12998 (N_12998,N_12701,N_12629);
and U12999 (N_12999,N_12757,N_12753);
xor U13000 (N_13000,N_12884,N_12926);
nand U13001 (N_13001,N_12937,N_12857);
xnor U13002 (N_13002,N_12994,N_12940);
xor U13003 (N_13003,N_12893,N_12837);
or U13004 (N_13004,N_12904,N_12887);
and U13005 (N_13005,N_12895,N_12865);
or U13006 (N_13006,N_12869,N_12906);
nand U13007 (N_13007,N_12945,N_12978);
and U13008 (N_13008,N_12800,N_12802);
nor U13009 (N_13009,N_12839,N_12901);
or U13010 (N_13010,N_12883,N_12987);
nor U13011 (N_13011,N_12949,N_12854);
xnor U13012 (N_13012,N_12976,N_12917);
nor U13013 (N_13013,N_12806,N_12850);
and U13014 (N_13014,N_12820,N_12822);
xor U13015 (N_13015,N_12810,N_12996);
or U13016 (N_13016,N_12928,N_12927);
or U13017 (N_13017,N_12871,N_12891);
xnor U13018 (N_13018,N_12860,N_12910);
or U13019 (N_13019,N_12878,N_12918);
or U13020 (N_13020,N_12916,N_12923);
and U13021 (N_13021,N_12914,N_12943);
xnor U13022 (N_13022,N_12919,N_12861);
nand U13023 (N_13023,N_12823,N_12817);
nor U13024 (N_13024,N_12954,N_12840);
nand U13025 (N_13025,N_12855,N_12858);
nand U13026 (N_13026,N_12847,N_12859);
xor U13027 (N_13027,N_12986,N_12947);
nand U13028 (N_13028,N_12932,N_12983);
and U13029 (N_13029,N_12842,N_12920);
or U13030 (N_13030,N_12812,N_12899);
nor U13031 (N_13031,N_12974,N_12845);
nor U13032 (N_13032,N_12818,N_12873);
xnor U13033 (N_13033,N_12921,N_12813);
or U13034 (N_13034,N_12912,N_12801);
xor U13035 (N_13035,N_12896,N_12825);
and U13036 (N_13036,N_12993,N_12991);
nand U13037 (N_13037,N_12881,N_12867);
nor U13038 (N_13038,N_12997,N_12956);
xnor U13039 (N_13039,N_12944,N_12852);
or U13040 (N_13040,N_12841,N_12853);
xor U13041 (N_13041,N_12815,N_12984);
nor U13042 (N_13042,N_12963,N_12948);
or U13043 (N_13043,N_12805,N_12870);
nand U13044 (N_13044,N_12811,N_12951);
nor U13045 (N_13045,N_12998,N_12875);
and U13046 (N_13046,N_12879,N_12888);
or U13047 (N_13047,N_12808,N_12957);
nor U13048 (N_13048,N_12941,N_12832);
xnor U13049 (N_13049,N_12925,N_12961);
or U13050 (N_13050,N_12897,N_12864);
or U13051 (N_13051,N_12868,N_12866);
nand U13052 (N_13052,N_12973,N_12824);
nand U13053 (N_13053,N_12826,N_12911);
xnor U13054 (N_13054,N_12863,N_12889);
or U13055 (N_13055,N_12851,N_12989);
or U13056 (N_13056,N_12969,N_12836);
nor U13057 (N_13057,N_12846,N_12913);
nand U13058 (N_13058,N_12939,N_12971);
nor U13059 (N_13059,N_12946,N_12807);
nor U13060 (N_13060,N_12999,N_12894);
xnor U13061 (N_13061,N_12804,N_12834);
or U13062 (N_13062,N_12882,N_12890);
and U13063 (N_13063,N_12975,N_12819);
nand U13064 (N_13064,N_12816,N_12924);
nand U13065 (N_13065,N_12843,N_12874);
xor U13066 (N_13066,N_12830,N_12835);
nand U13067 (N_13067,N_12872,N_12814);
or U13068 (N_13068,N_12905,N_12966);
nand U13069 (N_13069,N_12935,N_12931);
nor U13070 (N_13070,N_12990,N_12833);
nand U13071 (N_13071,N_12995,N_12915);
xor U13072 (N_13072,N_12933,N_12936);
nand U13073 (N_13073,N_12964,N_12955);
or U13074 (N_13074,N_12962,N_12900);
nand U13075 (N_13075,N_12992,N_12907);
nor U13076 (N_13076,N_12977,N_12982);
and U13077 (N_13077,N_12838,N_12965);
xnor U13078 (N_13078,N_12979,N_12981);
xnor U13079 (N_13079,N_12908,N_12953);
and U13080 (N_13080,N_12862,N_12828);
nor U13081 (N_13081,N_12960,N_12934);
xor U13082 (N_13082,N_12929,N_12950);
or U13083 (N_13083,N_12967,N_12980);
nand U13084 (N_13084,N_12988,N_12886);
nor U13085 (N_13085,N_12877,N_12930);
xnor U13086 (N_13086,N_12902,N_12809);
xnor U13087 (N_13087,N_12903,N_12880);
nand U13088 (N_13088,N_12959,N_12909);
xnor U13089 (N_13089,N_12803,N_12844);
nor U13090 (N_13090,N_12972,N_12968);
nand U13091 (N_13091,N_12876,N_12827);
nand U13092 (N_13092,N_12970,N_12821);
nor U13093 (N_13093,N_12942,N_12958);
nor U13094 (N_13094,N_12829,N_12848);
and U13095 (N_13095,N_12856,N_12849);
nand U13096 (N_13096,N_12938,N_12892);
xnor U13097 (N_13097,N_12831,N_12898);
and U13098 (N_13098,N_12885,N_12985);
xor U13099 (N_13099,N_12952,N_12922);
xnor U13100 (N_13100,N_12871,N_12813);
nand U13101 (N_13101,N_12811,N_12983);
nand U13102 (N_13102,N_12901,N_12988);
xnor U13103 (N_13103,N_12858,N_12911);
nor U13104 (N_13104,N_12859,N_12912);
nor U13105 (N_13105,N_12807,N_12886);
and U13106 (N_13106,N_12823,N_12859);
xnor U13107 (N_13107,N_12861,N_12876);
xor U13108 (N_13108,N_12979,N_12956);
xor U13109 (N_13109,N_12992,N_12931);
or U13110 (N_13110,N_12861,N_12986);
nand U13111 (N_13111,N_12911,N_12811);
or U13112 (N_13112,N_12913,N_12895);
or U13113 (N_13113,N_12812,N_12836);
xnor U13114 (N_13114,N_12985,N_12971);
nand U13115 (N_13115,N_12884,N_12818);
xnor U13116 (N_13116,N_12820,N_12861);
xnor U13117 (N_13117,N_12839,N_12949);
nand U13118 (N_13118,N_12878,N_12902);
and U13119 (N_13119,N_12941,N_12883);
or U13120 (N_13120,N_12859,N_12955);
or U13121 (N_13121,N_12920,N_12907);
xor U13122 (N_13122,N_12989,N_12921);
nor U13123 (N_13123,N_12871,N_12988);
xor U13124 (N_13124,N_12820,N_12832);
xor U13125 (N_13125,N_12916,N_12898);
and U13126 (N_13126,N_12989,N_12850);
xor U13127 (N_13127,N_12822,N_12911);
nand U13128 (N_13128,N_12885,N_12801);
nor U13129 (N_13129,N_12899,N_12896);
or U13130 (N_13130,N_12962,N_12857);
nand U13131 (N_13131,N_12993,N_12804);
and U13132 (N_13132,N_12965,N_12935);
xnor U13133 (N_13133,N_12826,N_12858);
nand U13134 (N_13134,N_12903,N_12955);
xnor U13135 (N_13135,N_12823,N_12950);
or U13136 (N_13136,N_12832,N_12852);
xnor U13137 (N_13137,N_12883,N_12865);
xnor U13138 (N_13138,N_12923,N_12866);
or U13139 (N_13139,N_12856,N_12829);
nand U13140 (N_13140,N_12804,N_12816);
nor U13141 (N_13141,N_12811,N_12990);
xor U13142 (N_13142,N_12818,N_12855);
and U13143 (N_13143,N_12878,N_12976);
or U13144 (N_13144,N_12881,N_12909);
nor U13145 (N_13145,N_12964,N_12875);
and U13146 (N_13146,N_12861,N_12854);
nand U13147 (N_13147,N_12921,N_12857);
xnor U13148 (N_13148,N_12930,N_12845);
xnor U13149 (N_13149,N_12839,N_12913);
nand U13150 (N_13150,N_12914,N_12920);
or U13151 (N_13151,N_12977,N_12946);
and U13152 (N_13152,N_12851,N_12987);
xor U13153 (N_13153,N_12954,N_12924);
xnor U13154 (N_13154,N_12800,N_12989);
nand U13155 (N_13155,N_12987,N_12893);
nor U13156 (N_13156,N_12945,N_12859);
nor U13157 (N_13157,N_12956,N_12951);
nor U13158 (N_13158,N_12916,N_12873);
nand U13159 (N_13159,N_12827,N_12961);
or U13160 (N_13160,N_12844,N_12839);
and U13161 (N_13161,N_12929,N_12985);
and U13162 (N_13162,N_12890,N_12881);
nand U13163 (N_13163,N_12923,N_12817);
nand U13164 (N_13164,N_12877,N_12974);
or U13165 (N_13165,N_12838,N_12950);
or U13166 (N_13166,N_12908,N_12961);
nand U13167 (N_13167,N_12842,N_12869);
and U13168 (N_13168,N_12969,N_12990);
xnor U13169 (N_13169,N_12835,N_12806);
nor U13170 (N_13170,N_12944,N_12890);
nor U13171 (N_13171,N_12986,N_12829);
and U13172 (N_13172,N_12972,N_12941);
or U13173 (N_13173,N_12950,N_12931);
nor U13174 (N_13174,N_12933,N_12988);
xor U13175 (N_13175,N_12940,N_12942);
xor U13176 (N_13176,N_12809,N_12951);
or U13177 (N_13177,N_12833,N_12936);
xnor U13178 (N_13178,N_12894,N_12856);
and U13179 (N_13179,N_12977,N_12965);
nor U13180 (N_13180,N_12986,N_12815);
or U13181 (N_13181,N_12823,N_12911);
or U13182 (N_13182,N_12813,N_12828);
xor U13183 (N_13183,N_12933,N_12991);
and U13184 (N_13184,N_12973,N_12970);
nand U13185 (N_13185,N_12926,N_12975);
and U13186 (N_13186,N_12847,N_12828);
nor U13187 (N_13187,N_12804,N_12941);
and U13188 (N_13188,N_12819,N_12874);
or U13189 (N_13189,N_12945,N_12826);
nand U13190 (N_13190,N_12947,N_12911);
or U13191 (N_13191,N_12819,N_12977);
and U13192 (N_13192,N_12810,N_12964);
nor U13193 (N_13193,N_12847,N_12975);
xnor U13194 (N_13194,N_12985,N_12899);
xor U13195 (N_13195,N_12896,N_12960);
or U13196 (N_13196,N_12924,N_12911);
or U13197 (N_13197,N_12923,N_12960);
and U13198 (N_13198,N_12814,N_12904);
nand U13199 (N_13199,N_12945,N_12909);
nor U13200 (N_13200,N_13155,N_13063);
or U13201 (N_13201,N_13187,N_13103);
or U13202 (N_13202,N_13127,N_13178);
nand U13203 (N_13203,N_13096,N_13046);
nor U13204 (N_13204,N_13016,N_13060);
nand U13205 (N_13205,N_13176,N_13186);
or U13206 (N_13206,N_13109,N_13115);
and U13207 (N_13207,N_13040,N_13168);
nand U13208 (N_13208,N_13067,N_13164);
nand U13209 (N_13209,N_13198,N_13089);
and U13210 (N_13210,N_13087,N_13024);
nor U13211 (N_13211,N_13041,N_13043);
and U13212 (N_13212,N_13083,N_13056);
nor U13213 (N_13213,N_13035,N_13153);
or U13214 (N_13214,N_13062,N_13125);
or U13215 (N_13215,N_13090,N_13112);
or U13216 (N_13216,N_13031,N_13033);
and U13217 (N_13217,N_13057,N_13172);
or U13218 (N_13218,N_13019,N_13078);
nor U13219 (N_13219,N_13054,N_13114);
nor U13220 (N_13220,N_13086,N_13123);
nor U13221 (N_13221,N_13138,N_13095);
nand U13222 (N_13222,N_13038,N_13120);
nor U13223 (N_13223,N_13161,N_13082);
nor U13224 (N_13224,N_13084,N_13199);
xnor U13225 (N_13225,N_13165,N_13130);
or U13226 (N_13226,N_13166,N_13000);
nor U13227 (N_13227,N_13070,N_13014);
nand U13228 (N_13228,N_13188,N_13009);
xnor U13229 (N_13229,N_13194,N_13018);
nand U13230 (N_13230,N_13162,N_13073);
or U13231 (N_13231,N_13049,N_13001);
and U13232 (N_13232,N_13119,N_13075);
nor U13233 (N_13233,N_13036,N_13011);
or U13234 (N_13234,N_13048,N_13159);
and U13235 (N_13235,N_13128,N_13197);
or U13236 (N_13236,N_13071,N_13160);
xnor U13237 (N_13237,N_13097,N_13034);
nor U13238 (N_13238,N_13196,N_13189);
nand U13239 (N_13239,N_13157,N_13131);
xor U13240 (N_13240,N_13021,N_13100);
or U13241 (N_13241,N_13044,N_13163);
nor U13242 (N_13242,N_13080,N_13136);
xor U13243 (N_13243,N_13173,N_13025);
xor U13244 (N_13244,N_13012,N_13190);
and U13245 (N_13245,N_13055,N_13066);
xnor U13246 (N_13246,N_13156,N_13051);
or U13247 (N_13247,N_13088,N_13076);
and U13248 (N_13248,N_13185,N_13013);
or U13249 (N_13249,N_13053,N_13126);
nor U13250 (N_13250,N_13068,N_13047);
nand U13251 (N_13251,N_13142,N_13171);
and U13252 (N_13252,N_13107,N_13027);
xor U13253 (N_13253,N_13004,N_13133);
nand U13254 (N_13254,N_13129,N_13079);
nor U13255 (N_13255,N_13145,N_13023);
xnor U13256 (N_13256,N_13132,N_13158);
or U13257 (N_13257,N_13069,N_13045);
and U13258 (N_13258,N_13101,N_13149);
or U13259 (N_13259,N_13144,N_13137);
or U13260 (N_13260,N_13008,N_13032);
and U13261 (N_13261,N_13140,N_13116);
nor U13262 (N_13262,N_13122,N_13192);
or U13263 (N_13263,N_13169,N_13072);
nand U13264 (N_13264,N_13118,N_13106);
nor U13265 (N_13265,N_13121,N_13177);
or U13266 (N_13266,N_13006,N_13147);
or U13267 (N_13267,N_13029,N_13028);
or U13268 (N_13268,N_13105,N_13113);
nand U13269 (N_13269,N_13065,N_13170);
or U13270 (N_13270,N_13058,N_13110);
and U13271 (N_13271,N_13030,N_13102);
xor U13272 (N_13272,N_13134,N_13050);
nor U13273 (N_13273,N_13150,N_13002);
xor U13274 (N_13274,N_13074,N_13085);
nor U13275 (N_13275,N_13026,N_13039);
and U13276 (N_13276,N_13174,N_13148);
nand U13277 (N_13277,N_13154,N_13003);
nor U13278 (N_13278,N_13146,N_13124);
nand U13279 (N_13279,N_13141,N_13052);
or U13280 (N_13280,N_13099,N_13117);
nor U13281 (N_13281,N_13017,N_13081);
nand U13282 (N_13282,N_13104,N_13010);
nor U13283 (N_13283,N_13037,N_13093);
xnor U13284 (N_13284,N_13181,N_13195);
xor U13285 (N_13285,N_13183,N_13059);
xnor U13286 (N_13286,N_13077,N_13167);
nand U13287 (N_13287,N_13061,N_13005);
xnor U13288 (N_13288,N_13175,N_13108);
xor U13289 (N_13289,N_13184,N_13015);
nor U13290 (N_13290,N_13098,N_13180);
xor U13291 (N_13291,N_13020,N_13143);
nand U13292 (N_13292,N_13193,N_13042);
nand U13293 (N_13293,N_13007,N_13135);
and U13294 (N_13294,N_13139,N_13094);
xor U13295 (N_13295,N_13064,N_13022);
nor U13296 (N_13296,N_13111,N_13191);
nor U13297 (N_13297,N_13151,N_13092);
or U13298 (N_13298,N_13152,N_13179);
and U13299 (N_13299,N_13182,N_13091);
and U13300 (N_13300,N_13025,N_13081);
nand U13301 (N_13301,N_13094,N_13087);
and U13302 (N_13302,N_13063,N_13001);
and U13303 (N_13303,N_13003,N_13192);
xnor U13304 (N_13304,N_13101,N_13181);
and U13305 (N_13305,N_13152,N_13133);
or U13306 (N_13306,N_13135,N_13011);
or U13307 (N_13307,N_13013,N_13153);
nor U13308 (N_13308,N_13053,N_13148);
and U13309 (N_13309,N_13114,N_13019);
and U13310 (N_13310,N_13159,N_13147);
or U13311 (N_13311,N_13083,N_13019);
nor U13312 (N_13312,N_13063,N_13062);
or U13313 (N_13313,N_13090,N_13075);
and U13314 (N_13314,N_13050,N_13136);
nand U13315 (N_13315,N_13162,N_13125);
or U13316 (N_13316,N_13119,N_13053);
nand U13317 (N_13317,N_13186,N_13078);
nand U13318 (N_13318,N_13191,N_13123);
nand U13319 (N_13319,N_13137,N_13054);
and U13320 (N_13320,N_13191,N_13151);
nand U13321 (N_13321,N_13003,N_13067);
nand U13322 (N_13322,N_13034,N_13031);
and U13323 (N_13323,N_13170,N_13154);
nor U13324 (N_13324,N_13027,N_13103);
xnor U13325 (N_13325,N_13171,N_13134);
nor U13326 (N_13326,N_13007,N_13171);
xor U13327 (N_13327,N_13021,N_13014);
nor U13328 (N_13328,N_13065,N_13035);
or U13329 (N_13329,N_13147,N_13183);
and U13330 (N_13330,N_13190,N_13106);
and U13331 (N_13331,N_13081,N_13072);
nor U13332 (N_13332,N_13012,N_13050);
or U13333 (N_13333,N_13173,N_13177);
nor U13334 (N_13334,N_13155,N_13057);
nor U13335 (N_13335,N_13150,N_13166);
nand U13336 (N_13336,N_13008,N_13017);
nand U13337 (N_13337,N_13141,N_13164);
and U13338 (N_13338,N_13199,N_13013);
or U13339 (N_13339,N_13013,N_13119);
nand U13340 (N_13340,N_13130,N_13005);
nand U13341 (N_13341,N_13138,N_13072);
and U13342 (N_13342,N_13136,N_13098);
xor U13343 (N_13343,N_13167,N_13034);
and U13344 (N_13344,N_13108,N_13012);
or U13345 (N_13345,N_13030,N_13156);
nand U13346 (N_13346,N_13182,N_13047);
and U13347 (N_13347,N_13073,N_13194);
nor U13348 (N_13348,N_13047,N_13008);
nand U13349 (N_13349,N_13187,N_13045);
xnor U13350 (N_13350,N_13027,N_13134);
nand U13351 (N_13351,N_13053,N_13142);
nor U13352 (N_13352,N_13100,N_13187);
nor U13353 (N_13353,N_13187,N_13197);
nor U13354 (N_13354,N_13049,N_13127);
xor U13355 (N_13355,N_13015,N_13164);
or U13356 (N_13356,N_13068,N_13169);
and U13357 (N_13357,N_13076,N_13014);
nand U13358 (N_13358,N_13100,N_13032);
nand U13359 (N_13359,N_13169,N_13041);
and U13360 (N_13360,N_13014,N_13063);
and U13361 (N_13361,N_13077,N_13123);
xor U13362 (N_13362,N_13092,N_13029);
nor U13363 (N_13363,N_13107,N_13022);
nand U13364 (N_13364,N_13094,N_13193);
and U13365 (N_13365,N_13027,N_13082);
nor U13366 (N_13366,N_13114,N_13081);
xor U13367 (N_13367,N_13049,N_13014);
or U13368 (N_13368,N_13064,N_13179);
nand U13369 (N_13369,N_13048,N_13049);
nor U13370 (N_13370,N_13007,N_13104);
xor U13371 (N_13371,N_13163,N_13111);
and U13372 (N_13372,N_13068,N_13140);
xor U13373 (N_13373,N_13195,N_13111);
xnor U13374 (N_13374,N_13032,N_13162);
or U13375 (N_13375,N_13034,N_13042);
nand U13376 (N_13376,N_13115,N_13008);
nor U13377 (N_13377,N_13100,N_13163);
xnor U13378 (N_13378,N_13132,N_13009);
nand U13379 (N_13379,N_13111,N_13030);
xor U13380 (N_13380,N_13165,N_13197);
and U13381 (N_13381,N_13114,N_13174);
or U13382 (N_13382,N_13050,N_13096);
and U13383 (N_13383,N_13152,N_13098);
nor U13384 (N_13384,N_13109,N_13052);
xnor U13385 (N_13385,N_13097,N_13179);
nand U13386 (N_13386,N_13026,N_13028);
xor U13387 (N_13387,N_13061,N_13054);
nand U13388 (N_13388,N_13063,N_13127);
nor U13389 (N_13389,N_13101,N_13029);
nand U13390 (N_13390,N_13038,N_13169);
or U13391 (N_13391,N_13192,N_13088);
nand U13392 (N_13392,N_13169,N_13015);
or U13393 (N_13393,N_13010,N_13158);
nand U13394 (N_13394,N_13116,N_13063);
nand U13395 (N_13395,N_13025,N_13146);
and U13396 (N_13396,N_13045,N_13171);
xor U13397 (N_13397,N_13008,N_13081);
and U13398 (N_13398,N_13152,N_13116);
xnor U13399 (N_13399,N_13148,N_13080);
nand U13400 (N_13400,N_13312,N_13386);
nor U13401 (N_13401,N_13376,N_13240);
nand U13402 (N_13402,N_13374,N_13215);
nand U13403 (N_13403,N_13286,N_13393);
nand U13404 (N_13404,N_13371,N_13293);
or U13405 (N_13405,N_13333,N_13235);
or U13406 (N_13406,N_13311,N_13256);
nand U13407 (N_13407,N_13261,N_13252);
xnor U13408 (N_13408,N_13216,N_13338);
or U13409 (N_13409,N_13309,N_13313);
or U13410 (N_13410,N_13296,N_13241);
nor U13411 (N_13411,N_13237,N_13272);
nand U13412 (N_13412,N_13279,N_13303);
nor U13413 (N_13413,N_13266,N_13213);
and U13414 (N_13414,N_13385,N_13399);
xnor U13415 (N_13415,N_13299,N_13326);
or U13416 (N_13416,N_13388,N_13322);
or U13417 (N_13417,N_13324,N_13221);
and U13418 (N_13418,N_13262,N_13327);
or U13419 (N_13419,N_13263,N_13288);
nand U13420 (N_13420,N_13206,N_13236);
and U13421 (N_13421,N_13225,N_13305);
nor U13422 (N_13422,N_13351,N_13378);
or U13423 (N_13423,N_13291,N_13223);
and U13424 (N_13424,N_13361,N_13227);
nor U13425 (N_13425,N_13356,N_13217);
nand U13426 (N_13426,N_13275,N_13325);
xnor U13427 (N_13427,N_13317,N_13255);
nor U13428 (N_13428,N_13392,N_13350);
or U13429 (N_13429,N_13258,N_13257);
or U13430 (N_13430,N_13287,N_13232);
nand U13431 (N_13431,N_13234,N_13273);
xnor U13432 (N_13432,N_13230,N_13364);
and U13433 (N_13433,N_13278,N_13316);
xor U13434 (N_13434,N_13251,N_13259);
nand U13435 (N_13435,N_13243,N_13253);
or U13436 (N_13436,N_13228,N_13250);
nand U13437 (N_13437,N_13211,N_13321);
or U13438 (N_13438,N_13360,N_13298);
or U13439 (N_13439,N_13348,N_13249);
and U13440 (N_13440,N_13319,N_13389);
or U13441 (N_13441,N_13233,N_13354);
and U13442 (N_13442,N_13334,N_13212);
xor U13443 (N_13443,N_13332,N_13290);
or U13444 (N_13444,N_13203,N_13379);
nand U13445 (N_13445,N_13384,N_13363);
nand U13446 (N_13446,N_13306,N_13245);
or U13447 (N_13447,N_13318,N_13294);
and U13448 (N_13448,N_13323,N_13390);
and U13449 (N_13449,N_13246,N_13274);
or U13450 (N_13450,N_13307,N_13345);
xor U13451 (N_13451,N_13229,N_13200);
xor U13452 (N_13452,N_13265,N_13289);
and U13453 (N_13453,N_13218,N_13396);
nor U13454 (N_13454,N_13283,N_13359);
nand U13455 (N_13455,N_13285,N_13397);
nor U13456 (N_13456,N_13387,N_13336);
nand U13457 (N_13457,N_13282,N_13244);
and U13458 (N_13458,N_13254,N_13207);
xor U13459 (N_13459,N_13368,N_13358);
nand U13460 (N_13460,N_13335,N_13373);
xnor U13461 (N_13461,N_13208,N_13310);
xor U13462 (N_13462,N_13284,N_13242);
xnor U13463 (N_13463,N_13281,N_13366);
nor U13464 (N_13464,N_13369,N_13268);
nand U13465 (N_13465,N_13238,N_13226);
nor U13466 (N_13466,N_13353,N_13224);
or U13467 (N_13467,N_13280,N_13301);
and U13468 (N_13468,N_13264,N_13343);
nand U13469 (N_13469,N_13300,N_13398);
nor U13470 (N_13470,N_13219,N_13346);
nand U13471 (N_13471,N_13204,N_13314);
and U13472 (N_13472,N_13362,N_13248);
or U13473 (N_13473,N_13395,N_13382);
xor U13474 (N_13474,N_13201,N_13381);
and U13475 (N_13475,N_13370,N_13367);
nand U13476 (N_13476,N_13260,N_13328);
xnor U13477 (N_13477,N_13375,N_13337);
nor U13478 (N_13478,N_13247,N_13270);
nand U13479 (N_13479,N_13357,N_13210);
nand U13480 (N_13480,N_13220,N_13341);
or U13481 (N_13481,N_13315,N_13269);
or U13482 (N_13482,N_13344,N_13271);
and U13483 (N_13483,N_13292,N_13339);
and U13484 (N_13484,N_13347,N_13365);
or U13485 (N_13485,N_13331,N_13383);
and U13486 (N_13486,N_13394,N_13372);
nor U13487 (N_13487,N_13205,N_13320);
xor U13488 (N_13488,N_13380,N_13209);
and U13489 (N_13489,N_13329,N_13276);
and U13490 (N_13490,N_13231,N_13340);
and U13491 (N_13491,N_13239,N_13349);
xnor U13492 (N_13492,N_13342,N_13267);
or U13493 (N_13493,N_13304,N_13222);
nand U13494 (N_13494,N_13295,N_13277);
and U13495 (N_13495,N_13330,N_13391);
nor U13496 (N_13496,N_13214,N_13352);
or U13497 (N_13497,N_13297,N_13355);
or U13498 (N_13498,N_13302,N_13308);
nor U13499 (N_13499,N_13202,N_13377);
nand U13500 (N_13500,N_13262,N_13205);
xor U13501 (N_13501,N_13236,N_13370);
and U13502 (N_13502,N_13396,N_13297);
or U13503 (N_13503,N_13233,N_13301);
and U13504 (N_13504,N_13222,N_13382);
nand U13505 (N_13505,N_13251,N_13345);
and U13506 (N_13506,N_13306,N_13355);
nor U13507 (N_13507,N_13209,N_13238);
nor U13508 (N_13508,N_13375,N_13204);
or U13509 (N_13509,N_13326,N_13247);
or U13510 (N_13510,N_13279,N_13334);
xor U13511 (N_13511,N_13206,N_13222);
or U13512 (N_13512,N_13359,N_13284);
nor U13513 (N_13513,N_13223,N_13297);
nor U13514 (N_13514,N_13350,N_13370);
and U13515 (N_13515,N_13217,N_13289);
nor U13516 (N_13516,N_13361,N_13295);
nor U13517 (N_13517,N_13371,N_13246);
or U13518 (N_13518,N_13267,N_13223);
nand U13519 (N_13519,N_13326,N_13390);
and U13520 (N_13520,N_13278,N_13262);
nor U13521 (N_13521,N_13359,N_13382);
or U13522 (N_13522,N_13287,N_13248);
nor U13523 (N_13523,N_13264,N_13360);
or U13524 (N_13524,N_13309,N_13299);
and U13525 (N_13525,N_13295,N_13342);
nor U13526 (N_13526,N_13364,N_13371);
nand U13527 (N_13527,N_13203,N_13243);
nor U13528 (N_13528,N_13214,N_13286);
nand U13529 (N_13529,N_13261,N_13362);
xnor U13530 (N_13530,N_13232,N_13263);
xor U13531 (N_13531,N_13288,N_13385);
or U13532 (N_13532,N_13252,N_13362);
or U13533 (N_13533,N_13313,N_13380);
nor U13534 (N_13534,N_13210,N_13330);
nand U13535 (N_13535,N_13264,N_13374);
or U13536 (N_13536,N_13269,N_13208);
and U13537 (N_13537,N_13372,N_13377);
nand U13538 (N_13538,N_13275,N_13278);
xor U13539 (N_13539,N_13245,N_13216);
nor U13540 (N_13540,N_13265,N_13332);
xnor U13541 (N_13541,N_13247,N_13310);
xnor U13542 (N_13542,N_13342,N_13261);
xor U13543 (N_13543,N_13329,N_13203);
xor U13544 (N_13544,N_13266,N_13273);
nor U13545 (N_13545,N_13213,N_13361);
nand U13546 (N_13546,N_13379,N_13303);
or U13547 (N_13547,N_13315,N_13372);
nand U13548 (N_13548,N_13348,N_13346);
or U13549 (N_13549,N_13335,N_13321);
nand U13550 (N_13550,N_13247,N_13299);
or U13551 (N_13551,N_13302,N_13394);
nor U13552 (N_13552,N_13218,N_13271);
xnor U13553 (N_13553,N_13393,N_13380);
xor U13554 (N_13554,N_13221,N_13323);
nand U13555 (N_13555,N_13228,N_13278);
nor U13556 (N_13556,N_13386,N_13381);
or U13557 (N_13557,N_13339,N_13224);
nor U13558 (N_13558,N_13326,N_13219);
and U13559 (N_13559,N_13392,N_13231);
xor U13560 (N_13560,N_13320,N_13242);
or U13561 (N_13561,N_13342,N_13304);
xor U13562 (N_13562,N_13328,N_13339);
nand U13563 (N_13563,N_13368,N_13393);
and U13564 (N_13564,N_13209,N_13328);
or U13565 (N_13565,N_13220,N_13278);
or U13566 (N_13566,N_13268,N_13229);
and U13567 (N_13567,N_13311,N_13351);
and U13568 (N_13568,N_13243,N_13364);
nand U13569 (N_13569,N_13383,N_13267);
xnor U13570 (N_13570,N_13263,N_13277);
and U13571 (N_13571,N_13250,N_13212);
nand U13572 (N_13572,N_13399,N_13214);
nand U13573 (N_13573,N_13201,N_13200);
and U13574 (N_13574,N_13369,N_13367);
nand U13575 (N_13575,N_13317,N_13284);
xor U13576 (N_13576,N_13262,N_13257);
xnor U13577 (N_13577,N_13319,N_13267);
or U13578 (N_13578,N_13397,N_13320);
nor U13579 (N_13579,N_13277,N_13353);
and U13580 (N_13580,N_13327,N_13236);
nor U13581 (N_13581,N_13372,N_13286);
or U13582 (N_13582,N_13227,N_13212);
nand U13583 (N_13583,N_13233,N_13293);
xor U13584 (N_13584,N_13268,N_13389);
nand U13585 (N_13585,N_13309,N_13371);
and U13586 (N_13586,N_13283,N_13257);
and U13587 (N_13587,N_13202,N_13281);
nand U13588 (N_13588,N_13307,N_13354);
or U13589 (N_13589,N_13356,N_13244);
nand U13590 (N_13590,N_13236,N_13376);
nand U13591 (N_13591,N_13215,N_13357);
or U13592 (N_13592,N_13227,N_13301);
and U13593 (N_13593,N_13265,N_13207);
nor U13594 (N_13594,N_13266,N_13392);
nand U13595 (N_13595,N_13290,N_13310);
and U13596 (N_13596,N_13368,N_13302);
or U13597 (N_13597,N_13231,N_13229);
and U13598 (N_13598,N_13215,N_13229);
or U13599 (N_13599,N_13211,N_13373);
or U13600 (N_13600,N_13490,N_13525);
xnor U13601 (N_13601,N_13463,N_13453);
nand U13602 (N_13602,N_13542,N_13509);
nand U13603 (N_13603,N_13593,N_13454);
xnor U13604 (N_13604,N_13414,N_13495);
nor U13605 (N_13605,N_13465,N_13592);
nor U13606 (N_13606,N_13496,N_13430);
nand U13607 (N_13607,N_13419,N_13477);
xor U13608 (N_13608,N_13591,N_13521);
or U13609 (N_13609,N_13505,N_13476);
nor U13610 (N_13610,N_13471,N_13508);
or U13611 (N_13611,N_13518,N_13451);
nor U13612 (N_13612,N_13533,N_13499);
and U13613 (N_13613,N_13551,N_13455);
xor U13614 (N_13614,N_13484,N_13578);
nand U13615 (N_13615,N_13532,N_13488);
xnor U13616 (N_13616,N_13581,N_13524);
or U13617 (N_13617,N_13552,N_13478);
xor U13618 (N_13618,N_13547,N_13522);
nand U13619 (N_13619,N_13571,N_13444);
and U13620 (N_13620,N_13489,N_13528);
or U13621 (N_13621,N_13580,N_13520);
nand U13622 (N_13622,N_13480,N_13437);
nor U13623 (N_13623,N_13565,N_13462);
xor U13624 (N_13624,N_13540,N_13497);
xor U13625 (N_13625,N_13573,N_13429);
and U13626 (N_13626,N_13426,N_13519);
nand U13627 (N_13627,N_13545,N_13410);
nor U13628 (N_13628,N_13411,N_13589);
or U13629 (N_13629,N_13594,N_13555);
xnor U13630 (N_13630,N_13510,N_13493);
xnor U13631 (N_13631,N_13539,N_13423);
or U13632 (N_13632,N_13424,N_13481);
xnor U13633 (N_13633,N_13598,N_13523);
nand U13634 (N_13634,N_13599,N_13404);
nor U13635 (N_13635,N_13527,N_13450);
or U13636 (N_13636,N_13553,N_13474);
nor U13637 (N_13637,N_13517,N_13575);
nor U13638 (N_13638,N_13473,N_13487);
xnor U13639 (N_13639,N_13469,N_13558);
and U13640 (N_13640,N_13550,N_13470);
xnor U13641 (N_13641,N_13407,N_13537);
nand U13642 (N_13642,N_13564,N_13427);
or U13643 (N_13643,N_13436,N_13452);
and U13644 (N_13644,N_13572,N_13428);
xor U13645 (N_13645,N_13443,N_13500);
nand U13646 (N_13646,N_13418,N_13595);
or U13647 (N_13647,N_13403,N_13447);
or U13648 (N_13648,N_13516,N_13590);
nand U13649 (N_13649,N_13439,N_13531);
xor U13650 (N_13650,N_13566,N_13502);
nor U13651 (N_13651,N_13467,N_13582);
nand U13652 (N_13652,N_13486,N_13538);
xnor U13653 (N_13653,N_13498,N_13422);
and U13654 (N_13654,N_13434,N_13460);
nand U13655 (N_13655,N_13507,N_13485);
and U13656 (N_13656,N_13492,N_13504);
nand U13657 (N_13657,N_13586,N_13503);
and U13658 (N_13658,N_13506,N_13468);
or U13659 (N_13659,N_13438,N_13416);
or U13660 (N_13660,N_13583,N_13431);
xor U13661 (N_13661,N_13546,N_13412);
nor U13662 (N_13662,N_13560,N_13458);
nand U13663 (N_13663,N_13570,N_13421);
nor U13664 (N_13664,N_13440,N_13466);
nand U13665 (N_13665,N_13456,N_13543);
and U13666 (N_13666,N_13442,N_13585);
nand U13667 (N_13667,N_13536,N_13475);
and U13668 (N_13668,N_13409,N_13483);
xnor U13669 (N_13669,N_13435,N_13514);
nor U13670 (N_13670,N_13515,N_13557);
nand U13671 (N_13671,N_13561,N_13491);
or U13672 (N_13672,N_13548,N_13544);
nand U13673 (N_13673,N_13568,N_13588);
xnor U13674 (N_13674,N_13464,N_13559);
or U13675 (N_13675,N_13441,N_13562);
nand U13676 (N_13676,N_13433,N_13401);
and U13677 (N_13677,N_13406,N_13529);
nor U13678 (N_13678,N_13526,N_13513);
and U13679 (N_13679,N_13494,N_13425);
nor U13680 (N_13680,N_13405,N_13549);
nand U13681 (N_13681,N_13512,N_13535);
nor U13682 (N_13682,N_13479,N_13402);
xnor U13683 (N_13683,N_13413,N_13569);
xor U13684 (N_13684,N_13556,N_13408);
nor U13685 (N_13685,N_13448,N_13511);
nand U13686 (N_13686,N_13587,N_13461);
or U13687 (N_13687,N_13459,N_13415);
or U13688 (N_13688,N_13482,N_13420);
and U13689 (N_13689,N_13596,N_13445);
nand U13690 (N_13690,N_13446,N_13501);
nor U13691 (N_13691,N_13534,N_13457);
nand U13692 (N_13692,N_13449,N_13432);
and U13693 (N_13693,N_13417,N_13597);
nor U13694 (N_13694,N_13541,N_13400);
and U13695 (N_13695,N_13574,N_13472);
nor U13696 (N_13696,N_13554,N_13563);
nor U13697 (N_13697,N_13584,N_13530);
nor U13698 (N_13698,N_13576,N_13567);
nor U13699 (N_13699,N_13579,N_13577);
xnor U13700 (N_13700,N_13556,N_13529);
and U13701 (N_13701,N_13409,N_13458);
or U13702 (N_13702,N_13556,N_13560);
and U13703 (N_13703,N_13498,N_13582);
nor U13704 (N_13704,N_13556,N_13527);
or U13705 (N_13705,N_13491,N_13419);
and U13706 (N_13706,N_13490,N_13402);
and U13707 (N_13707,N_13444,N_13577);
nor U13708 (N_13708,N_13578,N_13456);
nor U13709 (N_13709,N_13554,N_13484);
nand U13710 (N_13710,N_13456,N_13553);
xor U13711 (N_13711,N_13456,N_13486);
and U13712 (N_13712,N_13512,N_13446);
and U13713 (N_13713,N_13517,N_13484);
or U13714 (N_13714,N_13479,N_13503);
xor U13715 (N_13715,N_13416,N_13560);
or U13716 (N_13716,N_13554,N_13470);
or U13717 (N_13717,N_13515,N_13516);
or U13718 (N_13718,N_13491,N_13540);
nor U13719 (N_13719,N_13595,N_13562);
nor U13720 (N_13720,N_13571,N_13576);
or U13721 (N_13721,N_13557,N_13424);
nand U13722 (N_13722,N_13455,N_13574);
xnor U13723 (N_13723,N_13545,N_13530);
or U13724 (N_13724,N_13484,N_13560);
xor U13725 (N_13725,N_13582,N_13515);
nor U13726 (N_13726,N_13425,N_13557);
nor U13727 (N_13727,N_13521,N_13405);
nor U13728 (N_13728,N_13497,N_13449);
nor U13729 (N_13729,N_13550,N_13404);
or U13730 (N_13730,N_13479,N_13404);
xnor U13731 (N_13731,N_13585,N_13545);
nor U13732 (N_13732,N_13525,N_13518);
and U13733 (N_13733,N_13478,N_13507);
nand U13734 (N_13734,N_13572,N_13493);
xor U13735 (N_13735,N_13497,N_13567);
nand U13736 (N_13736,N_13481,N_13550);
and U13737 (N_13737,N_13526,N_13461);
or U13738 (N_13738,N_13568,N_13427);
nand U13739 (N_13739,N_13530,N_13572);
or U13740 (N_13740,N_13488,N_13596);
and U13741 (N_13741,N_13451,N_13455);
nor U13742 (N_13742,N_13534,N_13408);
nand U13743 (N_13743,N_13560,N_13489);
xnor U13744 (N_13744,N_13514,N_13412);
or U13745 (N_13745,N_13430,N_13465);
xor U13746 (N_13746,N_13457,N_13426);
or U13747 (N_13747,N_13595,N_13413);
xor U13748 (N_13748,N_13480,N_13473);
xnor U13749 (N_13749,N_13546,N_13411);
and U13750 (N_13750,N_13436,N_13450);
and U13751 (N_13751,N_13537,N_13571);
nor U13752 (N_13752,N_13530,N_13515);
nand U13753 (N_13753,N_13426,N_13565);
nor U13754 (N_13754,N_13550,N_13555);
xnor U13755 (N_13755,N_13567,N_13460);
nand U13756 (N_13756,N_13563,N_13527);
and U13757 (N_13757,N_13445,N_13567);
and U13758 (N_13758,N_13407,N_13547);
or U13759 (N_13759,N_13520,N_13431);
and U13760 (N_13760,N_13531,N_13538);
or U13761 (N_13761,N_13402,N_13404);
nand U13762 (N_13762,N_13472,N_13436);
and U13763 (N_13763,N_13449,N_13591);
xor U13764 (N_13764,N_13502,N_13422);
or U13765 (N_13765,N_13580,N_13420);
nand U13766 (N_13766,N_13585,N_13495);
nand U13767 (N_13767,N_13594,N_13447);
or U13768 (N_13768,N_13543,N_13564);
nor U13769 (N_13769,N_13412,N_13526);
xor U13770 (N_13770,N_13560,N_13434);
and U13771 (N_13771,N_13486,N_13429);
or U13772 (N_13772,N_13502,N_13426);
nand U13773 (N_13773,N_13471,N_13435);
and U13774 (N_13774,N_13492,N_13481);
nand U13775 (N_13775,N_13559,N_13513);
or U13776 (N_13776,N_13447,N_13582);
nand U13777 (N_13777,N_13581,N_13428);
or U13778 (N_13778,N_13525,N_13468);
nor U13779 (N_13779,N_13492,N_13431);
nand U13780 (N_13780,N_13424,N_13512);
xnor U13781 (N_13781,N_13554,N_13520);
or U13782 (N_13782,N_13518,N_13580);
nand U13783 (N_13783,N_13567,N_13511);
nor U13784 (N_13784,N_13586,N_13413);
and U13785 (N_13785,N_13416,N_13472);
nand U13786 (N_13786,N_13412,N_13467);
nand U13787 (N_13787,N_13597,N_13598);
or U13788 (N_13788,N_13580,N_13526);
and U13789 (N_13789,N_13537,N_13528);
xor U13790 (N_13790,N_13573,N_13463);
and U13791 (N_13791,N_13462,N_13577);
xor U13792 (N_13792,N_13497,N_13560);
xor U13793 (N_13793,N_13404,N_13566);
nand U13794 (N_13794,N_13467,N_13549);
xor U13795 (N_13795,N_13416,N_13405);
xnor U13796 (N_13796,N_13423,N_13416);
nor U13797 (N_13797,N_13416,N_13562);
or U13798 (N_13798,N_13497,N_13465);
nor U13799 (N_13799,N_13523,N_13476);
nand U13800 (N_13800,N_13604,N_13681);
or U13801 (N_13801,N_13605,N_13752);
and U13802 (N_13802,N_13626,N_13624);
xnor U13803 (N_13803,N_13747,N_13716);
xnor U13804 (N_13804,N_13691,N_13762);
and U13805 (N_13805,N_13650,N_13766);
or U13806 (N_13806,N_13619,N_13763);
nand U13807 (N_13807,N_13765,N_13699);
and U13808 (N_13808,N_13744,N_13780);
nand U13809 (N_13809,N_13761,N_13746);
or U13810 (N_13810,N_13674,N_13782);
or U13811 (N_13811,N_13729,N_13673);
nor U13812 (N_13812,N_13601,N_13771);
and U13813 (N_13813,N_13613,N_13730);
or U13814 (N_13814,N_13795,N_13634);
nand U13815 (N_13815,N_13748,N_13724);
or U13816 (N_13816,N_13631,N_13779);
or U13817 (N_13817,N_13714,N_13666);
or U13818 (N_13818,N_13687,N_13740);
or U13819 (N_13819,N_13715,N_13727);
or U13820 (N_13820,N_13722,N_13679);
nor U13821 (N_13821,N_13770,N_13788);
nor U13822 (N_13822,N_13647,N_13701);
nand U13823 (N_13823,N_13757,N_13657);
nor U13824 (N_13824,N_13649,N_13678);
nand U13825 (N_13825,N_13682,N_13753);
nor U13826 (N_13826,N_13713,N_13669);
nor U13827 (N_13827,N_13768,N_13670);
nand U13828 (N_13828,N_13690,N_13778);
xnor U13829 (N_13829,N_13789,N_13667);
xnor U13830 (N_13830,N_13602,N_13607);
and U13831 (N_13831,N_13772,N_13643);
nand U13832 (N_13832,N_13776,N_13775);
and U13833 (N_13833,N_13694,N_13630);
and U13834 (N_13834,N_13692,N_13709);
nor U13835 (N_13835,N_13790,N_13705);
and U13836 (N_13836,N_13660,N_13787);
xnor U13837 (N_13837,N_13668,N_13615);
xor U13838 (N_13838,N_13749,N_13664);
nor U13839 (N_13839,N_13783,N_13606);
nand U13840 (N_13840,N_13652,N_13756);
and U13841 (N_13841,N_13723,N_13791);
nor U13842 (N_13842,N_13629,N_13739);
xor U13843 (N_13843,N_13745,N_13616);
or U13844 (N_13844,N_13703,N_13720);
or U13845 (N_13845,N_13696,N_13659);
nor U13846 (N_13846,N_13797,N_13738);
nor U13847 (N_13847,N_13632,N_13702);
or U13848 (N_13848,N_13671,N_13640);
or U13849 (N_13849,N_13733,N_13612);
and U13850 (N_13850,N_13793,N_13654);
and U13851 (N_13851,N_13655,N_13689);
or U13852 (N_13852,N_13777,N_13697);
nand U13853 (N_13853,N_13620,N_13798);
or U13854 (N_13854,N_13618,N_13623);
and U13855 (N_13855,N_13611,N_13719);
or U13856 (N_13856,N_13760,N_13656);
nand U13857 (N_13857,N_13741,N_13755);
nand U13858 (N_13858,N_13698,N_13653);
nand U13859 (N_13859,N_13707,N_13717);
and U13860 (N_13860,N_13773,N_13711);
nand U13861 (N_13861,N_13665,N_13638);
xor U13862 (N_13862,N_13635,N_13710);
or U13863 (N_13863,N_13642,N_13675);
nor U13864 (N_13864,N_13636,N_13663);
and U13865 (N_13865,N_13651,N_13676);
xor U13866 (N_13866,N_13648,N_13695);
nor U13867 (N_13867,N_13683,N_13784);
nand U13868 (N_13868,N_13641,N_13743);
and U13869 (N_13869,N_13786,N_13700);
and U13870 (N_13870,N_13672,N_13637);
nor U13871 (N_13871,N_13628,N_13600);
xnor U13872 (N_13872,N_13658,N_13609);
nor U13873 (N_13873,N_13774,N_13685);
xor U13874 (N_13874,N_13767,N_13754);
xnor U13875 (N_13875,N_13610,N_13662);
nand U13876 (N_13876,N_13646,N_13799);
and U13877 (N_13877,N_13759,N_13645);
and U13878 (N_13878,N_13785,N_13684);
and U13879 (N_13879,N_13627,N_13621);
and U13880 (N_13880,N_13712,N_13680);
nor U13881 (N_13881,N_13794,N_13751);
xor U13882 (N_13882,N_13734,N_13758);
nor U13883 (N_13883,N_13677,N_13603);
xor U13884 (N_13884,N_13608,N_13750);
or U13885 (N_13885,N_13764,N_13639);
or U13886 (N_13886,N_13617,N_13735);
and U13887 (N_13887,N_13728,N_13693);
and U13888 (N_13888,N_13644,N_13725);
xor U13889 (N_13889,N_13726,N_13625);
and U13890 (N_13890,N_13633,N_13614);
xor U13891 (N_13891,N_13718,N_13792);
or U13892 (N_13892,N_13769,N_13721);
xnor U13893 (N_13893,N_13704,N_13731);
or U13894 (N_13894,N_13688,N_13622);
nor U13895 (N_13895,N_13732,N_13706);
or U13896 (N_13896,N_13686,N_13737);
nor U13897 (N_13897,N_13796,N_13736);
nor U13898 (N_13898,N_13708,N_13742);
or U13899 (N_13899,N_13781,N_13661);
or U13900 (N_13900,N_13649,N_13760);
nand U13901 (N_13901,N_13727,N_13618);
and U13902 (N_13902,N_13642,N_13631);
xnor U13903 (N_13903,N_13644,N_13767);
xor U13904 (N_13904,N_13721,N_13628);
nor U13905 (N_13905,N_13705,N_13700);
and U13906 (N_13906,N_13703,N_13629);
nor U13907 (N_13907,N_13735,N_13742);
nand U13908 (N_13908,N_13794,N_13671);
or U13909 (N_13909,N_13651,N_13653);
xor U13910 (N_13910,N_13644,N_13651);
or U13911 (N_13911,N_13619,N_13667);
nor U13912 (N_13912,N_13723,N_13653);
or U13913 (N_13913,N_13708,N_13755);
or U13914 (N_13914,N_13612,N_13634);
or U13915 (N_13915,N_13784,N_13627);
xnor U13916 (N_13916,N_13717,N_13792);
nand U13917 (N_13917,N_13765,N_13622);
nand U13918 (N_13918,N_13764,N_13638);
nand U13919 (N_13919,N_13738,N_13626);
nor U13920 (N_13920,N_13660,N_13614);
xnor U13921 (N_13921,N_13657,N_13676);
nand U13922 (N_13922,N_13752,N_13711);
or U13923 (N_13923,N_13649,N_13763);
xnor U13924 (N_13924,N_13699,N_13654);
nand U13925 (N_13925,N_13678,N_13696);
xnor U13926 (N_13926,N_13776,N_13655);
nor U13927 (N_13927,N_13757,N_13670);
and U13928 (N_13928,N_13652,N_13762);
or U13929 (N_13929,N_13671,N_13684);
nor U13930 (N_13930,N_13776,N_13651);
nor U13931 (N_13931,N_13673,N_13769);
or U13932 (N_13932,N_13715,N_13601);
or U13933 (N_13933,N_13681,N_13612);
nand U13934 (N_13934,N_13777,N_13635);
and U13935 (N_13935,N_13748,N_13713);
xnor U13936 (N_13936,N_13711,N_13600);
nand U13937 (N_13937,N_13606,N_13689);
nand U13938 (N_13938,N_13770,N_13657);
and U13939 (N_13939,N_13650,N_13647);
xor U13940 (N_13940,N_13782,N_13774);
or U13941 (N_13941,N_13657,N_13744);
nor U13942 (N_13942,N_13719,N_13730);
or U13943 (N_13943,N_13617,N_13642);
or U13944 (N_13944,N_13660,N_13714);
and U13945 (N_13945,N_13613,N_13717);
nand U13946 (N_13946,N_13682,N_13681);
nand U13947 (N_13947,N_13735,N_13670);
xnor U13948 (N_13948,N_13786,N_13659);
xor U13949 (N_13949,N_13677,N_13750);
nor U13950 (N_13950,N_13620,N_13687);
xor U13951 (N_13951,N_13675,N_13678);
nand U13952 (N_13952,N_13654,N_13719);
or U13953 (N_13953,N_13701,N_13745);
nand U13954 (N_13954,N_13769,N_13699);
nor U13955 (N_13955,N_13619,N_13656);
nor U13956 (N_13956,N_13649,N_13660);
or U13957 (N_13957,N_13704,N_13678);
xor U13958 (N_13958,N_13703,N_13635);
nor U13959 (N_13959,N_13723,N_13618);
or U13960 (N_13960,N_13606,N_13611);
nand U13961 (N_13961,N_13653,N_13713);
and U13962 (N_13962,N_13779,N_13652);
nor U13963 (N_13963,N_13646,N_13636);
nand U13964 (N_13964,N_13620,N_13735);
or U13965 (N_13965,N_13729,N_13661);
and U13966 (N_13966,N_13757,N_13678);
and U13967 (N_13967,N_13762,N_13636);
nand U13968 (N_13968,N_13623,N_13678);
nand U13969 (N_13969,N_13774,N_13719);
xnor U13970 (N_13970,N_13684,N_13750);
xor U13971 (N_13971,N_13675,N_13689);
or U13972 (N_13972,N_13765,N_13638);
xnor U13973 (N_13973,N_13644,N_13785);
nor U13974 (N_13974,N_13607,N_13608);
xor U13975 (N_13975,N_13725,N_13766);
xnor U13976 (N_13976,N_13757,N_13610);
xnor U13977 (N_13977,N_13601,N_13719);
or U13978 (N_13978,N_13768,N_13641);
nand U13979 (N_13979,N_13631,N_13680);
nand U13980 (N_13980,N_13789,N_13619);
and U13981 (N_13981,N_13628,N_13715);
and U13982 (N_13982,N_13780,N_13623);
nand U13983 (N_13983,N_13729,N_13676);
nand U13984 (N_13984,N_13767,N_13623);
xor U13985 (N_13985,N_13797,N_13640);
xnor U13986 (N_13986,N_13705,N_13702);
xor U13987 (N_13987,N_13794,N_13773);
xnor U13988 (N_13988,N_13624,N_13742);
or U13989 (N_13989,N_13712,N_13652);
nand U13990 (N_13990,N_13690,N_13651);
and U13991 (N_13991,N_13770,N_13653);
nor U13992 (N_13992,N_13622,N_13685);
or U13993 (N_13993,N_13732,N_13632);
nor U13994 (N_13994,N_13633,N_13684);
or U13995 (N_13995,N_13620,N_13691);
nor U13996 (N_13996,N_13794,N_13725);
nor U13997 (N_13997,N_13797,N_13647);
and U13998 (N_13998,N_13785,N_13660);
nand U13999 (N_13999,N_13734,N_13695);
xor U14000 (N_14000,N_13938,N_13990);
xnor U14001 (N_14001,N_13962,N_13986);
nand U14002 (N_14002,N_13993,N_13861);
nor U14003 (N_14003,N_13911,N_13954);
or U14004 (N_14004,N_13831,N_13974);
or U14005 (N_14005,N_13995,N_13916);
nand U14006 (N_14006,N_13926,N_13830);
or U14007 (N_14007,N_13818,N_13915);
xnor U14008 (N_14008,N_13906,N_13920);
xor U14009 (N_14009,N_13869,N_13876);
and U14010 (N_14010,N_13973,N_13883);
nor U14011 (N_14011,N_13900,N_13870);
and U14012 (N_14012,N_13866,N_13801);
and U14013 (N_14013,N_13820,N_13958);
and U14014 (N_14014,N_13942,N_13816);
and U14015 (N_14015,N_13997,N_13852);
and U14016 (N_14016,N_13940,N_13922);
or U14017 (N_14017,N_13827,N_13909);
xor U14018 (N_14018,N_13838,N_13889);
and U14019 (N_14019,N_13985,N_13821);
xnor U14020 (N_14020,N_13809,N_13982);
and U14021 (N_14021,N_13819,N_13892);
xor U14022 (N_14022,N_13865,N_13860);
nand U14023 (N_14023,N_13858,N_13951);
and U14024 (N_14024,N_13929,N_13934);
or U14025 (N_14025,N_13898,N_13989);
nand U14026 (N_14026,N_13914,N_13862);
and U14027 (N_14027,N_13825,N_13808);
nand U14028 (N_14028,N_13970,N_13833);
and U14029 (N_14029,N_13873,N_13853);
or U14030 (N_14030,N_13842,N_13921);
and U14031 (N_14031,N_13857,N_13882);
nand U14032 (N_14032,N_13885,N_13980);
nand U14033 (N_14033,N_13988,N_13810);
or U14034 (N_14034,N_13925,N_13859);
nand U14035 (N_14035,N_13987,N_13966);
and U14036 (N_14036,N_13991,N_13813);
and U14037 (N_14037,N_13981,N_13881);
and U14038 (N_14038,N_13978,N_13941);
nand U14039 (N_14039,N_13826,N_13891);
and U14040 (N_14040,N_13939,N_13868);
xor U14041 (N_14041,N_13895,N_13956);
and U14042 (N_14042,N_13888,N_13907);
xor U14043 (N_14043,N_13928,N_13967);
or U14044 (N_14044,N_13805,N_13975);
or U14045 (N_14045,N_13847,N_13935);
nand U14046 (N_14046,N_13824,N_13903);
or U14047 (N_14047,N_13912,N_13904);
or U14048 (N_14048,N_13930,N_13846);
nor U14049 (N_14049,N_13936,N_13945);
or U14050 (N_14050,N_13957,N_13984);
nand U14051 (N_14051,N_13812,N_13952);
xor U14052 (N_14052,N_13905,N_13843);
and U14053 (N_14053,N_13927,N_13815);
and U14054 (N_14054,N_13863,N_13834);
xor U14055 (N_14055,N_13976,N_13806);
xor U14056 (N_14056,N_13923,N_13851);
and U14057 (N_14057,N_13998,N_13867);
nor U14058 (N_14058,N_13800,N_13844);
nand U14059 (N_14059,N_13886,N_13959);
nor U14060 (N_14060,N_13880,N_13872);
and U14061 (N_14061,N_13999,N_13949);
nor U14062 (N_14062,N_13947,N_13807);
and U14063 (N_14063,N_13953,N_13965);
and U14064 (N_14064,N_13902,N_13878);
nand U14065 (N_14065,N_13823,N_13829);
or U14066 (N_14066,N_13811,N_13893);
and U14067 (N_14067,N_13964,N_13874);
and U14068 (N_14068,N_13943,N_13884);
nor U14069 (N_14069,N_13832,N_13828);
or U14070 (N_14070,N_13968,N_13899);
nor U14071 (N_14071,N_13850,N_13897);
nand U14072 (N_14072,N_13983,N_13854);
or U14073 (N_14073,N_13950,N_13937);
or U14074 (N_14074,N_13890,N_13817);
nor U14075 (N_14075,N_13996,N_13908);
or U14076 (N_14076,N_13960,N_13896);
nand U14077 (N_14077,N_13887,N_13932);
nand U14078 (N_14078,N_13979,N_13918);
or U14079 (N_14079,N_13848,N_13955);
and U14080 (N_14080,N_13835,N_13841);
xnor U14081 (N_14081,N_13845,N_13840);
nor U14082 (N_14082,N_13931,N_13910);
and U14083 (N_14083,N_13804,N_13877);
nand U14084 (N_14084,N_13864,N_13961);
or U14085 (N_14085,N_13901,N_13913);
xor U14086 (N_14086,N_13994,N_13879);
nor U14087 (N_14087,N_13871,N_13917);
and U14088 (N_14088,N_13977,N_13855);
nand U14089 (N_14089,N_13919,N_13836);
or U14090 (N_14090,N_13933,N_13875);
and U14091 (N_14091,N_13849,N_13839);
and U14092 (N_14092,N_13972,N_13814);
nand U14093 (N_14093,N_13894,N_13856);
xnor U14094 (N_14094,N_13969,N_13822);
and U14095 (N_14095,N_13944,N_13802);
nor U14096 (N_14096,N_13803,N_13971);
xor U14097 (N_14097,N_13963,N_13948);
or U14098 (N_14098,N_13946,N_13837);
xor U14099 (N_14099,N_13924,N_13992);
and U14100 (N_14100,N_13913,N_13927);
or U14101 (N_14101,N_13915,N_13886);
nor U14102 (N_14102,N_13887,N_13875);
and U14103 (N_14103,N_13867,N_13869);
nand U14104 (N_14104,N_13912,N_13833);
or U14105 (N_14105,N_13928,N_13981);
nand U14106 (N_14106,N_13901,N_13848);
and U14107 (N_14107,N_13947,N_13863);
nor U14108 (N_14108,N_13965,N_13856);
nor U14109 (N_14109,N_13971,N_13844);
xnor U14110 (N_14110,N_13824,N_13860);
nor U14111 (N_14111,N_13865,N_13811);
or U14112 (N_14112,N_13897,N_13932);
xnor U14113 (N_14113,N_13971,N_13996);
or U14114 (N_14114,N_13984,N_13982);
nand U14115 (N_14115,N_13805,N_13800);
xnor U14116 (N_14116,N_13814,N_13857);
or U14117 (N_14117,N_13947,N_13825);
nand U14118 (N_14118,N_13904,N_13973);
xor U14119 (N_14119,N_13818,N_13823);
xnor U14120 (N_14120,N_13884,N_13926);
nand U14121 (N_14121,N_13939,N_13886);
nor U14122 (N_14122,N_13930,N_13904);
nand U14123 (N_14123,N_13986,N_13842);
or U14124 (N_14124,N_13895,N_13896);
or U14125 (N_14125,N_13977,N_13973);
or U14126 (N_14126,N_13824,N_13851);
xor U14127 (N_14127,N_13816,N_13948);
nor U14128 (N_14128,N_13924,N_13833);
nand U14129 (N_14129,N_13872,N_13923);
nand U14130 (N_14130,N_13884,N_13982);
xor U14131 (N_14131,N_13994,N_13856);
or U14132 (N_14132,N_13926,N_13923);
xor U14133 (N_14133,N_13995,N_13852);
nor U14134 (N_14134,N_13887,N_13988);
and U14135 (N_14135,N_13901,N_13958);
xnor U14136 (N_14136,N_13928,N_13941);
or U14137 (N_14137,N_13803,N_13828);
nor U14138 (N_14138,N_13904,N_13939);
or U14139 (N_14139,N_13844,N_13872);
nand U14140 (N_14140,N_13950,N_13941);
and U14141 (N_14141,N_13980,N_13816);
nor U14142 (N_14142,N_13972,N_13865);
nand U14143 (N_14143,N_13961,N_13998);
xnor U14144 (N_14144,N_13996,N_13976);
and U14145 (N_14145,N_13815,N_13945);
nor U14146 (N_14146,N_13918,N_13861);
nor U14147 (N_14147,N_13842,N_13829);
xnor U14148 (N_14148,N_13925,N_13969);
xnor U14149 (N_14149,N_13981,N_13825);
and U14150 (N_14150,N_13889,N_13824);
and U14151 (N_14151,N_13874,N_13902);
or U14152 (N_14152,N_13978,N_13869);
or U14153 (N_14153,N_13900,N_13859);
nor U14154 (N_14154,N_13958,N_13982);
nand U14155 (N_14155,N_13963,N_13843);
nand U14156 (N_14156,N_13860,N_13830);
nor U14157 (N_14157,N_13889,N_13977);
nor U14158 (N_14158,N_13913,N_13892);
and U14159 (N_14159,N_13927,N_13985);
xor U14160 (N_14160,N_13949,N_13872);
nand U14161 (N_14161,N_13918,N_13947);
and U14162 (N_14162,N_13909,N_13911);
nor U14163 (N_14163,N_13963,N_13910);
or U14164 (N_14164,N_13872,N_13912);
nor U14165 (N_14165,N_13850,N_13967);
nand U14166 (N_14166,N_13887,N_13985);
xnor U14167 (N_14167,N_13978,N_13950);
and U14168 (N_14168,N_13936,N_13824);
nand U14169 (N_14169,N_13924,N_13918);
or U14170 (N_14170,N_13892,N_13846);
nor U14171 (N_14171,N_13989,N_13865);
xnor U14172 (N_14172,N_13928,N_13936);
and U14173 (N_14173,N_13976,N_13944);
and U14174 (N_14174,N_13876,N_13870);
nand U14175 (N_14175,N_13889,N_13890);
and U14176 (N_14176,N_13847,N_13944);
and U14177 (N_14177,N_13949,N_13986);
nand U14178 (N_14178,N_13960,N_13866);
nor U14179 (N_14179,N_13917,N_13947);
or U14180 (N_14180,N_13900,N_13960);
nand U14181 (N_14181,N_13959,N_13955);
and U14182 (N_14182,N_13819,N_13872);
nor U14183 (N_14183,N_13999,N_13976);
nand U14184 (N_14184,N_13983,N_13877);
xnor U14185 (N_14185,N_13996,N_13831);
nor U14186 (N_14186,N_13993,N_13839);
nor U14187 (N_14187,N_13980,N_13909);
xor U14188 (N_14188,N_13927,N_13947);
nand U14189 (N_14189,N_13898,N_13982);
and U14190 (N_14190,N_13977,N_13840);
nor U14191 (N_14191,N_13938,N_13892);
and U14192 (N_14192,N_13842,N_13957);
and U14193 (N_14193,N_13809,N_13987);
or U14194 (N_14194,N_13842,N_13904);
nand U14195 (N_14195,N_13862,N_13983);
xor U14196 (N_14196,N_13922,N_13880);
or U14197 (N_14197,N_13953,N_13856);
nand U14198 (N_14198,N_13820,N_13979);
and U14199 (N_14199,N_13879,N_13929);
xnor U14200 (N_14200,N_14063,N_14131);
or U14201 (N_14201,N_14195,N_14065);
nand U14202 (N_14202,N_14146,N_14070);
nor U14203 (N_14203,N_14079,N_14133);
nand U14204 (N_14204,N_14092,N_14023);
and U14205 (N_14205,N_14118,N_14190);
or U14206 (N_14206,N_14099,N_14106);
nand U14207 (N_14207,N_14179,N_14056);
and U14208 (N_14208,N_14198,N_14066);
nor U14209 (N_14209,N_14016,N_14164);
nand U14210 (N_14210,N_14017,N_14043);
xnor U14211 (N_14211,N_14059,N_14033);
and U14212 (N_14212,N_14109,N_14176);
or U14213 (N_14213,N_14135,N_14015);
and U14214 (N_14214,N_14058,N_14183);
nand U14215 (N_14215,N_14025,N_14018);
nand U14216 (N_14216,N_14062,N_14029);
nor U14217 (N_14217,N_14162,N_14104);
xor U14218 (N_14218,N_14119,N_14169);
nand U14219 (N_14219,N_14137,N_14101);
nor U14220 (N_14220,N_14021,N_14042);
xor U14221 (N_14221,N_14117,N_14088);
xnor U14222 (N_14222,N_14178,N_14161);
and U14223 (N_14223,N_14168,N_14089);
or U14224 (N_14224,N_14165,N_14108);
nor U14225 (N_14225,N_14091,N_14081);
or U14226 (N_14226,N_14160,N_14004);
xnor U14227 (N_14227,N_14075,N_14187);
nand U14228 (N_14228,N_14123,N_14036);
nor U14229 (N_14229,N_14115,N_14103);
and U14230 (N_14230,N_14124,N_14111);
or U14231 (N_14231,N_14053,N_14147);
xnor U14232 (N_14232,N_14002,N_14011);
xnor U14233 (N_14233,N_14170,N_14128);
or U14234 (N_14234,N_14148,N_14095);
and U14235 (N_14235,N_14048,N_14110);
or U14236 (N_14236,N_14193,N_14166);
xnor U14237 (N_14237,N_14113,N_14126);
nand U14238 (N_14238,N_14199,N_14076);
nor U14239 (N_14239,N_14112,N_14060);
and U14240 (N_14240,N_14151,N_14083);
nor U14241 (N_14241,N_14153,N_14097);
and U14242 (N_14242,N_14180,N_14082);
or U14243 (N_14243,N_14094,N_14055);
and U14244 (N_14244,N_14049,N_14030);
and U14245 (N_14245,N_14022,N_14090);
and U14246 (N_14246,N_14034,N_14039);
and U14247 (N_14247,N_14177,N_14144);
or U14248 (N_14248,N_14149,N_14035);
nand U14249 (N_14249,N_14116,N_14143);
or U14250 (N_14250,N_14172,N_14121);
xor U14251 (N_14251,N_14037,N_14105);
and U14252 (N_14252,N_14064,N_14085);
nor U14253 (N_14253,N_14073,N_14127);
nor U14254 (N_14254,N_14159,N_14173);
or U14255 (N_14255,N_14197,N_14132);
nor U14256 (N_14256,N_14031,N_14068);
or U14257 (N_14257,N_14093,N_14012);
nand U14258 (N_14258,N_14196,N_14040);
xor U14259 (N_14259,N_14071,N_14155);
xnor U14260 (N_14260,N_14057,N_14009);
nor U14261 (N_14261,N_14045,N_14100);
or U14262 (N_14262,N_14086,N_14019);
nand U14263 (N_14263,N_14005,N_14129);
and U14264 (N_14264,N_14114,N_14156);
and U14265 (N_14265,N_14051,N_14014);
or U14266 (N_14266,N_14098,N_14006);
nand U14267 (N_14267,N_14054,N_14158);
nand U14268 (N_14268,N_14167,N_14122);
or U14269 (N_14269,N_14084,N_14134);
nand U14270 (N_14270,N_14026,N_14181);
nor U14271 (N_14271,N_14182,N_14171);
nand U14272 (N_14272,N_14138,N_14069);
xnor U14273 (N_14273,N_14052,N_14154);
xor U14274 (N_14274,N_14067,N_14003);
nor U14275 (N_14275,N_14078,N_14087);
or U14276 (N_14276,N_14130,N_14008);
xnor U14277 (N_14277,N_14120,N_14136);
xnor U14278 (N_14278,N_14010,N_14024);
xnor U14279 (N_14279,N_14032,N_14044);
nand U14280 (N_14280,N_14185,N_14194);
nand U14281 (N_14281,N_14163,N_14020);
or U14282 (N_14282,N_14061,N_14077);
nor U14283 (N_14283,N_14028,N_14157);
xor U14284 (N_14284,N_14140,N_14184);
or U14285 (N_14285,N_14047,N_14152);
and U14286 (N_14286,N_14027,N_14041);
nor U14287 (N_14287,N_14150,N_14080);
nand U14288 (N_14288,N_14107,N_14072);
or U14289 (N_14289,N_14096,N_14000);
nor U14290 (N_14290,N_14007,N_14174);
nand U14291 (N_14291,N_14001,N_14189);
nor U14292 (N_14292,N_14013,N_14145);
or U14293 (N_14293,N_14192,N_14188);
and U14294 (N_14294,N_14125,N_14175);
xor U14295 (N_14295,N_14191,N_14046);
or U14296 (N_14296,N_14141,N_14139);
nor U14297 (N_14297,N_14142,N_14050);
and U14298 (N_14298,N_14102,N_14038);
or U14299 (N_14299,N_14186,N_14074);
nand U14300 (N_14300,N_14121,N_14049);
nand U14301 (N_14301,N_14199,N_14100);
xor U14302 (N_14302,N_14079,N_14131);
or U14303 (N_14303,N_14023,N_14153);
or U14304 (N_14304,N_14151,N_14082);
nand U14305 (N_14305,N_14003,N_14006);
xor U14306 (N_14306,N_14133,N_14138);
nor U14307 (N_14307,N_14183,N_14109);
or U14308 (N_14308,N_14046,N_14100);
and U14309 (N_14309,N_14090,N_14168);
xnor U14310 (N_14310,N_14135,N_14021);
nor U14311 (N_14311,N_14053,N_14025);
nor U14312 (N_14312,N_14167,N_14048);
nand U14313 (N_14313,N_14107,N_14047);
or U14314 (N_14314,N_14149,N_14031);
nand U14315 (N_14315,N_14052,N_14007);
nor U14316 (N_14316,N_14092,N_14160);
or U14317 (N_14317,N_14043,N_14141);
or U14318 (N_14318,N_14178,N_14194);
and U14319 (N_14319,N_14056,N_14172);
nand U14320 (N_14320,N_14110,N_14068);
nand U14321 (N_14321,N_14167,N_14187);
or U14322 (N_14322,N_14019,N_14008);
xnor U14323 (N_14323,N_14009,N_14131);
nor U14324 (N_14324,N_14104,N_14139);
nor U14325 (N_14325,N_14147,N_14197);
xnor U14326 (N_14326,N_14077,N_14043);
xnor U14327 (N_14327,N_14042,N_14176);
nand U14328 (N_14328,N_14021,N_14123);
nor U14329 (N_14329,N_14131,N_14024);
xor U14330 (N_14330,N_14034,N_14030);
or U14331 (N_14331,N_14139,N_14162);
nand U14332 (N_14332,N_14028,N_14138);
nand U14333 (N_14333,N_14019,N_14158);
or U14334 (N_14334,N_14123,N_14188);
nor U14335 (N_14335,N_14147,N_14049);
or U14336 (N_14336,N_14196,N_14000);
and U14337 (N_14337,N_14082,N_14190);
and U14338 (N_14338,N_14051,N_14117);
nor U14339 (N_14339,N_14071,N_14176);
nor U14340 (N_14340,N_14156,N_14138);
xnor U14341 (N_14341,N_14081,N_14042);
nor U14342 (N_14342,N_14089,N_14063);
nor U14343 (N_14343,N_14107,N_14086);
xor U14344 (N_14344,N_14132,N_14090);
nand U14345 (N_14345,N_14131,N_14029);
or U14346 (N_14346,N_14011,N_14194);
nand U14347 (N_14347,N_14099,N_14185);
or U14348 (N_14348,N_14157,N_14140);
nand U14349 (N_14349,N_14149,N_14170);
nand U14350 (N_14350,N_14192,N_14086);
or U14351 (N_14351,N_14150,N_14085);
xor U14352 (N_14352,N_14151,N_14004);
nor U14353 (N_14353,N_14046,N_14053);
xnor U14354 (N_14354,N_14024,N_14076);
and U14355 (N_14355,N_14103,N_14059);
xor U14356 (N_14356,N_14175,N_14036);
and U14357 (N_14357,N_14099,N_14033);
and U14358 (N_14358,N_14047,N_14121);
nor U14359 (N_14359,N_14186,N_14147);
and U14360 (N_14360,N_14194,N_14078);
nor U14361 (N_14361,N_14059,N_14003);
or U14362 (N_14362,N_14151,N_14180);
xnor U14363 (N_14363,N_14107,N_14192);
nor U14364 (N_14364,N_14067,N_14150);
or U14365 (N_14365,N_14085,N_14186);
nor U14366 (N_14366,N_14100,N_14036);
xor U14367 (N_14367,N_14036,N_14059);
or U14368 (N_14368,N_14188,N_14108);
and U14369 (N_14369,N_14160,N_14042);
xor U14370 (N_14370,N_14146,N_14017);
nand U14371 (N_14371,N_14186,N_14183);
nand U14372 (N_14372,N_14185,N_14064);
or U14373 (N_14373,N_14132,N_14066);
nor U14374 (N_14374,N_14073,N_14023);
xnor U14375 (N_14375,N_14109,N_14013);
xor U14376 (N_14376,N_14150,N_14090);
nand U14377 (N_14377,N_14055,N_14118);
and U14378 (N_14378,N_14107,N_14185);
or U14379 (N_14379,N_14198,N_14180);
and U14380 (N_14380,N_14130,N_14144);
nand U14381 (N_14381,N_14119,N_14041);
xor U14382 (N_14382,N_14140,N_14150);
nand U14383 (N_14383,N_14129,N_14039);
and U14384 (N_14384,N_14119,N_14187);
and U14385 (N_14385,N_14172,N_14116);
nor U14386 (N_14386,N_14127,N_14040);
nand U14387 (N_14387,N_14116,N_14101);
xnor U14388 (N_14388,N_14106,N_14019);
nor U14389 (N_14389,N_14061,N_14179);
or U14390 (N_14390,N_14106,N_14139);
or U14391 (N_14391,N_14058,N_14146);
nor U14392 (N_14392,N_14110,N_14047);
nand U14393 (N_14393,N_14103,N_14057);
xnor U14394 (N_14394,N_14173,N_14162);
xor U14395 (N_14395,N_14139,N_14199);
nor U14396 (N_14396,N_14117,N_14066);
nand U14397 (N_14397,N_14014,N_14155);
and U14398 (N_14398,N_14171,N_14032);
and U14399 (N_14399,N_14085,N_14013);
nand U14400 (N_14400,N_14230,N_14285);
xor U14401 (N_14401,N_14224,N_14214);
and U14402 (N_14402,N_14227,N_14378);
and U14403 (N_14403,N_14210,N_14320);
nor U14404 (N_14404,N_14390,N_14259);
nand U14405 (N_14405,N_14225,N_14267);
or U14406 (N_14406,N_14266,N_14352);
nand U14407 (N_14407,N_14382,N_14242);
or U14408 (N_14408,N_14358,N_14249);
nand U14409 (N_14409,N_14330,N_14340);
or U14410 (N_14410,N_14235,N_14391);
xnor U14411 (N_14411,N_14248,N_14346);
xnor U14412 (N_14412,N_14206,N_14331);
or U14413 (N_14413,N_14318,N_14322);
nor U14414 (N_14414,N_14361,N_14234);
and U14415 (N_14415,N_14363,N_14332);
xnor U14416 (N_14416,N_14294,N_14282);
or U14417 (N_14417,N_14395,N_14304);
nand U14418 (N_14418,N_14205,N_14243);
nor U14419 (N_14419,N_14386,N_14251);
and U14420 (N_14420,N_14238,N_14219);
nand U14421 (N_14421,N_14275,N_14292);
nand U14422 (N_14422,N_14376,N_14260);
nor U14423 (N_14423,N_14334,N_14208);
and U14424 (N_14424,N_14273,N_14308);
and U14425 (N_14425,N_14244,N_14222);
and U14426 (N_14426,N_14384,N_14204);
nand U14427 (N_14427,N_14231,N_14396);
or U14428 (N_14428,N_14217,N_14379);
nor U14429 (N_14429,N_14355,N_14311);
xor U14430 (N_14430,N_14293,N_14271);
and U14431 (N_14431,N_14344,N_14364);
nand U14432 (N_14432,N_14246,N_14220);
and U14433 (N_14433,N_14369,N_14255);
or U14434 (N_14434,N_14239,N_14365);
and U14435 (N_14435,N_14232,N_14223);
or U14436 (N_14436,N_14201,N_14336);
or U14437 (N_14437,N_14272,N_14348);
nor U14438 (N_14438,N_14302,N_14200);
or U14439 (N_14439,N_14342,N_14324);
nand U14440 (N_14440,N_14307,N_14221);
nand U14441 (N_14441,N_14269,N_14303);
xor U14442 (N_14442,N_14306,N_14247);
and U14443 (N_14443,N_14375,N_14368);
nand U14444 (N_14444,N_14281,N_14290);
and U14445 (N_14445,N_14398,N_14343);
nand U14446 (N_14446,N_14328,N_14264);
or U14447 (N_14447,N_14236,N_14256);
or U14448 (N_14448,N_14353,N_14357);
and U14449 (N_14449,N_14354,N_14257);
nor U14450 (N_14450,N_14211,N_14356);
or U14451 (N_14451,N_14359,N_14276);
nand U14452 (N_14452,N_14289,N_14349);
or U14453 (N_14453,N_14215,N_14370);
nor U14454 (N_14454,N_14245,N_14310);
nor U14455 (N_14455,N_14362,N_14263);
nand U14456 (N_14456,N_14202,N_14287);
or U14457 (N_14457,N_14323,N_14216);
nor U14458 (N_14458,N_14209,N_14270);
nor U14459 (N_14459,N_14397,N_14387);
nand U14460 (N_14460,N_14207,N_14284);
nand U14461 (N_14461,N_14291,N_14312);
xnor U14462 (N_14462,N_14277,N_14381);
and U14463 (N_14463,N_14262,N_14237);
xnor U14464 (N_14464,N_14258,N_14393);
or U14465 (N_14465,N_14288,N_14394);
nand U14466 (N_14466,N_14333,N_14351);
nor U14467 (N_14467,N_14228,N_14253);
or U14468 (N_14468,N_14229,N_14317);
nor U14469 (N_14469,N_14377,N_14241);
nor U14470 (N_14470,N_14297,N_14345);
or U14471 (N_14471,N_14374,N_14383);
or U14472 (N_14472,N_14389,N_14373);
xor U14473 (N_14473,N_14265,N_14233);
or U14474 (N_14474,N_14296,N_14326);
nand U14475 (N_14475,N_14321,N_14347);
nor U14476 (N_14476,N_14371,N_14315);
and U14477 (N_14477,N_14274,N_14240);
xnor U14478 (N_14478,N_14309,N_14341);
or U14479 (N_14479,N_14299,N_14298);
and U14480 (N_14480,N_14252,N_14337);
nor U14481 (N_14481,N_14329,N_14392);
nand U14482 (N_14482,N_14319,N_14305);
xnor U14483 (N_14483,N_14278,N_14366);
nor U14484 (N_14484,N_14250,N_14280);
xnor U14485 (N_14485,N_14279,N_14218);
nor U14486 (N_14486,N_14399,N_14372);
or U14487 (N_14487,N_14388,N_14226);
or U14488 (N_14488,N_14295,N_14385);
or U14489 (N_14489,N_14327,N_14261);
nor U14490 (N_14490,N_14360,N_14286);
xor U14491 (N_14491,N_14313,N_14380);
nor U14492 (N_14492,N_14213,N_14301);
or U14493 (N_14493,N_14335,N_14254);
nand U14494 (N_14494,N_14212,N_14367);
or U14495 (N_14495,N_14283,N_14316);
and U14496 (N_14496,N_14339,N_14350);
xnor U14497 (N_14497,N_14314,N_14268);
and U14498 (N_14498,N_14338,N_14325);
nand U14499 (N_14499,N_14203,N_14300);
nand U14500 (N_14500,N_14221,N_14341);
nand U14501 (N_14501,N_14298,N_14288);
nand U14502 (N_14502,N_14274,N_14337);
nand U14503 (N_14503,N_14330,N_14392);
nor U14504 (N_14504,N_14379,N_14265);
xnor U14505 (N_14505,N_14262,N_14217);
or U14506 (N_14506,N_14343,N_14242);
and U14507 (N_14507,N_14395,N_14305);
or U14508 (N_14508,N_14201,N_14259);
xnor U14509 (N_14509,N_14246,N_14309);
xnor U14510 (N_14510,N_14315,N_14369);
nand U14511 (N_14511,N_14302,N_14356);
xnor U14512 (N_14512,N_14396,N_14274);
nor U14513 (N_14513,N_14298,N_14321);
xnor U14514 (N_14514,N_14356,N_14374);
nor U14515 (N_14515,N_14349,N_14305);
nor U14516 (N_14516,N_14280,N_14349);
nand U14517 (N_14517,N_14301,N_14295);
and U14518 (N_14518,N_14399,N_14250);
xor U14519 (N_14519,N_14207,N_14327);
nor U14520 (N_14520,N_14280,N_14255);
nand U14521 (N_14521,N_14398,N_14328);
nor U14522 (N_14522,N_14362,N_14288);
nor U14523 (N_14523,N_14294,N_14359);
and U14524 (N_14524,N_14291,N_14268);
nand U14525 (N_14525,N_14345,N_14349);
nand U14526 (N_14526,N_14293,N_14371);
nand U14527 (N_14527,N_14296,N_14313);
or U14528 (N_14528,N_14220,N_14370);
or U14529 (N_14529,N_14371,N_14242);
or U14530 (N_14530,N_14320,N_14217);
nand U14531 (N_14531,N_14393,N_14280);
or U14532 (N_14532,N_14356,N_14328);
nand U14533 (N_14533,N_14354,N_14259);
nand U14534 (N_14534,N_14232,N_14250);
and U14535 (N_14535,N_14354,N_14269);
or U14536 (N_14536,N_14267,N_14395);
nor U14537 (N_14537,N_14281,N_14250);
nand U14538 (N_14538,N_14200,N_14393);
or U14539 (N_14539,N_14343,N_14372);
nand U14540 (N_14540,N_14388,N_14363);
xnor U14541 (N_14541,N_14272,N_14254);
xor U14542 (N_14542,N_14326,N_14353);
and U14543 (N_14543,N_14307,N_14235);
and U14544 (N_14544,N_14273,N_14390);
and U14545 (N_14545,N_14261,N_14365);
xor U14546 (N_14546,N_14385,N_14297);
and U14547 (N_14547,N_14366,N_14267);
or U14548 (N_14548,N_14344,N_14363);
or U14549 (N_14549,N_14236,N_14210);
nand U14550 (N_14550,N_14359,N_14397);
nor U14551 (N_14551,N_14211,N_14313);
or U14552 (N_14552,N_14361,N_14248);
nor U14553 (N_14553,N_14227,N_14365);
and U14554 (N_14554,N_14295,N_14205);
xnor U14555 (N_14555,N_14312,N_14384);
xor U14556 (N_14556,N_14205,N_14329);
and U14557 (N_14557,N_14249,N_14397);
and U14558 (N_14558,N_14330,N_14381);
or U14559 (N_14559,N_14262,N_14266);
and U14560 (N_14560,N_14396,N_14240);
nor U14561 (N_14561,N_14395,N_14229);
nor U14562 (N_14562,N_14394,N_14378);
and U14563 (N_14563,N_14255,N_14245);
nand U14564 (N_14564,N_14399,N_14214);
nor U14565 (N_14565,N_14279,N_14328);
xor U14566 (N_14566,N_14251,N_14235);
xor U14567 (N_14567,N_14338,N_14390);
xnor U14568 (N_14568,N_14233,N_14390);
or U14569 (N_14569,N_14233,N_14245);
xnor U14570 (N_14570,N_14301,N_14296);
and U14571 (N_14571,N_14323,N_14297);
and U14572 (N_14572,N_14240,N_14273);
nand U14573 (N_14573,N_14375,N_14366);
nor U14574 (N_14574,N_14322,N_14319);
or U14575 (N_14575,N_14239,N_14200);
nand U14576 (N_14576,N_14349,N_14355);
nor U14577 (N_14577,N_14254,N_14306);
or U14578 (N_14578,N_14214,N_14323);
or U14579 (N_14579,N_14382,N_14305);
nand U14580 (N_14580,N_14293,N_14300);
or U14581 (N_14581,N_14389,N_14261);
and U14582 (N_14582,N_14258,N_14326);
nand U14583 (N_14583,N_14296,N_14384);
xnor U14584 (N_14584,N_14231,N_14338);
xnor U14585 (N_14585,N_14235,N_14316);
or U14586 (N_14586,N_14340,N_14333);
xnor U14587 (N_14587,N_14284,N_14396);
nor U14588 (N_14588,N_14232,N_14237);
nor U14589 (N_14589,N_14233,N_14284);
and U14590 (N_14590,N_14305,N_14390);
nor U14591 (N_14591,N_14315,N_14234);
xnor U14592 (N_14592,N_14287,N_14324);
nand U14593 (N_14593,N_14328,N_14235);
or U14594 (N_14594,N_14277,N_14357);
or U14595 (N_14595,N_14228,N_14260);
nor U14596 (N_14596,N_14257,N_14260);
xnor U14597 (N_14597,N_14215,N_14242);
nor U14598 (N_14598,N_14337,N_14366);
xnor U14599 (N_14599,N_14392,N_14324);
xor U14600 (N_14600,N_14475,N_14413);
nand U14601 (N_14601,N_14449,N_14514);
nor U14602 (N_14602,N_14498,N_14567);
nor U14603 (N_14603,N_14452,N_14402);
nor U14604 (N_14604,N_14454,N_14532);
nor U14605 (N_14605,N_14459,N_14448);
xor U14606 (N_14606,N_14505,N_14584);
and U14607 (N_14607,N_14483,N_14519);
or U14608 (N_14608,N_14463,N_14527);
nand U14609 (N_14609,N_14491,N_14574);
xor U14610 (N_14610,N_14588,N_14530);
and U14611 (N_14611,N_14553,N_14556);
xnor U14612 (N_14612,N_14453,N_14548);
nor U14613 (N_14613,N_14416,N_14470);
nand U14614 (N_14614,N_14580,N_14420);
and U14615 (N_14615,N_14562,N_14407);
or U14616 (N_14616,N_14460,N_14433);
xor U14617 (N_14617,N_14465,N_14594);
or U14618 (N_14618,N_14510,N_14440);
nor U14619 (N_14619,N_14559,N_14573);
and U14620 (N_14620,N_14474,N_14587);
nor U14621 (N_14621,N_14598,N_14578);
and U14622 (N_14622,N_14495,N_14401);
xnor U14623 (N_14623,N_14496,N_14541);
xnor U14624 (N_14624,N_14473,N_14482);
and U14625 (N_14625,N_14409,N_14512);
nor U14626 (N_14626,N_14434,N_14583);
nor U14627 (N_14627,N_14403,N_14568);
nor U14628 (N_14628,N_14447,N_14599);
xnor U14629 (N_14629,N_14400,N_14561);
nand U14630 (N_14630,N_14435,N_14517);
or U14631 (N_14631,N_14456,N_14551);
xnor U14632 (N_14632,N_14441,N_14446);
xnor U14633 (N_14633,N_14444,N_14570);
nand U14634 (N_14634,N_14471,N_14438);
or U14635 (N_14635,N_14589,N_14513);
xor U14636 (N_14636,N_14545,N_14537);
xor U14637 (N_14637,N_14515,N_14468);
nand U14638 (N_14638,N_14565,N_14560);
and U14639 (N_14639,N_14550,N_14597);
and U14640 (N_14640,N_14536,N_14552);
nand U14641 (N_14641,N_14404,N_14442);
or U14642 (N_14642,N_14466,N_14430);
or U14643 (N_14643,N_14557,N_14581);
or U14644 (N_14644,N_14543,N_14590);
or U14645 (N_14645,N_14477,N_14423);
or U14646 (N_14646,N_14539,N_14542);
nand U14647 (N_14647,N_14439,N_14503);
xor U14648 (N_14648,N_14418,N_14526);
and U14649 (N_14649,N_14502,N_14585);
xnor U14650 (N_14650,N_14408,N_14499);
nand U14651 (N_14651,N_14500,N_14546);
or U14652 (N_14652,N_14428,N_14533);
xor U14653 (N_14653,N_14489,N_14593);
nor U14654 (N_14654,N_14436,N_14501);
xor U14655 (N_14655,N_14410,N_14595);
and U14656 (N_14656,N_14535,N_14476);
nor U14657 (N_14657,N_14531,N_14412);
nand U14658 (N_14658,N_14432,N_14571);
or U14659 (N_14659,N_14467,N_14455);
nor U14660 (N_14660,N_14511,N_14576);
nand U14661 (N_14661,N_14591,N_14586);
or U14662 (N_14662,N_14529,N_14426);
or U14663 (N_14663,N_14480,N_14525);
and U14664 (N_14664,N_14509,N_14577);
xnor U14665 (N_14665,N_14523,N_14528);
and U14666 (N_14666,N_14522,N_14461);
or U14667 (N_14667,N_14469,N_14566);
or U14668 (N_14668,N_14544,N_14554);
nand U14669 (N_14669,N_14485,N_14555);
or U14670 (N_14670,N_14445,N_14437);
and U14671 (N_14671,N_14479,N_14596);
nand U14672 (N_14672,N_14582,N_14406);
or U14673 (N_14673,N_14487,N_14464);
nor U14674 (N_14674,N_14457,N_14431);
xnor U14675 (N_14675,N_14488,N_14427);
nor U14676 (N_14676,N_14572,N_14486);
or U14677 (N_14677,N_14419,N_14425);
nand U14678 (N_14678,N_14506,N_14478);
and U14679 (N_14679,N_14472,N_14429);
nand U14680 (N_14680,N_14450,N_14504);
or U14681 (N_14681,N_14524,N_14462);
and U14682 (N_14682,N_14424,N_14492);
xnor U14683 (N_14683,N_14414,N_14508);
or U14684 (N_14684,N_14518,N_14516);
nand U14685 (N_14685,N_14411,N_14538);
nand U14686 (N_14686,N_14481,N_14417);
nand U14687 (N_14687,N_14415,N_14520);
xnor U14688 (N_14688,N_14497,N_14458);
nor U14689 (N_14689,N_14549,N_14422);
nand U14690 (N_14690,N_14569,N_14521);
nor U14691 (N_14691,N_14592,N_14494);
nand U14692 (N_14692,N_14547,N_14563);
and U14693 (N_14693,N_14421,N_14443);
and U14694 (N_14694,N_14405,N_14451);
and U14695 (N_14695,N_14493,N_14490);
nand U14696 (N_14696,N_14534,N_14575);
nand U14697 (N_14697,N_14540,N_14507);
nand U14698 (N_14698,N_14558,N_14579);
or U14699 (N_14699,N_14484,N_14564);
xnor U14700 (N_14700,N_14568,N_14590);
nand U14701 (N_14701,N_14520,N_14599);
nand U14702 (N_14702,N_14412,N_14409);
nor U14703 (N_14703,N_14410,N_14400);
or U14704 (N_14704,N_14509,N_14427);
nand U14705 (N_14705,N_14469,N_14498);
nand U14706 (N_14706,N_14412,N_14406);
nor U14707 (N_14707,N_14470,N_14433);
nor U14708 (N_14708,N_14581,N_14411);
or U14709 (N_14709,N_14490,N_14451);
nor U14710 (N_14710,N_14425,N_14415);
nand U14711 (N_14711,N_14572,N_14468);
nand U14712 (N_14712,N_14544,N_14430);
or U14713 (N_14713,N_14541,N_14464);
or U14714 (N_14714,N_14528,N_14461);
nor U14715 (N_14715,N_14452,N_14485);
nand U14716 (N_14716,N_14503,N_14485);
and U14717 (N_14717,N_14503,N_14467);
nor U14718 (N_14718,N_14554,N_14440);
or U14719 (N_14719,N_14576,N_14553);
and U14720 (N_14720,N_14475,N_14448);
xnor U14721 (N_14721,N_14478,N_14527);
and U14722 (N_14722,N_14529,N_14565);
nor U14723 (N_14723,N_14441,N_14404);
nand U14724 (N_14724,N_14507,N_14480);
xnor U14725 (N_14725,N_14512,N_14443);
nor U14726 (N_14726,N_14485,N_14537);
nor U14727 (N_14727,N_14432,N_14491);
nor U14728 (N_14728,N_14564,N_14500);
or U14729 (N_14729,N_14401,N_14434);
or U14730 (N_14730,N_14406,N_14455);
xor U14731 (N_14731,N_14508,N_14462);
nor U14732 (N_14732,N_14576,N_14571);
nand U14733 (N_14733,N_14523,N_14556);
xor U14734 (N_14734,N_14444,N_14565);
nor U14735 (N_14735,N_14544,N_14577);
and U14736 (N_14736,N_14409,N_14407);
xor U14737 (N_14737,N_14478,N_14569);
nor U14738 (N_14738,N_14572,N_14542);
nand U14739 (N_14739,N_14557,N_14520);
nor U14740 (N_14740,N_14443,N_14423);
xor U14741 (N_14741,N_14583,N_14447);
xor U14742 (N_14742,N_14522,N_14434);
nor U14743 (N_14743,N_14556,N_14454);
nand U14744 (N_14744,N_14514,N_14501);
and U14745 (N_14745,N_14584,N_14496);
xor U14746 (N_14746,N_14577,N_14479);
nor U14747 (N_14747,N_14598,N_14524);
and U14748 (N_14748,N_14424,N_14462);
xnor U14749 (N_14749,N_14501,N_14443);
xnor U14750 (N_14750,N_14563,N_14478);
nor U14751 (N_14751,N_14491,N_14503);
nor U14752 (N_14752,N_14477,N_14435);
nor U14753 (N_14753,N_14483,N_14568);
or U14754 (N_14754,N_14531,N_14474);
nor U14755 (N_14755,N_14473,N_14488);
nor U14756 (N_14756,N_14448,N_14584);
and U14757 (N_14757,N_14546,N_14543);
xnor U14758 (N_14758,N_14414,N_14443);
nor U14759 (N_14759,N_14565,N_14554);
nand U14760 (N_14760,N_14487,N_14576);
and U14761 (N_14761,N_14509,N_14567);
or U14762 (N_14762,N_14412,N_14503);
and U14763 (N_14763,N_14444,N_14503);
nor U14764 (N_14764,N_14553,N_14591);
or U14765 (N_14765,N_14455,N_14430);
xnor U14766 (N_14766,N_14505,N_14477);
xnor U14767 (N_14767,N_14434,N_14525);
nor U14768 (N_14768,N_14407,N_14583);
nand U14769 (N_14769,N_14415,N_14454);
or U14770 (N_14770,N_14478,N_14553);
nor U14771 (N_14771,N_14425,N_14498);
nand U14772 (N_14772,N_14405,N_14545);
or U14773 (N_14773,N_14491,N_14523);
nor U14774 (N_14774,N_14540,N_14483);
nor U14775 (N_14775,N_14453,N_14473);
and U14776 (N_14776,N_14510,N_14465);
xnor U14777 (N_14777,N_14423,N_14449);
xor U14778 (N_14778,N_14547,N_14565);
and U14779 (N_14779,N_14419,N_14541);
nor U14780 (N_14780,N_14521,N_14430);
xor U14781 (N_14781,N_14456,N_14584);
or U14782 (N_14782,N_14595,N_14474);
nor U14783 (N_14783,N_14423,N_14539);
nand U14784 (N_14784,N_14486,N_14548);
xnor U14785 (N_14785,N_14499,N_14581);
and U14786 (N_14786,N_14503,N_14463);
nand U14787 (N_14787,N_14598,N_14557);
xor U14788 (N_14788,N_14454,N_14553);
or U14789 (N_14789,N_14526,N_14424);
or U14790 (N_14790,N_14442,N_14441);
or U14791 (N_14791,N_14479,N_14569);
xnor U14792 (N_14792,N_14510,N_14512);
xor U14793 (N_14793,N_14462,N_14584);
nor U14794 (N_14794,N_14555,N_14501);
xnor U14795 (N_14795,N_14495,N_14503);
xnor U14796 (N_14796,N_14425,N_14574);
nor U14797 (N_14797,N_14543,N_14411);
nand U14798 (N_14798,N_14458,N_14496);
or U14799 (N_14799,N_14569,N_14482);
xor U14800 (N_14800,N_14722,N_14791);
or U14801 (N_14801,N_14797,N_14701);
nor U14802 (N_14802,N_14761,N_14643);
nand U14803 (N_14803,N_14630,N_14624);
or U14804 (N_14804,N_14638,N_14762);
nor U14805 (N_14805,N_14648,N_14778);
nor U14806 (N_14806,N_14769,N_14719);
and U14807 (N_14807,N_14755,N_14759);
nand U14808 (N_14808,N_14718,N_14772);
xnor U14809 (N_14809,N_14716,N_14708);
xor U14810 (N_14810,N_14647,N_14682);
xnor U14811 (N_14811,N_14736,N_14729);
xnor U14812 (N_14812,N_14745,N_14608);
or U14813 (N_14813,N_14795,N_14656);
xor U14814 (N_14814,N_14724,N_14607);
nand U14815 (N_14815,N_14730,N_14625);
or U14816 (N_14816,N_14785,N_14715);
xnor U14817 (N_14817,N_14694,N_14788);
nand U14818 (N_14818,N_14734,N_14726);
or U14819 (N_14819,N_14634,N_14741);
or U14820 (N_14820,N_14672,N_14752);
xnor U14821 (N_14821,N_14668,N_14602);
xor U14822 (N_14822,N_14646,N_14664);
nand U14823 (N_14823,N_14702,N_14740);
or U14824 (N_14824,N_14700,N_14766);
nor U14825 (N_14825,N_14774,N_14738);
nor U14826 (N_14826,N_14603,N_14787);
nand U14827 (N_14827,N_14721,N_14620);
nand U14828 (N_14828,N_14720,N_14610);
nor U14829 (N_14829,N_14675,N_14688);
or U14830 (N_14830,N_14611,N_14616);
xnor U14831 (N_14831,N_14784,N_14771);
xnor U14832 (N_14832,N_14711,N_14757);
nand U14833 (N_14833,N_14696,N_14677);
or U14834 (N_14834,N_14650,N_14614);
or U14835 (N_14835,N_14739,N_14623);
xnor U14836 (N_14836,N_14636,N_14793);
nand U14837 (N_14837,N_14657,N_14663);
and U14838 (N_14838,N_14669,N_14644);
and U14839 (N_14839,N_14645,N_14605);
and U14840 (N_14840,N_14737,N_14794);
xor U14841 (N_14841,N_14615,N_14609);
nand U14842 (N_14842,N_14728,N_14698);
and U14843 (N_14843,N_14622,N_14765);
nand U14844 (N_14844,N_14747,N_14627);
nor U14845 (N_14845,N_14786,N_14689);
nand U14846 (N_14846,N_14764,N_14684);
nor U14847 (N_14847,N_14683,N_14735);
or U14848 (N_14848,N_14639,N_14662);
or U14849 (N_14849,N_14732,N_14604);
xor U14850 (N_14850,N_14706,N_14796);
nand U14851 (N_14851,N_14792,N_14709);
nor U14852 (N_14852,N_14779,N_14703);
or U14853 (N_14853,N_14789,N_14676);
xnor U14854 (N_14854,N_14691,N_14723);
or U14855 (N_14855,N_14613,N_14748);
or U14856 (N_14856,N_14742,N_14665);
xnor U14857 (N_14857,N_14628,N_14758);
xor U14858 (N_14858,N_14621,N_14799);
xor U14859 (N_14859,N_14685,N_14617);
nor U14860 (N_14860,N_14775,N_14606);
nor U14861 (N_14861,N_14712,N_14690);
nor U14862 (N_14862,N_14670,N_14798);
nand U14863 (N_14863,N_14714,N_14781);
nand U14864 (N_14864,N_14653,N_14746);
and U14865 (N_14865,N_14705,N_14717);
or U14866 (N_14866,N_14671,N_14654);
xnor U14867 (N_14867,N_14743,N_14680);
or U14868 (N_14868,N_14655,N_14629);
nand U14869 (N_14869,N_14626,N_14649);
nand U14870 (N_14870,N_14707,N_14658);
and U14871 (N_14871,N_14601,N_14780);
or U14872 (N_14872,N_14635,N_14753);
or U14873 (N_14873,N_14699,N_14697);
nor U14874 (N_14874,N_14632,N_14618);
xnor U14875 (N_14875,N_14763,N_14612);
xor U14876 (N_14876,N_14686,N_14756);
and U14877 (N_14877,N_14600,N_14777);
or U14878 (N_14878,N_14687,N_14681);
or U14879 (N_14879,N_14750,N_14704);
xor U14880 (N_14880,N_14782,N_14674);
nand U14881 (N_14881,N_14733,N_14790);
and U14882 (N_14882,N_14661,N_14673);
nand U14883 (N_14883,N_14710,N_14783);
or U14884 (N_14884,N_14751,N_14749);
xor U14885 (N_14885,N_14659,N_14693);
xor U14886 (N_14886,N_14633,N_14744);
and U14887 (N_14887,N_14660,N_14642);
and U14888 (N_14888,N_14768,N_14727);
xnor U14889 (N_14889,N_14713,N_14695);
and U14890 (N_14890,N_14770,N_14725);
nor U14891 (N_14891,N_14651,N_14652);
and U14892 (N_14892,N_14678,N_14640);
or U14893 (N_14893,N_14760,N_14666);
xor U14894 (N_14894,N_14767,N_14679);
xor U14895 (N_14895,N_14776,N_14631);
xor U14896 (N_14896,N_14641,N_14773);
and U14897 (N_14897,N_14667,N_14637);
and U14898 (N_14898,N_14619,N_14731);
nand U14899 (N_14899,N_14692,N_14754);
nand U14900 (N_14900,N_14611,N_14718);
nand U14901 (N_14901,N_14747,N_14635);
and U14902 (N_14902,N_14660,N_14762);
or U14903 (N_14903,N_14696,N_14644);
and U14904 (N_14904,N_14773,N_14717);
nor U14905 (N_14905,N_14632,N_14705);
and U14906 (N_14906,N_14772,N_14790);
nand U14907 (N_14907,N_14794,N_14620);
nor U14908 (N_14908,N_14669,N_14702);
xnor U14909 (N_14909,N_14671,N_14754);
and U14910 (N_14910,N_14773,N_14659);
nand U14911 (N_14911,N_14694,N_14690);
and U14912 (N_14912,N_14607,N_14789);
nor U14913 (N_14913,N_14728,N_14694);
or U14914 (N_14914,N_14760,N_14701);
xor U14915 (N_14915,N_14741,N_14703);
nor U14916 (N_14916,N_14616,N_14727);
nand U14917 (N_14917,N_14652,N_14663);
and U14918 (N_14918,N_14755,N_14686);
nand U14919 (N_14919,N_14684,N_14734);
and U14920 (N_14920,N_14740,N_14788);
or U14921 (N_14921,N_14775,N_14634);
nor U14922 (N_14922,N_14646,N_14715);
nor U14923 (N_14923,N_14772,N_14624);
xor U14924 (N_14924,N_14630,N_14765);
or U14925 (N_14925,N_14725,N_14636);
nor U14926 (N_14926,N_14705,N_14635);
and U14927 (N_14927,N_14796,N_14630);
nor U14928 (N_14928,N_14668,N_14715);
xor U14929 (N_14929,N_14779,N_14657);
xor U14930 (N_14930,N_14704,N_14758);
nand U14931 (N_14931,N_14768,N_14615);
or U14932 (N_14932,N_14680,N_14770);
xor U14933 (N_14933,N_14714,N_14733);
xor U14934 (N_14934,N_14608,N_14756);
or U14935 (N_14935,N_14687,N_14675);
nor U14936 (N_14936,N_14787,N_14742);
nor U14937 (N_14937,N_14757,N_14730);
nor U14938 (N_14938,N_14768,N_14750);
nor U14939 (N_14939,N_14656,N_14704);
or U14940 (N_14940,N_14721,N_14660);
xnor U14941 (N_14941,N_14601,N_14747);
and U14942 (N_14942,N_14639,N_14641);
or U14943 (N_14943,N_14614,N_14610);
nor U14944 (N_14944,N_14733,N_14698);
nor U14945 (N_14945,N_14769,N_14782);
and U14946 (N_14946,N_14739,N_14744);
nor U14947 (N_14947,N_14693,N_14676);
and U14948 (N_14948,N_14631,N_14652);
xor U14949 (N_14949,N_14699,N_14664);
nor U14950 (N_14950,N_14723,N_14703);
xnor U14951 (N_14951,N_14682,N_14776);
xor U14952 (N_14952,N_14730,N_14754);
nand U14953 (N_14953,N_14672,N_14637);
and U14954 (N_14954,N_14675,N_14667);
xnor U14955 (N_14955,N_14699,N_14746);
or U14956 (N_14956,N_14793,N_14702);
xor U14957 (N_14957,N_14631,N_14620);
nand U14958 (N_14958,N_14799,N_14749);
nor U14959 (N_14959,N_14678,N_14643);
or U14960 (N_14960,N_14769,N_14658);
nand U14961 (N_14961,N_14792,N_14687);
nand U14962 (N_14962,N_14689,N_14692);
or U14963 (N_14963,N_14744,N_14680);
nor U14964 (N_14964,N_14666,N_14739);
xor U14965 (N_14965,N_14638,N_14618);
nand U14966 (N_14966,N_14704,N_14770);
or U14967 (N_14967,N_14704,N_14759);
nand U14968 (N_14968,N_14732,N_14645);
nand U14969 (N_14969,N_14609,N_14725);
and U14970 (N_14970,N_14767,N_14790);
nand U14971 (N_14971,N_14704,N_14689);
nand U14972 (N_14972,N_14602,N_14798);
xor U14973 (N_14973,N_14674,N_14693);
xor U14974 (N_14974,N_14664,N_14641);
nand U14975 (N_14975,N_14663,N_14613);
xnor U14976 (N_14976,N_14772,N_14646);
xor U14977 (N_14977,N_14753,N_14737);
or U14978 (N_14978,N_14798,N_14632);
or U14979 (N_14979,N_14759,N_14639);
xor U14980 (N_14980,N_14718,N_14659);
xor U14981 (N_14981,N_14768,N_14630);
and U14982 (N_14982,N_14718,N_14696);
nand U14983 (N_14983,N_14616,N_14769);
xnor U14984 (N_14984,N_14645,N_14619);
nand U14985 (N_14985,N_14614,N_14789);
nor U14986 (N_14986,N_14772,N_14677);
or U14987 (N_14987,N_14691,N_14646);
xnor U14988 (N_14988,N_14673,N_14731);
or U14989 (N_14989,N_14675,N_14655);
and U14990 (N_14990,N_14660,N_14728);
nor U14991 (N_14991,N_14705,N_14641);
nand U14992 (N_14992,N_14798,N_14623);
and U14993 (N_14993,N_14796,N_14635);
and U14994 (N_14994,N_14684,N_14698);
and U14995 (N_14995,N_14602,N_14797);
and U14996 (N_14996,N_14700,N_14634);
xnor U14997 (N_14997,N_14743,N_14771);
and U14998 (N_14998,N_14759,N_14763);
or U14999 (N_14999,N_14645,N_14609);
nand U15000 (N_15000,N_14882,N_14802);
or U15001 (N_15001,N_14954,N_14889);
and U15002 (N_15002,N_14934,N_14881);
nor U15003 (N_15003,N_14839,N_14949);
nor U15004 (N_15004,N_14969,N_14824);
and U15005 (N_15005,N_14885,N_14847);
nand U15006 (N_15006,N_14870,N_14876);
or U15007 (N_15007,N_14859,N_14912);
xnor U15008 (N_15008,N_14937,N_14895);
and U15009 (N_15009,N_14922,N_14932);
or U15010 (N_15010,N_14942,N_14936);
nand U15011 (N_15011,N_14930,N_14967);
xnor U15012 (N_15012,N_14975,N_14990);
nand U15013 (N_15013,N_14856,N_14863);
nand U15014 (N_15014,N_14901,N_14924);
nand U15015 (N_15015,N_14872,N_14846);
or U15016 (N_15016,N_14943,N_14928);
xor U15017 (N_15017,N_14807,N_14850);
or U15018 (N_15018,N_14945,N_14997);
nand U15019 (N_15019,N_14831,N_14985);
xnor U15020 (N_15020,N_14820,N_14965);
or U15021 (N_15021,N_14808,N_14981);
or U15022 (N_15022,N_14804,N_14926);
or U15023 (N_15023,N_14995,N_14964);
nand U15024 (N_15024,N_14857,N_14869);
nor U15025 (N_15025,N_14817,N_14883);
or U15026 (N_15026,N_14845,N_14933);
and U15027 (N_15027,N_14812,N_14991);
nor U15028 (N_15028,N_14838,N_14830);
or U15029 (N_15029,N_14993,N_14871);
nand U15030 (N_15030,N_14987,N_14904);
xnor U15031 (N_15031,N_14910,N_14874);
or U15032 (N_15032,N_14955,N_14862);
xor U15033 (N_15033,N_14832,N_14966);
xor U15034 (N_15034,N_14849,N_14815);
or U15035 (N_15035,N_14896,N_14983);
or U15036 (N_15036,N_14984,N_14880);
nand U15037 (N_15037,N_14890,N_14811);
and U15038 (N_15038,N_14829,N_14888);
xnor U15039 (N_15039,N_14826,N_14897);
and U15040 (N_15040,N_14810,N_14825);
nor U15041 (N_15041,N_14900,N_14854);
nor U15042 (N_15042,N_14914,N_14877);
and U15043 (N_15043,N_14822,N_14861);
nor U15044 (N_15044,N_14913,N_14858);
nor U15045 (N_15045,N_14931,N_14974);
and U15046 (N_15046,N_14918,N_14844);
xnor U15047 (N_15047,N_14879,N_14827);
or U15048 (N_15048,N_14868,N_14961);
nor U15049 (N_15049,N_14968,N_14988);
xnor U15050 (N_15050,N_14873,N_14977);
or U15051 (N_15051,N_14905,N_14999);
or U15052 (N_15052,N_14998,N_14842);
and U15053 (N_15053,N_14853,N_14814);
and U15054 (N_15054,N_14894,N_14806);
xnor U15055 (N_15055,N_14833,N_14892);
and U15056 (N_15056,N_14986,N_14944);
nand U15057 (N_15057,N_14891,N_14927);
nor U15058 (N_15058,N_14813,N_14976);
xor U15059 (N_15059,N_14925,N_14818);
or U15060 (N_15060,N_14941,N_14970);
nor U15061 (N_15061,N_14855,N_14851);
and U15062 (N_15062,N_14887,N_14956);
nand U15063 (N_15063,N_14886,N_14982);
nor U15064 (N_15064,N_14948,N_14898);
nand U15065 (N_15065,N_14803,N_14920);
nand U15066 (N_15066,N_14963,N_14950);
or U15067 (N_15067,N_14878,N_14951);
xor U15068 (N_15068,N_14805,N_14903);
nand U15069 (N_15069,N_14908,N_14801);
or U15070 (N_15070,N_14837,N_14836);
nand U15071 (N_15071,N_14989,N_14958);
nand U15072 (N_15072,N_14940,N_14972);
nand U15073 (N_15073,N_14841,N_14800);
nand U15074 (N_15074,N_14909,N_14907);
nor U15075 (N_15075,N_14921,N_14884);
or U15076 (N_15076,N_14959,N_14902);
or U15077 (N_15077,N_14980,N_14971);
or U15078 (N_15078,N_14865,N_14979);
nor U15079 (N_15079,N_14875,N_14821);
or U15080 (N_15080,N_14819,N_14962);
xnor U15081 (N_15081,N_14866,N_14992);
nand U15082 (N_15082,N_14952,N_14834);
xor U15083 (N_15083,N_14867,N_14860);
and U15084 (N_15084,N_14828,N_14816);
nor U15085 (N_15085,N_14953,N_14923);
xnor U15086 (N_15086,N_14947,N_14929);
xor U15087 (N_15087,N_14996,N_14899);
and U15088 (N_15088,N_14893,N_14978);
and U15089 (N_15089,N_14911,N_14916);
nand U15090 (N_15090,N_14994,N_14935);
nand U15091 (N_15091,N_14946,N_14915);
or U15092 (N_15092,N_14848,N_14852);
and U15093 (N_15093,N_14960,N_14919);
nand U15094 (N_15094,N_14957,N_14938);
xor U15095 (N_15095,N_14823,N_14840);
and U15096 (N_15096,N_14973,N_14939);
and U15097 (N_15097,N_14864,N_14835);
xor U15098 (N_15098,N_14917,N_14843);
or U15099 (N_15099,N_14906,N_14809);
or U15100 (N_15100,N_14819,N_14924);
xor U15101 (N_15101,N_14911,N_14956);
and U15102 (N_15102,N_14997,N_14907);
and U15103 (N_15103,N_14947,N_14973);
and U15104 (N_15104,N_14817,N_14853);
or U15105 (N_15105,N_14972,N_14881);
xnor U15106 (N_15106,N_14824,N_14945);
nor U15107 (N_15107,N_14836,N_14819);
nor U15108 (N_15108,N_14953,N_14935);
nor U15109 (N_15109,N_14845,N_14985);
nand U15110 (N_15110,N_14982,N_14848);
nand U15111 (N_15111,N_14987,N_14860);
nand U15112 (N_15112,N_14831,N_14871);
nor U15113 (N_15113,N_14801,N_14879);
and U15114 (N_15114,N_14919,N_14830);
and U15115 (N_15115,N_14907,N_14934);
or U15116 (N_15116,N_14845,N_14817);
and U15117 (N_15117,N_14858,N_14911);
nor U15118 (N_15118,N_14817,N_14941);
and U15119 (N_15119,N_14892,N_14942);
or U15120 (N_15120,N_14925,N_14971);
or U15121 (N_15121,N_14919,N_14882);
and U15122 (N_15122,N_14811,N_14924);
or U15123 (N_15123,N_14832,N_14946);
nor U15124 (N_15124,N_14801,N_14954);
or U15125 (N_15125,N_14859,N_14869);
and U15126 (N_15126,N_14898,N_14943);
or U15127 (N_15127,N_14866,N_14822);
and U15128 (N_15128,N_14999,N_14875);
xor U15129 (N_15129,N_14816,N_14977);
and U15130 (N_15130,N_14929,N_14984);
xor U15131 (N_15131,N_14855,N_14920);
nand U15132 (N_15132,N_14964,N_14942);
nor U15133 (N_15133,N_14971,N_14943);
nand U15134 (N_15134,N_14882,N_14930);
xnor U15135 (N_15135,N_14996,N_14833);
nand U15136 (N_15136,N_14981,N_14850);
xnor U15137 (N_15137,N_14917,N_14828);
xnor U15138 (N_15138,N_14852,N_14902);
nand U15139 (N_15139,N_14838,N_14930);
or U15140 (N_15140,N_14965,N_14838);
xnor U15141 (N_15141,N_14918,N_14853);
or U15142 (N_15142,N_14888,N_14881);
nand U15143 (N_15143,N_14911,N_14874);
nor U15144 (N_15144,N_14890,N_14833);
nand U15145 (N_15145,N_14973,N_14866);
nor U15146 (N_15146,N_14873,N_14985);
nor U15147 (N_15147,N_14848,N_14941);
and U15148 (N_15148,N_14839,N_14902);
or U15149 (N_15149,N_14932,N_14848);
and U15150 (N_15150,N_14847,N_14824);
xnor U15151 (N_15151,N_14980,N_14808);
or U15152 (N_15152,N_14915,N_14912);
and U15153 (N_15153,N_14983,N_14862);
xor U15154 (N_15154,N_14877,N_14929);
nand U15155 (N_15155,N_14937,N_14978);
or U15156 (N_15156,N_14921,N_14959);
or U15157 (N_15157,N_14809,N_14931);
or U15158 (N_15158,N_14976,N_14978);
or U15159 (N_15159,N_14880,N_14892);
nor U15160 (N_15160,N_14970,N_14992);
nor U15161 (N_15161,N_14954,N_14845);
nand U15162 (N_15162,N_14920,N_14992);
or U15163 (N_15163,N_14945,N_14955);
or U15164 (N_15164,N_14938,N_14880);
nor U15165 (N_15165,N_14926,N_14833);
and U15166 (N_15166,N_14911,N_14834);
nor U15167 (N_15167,N_14836,N_14811);
xnor U15168 (N_15168,N_14817,N_14977);
or U15169 (N_15169,N_14832,N_14973);
nor U15170 (N_15170,N_14952,N_14891);
nor U15171 (N_15171,N_14828,N_14931);
nand U15172 (N_15172,N_14908,N_14951);
nand U15173 (N_15173,N_14894,N_14906);
and U15174 (N_15174,N_14800,N_14934);
nand U15175 (N_15175,N_14912,N_14911);
and U15176 (N_15176,N_14906,N_14997);
nand U15177 (N_15177,N_14823,N_14901);
nand U15178 (N_15178,N_14821,N_14850);
nor U15179 (N_15179,N_14899,N_14894);
and U15180 (N_15180,N_14928,N_14994);
or U15181 (N_15181,N_14872,N_14949);
and U15182 (N_15182,N_14963,N_14946);
and U15183 (N_15183,N_14841,N_14869);
nand U15184 (N_15184,N_14800,N_14900);
xor U15185 (N_15185,N_14980,N_14894);
nor U15186 (N_15186,N_14989,N_14930);
and U15187 (N_15187,N_14856,N_14808);
and U15188 (N_15188,N_14808,N_14960);
and U15189 (N_15189,N_14975,N_14865);
xnor U15190 (N_15190,N_14974,N_14897);
nand U15191 (N_15191,N_14880,N_14813);
and U15192 (N_15192,N_14931,N_14906);
xnor U15193 (N_15193,N_14810,N_14945);
and U15194 (N_15194,N_14967,N_14945);
nor U15195 (N_15195,N_14889,N_14894);
xnor U15196 (N_15196,N_14952,N_14959);
or U15197 (N_15197,N_14832,N_14887);
and U15198 (N_15198,N_14841,N_14901);
nand U15199 (N_15199,N_14897,N_14867);
nand U15200 (N_15200,N_15182,N_15083);
or U15201 (N_15201,N_15048,N_15062);
and U15202 (N_15202,N_15154,N_15135);
xor U15203 (N_15203,N_15053,N_15027);
and U15204 (N_15204,N_15005,N_15037);
xnor U15205 (N_15205,N_15124,N_15078);
nor U15206 (N_15206,N_15186,N_15009);
or U15207 (N_15207,N_15107,N_15011);
or U15208 (N_15208,N_15170,N_15003);
nand U15209 (N_15209,N_15167,N_15125);
nand U15210 (N_15210,N_15067,N_15114);
nor U15211 (N_15211,N_15128,N_15143);
or U15212 (N_15212,N_15144,N_15150);
nand U15213 (N_15213,N_15036,N_15021);
xor U15214 (N_15214,N_15072,N_15096);
nor U15215 (N_15215,N_15134,N_15147);
and U15216 (N_15216,N_15018,N_15120);
xor U15217 (N_15217,N_15031,N_15174);
or U15218 (N_15218,N_15105,N_15051);
nand U15219 (N_15219,N_15157,N_15152);
or U15220 (N_15220,N_15195,N_15085);
or U15221 (N_15221,N_15099,N_15191);
nor U15222 (N_15222,N_15029,N_15142);
and U15223 (N_15223,N_15073,N_15104);
or U15224 (N_15224,N_15007,N_15016);
nor U15225 (N_15225,N_15022,N_15175);
or U15226 (N_15226,N_15043,N_15193);
and U15227 (N_15227,N_15102,N_15091);
or U15228 (N_15228,N_15189,N_15004);
xor U15229 (N_15229,N_15145,N_15132);
xor U15230 (N_15230,N_15086,N_15192);
nor U15231 (N_15231,N_15118,N_15041);
nor U15232 (N_15232,N_15057,N_15155);
nand U15233 (N_15233,N_15045,N_15087);
xnor U15234 (N_15234,N_15133,N_15024);
or U15235 (N_15235,N_15110,N_15071);
xnor U15236 (N_15236,N_15176,N_15017);
xor U15237 (N_15237,N_15180,N_15109);
xnor U15238 (N_15238,N_15177,N_15127);
xor U15239 (N_15239,N_15137,N_15050);
or U15240 (N_15240,N_15098,N_15034);
nand U15241 (N_15241,N_15077,N_15030);
nand U15242 (N_15242,N_15151,N_15090);
nand U15243 (N_15243,N_15093,N_15158);
or U15244 (N_15244,N_15126,N_15046);
nor U15245 (N_15245,N_15140,N_15079);
nor U15246 (N_15246,N_15089,N_15198);
xor U15247 (N_15247,N_15061,N_15012);
nand U15248 (N_15248,N_15023,N_15032);
or U15249 (N_15249,N_15117,N_15197);
and U15250 (N_15250,N_15130,N_15166);
nor U15251 (N_15251,N_15123,N_15122);
nand U15252 (N_15252,N_15076,N_15040);
nand U15253 (N_15253,N_15113,N_15172);
and U15254 (N_15254,N_15131,N_15052);
or U15255 (N_15255,N_15121,N_15000);
and U15256 (N_15256,N_15165,N_15162);
nor U15257 (N_15257,N_15138,N_15171);
or U15258 (N_15258,N_15059,N_15173);
xor U15259 (N_15259,N_15010,N_15196);
and U15260 (N_15260,N_15056,N_15035);
and U15261 (N_15261,N_15136,N_15013);
or U15262 (N_15262,N_15161,N_15070);
and U15263 (N_15263,N_15181,N_15008);
or U15264 (N_15264,N_15006,N_15178);
nor U15265 (N_15265,N_15002,N_15014);
nor U15266 (N_15266,N_15097,N_15088);
nor U15267 (N_15267,N_15156,N_15084);
nand U15268 (N_15268,N_15141,N_15163);
nand U15269 (N_15269,N_15060,N_15015);
nand U15270 (N_15270,N_15179,N_15001);
or U15271 (N_15271,N_15025,N_15075);
nand U15272 (N_15272,N_15047,N_15168);
and U15273 (N_15273,N_15054,N_15069);
nor U15274 (N_15274,N_15055,N_15074);
or U15275 (N_15275,N_15020,N_15185);
and U15276 (N_15276,N_15065,N_15183);
or U15277 (N_15277,N_15044,N_15153);
or U15278 (N_15278,N_15184,N_15080);
nor U15279 (N_15279,N_15116,N_15129);
and U15280 (N_15280,N_15188,N_15190);
and U15281 (N_15281,N_15033,N_15064);
xnor U15282 (N_15282,N_15139,N_15106);
nor U15283 (N_15283,N_15187,N_15169);
or U15284 (N_15284,N_15019,N_15199);
and U15285 (N_15285,N_15146,N_15026);
xor U15286 (N_15286,N_15095,N_15066);
nand U15287 (N_15287,N_15115,N_15094);
or U15288 (N_15288,N_15058,N_15100);
nand U15289 (N_15289,N_15049,N_15119);
and U15290 (N_15290,N_15103,N_15082);
and U15291 (N_15291,N_15194,N_15108);
nand U15292 (N_15292,N_15038,N_15101);
or U15293 (N_15293,N_15112,N_15042);
nor U15294 (N_15294,N_15111,N_15148);
xnor U15295 (N_15295,N_15063,N_15159);
nor U15296 (N_15296,N_15081,N_15068);
or U15297 (N_15297,N_15149,N_15160);
xnor U15298 (N_15298,N_15164,N_15039);
and U15299 (N_15299,N_15028,N_15092);
nand U15300 (N_15300,N_15001,N_15142);
or U15301 (N_15301,N_15171,N_15080);
or U15302 (N_15302,N_15009,N_15055);
nand U15303 (N_15303,N_15175,N_15144);
or U15304 (N_15304,N_15128,N_15112);
nand U15305 (N_15305,N_15137,N_15132);
nand U15306 (N_15306,N_15015,N_15016);
or U15307 (N_15307,N_15118,N_15197);
nand U15308 (N_15308,N_15173,N_15047);
xnor U15309 (N_15309,N_15095,N_15041);
nor U15310 (N_15310,N_15070,N_15054);
or U15311 (N_15311,N_15037,N_15197);
xnor U15312 (N_15312,N_15148,N_15136);
nor U15313 (N_15313,N_15065,N_15178);
or U15314 (N_15314,N_15078,N_15000);
xnor U15315 (N_15315,N_15162,N_15065);
nor U15316 (N_15316,N_15002,N_15036);
nor U15317 (N_15317,N_15068,N_15087);
nor U15318 (N_15318,N_15168,N_15093);
and U15319 (N_15319,N_15141,N_15090);
xnor U15320 (N_15320,N_15066,N_15087);
nor U15321 (N_15321,N_15101,N_15142);
or U15322 (N_15322,N_15119,N_15132);
xor U15323 (N_15323,N_15185,N_15116);
xnor U15324 (N_15324,N_15101,N_15058);
nor U15325 (N_15325,N_15061,N_15195);
or U15326 (N_15326,N_15059,N_15128);
nor U15327 (N_15327,N_15000,N_15050);
or U15328 (N_15328,N_15101,N_15179);
nand U15329 (N_15329,N_15128,N_15023);
xnor U15330 (N_15330,N_15002,N_15052);
xor U15331 (N_15331,N_15116,N_15067);
nand U15332 (N_15332,N_15043,N_15175);
xnor U15333 (N_15333,N_15164,N_15185);
nor U15334 (N_15334,N_15085,N_15138);
or U15335 (N_15335,N_15196,N_15136);
or U15336 (N_15336,N_15000,N_15187);
or U15337 (N_15337,N_15074,N_15180);
and U15338 (N_15338,N_15006,N_15142);
or U15339 (N_15339,N_15116,N_15040);
nor U15340 (N_15340,N_15107,N_15127);
and U15341 (N_15341,N_15188,N_15082);
and U15342 (N_15342,N_15163,N_15106);
xnor U15343 (N_15343,N_15141,N_15134);
or U15344 (N_15344,N_15002,N_15163);
and U15345 (N_15345,N_15118,N_15141);
and U15346 (N_15346,N_15130,N_15008);
xnor U15347 (N_15347,N_15139,N_15078);
and U15348 (N_15348,N_15077,N_15187);
or U15349 (N_15349,N_15031,N_15022);
xor U15350 (N_15350,N_15188,N_15043);
nand U15351 (N_15351,N_15041,N_15028);
nand U15352 (N_15352,N_15127,N_15187);
and U15353 (N_15353,N_15082,N_15087);
or U15354 (N_15354,N_15163,N_15111);
nor U15355 (N_15355,N_15135,N_15012);
nor U15356 (N_15356,N_15053,N_15104);
xor U15357 (N_15357,N_15152,N_15092);
and U15358 (N_15358,N_15036,N_15098);
xnor U15359 (N_15359,N_15122,N_15189);
nand U15360 (N_15360,N_15047,N_15137);
or U15361 (N_15361,N_15072,N_15165);
xnor U15362 (N_15362,N_15021,N_15020);
nor U15363 (N_15363,N_15076,N_15067);
nor U15364 (N_15364,N_15023,N_15005);
or U15365 (N_15365,N_15103,N_15013);
or U15366 (N_15366,N_15132,N_15161);
nand U15367 (N_15367,N_15037,N_15023);
nand U15368 (N_15368,N_15121,N_15143);
and U15369 (N_15369,N_15143,N_15075);
or U15370 (N_15370,N_15170,N_15098);
nand U15371 (N_15371,N_15156,N_15178);
and U15372 (N_15372,N_15065,N_15115);
and U15373 (N_15373,N_15136,N_15126);
nor U15374 (N_15374,N_15098,N_15050);
nand U15375 (N_15375,N_15026,N_15147);
nand U15376 (N_15376,N_15194,N_15121);
or U15377 (N_15377,N_15002,N_15069);
nor U15378 (N_15378,N_15140,N_15093);
nand U15379 (N_15379,N_15032,N_15046);
xnor U15380 (N_15380,N_15143,N_15067);
nand U15381 (N_15381,N_15195,N_15094);
xnor U15382 (N_15382,N_15002,N_15125);
or U15383 (N_15383,N_15078,N_15057);
or U15384 (N_15384,N_15129,N_15077);
nand U15385 (N_15385,N_15053,N_15013);
xnor U15386 (N_15386,N_15148,N_15079);
nand U15387 (N_15387,N_15047,N_15051);
xnor U15388 (N_15388,N_15175,N_15124);
nand U15389 (N_15389,N_15027,N_15109);
and U15390 (N_15390,N_15179,N_15008);
and U15391 (N_15391,N_15053,N_15184);
nand U15392 (N_15392,N_15143,N_15100);
or U15393 (N_15393,N_15022,N_15026);
xor U15394 (N_15394,N_15091,N_15038);
nor U15395 (N_15395,N_15178,N_15182);
xnor U15396 (N_15396,N_15002,N_15067);
nand U15397 (N_15397,N_15068,N_15067);
and U15398 (N_15398,N_15078,N_15111);
and U15399 (N_15399,N_15050,N_15073);
or U15400 (N_15400,N_15360,N_15211);
and U15401 (N_15401,N_15225,N_15291);
xor U15402 (N_15402,N_15227,N_15299);
nand U15403 (N_15403,N_15221,N_15239);
nor U15404 (N_15404,N_15255,N_15269);
and U15405 (N_15405,N_15293,N_15363);
nor U15406 (N_15406,N_15367,N_15378);
or U15407 (N_15407,N_15246,N_15341);
nand U15408 (N_15408,N_15265,N_15354);
nor U15409 (N_15409,N_15216,N_15310);
nor U15410 (N_15410,N_15257,N_15296);
and U15411 (N_15411,N_15348,N_15351);
nand U15412 (N_15412,N_15364,N_15284);
nor U15413 (N_15413,N_15346,N_15350);
and U15414 (N_15414,N_15277,N_15306);
nor U15415 (N_15415,N_15386,N_15353);
and U15416 (N_15416,N_15251,N_15218);
or U15417 (N_15417,N_15315,N_15394);
or U15418 (N_15418,N_15336,N_15314);
and U15419 (N_15419,N_15254,N_15243);
or U15420 (N_15420,N_15339,N_15248);
or U15421 (N_15421,N_15381,N_15222);
nor U15422 (N_15422,N_15259,N_15202);
nand U15423 (N_15423,N_15332,N_15223);
xor U15424 (N_15424,N_15272,N_15256);
nor U15425 (N_15425,N_15266,N_15334);
and U15426 (N_15426,N_15396,N_15304);
nor U15427 (N_15427,N_15333,N_15313);
and U15428 (N_15428,N_15281,N_15365);
xor U15429 (N_15429,N_15379,N_15327);
nand U15430 (N_15430,N_15276,N_15324);
or U15431 (N_15431,N_15374,N_15268);
and U15432 (N_15432,N_15279,N_15377);
nand U15433 (N_15433,N_15358,N_15236);
and U15434 (N_15434,N_15282,N_15275);
nor U15435 (N_15435,N_15229,N_15270);
and U15436 (N_15436,N_15340,N_15330);
or U15437 (N_15437,N_15298,N_15263);
nand U15438 (N_15438,N_15344,N_15212);
and U15439 (N_15439,N_15321,N_15375);
or U15440 (N_15440,N_15214,N_15205);
xor U15441 (N_15441,N_15385,N_15283);
nand U15442 (N_15442,N_15397,N_15390);
nand U15443 (N_15443,N_15368,N_15372);
nand U15444 (N_15444,N_15206,N_15247);
nor U15445 (N_15445,N_15305,N_15217);
and U15446 (N_15446,N_15231,N_15398);
xnor U15447 (N_15447,N_15343,N_15326);
or U15448 (N_15448,N_15307,N_15235);
and U15449 (N_15449,N_15280,N_15319);
xnor U15450 (N_15450,N_15253,N_15380);
or U15451 (N_15451,N_15383,N_15328);
xnor U15452 (N_15452,N_15242,N_15320);
and U15453 (N_15453,N_15311,N_15317);
xnor U15454 (N_15454,N_15342,N_15384);
nand U15455 (N_15455,N_15271,N_15287);
nand U15456 (N_15456,N_15244,N_15369);
xor U15457 (N_15457,N_15207,N_15261);
and U15458 (N_15458,N_15387,N_15215);
xor U15459 (N_15459,N_15349,N_15219);
nand U15460 (N_15460,N_15258,N_15308);
or U15461 (N_15461,N_15382,N_15295);
nor U15462 (N_15462,N_15399,N_15201);
xnor U15463 (N_15463,N_15392,N_15371);
nand U15464 (N_15464,N_15335,N_15210);
nor U15465 (N_15465,N_15357,N_15240);
nor U15466 (N_15466,N_15347,N_15355);
xor U15467 (N_15467,N_15331,N_15370);
nor U15468 (N_15468,N_15388,N_15323);
and U15469 (N_15469,N_15318,N_15262);
nand U15470 (N_15470,N_15252,N_15273);
and U15471 (N_15471,N_15264,N_15389);
nor U15472 (N_15472,N_15267,N_15285);
nor U15473 (N_15473,N_15274,N_15294);
nand U15474 (N_15474,N_15312,N_15373);
or U15475 (N_15475,N_15292,N_15316);
and U15476 (N_15476,N_15220,N_15376);
nand U15477 (N_15477,N_15224,N_15391);
and U15478 (N_15478,N_15359,N_15232);
xor U15479 (N_15479,N_15322,N_15200);
or U15480 (N_15480,N_15356,N_15338);
or U15481 (N_15481,N_15288,N_15226);
and U15482 (N_15482,N_15337,N_15228);
and U15483 (N_15483,N_15237,N_15245);
nor U15484 (N_15484,N_15289,N_15249);
nand U15485 (N_15485,N_15241,N_15362);
xor U15486 (N_15486,N_15352,N_15290);
nor U15487 (N_15487,N_15230,N_15301);
xnor U15488 (N_15488,N_15203,N_15204);
or U15489 (N_15489,N_15366,N_15233);
and U15490 (N_15490,N_15234,N_15300);
or U15491 (N_15491,N_15303,N_15395);
nand U15492 (N_15492,N_15250,N_15345);
or U15493 (N_15493,N_15325,N_15329);
nor U15494 (N_15494,N_15278,N_15238);
and U15495 (N_15495,N_15208,N_15286);
or U15496 (N_15496,N_15309,N_15260);
and U15497 (N_15497,N_15393,N_15213);
nand U15498 (N_15498,N_15209,N_15297);
nand U15499 (N_15499,N_15302,N_15361);
or U15500 (N_15500,N_15327,N_15265);
or U15501 (N_15501,N_15392,N_15257);
and U15502 (N_15502,N_15256,N_15292);
or U15503 (N_15503,N_15368,N_15362);
xor U15504 (N_15504,N_15259,N_15360);
nor U15505 (N_15505,N_15366,N_15213);
or U15506 (N_15506,N_15216,N_15265);
xor U15507 (N_15507,N_15380,N_15333);
xnor U15508 (N_15508,N_15307,N_15211);
xor U15509 (N_15509,N_15284,N_15295);
nand U15510 (N_15510,N_15210,N_15319);
xor U15511 (N_15511,N_15268,N_15214);
or U15512 (N_15512,N_15274,N_15283);
or U15513 (N_15513,N_15275,N_15319);
xnor U15514 (N_15514,N_15202,N_15326);
xnor U15515 (N_15515,N_15321,N_15254);
nand U15516 (N_15516,N_15381,N_15261);
xnor U15517 (N_15517,N_15228,N_15393);
nand U15518 (N_15518,N_15234,N_15301);
nand U15519 (N_15519,N_15296,N_15333);
nor U15520 (N_15520,N_15222,N_15357);
and U15521 (N_15521,N_15276,N_15367);
nand U15522 (N_15522,N_15290,N_15368);
nor U15523 (N_15523,N_15266,N_15331);
nor U15524 (N_15524,N_15267,N_15369);
and U15525 (N_15525,N_15315,N_15314);
nand U15526 (N_15526,N_15236,N_15375);
or U15527 (N_15527,N_15282,N_15265);
nand U15528 (N_15528,N_15303,N_15331);
nand U15529 (N_15529,N_15323,N_15212);
nor U15530 (N_15530,N_15278,N_15219);
nand U15531 (N_15531,N_15393,N_15382);
nand U15532 (N_15532,N_15247,N_15245);
or U15533 (N_15533,N_15306,N_15372);
nor U15534 (N_15534,N_15270,N_15385);
or U15535 (N_15535,N_15232,N_15368);
xor U15536 (N_15536,N_15237,N_15243);
and U15537 (N_15537,N_15230,N_15276);
and U15538 (N_15538,N_15259,N_15204);
nand U15539 (N_15539,N_15269,N_15214);
xor U15540 (N_15540,N_15348,N_15361);
nor U15541 (N_15541,N_15241,N_15265);
xor U15542 (N_15542,N_15239,N_15215);
and U15543 (N_15543,N_15307,N_15368);
xor U15544 (N_15544,N_15341,N_15344);
nor U15545 (N_15545,N_15373,N_15211);
nor U15546 (N_15546,N_15308,N_15267);
and U15547 (N_15547,N_15216,N_15239);
nand U15548 (N_15548,N_15284,N_15346);
and U15549 (N_15549,N_15361,N_15207);
nand U15550 (N_15550,N_15310,N_15321);
and U15551 (N_15551,N_15352,N_15284);
and U15552 (N_15552,N_15293,N_15228);
or U15553 (N_15553,N_15304,N_15328);
nor U15554 (N_15554,N_15296,N_15208);
and U15555 (N_15555,N_15291,N_15200);
and U15556 (N_15556,N_15269,N_15343);
nor U15557 (N_15557,N_15218,N_15256);
or U15558 (N_15558,N_15233,N_15224);
or U15559 (N_15559,N_15264,N_15379);
and U15560 (N_15560,N_15361,N_15290);
nor U15561 (N_15561,N_15274,N_15394);
nand U15562 (N_15562,N_15353,N_15349);
or U15563 (N_15563,N_15361,N_15389);
nor U15564 (N_15564,N_15331,N_15304);
and U15565 (N_15565,N_15358,N_15272);
nor U15566 (N_15566,N_15343,N_15351);
nand U15567 (N_15567,N_15353,N_15339);
nor U15568 (N_15568,N_15339,N_15287);
nand U15569 (N_15569,N_15281,N_15266);
and U15570 (N_15570,N_15202,N_15374);
nand U15571 (N_15571,N_15229,N_15346);
xor U15572 (N_15572,N_15367,N_15317);
or U15573 (N_15573,N_15394,N_15293);
or U15574 (N_15574,N_15291,N_15389);
and U15575 (N_15575,N_15369,N_15347);
or U15576 (N_15576,N_15336,N_15266);
or U15577 (N_15577,N_15207,N_15239);
nand U15578 (N_15578,N_15324,N_15257);
and U15579 (N_15579,N_15347,N_15338);
xnor U15580 (N_15580,N_15285,N_15386);
nor U15581 (N_15581,N_15392,N_15208);
nand U15582 (N_15582,N_15282,N_15383);
and U15583 (N_15583,N_15360,N_15352);
and U15584 (N_15584,N_15307,N_15234);
nand U15585 (N_15585,N_15312,N_15345);
nor U15586 (N_15586,N_15240,N_15232);
nand U15587 (N_15587,N_15235,N_15352);
or U15588 (N_15588,N_15258,N_15333);
nor U15589 (N_15589,N_15315,N_15329);
xor U15590 (N_15590,N_15387,N_15279);
xor U15591 (N_15591,N_15339,N_15270);
nor U15592 (N_15592,N_15388,N_15390);
or U15593 (N_15593,N_15290,N_15327);
nand U15594 (N_15594,N_15332,N_15399);
nor U15595 (N_15595,N_15266,N_15298);
or U15596 (N_15596,N_15205,N_15374);
or U15597 (N_15597,N_15336,N_15396);
xnor U15598 (N_15598,N_15392,N_15220);
and U15599 (N_15599,N_15357,N_15259);
or U15600 (N_15600,N_15536,N_15462);
or U15601 (N_15601,N_15418,N_15436);
nor U15602 (N_15602,N_15444,N_15556);
nor U15603 (N_15603,N_15598,N_15498);
and U15604 (N_15604,N_15403,N_15544);
xnor U15605 (N_15605,N_15596,N_15489);
or U15606 (N_15606,N_15542,N_15594);
or U15607 (N_15607,N_15560,N_15409);
or U15608 (N_15608,N_15460,N_15518);
nor U15609 (N_15609,N_15591,N_15589);
xnor U15610 (N_15610,N_15561,N_15491);
xor U15611 (N_15611,N_15547,N_15475);
and U15612 (N_15612,N_15463,N_15527);
xnor U15613 (N_15613,N_15434,N_15582);
xnor U15614 (N_15614,N_15538,N_15555);
nand U15615 (N_15615,N_15511,N_15412);
or U15616 (N_15616,N_15474,N_15421);
nor U15617 (N_15617,N_15587,N_15401);
or U15618 (N_15618,N_15593,N_15530);
xnor U15619 (N_15619,N_15445,N_15437);
nand U15620 (N_15620,N_15514,N_15459);
or U15621 (N_15621,N_15422,N_15519);
and U15622 (N_15622,N_15599,N_15590);
nor U15623 (N_15623,N_15515,N_15573);
xor U15624 (N_15624,N_15488,N_15465);
nand U15625 (N_15625,N_15579,N_15427);
or U15626 (N_15626,N_15513,N_15402);
nor U15627 (N_15627,N_15477,N_15446);
xnor U15628 (N_15628,N_15450,N_15563);
nand U15629 (N_15629,N_15578,N_15440);
and U15630 (N_15630,N_15490,N_15423);
xor U15631 (N_15631,N_15505,N_15535);
xnor U15632 (N_15632,N_15497,N_15478);
and U15633 (N_15633,N_15433,N_15453);
xnor U15634 (N_15634,N_15520,N_15583);
and U15635 (N_15635,N_15439,N_15580);
xnor U15636 (N_15636,N_15565,N_15558);
or U15637 (N_15637,N_15476,N_15549);
and U15638 (N_15638,N_15562,N_15410);
and U15639 (N_15639,N_15567,N_15471);
xnor U15640 (N_15640,N_15571,N_15577);
nand U15641 (N_15641,N_15419,N_15479);
xor U15642 (N_15642,N_15552,N_15415);
nor U15643 (N_15643,N_15493,N_15575);
or U15644 (N_15644,N_15508,N_15526);
xor U15645 (N_15645,N_15458,N_15597);
and U15646 (N_15646,N_15443,N_15408);
or U15647 (N_15647,N_15554,N_15503);
and U15648 (N_15648,N_15470,N_15537);
xor U15649 (N_15649,N_15539,N_15523);
nand U15650 (N_15650,N_15425,N_15411);
xnor U15651 (N_15651,N_15550,N_15559);
xor U15652 (N_15652,N_15532,N_15522);
nor U15653 (N_15653,N_15502,N_15473);
nand U15654 (N_15654,N_15517,N_15533);
and U15655 (N_15655,N_15551,N_15595);
and U15656 (N_15656,N_15507,N_15495);
nand U15657 (N_15657,N_15510,N_15414);
and U15658 (N_15658,N_15413,N_15420);
xnor U15659 (N_15659,N_15428,N_15442);
xnor U15660 (N_15660,N_15405,N_15480);
xnor U15661 (N_15661,N_15592,N_15521);
or U15662 (N_15662,N_15456,N_15528);
or U15663 (N_15663,N_15529,N_15586);
nor U15664 (N_15664,N_15564,N_15534);
nor U15665 (N_15665,N_15492,N_15501);
nand U15666 (N_15666,N_15481,N_15404);
and U15667 (N_15667,N_15438,N_15452);
xor U15668 (N_15668,N_15531,N_15569);
and U15669 (N_15669,N_15540,N_15457);
nand U15670 (N_15670,N_15432,N_15572);
nor U15671 (N_15671,N_15429,N_15499);
nor U15672 (N_15672,N_15487,N_15543);
xnor U15673 (N_15673,N_15417,N_15461);
nand U15674 (N_15674,N_15504,N_15426);
or U15675 (N_15675,N_15576,N_15400);
nor U15676 (N_15676,N_15566,N_15449);
nor U15677 (N_15677,N_15451,N_15570);
xnor U15678 (N_15678,N_15574,N_15455);
nand U15679 (N_15679,N_15509,N_15406);
or U15680 (N_15680,N_15512,N_15525);
nor U15681 (N_15681,N_15584,N_15545);
or U15682 (N_15682,N_15541,N_15467);
nor U15683 (N_15683,N_15407,N_15466);
or U15684 (N_15684,N_15485,N_15430);
nand U15685 (N_15685,N_15516,N_15416);
nand U15686 (N_15686,N_15486,N_15506);
nand U15687 (N_15687,N_15585,N_15431);
nand U15688 (N_15688,N_15482,N_15424);
nor U15689 (N_15689,N_15472,N_15557);
nand U15690 (N_15690,N_15448,N_15581);
and U15691 (N_15691,N_15546,N_15524);
nand U15692 (N_15692,N_15484,N_15468);
xor U15693 (N_15693,N_15469,N_15483);
nand U15694 (N_15694,N_15435,N_15588);
nor U15695 (N_15695,N_15454,N_15464);
and U15696 (N_15696,N_15568,N_15496);
or U15697 (N_15697,N_15441,N_15553);
or U15698 (N_15698,N_15500,N_15494);
nand U15699 (N_15699,N_15447,N_15548);
or U15700 (N_15700,N_15522,N_15517);
nand U15701 (N_15701,N_15534,N_15561);
or U15702 (N_15702,N_15571,N_15497);
xor U15703 (N_15703,N_15517,N_15492);
xnor U15704 (N_15704,N_15599,N_15596);
nand U15705 (N_15705,N_15531,N_15586);
xnor U15706 (N_15706,N_15596,N_15460);
xnor U15707 (N_15707,N_15413,N_15408);
nor U15708 (N_15708,N_15570,N_15550);
and U15709 (N_15709,N_15569,N_15453);
xnor U15710 (N_15710,N_15523,N_15439);
or U15711 (N_15711,N_15460,N_15548);
nand U15712 (N_15712,N_15494,N_15513);
nor U15713 (N_15713,N_15550,N_15546);
and U15714 (N_15714,N_15412,N_15456);
nand U15715 (N_15715,N_15590,N_15531);
nand U15716 (N_15716,N_15491,N_15520);
or U15717 (N_15717,N_15501,N_15512);
and U15718 (N_15718,N_15517,N_15503);
nand U15719 (N_15719,N_15487,N_15493);
nor U15720 (N_15720,N_15464,N_15482);
or U15721 (N_15721,N_15418,N_15408);
and U15722 (N_15722,N_15414,N_15440);
xor U15723 (N_15723,N_15436,N_15433);
xor U15724 (N_15724,N_15413,N_15439);
xor U15725 (N_15725,N_15423,N_15463);
nor U15726 (N_15726,N_15505,N_15453);
xor U15727 (N_15727,N_15486,N_15511);
and U15728 (N_15728,N_15408,N_15415);
nand U15729 (N_15729,N_15567,N_15584);
and U15730 (N_15730,N_15560,N_15582);
nand U15731 (N_15731,N_15579,N_15495);
xor U15732 (N_15732,N_15410,N_15542);
xor U15733 (N_15733,N_15597,N_15498);
nand U15734 (N_15734,N_15483,N_15412);
or U15735 (N_15735,N_15506,N_15517);
nand U15736 (N_15736,N_15447,N_15481);
nor U15737 (N_15737,N_15414,N_15542);
and U15738 (N_15738,N_15522,N_15446);
nand U15739 (N_15739,N_15518,N_15488);
nand U15740 (N_15740,N_15585,N_15533);
nand U15741 (N_15741,N_15456,N_15557);
nor U15742 (N_15742,N_15447,N_15445);
and U15743 (N_15743,N_15536,N_15401);
and U15744 (N_15744,N_15446,N_15464);
and U15745 (N_15745,N_15584,N_15465);
nand U15746 (N_15746,N_15557,N_15420);
nor U15747 (N_15747,N_15511,N_15493);
nand U15748 (N_15748,N_15511,N_15452);
and U15749 (N_15749,N_15532,N_15485);
and U15750 (N_15750,N_15514,N_15434);
and U15751 (N_15751,N_15432,N_15418);
xnor U15752 (N_15752,N_15551,N_15498);
nor U15753 (N_15753,N_15581,N_15514);
nand U15754 (N_15754,N_15494,N_15462);
nor U15755 (N_15755,N_15568,N_15558);
and U15756 (N_15756,N_15482,N_15415);
nor U15757 (N_15757,N_15475,N_15407);
nand U15758 (N_15758,N_15577,N_15430);
nand U15759 (N_15759,N_15594,N_15586);
and U15760 (N_15760,N_15586,N_15423);
xnor U15761 (N_15761,N_15470,N_15589);
or U15762 (N_15762,N_15439,N_15500);
and U15763 (N_15763,N_15549,N_15414);
and U15764 (N_15764,N_15473,N_15577);
or U15765 (N_15765,N_15525,N_15538);
nand U15766 (N_15766,N_15526,N_15518);
nand U15767 (N_15767,N_15459,N_15531);
xnor U15768 (N_15768,N_15586,N_15472);
nor U15769 (N_15769,N_15510,N_15440);
nand U15770 (N_15770,N_15483,N_15486);
or U15771 (N_15771,N_15575,N_15475);
nor U15772 (N_15772,N_15404,N_15505);
nor U15773 (N_15773,N_15472,N_15530);
xnor U15774 (N_15774,N_15505,N_15599);
nor U15775 (N_15775,N_15404,N_15437);
xnor U15776 (N_15776,N_15529,N_15520);
or U15777 (N_15777,N_15417,N_15504);
xor U15778 (N_15778,N_15415,N_15457);
nor U15779 (N_15779,N_15541,N_15446);
nand U15780 (N_15780,N_15507,N_15577);
xor U15781 (N_15781,N_15508,N_15465);
and U15782 (N_15782,N_15569,N_15479);
nor U15783 (N_15783,N_15500,N_15592);
nand U15784 (N_15784,N_15565,N_15562);
and U15785 (N_15785,N_15487,N_15459);
nand U15786 (N_15786,N_15579,N_15589);
nor U15787 (N_15787,N_15404,N_15467);
or U15788 (N_15788,N_15495,N_15450);
or U15789 (N_15789,N_15508,N_15517);
xor U15790 (N_15790,N_15523,N_15519);
and U15791 (N_15791,N_15533,N_15430);
or U15792 (N_15792,N_15591,N_15487);
nor U15793 (N_15793,N_15511,N_15502);
or U15794 (N_15794,N_15573,N_15542);
xor U15795 (N_15795,N_15556,N_15438);
and U15796 (N_15796,N_15470,N_15500);
nor U15797 (N_15797,N_15406,N_15473);
and U15798 (N_15798,N_15431,N_15470);
nand U15799 (N_15799,N_15457,N_15402);
nand U15800 (N_15800,N_15600,N_15605);
xnor U15801 (N_15801,N_15711,N_15622);
or U15802 (N_15802,N_15736,N_15710);
or U15803 (N_15803,N_15760,N_15649);
or U15804 (N_15804,N_15731,N_15657);
nor U15805 (N_15805,N_15708,N_15721);
nor U15806 (N_15806,N_15735,N_15677);
nand U15807 (N_15807,N_15637,N_15653);
xnor U15808 (N_15808,N_15730,N_15781);
and U15809 (N_15809,N_15686,N_15696);
nor U15810 (N_15810,N_15739,N_15672);
nand U15811 (N_15811,N_15723,N_15635);
nand U15812 (N_15812,N_15674,N_15770);
or U15813 (N_15813,N_15787,N_15669);
and U15814 (N_15814,N_15729,N_15722);
nand U15815 (N_15815,N_15684,N_15749);
nor U15816 (N_15816,N_15790,N_15639);
and U15817 (N_15817,N_15705,N_15642);
and U15818 (N_15818,N_15706,N_15695);
nor U15819 (N_15819,N_15606,N_15691);
nor U15820 (N_15820,N_15659,N_15614);
nor U15821 (N_15821,N_15631,N_15772);
or U15822 (N_15822,N_15699,N_15636);
xor U15823 (N_15823,N_15746,N_15685);
nor U15824 (N_15824,N_15757,N_15724);
nand U15825 (N_15825,N_15681,N_15655);
nor U15826 (N_15826,N_15633,N_15626);
nor U15827 (N_15827,N_15741,N_15785);
and U15828 (N_15828,N_15767,N_15717);
and U15829 (N_15829,N_15630,N_15713);
xor U15830 (N_15830,N_15640,N_15766);
or U15831 (N_15831,N_15628,N_15701);
nor U15832 (N_15832,N_15698,N_15732);
and U15833 (N_15833,N_15678,N_15758);
nor U15834 (N_15834,N_15765,N_15603);
and U15835 (N_15835,N_15769,N_15641);
nor U15836 (N_15836,N_15777,N_15668);
and U15837 (N_15837,N_15661,N_15750);
or U15838 (N_15838,N_15703,N_15646);
nor U15839 (N_15839,N_15658,N_15793);
nor U15840 (N_15840,N_15602,N_15704);
nor U15841 (N_15841,N_15795,N_15715);
or U15842 (N_15842,N_15733,N_15670);
and U15843 (N_15843,N_15617,N_15762);
and U15844 (N_15844,N_15656,N_15634);
or U15845 (N_15845,N_15747,N_15745);
or U15846 (N_15846,N_15783,N_15612);
nor U15847 (N_15847,N_15780,N_15676);
xnor U15848 (N_15848,N_15654,N_15725);
nand U15849 (N_15849,N_15697,N_15738);
or U15850 (N_15850,N_15751,N_15682);
nand U15851 (N_15851,N_15671,N_15687);
nor U15852 (N_15852,N_15629,N_15776);
or U15853 (N_15853,N_15719,N_15615);
xnor U15854 (N_15854,N_15768,N_15752);
xnor U15855 (N_15855,N_15726,N_15618);
or U15856 (N_15856,N_15782,N_15619);
nand U15857 (N_15857,N_15779,N_15673);
or U15858 (N_15858,N_15644,N_15647);
xor U15859 (N_15859,N_15643,N_15693);
or U15860 (N_15860,N_15601,N_15609);
nor U15861 (N_15861,N_15675,N_15796);
xnor U15862 (N_15862,N_15788,N_15786);
nor U15863 (N_15863,N_15611,N_15728);
nor U15864 (N_15864,N_15727,N_15616);
nand U15865 (N_15865,N_15666,N_15620);
nor U15866 (N_15866,N_15761,N_15667);
or U15867 (N_15867,N_15755,N_15700);
or U15868 (N_15868,N_15664,N_15638);
and U15869 (N_15869,N_15789,N_15742);
and U15870 (N_15870,N_15688,N_15756);
nor U15871 (N_15871,N_15709,N_15692);
nand U15872 (N_15872,N_15798,N_15625);
xnor U15873 (N_15873,N_15716,N_15702);
and U15874 (N_15874,N_15740,N_15771);
nand U15875 (N_15875,N_15748,N_15712);
xnor U15876 (N_15876,N_15683,N_15707);
nand U15877 (N_15877,N_15799,N_15623);
nor U15878 (N_15878,N_15794,N_15784);
and U15879 (N_15879,N_15763,N_15651);
nand U15880 (N_15880,N_15662,N_15791);
xor U15881 (N_15881,N_15753,N_15680);
and U15882 (N_15882,N_15652,N_15775);
nand U15883 (N_15883,N_15660,N_15663);
nand U15884 (N_15884,N_15754,N_15774);
or U15885 (N_15885,N_15624,N_15632);
and U15886 (N_15886,N_15743,N_15650);
xnor U15887 (N_15887,N_15714,N_15613);
nor U15888 (N_15888,N_15621,N_15665);
xnor U15889 (N_15889,N_15734,N_15645);
and U15890 (N_15890,N_15720,N_15773);
or U15891 (N_15891,N_15604,N_15694);
nand U15892 (N_15892,N_15718,N_15737);
nor U15893 (N_15893,N_15689,N_15679);
or U15894 (N_15894,N_15759,N_15797);
or U15895 (N_15895,N_15610,N_15690);
or U15896 (N_15896,N_15764,N_15778);
and U15897 (N_15897,N_15744,N_15627);
and U15898 (N_15898,N_15648,N_15792);
and U15899 (N_15899,N_15608,N_15607);
nand U15900 (N_15900,N_15672,N_15772);
xnor U15901 (N_15901,N_15784,N_15658);
and U15902 (N_15902,N_15760,N_15752);
xnor U15903 (N_15903,N_15703,N_15632);
nor U15904 (N_15904,N_15621,N_15687);
nor U15905 (N_15905,N_15644,N_15737);
nand U15906 (N_15906,N_15690,N_15689);
nand U15907 (N_15907,N_15742,N_15786);
or U15908 (N_15908,N_15731,N_15699);
nor U15909 (N_15909,N_15691,N_15793);
xnor U15910 (N_15910,N_15601,N_15641);
nor U15911 (N_15911,N_15635,N_15797);
xnor U15912 (N_15912,N_15754,N_15669);
nand U15913 (N_15913,N_15723,N_15704);
xnor U15914 (N_15914,N_15713,N_15737);
and U15915 (N_15915,N_15699,N_15727);
and U15916 (N_15916,N_15613,N_15635);
or U15917 (N_15917,N_15602,N_15740);
nor U15918 (N_15918,N_15762,N_15681);
xnor U15919 (N_15919,N_15794,N_15654);
nand U15920 (N_15920,N_15641,N_15667);
nand U15921 (N_15921,N_15727,N_15637);
or U15922 (N_15922,N_15770,N_15769);
nand U15923 (N_15923,N_15728,N_15633);
or U15924 (N_15924,N_15757,N_15702);
nor U15925 (N_15925,N_15651,N_15738);
and U15926 (N_15926,N_15749,N_15704);
or U15927 (N_15927,N_15797,N_15640);
nor U15928 (N_15928,N_15773,N_15695);
or U15929 (N_15929,N_15740,N_15759);
or U15930 (N_15930,N_15682,N_15782);
and U15931 (N_15931,N_15668,N_15758);
and U15932 (N_15932,N_15792,N_15639);
nor U15933 (N_15933,N_15760,N_15786);
xnor U15934 (N_15934,N_15604,N_15625);
nand U15935 (N_15935,N_15674,N_15754);
nand U15936 (N_15936,N_15738,N_15670);
or U15937 (N_15937,N_15622,N_15675);
nand U15938 (N_15938,N_15723,N_15779);
and U15939 (N_15939,N_15755,N_15716);
or U15940 (N_15940,N_15660,N_15694);
xnor U15941 (N_15941,N_15733,N_15616);
and U15942 (N_15942,N_15762,N_15746);
and U15943 (N_15943,N_15772,N_15755);
and U15944 (N_15944,N_15766,N_15716);
nor U15945 (N_15945,N_15743,N_15689);
nor U15946 (N_15946,N_15694,N_15671);
nand U15947 (N_15947,N_15612,N_15604);
xor U15948 (N_15948,N_15600,N_15748);
xnor U15949 (N_15949,N_15698,N_15795);
or U15950 (N_15950,N_15752,N_15736);
and U15951 (N_15951,N_15606,N_15669);
nand U15952 (N_15952,N_15746,N_15710);
or U15953 (N_15953,N_15624,N_15731);
xnor U15954 (N_15954,N_15727,N_15681);
or U15955 (N_15955,N_15764,N_15687);
xnor U15956 (N_15956,N_15651,N_15707);
or U15957 (N_15957,N_15778,N_15707);
nand U15958 (N_15958,N_15661,N_15782);
nand U15959 (N_15959,N_15705,N_15717);
xor U15960 (N_15960,N_15622,N_15798);
nand U15961 (N_15961,N_15703,N_15778);
xor U15962 (N_15962,N_15638,N_15789);
and U15963 (N_15963,N_15678,N_15663);
nor U15964 (N_15964,N_15788,N_15694);
or U15965 (N_15965,N_15649,N_15717);
or U15966 (N_15966,N_15692,N_15708);
or U15967 (N_15967,N_15728,N_15675);
xor U15968 (N_15968,N_15777,N_15795);
nand U15969 (N_15969,N_15762,N_15726);
xor U15970 (N_15970,N_15717,N_15768);
xnor U15971 (N_15971,N_15707,N_15769);
or U15972 (N_15972,N_15790,N_15779);
nor U15973 (N_15973,N_15718,N_15662);
nor U15974 (N_15974,N_15772,N_15680);
xor U15975 (N_15975,N_15639,N_15653);
or U15976 (N_15976,N_15611,N_15627);
xnor U15977 (N_15977,N_15675,N_15766);
xor U15978 (N_15978,N_15677,N_15682);
or U15979 (N_15979,N_15702,N_15763);
and U15980 (N_15980,N_15786,N_15796);
and U15981 (N_15981,N_15654,N_15768);
nand U15982 (N_15982,N_15778,N_15646);
xor U15983 (N_15983,N_15798,N_15720);
xor U15984 (N_15984,N_15724,N_15778);
or U15985 (N_15985,N_15634,N_15767);
nand U15986 (N_15986,N_15682,N_15643);
nor U15987 (N_15987,N_15799,N_15696);
xnor U15988 (N_15988,N_15607,N_15753);
xnor U15989 (N_15989,N_15602,N_15765);
nand U15990 (N_15990,N_15690,N_15749);
nand U15991 (N_15991,N_15645,N_15658);
xnor U15992 (N_15992,N_15600,N_15633);
or U15993 (N_15993,N_15734,N_15798);
and U15994 (N_15994,N_15736,N_15682);
xor U15995 (N_15995,N_15749,N_15632);
xnor U15996 (N_15996,N_15651,N_15760);
xnor U15997 (N_15997,N_15711,N_15745);
xor U15998 (N_15998,N_15724,N_15657);
nand U15999 (N_15999,N_15697,N_15668);
and U16000 (N_16000,N_15828,N_15894);
and U16001 (N_16001,N_15815,N_15857);
or U16002 (N_16002,N_15935,N_15985);
nor U16003 (N_16003,N_15836,N_15956);
nand U16004 (N_16004,N_15909,N_15991);
and U16005 (N_16005,N_15976,N_15879);
or U16006 (N_16006,N_15918,N_15937);
or U16007 (N_16007,N_15930,N_15814);
and U16008 (N_16008,N_15870,N_15950);
nor U16009 (N_16009,N_15901,N_15801);
nor U16010 (N_16010,N_15912,N_15876);
and U16011 (N_16011,N_15844,N_15917);
xnor U16012 (N_16012,N_15943,N_15819);
and U16013 (N_16013,N_15959,N_15978);
and U16014 (N_16014,N_15858,N_15885);
and U16015 (N_16015,N_15804,N_15942);
nand U16016 (N_16016,N_15924,N_15896);
and U16017 (N_16017,N_15877,N_15954);
nor U16018 (N_16018,N_15975,N_15986);
or U16019 (N_16019,N_15981,N_15899);
xor U16020 (N_16020,N_15977,N_15931);
nor U16021 (N_16021,N_15852,N_15854);
nor U16022 (N_16022,N_15862,N_15875);
or U16023 (N_16023,N_15968,N_15808);
or U16024 (N_16024,N_15970,N_15921);
or U16025 (N_16025,N_15940,N_15897);
and U16026 (N_16026,N_15973,N_15802);
nor U16027 (N_16027,N_15847,N_15972);
and U16028 (N_16028,N_15997,N_15998);
nand U16029 (N_16029,N_15961,N_15807);
and U16030 (N_16030,N_15927,N_15872);
nor U16031 (N_16031,N_15829,N_15925);
or U16032 (N_16032,N_15929,N_15895);
or U16033 (N_16033,N_15869,N_15955);
or U16034 (N_16034,N_15818,N_15945);
xnor U16035 (N_16035,N_15920,N_15884);
and U16036 (N_16036,N_15850,N_15839);
xor U16037 (N_16037,N_15987,N_15800);
xnor U16038 (N_16038,N_15989,N_15845);
xnor U16039 (N_16039,N_15810,N_15892);
or U16040 (N_16040,N_15873,N_15840);
nor U16041 (N_16041,N_15880,N_15837);
and U16042 (N_16042,N_15910,N_15886);
or U16043 (N_16043,N_15992,N_15883);
xnor U16044 (N_16044,N_15851,N_15971);
nor U16045 (N_16045,N_15824,N_15865);
nor U16046 (N_16046,N_15887,N_15835);
xnor U16047 (N_16047,N_15821,N_15965);
and U16048 (N_16048,N_15932,N_15962);
nor U16049 (N_16049,N_15980,N_15947);
and U16050 (N_16050,N_15830,N_15881);
or U16051 (N_16051,N_15904,N_15860);
nand U16052 (N_16052,N_15826,N_15934);
and U16053 (N_16053,N_15933,N_15966);
or U16054 (N_16054,N_15906,N_15898);
nand U16055 (N_16055,N_15939,N_15949);
nor U16056 (N_16056,N_15900,N_15936);
xnor U16057 (N_16057,N_15984,N_15964);
nor U16058 (N_16058,N_15866,N_15834);
nand U16059 (N_16059,N_15915,N_15832);
nand U16060 (N_16060,N_15893,N_15805);
nand U16061 (N_16061,N_15831,N_15817);
nand U16062 (N_16062,N_15864,N_15946);
or U16063 (N_16063,N_15994,N_15841);
nand U16064 (N_16064,N_15843,N_15948);
and U16065 (N_16065,N_15952,N_15913);
and U16066 (N_16066,N_15902,N_15833);
or U16067 (N_16067,N_15996,N_15960);
nor U16068 (N_16068,N_15905,N_15811);
nand U16069 (N_16069,N_15867,N_15983);
and U16070 (N_16070,N_15907,N_15812);
xnor U16071 (N_16071,N_15903,N_15982);
nor U16072 (N_16072,N_15914,N_15846);
and U16073 (N_16073,N_15820,N_15974);
and U16074 (N_16074,N_15813,N_15838);
nand U16075 (N_16075,N_15859,N_15938);
nor U16076 (N_16076,N_15855,N_15889);
nand U16077 (N_16077,N_15891,N_15923);
and U16078 (N_16078,N_15908,N_15988);
or U16079 (N_16079,N_15919,N_15827);
nand U16080 (N_16080,N_15848,N_15941);
or U16081 (N_16081,N_15922,N_15911);
or U16082 (N_16082,N_15944,N_15963);
nand U16083 (N_16083,N_15957,N_15842);
and U16084 (N_16084,N_15878,N_15823);
xor U16085 (N_16085,N_15809,N_15993);
nor U16086 (N_16086,N_15882,N_15999);
xnor U16087 (N_16087,N_15803,N_15958);
nand U16088 (N_16088,N_15806,N_15969);
nand U16089 (N_16089,N_15822,N_15916);
xnor U16090 (N_16090,N_15816,N_15928);
nand U16091 (N_16091,N_15953,N_15853);
nor U16092 (N_16092,N_15967,N_15861);
or U16093 (N_16093,N_15995,N_15951);
xor U16094 (N_16094,N_15926,N_15888);
nor U16095 (N_16095,N_15849,N_15874);
and U16096 (N_16096,N_15863,N_15979);
nor U16097 (N_16097,N_15990,N_15890);
nand U16098 (N_16098,N_15868,N_15825);
and U16099 (N_16099,N_15856,N_15871);
or U16100 (N_16100,N_15986,N_15963);
xnor U16101 (N_16101,N_15929,N_15905);
or U16102 (N_16102,N_15979,N_15865);
xor U16103 (N_16103,N_15816,N_15955);
or U16104 (N_16104,N_15975,N_15869);
nor U16105 (N_16105,N_15979,N_15819);
nor U16106 (N_16106,N_15822,N_15888);
and U16107 (N_16107,N_15828,N_15809);
xor U16108 (N_16108,N_15964,N_15804);
or U16109 (N_16109,N_15869,N_15935);
and U16110 (N_16110,N_15872,N_15933);
nor U16111 (N_16111,N_15819,N_15882);
nand U16112 (N_16112,N_15868,N_15802);
xnor U16113 (N_16113,N_15887,N_15813);
nand U16114 (N_16114,N_15924,N_15811);
nor U16115 (N_16115,N_15923,N_15918);
and U16116 (N_16116,N_15852,N_15973);
or U16117 (N_16117,N_15926,N_15860);
and U16118 (N_16118,N_15927,N_15822);
nand U16119 (N_16119,N_15862,N_15840);
nor U16120 (N_16120,N_15880,N_15819);
nor U16121 (N_16121,N_15967,N_15908);
or U16122 (N_16122,N_15908,N_15994);
xnor U16123 (N_16123,N_15981,N_15881);
nand U16124 (N_16124,N_15844,N_15921);
nand U16125 (N_16125,N_15964,N_15992);
or U16126 (N_16126,N_15932,N_15809);
nor U16127 (N_16127,N_15871,N_15972);
xnor U16128 (N_16128,N_15881,N_15999);
nand U16129 (N_16129,N_15894,N_15857);
or U16130 (N_16130,N_15874,N_15881);
nor U16131 (N_16131,N_15840,N_15883);
xnor U16132 (N_16132,N_15877,N_15914);
nor U16133 (N_16133,N_15872,N_15838);
and U16134 (N_16134,N_15977,N_15915);
xor U16135 (N_16135,N_15828,N_15999);
nor U16136 (N_16136,N_15983,N_15878);
nor U16137 (N_16137,N_15821,N_15854);
or U16138 (N_16138,N_15936,N_15801);
nand U16139 (N_16139,N_15840,N_15893);
nor U16140 (N_16140,N_15903,N_15800);
xnor U16141 (N_16141,N_15863,N_15987);
or U16142 (N_16142,N_15862,N_15870);
nor U16143 (N_16143,N_15808,N_15846);
nand U16144 (N_16144,N_15829,N_15869);
xnor U16145 (N_16145,N_15893,N_15928);
nand U16146 (N_16146,N_15883,N_15956);
and U16147 (N_16147,N_15865,N_15859);
xor U16148 (N_16148,N_15906,N_15801);
or U16149 (N_16149,N_15889,N_15964);
or U16150 (N_16150,N_15851,N_15936);
or U16151 (N_16151,N_15888,N_15997);
nor U16152 (N_16152,N_15873,N_15813);
or U16153 (N_16153,N_15987,N_15940);
xor U16154 (N_16154,N_15841,N_15843);
and U16155 (N_16155,N_15996,N_15844);
and U16156 (N_16156,N_15833,N_15959);
or U16157 (N_16157,N_15890,N_15838);
and U16158 (N_16158,N_15970,N_15910);
or U16159 (N_16159,N_15936,N_15878);
nor U16160 (N_16160,N_15848,N_15870);
and U16161 (N_16161,N_15939,N_15857);
nor U16162 (N_16162,N_15923,N_15816);
and U16163 (N_16163,N_15826,N_15841);
xnor U16164 (N_16164,N_15819,N_15849);
nor U16165 (N_16165,N_15905,N_15956);
or U16166 (N_16166,N_15922,N_15923);
or U16167 (N_16167,N_15926,N_15820);
or U16168 (N_16168,N_15931,N_15868);
xor U16169 (N_16169,N_15802,N_15819);
and U16170 (N_16170,N_15809,N_15983);
xnor U16171 (N_16171,N_15828,N_15879);
nor U16172 (N_16172,N_15928,N_15892);
and U16173 (N_16173,N_15832,N_15903);
or U16174 (N_16174,N_15974,N_15960);
xor U16175 (N_16175,N_15982,N_15808);
or U16176 (N_16176,N_15811,N_15925);
or U16177 (N_16177,N_15929,N_15917);
xor U16178 (N_16178,N_15810,N_15883);
nand U16179 (N_16179,N_15831,N_15879);
nor U16180 (N_16180,N_15858,N_15835);
xnor U16181 (N_16181,N_15911,N_15915);
xor U16182 (N_16182,N_15828,N_15951);
nor U16183 (N_16183,N_15883,N_15965);
nor U16184 (N_16184,N_15950,N_15939);
nor U16185 (N_16185,N_15831,N_15979);
nand U16186 (N_16186,N_15842,N_15917);
or U16187 (N_16187,N_15907,N_15813);
nor U16188 (N_16188,N_15841,N_15802);
nor U16189 (N_16189,N_15972,N_15924);
nand U16190 (N_16190,N_15865,N_15990);
and U16191 (N_16191,N_15994,N_15826);
nand U16192 (N_16192,N_15917,N_15972);
nor U16193 (N_16193,N_15964,N_15820);
xor U16194 (N_16194,N_15929,N_15872);
and U16195 (N_16195,N_15939,N_15984);
and U16196 (N_16196,N_15829,N_15919);
xnor U16197 (N_16197,N_15816,N_15836);
nand U16198 (N_16198,N_15887,N_15811);
nor U16199 (N_16199,N_15904,N_15992);
or U16200 (N_16200,N_16173,N_16168);
or U16201 (N_16201,N_16015,N_16037);
xnor U16202 (N_16202,N_16097,N_16105);
nor U16203 (N_16203,N_16196,N_16134);
xnor U16204 (N_16204,N_16121,N_16058);
nand U16205 (N_16205,N_16065,N_16172);
nand U16206 (N_16206,N_16135,N_16125);
nand U16207 (N_16207,N_16059,N_16090);
or U16208 (N_16208,N_16195,N_16091);
and U16209 (N_16209,N_16095,N_16154);
or U16210 (N_16210,N_16141,N_16166);
or U16211 (N_16211,N_16063,N_16006);
or U16212 (N_16212,N_16061,N_16016);
nand U16213 (N_16213,N_16084,N_16187);
nor U16214 (N_16214,N_16115,N_16012);
and U16215 (N_16215,N_16126,N_16174);
nand U16216 (N_16216,N_16101,N_16169);
nor U16217 (N_16217,N_16096,N_16033);
and U16218 (N_16218,N_16040,N_16157);
xnor U16219 (N_16219,N_16041,N_16177);
nor U16220 (N_16220,N_16048,N_16190);
nor U16221 (N_16221,N_16165,N_16044);
nor U16222 (N_16222,N_16087,N_16122);
xor U16223 (N_16223,N_16132,N_16027);
nand U16224 (N_16224,N_16034,N_16054);
xnor U16225 (N_16225,N_16074,N_16197);
or U16226 (N_16226,N_16019,N_16124);
and U16227 (N_16227,N_16194,N_16029);
and U16228 (N_16228,N_16158,N_16103);
xor U16229 (N_16229,N_16171,N_16147);
nor U16230 (N_16230,N_16053,N_16070);
or U16231 (N_16231,N_16002,N_16080);
and U16232 (N_16232,N_16180,N_16017);
nand U16233 (N_16233,N_16039,N_16024);
nor U16234 (N_16234,N_16185,N_16081);
and U16235 (N_16235,N_16057,N_16131);
nand U16236 (N_16236,N_16191,N_16104);
nor U16237 (N_16237,N_16139,N_16077);
nand U16238 (N_16238,N_16127,N_16159);
nand U16239 (N_16239,N_16099,N_16082);
nor U16240 (N_16240,N_16123,N_16162);
and U16241 (N_16241,N_16178,N_16183);
xor U16242 (N_16242,N_16003,N_16170);
nand U16243 (N_16243,N_16140,N_16184);
nand U16244 (N_16244,N_16075,N_16021);
xnor U16245 (N_16245,N_16148,N_16193);
xor U16246 (N_16246,N_16026,N_16025);
xor U16247 (N_16247,N_16130,N_16102);
and U16248 (N_16248,N_16023,N_16085);
and U16249 (N_16249,N_16051,N_16013);
nor U16250 (N_16250,N_16004,N_16118);
nor U16251 (N_16251,N_16066,N_16011);
and U16252 (N_16252,N_16128,N_16000);
xor U16253 (N_16253,N_16056,N_16093);
nand U16254 (N_16254,N_16167,N_16129);
xnor U16255 (N_16255,N_16142,N_16146);
or U16256 (N_16256,N_16109,N_16144);
xor U16257 (N_16257,N_16164,N_16073);
nand U16258 (N_16258,N_16119,N_16107);
or U16259 (N_16259,N_16062,N_16050);
nor U16260 (N_16260,N_16067,N_16161);
nand U16261 (N_16261,N_16098,N_16116);
or U16262 (N_16262,N_16133,N_16136);
and U16263 (N_16263,N_16114,N_16078);
nor U16264 (N_16264,N_16181,N_16117);
or U16265 (N_16265,N_16176,N_16089);
xnor U16266 (N_16266,N_16001,N_16182);
and U16267 (N_16267,N_16031,N_16072);
or U16268 (N_16268,N_16138,N_16186);
xnor U16269 (N_16269,N_16088,N_16110);
nand U16270 (N_16270,N_16179,N_16064);
nor U16271 (N_16271,N_16156,N_16155);
and U16272 (N_16272,N_16137,N_16199);
or U16273 (N_16273,N_16149,N_16153);
or U16274 (N_16274,N_16175,N_16188);
xnor U16275 (N_16275,N_16032,N_16045);
xnor U16276 (N_16276,N_16092,N_16108);
or U16277 (N_16277,N_16068,N_16160);
nand U16278 (N_16278,N_16111,N_16192);
xnor U16279 (N_16279,N_16047,N_16055);
and U16280 (N_16280,N_16009,N_16152);
nor U16281 (N_16281,N_16106,N_16018);
nand U16282 (N_16282,N_16083,N_16010);
nand U16283 (N_16283,N_16049,N_16069);
nand U16284 (N_16284,N_16060,N_16113);
xnor U16285 (N_16285,N_16071,N_16007);
or U16286 (N_16286,N_16151,N_16100);
nand U16287 (N_16287,N_16038,N_16042);
and U16288 (N_16288,N_16189,N_16030);
nor U16289 (N_16289,N_16112,N_16163);
and U16290 (N_16290,N_16036,N_16005);
nand U16291 (N_16291,N_16020,N_16120);
xnor U16292 (N_16292,N_16014,N_16076);
or U16293 (N_16293,N_16043,N_16079);
nor U16294 (N_16294,N_16052,N_16094);
or U16295 (N_16295,N_16086,N_16145);
xnor U16296 (N_16296,N_16022,N_16143);
nand U16297 (N_16297,N_16008,N_16046);
nand U16298 (N_16298,N_16150,N_16028);
or U16299 (N_16299,N_16035,N_16198);
nand U16300 (N_16300,N_16074,N_16135);
nor U16301 (N_16301,N_16164,N_16076);
or U16302 (N_16302,N_16047,N_16043);
nand U16303 (N_16303,N_16192,N_16083);
nand U16304 (N_16304,N_16082,N_16073);
or U16305 (N_16305,N_16129,N_16174);
or U16306 (N_16306,N_16106,N_16009);
nand U16307 (N_16307,N_16013,N_16085);
or U16308 (N_16308,N_16036,N_16188);
nor U16309 (N_16309,N_16020,N_16076);
nand U16310 (N_16310,N_16179,N_16126);
nor U16311 (N_16311,N_16193,N_16014);
nand U16312 (N_16312,N_16161,N_16182);
nand U16313 (N_16313,N_16031,N_16166);
xor U16314 (N_16314,N_16089,N_16132);
nand U16315 (N_16315,N_16094,N_16198);
nor U16316 (N_16316,N_16163,N_16078);
xnor U16317 (N_16317,N_16102,N_16116);
and U16318 (N_16318,N_16125,N_16188);
xor U16319 (N_16319,N_16135,N_16001);
and U16320 (N_16320,N_16030,N_16040);
xor U16321 (N_16321,N_16159,N_16192);
xnor U16322 (N_16322,N_16065,N_16174);
xor U16323 (N_16323,N_16099,N_16134);
xnor U16324 (N_16324,N_16050,N_16118);
nand U16325 (N_16325,N_16192,N_16107);
nand U16326 (N_16326,N_16033,N_16186);
nand U16327 (N_16327,N_16082,N_16153);
nor U16328 (N_16328,N_16064,N_16198);
nand U16329 (N_16329,N_16126,N_16051);
or U16330 (N_16330,N_16181,N_16185);
nand U16331 (N_16331,N_16069,N_16078);
xnor U16332 (N_16332,N_16035,N_16047);
nand U16333 (N_16333,N_16138,N_16182);
or U16334 (N_16334,N_16111,N_16167);
nor U16335 (N_16335,N_16096,N_16045);
nand U16336 (N_16336,N_16023,N_16028);
nand U16337 (N_16337,N_16044,N_16124);
nor U16338 (N_16338,N_16052,N_16060);
and U16339 (N_16339,N_16020,N_16191);
nor U16340 (N_16340,N_16113,N_16190);
or U16341 (N_16341,N_16110,N_16040);
nor U16342 (N_16342,N_16194,N_16152);
or U16343 (N_16343,N_16012,N_16016);
or U16344 (N_16344,N_16032,N_16099);
nor U16345 (N_16345,N_16179,N_16016);
and U16346 (N_16346,N_16075,N_16011);
or U16347 (N_16347,N_16075,N_16103);
and U16348 (N_16348,N_16098,N_16021);
nor U16349 (N_16349,N_16153,N_16041);
xnor U16350 (N_16350,N_16053,N_16061);
nor U16351 (N_16351,N_16127,N_16107);
and U16352 (N_16352,N_16057,N_16090);
xor U16353 (N_16353,N_16057,N_16029);
xor U16354 (N_16354,N_16095,N_16086);
xor U16355 (N_16355,N_16097,N_16011);
nand U16356 (N_16356,N_16188,N_16026);
nand U16357 (N_16357,N_16174,N_16106);
xor U16358 (N_16358,N_16134,N_16127);
and U16359 (N_16359,N_16158,N_16136);
nand U16360 (N_16360,N_16056,N_16181);
and U16361 (N_16361,N_16046,N_16053);
xor U16362 (N_16362,N_16195,N_16181);
and U16363 (N_16363,N_16074,N_16055);
xor U16364 (N_16364,N_16061,N_16070);
nand U16365 (N_16365,N_16081,N_16040);
and U16366 (N_16366,N_16119,N_16114);
and U16367 (N_16367,N_16135,N_16117);
xor U16368 (N_16368,N_16019,N_16155);
and U16369 (N_16369,N_16195,N_16191);
nor U16370 (N_16370,N_16063,N_16040);
and U16371 (N_16371,N_16132,N_16079);
or U16372 (N_16372,N_16155,N_16110);
and U16373 (N_16373,N_16043,N_16108);
nor U16374 (N_16374,N_16133,N_16171);
or U16375 (N_16375,N_16078,N_16038);
and U16376 (N_16376,N_16182,N_16193);
nand U16377 (N_16377,N_16048,N_16027);
nand U16378 (N_16378,N_16061,N_16067);
or U16379 (N_16379,N_16091,N_16071);
xnor U16380 (N_16380,N_16040,N_16098);
and U16381 (N_16381,N_16083,N_16072);
or U16382 (N_16382,N_16181,N_16199);
or U16383 (N_16383,N_16154,N_16188);
or U16384 (N_16384,N_16198,N_16133);
nor U16385 (N_16385,N_16050,N_16110);
or U16386 (N_16386,N_16062,N_16192);
xnor U16387 (N_16387,N_16183,N_16102);
and U16388 (N_16388,N_16168,N_16000);
and U16389 (N_16389,N_16127,N_16045);
or U16390 (N_16390,N_16018,N_16083);
nor U16391 (N_16391,N_16053,N_16097);
nand U16392 (N_16392,N_16072,N_16131);
xnor U16393 (N_16393,N_16084,N_16164);
and U16394 (N_16394,N_16107,N_16051);
and U16395 (N_16395,N_16025,N_16198);
nor U16396 (N_16396,N_16169,N_16009);
xnor U16397 (N_16397,N_16129,N_16198);
and U16398 (N_16398,N_16117,N_16009);
xnor U16399 (N_16399,N_16172,N_16057);
nor U16400 (N_16400,N_16375,N_16259);
and U16401 (N_16401,N_16233,N_16371);
nand U16402 (N_16402,N_16367,N_16247);
and U16403 (N_16403,N_16268,N_16280);
or U16404 (N_16404,N_16267,N_16354);
nor U16405 (N_16405,N_16316,N_16288);
nand U16406 (N_16406,N_16313,N_16258);
xnor U16407 (N_16407,N_16369,N_16349);
nor U16408 (N_16408,N_16332,N_16292);
or U16409 (N_16409,N_16307,N_16276);
xnor U16410 (N_16410,N_16327,N_16309);
and U16411 (N_16411,N_16356,N_16261);
or U16412 (N_16412,N_16346,N_16253);
xor U16413 (N_16413,N_16294,N_16363);
nor U16414 (N_16414,N_16388,N_16290);
and U16415 (N_16415,N_16321,N_16336);
nand U16416 (N_16416,N_16232,N_16291);
nand U16417 (N_16417,N_16302,N_16240);
nand U16418 (N_16418,N_16330,N_16335);
xnor U16419 (N_16419,N_16379,N_16383);
xnor U16420 (N_16420,N_16359,N_16256);
xor U16421 (N_16421,N_16389,N_16378);
or U16422 (N_16422,N_16236,N_16324);
or U16423 (N_16423,N_16216,N_16250);
or U16424 (N_16424,N_16339,N_16285);
and U16425 (N_16425,N_16395,N_16220);
nand U16426 (N_16426,N_16275,N_16281);
nor U16427 (N_16427,N_16273,N_16278);
nand U16428 (N_16428,N_16239,N_16318);
nand U16429 (N_16429,N_16264,N_16352);
xnor U16430 (N_16430,N_16237,N_16394);
nand U16431 (N_16431,N_16365,N_16252);
or U16432 (N_16432,N_16331,N_16387);
and U16433 (N_16433,N_16235,N_16296);
nor U16434 (N_16434,N_16202,N_16211);
and U16435 (N_16435,N_16301,N_16283);
or U16436 (N_16436,N_16212,N_16377);
or U16437 (N_16437,N_16209,N_16362);
nand U16438 (N_16438,N_16345,N_16266);
nand U16439 (N_16439,N_16295,N_16231);
and U16440 (N_16440,N_16246,N_16217);
nor U16441 (N_16441,N_16344,N_16287);
nand U16442 (N_16442,N_16263,N_16355);
nor U16443 (N_16443,N_16201,N_16226);
nand U16444 (N_16444,N_16257,N_16244);
nor U16445 (N_16445,N_16329,N_16342);
and U16446 (N_16446,N_16300,N_16376);
nor U16447 (N_16447,N_16282,N_16380);
and U16448 (N_16448,N_16373,N_16262);
and U16449 (N_16449,N_16277,N_16338);
nor U16450 (N_16450,N_16357,N_16207);
or U16451 (N_16451,N_16360,N_16299);
and U16452 (N_16452,N_16306,N_16272);
xor U16453 (N_16453,N_16254,N_16218);
and U16454 (N_16454,N_16398,N_16350);
or U16455 (N_16455,N_16286,N_16242);
or U16456 (N_16456,N_16390,N_16297);
or U16457 (N_16457,N_16279,N_16319);
xor U16458 (N_16458,N_16347,N_16308);
nor U16459 (N_16459,N_16215,N_16238);
xor U16460 (N_16460,N_16341,N_16314);
and U16461 (N_16461,N_16311,N_16241);
or U16462 (N_16462,N_16289,N_16204);
nand U16463 (N_16463,N_16221,N_16393);
nand U16464 (N_16464,N_16213,N_16312);
nor U16465 (N_16465,N_16337,N_16274);
xor U16466 (N_16466,N_16385,N_16391);
or U16467 (N_16467,N_16225,N_16223);
or U16468 (N_16468,N_16219,N_16234);
xnor U16469 (N_16469,N_16323,N_16305);
nor U16470 (N_16470,N_16205,N_16243);
and U16471 (N_16471,N_16298,N_16397);
and U16472 (N_16472,N_16326,N_16228);
nor U16473 (N_16473,N_16353,N_16333);
and U16474 (N_16474,N_16200,N_16251);
nor U16475 (N_16475,N_16304,N_16374);
nor U16476 (N_16476,N_16269,N_16271);
nand U16477 (N_16477,N_16399,N_16325);
nand U16478 (N_16478,N_16203,N_16224);
xnor U16479 (N_16479,N_16248,N_16364);
or U16480 (N_16480,N_16293,N_16265);
xor U16481 (N_16481,N_16372,N_16208);
nor U16482 (N_16482,N_16386,N_16229);
nand U16483 (N_16483,N_16361,N_16366);
nand U16484 (N_16484,N_16222,N_16284);
nand U16485 (N_16485,N_16255,N_16343);
or U16486 (N_16486,N_16310,N_16351);
nor U16487 (N_16487,N_16227,N_16245);
xor U16488 (N_16488,N_16340,N_16249);
or U16489 (N_16489,N_16322,N_16303);
and U16490 (N_16490,N_16315,N_16230);
xor U16491 (N_16491,N_16370,N_16270);
nand U16492 (N_16492,N_16358,N_16348);
nor U16493 (N_16493,N_16206,N_16382);
xnor U16494 (N_16494,N_16381,N_16334);
or U16495 (N_16495,N_16214,N_16392);
or U16496 (N_16496,N_16396,N_16384);
and U16497 (N_16497,N_16320,N_16210);
nand U16498 (N_16498,N_16368,N_16328);
xnor U16499 (N_16499,N_16260,N_16317);
or U16500 (N_16500,N_16321,N_16233);
or U16501 (N_16501,N_16396,N_16381);
nor U16502 (N_16502,N_16342,N_16290);
or U16503 (N_16503,N_16298,N_16271);
nor U16504 (N_16504,N_16387,N_16226);
nor U16505 (N_16505,N_16289,N_16224);
nor U16506 (N_16506,N_16284,N_16382);
nand U16507 (N_16507,N_16336,N_16262);
and U16508 (N_16508,N_16254,N_16284);
or U16509 (N_16509,N_16358,N_16302);
nor U16510 (N_16510,N_16249,N_16279);
or U16511 (N_16511,N_16228,N_16218);
and U16512 (N_16512,N_16296,N_16389);
nor U16513 (N_16513,N_16328,N_16389);
or U16514 (N_16514,N_16232,N_16272);
nand U16515 (N_16515,N_16358,N_16237);
nand U16516 (N_16516,N_16321,N_16339);
nand U16517 (N_16517,N_16329,N_16350);
xnor U16518 (N_16518,N_16398,N_16304);
and U16519 (N_16519,N_16283,N_16240);
nand U16520 (N_16520,N_16351,N_16221);
nor U16521 (N_16521,N_16398,N_16390);
or U16522 (N_16522,N_16392,N_16377);
and U16523 (N_16523,N_16320,N_16286);
xor U16524 (N_16524,N_16248,N_16280);
nor U16525 (N_16525,N_16343,N_16367);
or U16526 (N_16526,N_16350,N_16225);
or U16527 (N_16527,N_16363,N_16226);
and U16528 (N_16528,N_16243,N_16286);
nand U16529 (N_16529,N_16254,N_16288);
nor U16530 (N_16530,N_16213,N_16304);
and U16531 (N_16531,N_16375,N_16333);
and U16532 (N_16532,N_16253,N_16345);
xnor U16533 (N_16533,N_16298,N_16311);
nor U16534 (N_16534,N_16268,N_16285);
or U16535 (N_16535,N_16367,N_16238);
nor U16536 (N_16536,N_16252,N_16339);
nand U16537 (N_16537,N_16236,N_16278);
nor U16538 (N_16538,N_16323,N_16294);
nor U16539 (N_16539,N_16331,N_16263);
xor U16540 (N_16540,N_16239,N_16366);
nand U16541 (N_16541,N_16362,N_16375);
nor U16542 (N_16542,N_16312,N_16323);
nor U16543 (N_16543,N_16279,N_16250);
nand U16544 (N_16544,N_16225,N_16360);
or U16545 (N_16545,N_16306,N_16275);
or U16546 (N_16546,N_16278,N_16261);
nand U16547 (N_16547,N_16395,N_16310);
xnor U16548 (N_16548,N_16320,N_16253);
and U16549 (N_16549,N_16260,N_16375);
and U16550 (N_16550,N_16307,N_16321);
or U16551 (N_16551,N_16364,N_16356);
xnor U16552 (N_16552,N_16218,N_16246);
or U16553 (N_16553,N_16326,N_16238);
nor U16554 (N_16554,N_16256,N_16217);
xor U16555 (N_16555,N_16276,N_16300);
and U16556 (N_16556,N_16364,N_16218);
or U16557 (N_16557,N_16292,N_16365);
or U16558 (N_16558,N_16308,N_16284);
or U16559 (N_16559,N_16315,N_16251);
and U16560 (N_16560,N_16261,N_16245);
nor U16561 (N_16561,N_16224,N_16348);
and U16562 (N_16562,N_16310,N_16274);
or U16563 (N_16563,N_16230,N_16390);
or U16564 (N_16564,N_16330,N_16288);
xor U16565 (N_16565,N_16245,N_16291);
nor U16566 (N_16566,N_16377,N_16200);
nand U16567 (N_16567,N_16296,N_16242);
xnor U16568 (N_16568,N_16335,N_16210);
xnor U16569 (N_16569,N_16348,N_16375);
xor U16570 (N_16570,N_16274,N_16284);
xor U16571 (N_16571,N_16333,N_16218);
xnor U16572 (N_16572,N_16254,N_16268);
or U16573 (N_16573,N_16259,N_16293);
nor U16574 (N_16574,N_16371,N_16311);
or U16575 (N_16575,N_16368,N_16216);
and U16576 (N_16576,N_16297,N_16250);
nand U16577 (N_16577,N_16279,N_16358);
nand U16578 (N_16578,N_16364,N_16278);
nor U16579 (N_16579,N_16332,N_16274);
xor U16580 (N_16580,N_16245,N_16308);
nand U16581 (N_16581,N_16293,N_16268);
and U16582 (N_16582,N_16392,N_16348);
nand U16583 (N_16583,N_16227,N_16317);
or U16584 (N_16584,N_16226,N_16355);
nor U16585 (N_16585,N_16317,N_16364);
and U16586 (N_16586,N_16226,N_16364);
nor U16587 (N_16587,N_16211,N_16254);
nand U16588 (N_16588,N_16214,N_16237);
nor U16589 (N_16589,N_16253,N_16340);
nand U16590 (N_16590,N_16366,N_16207);
or U16591 (N_16591,N_16375,N_16281);
nor U16592 (N_16592,N_16238,N_16277);
nor U16593 (N_16593,N_16228,N_16225);
and U16594 (N_16594,N_16321,N_16228);
nor U16595 (N_16595,N_16325,N_16266);
nor U16596 (N_16596,N_16363,N_16202);
or U16597 (N_16597,N_16382,N_16390);
xnor U16598 (N_16598,N_16215,N_16362);
nor U16599 (N_16599,N_16273,N_16316);
or U16600 (N_16600,N_16592,N_16412);
xor U16601 (N_16601,N_16548,N_16468);
xor U16602 (N_16602,N_16541,N_16529);
and U16603 (N_16603,N_16503,N_16436);
or U16604 (N_16604,N_16440,N_16465);
or U16605 (N_16605,N_16509,N_16579);
and U16606 (N_16606,N_16535,N_16450);
xnor U16607 (N_16607,N_16558,N_16499);
or U16608 (N_16608,N_16464,N_16457);
and U16609 (N_16609,N_16447,N_16474);
xnor U16610 (N_16610,N_16595,N_16556);
nand U16611 (N_16611,N_16437,N_16476);
xnor U16612 (N_16612,N_16555,N_16434);
nand U16613 (N_16613,N_16430,N_16431);
or U16614 (N_16614,N_16545,N_16517);
and U16615 (N_16615,N_16415,N_16526);
xor U16616 (N_16616,N_16454,N_16534);
nor U16617 (N_16617,N_16574,N_16424);
nor U16618 (N_16618,N_16439,N_16432);
nor U16619 (N_16619,N_16562,N_16533);
nand U16620 (N_16620,N_16513,N_16570);
nand U16621 (N_16621,N_16560,N_16504);
and U16622 (N_16622,N_16527,N_16467);
and U16623 (N_16623,N_16404,N_16460);
or U16624 (N_16624,N_16400,N_16403);
or U16625 (N_16625,N_16530,N_16470);
or U16626 (N_16626,N_16572,N_16566);
nor U16627 (N_16627,N_16591,N_16512);
or U16628 (N_16628,N_16571,N_16428);
and U16629 (N_16629,N_16506,N_16448);
xnor U16630 (N_16630,N_16563,N_16525);
nor U16631 (N_16631,N_16475,N_16473);
and U16632 (N_16632,N_16542,N_16588);
or U16633 (N_16633,N_16416,N_16502);
xor U16634 (N_16634,N_16401,N_16443);
and U16635 (N_16635,N_16406,N_16564);
or U16636 (N_16636,N_16445,N_16480);
nand U16637 (N_16637,N_16441,N_16472);
nor U16638 (N_16638,N_16522,N_16510);
or U16639 (N_16639,N_16586,N_16455);
xor U16640 (N_16640,N_16422,N_16581);
nor U16641 (N_16641,N_16553,N_16420);
nand U16642 (N_16642,N_16575,N_16557);
nor U16643 (N_16643,N_16459,N_16429);
nor U16644 (N_16644,N_16584,N_16521);
nor U16645 (N_16645,N_16461,N_16410);
or U16646 (N_16646,N_16550,N_16485);
nand U16647 (N_16647,N_16539,N_16484);
nor U16648 (N_16648,N_16407,N_16402);
nand U16649 (N_16649,N_16554,N_16446);
nor U16650 (N_16650,N_16479,N_16515);
nor U16651 (N_16651,N_16507,N_16598);
and U16652 (N_16652,N_16537,N_16419);
xor U16653 (N_16653,N_16456,N_16466);
nor U16654 (N_16654,N_16453,N_16409);
xor U16655 (N_16655,N_16489,N_16481);
nor U16656 (N_16656,N_16451,N_16494);
and U16657 (N_16657,N_16486,N_16421);
xnor U16658 (N_16658,N_16577,N_16496);
and U16659 (N_16659,N_16435,N_16508);
xnor U16660 (N_16660,N_16552,N_16546);
and U16661 (N_16661,N_16549,N_16589);
and U16662 (N_16662,N_16491,N_16559);
nand U16663 (N_16663,N_16565,N_16569);
and U16664 (N_16664,N_16442,N_16423);
nor U16665 (N_16665,N_16493,N_16418);
xor U16666 (N_16666,N_16543,N_16590);
nand U16667 (N_16667,N_16544,N_16417);
nand U16668 (N_16668,N_16599,N_16452);
nor U16669 (N_16669,N_16462,N_16488);
and U16670 (N_16670,N_16408,N_16578);
and U16671 (N_16671,N_16532,N_16528);
nand U16672 (N_16672,N_16449,N_16501);
xnor U16673 (N_16673,N_16413,N_16444);
and U16674 (N_16674,N_16523,N_16478);
nand U16675 (N_16675,N_16568,N_16538);
or U16676 (N_16676,N_16540,N_16483);
xnor U16677 (N_16677,N_16585,N_16433);
and U16678 (N_16678,N_16438,N_16547);
and U16679 (N_16679,N_16500,N_16593);
or U16680 (N_16680,N_16531,N_16458);
and U16681 (N_16681,N_16427,N_16519);
nor U16682 (N_16682,N_16597,N_16520);
and U16683 (N_16683,N_16469,N_16536);
or U16684 (N_16684,N_16411,N_16573);
or U16685 (N_16685,N_16587,N_16505);
nand U16686 (N_16686,N_16582,N_16490);
nand U16687 (N_16687,N_16487,N_16498);
nor U16688 (N_16688,N_16463,N_16567);
nand U16689 (N_16689,N_16583,N_16596);
nand U16690 (N_16690,N_16551,N_16561);
and U16691 (N_16691,N_16495,N_16477);
and U16692 (N_16692,N_16511,N_16594);
or U16693 (N_16693,N_16514,N_16516);
nand U16694 (N_16694,N_16524,N_16580);
nor U16695 (N_16695,N_16471,N_16576);
and U16696 (N_16696,N_16518,N_16497);
or U16697 (N_16697,N_16425,N_16405);
nor U16698 (N_16698,N_16482,N_16414);
and U16699 (N_16699,N_16426,N_16492);
xor U16700 (N_16700,N_16462,N_16434);
and U16701 (N_16701,N_16577,N_16567);
nor U16702 (N_16702,N_16545,N_16535);
or U16703 (N_16703,N_16573,N_16496);
and U16704 (N_16704,N_16470,N_16414);
xor U16705 (N_16705,N_16599,N_16402);
nand U16706 (N_16706,N_16479,N_16540);
nand U16707 (N_16707,N_16533,N_16461);
nand U16708 (N_16708,N_16502,N_16521);
or U16709 (N_16709,N_16420,N_16514);
nor U16710 (N_16710,N_16509,N_16594);
or U16711 (N_16711,N_16436,N_16514);
or U16712 (N_16712,N_16544,N_16492);
and U16713 (N_16713,N_16599,N_16411);
and U16714 (N_16714,N_16453,N_16408);
or U16715 (N_16715,N_16472,N_16442);
or U16716 (N_16716,N_16413,N_16400);
nand U16717 (N_16717,N_16583,N_16519);
nor U16718 (N_16718,N_16442,N_16530);
and U16719 (N_16719,N_16576,N_16434);
xnor U16720 (N_16720,N_16435,N_16556);
nor U16721 (N_16721,N_16590,N_16575);
nand U16722 (N_16722,N_16545,N_16431);
xnor U16723 (N_16723,N_16430,N_16408);
xor U16724 (N_16724,N_16422,N_16409);
nor U16725 (N_16725,N_16502,N_16571);
nor U16726 (N_16726,N_16409,N_16561);
xor U16727 (N_16727,N_16430,N_16559);
nor U16728 (N_16728,N_16517,N_16427);
nor U16729 (N_16729,N_16441,N_16452);
xor U16730 (N_16730,N_16516,N_16406);
nor U16731 (N_16731,N_16441,N_16456);
and U16732 (N_16732,N_16501,N_16513);
nand U16733 (N_16733,N_16434,N_16509);
nor U16734 (N_16734,N_16542,N_16568);
or U16735 (N_16735,N_16590,N_16514);
and U16736 (N_16736,N_16515,N_16566);
nand U16737 (N_16737,N_16419,N_16560);
and U16738 (N_16738,N_16546,N_16496);
nor U16739 (N_16739,N_16448,N_16543);
and U16740 (N_16740,N_16544,N_16511);
or U16741 (N_16741,N_16420,N_16558);
nor U16742 (N_16742,N_16592,N_16568);
nand U16743 (N_16743,N_16567,N_16459);
and U16744 (N_16744,N_16440,N_16526);
xor U16745 (N_16745,N_16562,N_16559);
and U16746 (N_16746,N_16455,N_16488);
or U16747 (N_16747,N_16451,N_16454);
and U16748 (N_16748,N_16444,N_16476);
and U16749 (N_16749,N_16576,N_16444);
xor U16750 (N_16750,N_16574,N_16405);
and U16751 (N_16751,N_16475,N_16415);
nand U16752 (N_16752,N_16596,N_16448);
xor U16753 (N_16753,N_16473,N_16545);
nand U16754 (N_16754,N_16573,N_16480);
xor U16755 (N_16755,N_16596,N_16552);
xnor U16756 (N_16756,N_16539,N_16488);
xnor U16757 (N_16757,N_16561,N_16555);
and U16758 (N_16758,N_16485,N_16446);
nor U16759 (N_16759,N_16586,N_16564);
nor U16760 (N_16760,N_16576,N_16486);
nand U16761 (N_16761,N_16573,N_16515);
nor U16762 (N_16762,N_16402,N_16416);
or U16763 (N_16763,N_16505,N_16523);
and U16764 (N_16764,N_16498,N_16574);
and U16765 (N_16765,N_16521,N_16505);
nor U16766 (N_16766,N_16473,N_16530);
or U16767 (N_16767,N_16541,N_16599);
nor U16768 (N_16768,N_16520,N_16514);
nand U16769 (N_16769,N_16521,N_16513);
xnor U16770 (N_16770,N_16564,N_16503);
and U16771 (N_16771,N_16581,N_16536);
nor U16772 (N_16772,N_16437,N_16416);
xor U16773 (N_16773,N_16453,N_16593);
nor U16774 (N_16774,N_16438,N_16536);
or U16775 (N_16775,N_16579,N_16462);
or U16776 (N_16776,N_16494,N_16427);
nor U16777 (N_16777,N_16420,N_16415);
nor U16778 (N_16778,N_16527,N_16414);
nor U16779 (N_16779,N_16522,N_16495);
nor U16780 (N_16780,N_16431,N_16406);
xnor U16781 (N_16781,N_16409,N_16448);
or U16782 (N_16782,N_16482,N_16551);
and U16783 (N_16783,N_16450,N_16581);
and U16784 (N_16784,N_16578,N_16503);
xnor U16785 (N_16785,N_16553,N_16446);
xnor U16786 (N_16786,N_16410,N_16541);
nand U16787 (N_16787,N_16543,N_16574);
or U16788 (N_16788,N_16465,N_16454);
xor U16789 (N_16789,N_16498,N_16545);
nor U16790 (N_16790,N_16479,N_16459);
nand U16791 (N_16791,N_16541,N_16423);
and U16792 (N_16792,N_16508,N_16412);
xor U16793 (N_16793,N_16505,N_16558);
nand U16794 (N_16794,N_16496,N_16501);
nand U16795 (N_16795,N_16521,N_16489);
nand U16796 (N_16796,N_16507,N_16561);
xnor U16797 (N_16797,N_16474,N_16542);
nor U16798 (N_16798,N_16563,N_16460);
or U16799 (N_16799,N_16543,N_16562);
nor U16800 (N_16800,N_16777,N_16726);
xor U16801 (N_16801,N_16663,N_16637);
nand U16802 (N_16802,N_16759,N_16639);
or U16803 (N_16803,N_16679,N_16641);
nand U16804 (N_16804,N_16769,N_16657);
xor U16805 (N_16805,N_16647,N_16733);
and U16806 (N_16806,N_16660,N_16666);
xnor U16807 (N_16807,N_16682,N_16675);
nor U16808 (N_16808,N_16686,N_16772);
xor U16809 (N_16809,N_16738,N_16775);
xor U16810 (N_16810,N_16692,N_16767);
or U16811 (N_16811,N_16763,N_16762);
and U16812 (N_16812,N_16753,N_16618);
or U16813 (N_16813,N_16701,N_16783);
nand U16814 (N_16814,N_16799,N_16661);
nor U16815 (N_16815,N_16635,N_16620);
or U16816 (N_16816,N_16626,N_16795);
nor U16817 (N_16817,N_16741,N_16774);
nor U16818 (N_16818,N_16765,N_16751);
nor U16819 (N_16819,N_16724,N_16625);
nand U16820 (N_16820,N_16739,N_16685);
nand U16821 (N_16821,N_16671,N_16714);
nor U16822 (N_16822,N_16691,N_16720);
and U16823 (N_16823,N_16645,N_16782);
nand U16824 (N_16824,N_16735,N_16638);
or U16825 (N_16825,N_16667,N_16621);
nor U16826 (N_16826,N_16788,N_16622);
nor U16827 (N_16827,N_16796,N_16707);
nand U16828 (N_16828,N_16601,N_16676);
nand U16829 (N_16829,N_16728,N_16611);
nor U16830 (N_16830,N_16754,N_16654);
or U16831 (N_16831,N_16662,N_16732);
nor U16832 (N_16832,N_16764,N_16719);
nor U16833 (N_16833,N_16604,N_16652);
or U16834 (N_16834,N_16656,N_16619);
nand U16835 (N_16835,N_16697,N_16655);
nor U16836 (N_16836,N_16642,N_16624);
or U16837 (N_16837,N_16602,N_16628);
nand U16838 (N_16838,N_16756,N_16723);
and U16839 (N_16839,N_16630,N_16790);
nor U16840 (N_16840,N_16784,N_16718);
and U16841 (N_16841,N_16649,N_16646);
and U16842 (N_16842,N_16644,N_16722);
and U16843 (N_16843,N_16704,N_16617);
or U16844 (N_16844,N_16731,N_16632);
and U16845 (N_16845,N_16746,N_16768);
and U16846 (N_16846,N_16750,N_16710);
or U16847 (N_16847,N_16658,N_16648);
and U16848 (N_16848,N_16672,N_16789);
or U16849 (N_16849,N_16687,N_16740);
and U16850 (N_16850,N_16744,N_16755);
and U16851 (N_16851,N_16778,N_16605);
nand U16852 (N_16852,N_16794,N_16716);
and U16853 (N_16853,N_16757,N_16627);
nand U16854 (N_16854,N_16677,N_16608);
nor U16855 (N_16855,N_16695,N_16609);
nand U16856 (N_16856,N_16737,N_16792);
or U16857 (N_16857,N_16631,N_16734);
nand U16858 (N_16858,N_16725,N_16636);
nor U16859 (N_16859,N_16643,N_16706);
nand U16860 (N_16860,N_16702,N_16694);
nand U16861 (N_16861,N_16696,N_16700);
nand U16862 (N_16862,N_16779,N_16607);
nor U16863 (N_16863,N_16717,N_16758);
or U16864 (N_16864,N_16711,N_16708);
nor U16865 (N_16865,N_16773,N_16771);
nand U16866 (N_16866,N_16776,N_16729);
xnor U16867 (N_16867,N_16681,N_16747);
nor U16868 (N_16868,N_16673,N_16743);
nor U16869 (N_16869,N_16623,N_16703);
xnor U16870 (N_16870,N_16610,N_16709);
nor U16871 (N_16871,N_16651,N_16640);
xnor U16872 (N_16872,N_16705,N_16749);
or U16873 (N_16873,N_16606,N_16785);
xnor U16874 (N_16874,N_16633,N_16698);
or U16875 (N_16875,N_16787,N_16665);
and U16876 (N_16876,N_16727,N_16693);
or U16877 (N_16877,N_16791,N_16683);
xnor U16878 (N_16878,N_16684,N_16634);
nand U16879 (N_16879,N_16670,N_16615);
xor U16880 (N_16880,N_16600,N_16650);
and U16881 (N_16881,N_16664,N_16699);
or U16882 (N_16882,N_16786,N_16668);
nor U16883 (N_16883,N_16674,N_16669);
xor U16884 (N_16884,N_16742,N_16616);
xor U16885 (N_16885,N_16730,N_16793);
nand U16886 (N_16886,N_16770,N_16612);
xnor U16887 (N_16887,N_16712,N_16659);
and U16888 (N_16888,N_16736,N_16745);
nand U16889 (N_16889,N_16761,N_16766);
nor U16890 (N_16890,N_16798,N_16613);
xor U16891 (N_16891,N_16781,N_16680);
nand U16892 (N_16892,N_16688,N_16614);
or U16893 (N_16893,N_16748,N_16678);
nand U16894 (N_16894,N_16752,N_16689);
xnor U16895 (N_16895,N_16713,N_16690);
nor U16896 (N_16896,N_16780,N_16797);
xor U16897 (N_16897,N_16629,N_16603);
or U16898 (N_16898,N_16721,N_16715);
nor U16899 (N_16899,N_16653,N_16760);
nor U16900 (N_16900,N_16741,N_16743);
or U16901 (N_16901,N_16747,N_16684);
nor U16902 (N_16902,N_16630,N_16622);
xor U16903 (N_16903,N_16721,N_16767);
xnor U16904 (N_16904,N_16782,N_16634);
and U16905 (N_16905,N_16690,N_16665);
or U16906 (N_16906,N_16710,N_16726);
nor U16907 (N_16907,N_16699,N_16644);
or U16908 (N_16908,N_16764,N_16767);
or U16909 (N_16909,N_16755,N_16618);
xor U16910 (N_16910,N_16708,N_16608);
xnor U16911 (N_16911,N_16768,N_16662);
nor U16912 (N_16912,N_16652,N_16720);
or U16913 (N_16913,N_16620,N_16757);
and U16914 (N_16914,N_16645,N_16630);
nand U16915 (N_16915,N_16786,N_16771);
nand U16916 (N_16916,N_16686,N_16670);
or U16917 (N_16917,N_16769,N_16740);
xnor U16918 (N_16918,N_16735,N_16696);
nor U16919 (N_16919,N_16730,N_16768);
xor U16920 (N_16920,N_16791,N_16626);
nand U16921 (N_16921,N_16634,N_16762);
and U16922 (N_16922,N_16619,N_16620);
or U16923 (N_16923,N_16770,N_16696);
xor U16924 (N_16924,N_16627,N_16662);
xnor U16925 (N_16925,N_16779,N_16675);
nor U16926 (N_16926,N_16636,N_16733);
xor U16927 (N_16927,N_16780,N_16675);
nand U16928 (N_16928,N_16644,N_16696);
nor U16929 (N_16929,N_16788,N_16694);
and U16930 (N_16930,N_16720,N_16722);
xnor U16931 (N_16931,N_16612,N_16775);
xor U16932 (N_16932,N_16650,N_16632);
or U16933 (N_16933,N_16659,N_16717);
or U16934 (N_16934,N_16792,N_16794);
nor U16935 (N_16935,N_16667,N_16642);
and U16936 (N_16936,N_16761,N_16665);
nand U16937 (N_16937,N_16709,N_16724);
or U16938 (N_16938,N_16629,N_16743);
nor U16939 (N_16939,N_16621,N_16672);
nor U16940 (N_16940,N_16634,N_16796);
nor U16941 (N_16941,N_16776,N_16631);
nand U16942 (N_16942,N_16643,N_16738);
nor U16943 (N_16943,N_16752,N_16624);
or U16944 (N_16944,N_16691,N_16791);
nand U16945 (N_16945,N_16672,N_16632);
or U16946 (N_16946,N_16688,N_16726);
xor U16947 (N_16947,N_16738,N_16642);
nor U16948 (N_16948,N_16769,N_16702);
xnor U16949 (N_16949,N_16795,N_16647);
or U16950 (N_16950,N_16603,N_16663);
or U16951 (N_16951,N_16642,N_16634);
and U16952 (N_16952,N_16621,N_16724);
nor U16953 (N_16953,N_16656,N_16691);
nor U16954 (N_16954,N_16748,N_16766);
nand U16955 (N_16955,N_16714,N_16720);
or U16956 (N_16956,N_16778,N_16666);
nand U16957 (N_16957,N_16660,N_16759);
xor U16958 (N_16958,N_16767,N_16671);
nand U16959 (N_16959,N_16714,N_16624);
nand U16960 (N_16960,N_16629,N_16694);
xnor U16961 (N_16961,N_16636,N_16797);
nor U16962 (N_16962,N_16790,N_16703);
nor U16963 (N_16963,N_16601,N_16641);
or U16964 (N_16964,N_16617,N_16691);
nand U16965 (N_16965,N_16685,N_16733);
nor U16966 (N_16966,N_16665,N_16758);
xor U16967 (N_16967,N_16758,N_16790);
nand U16968 (N_16968,N_16638,N_16673);
nor U16969 (N_16969,N_16643,N_16600);
xor U16970 (N_16970,N_16623,N_16727);
nor U16971 (N_16971,N_16723,N_16604);
or U16972 (N_16972,N_16655,N_16680);
nand U16973 (N_16973,N_16671,N_16756);
and U16974 (N_16974,N_16655,N_16760);
or U16975 (N_16975,N_16634,N_16670);
or U16976 (N_16976,N_16641,N_16736);
and U16977 (N_16977,N_16777,N_16704);
nor U16978 (N_16978,N_16640,N_16702);
nand U16979 (N_16979,N_16799,N_16736);
or U16980 (N_16980,N_16616,N_16608);
and U16981 (N_16981,N_16745,N_16616);
nand U16982 (N_16982,N_16791,N_16718);
xor U16983 (N_16983,N_16776,N_16778);
nand U16984 (N_16984,N_16772,N_16607);
nand U16985 (N_16985,N_16737,N_16640);
nand U16986 (N_16986,N_16665,N_16735);
xor U16987 (N_16987,N_16680,N_16763);
or U16988 (N_16988,N_16666,N_16674);
nand U16989 (N_16989,N_16604,N_16655);
nand U16990 (N_16990,N_16733,N_16762);
and U16991 (N_16991,N_16790,N_16781);
xor U16992 (N_16992,N_16709,N_16700);
nor U16993 (N_16993,N_16772,N_16688);
xnor U16994 (N_16994,N_16756,N_16780);
nand U16995 (N_16995,N_16610,N_16663);
xor U16996 (N_16996,N_16734,N_16743);
nand U16997 (N_16997,N_16604,N_16660);
xor U16998 (N_16998,N_16782,N_16779);
nor U16999 (N_16999,N_16708,N_16605);
xnor U17000 (N_17000,N_16819,N_16992);
nand U17001 (N_17001,N_16919,N_16849);
and U17002 (N_17002,N_16874,N_16808);
nor U17003 (N_17003,N_16902,N_16830);
or U17004 (N_17004,N_16951,N_16876);
or U17005 (N_17005,N_16920,N_16841);
nor U17006 (N_17006,N_16944,N_16851);
xnor U17007 (N_17007,N_16837,N_16866);
or U17008 (N_17008,N_16893,N_16887);
nor U17009 (N_17009,N_16987,N_16946);
nand U17010 (N_17010,N_16848,N_16958);
xor U17011 (N_17011,N_16882,N_16976);
nor U17012 (N_17012,N_16910,N_16859);
xnor U17013 (N_17013,N_16969,N_16817);
and U17014 (N_17014,N_16991,N_16818);
or U17015 (N_17015,N_16840,N_16867);
xor U17016 (N_17016,N_16843,N_16947);
or U17017 (N_17017,N_16993,N_16900);
nor U17018 (N_17018,N_16803,N_16895);
and U17019 (N_17019,N_16928,N_16988);
and U17020 (N_17020,N_16917,N_16941);
xnor U17021 (N_17021,N_16875,N_16839);
nor U17022 (N_17022,N_16945,N_16989);
and U17023 (N_17023,N_16912,N_16929);
xor U17024 (N_17024,N_16968,N_16978);
or U17025 (N_17025,N_16967,N_16909);
xnor U17026 (N_17026,N_16986,N_16926);
nor U17027 (N_17027,N_16886,N_16800);
nand U17028 (N_17028,N_16956,N_16964);
and U17029 (N_17029,N_16975,N_16972);
or U17030 (N_17030,N_16854,N_16970);
nor U17031 (N_17031,N_16834,N_16889);
nand U17032 (N_17032,N_16911,N_16881);
xor U17033 (N_17033,N_16921,N_16804);
or U17034 (N_17034,N_16953,N_16807);
and U17035 (N_17035,N_16943,N_16813);
nand U17036 (N_17036,N_16828,N_16927);
nand U17037 (N_17037,N_16961,N_16995);
nor U17038 (N_17038,N_16864,N_16999);
nor U17039 (N_17039,N_16857,N_16948);
xnor U17040 (N_17040,N_16997,N_16963);
xnor U17041 (N_17041,N_16855,N_16858);
and U17042 (N_17042,N_16957,N_16962);
nor U17043 (N_17043,N_16979,N_16844);
nand U17044 (N_17044,N_16907,N_16905);
xnor U17045 (N_17045,N_16934,N_16894);
xnor U17046 (N_17046,N_16810,N_16823);
xnor U17047 (N_17047,N_16838,N_16884);
and U17048 (N_17048,N_16862,N_16896);
and U17049 (N_17049,N_16842,N_16960);
or U17050 (N_17050,N_16850,N_16890);
and U17051 (N_17051,N_16996,N_16897);
nand U17052 (N_17052,N_16801,N_16899);
and U17053 (N_17053,N_16936,N_16846);
nor U17054 (N_17054,N_16898,N_16878);
nor U17055 (N_17055,N_16816,N_16952);
nand U17056 (N_17056,N_16901,N_16809);
and U17057 (N_17057,N_16937,N_16935);
or U17058 (N_17058,N_16938,N_16932);
nand U17059 (N_17059,N_16994,N_16930);
nand U17060 (N_17060,N_16853,N_16959);
xnor U17061 (N_17061,N_16802,N_16922);
nand U17062 (N_17062,N_16847,N_16832);
or U17063 (N_17063,N_16871,N_16868);
nor U17064 (N_17064,N_16998,N_16990);
and U17065 (N_17065,N_16860,N_16865);
or U17066 (N_17066,N_16981,N_16908);
xnor U17067 (N_17067,N_16833,N_16852);
nand U17068 (N_17068,N_16820,N_16913);
nor U17069 (N_17069,N_16982,N_16915);
xnor U17070 (N_17070,N_16924,N_16955);
xnor U17071 (N_17071,N_16931,N_16892);
or U17072 (N_17072,N_16845,N_16836);
and U17073 (N_17073,N_16906,N_16983);
nor U17074 (N_17074,N_16873,N_16984);
nand U17075 (N_17075,N_16950,N_16940);
nand U17076 (N_17076,N_16806,N_16965);
nand U17077 (N_17077,N_16966,N_16904);
and U17078 (N_17078,N_16980,N_16916);
nand U17079 (N_17079,N_16914,N_16933);
xnor U17080 (N_17080,N_16925,N_16821);
and U17081 (N_17081,N_16877,N_16835);
xor U17082 (N_17082,N_16880,N_16977);
nor U17083 (N_17083,N_16923,N_16826);
or U17084 (N_17084,N_16815,N_16973);
xor U17085 (N_17085,N_16812,N_16971);
nor U17086 (N_17086,N_16861,N_16939);
xor U17087 (N_17087,N_16811,N_16856);
nor U17088 (N_17088,N_16824,N_16872);
nand U17089 (N_17089,N_16974,N_16891);
or U17090 (N_17090,N_16827,N_16825);
nand U17091 (N_17091,N_16954,N_16883);
or U17092 (N_17092,N_16903,N_16869);
or U17093 (N_17093,N_16879,N_16985);
and U17094 (N_17094,N_16829,N_16831);
nand U17095 (N_17095,N_16805,N_16863);
xnor U17096 (N_17096,N_16918,N_16949);
xor U17097 (N_17097,N_16885,N_16888);
xor U17098 (N_17098,N_16822,N_16942);
or U17099 (N_17099,N_16814,N_16870);
nand U17100 (N_17100,N_16920,N_16888);
or U17101 (N_17101,N_16878,N_16972);
or U17102 (N_17102,N_16973,N_16978);
and U17103 (N_17103,N_16900,N_16894);
nand U17104 (N_17104,N_16876,N_16903);
or U17105 (N_17105,N_16817,N_16821);
or U17106 (N_17106,N_16828,N_16860);
nand U17107 (N_17107,N_16853,N_16988);
and U17108 (N_17108,N_16854,N_16828);
nor U17109 (N_17109,N_16932,N_16887);
and U17110 (N_17110,N_16890,N_16847);
nor U17111 (N_17111,N_16882,N_16958);
xor U17112 (N_17112,N_16887,N_16934);
or U17113 (N_17113,N_16981,N_16970);
nand U17114 (N_17114,N_16942,N_16851);
and U17115 (N_17115,N_16966,N_16864);
and U17116 (N_17116,N_16869,N_16820);
nor U17117 (N_17117,N_16906,N_16804);
and U17118 (N_17118,N_16812,N_16928);
and U17119 (N_17119,N_16885,N_16855);
or U17120 (N_17120,N_16921,N_16892);
nor U17121 (N_17121,N_16893,N_16979);
xnor U17122 (N_17122,N_16914,N_16840);
nand U17123 (N_17123,N_16830,N_16834);
nor U17124 (N_17124,N_16844,N_16806);
and U17125 (N_17125,N_16863,N_16976);
xor U17126 (N_17126,N_16979,N_16859);
and U17127 (N_17127,N_16870,N_16918);
and U17128 (N_17128,N_16833,N_16930);
and U17129 (N_17129,N_16969,N_16944);
nand U17130 (N_17130,N_16895,N_16842);
and U17131 (N_17131,N_16813,N_16921);
nand U17132 (N_17132,N_16951,N_16910);
nand U17133 (N_17133,N_16967,N_16807);
or U17134 (N_17134,N_16808,N_16806);
nor U17135 (N_17135,N_16818,N_16894);
nor U17136 (N_17136,N_16916,N_16882);
nand U17137 (N_17137,N_16932,N_16927);
and U17138 (N_17138,N_16887,N_16818);
xor U17139 (N_17139,N_16882,N_16872);
or U17140 (N_17140,N_16839,N_16993);
or U17141 (N_17141,N_16878,N_16994);
and U17142 (N_17142,N_16930,N_16855);
nor U17143 (N_17143,N_16822,N_16923);
xnor U17144 (N_17144,N_16946,N_16913);
nand U17145 (N_17145,N_16967,N_16800);
or U17146 (N_17146,N_16961,N_16956);
nor U17147 (N_17147,N_16843,N_16952);
and U17148 (N_17148,N_16954,N_16996);
or U17149 (N_17149,N_16926,N_16946);
nand U17150 (N_17150,N_16863,N_16830);
nand U17151 (N_17151,N_16855,N_16903);
xor U17152 (N_17152,N_16862,N_16866);
xnor U17153 (N_17153,N_16918,N_16877);
nor U17154 (N_17154,N_16827,N_16805);
nand U17155 (N_17155,N_16834,N_16969);
or U17156 (N_17156,N_16914,N_16874);
nor U17157 (N_17157,N_16972,N_16933);
nand U17158 (N_17158,N_16885,N_16886);
nor U17159 (N_17159,N_16803,N_16923);
or U17160 (N_17160,N_16868,N_16907);
nand U17161 (N_17161,N_16980,N_16823);
xor U17162 (N_17162,N_16848,N_16820);
or U17163 (N_17163,N_16978,N_16809);
nand U17164 (N_17164,N_16844,N_16913);
and U17165 (N_17165,N_16934,N_16944);
xnor U17166 (N_17166,N_16909,N_16970);
and U17167 (N_17167,N_16959,N_16806);
or U17168 (N_17168,N_16906,N_16835);
nor U17169 (N_17169,N_16957,N_16828);
nor U17170 (N_17170,N_16903,N_16910);
xor U17171 (N_17171,N_16812,N_16804);
or U17172 (N_17172,N_16905,N_16957);
or U17173 (N_17173,N_16935,N_16883);
or U17174 (N_17174,N_16886,N_16905);
or U17175 (N_17175,N_16815,N_16928);
or U17176 (N_17176,N_16810,N_16839);
nand U17177 (N_17177,N_16869,N_16990);
and U17178 (N_17178,N_16990,N_16843);
nor U17179 (N_17179,N_16981,N_16840);
xnor U17180 (N_17180,N_16940,N_16866);
xor U17181 (N_17181,N_16886,N_16992);
or U17182 (N_17182,N_16824,N_16930);
nand U17183 (N_17183,N_16833,N_16953);
and U17184 (N_17184,N_16867,N_16804);
and U17185 (N_17185,N_16991,N_16905);
xor U17186 (N_17186,N_16957,N_16890);
nand U17187 (N_17187,N_16835,N_16833);
xnor U17188 (N_17188,N_16926,N_16863);
and U17189 (N_17189,N_16968,N_16871);
and U17190 (N_17190,N_16898,N_16984);
xor U17191 (N_17191,N_16928,N_16927);
nand U17192 (N_17192,N_16860,N_16819);
xor U17193 (N_17193,N_16916,N_16965);
or U17194 (N_17194,N_16893,N_16996);
nand U17195 (N_17195,N_16976,N_16851);
nand U17196 (N_17196,N_16948,N_16885);
nand U17197 (N_17197,N_16804,N_16855);
or U17198 (N_17198,N_16871,N_16867);
xnor U17199 (N_17199,N_16933,N_16909);
xor U17200 (N_17200,N_17106,N_17121);
and U17201 (N_17201,N_17104,N_17110);
nor U17202 (N_17202,N_17012,N_17189);
xnor U17203 (N_17203,N_17082,N_17063);
and U17204 (N_17204,N_17031,N_17034);
nand U17205 (N_17205,N_17113,N_17092);
nand U17206 (N_17206,N_17051,N_17125);
and U17207 (N_17207,N_17075,N_17022);
nand U17208 (N_17208,N_17112,N_17146);
nand U17209 (N_17209,N_17054,N_17001);
xnor U17210 (N_17210,N_17013,N_17118);
and U17211 (N_17211,N_17158,N_17002);
nor U17212 (N_17212,N_17066,N_17008);
or U17213 (N_17213,N_17076,N_17058);
nor U17214 (N_17214,N_17086,N_17103);
xor U17215 (N_17215,N_17045,N_17087);
nor U17216 (N_17216,N_17175,N_17192);
xnor U17217 (N_17217,N_17043,N_17027);
and U17218 (N_17218,N_17056,N_17047);
and U17219 (N_17219,N_17028,N_17078);
nor U17220 (N_17220,N_17041,N_17156);
xor U17221 (N_17221,N_17074,N_17138);
nand U17222 (N_17222,N_17169,N_17162);
nor U17223 (N_17223,N_17036,N_17044);
nor U17224 (N_17224,N_17049,N_17166);
nand U17225 (N_17225,N_17065,N_17159);
and U17226 (N_17226,N_17079,N_17141);
nand U17227 (N_17227,N_17177,N_17186);
and U17228 (N_17228,N_17135,N_17130);
or U17229 (N_17229,N_17137,N_17193);
xnor U17230 (N_17230,N_17160,N_17199);
or U17231 (N_17231,N_17173,N_17139);
xnor U17232 (N_17232,N_17010,N_17134);
and U17233 (N_17233,N_17144,N_17070);
xnor U17234 (N_17234,N_17191,N_17014);
nand U17235 (N_17235,N_17198,N_17009);
or U17236 (N_17236,N_17029,N_17185);
nor U17237 (N_17237,N_17196,N_17171);
or U17238 (N_17238,N_17060,N_17107);
xor U17239 (N_17239,N_17163,N_17046);
or U17240 (N_17240,N_17083,N_17108);
and U17241 (N_17241,N_17181,N_17197);
and U17242 (N_17242,N_17109,N_17064);
and U17243 (N_17243,N_17088,N_17085);
or U17244 (N_17244,N_17072,N_17111);
or U17245 (N_17245,N_17055,N_17168);
nand U17246 (N_17246,N_17006,N_17155);
nor U17247 (N_17247,N_17067,N_17127);
nand U17248 (N_17248,N_17039,N_17030);
and U17249 (N_17249,N_17164,N_17021);
or U17250 (N_17250,N_17093,N_17061);
nor U17251 (N_17251,N_17000,N_17119);
nor U17252 (N_17252,N_17182,N_17132);
nor U17253 (N_17253,N_17140,N_17099);
nand U17254 (N_17254,N_17004,N_17142);
xnor U17255 (N_17255,N_17151,N_17037);
xor U17256 (N_17256,N_17080,N_17183);
and U17257 (N_17257,N_17091,N_17069);
or U17258 (N_17258,N_17025,N_17084);
nand U17259 (N_17259,N_17023,N_17005);
and U17260 (N_17260,N_17120,N_17026);
xnor U17261 (N_17261,N_17090,N_17187);
xnor U17262 (N_17262,N_17143,N_17167);
nand U17263 (N_17263,N_17035,N_17117);
and U17264 (N_17264,N_17095,N_17170);
xor U17265 (N_17265,N_17101,N_17032);
nand U17266 (N_17266,N_17020,N_17015);
nor U17267 (N_17267,N_17100,N_17194);
nand U17268 (N_17268,N_17161,N_17081);
nand U17269 (N_17269,N_17126,N_17073);
nand U17270 (N_17270,N_17068,N_17042);
nand U17271 (N_17271,N_17048,N_17102);
nor U17272 (N_17272,N_17153,N_17131);
or U17273 (N_17273,N_17003,N_17180);
and U17274 (N_17274,N_17040,N_17178);
nor U17275 (N_17275,N_17007,N_17129);
nand U17276 (N_17276,N_17053,N_17097);
nand U17277 (N_17277,N_17059,N_17077);
xor U17278 (N_17278,N_17024,N_17145);
or U17279 (N_17279,N_17157,N_17115);
and U17280 (N_17280,N_17184,N_17174);
nand U17281 (N_17281,N_17147,N_17172);
nand U17282 (N_17282,N_17116,N_17050);
nand U17283 (N_17283,N_17190,N_17122);
xor U17284 (N_17284,N_17057,N_17128);
and U17285 (N_17285,N_17089,N_17123);
and U17286 (N_17286,N_17136,N_17154);
or U17287 (N_17287,N_17038,N_17176);
and U17288 (N_17288,N_17150,N_17017);
or U17289 (N_17289,N_17149,N_17033);
xnor U17290 (N_17290,N_17165,N_17124);
and U17291 (N_17291,N_17114,N_17195);
or U17292 (N_17292,N_17098,N_17188);
nand U17293 (N_17293,N_17152,N_17052);
nand U17294 (N_17294,N_17105,N_17071);
and U17295 (N_17295,N_17148,N_17018);
nand U17296 (N_17296,N_17133,N_17062);
or U17297 (N_17297,N_17016,N_17179);
nand U17298 (N_17298,N_17096,N_17011);
and U17299 (N_17299,N_17094,N_17019);
nor U17300 (N_17300,N_17198,N_17160);
or U17301 (N_17301,N_17101,N_17172);
or U17302 (N_17302,N_17192,N_17051);
xnor U17303 (N_17303,N_17042,N_17152);
nand U17304 (N_17304,N_17117,N_17063);
or U17305 (N_17305,N_17123,N_17022);
or U17306 (N_17306,N_17111,N_17089);
xnor U17307 (N_17307,N_17057,N_17180);
or U17308 (N_17308,N_17045,N_17040);
and U17309 (N_17309,N_17096,N_17104);
or U17310 (N_17310,N_17067,N_17142);
xnor U17311 (N_17311,N_17161,N_17186);
xnor U17312 (N_17312,N_17072,N_17050);
nor U17313 (N_17313,N_17012,N_17106);
or U17314 (N_17314,N_17127,N_17074);
xor U17315 (N_17315,N_17064,N_17189);
or U17316 (N_17316,N_17165,N_17075);
and U17317 (N_17317,N_17097,N_17190);
xor U17318 (N_17318,N_17049,N_17143);
xnor U17319 (N_17319,N_17159,N_17007);
and U17320 (N_17320,N_17013,N_17149);
nand U17321 (N_17321,N_17086,N_17017);
or U17322 (N_17322,N_17020,N_17116);
xnor U17323 (N_17323,N_17172,N_17103);
or U17324 (N_17324,N_17004,N_17191);
xor U17325 (N_17325,N_17025,N_17138);
or U17326 (N_17326,N_17061,N_17083);
and U17327 (N_17327,N_17018,N_17086);
nor U17328 (N_17328,N_17103,N_17097);
nor U17329 (N_17329,N_17022,N_17163);
nor U17330 (N_17330,N_17048,N_17069);
and U17331 (N_17331,N_17033,N_17160);
xor U17332 (N_17332,N_17099,N_17094);
or U17333 (N_17333,N_17142,N_17171);
nand U17334 (N_17334,N_17147,N_17048);
and U17335 (N_17335,N_17183,N_17184);
or U17336 (N_17336,N_17053,N_17178);
nor U17337 (N_17337,N_17092,N_17147);
xor U17338 (N_17338,N_17095,N_17189);
and U17339 (N_17339,N_17066,N_17006);
nor U17340 (N_17340,N_17155,N_17048);
nand U17341 (N_17341,N_17077,N_17076);
and U17342 (N_17342,N_17193,N_17036);
nor U17343 (N_17343,N_17069,N_17112);
or U17344 (N_17344,N_17067,N_17198);
and U17345 (N_17345,N_17087,N_17068);
nor U17346 (N_17346,N_17150,N_17193);
nand U17347 (N_17347,N_17150,N_17174);
nor U17348 (N_17348,N_17113,N_17142);
and U17349 (N_17349,N_17035,N_17149);
nor U17350 (N_17350,N_17071,N_17114);
xor U17351 (N_17351,N_17090,N_17149);
or U17352 (N_17352,N_17091,N_17005);
nand U17353 (N_17353,N_17113,N_17052);
or U17354 (N_17354,N_17134,N_17153);
nor U17355 (N_17355,N_17165,N_17121);
xor U17356 (N_17356,N_17057,N_17110);
and U17357 (N_17357,N_17176,N_17167);
or U17358 (N_17358,N_17048,N_17043);
xnor U17359 (N_17359,N_17123,N_17186);
and U17360 (N_17360,N_17150,N_17133);
or U17361 (N_17361,N_17051,N_17179);
xor U17362 (N_17362,N_17165,N_17022);
and U17363 (N_17363,N_17087,N_17106);
or U17364 (N_17364,N_17129,N_17120);
xor U17365 (N_17365,N_17185,N_17140);
xor U17366 (N_17366,N_17155,N_17037);
or U17367 (N_17367,N_17083,N_17137);
xnor U17368 (N_17368,N_17056,N_17148);
or U17369 (N_17369,N_17017,N_17173);
nand U17370 (N_17370,N_17075,N_17120);
xor U17371 (N_17371,N_17116,N_17102);
or U17372 (N_17372,N_17144,N_17059);
or U17373 (N_17373,N_17029,N_17015);
nor U17374 (N_17374,N_17190,N_17038);
xnor U17375 (N_17375,N_17139,N_17022);
nor U17376 (N_17376,N_17005,N_17077);
or U17377 (N_17377,N_17031,N_17111);
nand U17378 (N_17378,N_17084,N_17110);
or U17379 (N_17379,N_17143,N_17067);
xnor U17380 (N_17380,N_17102,N_17157);
nand U17381 (N_17381,N_17070,N_17078);
and U17382 (N_17382,N_17141,N_17033);
nor U17383 (N_17383,N_17034,N_17029);
nand U17384 (N_17384,N_17102,N_17089);
nor U17385 (N_17385,N_17177,N_17141);
nor U17386 (N_17386,N_17104,N_17199);
or U17387 (N_17387,N_17161,N_17195);
xnor U17388 (N_17388,N_17130,N_17093);
and U17389 (N_17389,N_17129,N_17143);
nand U17390 (N_17390,N_17005,N_17012);
and U17391 (N_17391,N_17128,N_17129);
or U17392 (N_17392,N_17165,N_17047);
xnor U17393 (N_17393,N_17137,N_17021);
nor U17394 (N_17394,N_17014,N_17138);
nand U17395 (N_17395,N_17162,N_17066);
or U17396 (N_17396,N_17122,N_17036);
xor U17397 (N_17397,N_17068,N_17063);
or U17398 (N_17398,N_17193,N_17039);
nand U17399 (N_17399,N_17037,N_17043);
xor U17400 (N_17400,N_17370,N_17337);
nand U17401 (N_17401,N_17314,N_17395);
nor U17402 (N_17402,N_17378,N_17359);
xnor U17403 (N_17403,N_17248,N_17243);
nand U17404 (N_17404,N_17207,N_17204);
nand U17405 (N_17405,N_17299,N_17300);
nand U17406 (N_17406,N_17317,N_17377);
nor U17407 (N_17407,N_17316,N_17352);
xor U17408 (N_17408,N_17290,N_17350);
and U17409 (N_17409,N_17227,N_17263);
nor U17410 (N_17410,N_17323,N_17235);
nor U17411 (N_17411,N_17387,N_17342);
nand U17412 (N_17412,N_17238,N_17222);
and U17413 (N_17413,N_17333,N_17216);
or U17414 (N_17414,N_17285,N_17247);
xor U17415 (N_17415,N_17295,N_17205);
and U17416 (N_17416,N_17324,N_17214);
xor U17417 (N_17417,N_17381,N_17393);
nand U17418 (N_17418,N_17312,N_17375);
and U17419 (N_17419,N_17327,N_17215);
or U17420 (N_17420,N_17209,N_17362);
nor U17421 (N_17421,N_17335,N_17201);
nand U17422 (N_17422,N_17261,N_17355);
or U17423 (N_17423,N_17357,N_17231);
xnor U17424 (N_17424,N_17360,N_17331);
nor U17425 (N_17425,N_17294,N_17217);
nand U17426 (N_17426,N_17341,N_17384);
nand U17427 (N_17427,N_17250,N_17276);
xnor U17428 (N_17428,N_17218,N_17274);
and U17429 (N_17429,N_17221,N_17275);
or U17430 (N_17430,N_17332,N_17338);
nand U17431 (N_17431,N_17347,N_17219);
nand U17432 (N_17432,N_17373,N_17344);
nor U17433 (N_17433,N_17225,N_17311);
and U17434 (N_17434,N_17380,N_17367);
and U17435 (N_17435,N_17330,N_17297);
nand U17436 (N_17436,N_17315,N_17226);
or U17437 (N_17437,N_17280,N_17291);
nor U17438 (N_17438,N_17394,N_17246);
nand U17439 (N_17439,N_17282,N_17202);
xnor U17440 (N_17440,N_17266,N_17322);
xnor U17441 (N_17441,N_17346,N_17211);
or U17442 (N_17442,N_17281,N_17398);
xor U17443 (N_17443,N_17302,N_17309);
nand U17444 (N_17444,N_17369,N_17329);
and U17445 (N_17445,N_17240,N_17307);
and U17446 (N_17446,N_17364,N_17358);
and U17447 (N_17447,N_17265,N_17392);
nor U17448 (N_17448,N_17348,N_17228);
nand U17449 (N_17449,N_17289,N_17356);
nor U17450 (N_17450,N_17249,N_17339);
and U17451 (N_17451,N_17366,N_17229);
or U17452 (N_17452,N_17328,N_17386);
or U17453 (N_17453,N_17257,N_17340);
nor U17454 (N_17454,N_17354,N_17223);
or U17455 (N_17455,N_17368,N_17382);
xor U17456 (N_17456,N_17371,N_17365);
nor U17457 (N_17457,N_17208,N_17230);
or U17458 (N_17458,N_17267,N_17212);
and U17459 (N_17459,N_17255,N_17391);
nor U17460 (N_17460,N_17353,N_17272);
nor U17461 (N_17461,N_17237,N_17220);
xnor U17462 (N_17462,N_17308,N_17304);
nand U17463 (N_17463,N_17376,N_17251);
and U17464 (N_17464,N_17320,N_17245);
or U17465 (N_17465,N_17306,N_17264);
nand U17466 (N_17466,N_17241,N_17279);
nor U17467 (N_17467,N_17325,N_17236);
nand U17468 (N_17468,N_17396,N_17349);
xor U17469 (N_17469,N_17262,N_17200);
nor U17470 (N_17470,N_17379,N_17234);
nor U17471 (N_17471,N_17292,N_17305);
or U17472 (N_17472,N_17390,N_17326);
nor U17473 (N_17473,N_17287,N_17210);
nor U17474 (N_17474,N_17372,N_17318);
or U17475 (N_17475,N_17239,N_17268);
nand U17476 (N_17476,N_17258,N_17363);
nand U17477 (N_17477,N_17397,N_17233);
nor U17478 (N_17478,N_17389,N_17343);
nand U17479 (N_17479,N_17303,N_17399);
and U17480 (N_17480,N_17313,N_17345);
nor U17481 (N_17481,N_17259,N_17361);
xnor U17482 (N_17482,N_17277,N_17224);
xnor U17483 (N_17483,N_17269,N_17203);
nand U17484 (N_17484,N_17213,N_17301);
and U17485 (N_17485,N_17244,N_17283);
xnor U17486 (N_17486,N_17284,N_17252);
and U17487 (N_17487,N_17310,N_17288);
or U17488 (N_17488,N_17383,N_17374);
or U17489 (N_17489,N_17298,N_17351);
or U17490 (N_17490,N_17242,N_17385);
xnor U17491 (N_17491,N_17278,N_17296);
and U17492 (N_17492,N_17336,N_17319);
nor U17493 (N_17493,N_17270,N_17260);
xor U17494 (N_17494,N_17256,N_17206);
xor U17495 (N_17495,N_17286,N_17334);
nand U17496 (N_17496,N_17271,N_17293);
and U17497 (N_17497,N_17253,N_17388);
nand U17498 (N_17498,N_17273,N_17254);
or U17499 (N_17499,N_17232,N_17321);
nand U17500 (N_17500,N_17366,N_17397);
nand U17501 (N_17501,N_17267,N_17286);
nand U17502 (N_17502,N_17393,N_17289);
nor U17503 (N_17503,N_17286,N_17332);
nor U17504 (N_17504,N_17353,N_17204);
and U17505 (N_17505,N_17359,N_17351);
or U17506 (N_17506,N_17269,N_17370);
xor U17507 (N_17507,N_17305,N_17375);
nand U17508 (N_17508,N_17257,N_17366);
nor U17509 (N_17509,N_17228,N_17396);
or U17510 (N_17510,N_17222,N_17205);
nand U17511 (N_17511,N_17286,N_17333);
nor U17512 (N_17512,N_17347,N_17324);
and U17513 (N_17513,N_17307,N_17232);
nand U17514 (N_17514,N_17264,N_17325);
xor U17515 (N_17515,N_17273,N_17232);
nor U17516 (N_17516,N_17251,N_17230);
xor U17517 (N_17517,N_17298,N_17221);
nand U17518 (N_17518,N_17344,N_17298);
xor U17519 (N_17519,N_17389,N_17232);
nor U17520 (N_17520,N_17222,N_17231);
nor U17521 (N_17521,N_17279,N_17349);
xnor U17522 (N_17522,N_17380,N_17294);
or U17523 (N_17523,N_17315,N_17271);
and U17524 (N_17524,N_17282,N_17359);
nand U17525 (N_17525,N_17384,N_17328);
nor U17526 (N_17526,N_17218,N_17280);
xnor U17527 (N_17527,N_17296,N_17386);
and U17528 (N_17528,N_17220,N_17353);
xor U17529 (N_17529,N_17243,N_17327);
and U17530 (N_17530,N_17380,N_17314);
nor U17531 (N_17531,N_17314,N_17324);
nand U17532 (N_17532,N_17319,N_17299);
and U17533 (N_17533,N_17242,N_17266);
and U17534 (N_17534,N_17355,N_17393);
and U17535 (N_17535,N_17399,N_17204);
nor U17536 (N_17536,N_17213,N_17345);
nand U17537 (N_17537,N_17200,N_17214);
and U17538 (N_17538,N_17397,N_17241);
nand U17539 (N_17539,N_17217,N_17277);
nor U17540 (N_17540,N_17385,N_17205);
and U17541 (N_17541,N_17227,N_17220);
nor U17542 (N_17542,N_17391,N_17341);
nor U17543 (N_17543,N_17297,N_17226);
or U17544 (N_17544,N_17275,N_17358);
nand U17545 (N_17545,N_17330,N_17271);
or U17546 (N_17546,N_17265,N_17365);
nand U17547 (N_17547,N_17341,N_17356);
nor U17548 (N_17548,N_17282,N_17394);
or U17549 (N_17549,N_17384,N_17343);
and U17550 (N_17550,N_17317,N_17316);
xor U17551 (N_17551,N_17241,N_17366);
nand U17552 (N_17552,N_17222,N_17279);
nand U17553 (N_17553,N_17212,N_17225);
xor U17554 (N_17554,N_17298,N_17347);
nor U17555 (N_17555,N_17306,N_17252);
nand U17556 (N_17556,N_17239,N_17345);
nor U17557 (N_17557,N_17352,N_17231);
nand U17558 (N_17558,N_17297,N_17263);
or U17559 (N_17559,N_17273,N_17356);
xor U17560 (N_17560,N_17303,N_17261);
and U17561 (N_17561,N_17319,N_17284);
xor U17562 (N_17562,N_17275,N_17249);
nand U17563 (N_17563,N_17227,N_17266);
and U17564 (N_17564,N_17209,N_17288);
or U17565 (N_17565,N_17283,N_17371);
nor U17566 (N_17566,N_17340,N_17384);
or U17567 (N_17567,N_17324,N_17282);
and U17568 (N_17568,N_17314,N_17292);
and U17569 (N_17569,N_17359,N_17330);
nand U17570 (N_17570,N_17313,N_17247);
nand U17571 (N_17571,N_17304,N_17290);
nor U17572 (N_17572,N_17317,N_17239);
xor U17573 (N_17573,N_17291,N_17273);
or U17574 (N_17574,N_17265,N_17282);
xnor U17575 (N_17575,N_17229,N_17394);
nand U17576 (N_17576,N_17267,N_17399);
xor U17577 (N_17577,N_17272,N_17342);
nand U17578 (N_17578,N_17310,N_17337);
nor U17579 (N_17579,N_17399,N_17222);
nand U17580 (N_17580,N_17332,N_17310);
and U17581 (N_17581,N_17283,N_17297);
xor U17582 (N_17582,N_17319,N_17255);
and U17583 (N_17583,N_17254,N_17238);
nor U17584 (N_17584,N_17235,N_17319);
nor U17585 (N_17585,N_17286,N_17346);
or U17586 (N_17586,N_17335,N_17255);
and U17587 (N_17587,N_17282,N_17355);
xor U17588 (N_17588,N_17346,N_17290);
or U17589 (N_17589,N_17384,N_17267);
and U17590 (N_17590,N_17380,N_17372);
nand U17591 (N_17591,N_17282,N_17205);
or U17592 (N_17592,N_17282,N_17354);
or U17593 (N_17593,N_17312,N_17323);
nor U17594 (N_17594,N_17333,N_17319);
nand U17595 (N_17595,N_17315,N_17258);
and U17596 (N_17596,N_17232,N_17395);
nand U17597 (N_17597,N_17243,N_17384);
or U17598 (N_17598,N_17325,N_17334);
nor U17599 (N_17599,N_17354,N_17362);
nor U17600 (N_17600,N_17529,N_17434);
or U17601 (N_17601,N_17401,N_17427);
nor U17602 (N_17602,N_17483,N_17486);
nand U17603 (N_17603,N_17585,N_17597);
or U17604 (N_17604,N_17418,N_17420);
nand U17605 (N_17605,N_17556,N_17506);
xor U17606 (N_17606,N_17410,N_17553);
nand U17607 (N_17607,N_17503,N_17587);
nor U17608 (N_17608,N_17572,N_17406);
nand U17609 (N_17609,N_17546,N_17534);
or U17610 (N_17610,N_17538,N_17424);
nand U17611 (N_17611,N_17568,N_17554);
or U17612 (N_17612,N_17552,N_17471);
nand U17613 (N_17613,N_17561,N_17579);
and U17614 (N_17614,N_17594,N_17555);
nor U17615 (N_17615,N_17515,N_17576);
nand U17616 (N_17616,N_17590,N_17468);
nand U17617 (N_17617,N_17445,N_17516);
xnor U17618 (N_17618,N_17433,N_17425);
nand U17619 (N_17619,N_17584,N_17415);
nor U17620 (N_17620,N_17484,N_17409);
xor U17621 (N_17621,N_17442,N_17599);
nand U17622 (N_17622,N_17545,N_17493);
or U17623 (N_17623,N_17480,N_17520);
and U17624 (N_17624,N_17531,N_17522);
and U17625 (N_17625,N_17446,N_17513);
or U17626 (N_17626,N_17500,N_17492);
and U17627 (N_17627,N_17537,N_17494);
xnor U17628 (N_17628,N_17559,N_17571);
nand U17629 (N_17629,N_17426,N_17472);
xnor U17630 (N_17630,N_17477,N_17439);
nor U17631 (N_17631,N_17595,N_17438);
nand U17632 (N_17632,N_17535,N_17449);
nor U17633 (N_17633,N_17466,N_17532);
or U17634 (N_17634,N_17491,N_17527);
nor U17635 (N_17635,N_17470,N_17586);
nor U17636 (N_17636,N_17578,N_17429);
or U17637 (N_17637,N_17573,N_17588);
or U17638 (N_17638,N_17411,N_17521);
xor U17639 (N_17639,N_17509,N_17465);
and U17640 (N_17640,N_17510,N_17469);
nand U17641 (N_17641,N_17455,N_17569);
and U17642 (N_17642,N_17505,N_17580);
nand U17643 (N_17643,N_17489,N_17575);
or U17644 (N_17644,N_17462,N_17591);
xor U17645 (N_17645,N_17478,N_17453);
and U17646 (N_17646,N_17400,N_17541);
nand U17647 (N_17647,N_17507,N_17593);
nor U17648 (N_17648,N_17524,N_17536);
xor U17649 (N_17649,N_17581,N_17560);
nand U17650 (N_17650,N_17540,N_17460);
nor U17651 (N_17651,N_17511,N_17435);
or U17652 (N_17652,N_17564,N_17436);
nand U17653 (N_17653,N_17430,N_17502);
or U17654 (N_17654,N_17562,N_17563);
nor U17655 (N_17655,N_17582,N_17499);
xor U17656 (N_17656,N_17421,N_17539);
nor U17657 (N_17657,N_17475,N_17543);
nor U17658 (N_17658,N_17551,N_17598);
xnor U17659 (N_17659,N_17482,N_17452);
or U17660 (N_17660,N_17405,N_17495);
nand U17661 (N_17661,N_17428,N_17577);
or U17662 (N_17662,N_17432,N_17403);
or U17663 (N_17663,N_17416,N_17451);
and U17664 (N_17664,N_17419,N_17504);
nor U17665 (N_17665,N_17414,N_17437);
xnor U17666 (N_17666,N_17558,N_17565);
nor U17667 (N_17667,N_17431,N_17530);
and U17668 (N_17668,N_17557,N_17518);
nand U17669 (N_17669,N_17574,N_17407);
or U17670 (N_17670,N_17456,N_17450);
nand U17671 (N_17671,N_17498,N_17473);
nand U17672 (N_17672,N_17547,N_17501);
nand U17673 (N_17673,N_17461,N_17549);
xnor U17674 (N_17674,N_17496,N_17544);
nor U17675 (N_17675,N_17443,N_17458);
nand U17676 (N_17676,N_17404,N_17441);
nand U17677 (N_17677,N_17519,N_17447);
nand U17678 (N_17678,N_17474,N_17454);
nor U17679 (N_17679,N_17481,N_17567);
nor U17680 (N_17680,N_17533,N_17589);
or U17681 (N_17681,N_17417,N_17596);
xor U17682 (N_17682,N_17592,N_17570);
xor U17683 (N_17683,N_17542,N_17423);
or U17684 (N_17684,N_17467,N_17517);
nor U17685 (N_17685,N_17525,N_17459);
nor U17686 (N_17686,N_17479,N_17550);
nand U17687 (N_17687,N_17487,N_17523);
and U17688 (N_17688,N_17408,N_17412);
nor U17689 (N_17689,N_17583,N_17402);
and U17690 (N_17690,N_17464,N_17457);
xor U17691 (N_17691,N_17476,N_17490);
nor U17692 (N_17692,N_17514,N_17413);
or U17693 (N_17693,N_17497,N_17548);
xnor U17694 (N_17694,N_17444,N_17566);
nor U17695 (N_17695,N_17512,N_17526);
nor U17696 (N_17696,N_17508,N_17463);
nand U17697 (N_17697,N_17440,N_17488);
nor U17698 (N_17698,N_17485,N_17422);
nand U17699 (N_17699,N_17528,N_17448);
or U17700 (N_17700,N_17562,N_17551);
nand U17701 (N_17701,N_17512,N_17508);
xor U17702 (N_17702,N_17450,N_17497);
nor U17703 (N_17703,N_17402,N_17469);
or U17704 (N_17704,N_17477,N_17409);
nor U17705 (N_17705,N_17556,N_17593);
nor U17706 (N_17706,N_17592,N_17523);
xor U17707 (N_17707,N_17400,N_17470);
nand U17708 (N_17708,N_17505,N_17576);
and U17709 (N_17709,N_17566,N_17555);
xnor U17710 (N_17710,N_17599,N_17415);
and U17711 (N_17711,N_17410,N_17421);
and U17712 (N_17712,N_17454,N_17494);
nor U17713 (N_17713,N_17568,N_17561);
and U17714 (N_17714,N_17410,N_17481);
or U17715 (N_17715,N_17592,N_17526);
nand U17716 (N_17716,N_17481,N_17543);
nand U17717 (N_17717,N_17571,N_17537);
xnor U17718 (N_17718,N_17417,N_17581);
xor U17719 (N_17719,N_17561,N_17443);
nand U17720 (N_17720,N_17446,N_17452);
or U17721 (N_17721,N_17409,N_17533);
or U17722 (N_17722,N_17440,N_17529);
nor U17723 (N_17723,N_17494,N_17582);
nor U17724 (N_17724,N_17595,N_17511);
nand U17725 (N_17725,N_17433,N_17589);
or U17726 (N_17726,N_17556,N_17425);
nand U17727 (N_17727,N_17515,N_17407);
nor U17728 (N_17728,N_17401,N_17426);
nand U17729 (N_17729,N_17559,N_17538);
nor U17730 (N_17730,N_17443,N_17553);
nand U17731 (N_17731,N_17450,N_17452);
and U17732 (N_17732,N_17479,N_17488);
xor U17733 (N_17733,N_17464,N_17561);
xnor U17734 (N_17734,N_17577,N_17405);
or U17735 (N_17735,N_17400,N_17543);
nor U17736 (N_17736,N_17415,N_17503);
and U17737 (N_17737,N_17483,N_17580);
nand U17738 (N_17738,N_17403,N_17429);
nor U17739 (N_17739,N_17575,N_17447);
nand U17740 (N_17740,N_17448,N_17553);
or U17741 (N_17741,N_17534,N_17522);
nor U17742 (N_17742,N_17487,N_17430);
nor U17743 (N_17743,N_17596,N_17510);
nor U17744 (N_17744,N_17480,N_17552);
or U17745 (N_17745,N_17541,N_17501);
xor U17746 (N_17746,N_17556,N_17580);
or U17747 (N_17747,N_17529,N_17563);
nand U17748 (N_17748,N_17475,N_17585);
xor U17749 (N_17749,N_17474,N_17480);
nor U17750 (N_17750,N_17579,N_17400);
xor U17751 (N_17751,N_17568,N_17483);
or U17752 (N_17752,N_17597,N_17497);
and U17753 (N_17753,N_17479,N_17572);
and U17754 (N_17754,N_17451,N_17417);
xnor U17755 (N_17755,N_17414,N_17595);
or U17756 (N_17756,N_17468,N_17577);
or U17757 (N_17757,N_17560,N_17428);
xnor U17758 (N_17758,N_17536,N_17504);
nor U17759 (N_17759,N_17536,N_17532);
or U17760 (N_17760,N_17450,N_17501);
nand U17761 (N_17761,N_17418,N_17402);
or U17762 (N_17762,N_17478,N_17580);
nand U17763 (N_17763,N_17433,N_17565);
nor U17764 (N_17764,N_17556,N_17413);
nor U17765 (N_17765,N_17491,N_17441);
or U17766 (N_17766,N_17416,N_17489);
and U17767 (N_17767,N_17524,N_17493);
nor U17768 (N_17768,N_17513,N_17449);
nand U17769 (N_17769,N_17404,N_17423);
nand U17770 (N_17770,N_17554,N_17591);
or U17771 (N_17771,N_17519,N_17589);
and U17772 (N_17772,N_17532,N_17571);
xnor U17773 (N_17773,N_17428,N_17424);
nor U17774 (N_17774,N_17421,N_17566);
xnor U17775 (N_17775,N_17457,N_17551);
nand U17776 (N_17776,N_17584,N_17465);
nor U17777 (N_17777,N_17523,N_17453);
or U17778 (N_17778,N_17509,N_17472);
xor U17779 (N_17779,N_17563,N_17555);
or U17780 (N_17780,N_17592,N_17559);
xnor U17781 (N_17781,N_17436,N_17410);
or U17782 (N_17782,N_17522,N_17438);
xnor U17783 (N_17783,N_17474,N_17523);
nor U17784 (N_17784,N_17558,N_17540);
and U17785 (N_17785,N_17559,N_17496);
or U17786 (N_17786,N_17539,N_17413);
and U17787 (N_17787,N_17577,N_17488);
or U17788 (N_17788,N_17504,N_17598);
xnor U17789 (N_17789,N_17587,N_17443);
or U17790 (N_17790,N_17594,N_17478);
or U17791 (N_17791,N_17591,N_17482);
nor U17792 (N_17792,N_17419,N_17499);
or U17793 (N_17793,N_17537,N_17518);
nand U17794 (N_17794,N_17595,N_17461);
xnor U17795 (N_17795,N_17501,N_17598);
or U17796 (N_17796,N_17419,N_17563);
nor U17797 (N_17797,N_17594,N_17472);
xnor U17798 (N_17798,N_17532,N_17503);
xnor U17799 (N_17799,N_17591,N_17436);
and U17800 (N_17800,N_17619,N_17705);
and U17801 (N_17801,N_17794,N_17731);
or U17802 (N_17802,N_17634,N_17689);
and U17803 (N_17803,N_17665,N_17788);
nand U17804 (N_17804,N_17655,N_17703);
and U17805 (N_17805,N_17625,N_17684);
or U17806 (N_17806,N_17606,N_17793);
xor U17807 (N_17807,N_17774,N_17771);
or U17808 (N_17808,N_17629,N_17679);
nand U17809 (N_17809,N_17601,N_17734);
nand U17810 (N_17810,N_17709,N_17658);
or U17811 (N_17811,N_17730,N_17674);
xnor U17812 (N_17812,N_17692,N_17700);
nor U17813 (N_17813,N_17789,N_17779);
nor U17814 (N_17814,N_17715,N_17657);
or U17815 (N_17815,N_17786,N_17668);
and U17816 (N_17816,N_17639,N_17670);
xnor U17817 (N_17817,N_17701,N_17790);
xnor U17818 (N_17818,N_17773,N_17682);
or U17819 (N_17819,N_17732,N_17743);
or U17820 (N_17820,N_17662,N_17776);
nand U17821 (N_17821,N_17765,N_17714);
nor U17822 (N_17822,N_17627,N_17744);
xnor U17823 (N_17823,N_17772,N_17628);
nor U17824 (N_17824,N_17726,N_17775);
and U17825 (N_17825,N_17667,N_17638);
xnor U17826 (N_17826,N_17623,N_17747);
nor U17827 (N_17827,N_17752,N_17769);
xnor U17828 (N_17828,N_17751,N_17637);
nor U17829 (N_17829,N_17748,N_17608);
nor U17830 (N_17830,N_17615,N_17650);
nand U17831 (N_17831,N_17652,N_17741);
or U17832 (N_17832,N_17621,N_17706);
nor U17833 (N_17833,N_17719,N_17739);
nand U17834 (N_17834,N_17704,N_17605);
nand U17835 (N_17835,N_17759,N_17720);
xor U17836 (N_17836,N_17713,N_17604);
nor U17837 (N_17837,N_17767,N_17737);
or U17838 (N_17838,N_17622,N_17696);
xnor U17839 (N_17839,N_17617,N_17718);
and U17840 (N_17840,N_17760,N_17660);
nand U17841 (N_17841,N_17653,N_17763);
and U17842 (N_17842,N_17795,N_17626);
or U17843 (N_17843,N_17644,N_17764);
nand U17844 (N_17844,N_17612,N_17680);
and U17845 (N_17845,N_17610,N_17745);
nand U17846 (N_17846,N_17783,N_17651);
and U17847 (N_17847,N_17781,N_17678);
and U17848 (N_17848,N_17780,N_17681);
or U17849 (N_17849,N_17746,N_17784);
nor U17850 (N_17850,N_17614,N_17699);
nand U17851 (N_17851,N_17787,N_17685);
xor U17852 (N_17852,N_17756,N_17636);
and U17853 (N_17853,N_17691,N_17641);
nor U17854 (N_17854,N_17669,N_17716);
xnor U17855 (N_17855,N_17796,N_17602);
or U17856 (N_17856,N_17698,N_17697);
nand U17857 (N_17857,N_17742,N_17710);
nor U17858 (N_17858,N_17792,N_17724);
and U17859 (N_17859,N_17757,N_17620);
nand U17860 (N_17860,N_17768,N_17624);
xor U17861 (N_17861,N_17717,N_17673);
or U17862 (N_17862,N_17675,N_17687);
xnor U17863 (N_17863,N_17750,N_17755);
xnor U17864 (N_17864,N_17762,N_17609);
nand U17865 (N_17865,N_17613,N_17671);
and U17866 (N_17866,N_17611,N_17708);
nand U17867 (N_17867,N_17648,N_17722);
and U17868 (N_17868,N_17618,N_17738);
xor U17869 (N_17869,N_17702,N_17753);
or U17870 (N_17870,N_17690,N_17616);
nand U17871 (N_17871,N_17729,N_17683);
nor U17872 (N_17872,N_17791,N_17666);
nand U17873 (N_17873,N_17646,N_17640);
xnor U17874 (N_17874,N_17642,N_17733);
or U17875 (N_17875,N_17631,N_17725);
or U17876 (N_17876,N_17676,N_17727);
or U17877 (N_17877,N_17607,N_17659);
xor U17878 (N_17878,N_17761,N_17600);
nand U17879 (N_17879,N_17695,N_17778);
and U17880 (N_17880,N_17677,N_17649);
nand U17881 (N_17881,N_17632,N_17693);
or U17882 (N_17882,N_17785,N_17643);
or U17883 (N_17883,N_17664,N_17712);
xor U17884 (N_17884,N_17688,N_17797);
xor U17885 (N_17885,N_17661,N_17603);
xnor U17886 (N_17886,N_17647,N_17723);
xor U17887 (N_17887,N_17758,N_17782);
and U17888 (N_17888,N_17694,N_17635);
nand U17889 (N_17889,N_17707,N_17770);
nand U17890 (N_17890,N_17777,N_17711);
xor U17891 (N_17891,N_17672,N_17740);
xor U17892 (N_17892,N_17736,N_17721);
xnor U17893 (N_17893,N_17728,N_17656);
nor U17894 (N_17894,N_17766,N_17630);
nand U17895 (N_17895,N_17654,N_17735);
nor U17896 (N_17896,N_17663,N_17686);
or U17897 (N_17897,N_17798,N_17749);
nand U17898 (N_17898,N_17645,N_17799);
xnor U17899 (N_17899,N_17633,N_17754);
and U17900 (N_17900,N_17698,N_17743);
nor U17901 (N_17901,N_17688,N_17645);
nor U17902 (N_17902,N_17747,N_17710);
nor U17903 (N_17903,N_17678,N_17790);
and U17904 (N_17904,N_17626,N_17639);
nor U17905 (N_17905,N_17715,N_17627);
nand U17906 (N_17906,N_17735,N_17646);
or U17907 (N_17907,N_17693,N_17792);
and U17908 (N_17908,N_17618,N_17620);
nor U17909 (N_17909,N_17731,N_17793);
xor U17910 (N_17910,N_17756,N_17767);
xor U17911 (N_17911,N_17693,N_17764);
nor U17912 (N_17912,N_17618,N_17735);
xor U17913 (N_17913,N_17708,N_17773);
nand U17914 (N_17914,N_17674,N_17627);
and U17915 (N_17915,N_17760,N_17604);
and U17916 (N_17916,N_17642,N_17724);
nor U17917 (N_17917,N_17641,N_17655);
nor U17918 (N_17918,N_17771,N_17790);
or U17919 (N_17919,N_17745,N_17726);
and U17920 (N_17920,N_17646,N_17687);
or U17921 (N_17921,N_17664,N_17741);
nor U17922 (N_17922,N_17764,N_17735);
nor U17923 (N_17923,N_17622,N_17733);
nand U17924 (N_17924,N_17674,N_17645);
or U17925 (N_17925,N_17646,N_17747);
nor U17926 (N_17926,N_17702,N_17736);
and U17927 (N_17927,N_17610,N_17622);
nand U17928 (N_17928,N_17600,N_17759);
nor U17929 (N_17929,N_17691,N_17707);
xnor U17930 (N_17930,N_17627,N_17702);
or U17931 (N_17931,N_17758,N_17676);
nor U17932 (N_17932,N_17706,N_17604);
nand U17933 (N_17933,N_17686,N_17773);
or U17934 (N_17934,N_17714,N_17693);
or U17935 (N_17935,N_17735,N_17727);
nor U17936 (N_17936,N_17718,N_17674);
nand U17937 (N_17937,N_17747,N_17712);
nor U17938 (N_17938,N_17635,N_17710);
xnor U17939 (N_17939,N_17623,N_17613);
or U17940 (N_17940,N_17716,N_17754);
nand U17941 (N_17941,N_17602,N_17770);
nor U17942 (N_17942,N_17667,N_17754);
nand U17943 (N_17943,N_17613,N_17642);
nor U17944 (N_17944,N_17770,N_17630);
xnor U17945 (N_17945,N_17715,N_17738);
nor U17946 (N_17946,N_17748,N_17644);
or U17947 (N_17947,N_17717,N_17601);
and U17948 (N_17948,N_17743,N_17632);
xor U17949 (N_17949,N_17712,N_17762);
xor U17950 (N_17950,N_17751,N_17710);
nand U17951 (N_17951,N_17719,N_17767);
or U17952 (N_17952,N_17761,N_17714);
and U17953 (N_17953,N_17741,N_17759);
xor U17954 (N_17954,N_17797,N_17608);
nor U17955 (N_17955,N_17720,N_17797);
nand U17956 (N_17956,N_17665,N_17787);
xnor U17957 (N_17957,N_17604,N_17733);
xor U17958 (N_17958,N_17787,N_17713);
and U17959 (N_17959,N_17641,N_17620);
nand U17960 (N_17960,N_17671,N_17752);
xor U17961 (N_17961,N_17732,N_17683);
or U17962 (N_17962,N_17628,N_17653);
xor U17963 (N_17963,N_17751,N_17683);
and U17964 (N_17964,N_17749,N_17799);
nand U17965 (N_17965,N_17660,N_17618);
or U17966 (N_17966,N_17674,N_17687);
xor U17967 (N_17967,N_17672,N_17649);
or U17968 (N_17968,N_17785,N_17738);
nand U17969 (N_17969,N_17723,N_17725);
and U17970 (N_17970,N_17715,N_17766);
nand U17971 (N_17971,N_17778,N_17688);
or U17972 (N_17972,N_17622,N_17701);
nand U17973 (N_17973,N_17778,N_17667);
or U17974 (N_17974,N_17789,N_17733);
xnor U17975 (N_17975,N_17707,N_17789);
nor U17976 (N_17976,N_17798,N_17733);
and U17977 (N_17977,N_17611,N_17765);
xor U17978 (N_17978,N_17715,N_17705);
or U17979 (N_17979,N_17728,N_17709);
or U17980 (N_17980,N_17710,N_17752);
xnor U17981 (N_17981,N_17753,N_17669);
nor U17982 (N_17982,N_17706,N_17665);
nor U17983 (N_17983,N_17637,N_17692);
or U17984 (N_17984,N_17671,N_17743);
nor U17985 (N_17985,N_17793,N_17757);
or U17986 (N_17986,N_17629,N_17726);
or U17987 (N_17987,N_17792,N_17698);
or U17988 (N_17988,N_17736,N_17606);
and U17989 (N_17989,N_17792,N_17692);
xor U17990 (N_17990,N_17650,N_17750);
and U17991 (N_17991,N_17751,N_17618);
xnor U17992 (N_17992,N_17752,N_17613);
and U17993 (N_17993,N_17741,N_17610);
nor U17994 (N_17994,N_17665,N_17662);
xnor U17995 (N_17995,N_17625,N_17719);
nor U17996 (N_17996,N_17698,N_17652);
and U17997 (N_17997,N_17797,N_17708);
nand U17998 (N_17998,N_17635,N_17650);
nor U17999 (N_17999,N_17622,N_17732);
xor U18000 (N_18000,N_17983,N_17898);
nor U18001 (N_18001,N_17840,N_17977);
xor U18002 (N_18002,N_17826,N_17903);
or U18003 (N_18003,N_17976,N_17959);
or U18004 (N_18004,N_17964,N_17955);
nand U18005 (N_18005,N_17966,N_17820);
xor U18006 (N_18006,N_17886,N_17892);
nor U18007 (N_18007,N_17878,N_17857);
nor U18008 (N_18008,N_17984,N_17987);
xnor U18009 (N_18009,N_17861,N_17875);
nand U18010 (N_18010,N_17910,N_17991);
xor U18011 (N_18011,N_17981,N_17906);
nand U18012 (N_18012,N_17992,N_17894);
nor U18013 (N_18013,N_17879,N_17994);
nor U18014 (N_18014,N_17927,N_17940);
or U18015 (N_18015,N_17869,N_17934);
and U18016 (N_18016,N_17831,N_17839);
nand U18017 (N_18017,N_17952,N_17924);
and U18018 (N_18018,N_17834,N_17939);
xnor U18019 (N_18019,N_17997,N_17816);
nand U18020 (N_18020,N_17823,N_17916);
nand U18021 (N_18021,N_17998,N_17859);
nand U18022 (N_18022,N_17836,N_17855);
or U18023 (N_18023,N_17872,N_17996);
xor U18024 (N_18024,N_17914,N_17922);
and U18025 (N_18025,N_17958,N_17841);
and U18026 (N_18026,N_17866,N_17812);
nor U18027 (N_18027,N_17936,N_17860);
nor U18028 (N_18028,N_17933,N_17900);
xor U18029 (N_18029,N_17979,N_17961);
or U18030 (N_18030,N_17871,N_17912);
nand U18031 (N_18031,N_17905,N_17867);
nand U18032 (N_18032,N_17901,N_17851);
nand U18033 (N_18033,N_17808,N_17971);
or U18034 (N_18034,N_17822,N_17956);
xnor U18035 (N_18035,N_17835,N_17809);
xnor U18036 (N_18036,N_17853,N_17868);
or U18037 (N_18037,N_17881,N_17837);
or U18038 (N_18038,N_17908,N_17990);
or U18039 (N_18039,N_17844,N_17909);
nor U18040 (N_18040,N_17843,N_17965);
xnor U18041 (N_18041,N_17802,N_17953);
xor U18042 (N_18042,N_17941,N_17932);
and U18043 (N_18043,N_17923,N_17858);
nor U18044 (N_18044,N_17842,N_17846);
or U18045 (N_18045,N_17832,N_17970);
nor U18046 (N_18046,N_17813,N_17804);
xor U18047 (N_18047,N_17899,N_17968);
xor U18048 (N_18048,N_17806,N_17951);
nand U18049 (N_18049,N_17810,N_17895);
and U18050 (N_18050,N_17944,N_17938);
xnor U18051 (N_18051,N_17975,N_17967);
xor U18052 (N_18052,N_17918,N_17830);
nor U18053 (N_18053,N_17978,N_17969);
nor U18054 (N_18054,N_17995,N_17888);
nand U18055 (N_18055,N_17874,N_17920);
and U18056 (N_18056,N_17849,N_17887);
xnor U18057 (N_18057,N_17930,N_17937);
nor U18058 (N_18058,N_17882,N_17856);
nor U18059 (N_18059,N_17960,N_17986);
xnor U18060 (N_18060,N_17957,N_17943);
nor U18061 (N_18061,N_17880,N_17948);
xnor U18062 (N_18062,N_17917,N_17902);
xor U18063 (N_18063,N_17974,N_17864);
or U18064 (N_18064,N_17825,N_17942);
and U18065 (N_18065,N_17931,N_17877);
xnor U18066 (N_18066,N_17876,N_17921);
and U18067 (N_18067,N_17985,N_17949);
and U18068 (N_18068,N_17817,N_17827);
and U18069 (N_18069,N_17862,N_17911);
nand U18070 (N_18070,N_17807,N_17821);
nor U18071 (N_18071,N_17854,N_17999);
nand U18072 (N_18072,N_17847,N_17973);
nor U18073 (N_18073,N_17889,N_17950);
and U18074 (N_18074,N_17838,N_17885);
nor U18075 (N_18075,N_17870,N_17865);
nand U18076 (N_18076,N_17926,N_17989);
nand U18077 (N_18077,N_17819,N_17891);
nand U18078 (N_18078,N_17852,N_17893);
nand U18079 (N_18079,N_17850,N_17980);
xnor U18080 (N_18080,N_17803,N_17845);
nor U18081 (N_18081,N_17815,N_17945);
and U18082 (N_18082,N_17824,N_17818);
nor U18083 (N_18083,N_17962,N_17925);
nand U18084 (N_18084,N_17801,N_17897);
or U18085 (N_18085,N_17873,N_17963);
xnor U18086 (N_18086,N_17929,N_17814);
and U18087 (N_18087,N_17833,N_17919);
nand U18088 (N_18088,N_17972,N_17883);
or U18089 (N_18089,N_17800,N_17863);
and U18090 (N_18090,N_17913,N_17993);
or U18091 (N_18091,N_17946,N_17988);
nand U18092 (N_18092,N_17805,N_17907);
xnor U18093 (N_18093,N_17884,N_17928);
or U18094 (N_18094,N_17848,N_17896);
nand U18095 (N_18095,N_17935,N_17811);
or U18096 (N_18096,N_17982,N_17954);
nand U18097 (N_18097,N_17904,N_17947);
or U18098 (N_18098,N_17915,N_17890);
and U18099 (N_18099,N_17828,N_17829);
nand U18100 (N_18100,N_17827,N_17948);
xor U18101 (N_18101,N_17819,N_17912);
and U18102 (N_18102,N_17818,N_17911);
nor U18103 (N_18103,N_17871,N_17800);
xnor U18104 (N_18104,N_17878,N_17975);
and U18105 (N_18105,N_17905,N_17819);
xor U18106 (N_18106,N_17835,N_17949);
and U18107 (N_18107,N_17803,N_17828);
or U18108 (N_18108,N_17841,N_17905);
or U18109 (N_18109,N_17956,N_17821);
and U18110 (N_18110,N_17808,N_17911);
nand U18111 (N_18111,N_17821,N_17892);
xor U18112 (N_18112,N_17889,N_17831);
nand U18113 (N_18113,N_17904,N_17984);
nand U18114 (N_18114,N_17908,N_17946);
nor U18115 (N_18115,N_17901,N_17939);
nand U18116 (N_18116,N_17804,N_17807);
nand U18117 (N_18117,N_17987,N_17883);
or U18118 (N_18118,N_17889,N_17892);
or U18119 (N_18119,N_17848,N_17814);
nand U18120 (N_18120,N_17815,N_17968);
nand U18121 (N_18121,N_17805,N_17917);
and U18122 (N_18122,N_17916,N_17892);
or U18123 (N_18123,N_17871,N_17835);
xor U18124 (N_18124,N_17899,N_17830);
nor U18125 (N_18125,N_17998,N_17946);
and U18126 (N_18126,N_17809,N_17967);
xnor U18127 (N_18127,N_17840,N_17950);
nand U18128 (N_18128,N_17959,N_17867);
or U18129 (N_18129,N_17941,N_17977);
nand U18130 (N_18130,N_17822,N_17907);
and U18131 (N_18131,N_17953,N_17862);
xnor U18132 (N_18132,N_17967,N_17880);
nand U18133 (N_18133,N_17995,N_17920);
or U18134 (N_18134,N_17978,N_17930);
nand U18135 (N_18135,N_17888,N_17880);
or U18136 (N_18136,N_17959,N_17898);
nand U18137 (N_18137,N_17853,N_17862);
nor U18138 (N_18138,N_17806,N_17873);
xor U18139 (N_18139,N_17961,N_17850);
nand U18140 (N_18140,N_17974,N_17921);
nand U18141 (N_18141,N_17928,N_17860);
nor U18142 (N_18142,N_17876,N_17843);
and U18143 (N_18143,N_17948,N_17851);
nand U18144 (N_18144,N_17928,N_17839);
or U18145 (N_18145,N_17963,N_17824);
nor U18146 (N_18146,N_17818,N_17803);
nor U18147 (N_18147,N_17951,N_17878);
nor U18148 (N_18148,N_17981,N_17878);
nor U18149 (N_18149,N_17921,N_17973);
or U18150 (N_18150,N_17860,N_17901);
nand U18151 (N_18151,N_17826,N_17861);
nand U18152 (N_18152,N_17802,N_17814);
nand U18153 (N_18153,N_17959,N_17830);
or U18154 (N_18154,N_17818,N_17826);
or U18155 (N_18155,N_17996,N_17886);
or U18156 (N_18156,N_17897,N_17959);
nor U18157 (N_18157,N_17925,N_17907);
nor U18158 (N_18158,N_17887,N_17846);
and U18159 (N_18159,N_17887,N_17999);
nor U18160 (N_18160,N_17812,N_17822);
xnor U18161 (N_18161,N_17972,N_17912);
or U18162 (N_18162,N_17854,N_17860);
nor U18163 (N_18163,N_17869,N_17836);
nor U18164 (N_18164,N_17871,N_17883);
nor U18165 (N_18165,N_17843,N_17879);
xor U18166 (N_18166,N_17988,N_17955);
nor U18167 (N_18167,N_17955,N_17808);
xnor U18168 (N_18168,N_17899,N_17824);
or U18169 (N_18169,N_17918,N_17837);
nor U18170 (N_18170,N_17801,N_17882);
and U18171 (N_18171,N_17849,N_17901);
nor U18172 (N_18172,N_17961,N_17814);
nor U18173 (N_18173,N_17933,N_17953);
or U18174 (N_18174,N_17805,N_17971);
nor U18175 (N_18175,N_17993,N_17816);
nand U18176 (N_18176,N_17980,N_17910);
xnor U18177 (N_18177,N_17867,N_17883);
nand U18178 (N_18178,N_17937,N_17808);
and U18179 (N_18179,N_17951,N_17950);
and U18180 (N_18180,N_17993,N_17809);
nor U18181 (N_18181,N_17967,N_17925);
nor U18182 (N_18182,N_17802,N_17801);
or U18183 (N_18183,N_17936,N_17998);
and U18184 (N_18184,N_17974,N_17846);
or U18185 (N_18185,N_17958,N_17892);
or U18186 (N_18186,N_17976,N_17803);
xnor U18187 (N_18187,N_17822,N_17944);
or U18188 (N_18188,N_17839,N_17939);
xor U18189 (N_18189,N_17917,N_17852);
and U18190 (N_18190,N_17859,N_17923);
nand U18191 (N_18191,N_17997,N_17979);
nor U18192 (N_18192,N_17869,N_17958);
xnor U18193 (N_18193,N_17991,N_17937);
nor U18194 (N_18194,N_17822,N_17849);
xnor U18195 (N_18195,N_17831,N_17964);
and U18196 (N_18196,N_17836,N_17963);
or U18197 (N_18197,N_17995,N_17974);
nand U18198 (N_18198,N_17989,N_17907);
nor U18199 (N_18199,N_17846,N_17937);
nand U18200 (N_18200,N_18111,N_18060);
and U18201 (N_18201,N_18101,N_18071);
xnor U18202 (N_18202,N_18154,N_18122);
nor U18203 (N_18203,N_18051,N_18164);
and U18204 (N_18204,N_18123,N_18087);
nand U18205 (N_18205,N_18094,N_18153);
and U18206 (N_18206,N_18131,N_18142);
nor U18207 (N_18207,N_18088,N_18081);
or U18208 (N_18208,N_18078,N_18039);
xor U18209 (N_18209,N_18112,N_18107);
and U18210 (N_18210,N_18037,N_18083);
xnor U18211 (N_18211,N_18196,N_18013);
nand U18212 (N_18212,N_18002,N_18027);
xor U18213 (N_18213,N_18089,N_18188);
and U18214 (N_18214,N_18128,N_18025);
or U18215 (N_18215,N_18029,N_18124);
or U18216 (N_18216,N_18022,N_18085);
or U18217 (N_18217,N_18052,N_18145);
and U18218 (N_18218,N_18017,N_18006);
and U18219 (N_18219,N_18189,N_18148);
xor U18220 (N_18220,N_18009,N_18158);
nor U18221 (N_18221,N_18028,N_18197);
or U18222 (N_18222,N_18199,N_18125);
or U18223 (N_18223,N_18066,N_18091);
or U18224 (N_18224,N_18067,N_18047);
or U18225 (N_18225,N_18043,N_18015);
and U18226 (N_18226,N_18135,N_18130);
nor U18227 (N_18227,N_18056,N_18177);
nor U18228 (N_18228,N_18031,N_18116);
nand U18229 (N_18229,N_18127,N_18173);
or U18230 (N_18230,N_18152,N_18044);
xor U18231 (N_18231,N_18167,N_18129);
and U18232 (N_18232,N_18098,N_18159);
nand U18233 (N_18233,N_18095,N_18151);
or U18234 (N_18234,N_18076,N_18113);
nor U18235 (N_18235,N_18042,N_18041);
and U18236 (N_18236,N_18063,N_18149);
and U18237 (N_18237,N_18054,N_18169);
xor U18238 (N_18238,N_18139,N_18046);
nand U18239 (N_18239,N_18133,N_18048);
xor U18240 (N_18240,N_18090,N_18064);
or U18241 (N_18241,N_18162,N_18163);
xnor U18242 (N_18242,N_18073,N_18117);
or U18243 (N_18243,N_18012,N_18156);
nor U18244 (N_18244,N_18141,N_18120);
or U18245 (N_18245,N_18126,N_18062);
or U18246 (N_18246,N_18018,N_18184);
or U18247 (N_18247,N_18106,N_18097);
xor U18248 (N_18248,N_18082,N_18070);
xnor U18249 (N_18249,N_18144,N_18166);
nor U18250 (N_18250,N_18058,N_18003);
and U18251 (N_18251,N_18165,N_18086);
xnor U18252 (N_18252,N_18143,N_18035);
and U18253 (N_18253,N_18157,N_18061);
xnor U18254 (N_18254,N_18121,N_18140);
nor U18255 (N_18255,N_18033,N_18170);
and U18256 (N_18256,N_18069,N_18146);
or U18257 (N_18257,N_18068,N_18194);
nor U18258 (N_18258,N_18072,N_18055);
and U18259 (N_18259,N_18036,N_18136);
nand U18260 (N_18260,N_18053,N_18079);
xor U18261 (N_18261,N_18134,N_18103);
xnor U18262 (N_18262,N_18114,N_18138);
nor U18263 (N_18263,N_18032,N_18110);
or U18264 (N_18264,N_18115,N_18172);
xnor U18265 (N_18265,N_18049,N_18174);
or U18266 (N_18266,N_18010,N_18118);
nand U18267 (N_18267,N_18045,N_18092);
or U18268 (N_18268,N_18147,N_18161);
xnor U18269 (N_18269,N_18004,N_18019);
xor U18270 (N_18270,N_18183,N_18191);
or U18271 (N_18271,N_18007,N_18180);
nand U18272 (N_18272,N_18150,N_18195);
and U18273 (N_18273,N_18011,N_18001);
xor U18274 (N_18274,N_18026,N_18193);
nor U18275 (N_18275,N_18020,N_18005);
nor U18276 (N_18276,N_18109,N_18059);
nor U18277 (N_18277,N_18077,N_18137);
nor U18278 (N_18278,N_18096,N_18187);
nor U18279 (N_18279,N_18168,N_18155);
nand U18280 (N_18280,N_18171,N_18016);
xor U18281 (N_18281,N_18023,N_18176);
nor U18282 (N_18282,N_18102,N_18014);
nor U18283 (N_18283,N_18099,N_18080);
nand U18284 (N_18284,N_18132,N_18057);
or U18285 (N_18285,N_18038,N_18050);
xnor U18286 (N_18286,N_18040,N_18160);
xnor U18287 (N_18287,N_18084,N_18198);
and U18288 (N_18288,N_18192,N_18021);
xor U18289 (N_18289,N_18105,N_18104);
nand U18290 (N_18290,N_18181,N_18030);
and U18291 (N_18291,N_18100,N_18074);
nand U18292 (N_18292,N_18075,N_18093);
and U18293 (N_18293,N_18008,N_18000);
xnor U18294 (N_18294,N_18179,N_18186);
xor U18295 (N_18295,N_18024,N_18178);
xnor U18296 (N_18296,N_18190,N_18185);
and U18297 (N_18297,N_18065,N_18034);
and U18298 (N_18298,N_18175,N_18119);
or U18299 (N_18299,N_18108,N_18182);
and U18300 (N_18300,N_18079,N_18067);
nor U18301 (N_18301,N_18121,N_18055);
nand U18302 (N_18302,N_18059,N_18180);
nand U18303 (N_18303,N_18058,N_18066);
nand U18304 (N_18304,N_18150,N_18069);
or U18305 (N_18305,N_18016,N_18040);
nor U18306 (N_18306,N_18044,N_18127);
nand U18307 (N_18307,N_18048,N_18197);
and U18308 (N_18308,N_18115,N_18061);
or U18309 (N_18309,N_18022,N_18145);
or U18310 (N_18310,N_18195,N_18122);
xnor U18311 (N_18311,N_18002,N_18116);
nand U18312 (N_18312,N_18025,N_18019);
nand U18313 (N_18313,N_18043,N_18092);
xnor U18314 (N_18314,N_18135,N_18094);
or U18315 (N_18315,N_18087,N_18137);
and U18316 (N_18316,N_18061,N_18070);
nor U18317 (N_18317,N_18190,N_18074);
or U18318 (N_18318,N_18117,N_18164);
and U18319 (N_18319,N_18050,N_18182);
nor U18320 (N_18320,N_18057,N_18108);
nor U18321 (N_18321,N_18052,N_18006);
or U18322 (N_18322,N_18011,N_18142);
or U18323 (N_18323,N_18160,N_18032);
nand U18324 (N_18324,N_18193,N_18019);
xnor U18325 (N_18325,N_18129,N_18008);
xor U18326 (N_18326,N_18173,N_18138);
nand U18327 (N_18327,N_18017,N_18089);
and U18328 (N_18328,N_18023,N_18039);
and U18329 (N_18329,N_18091,N_18019);
nand U18330 (N_18330,N_18029,N_18119);
nor U18331 (N_18331,N_18054,N_18058);
nand U18332 (N_18332,N_18087,N_18048);
or U18333 (N_18333,N_18182,N_18186);
nor U18334 (N_18334,N_18169,N_18113);
nor U18335 (N_18335,N_18093,N_18088);
nand U18336 (N_18336,N_18087,N_18055);
xor U18337 (N_18337,N_18090,N_18040);
nor U18338 (N_18338,N_18029,N_18096);
nand U18339 (N_18339,N_18112,N_18163);
or U18340 (N_18340,N_18165,N_18073);
nor U18341 (N_18341,N_18089,N_18038);
nor U18342 (N_18342,N_18147,N_18062);
nand U18343 (N_18343,N_18044,N_18183);
xor U18344 (N_18344,N_18037,N_18130);
or U18345 (N_18345,N_18114,N_18148);
nor U18346 (N_18346,N_18039,N_18050);
nand U18347 (N_18347,N_18124,N_18175);
xnor U18348 (N_18348,N_18108,N_18162);
nand U18349 (N_18349,N_18004,N_18126);
xor U18350 (N_18350,N_18017,N_18100);
nand U18351 (N_18351,N_18175,N_18029);
nor U18352 (N_18352,N_18014,N_18096);
xnor U18353 (N_18353,N_18183,N_18010);
and U18354 (N_18354,N_18106,N_18017);
or U18355 (N_18355,N_18114,N_18155);
nand U18356 (N_18356,N_18098,N_18074);
nor U18357 (N_18357,N_18110,N_18147);
and U18358 (N_18358,N_18171,N_18176);
nor U18359 (N_18359,N_18037,N_18199);
nand U18360 (N_18360,N_18027,N_18073);
nand U18361 (N_18361,N_18116,N_18151);
nor U18362 (N_18362,N_18016,N_18170);
xor U18363 (N_18363,N_18189,N_18185);
xnor U18364 (N_18364,N_18159,N_18039);
xnor U18365 (N_18365,N_18112,N_18110);
nor U18366 (N_18366,N_18192,N_18116);
nand U18367 (N_18367,N_18022,N_18116);
nor U18368 (N_18368,N_18023,N_18106);
or U18369 (N_18369,N_18019,N_18096);
and U18370 (N_18370,N_18099,N_18138);
xnor U18371 (N_18371,N_18154,N_18113);
xor U18372 (N_18372,N_18105,N_18170);
and U18373 (N_18373,N_18124,N_18197);
nand U18374 (N_18374,N_18001,N_18174);
xnor U18375 (N_18375,N_18174,N_18178);
xor U18376 (N_18376,N_18103,N_18155);
nor U18377 (N_18377,N_18107,N_18048);
and U18378 (N_18378,N_18138,N_18081);
and U18379 (N_18379,N_18031,N_18166);
or U18380 (N_18380,N_18026,N_18177);
nor U18381 (N_18381,N_18138,N_18191);
nand U18382 (N_18382,N_18109,N_18080);
xor U18383 (N_18383,N_18007,N_18078);
nand U18384 (N_18384,N_18019,N_18011);
and U18385 (N_18385,N_18086,N_18111);
nor U18386 (N_18386,N_18132,N_18134);
nor U18387 (N_18387,N_18158,N_18139);
or U18388 (N_18388,N_18145,N_18020);
nand U18389 (N_18389,N_18146,N_18178);
nor U18390 (N_18390,N_18141,N_18057);
or U18391 (N_18391,N_18178,N_18002);
nor U18392 (N_18392,N_18151,N_18078);
and U18393 (N_18393,N_18109,N_18072);
xor U18394 (N_18394,N_18124,N_18163);
nand U18395 (N_18395,N_18079,N_18161);
xor U18396 (N_18396,N_18063,N_18021);
nand U18397 (N_18397,N_18024,N_18153);
nor U18398 (N_18398,N_18033,N_18059);
and U18399 (N_18399,N_18098,N_18133);
nand U18400 (N_18400,N_18283,N_18306);
nand U18401 (N_18401,N_18243,N_18264);
and U18402 (N_18402,N_18378,N_18382);
or U18403 (N_18403,N_18200,N_18330);
nor U18404 (N_18404,N_18394,N_18300);
nand U18405 (N_18405,N_18251,N_18312);
and U18406 (N_18406,N_18343,N_18244);
nand U18407 (N_18407,N_18228,N_18274);
and U18408 (N_18408,N_18233,N_18298);
xnor U18409 (N_18409,N_18259,N_18342);
nor U18410 (N_18410,N_18326,N_18311);
nor U18411 (N_18411,N_18374,N_18285);
and U18412 (N_18412,N_18221,N_18208);
nor U18413 (N_18413,N_18230,N_18246);
nand U18414 (N_18414,N_18332,N_18391);
nor U18415 (N_18415,N_18212,N_18393);
nand U18416 (N_18416,N_18210,N_18370);
nand U18417 (N_18417,N_18254,N_18392);
or U18418 (N_18418,N_18341,N_18286);
nor U18419 (N_18419,N_18361,N_18376);
or U18420 (N_18420,N_18294,N_18339);
nand U18421 (N_18421,N_18270,N_18227);
nand U18422 (N_18422,N_18271,N_18331);
xnor U18423 (N_18423,N_18275,N_18262);
and U18424 (N_18424,N_18211,N_18247);
nor U18425 (N_18425,N_18303,N_18380);
nand U18426 (N_18426,N_18204,N_18325);
xor U18427 (N_18427,N_18241,N_18359);
or U18428 (N_18428,N_18284,N_18333);
or U18429 (N_18429,N_18201,N_18371);
nor U18430 (N_18430,N_18358,N_18373);
and U18431 (N_18431,N_18335,N_18323);
nand U18432 (N_18432,N_18320,N_18362);
nor U18433 (N_18433,N_18318,N_18209);
nand U18434 (N_18434,N_18266,N_18344);
or U18435 (N_18435,N_18304,N_18290);
or U18436 (N_18436,N_18322,N_18203);
or U18437 (N_18437,N_18336,N_18305);
and U18438 (N_18438,N_18231,N_18364);
xor U18439 (N_18439,N_18279,N_18349);
xnor U18440 (N_18440,N_18225,N_18346);
nand U18441 (N_18441,N_18315,N_18287);
or U18442 (N_18442,N_18218,N_18268);
xor U18443 (N_18443,N_18240,N_18272);
nand U18444 (N_18444,N_18278,N_18387);
or U18445 (N_18445,N_18396,N_18277);
and U18446 (N_18446,N_18232,N_18385);
or U18447 (N_18447,N_18206,N_18334);
or U18448 (N_18448,N_18224,N_18289);
nor U18449 (N_18449,N_18293,N_18355);
xor U18450 (N_18450,N_18309,N_18239);
xor U18451 (N_18451,N_18217,N_18310);
or U18452 (N_18452,N_18263,N_18255);
nand U18453 (N_18453,N_18337,N_18252);
and U18454 (N_18454,N_18237,N_18367);
and U18455 (N_18455,N_18213,N_18234);
xor U18456 (N_18456,N_18276,N_18345);
or U18457 (N_18457,N_18249,N_18398);
nor U18458 (N_18458,N_18329,N_18223);
nand U18459 (N_18459,N_18229,N_18356);
nand U18460 (N_18460,N_18348,N_18360);
nand U18461 (N_18461,N_18314,N_18395);
or U18462 (N_18462,N_18390,N_18377);
nor U18463 (N_18463,N_18316,N_18250);
nor U18464 (N_18464,N_18386,N_18215);
nand U18465 (N_18465,N_18226,N_18399);
nor U18466 (N_18466,N_18328,N_18301);
xor U18467 (N_18467,N_18384,N_18258);
nand U18468 (N_18468,N_18280,N_18256);
or U18469 (N_18469,N_18307,N_18257);
xnor U18470 (N_18470,N_18321,N_18340);
and U18471 (N_18471,N_18324,N_18375);
nor U18472 (N_18472,N_18269,N_18291);
and U18473 (N_18473,N_18261,N_18363);
or U18474 (N_18474,N_18368,N_18282);
nor U18475 (N_18475,N_18273,N_18296);
nor U18476 (N_18476,N_18216,N_18292);
and U18477 (N_18477,N_18260,N_18347);
or U18478 (N_18478,N_18338,N_18235);
nand U18479 (N_18479,N_18248,N_18288);
nand U18480 (N_18480,N_18353,N_18245);
and U18481 (N_18481,N_18319,N_18219);
and U18482 (N_18482,N_18205,N_18207);
nor U18483 (N_18483,N_18351,N_18295);
xnor U18484 (N_18484,N_18299,N_18267);
nand U18485 (N_18485,N_18297,N_18238);
or U18486 (N_18486,N_18222,N_18302);
xnor U18487 (N_18487,N_18383,N_18357);
nor U18488 (N_18488,N_18397,N_18281);
nand U18489 (N_18489,N_18365,N_18389);
nand U18490 (N_18490,N_18366,N_18214);
nor U18491 (N_18491,N_18327,N_18202);
nor U18492 (N_18492,N_18317,N_18253);
and U18493 (N_18493,N_18352,N_18381);
xnor U18494 (N_18494,N_18354,N_18369);
nor U18495 (N_18495,N_18220,N_18236);
xor U18496 (N_18496,N_18379,N_18308);
nand U18497 (N_18497,N_18388,N_18265);
nor U18498 (N_18498,N_18313,N_18242);
nand U18499 (N_18499,N_18350,N_18372);
nand U18500 (N_18500,N_18226,N_18391);
or U18501 (N_18501,N_18251,N_18217);
nor U18502 (N_18502,N_18398,N_18202);
nand U18503 (N_18503,N_18367,N_18203);
or U18504 (N_18504,N_18356,N_18237);
and U18505 (N_18505,N_18286,N_18214);
nor U18506 (N_18506,N_18283,N_18274);
or U18507 (N_18507,N_18261,N_18379);
xor U18508 (N_18508,N_18230,N_18281);
nand U18509 (N_18509,N_18362,N_18236);
nor U18510 (N_18510,N_18308,N_18289);
nor U18511 (N_18511,N_18240,N_18277);
or U18512 (N_18512,N_18222,N_18390);
nor U18513 (N_18513,N_18306,N_18302);
and U18514 (N_18514,N_18374,N_18299);
or U18515 (N_18515,N_18239,N_18219);
nor U18516 (N_18516,N_18200,N_18313);
nor U18517 (N_18517,N_18231,N_18218);
nor U18518 (N_18518,N_18217,N_18335);
xnor U18519 (N_18519,N_18319,N_18281);
or U18520 (N_18520,N_18237,N_18388);
and U18521 (N_18521,N_18335,N_18371);
nor U18522 (N_18522,N_18275,N_18226);
and U18523 (N_18523,N_18377,N_18243);
and U18524 (N_18524,N_18234,N_18252);
xnor U18525 (N_18525,N_18328,N_18348);
nor U18526 (N_18526,N_18275,N_18210);
nand U18527 (N_18527,N_18281,N_18347);
nand U18528 (N_18528,N_18309,N_18280);
nor U18529 (N_18529,N_18275,N_18261);
xor U18530 (N_18530,N_18378,N_18345);
nor U18531 (N_18531,N_18237,N_18281);
xor U18532 (N_18532,N_18301,N_18325);
or U18533 (N_18533,N_18309,N_18278);
or U18534 (N_18534,N_18357,N_18237);
or U18535 (N_18535,N_18385,N_18302);
nor U18536 (N_18536,N_18394,N_18350);
and U18537 (N_18537,N_18296,N_18287);
or U18538 (N_18538,N_18248,N_18270);
nor U18539 (N_18539,N_18369,N_18277);
nor U18540 (N_18540,N_18225,N_18388);
or U18541 (N_18541,N_18216,N_18312);
or U18542 (N_18542,N_18238,N_18318);
or U18543 (N_18543,N_18222,N_18303);
or U18544 (N_18544,N_18220,N_18266);
xor U18545 (N_18545,N_18370,N_18386);
xor U18546 (N_18546,N_18347,N_18372);
nor U18547 (N_18547,N_18358,N_18303);
and U18548 (N_18548,N_18297,N_18267);
or U18549 (N_18549,N_18372,N_18307);
and U18550 (N_18550,N_18374,N_18235);
or U18551 (N_18551,N_18356,N_18262);
and U18552 (N_18552,N_18399,N_18370);
and U18553 (N_18553,N_18393,N_18346);
nand U18554 (N_18554,N_18341,N_18239);
and U18555 (N_18555,N_18260,N_18300);
nand U18556 (N_18556,N_18358,N_18379);
and U18557 (N_18557,N_18228,N_18275);
nand U18558 (N_18558,N_18343,N_18305);
and U18559 (N_18559,N_18364,N_18212);
or U18560 (N_18560,N_18272,N_18294);
or U18561 (N_18561,N_18349,N_18211);
nor U18562 (N_18562,N_18260,N_18359);
nor U18563 (N_18563,N_18381,N_18294);
nand U18564 (N_18564,N_18254,N_18351);
and U18565 (N_18565,N_18289,N_18311);
xnor U18566 (N_18566,N_18356,N_18399);
or U18567 (N_18567,N_18268,N_18308);
xnor U18568 (N_18568,N_18291,N_18360);
and U18569 (N_18569,N_18285,N_18399);
or U18570 (N_18570,N_18213,N_18252);
xnor U18571 (N_18571,N_18265,N_18263);
nand U18572 (N_18572,N_18285,N_18348);
xor U18573 (N_18573,N_18350,N_18292);
and U18574 (N_18574,N_18215,N_18297);
xor U18575 (N_18575,N_18273,N_18218);
and U18576 (N_18576,N_18210,N_18356);
and U18577 (N_18577,N_18339,N_18285);
and U18578 (N_18578,N_18356,N_18263);
nand U18579 (N_18579,N_18325,N_18310);
xnor U18580 (N_18580,N_18262,N_18216);
xnor U18581 (N_18581,N_18316,N_18398);
xnor U18582 (N_18582,N_18277,N_18321);
or U18583 (N_18583,N_18290,N_18296);
and U18584 (N_18584,N_18317,N_18275);
or U18585 (N_18585,N_18217,N_18358);
nor U18586 (N_18586,N_18341,N_18289);
nand U18587 (N_18587,N_18325,N_18217);
nand U18588 (N_18588,N_18382,N_18200);
xor U18589 (N_18589,N_18230,N_18348);
and U18590 (N_18590,N_18385,N_18292);
nor U18591 (N_18591,N_18345,N_18318);
xnor U18592 (N_18592,N_18330,N_18314);
nor U18593 (N_18593,N_18242,N_18220);
nand U18594 (N_18594,N_18287,N_18394);
xnor U18595 (N_18595,N_18273,N_18377);
and U18596 (N_18596,N_18327,N_18240);
or U18597 (N_18597,N_18290,N_18302);
or U18598 (N_18598,N_18356,N_18216);
nor U18599 (N_18599,N_18220,N_18341);
or U18600 (N_18600,N_18503,N_18546);
xnor U18601 (N_18601,N_18463,N_18530);
nor U18602 (N_18602,N_18455,N_18457);
and U18603 (N_18603,N_18476,N_18465);
and U18604 (N_18604,N_18513,N_18494);
nor U18605 (N_18605,N_18512,N_18484);
xnor U18606 (N_18606,N_18539,N_18496);
xor U18607 (N_18607,N_18436,N_18551);
and U18608 (N_18608,N_18557,N_18485);
or U18609 (N_18609,N_18556,N_18590);
and U18610 (N_18610,N_18450,N_18427);
and U18611 (N_18611,N_18423,N_18550);
xnor U18612 (N_18612,N_18477,N_18458);
and U18613 (N_18613,N_18489,N_18569);
and U18614 (N_18614,N_18573,N_18502);
nor U18615 (N_18615,N_18438,N_18425);
or U18616 (N_18616,N_18483,N_18522);
and U18617 (N_18617,N_18412,N_18426);
and U18618 (N_18618,N_18461,N_18584);
and U18619 (N_18619,N_18456,N_18531);
nor U18620 (N_18620,N_18408,N_18442);
and U18621 (N_18621,N_18469,N_18521);
or U18622 (N_18622,N_18549,N_18444);
nand U18623 (N_18623,N_18419,N_18571);
xnor U18624 (N_18624,N_18529,N_18534);
or U18625 (N_18625,N_18588,N_18559);
nor U18626 (N_18626,N_18555,N_18533);
nand U18627 (N_18627,N_18525,N_18500);
nand U18628 (N_18628,N_18583,N_18479);
or U18629 (N_18629,N_18422,N_18424);
or U18630 (N_18630,N_18597,N_18413);
nand U18631 (N_18631,N_18577,N_18486);
nor U18632 (N_18632,N_18474,N_18405);
xnor U18633 (N_18633,N_18542,N_18586);
and U18634 (N_18634,N_18574,N_18429);
nor U18635 (N_18635,N_18575,N_18493);
nor U18636 (N_18636,N_18468,N_18585);
nand U18637 (N_18637,N_18414,N_18596);
nand U18638 (N_18638,N_18526,N_18464);
and U18639 (N_18639,N_18421,N_18454);
or U18640 (N_18640,N_18443,N_18440);
nand U18641 (N_18641,N_18417,N_18580);
and U18642 (N_18642,N_18451,N_18568);
nor U18643 (N_18643,N_18431,N_18448);
or U18644 (N_18644,N_18558,N_18501);
nand U18645 (N_18645,N_18487,N_18506);
and U18646 (N_18646,N_18466,N_18581);
nor U18647 (N_18647,N_18570,N_18401);
nand U18648 (N_18648,N_18517,N_18540);
or U18649 (N_18649,N_18488,N_18491);
nand U18650 (N_18650,N_18579,N_18473);
nor U18651 (N_18651,N_18562,N_18402);
nand U18652 (N_18652,N_18428,N_18508);
xnor U18653 (N_18653,N_18409,N_18434);
nor U18654 (N_18654,N_18563,N_18439);
xor U18655 (N_18655,N_18591,N_18537);
nor U18656 (N_18656,N_18576,N_18518);
nor U18657 (N_18657,N_18509,N_18564);
nand U18658 (N_18658,N_18411,N_18516);
nand U18659 (N_18659,N_18482,N_18433);
nor U18660 (N_18660,N_18460,N_18447);
and U18661 (N_18661,N_18524,N_18453);
nand U18662 (N_18662,N_18527,N_18470);
nor U18663 (N_18663,N_18554,N_18415);
or U18664 (N_18664,N_18553,N_18481);
nor U18665 (N_18665,N_18407,N_18599);
nand U18666 (N_18666,N_18592,N_18535);
or U18667 (N_18667,N_18572,N_18510);
nand U18668 (N_18668,N_18441,N_18548);
xor U18669 (N_18669,N_18449,N_18404);
nand U18670 (N_18670,N_18547,N_18514);
and U18671 (N_18671,N_18490,N_18536);
nor U18672 (N_18672,N_18594,N_18567);
nor U18673 (N_18673,N_18587,N_18459);
nor U18674 (N_18674,N_18532,N_18515);
and U18675 (N_18675,N_18452,N_18437);
nor U18676 (N_18676,N_18418,N_18430);
nor U18677 (N_18677,N_18462,N_18561);
nand U18678 (N_18678,N_18560,N_18435);
nand U18679 (N_18679,N_18480,N_18504);
and U18680 (N_18680,N_18520,N_18519);
or U18681 (N_18681,N_18472,N_18400);
and U18682 (N_18682,N_18507,N_18499);
or U18683 (N_18683,N_18445,N_18432);
or U18684 (N_18684,N_18495,N_18416);
and U18685 (N_18685,N_18410,N_18471);
or U18686 (N_18686,N_18492,N_18505);
nand U18687 (N_18687,N_18543,N_18523);
and U18688 (N_18688,N_18589,N_18497);
xor U18689 (N_18689,N_18478,N_18406);
nor U18690 (N_18690,N_18511,N_18552);
or U18691 (N_18691,N_18578,N_18565);
xor U18692 (N_18692,N_18593,N_18420);
or U18693 (N_18693,N_18566,N_18541);
nor U18694 (N_18694,N_18538,N_18544);
xnor U18695 (N_18695,N_18598,N_18582);
nand U18696 (N_18696,N_18403,N_18528);
nor U18697 (N_18697,N_18595,N_18545);
or U18698 (N_18698,N_18498,N_18467);
or U18699 (N_18699,N_18446,N_18475);
nor U18700 (N_18700,N_18472,N_18575);
or U18701 (N_18701,N_18480,N_18472);
nor U18702 (N_18702,N_18437,N_18476);
nor U18703 (N_18703,N_18489,N_18514);
xnor U18704 (N_18704,N_18427,N_18558);
and U18705 (N_18705,N_18565,N_18454);
xor U18706 (N_18706,N_18599,N_18437);
and U18707 (N_18707,N_18407,N_18592);
and U18708 (N_18708,N_18438,N_18452);
nor U18709 (N_18709,N_18476,N_18454);
xor U18710 (N_18710,N_18573,N_18496);
nor U18711 (N_18711,N_18598,N_18509);
nand U18712 (N_18712,N_18490,N_18574);
nor U18713 (N_18713,N_18510,N_18583);
nand U18714 (N_18714,N_18597,N_18506);
nor U18715 (N_18715,N_18578,N_18521);
nand U18716 (N_18716,N_18417,N_18590);
and U18717 (N_18717,N_18418,N_18577);
and U18718 (N_18718,N_18417,N_18490);
nand U18719 (N_18719,N_18505,N_18599);
and U18720 (N_18720,N_18555,N_18445);
xnor U18721 (N_18721,N_18420,N_18520);
xnor U18722 (N_18722,N_18564,N_18512);
nor U18723 (N_18723,N_18546,N_18471);
and U18724 (N_18724,N_18593,N_18590);
nor U18725 (N_18725,N_18481,N_18508);
nand U18726 (N_18726,N_18533,N_18406);
xor U18727 (N_18727,N_18430,N_18454);
and U18728 (N_18728,N_18586,N_18490);
nand U18729 (N_18729,N_18464,N_18548);
nor U18730 (N_18730,N_18525,N_18476);
or U18731 (N_18731,N_18425,N_18483);
xnor U18732 (N_18732,N_18523,N_18563);
nand U18733 (N_18733,N_18509,N_18449);
xor U18734 (N_18734,N_18517,N_18464);
or U18735 (N_18735,N_18580,N_18507);
nor U18736 (N_18736,N_18576,N_18402);
nand U18737 (N_18737,N_18535,N_18573);
or U18738 (N_18738,N_18499,N_18471);
xnor U18739 (N_18739,N_18449,N_18474);
nand U18740 (N_18740,N_18453,N_18446);
xnor U18741 (N_18741,N_18428,N_18427);
nand U18742 (N_18742,N_18538,N_18448);
xor U18743 (N_18743,N_18549,N_18597);
xor U18744 (N_18744,N_18527,N_18466);
or U18745 (N_18745,N_18468,N_18449);
nand U18746 (N_18746,N_18599,N_18532);
xnor U18747 (N_18747,N_18408,N_18598);
nand U18748 (N_18748,N_18459,N_18497);
xnor U18749 (N_18749,N_18464,N_18562);
nand U18750 (N_18750,N_18591,N_18406);
nand U18751 (N_18751,N_18423,N_18420);
nand U18752 (N_18752,N_18532,N_18578);
or U18753 (N_18753,N_18406,N_18596);
and U18754 (N_18754,N_18583,N_18402);
nor U18755 (N_18755,N_18429,N_18459);
xnor U18756 (N_18756,N_18418,N_18401);
or U18757 (N_18757,N_18538,N_18409);
nand U18758 (N_18758,N_18407,N_18466);
xor U18759 (N_18759,N_18536,N_18590);
nand U18760 (N_18760,N_18598,N_18422);
xor U18761 (N_18761,N_18409,N_18412);
and U18762 (N_18762,N_18417,N_18474);
or U18763 (N_18763,N_18415,N_18487);
xor U18764 (N_18764,N_18414,N_18589);
nand U18765 (N_18765,N_18493,N_18419);
or U18766 (N_18766,N_18567,N_18453);
or U18767 (N_18767,N_18513,N_18589);
or U18768 (N_18768,N_18456,N_18492);
nor U18769 (N_18769,N_18558,N_18458);
nor U18770 (N_18770,N_18491,N_18556);
or U18771 (N_18771,N_18485,N_18434);
or U18772 (N_18772,N_18467,N_18536);
nor U18773 (N_18773,N_18582,N_18451);
nand U18774 (N_18774,N_18417,N_18597);
and U18775 (N_18775,N_18502,N_18454);
or U18776 (N_18776,N_18544,N_18536);
nor U18777 (N_18777,N_18499,N_18575);
xnor U18778 (N_18778,N_18484,N_18431);
or U18779 (N_18779,N_18415,N_18525);
and U18780 (N_18780,N_18580,N_18429);
and U18781 (N_18781,N_18440,N_18559);
nor U18782 (N_18782,N_18533,N_18519);
nand U18783 (N_18783,N_18475,N_18560);
nand U18784 (N_18784,N_18493,N_18461);
nor U18785 (N_18785,N_18462,N_18507);
nor U18786 (N_18786,N_18596,N_18445);
and U18787 (N_18787,N_18597,N_18496);
xnor U18788 (N_18788,N_18419,N_18579);
nor U18789 (N_18789,N_18551,N_18418);
nor U18790 (N_18790,N_18587,N_18547);
xnor U18791 (N_18791,N_18409,N_18478);
nor U18792 (N_18792,N_18417,N_18483);
and U18793 (N_18793,N_18461,N_18400);
or U18794 (N_18794,N_18445,N_18599);
or U18795 (N_18795,N_18567,N_18413);
nand U18796 (N_18796,N_18484,N_18549);
nand U18797 (N_18797,N_18525,N_18510);
nor U18798 (N_18798,N_18505,N_18591);
xor U18799 (N_18799,N_18584,N_18435);
nor U18800 (N_18800,N_18679,N_18697);
nand U18801 (N_18801,N_18618,N_18779);
and U18802 (N_18802,N_18756,N_18704);
xnor U18803 (N_18803,N_18726,N_18735);
nor U18804 (N_18804,N_18622,N_18693);
nand U18805 (N_18805,N_18714,N_18736);
nor U18806 (N_18806,N_18738,N_18600);
or U18807 (N_18807,N_18629,N_18750);
xor U18808 (N_18808,N_18631,N_18712);
nor U18809 (N_18809,N_18776,N_18604);
and U18810 (N_18810,N_18690,N_18689);
nor U18811 (N_18811,N_18683,N_18728);
xnor U18812 (N_18812,N_18734,N_18682);
or U18813 (N_18813,N_18639,N_18731);
or U18814 (N_18814,N_18782,N_18638);
or U18815 (N_18815,N_18640,N_18651);
xor U18816 (N_18816,N_18632,N_18793);
and U18817 (N_18817,N_18785,N_18650);
or U18818 (N_18818,N_18743,N_18769);
xor U18819 (N_18819,N_18752,N_18602);
xor U18820 (N_18820,N_18794,N_18724);
xnor U18821 (N_18821,N_18771,N_18661);
and U18822 (N_18822,N_18788,N_18627);
or U18823 (N_18823,N_18775,N_18706);
and U18824 (N_18824,N_18646,N_18616);
nand U18825 (N_18825,N_18680,N_18666);
xnor U18826 (N_18826,N_18740,N_18745);
nor U18827 (N_18827,N_18777,N_18623);
or U18828 (N_18828,N_18614,N_18705);
and U18829 (N_18829,N_18720,N_18737);
and U18830 (N_18830,N_18677,N_18798);
nor U18831 (N_18831,N_18762,N_18607);
nor U18832 (N_18832,N_18628,N_18685);
xor U18833 (N_18833,N_18643,N_18727);
or U18834 (N_18834,N_18605,N_18630);
nor U18835 (N_18835,N_18606,N_18626);
nand U18836 (N_18836,N_18636,N_18708);
nor U18837 (N_18837,N_18796,N_18687);
nor U18838 (N_18838,N_18755,N_18778);
or U18839 (N_18839,N_18676,N_18768);
or U18840 (N_18840,N_18733,N_18665);
or U18841 (N_18841,N_18730,N_18701);
nor U18842 (N_18842,N_18718,N_18688);
nor U18843 (N_18843,N_18649,N_18721);
nand U18844 (N_18844,N_18773,N_18786);
xor U18845 (N_18845,N_18692,N_18635);
nor U18846 (N_18846,N_18664,N_18767);
nand U18847 (N_18847,N_18648,N_18633);
nor U18848 (N_18848,N_18619,N_18671);
and U18849 (N_18849,N_18765,N_18624);
nor U18850 (N_18850,N_18699,N_18610);
nor U18851 (N_18851,N_18723,N_18662);
and U18852 (N_18852,N_18797,N_18757);
nor U18853 (N_18853,N_18764,N_18642);
or U18854 (N_18854,N_18657,N_18789);
or U18855 (N_18855,N_18625,N_18783);
nand U18856 (N_18856,N_18791,N_18641);
xor U18857 (N_18857,N_18603,N_18725);
nand U18858 (N_18858,N_18644,N_18751);
nor U18859 (N_18859,N_18670,N_18790);
or U18860 (N_18860,N_18621,N_18686);
or U18861 (N_18861,N_18795,N_18715);
nand U18862 (N_18862,N_18758,N_18684);
and U18863 (N_18863,N_18647,N_18601);
or U18864 (N_18864,N_18645,N_18617);
xnor U18865 (N_18865,N_18674,N_18620);
xor U18866 (N_18866,N_18754,N_18700);
xor U18867 (N_18867,N_18709,N_18652);
or U18868 (N_18868,N_18763,N_18669);
xnor U18869 (N_18869,N_18656,N_18612);
and U18870 (N_18870,N_18702,N_18717);
nand U18871 (N_18871,N_18710,N_18781);
and U18872 (N_18872,N_18694,N_18654);
xnor U18873 (N_18873,N_18707,N_18716);
nand U18874 (N_18874,N_18766,N_18659);
nand U18875 (N_18875,N_18739,N_18637);
xnor U18876 (N_18876,N_18784,N_18655);
xor U18877 (N_18877,N_18753,N_18770);
and U18878 (N_18878,N_18634,N_18678);
xnor U18879 (N_18879,N_18703,N_18759);
and U18880 (N_18880,N_18729,N_18713);
or U18881 (N_18881,N_18742,N_18660);
and U18882 (N_18882,N_18749,N_18787);
or U18883 (N_18883,N_18780,N_18760);
nand U18884 (N_18884,N_18608,N_18711);
nor U18885 (N_18885,N_18772,N_18744);
or U18886 (N_18886,N_18696,N_18681);
and U18887 (N_18887,N_18746,N_18747);
nand U18888 (N_18888,N_18722,N_18774);
or U18889 (N_18889,N_18611,N_18792);
nand U18890 (N_18890,N_18667,N_18663);
xor U18891 (N_18891,N_18658,N_18799);
nand U18892 (N_18892,N_18761,N_18695);
nand U18893 (N_18893,N_18609,N_18719);
nor U18894 (N_18894,N_18613,N_18673);
nor U18895 (N_18895,N_18732,N_18615);
and U18896 (N_18896,N_18691,N_18672);
nand U18897 (N_18897,N_18741,N_18653);
nand U18898 (N_18898,N_18675,N_18668);
nor U18899 (N_18899,N_18748,N_18698);
nand U18900 (N_18900,N_18639,N_18680);
xnor U18901 (N_18901,N_18637,N_18609);
and U18902 (N_18902,N_18708,N_18639);
or U18903 (N_18903,N_18666,N_18677);
or U18904 (N_18904,N_18669,N_18650);
nand U18905 (N_18905,N_18649,N_18773);
nand U18906 (N_18906,N_18702,N_18623);
or U18907 (N_18907,N_18767,N_18618);
xor U18908 (N_18908,N_18725,N_18640);
xor U18909 (N_18909,N_18682,N_18726);
nor U18910 (N_18910,N_18727,N_18763);
nand U18911 (N_18911,N_18668,N_18644);
nand U18912 (N_18912,N_18676,N_18698);
nor U18913 (N_18913,N_18743,N_18780);
or U18914 (N_18914,N_18650,N_18666);
nor U18915 (N_18915,N_18686,N_18709);
xor U18916 (N_18916,N_18747,N_18710);
or U18917 (N_18917,N_18696,N_18687);
xnor U18918 (N_18918,N_18683,N_18658);
or U18919 (N_18919,N_18676,N_18695);
nand U18920 (N_18920,N_18642,N_18716);
and U18921 (N_18921,N_18727,N_18612);
and U18922 (N_18922,N_18641,N_18718);
nand U18923 (N_18923,N_18797,N_18702);
or U18924 (N_18924,N_18723,N_18714);
and U18925 (N_18925,N_18770,N_18660);
or U18926 (N_18926,N_18690,N_18682);
xnor U18927 (N_18927,N_18778,N_18789);
and U18928 (N_18928,N_18673,N_18651);
and U18929 (N_18929,N_18644,N_18739);
and U18930 (N_18930,N_18752,N_18739);
and U18931 (N_18931,N_18658,N_18754);
or U18932 (N_18932,N_18606,N_18666);
and U18933 (N_18933,N_18747,N_18675);
xnor U18934 (N_18934,N_18731,N_18727);
or U18935 (N_18935,N_18674,N_18657);
or U18936 (N_18936,N_18737,N_18726);
xnor U18937 (N_18937,N_18636,N_18769);
or U18938 (N_18938,N_18785,N_18748);
or U18939 (N_18939,N_18669,N_18603);
nor U18940 (N_18940,N_18794,N_18730);
nor U18941 (N_18941,N_18707,N_18772);
or U18942 (N_18942,N_18669,N_18612);
xor U18943 (N_18943,N_18727,N_18732);
or U18944 (N_18944,N_18753,N_18796);
nor U18945 (N_18945,N_18628,N_18776);
and U18946 (N_18946,N_18629,N_18796);
or U18947 (N_18947,N_18650,N_18688);
and U18948 (N_18948,N_18671,N_18736);
or U18949 (N_18949,N_18770,N_18625);
nor U18950 (N_18950,N_18600,N_18724);
nand U18951 (N_18951,N_18722,N_18793);
xnor U18952 (N_18952,N_18673,N_18749);
or U18953 (N_18953,N_18766,N_18697);
and U18954 (N_18954,N_18690,N_18647);
xor U18955 (N_18955,N_18678,N_18779);
nand U18956 (N_18956,N_18736,N_18696);
or U18957 (N_18957,N_18627,N_18734);
nand U18958 (N_18958,N_18665,N_18717);
and U18959 (N_18959,N_18719,N_18755);
or U18960 (N_18960,N_18634,N_18768);
nand U18961 (N_18961,N_18672,N_18711);
nor U18962 (N_18962,N_18700,N_18751);
xnor U18963 (N_18963,N_18656,N_18789);
and U18964 (N_18964,N_18690,N_18703);
or U18965 (N_18965,N_18742,N_18736);
and U18966 (N_18966,N_18692,N_18731);
nor U18967 (N_18967,N_18716,N_18784);
nand U18968 (N_18968,N_18666,N_18794);
and U18969 (N_18969,N_18769,N_18651);
nand U18970 (N_18970,N_18670,N_18607);
and U18971 (N_18971,N_18762,N_18679);
xnor U18972 (N_18972,N_18623,N_18703);
and U18973 (N_18973,N_18642,N_18748);
nor U18974 (N_18974,N_18671,N_18700);
nor U18975 (N_18975,N_18798,N_18758);
nand U18976 (N_18976,N_18782,N_18675);
nor U18977 (N_18977,N_18610,N_18713);
nor U18978 (N_18978,N_18781,N_18613);
nand U18979 (N_18979,N_18709,N_18703);
or U18980 (N_18980,N_18698,N_18732);
nor U18981 (N_18981,N_18711,N_18643);
or U18982 (N_18982,N_18797,N_18762);
and U18983 (N_18983,N_18601,N_18752);
nand U18984 (N_18984,N_18626,N_18629);
or U18985 (N_18985,N_18700,N_18740);
or U18986 (N_18986,N_18659,N_18721);
nor U18987 (N_18987,N_18712,N_18761);
and U18988 (N_18988,N_18702,N_18644);
nor U18989 (N_18989,N_18741,N_18718);
nand U18990 (N_18990,N_18668,N_18603);
nand U18991 (N_18991,N_18782,N_18645);
nand U18992 (N_18992,N_18766,N_18791);
nand U18993 (N_18993,N_18753,N_18692);
nor U18994 (N_18994,N_18662,N_18719);
or U18995 (N_18995,N_18602,N_18627);
nor U18996 (N_18996,N_18629,N_18650);
and U18997 (N_18997,N_18785,N_18770);
nor U18998 (N_18998,N_18725,N_18641);
nor U18999 (N_18999,N_18763,N_18660);
or U19000 (N_19000,N_18884,N_18908);
or U19001 (N_19001,N_18922,N_18904);
and U19002 (N_19002,N_18949,N_18984);
xnor U19003 (N_19003,N_18835,N_18851);
and U19004 (N_19004,N_18878,N_18981);
and U19005 (N_19005,N_18823,N_18850);
xnor U19006 (N_19006,N_18986,N_18971);
or U19007 (N_19007,N_18910,N_18913);
nor U19008 (N_19008,N_18834,N_18839);
and U19009 (N_19009,N_18988,N_18818);
nor U19010 (N_19010,N_18927,N_18975);
or U19011 (N_19011,N_18974,N_18942);
or U19012 (N_19012,N_18808,N_18865);
and U19013 (N_19013,N_18929,N_18995);
xor U19014 (N_19014,N_18862,N_18859);
xnor U19015 (N_19015,N_18821,N_18939);
nand U19016 (N_19016,N_18882,N_18963);
xor U19017 (N_19017,N_18985,N_18833);
xor U19018 (N_19018,N_18830,N_18936);
xnor U19019 (N_19019,N_18940,N_18982);
nor U19020 (N_19020,N_18806,N_18919);
nand U19021 (N_19021,N_18816,N_18979);
nor U19022 (N_19022,N_18809,N_18888);
xnor U19023 (N_19023,N_18915,N_18832);
xor U19024 (N_19024,N_18872,N_18935);
nand U19025 (N_19025,N_18905,N_18914);
nand U19026 (N_19026,N_18909,N_18967);
xor U19027 (N_19027,N_18814,N_18869);
nor U19028 (N_19028,N_18920,N_18932);
nand U19029 (N_19029,N_18838,N_18893);
or U19030 (N_19030,N_18897,N_18828);
nor U19031 (N_19031,N_18894,N_18848);
and U19032 (N_19032,N_18877,N_18976);
or U19033 (N_19033,N_18863,N_18885);
nand U19034 (N_19034,N_18958,N_18966);
xor U19035 (N_19035,N_18965,N_18956);
nand U19036 (N_19036,N_18868,N_18951);
and U19037 (N_19037,N_18934,N_18998);
or U19038 (N_19038,N_18997,N_18871);
and U19039 (N_19039,N_18824,N_18944);
nand U19040 (N_19040,N_18961,N_18802);
and U19041 (N_19041,N_18970,N_18836);
nand U19042 (N_19042,N_18968,N_18898);
nor U19043 (N_19043,N_18918,N_18805);
and U19044 (N_19044,N_18917,N_18937);
nor U19045 (N_19045,N_18957,N_18827);
and U19046 (N_19046,N_18887,N_18807);
xor U19047 (N_19047,N_18943,N_18916);
or U19048 (N_19048,N_18858,N_18879);
nand U19049 (N_19049,N_18962,N_18912);
and U19050 (N_19050,N_18901,N_18954);
and U19051 (N_19051,N_18886,N_18825);
or U19052 (N_19052,N_18964,N_18837);
nand U19053 (N_19053,N_18911,N_18946);
nand U19054 (N_19054,N_18803,N_18953);
xnor U19055 (N_19055,N_18867,N_18813);
nor U19056 (N_19056,N_18969,N_18841);
or U19057 (N_19057,N_18804,N_18800);
and U19058 (N_19058,N_18955,N_18812);
nor U19059 (N_19059,N_18810,N_18931);
xnor U19060 (N_19060,N_18928,N_18892);
or U19061 (N_19061,N_18801,N_18923);
or U19062 (N_19062,N_18989,N_18817);
nor U19063 (N_19063,N_18852,N_18960);
or U19064 (N_19064,N_18847,N_18891);
nor U19065 (N_19065,N_18948,N_18857);
xor U19066 (N_19066,N_18843,N_18972);
and U19067 (N_19067,N_18993,N_18903);
or U19068 (N_19068,N_18980,N_18831);
nor U19069 (N_19069,N_18926,N_18846);
xor U19070 (N_19070,N_18866,N_18820);
or U19071 (N_19071,N_18811,N_18959);
and U19072 (N_19072,N_18895,N_18856);
nor U19073 (N_19073,N_18815,N_18881);
or U19074 (N_19074,N_18822,N_18996);
nor U19075 (N_19075,N_18977,N_18941);
and U19076 (N_19076,N_18978,N_18842);
xnor U19077 (N_19077,N_18991,N_18876);
and U19078 (N_19078,N_18870,N_18861);
and U19079 (N_19079,N_18947,N_18952);
xnor U19080 (N_19080,N_18875,N_18994);
nor U19081 (N_19081,N_18990,N_18845);
or U19082 (N_19082,N_18983,N_18921);
nor U19083 (N_19083,N_18819,N_18829);
and U19084 (N_19084,N_18860,N_18844);
xnor U19085 (N_19085,N_18945,N_18999);
nand U19086 (N_19086,N_18855,N_18854);
and U19087 (N_19087,N_18930,N_18873);
nand U19088 (N_19088,N_18883,N_18973);
nand U19089 (N_19089,N_18899,N_18849);
and U19090 (N_19090,N_18938,N_18933);
nor U19091 (N_19091,N_18896,N_18889);
or U19092 (N_19092,N_18924,N_18853);
or U19093 (N_19093,N_18826,N_18992);
nor U19094 (N_19094,N_18890,N_18864);
or U19095 (N_19095,N_18987,N_18902);
nor U19096 (N_19096,N_18900,N_18907);
xnor U19097 (N_19097,N_18950,N_18840);
or U19098 (N_19098,N_18925,N_18874);
and U19099 (N_19099,N_18906,N_18880);
xor U19100 (N_19100,N_18868,N_18977);
nor U19101 (N_19101,N_18909,N_18872);
and U19102 (N_19102,N_18958,N_18977);
and U19103 (N_19103,N_18806,N_18888);
or U19104 (N_19104,N_18828,N_18970);
and U19105 (N_19105,N_18890,N_18850);
and U19106 (N_19106,N_18816,N_18881);
xor U19107 (N_19107,N_18927,N_18850);
and U19108 (N_19108,N_18837,N_18889);
nor U19109 (N_19109,N_18909,N_18987);
or U19110 (N_19110,N_18953,N_18883);
nand U19111 (N_19111,N_18925,N_18960);
or U19112 (N_19112,N_18995,N_18951);
nand U19113 (N_19113,N_18941,N_18805);
nand U19114 (N_19114,N_18992,N_18978);
xor U19115 (N_19115,N_18806,N_18973);
nor U19116 (N_19116,N_18801,N_18999);
xnor U19117 (N_19117,N_18946,N_18846);
nor U19118 (N_19118,N_18872,N_18895);
xnor U19119 (N_19119,N_18987,N_18849);
nand U19120 (N_19120,N_18977,N_18900);
nor U19121 (N_19121,N_18823,N_18872);
xor U19122 (N_19122,N_18972,N_18999);
nor U19123 (N_19123,N_18928,N_18845);
nand U19124 (N_19124,N_18857,N_18963);
nand U19125 (N_19125,N_18803,N_18905);
xnor U19126 (N_19126,N_18830,N_18975);
nor U19127 (N_19127,N_18960,N_18856);
and U19128 (N_19128,N_18812,N_18921);
or U19129 (N_19129,N_18809,N_18967);
or U19130 (N_19130,N_18863,N_18994);
nor U19131 (N_19131,N_18953,N_18860);
or U19132 (N_19132,N_18893,N_18989);
or U19133 (N_19133,N_18973,N_18868);
nand U19134 (N_19134,N_18996,N_18842);
nor U19135 (N_19135,N_18846,N_18804);
nor U19136 (N_19136,N_18998,N_18848);
nor U19137 (N_19137,N_18921,N_18863);
or U19138 (N_19138,N_18829,N_18883);
xor U19139 (N_19139,N_18838,N_18846);
nor U19140 (N_19140,N_18914,N_18874);
xnor U19141 (N_19141,N_18919,N_18826);
nor U19142 (N_19142,N_18983,N_18809);
nor U19143 (N_19143,N_18900,N_18945);
or U19144 (N_19144,N_18977,N_18949);
or U19145 (N_19145,N_18956,N_18902);
and U19146 (N_19146,N_18932,N_18965);
xor U19147 (N_19147,N_18985,N_18945);
or U19148 (N_19148,N_18824,N_18886);
xor U19149 (N_19149,N_18978,N_18813);
nand U19150 (N_19150,N_18945,N_18855);
nand U19151 (N_19151,N_18811,N_18819);
xor U19152 (N_19152,N_18970,N_18984);
or U19153 (N_19153,N_18806,N_18921);
nor U19154 (N_19154,N_18846,N_18825);
or U19155 (N_19155,N_18836,N_18877);
xor U19156 (N_19156,N_18868,N_18825);
nand U19157 (N_19157,N_18957,N_18872);
nor U19158 (N_19158,N_18986,N_18927);
xnor U19159 (N_19159,N_18830,N_18875);
and U19160 (N_19160,N_18892,N_18979);
or U19161 (N_19161,N_18928,N_18975);
or U19162 (N_19162,N_18941,N_18898);
nand U19163 (N_19163,N_18954,N_18986);
and U19164 (N_19164,N_18943,N_18833);
xor U19165 (N_19165,N_18965,N_18833);
nand U19166 (N_19166,N_18955,N_18945);
or U19167 (N_19167,N_18891,N_18883);
xor U19168 (N_19168,N_18888,N_18887);
nor U19169 (N_19169,N_18852,N_18975);
or U19170 (N_19170,N_18950,N_18832);
nor U19171 (N_19171,N_18984,N_18922);
nand U19172 (N_19172,N_18989,N_18887);
and U19173 (N_19173,N_18873,N_18911);
xnor U19174 (N_19174,N_18898,N_18962);
nor U19175 (N_19175,N_18979,N_18985);
nand U19176 (N_19176,N_18865,N_18902);
nor U19177 (N_19177,N_18968,N_18805);
and U19178 (N_19178,N_18991,N_18920);
or U19179 (N_19179,N_18805,N_18824);
nor U19180 (N_19180,N_18907,N_18985);
xnor U19181 (N_19181,N_18964,N_18881);
nor U19182 (N_19182,N_18890,N_18976);
nor U19183 (N_19183,N_18830,N_18977);
nand U19184 (N_19184,N_18870,N_18904);
and U19185 (N_19185,N_18836,N_18928);
or U19186 (N_19186,N_18991,N_18965);
and U19187 (N_19187,N_18988,N_18810);
or U19188 (N_19188,N_18844,N_18826);
or U19189 (N_19189,N_18952,N_18981);
or U19190 (N_19190,N_18944,N_18822);
xor U19191 (N_19191,N_18853,N_18912);
or U19192 (N_19192,N_18806,N_18829);
nor U19193 (N_19193,N_18934,N_18953);
and U19194 (N_19194,N_18845,N_18970);
nand U19195 (N_19195,N_18872,N_18900);
or U19196 (N_19196,N_18922,N_18932);
xnor U19197 (N_19197,N_18814,N_18846);
or U19198 (N_19198,N_18805,N_18914);
nand U19199 (N_19199,N_18980,N_18899);
nand U19200 (N_19200,N_19078,N_19151);
nand U19201 (N_19201,N_19158,N_19000);
and U19202 (N_19202,N_19090,N_19176);
and U19203 (N_19203,N_19142,N_19192);
and U19204 (N_19204,N_19047,N_19022);
nand U19205 (N_19205,N_19074,N_19025);
nor U19206 (N_19206,N_19164,N_19171);
and U19207 (N_19207,N_19070,N_19177);
xnor U19208 (N_19208,N_19133,N_19028);
nor U19209 (N_19209,N_19137,N_19053);
and U19210 (N_19210,N_19087,N_19084);
nand U19211 (N_19211,N_19049,N_19165);
or U19212 (N_19212,N_19135,N_19129);
and U19213 (N_19213,N_19170,N_19037);
nor U19214 (N_19214,N_19172,N_19120);
xor U19215 (N_19215,N_19175,N_19033);
and U19216 (N_19216,N_19122,N_19190);
nand U19217 (N_19217,N_19044,N_19174);
xor U19218 (N_19218,N_19160,N_19054);
or U19219 (N_19219,N_19157,N_19008);
and U19220 (N_19220,N_19071,N_19094);
nand U19221 (N_19221,N_19099,N_19132);
xnor U19222 (N_19222,N_19154,N_19155);
nor U19223 (N_19223,N_19046,N_19145);
nand U19224 (N_19224,N_19061,N_19167);
nor U19225 (N_19225,N_19002,N_19141);
and U19226 (N_19226,N_19178,N_19086);
or U19227 (N_19227,N_19100,N_19196);
or U19228 (N_19228,N_19005,N_19199);
nand U19229 (N_19229,N_19184,N_19095);
xnor U19230 (N_19230,N_19194,N_19089);
or U19231 (N_19231,N_19088,N_19106);
or U19232 (N_19232,N_19015,N_19065);
and U19233 (N_19233,N_19161,N_19169);
nor U19234 (N_19234,N_19032,N_19007);
and U19235 (N_19235,N_19064,N_19105);
and U19236 (N_19236,N_19055,N_19068);
and U19237 (N_19237,N_19188,N_19117);
nor U19238 (N_19238,N_19042,N_19051);
nor U19239 (N_19239,N_19052,N_19163);
nor U19240 (N_19240,N_19104,N_19183);
nand U19241 (N_19241,N_19026,N_19111);
or U19242 (N_19242,N_19024,N_19128);
nand U19243 (N_19243,N_19112,N_19050);
nand U19244 (N_19244,N_19031,N_19080);
or U19245 (N_19245,N_19118,N_19072);
xor U19246 (N_19246,N_19166,N_19168);
nor U19247 (N_19247,N_19082,N_19077);
or U19248 (N_19248,N_19043,N_19110);
nand U19249 (N_19249,N_19010,N_19138);
or U19250 (N_19250,N_19126,N_19108);
and U19251 (N_19251,N_19181,N_19143);
xor U19252 (N_19252,N_19107,N_19123);
and U19253 (N_19253,N_19017,N_19013);
or U19254 (N_19254,N_19030,N_19062);
and U19255 (N_19255,N_19144,N_19149);
xnor U19256 (N_19256,N_19009,N_19011);
or U19257 (N_19257,N_19125,N_19085);
xnor U19258 (N_19258,N_19036,N_19131);
xor U19259 (N_19259,N_19197,N_19034);
and U19260 (N_19260,N_19029,N_19198);
nand U19261 (N_19261,N_19060,N_19140);
and U19262 (N_19262,N_19098,N_19038);
xor U19263 (N_19263,N_19021,N_19162);
xnor U19264 (N_19264,N_19114,N_19136);
xnor U19265 (N_19265,N_19040,N_19187);
nor U19266 (N_19266,N_19076,N_19102);
nand U19267 (N_19267,N_19004,N_19139);
and U19268 (N_19268,N_19073,N_19093);
xor U19269 (N_19269,N_19014,N_19016);
nor U19270 (N_19270,N_19191,N_19091);
or U19271 (N_19271,N_19182,N_19159);
and U19272 (N_19272,N_19067,N_19103);
or U19273 (N_19273,N_19124,N_19109);
xor U19274 (N_19274,N_19039,N_19035);
nand U19275 (N_19275,N_19127,N_19018);
xor U19276 (N_19276,N_19130,N_19186);
or U19277 (N_19277,N_19134,N_19048);
xnor U19278 (N_19278,N_19179,N_19113);
and U19279 (N_19279,N_19069,N_19189);
or U19280 (N_19280,N_19023,N_19075);
or U19281 (N_19281,N_19045,N_19146);
or U19282 (N_19282,N_19101,N_19092);
nand U19283 (N_19283,N_19059,N_19153);
xnor U19284 (N_19284,N_19147,N_19116);
nor U19285 (N_19285,N_19019,N_19003);
xor U19286 (N_19286,N_19058,N_19012);
and U19287 (N_19287,N_19041,N_19195);
and U19288 (N_19288,N_19150,N_19057);
xor U19289 (N_19289,N_19066,N_19056);
xor U19290 (N_19290,N_19027,N_19156);
xnor U19291 (N_19291,N_19193,N_19180);
or U19292 (N_19292,N_19063,N_19121);
xor U19293 (N_19293,N_19079,N_19083);
nor U19294 (N_19294,N_19001,N_19096);
xor U19295 (N_19295,N_19173,N_19119);
and U19296 (N_19296,N_19097,N_19185);
or U19297 (N_19297,N_19115,N_19152);
xor U19298 (N_19298,N_19020,N_19006);
or U19299 (N_19299,N_19148,N_19081);
nor U19300 (N_19300,N_19177,N_19001);
and U19301 (N_19301,N_19071,N_19067);
xnor U19302 (N_19302,N_19027,N_19043);
xnor U19303 (N_19303,N_19142,N_19014);
nor U19304 (N_19304,N_19090,N_19034);
nor U19305 (N_19305,N_19134,N_19156);
xnor U19306 (N_19306,N_19104,N_19047);
or U19307 (N_19307,N_19147,N_19027);
nand U19308 (N_19308,N_19152,N_19127);
and U19309 (N_19309,N_19161,N_19093);
and U19310 (N_19310,N_19069,N_19012);
nor U19311 (N_19311,N_19047,N_19074);
or U19312 (N_19312,N_19039,N_19012);
nor U19313 (N_19313,N_19006,N_19015);
xnor U19314 (N_19314,N_19028,N_19030);
and U19315 (N_19315,N_19199,N_19185);
or U19316 (N_19316,N_19170,N_19149);
or U19317 (N_19317,N_19023,N_19162);
and U19318 (N_19318,N_19080,N_19052);
and U19319 (N_19319,N_19076,N_19108);
xor U19320 (N_19320,N_19056,N_19021);
or U19321 (N_19321,N_19047,N_19146);
nand U19322 (N_19322,N_19184,N_19173);
nand U19323 (N_19323,N_19169,N_19005);
or U19324 (N_19324,N_19110,N_19151);
nand U19325 (N_19325,N_19080,N_19082);
or U19326 (N_19326,N_19041,N_19024);
nand U19327 (N_19327,N_19078,N_19153);
nor U19328 (N_19328,N_19138,N_19145);
or U19329 (N_19329,N_19169,N_19110);
nor U19330 (N_19330,N_19140,N_19112);
nor U19331 (N_19331,N_19102,N_19027);
nand U19332 (N_19332,N_19075,N_19162);
nand U19333 (N_19333,N_19074,N_19179);
and U19334 (N_19334,N_19064,N_19016);
and U19335 (N_19335,N_19185,N_19003);
xor U19336 (N_19336,N_19177,N_19074);
nor U19337 (N_19337,N_19148,N_19188);
xnor U19338 (N_19338,N_19181,N_19011);
or U19339 (N_19339,N_19003,N_19072);
nor U19340 (N_19340,N_19172,N_19134);
nor U19341 (N_19341,N_19100,N_19180);
or U19342 (N_19342,N_19096,N_19013);
nand U19343 (N_19343,N_19006,N_19132);
xor U19344 (N_19344,N_19149,N_19125);
xnor U19345 (N_19345,N_19162,N_19097);
xnor U19346 (N_19346,N_19112,N_19183);
nor U19347 (N_19347,N_19152,N_19079);
nand U19348 (N_19348,N_19070,N_19199);
nand U19349 (N_19349,N_19119,N_19010);
or U19350 (N_19350,N_19061,N_19103);
and U19351 (N_19351,N_19007,N_19042);
or U19352 (N_19352,N_19045,N_19011);
and U19353 (N_19353,N_19004,N_19089);
nand U19354 (N_19354,N_19192,N_19160);
nor U19355 (N_19355,N_19068,N_19034);
or U19356 (N_19356,N_19078,N_19177);
nand U19357 (N_19357,N_19079,N_19004);
or U19358 (N_19358,N_19025,N_19156);
xnor U19359 (N_19359,N_19170,N_19155);
and U19360 (N_19360,N_19161,N_19198);
and U19361 (N_19361,N_19080,N_19152);
and U19362 (N_19362,N_19137,N_19112);
xor U19363 (N_19363,N_19196,N_19148);
xnor U19364 (N_19364,N_19117,N_19178);
and U19365 (N_19365,N_19062,N_19122);
nand U19366 (N_19366,N_19108,N_19157);
or U19367 (N_19367,N_19123,N_19139);
or U19368 (N_19368,N_19066,N_19177);
xor U19369 (N_19369,N_19004,N_19164);
or U19370 (N_19370,N_19087,N_19174);
or U19371 (N_19371,N_19074,N_19135);
xor U19372 (N_19372,N_19128,N_19051);
xor U19373 (N_19373,N_19013,N_19050);
xor U19374 (N_19374,N_19110,N_19089);
nor U19375 (N_19375,N_19001,N_19154);
or U19376 (N_19376,N_19032,N_19100);
xnor U19377 (N_19377,N_19094,N_19189);
nor U19378 (N_19378,N_19118,N_19086);
nand U19379 (N_19379,N_19047,N_19045);
or U19380 (N_19380,N_19147,N_19002);
and U19381 (N_19381,N_19095,N_19156);
nor U19382 (N_19382,N_19060,N_19070);
nor U19383 (N_19383,N_19028,N_19123);
or U19384 (N_19384,N_19100,N_19016);
nor U19385 (N_19385,N_19079,N_19101);
nand U19386 (N_19386,N_19179,N_19147);
nor U19387 (N_19387,N_19086,N_19171);
nor U19388 (N_19388,N_19028,N_19085);
nand U19389 (N_19389,N_19176,N_19018);
nor U19390 (N_19390,N_19131,N_19016);
nor U19391 (N_19391,N_19089,N_19170);
xor U19392 (N_19392,N_19017,N_19035);
or U19393 (N_19393,N_19159,N_19041);
nand U19394 (N_19394,N_19169,N_19121);
or U19395 (N_19395,N_19134,N_19050);
and U19396 (N_19396,N_19042,N_19146);
or U19397 (N_19397,N_19093,N_19001);
xor U19398 (N_19398,N_19072,N_19162);
and U19399 (N_19399,N_19134,N_19133);
nor U19400 (N_19400,N_19376,N_19361);
or U19401 (N_19401,N_19340,N_19231);
xor U19402 (N_19402,N_19305,N_19389);
xnor U19403 (N_19403,N_19239,N_19354);
and U19404 (N_19404,N_19212,N_19281);
nor U19405 (N_19405,N_19312,N_19228);
or U19406 (N_19406,N_19217,N_19315);
and U19407 (N_19407,N_19328,N_19223);
or U19408 (N_19408,N_19370,N_19313);
and U19409 (N_19409,N_19381,N_19369);
or U19410 (N_19410,N_19353,N_19234);
nor U19411 (N_19411,N_19259,N_19248);
nand U19412 (N_19412,N_19200,N_19351);
or U19413 (N_19413,N_19268,N_19262);
nor U19414 (N_19414,N_19392,N_19277);
and U19415 (N_19415,N_19338,N_19350);
nand U19416 (N_19416,N_19393,N_19276);
nand U19417 (N_19417,N_19334,N_19273);
or U19418 (N_19418,N_19310,N_19347);
nor U19419 (N_19419,N_19318,N_19289);
or U19420 (N_19420,N_19294,N_19357);
and U19421 (N_19421,N_19220,N_19304);
and U19422 (N_19422,N_19321,N_19386);
and U19423 (N_19423,N_19319,N_19226);
nand U19424 (N_19424,N_19307,N_19385);
nor U19425 (N_19425,N_19271,N_19378);
or U19426 (N_19426,N_19325,N_19291);
nand U19427 (N_19427,N_19395,N_19383);
and U19428 (N_19428,N_19363,N_19208);
nand U19429 (N_19429,N_19394,N_19269);
or U19430 (N_19430,N_19348,N_19374);
and U19431 (N_19431,N_19205,N_19298);
and U19432 (N_19432,N_19341,N_19331);
xor U19433 (N_19433,N_19222,N_19266);
or U19434 (N_19434,N_19355,N_19290);
nor U19435 (N_19435,N_19240,N_19275);
nor U19436 (N_19436,N_19251,N_19286);
or U19437 (N_19437,N_19206,N_19218);
nand U19438 (N_19438,N_19336,N_19380);
or U19439 (N_19439,N_19301,N_19261);
nand U19440 (N_19440,N_19390,N_19322);
nor U19441 (N_19441,N_19326,N_19241);
nor U19442 (N_19442,N_19254,N_19372);
or U19443 (N_19443,N_19246,N_19335);
nand U19444 (N_19444,N_19202,N_19243);
xor U19445 (N_19445,N_19391,N_19309);
xnor U19446 (N_19446,N_19210,N_19256);
xnor U19447 (N_19447,N_19229,N_19329);
or U19448 (N_19448,N_19213,N_19365);
nor U19449 (N_19449,N_19300,N_19283);
nor U19450 (N_19450,N_19252,N_19352);
xnor U19451 (N_19451,N_19219,N_19373);
or U19452 (N_19452,N_19364,N_19270);
and U19453 (N_19453,N_19201,N_19356);
xnor U19454 (N_19454,N_19204,N_19302);
nand U19455 (N_19455,N_19387,N_19396);
or U19456 (N_19456,N_19267,N_19368);
nor U19457 (N_19457,N_19296,N_19238);
nand U19458 (N_19458,N_19257,N_19299);
nand U19459 (N_19459,N_19255,N_19343);
nor U19460 (N_19460,N_19211,N_19264);
nand U19461 (N_19461,N_19253,N_19303);
nand U19462 (N_19462,N_19282,N_19382);
nand U19463 (N_19463,N_19327,N_19245);
and U19464 (N_19464,N_19339,N_19379);
nand U19465 (N_19465,N_19371,N_19209);
and U19466 (N_19466,N_19332,N_19366);
and U19467 (N_19467,N_19388,N_19250);
and U19468 (N_19468,N_19280,N_19237);
nor U19469 (N_19469,N_19375,N_19362);
nor U19470 (N_19470,N_19384,N_19346);
nor U19471 (N_19471,N_19295,N_19244);
and U19472 (N_19472,N_19342,N_19288);
or U19473 (N_19473,N_19265,N_19214);
nand U19474 (N_19474,N_19263,N_19233);
xnor U19475 (N_19475,N_19278,N_19324);
or U19476 (N_19476,N_19258,N_19330);
xnor U19477 (N_19477,N_19225,N_19232);
nand U19478 (N_19478,N_19221,N_19317);
nand U19479 (N_19479,N_19249,N_19397);
nand U19480 (N_19480,N_19230,N_19399);
nand U19481 (N_19481,N_19297,N_19216);
xor U19482 (N_19482,N_19285,N_19287);
and U19483 (N_19483,N_19235,N_19323);
nor U19484 (N_19484,N_19242,N_19260);
or U19485 (N_19485,N_19308,N_19337);
xnor U19486 (N_19486,N_19284,N_19398);
or U19487 (N_19487,N_19247,N_19203);
nor U19488 (N_19488,N_19215,N_19316);
or U19489 (N_19489,N_19311,N_19227);
nand U19490 (N_19490,N_19359,N_19279);
nor U19491 (N_19491,N_19207,N_19236);
xnor U19492 (N_19492,N_19292,N_19274);
nor U19493 (N_19493,N_19344,N_19377);
and U19494 (N_19494,N_19333,N_19224);
xnor U19495 (N_19495,N_19349,N_19367);
nor U19496 (N_19496,N_19306,N_19272);
nor U19497 (N_19497,N_19360,N_19358);
and U19498 (N_19498,N_19320,N_19293);
nand U19499 (N_19499,N_19314,N_19345);
nor U19500 (N_19500,N_19270,N_19284);
or U19501 (N_19501,N_19372,N_19226);
or U19502 (N_19502,N_19366,N_19373);
nor U19503 (N_19503,N_19297,N_19256);
or U19504 (N_19504,N_19351,N_19326);
nand U19505 (N_19505,N_19206,N_19351);
and U19506 (N_19506,N_19339,N_19399);
and U19507 (N_19507,N_19234,N_19320);
nor U19508 (N_19508,N_19280,N_19316);
and U19509 (N_19509,N_19234,N_19210);
xor U19510 (N_19510,N_19327,N_19289);
or U19511 (N_19511,N_19310,N_19275);
and U19512 (N_19512,N_19343,N_19305);
xnor U19513 (N_19513,N_19364,N_19384);
nand U19514 (N_19514,N_19262,N_19230);
nand U19515 (N_19515,N_19275,N_19214);
or U19516 (N_19516,N_19277,N_19298);
nor U19517 (N_19517,N_19332,N_19323);
nand U19518 (N_19518,N_19210,N_19398);
nor U19519 (N_19519,N_19219,N_19385);
xor U19520 (N_19520,N_19207,N_19260);
nand U19521 (N_19521,N_19300,N_19286);
or U19522 (N_19522,N_19202,N_19283);
and U19523 (N_19523,N_19236,N_19290);
and U19524 (N_19524,N_19226,N_19208);
nand U19525 (N_19525,N_19303,N_19244);
xnor U19526 (N_19526,N_19287,N_19379);
or U19527 (N_19527,N_19372,N_19309);
nand U19528 (N_19528,N_19253,N_19381);
nand U19529 (N_19529,N_19395,N_19298);
nor U19530 (N_19530,N_19233,N_19260);
and U19531 (N_19531,N_19246,N_19385);
and U19532 (N_19532,N_19365,N_19254);
and U19533 (N_19533,N_19250,N_19307);
nand U19534 (N_19534,N_19358,N_19264);
nor U19535 (N_19535,N_19211,N_19360);
and U19536 (N_19536,N_19207,N_19304);
or U19537 (N_19537,N_19344,N_19285);
and U19538 (N_19538,N_19207,N_19226);
or U19539 (N_19539,N_19255,N_19349);
or U19540 (N_19540,N_19369,N_19310);
nor U19541 (N_19541,N_19209,N_19218);
or U19542 (N_19542,N_19215,N_19399);
and U19543 (N_19543,N_19319,N_19239);
nand U19544 (N_19544,N_19254,N_19233);
nor U19545 (N_19545,N_19282,N_19375);
nand U19546 (N_19546,N_19211,N_19337);
xor U19547 (N_19547,N_19250,N_19357);
nor U19548 (N_19548,N_19387,N_19364);
nor U19549 (N_19549,N_19348,N_19399);
xnor U19550 (N_19550,N_19375,N_19275);
and U19551 (N_19551,N_19244,N_19358);
and U19552 (N_19552,N_19346,N_19269);
nand U19553 (N_19553,N_19363,N_19354);
and U19554 (N_19554,N_19371,N_19264);
or U19555 (N_19555,N_19284,N_19295);
or U19556 (N_19556,N_19235,N_19300);
nor U19557 (N_19557,N_19398,N_19374);
and U19558 (N_19558,N_19312,N_19250);
nand U19559 (N_19559,N_19231,N_19385);
nor U19560 (N_19560,N_19321,N_19390);
xnor U19561 (N_19561,N_19398,N_19291);
or U19562 (N_19562,N_19297,N_19320);
or U19563 (N_19563,N_19366,N_19277);
and U19564 (N_19564,N_19200,N_19231);
or U19565 (N_19565,N_19253,N_19230);
and U19566 (N_19566,N_19237,N_19224);
nand U19567 (N_19567,N_19382,N_19325);
xnor U19568 (N_19568,N_19391,N_19336);
or U19569 (N_19569,N_19271,N_19391);
xnor U19570 (N_19570,N_19236,N_19258);
or U19571 (N_19571,N_19374,N_19246);
and U19572 (N_19572,N_19372,N_19282);
xnor U19573 (N_19573,N_19232,N_19229);
or U19574 (N_19574,N_19280,N_19365);
or U19575 (N_19575,N_19280,N_19262);
nor U19576 (N_19576,N_19397,N_19279);
nor U19577 (N_19577,N_19213,N_19272);
or U19578 (N_19578,N_19245,N_19271);
nor U19579 (N_19579,N_19332,N_19368);
nor U19580 (N_19580,N_19256,N_19343);
or U19581 (N_19581,N_19321,N_19373);
and U19582 (N_19582,N_19285,N_19247);
and U19583 (N_19583,N_19237,N_19265);
nor U19584 (N_19584,N_19375,N_19255);
nor U19585 (N_19585,N_19319,N_19261);
nand U19586 (N_19586,N_19388,N_19276);
xor U19587 (N_19587,N_19313,N_19226);
nand U19588 (N_19588,N_19391,N_19267);
nor U19589 (N_19589,N_19339,N_19227);
xor U19590 (N_19590,N_19283,N_19391);
nor U19591 (N_19591,N_19220,N_19280);
nand U19592 (N_19592,N_19299,N_19252);
xor U19593 (N_19593,N_19379,N_19350);
nor U19594 (N_19594,N_19316,N_19344);
and U19595 (N_19595,N_19241,N_19211);
nand U19596 (N_19596,N_19330,N_19391);
nand U19597 (N_19597,N_19351,N_19215);
nor U19598 (N_19598,N_19388,N_19253);
and U19599 (N_19599,N_19241,N_19222);
and U19600 (N_19600,N_19450,N_19446);
and U19601 (N_19601,N_19421,N_19560);
nor U19602 (N_19602,N_19443,N_19423);
or U19603 (N_19603,N_19461,N_19478);
and U19604 (N_19604,N_19514,N_19437);
nor U19605 (N_19605,N_19508,N_19528);
nor U19606 (N_19606,N_19559,N_19473);
and U19607 (N_19607,N_19518,N_19536);
and U19608 (N_19608,N_19438,N_19474);
xor U19609 (N_19609,N_19400,N_19532);
and U19610 (N_19610,N_19415,N_19545);
xor U19611 (N_19611,N_19599,N_19554);
nor U19612 (N_19612,N_19422,N_19420);
and U19613 (N_19613,N_19491,N_19529);
and U19614 (N_19614,N_19572,N_19431);
and U19615 (N_19615,N_19436,N_19577);
xor U19616 (N_19616,N_19558,N_19569);
nor U19617 (N_19617,N_19439,N_19496);
nor U19618 (N_19618,N_19494,N_19477);
nand U19619 (N_19619,N_19495,N_19499);
or U19620 (N_19620,N_19588,N_19406);
or U19621 (N_19621,N_19498,N_19425);
xnor U19622 (N_19622,N_19482,N_19523);
or U19623 (N_19623,N_19540,N_19480);
nor U19624 (N_19624,N_19410,N_19463);
nor U19625 (N_19625,N_19427,N_19513);
nand U19626 (N_19626,N_19505,N_19575);
or U19627 (N_19627,N_19527,N_19485);
or U19628 (N_19628,N_19563,N_19549);
and U19629 (N_19629,N_19530,N_19489);
nor U19630 (N_19630,N_19497,N_19409);
xor U19631 (N_19631,N_19565,N_19592);
and U19632 (N_19632,N_19524,N_19441);
nand U19633 (N_19633,N_19598,N_19465);
nand U19634 (N_19634,N_19475,N_19571);
xnor U19635 (N_19635,N_19447,N_19542);
xnor U19636 (N_19636,N_19506,N_19457);
nand U19637 (N_19637,N_19416,N_19411);
nand U19638 (N_19638,N_19589,N_19580);
xor U19639 (N_19639,N_19511,N_19440);
xnor U19640 (N_19640,N_19552,N_19404);
nand U19641 (N_19641,N_19548,N_19471);
xnor U19642 (N_19642,N_19551,N_19403);
nor U19643 (N_19643,N_19476,N_19417);
or U19644 (N_19644,N_19526,N_19566);
nand U19645 (N_19645,N_19553,N_19525);
or U19646 (N_19646,N_19546,N_19587);
nor U19647 (N_19647,N_19591,N_19585);
nor U19648 (N_19648,N_19493,N_19504);
xor U19649 (N_19649,N_19466,N_19573);
or U19650 (N_19650,N_19462,N_19448);
and U19651 (N_19651,N_19509,N_19490);
nor U19652 (N_19652,N_19481,N_19444);
and U19653 (N_19653,N_19539,N_19564);
xnor U19654 (N_19654,N_19533,N_19512);
and U19655 (N_19655,N_19574,N_19576);
xnor U19656 (N_19656,N_19453,N_19584);
nor U19657 (N_19657,N_19555,N_19405);
and U19658 (N_19658,N_19593,N_19556);
or U19659 (N_19659,N_19590,N_19483);
and U19660 (N_19660,N_19412,N_19451);
or U19661 (N_19661,N_19517,N_19429);
nand U19662 (N_19662,N_19586,N_19547);
or U19663 (N_19663,N_19428,N_19492);
nor U19664 (N_19664,N_19487,N_19522);
and U19665 (N_19665,N_19435,N_19433);
and U19666 (N_19666,N_19458,N_19583);
nor U19667 (N_19667,N_19541,N_19596);
and U19668 (N_19668,N_19515,N_19452);
nand U19669 (N_19669,N_19460,N_19470);
or U19670 (N_19670,N_19418,N_19455);
nand U19671 (N_19671,N_19402,N_19501);
or U19672 (N_19672,N_19567,N_19516);
and U19673 (N_19673,N_19503,N_19520);
or U19674 (N_19674,N_19432,N_19484);
and U19675 (N_19675,N_19449,N_19500);
nor U19676 (N_19676,N_19595,N_19456);
xnor U19677 (N_19677,N_19519,N_19543);
nor U19678 (N_19678,N_19434,N_19582);
nand U19679 (N_19679,N_19568,N_19464);
and U19680 (N_19680,N_19561,N_19510);
or U19681 (N_19681,N_19413,N_19454);
nor U19682 (N_19682,N_19579,N_19581);
xnor U19683 (N_19683,N_19430,N_19537);
or U19684 (N_19684,N_19424,N_19414);
and U19685 (N_19685,N_19468,N_19538);
nand U19686 (N_19686,N_19597,N_19488);
nand U19687 (N_19687,N_19507,N_19459);
nand U19688 (N_19688,N_19467,N_19426);
xnor U19689 (N_19689,N_19419,N_19534);
xnor U19690 (N_19690,N_19521,N_19557);
or U19691 (N_19691,N_19442,N_19445);
xnor U19692 (N_19692,N_19472,N_19479);
or U19693 (N_19693,N_19486,N_19469);
xnor U19694 (N_19694,N_19544,N_19550);
nor U19695 (N_19695,N_19408,N_19594);
and U19696 (N_19696,N_19531,N_19502);
nand U19697 (N_19697,N_19535,N_19407);
xor U19698 (N_19698,N_19562,N_19570);
and U19699 (N_19699,N_19401,N_19578);
xnor U19700 (N_19700,N_19407,N_19423);
xor U19701 (N_19701,N_19517,N_19402);
nor U19702 (N_19702,N_19599,N_19585);
or U19703 (N_19703,N_19474,N_19533);
and U19704 (N_19704,N_19566,N_19518);
xnor U19705 (N_19705,N_19445,N_19549);
and U19706 (N_19706,N_19454,N_19440);
and U19707 (N_19707,N_19400,N_19439);
and U19708 (N_19708,N_19538,N_19557);
or U19709 (N_19709,N_19488,N_19430);
or U19710 (N_19710,N_19562,N_19569);
nand U19711 (N_19711,N_19597,N_19507);
xnor U19712 (N_19712,N_19421,N_19456);
and U19713 (N_19713,N_19570,N_19455);
and U19714 (N_19714,N_19564,N_19583);
or U19715 (N_19715,N_19461,N_19546);
or U19716 (N_19716,N_19422,N_19459);
or U19717 (N_19717,N_19449,N_19472);
xor U19718 (N_19718,N_19448,N_19456);
nand U19719 (N_19719,N_19527,N_19549);
nand U19720 (N_19720,N_19598,N_19477);
xor U19721 (N_19721,N_19506,N_19545);
nand U19722 (N_19722,N_19510,N_19477);
or U19723 (N_19723,N_19403,N_19404);
nor U19724 (N_19724,N_19510,N_19586);
or U19725 (N_19725,N_19537,N_19472);
nor U19726 (N_19726,N_19574,N_19571);
xnor U19727 (N_19727,N_19540,N_19539);
xnor U19728 (N_19728,N_19495,N_19468);
xnor U19729 (N_19729,N_19429,N_19560);
or U19730 (N_19730,N_19468,N_19471);
nand U19731 (N_19731,N_19527,N_19430);
nor U19732 (N_19732,N_19593,N_19481);
and U19733 (N_19733,N_19562,N_19542);
or U19734 (N_19734,N_19558,N_19430);
or U19735 (N_19735,N_19497,N_19566);
xor U19736 (N_19736,N_19574,N_19419);
nor U19737 (N_19737,N_19546,N_19552);
and U19738 (N_19738,N_19554,N_19498);
nand U19739 (N_19739,N_19567,N_19407);
xor U19740 (N_19740,N_19502,N_19493);
nor U19741 (N_19741,N_19513,N_19410);
and U19742 (N_19742,N_19533,N_19444);
nand U19743 (N_19743,N_19564,N_19453);
xnor U19744 (N_19744,N_19489,N_19552);
nor U19745 (N_19745,N_19419,N_19570);
or U19746 (N_19746,N_19460,N_19550);
nand U19747 (N_19747,N_19514,N_19455);
or U19748 (N_19748,N_19584,N_19409);
nor U19749 (N_19749,N_19440,N_19529);
nand U19750 (N_19750,N_19552,N_19469);
nand U19751 (N_19751,N_19516,N_19495);
and U19752 (N_19752,N_19435,N_19475);
nand U19753 (N_19753,N_19544,N_19478);
or U19754 (N_19754,N_19523,N_19521);
nor U19755 (N_19755,N_19569,N_19454);
nand U19756 (N_19756,N_19485,N_19500);
nand U19757 (N_19757,N_19455,N_19583);
and U19758 (N_19758,N_19588,N_19404);
nor U19759 (N_19759,N_19401,N_19529);
nand U19760 (N_19760,N_19583,N_19430);
or U19761 (N_19761,N_19449,N_19593);
nand U19762 (N_19762,N_19479,N_19540);
and U19763 (N_19763,N_19587,N_19549);
and U19764 (N_19764,N_19434,N_19448);
or U19765 (N_19765,N_19484,N_19557);
and U19766 (N_19766,N_19488,N_19591);
xnor U19767 (N_19767,N_19433,N_19539);
nor U19768 (N_19768,N_19416,N_19510);
or U19769 (N_19769,N_19452,N_19451);
or U19770 (N_19770,N_19592,N_19573);
nor U19771 (N_19771,N_19543,N_19563);
and U19772 (N_19772,N_19447,N_19552);
xor U19773 (N_19773,N_19449,N_19436);
xor U19774 (N_19774,N_19507,N_19530);
and U19775 (N_19775,N_19518,N_19465);
xor U19776 (N_19776,N_19571,N_19521);
nor U19777 (N_19777,N_19442,N_19538);
nor U19778 (N_19778,N_19516,N_19520);
xor U19779 (N_19779,N_19574,N_19424);
nand U19780 (N_19780,N_19428,N_19404);
or U19781 (N_19781,N_19553,N_19478);
or U19782 (N_19782,N_19536,N_19500);
xnor U19783 (N_19783,N_19479,N_19474);
xor U19784 (N_19784,N_19437,N_19492);
nand U19785 (N_19785,N_19441,N_19434);
nor U19786 (N_19786,N_19485,N_19458);
nand U19787 (N_19787,N_19414,N_19401);
and U19788 (N_19788,N_19482,N_19430);
nand U19789 (N_19789,N_19428,N_19539);
and U19790 (N_19790,N_19526,N_19439);
nor U19791 (N_19791,N_19420,N_19555);
and U19792 (N_19792,N_19434,N_19497);
and U19793 (N_19793,N_19442,N_19431);
nand U19794 (N_19794,N_19526,N_19425);
xnor U19795 (N_19795,N_19576,N_19481);
and U19796 (N_19796,N_19442,N_19482);
and U19797 (N_19797,N_19564,N_19472);
nor U19798 (N_19798,N_19401,N_19446);
nand U19799 (N_19799,N_19425,N_19521);
xor U19800 (N_19800,N_19655,N_19658);
xor U19801 (N_19801,N_19755,N_19652);
nor U19802 (N_19802,N_19684,N_19646);
and U19803 (N_19803,N_19781,N_19709);
nand U19804 (N_19804,N_19644,N_19727);
and U19805 (N_19805,N_19676,N_19793);
xnor U19806 (N_19806,N_19777,N_19617);
nand U19807 (N_19807,N_19724,N_19687);
nor U19808 (N_19808,N_19739,N_19673);
xnor U19809 (N_19809,N_19651,N_19785);
nor U19810 (N_19810,N_19650,N_19730);
and U19811 (N_19811,N_19647,N_19678);
nand U19812 (N_19812,N_19754,N_19633);
or U19813 (N_19813,N_19604,N_19728);
xor U19814 (N_19814,N_19677,N_19792);
or U19815 (N_19815,N_19611,N_19758);
nor U19816 (N_19816,N_19714,N_19643);
and U19817 (N_19817,N_19613,N_19787);
xor U19818 (N_19818,N_19736,N_19697);
xnor U19819 (N_19819,N_19671,N_19774);
and U19820 (N_19820,N_19693,N_19608);
nor U19821 (N_19821,N_19699,N_19723);
nand U19822 (N_19822,N_19675,N_19601);
or U19823 (N_19823,N_19745,N_19702);
nand U19824 (N_19824,N_19708,N_19635);
and U19825 (N_19825,N_19737,N_19609);
nand U19826 (N_19826,N_19649,N_19600);
and U19827 (N_19827,N_19603,N_19701);
or U19828 (N_19828,N_19641,N_19756);
or U19829 (N_19829,N_19784,N_19744);
nand U19830 (N_19830,N_19731,N_19732);
or U19831 (N_19831,N_19757,N_19707);
or U19832 (N_19832,N_19624,N_19686);
or U19833 (N_19833,N_19768,N_19656);
and U19834 (N_19834,N_19639,N_19782);
nor U19835 (N_19835,N_19743,N_19668);
or U19836 (N_19836,N_19704,N_19741);
nand U19837 (N_19837,N_19796,N_19627);
and U19838 (N_19838,N_19630,N_19778);
and U19839 (N_19839,N_19761,N_19621);
nand U19840 (N_19840,N_19672,N_19626);
xor U19841 (N_19841,N_19753,N_19712);
and U19842 (N_19842,N_19645,N_19640);
nor U19843 (N_19843,N_19716,N_19713);
and U19844 (N_19844,N_19762,N_19666);
nand U19845 (N_19845,N_19706,N_19629);
nor U19846 (N_19846,N_19726,N_19663);
xnor U19847 (N_19847,N_19606,N_19694);
nand U19848 (N_19848,N_19794,N_19715);
nor U19849 (N_19849,N_19789,N_19729);
or U19850 (N_19850,N_19690,N_19700);
nor U19851 (N_19851,N_19660,N_19773);
or U19852 (N_19852,N_19740,N_19692);
and U19853 (N_19853,N_19725,N_19642);
xor U19854 (N_19854,N_19669,N_19685);
nor U19855 (N_19855,N_19764,N_19683);
or U19856 (N_19856,N_19602,N_19711);
xnor U19857 (N_19857,N_19664,N_19798);
or U19858 (N_19858,N_19797,N_19760);
and U19859 (N_19859,N_19619,N_19628);
xor U19860 (N_19860,N_19657,N_19667);
or U19861 (N_19861,N_19654,N_19780);
nor U19862 (N_19862,N_19623,N_19747);
nand U19863 (N_19863,N_19665,N_19607);
or U19864 (N_19864,N_19662,N_19636);
and U19865 (N_19865,N_19682,N_19750);
and U19866 (N_19866,N_19696,N_19634);
nor U19867 (N_19867,N_19795,N_19612);
xnor U19868 (N_19868,N_19749,N_19772);
and U19869 (N_19869,N_19638,N_19766);
or U19870 (N_19870,N_19738,N_19679);
and U19871 (N_19871,N_19615,N_19763);
or U19872 (N_19872,N_19614,N_19681);
nand U19873 (N_19873,N_19776,N_19653);
or U19874 (N_19874,N_19670,N_19661);
and U19875 (N_19875,N_19786,N_19748);
nand U19876 (N_19876,N_19721,N_19735);
xnor U19877 (N_19877,N_19703,N_19746);
or U19878 (N_19878,N_19659,N_19717);
or U19879 (N_19879,N_19759,N_19783);
nand U19880 (N_19880,N_19698,N_19771);
and U19881 (N_19881,N_19791,N_19720);
nor U19882 (N_19882,N_19674,N_19637);
nor U19883 (N_19883,N_19742,N_19734);
and U19884 (N_19884,N_19616,N_19775);
xor U19885 (N_19885,N_19790,N_19769);
or U19886 (N_19886,N_19689,N_19765);
nand U19887 (N_19887,N_19719,N_19620);
or U19888 (N_19888,N_19722,N_19788);
or U19889 (N_19889,N_19631,N_19733);
xnor U19890 (N_19890,N_19752,N_19770);
xor U19891 (N_19891,N_19610,N_19688);
and U19892 (N_19892,N_19695,N_19705);
and U19893 (N_19893,N_19618,N_19622);
or U19894 (N_19894,N_19779,N_19632);
nand U19895 (N_19895,N_19718,N_19680);
nor U19896 (N_19896,N_19767,N_19710);
xor U19897 (N_19897,N_19799,N_19751);
xnor U19898 (N_19898,N_19605,N_19691);
or U19899 (N_19899,N_19625,N_19648);
or U19900 (N_19900,N_19633,N_19654);
and U19901 (N_19901,N_19604,N_19726);
nor U19902 (N_19902,N_19763,N_19625);
xnor U19903 (N_19903,N_19642,N_19631);
nor U19904 (N_19904,N_19663,N_19795);
nand U19905 (N_19905,N_19712,N_19690);
nor U19906 (N_19906,N_19674,N_19731);
nor U19907 (N_19907,N_19649,N_19615);
xnor U19908 (N_19908,N_19758,N_19735);
or U19909 (N_19909,N_19644,N_19602);
nand U19910 (N_19910,N_19728,N_19791);
nand U19911 (N_19911,N_19718,N_19708);
nand U19912 (N_19912,N_19714,N_19691);
or U19913 (N_19913,N_19606,N_19619);
nor U19914 (N_19914,N_19663,N_19790);
nor U19915 (N_19915,N_19662,N_19706);
or U19916 (N_19916,N_19714,N_19793);
nor U19917 (N_19917,N_19620,N_19654);
or U19918 (N_19918,N_19666,N_19600);
nand U19919 (N_19919,N_19662,N_19638);
or U19920 (N_19920,N_19769,N_19627);
or U19921 (N_19921,N_19658,N_19723);
nand U19922 (N_19922,N_19723,N_19725);
nor U19923 (N_19923,N_19796,N_19781);
nor U19924 (N_19924,N_19741,N_19734);
xor U19925 (N_19925,N_19786,N_19608);
or U19926 (N_19926,N_19785,N_19722);
nand U19927 (N_19927,N_19716,N_19773);
nand U19928 (N_19928,N_19732,N_19707);
and U19929 (N_19929,N_19659,N_19611);
xnor U19930 (N_19930,N_19695,N_19724);
nor U19931 (N_19931,N_19673,N_19729);
nand U19932 (N_19932,N_19766,N_19736);
nand U19933 (N_19933,N_19757,N_19681);
and U19934 (N_19934,N_19604,N_19732);
and U19935 (N_19935,N_19680,N_19640);
nand U19936 (N_19936,N_19757,N_19732);
nand U19937 (N_19937,N_19693,N_19705);
or U19938 (N_19938,N_19610,N_19789);
and U19939 (N_19939,N_19718,N_19694);
nand U19940 (N_19940,N_19611,N_19715);
nor U19941 (N_19941,N_19639,N_19758);
nor U19942 (N_19942,N_19699,N_19766);
nor U19943 (N_19943,N_19712,N_19662);
or U19944 (N_19944,N_19792,N_19614);
and U19945 (N_19945,N_19616,N_19759);
nor U19946 (N_19946,N_19753,N_19686);
or U19947 (N_19947,N_19750,N_19763);
nand U19948 (N_19948,N_19785,N_19793);
xnor U19949 (N_19949,N_19692,N_19687);
and U19950 (N_19950,N_19691,N_19628);
xnor U19951 (N_19951,N_19628,N_19716);
or U19952 (N_19952,N_19641,N_19628);
nor U19953 (N_19953,N_19766,N_19612);
or U19954 (N_19954,N_19737,N_19694);
and U19955 (N_19955,N_19770,N_19620);
xnor U19956 (N_19956,N_19627,N_19790);
nor U19957 (N_19957,N_19661,N_19776);
nand U19958 (N_19958,N_19779,N_19765);
xnor U19959 (N_19959,N_19711,N_19655);
or U19960 (N_19960,N_19717,N_19676);
nor U19961 (N_19961,N_19629,N_19618);
and U19962 (N_19962,N_19628,N_19624);
xor U19963 (N_19963,N_19730,N_19710);
nand U19964 (N_19964,N_19617,N_19772);
and U19965 (N_19965,N_19730,N_19720);
nor U19966 (N_19966,N_19794,N_19615);
or U19967 (N_19967,N_19623,N_19602);
nand U19968 (N_19968,N_19669,N_19688);
and U19969 (N_19969,N_19755,N_19697);
nand U19970 (N_19970,N_19708,N_19668);
xnor U19971 (N_19971,N_19748,N_19696);
xor U19972 (N_19972,N_19785,N_19611);
nor U19973 (N_19973,N_19772,N_19670);
and U19974 (N_19974,N_19650,N_19627);
xor U19975 (N_19975,N_19787,N_19749);
nor U19976 (N_19976,N_19603,N_19784);
nand U19977 (N_19977,N_19639,N_19727);
nand U19978 (N_19978,N_19696,N_19765);
xnor U19979 (N_19979,N_19771,N_19657);
or U19980 (N_19980,N_19700,N_19764);
nand U19981 (N_19981,N_19640,N_19728);
nor U19982 (N_19982,N_19701,N_19711);
nor U19983 (N_19983,N_19669,N_19698);
or U19984 (N_19984,N_19705,N_19760);
nand U19985 (N_19985,N_19678,N_19736);
nand U19986 (N_19986,N_19760,N_19656);
or U19987 (N_19987,N_19633,N_19712);
xor U19988 (N_19988,N_19743,N_19752);
nor U19989 (N_19989,N_19740,N_19774);
xor U19990 (N_19990,N_19631,N_19650);
nor U19991 (N_19991,N_19742,N_19660);
xnor U19992 (N_19992,N_19774,N_19709);
nor U19993 (N_19993,N_19698,N_19665);
xnor U19994 (N_19994,N_19623,N_19613);
nand U19995 (N_19995,N_19643,N_19780);
and U19996 (N_19996,N_19744,N_19713);
and U19997 (N_19997,N_19600,N_19607);
and U19998 (N_19998,N_19785,N_19704);
nor U19999 (N_19999,N_19667,N_19701);
or U20000 (N_20000,N_19898,N_19875);
nor U20001 (N_20001,N_19928,N_19947);
or U20002 (N_20002,N_19888,N_19852);
and U20003 (N_20003,N_19800,N_19986);
nand U20004 (N_20004,N_19809,N_19886);
and U20005 (N_20005,N_19818,N_19835);
nand U20006 (N_20006,N_19938,N_19868);
and U20007 (N_20007,N_19906,N_19833);
nor U20008 (N_20008,N_19870,N_19806);
xor U20009 (N_20009,N_19950,N_19953);
and U20010 (N_20010,N_19987,N_19983);
and U20011 (N_20011,N_19879,N_19894);
or U20012 (N_20012,N_19940,N_19854);
xnor U20013 (N_20013,N_19831,N_19982);
or U20014 (N_20014,N_19985,N_19805);
or U20015 (N_20015,N_19922,N_19810);
xor U20016 (N_20016,N_19943,N_19874);
nand U20017 (N_20017,N_19878,N_19801);
and U20018 (N_20018,N_19964,N_19904);
or U20019 (N_20019,N_19827,N_19908);
and U20020 (N_20020,N_19944,N_19926);
nand U20021 (N_20021,N_19816,N_19889);
nor U20022 (N_20022,N_19897,N_19814);
nor U20023 (N_20023,N_19837,N_19841);
xor U20024 (N_20024,N_19887,N_19861);
and U20025 (N_20025,N_19895,N_19807);
or U20026 (N_20026,N_19804,N_19910);
nand U20027 (N_20027,N_19939,N_19951);
xor U20028 (N_20028,N_19994,N_19933);
xor U20029 (N_20029,N_19975,N_19960);
nand U20030 (N_20030,N_19919,N_19967);
nand U20031 (N_20031,N_19976,N_19920);
nor U20032 (N_20032,N_19819,N_19932);
xor U20033 (N_20033,N_19851,N_19813);
nand U20034 (N_20034,N_19902,N_19823);
or U20035 (N_20035,N_19996,N_19999);
xnor U20036 (N_20036,N_19912,N_19812);
nor U20037 (N_20037,N_19963,N_19839);
nand U20038 (N_20038,N_19990,N_19991);
nand U20039 (N_20039,N_19855,N_19873);
and U20040 (N_20040,N_19821,N_19826);
nand U20041 (N_20041,N_19907,N_19829);
and U20042 (N_20042,N_19850,N_19853);
xnor U20043 (N_20043,N_19952,N_19915);
and U20044 (N_20044,N_19803,N_19935);
xor U20045 (N_20045,N_19825,N_19890);
or U20046 (N_20046,N_19929,N_19942);
nor U20047 (N_20047,N_19838,N_19927);
nand U20048 (N_20048,N_19941,N_19903);
or U20049 (N_20049,N_19884,N_19974);
nor U20050 (N_20050,N_19867,N_19840);
or U20051 (N_20051,N_19900,N_19844);
or U20052 (N_20052,N_19945,N_19980);
xor U20053 (N_20053,N_19877,N_19989);
nand U20054 (N_20054,N_19899,N_19828);
and U20055 (N_20055,N_19917,N_19862);
xor U20056 (N_20056,N_19923,N_19857);
nor U20057 (N_20057,N_19968,N_19921);
nand U20058 (N_20058,N_19859,N_19824);
xnor U20059 (N_20059,N_19811,N_19865);
or U20060 (N_20060,N_19965,N_19891);
and U20061 (N_20061,N_19869,N_19988);
or U20062 (N_20062,N_19843,N_19849);
nand U20063 (N_20063,N_19957,N_19918);
xnor U20064 (N_20064,N_19970,N_19848);
xnor U20065 (N_20065,N_19836,N_19961);
nand U20066 (N_20066,N_19820,N_19832);
xnor U20067 (N_20067,N_19883,N_19866);
or U20068 (N_20068,N_19981,N_19893);
or U20069 (N_20069,N_19872,N_19969);
nor U20070 (N_20070,N_19949,N_19937);
xor U20071 (N_20071,N_19934,N_19973);
xnor U20072 (N_20072,N_19846,N_19930);
nand U20073 (N_20073,N_19822,N_19905);
nor U20074 (N_20074,N_19880,N_19931);
and U20075 (N_20075,N_19842,N_19864);
nand U20076 (N_20076,N_19966,N_19909);
nor U20077 (N_20077,N_19863,N_19911);
xnor U20078 (N_20078,N_19815,N_19858);
nand U20079 (N_20079,N_19992,N_19972);
and U20080 (N_20080,N_19955,N_19896);
nand U20081 (N_20081,N_19881,N_19871);
nand U20082 (N_20082,N_19856,N_19808);
or U20083 (N_20083,N_19847,N_19830);
or U20084 (N_20084,N_19882,N_19916);
xor U20085 (N_20085,N_19925,N_19914);
or U20086 (N_20086,N_19971,N_19948);
nor U20087 (N_20087,N_19995,N_19901);
xnor U20088 (N_20088,N_19998,N_19913);
nor U20089 (N_20089,N_19984,N_19892);
xnor U20090 (N_20090,N_19924,N_19977);
xnor U20091 (N_20091,N_19979,N_19834);
nand U20092 (N_20092,N_19997,N_19860);
and U20093 (N_20093,N_19959,N_19958);
or U20094 (N_20094,N_19993,N_19802);
xor U20095 (N_20095,N_19946,N_19817);
and U20096 (N_20096,N_19936,N_19956);
or U20097 (N_20097,N_19885,N_19978);
nor U20098 (N_20098,N_19954,N_19845);
nor U20099 (N_20099,N_19876,N_19962);
or U20100 (N_20100,N_19805,N_19878);
and U20101 (N_20101,N_19924,N_19968);
nand U20102 (N_20102,N_19820,N_19840);
and U20103 (N_20103,N_19812,N_19864);
or U20104 (N_20104,N_19980,N_19865);
nor U20105 (N_20105,N_19937,N_19924);
xor U20106 (N_20106,N_19982,N_19941);
or U20107 (N_20107,N_19888,N_19997);
and U20108 (N_20108,N_19866,N_19824);
and U20109 (N_20109,N_19805,N_19809);
or U20110 (N_20110,N_19848,N_19924);
or U20111 (N_20111,N_19814,N_19856);
and U20112 (N_20112,N_19808,N_19985);
xor U20113 (N_20113,N_19899,N_19975);
nand U20114 (N_20114,N_19892,N_19916);
nor U20115 (N_20115,N_19901,N_19953);
and U20116 (N_20116,N_19868,N_19947);
and U20117 (N_20117,N_19879,N_19966);
nand U20118 (N_20118,N_19978,N_19853);
nand U20119 (N_20119,N_19926,N_19941);
and U20120 (N_20120,N_19933,N_19822);
and U20121 (N_20121,N_19812,N_19844);
or U20122 (N_20122,N_19897,N_19921);
xor U20123 (N_20123,N_19959,N_19818);
nor U20124 (N_20124,N_19811,N_19804);
or U20125 (N_20125,N_19902,N_19809);
nand U20126 (N_20126,N_19931,N_19884);
nor U20127 (N_20127,N_19891,N_19915);
nand U20128 (N_20128,N_19957,N_19926);
xnor U20129 (N_20129,N_19980,N_19891);
xnor U20130 (N_20130,N_19937,N_19999);
and U20131 (N_20131,N_19910,N_19933);
and U20132 (N_20132,N_19859,N_19894);
nor U20133 (N_20133,N_19965,N_19827);
or U20134 (N_20134,N_19901,N_19998);
and U20135 (N_20135,N_19951,N_19959);
or U20136 (N_20136,N_19983,N_19932);
nand U20137 (N_20137,N_19831,N_19859);
xor U20138 (N_20138,N_19956,N_19870);
nor U20139 (N_20139,N_19841,N_19931);
and U20140 (N_20140,N_19864,N_19804);
nor U20141 (N_20141,N_19912,N_19930);
or U20142 (N_20142,N_19958,N_19915);
xor U20143 (N_20143,N_19930,N_19878);
nand U20144 (N_20144,N_19987,N_19843);
xor U20145 (N_20145,N_19804,N_19959);
nand U20146 (N_20146,N_19956,N_19992);
or U20147 (N_20147,N_19863,N_19879);
nand U20148 (N_20148,N_19922,N_19872);
nor U20149 (N_20149,N_19922,N_19921);
nand U20150 (N_20150,N_19877,N_19823);
xnor U20151 (N_20151,N_19855,N_19918);
or U20152 (N_20152,N_19803,N_19924);
and U20153 (N_20153,N_19956,N_19803);
or U20154 (N_20154,N_19839,N_19882);
or U20155 (N_20155,N_19946,N_19834);
nor U20156 (N_20156,N_19853,N_19875);
xnor U20157 (N_20157,N_19885,N_19973);
xnor U20158 (N_20158,N_19891,N_19816);
nor U20159 (N_20159,N_19924,N_19852);
xor U20160 (N_20160,N_19807,N_19892);
xor U20161 (N_20161,N_19908,N_19894);
xor U20162 (N_20162,N_19949,N_19870);
xor U20163 (N_20163,N_19874,N_19902);
xnor U20164 (N_20164,N_19954,N_19984);
or U20165 (N_20165,N_19852,N_19940);
nand U20166 (N_20166,N_19883,N_19948);
or U20167 (N_20167,N_19962,N_19848);
xor U20168 (N_20168,N_19976,N_19882);
and U20169 (N_20169,N_19940,N_19902);
and U20170 (N_20170,N_19968,N_19891);
and U20171 (N_20171,N_19965,N_19895);
nor U20172 (N_20172,N_19898,N_19961);
nor U20173 (N_20173,N_19999,N_19916);
nor U20174 (N_20174,N_19854,N_19857);
xnor U20175 (N_20175,N_19937,N_19863);
or U20176 (N_20176,N_19802,N_19946);
nor U20177 (N_20177,N_19807,N_19918);
nand U20178 (N_20178,N_19955,N_19830);
nand U20179 (N_20179,N_19881,N_19831);
xor U20180 (N_20180,N_19969,N_19997);
nor U20181 (N_20181,N_19887,N_19976);
or U20182 (N_20182,N_19816,N_19809);
nand U20183 (N_20183,N_19930,N_19808);
and U20184 (N_20184,N_19901,N_19913);
nor U20185 (N_20185,N_19989,N_19814);
xor U20186 (N_20186,N_19868,N_19934);
xor U20187 (N_20187,N_19845,N_19935);
and U20188 (N_20188,N_19926,N_19815);
or U20189 (N_20189,N_19974,N_19853);
xor U20190 (N_20190,N_19872,N_19905);
or U20191 (N_20191,N_19901,N_19882);
xnor U20192 (N_20192,N_19946,N_19941);
nand U20193 (N_20193,N_19862,N_19909);
nor U20194 (N_20194,N_19985,N_19828);
or U20195 (N_20195,N_19861,N_19865);
nand U20196 (N_20196,N_19837,N_19987);
nand U20197 (N_20197,N_19932,N_19955);
nand U20198 (N_20198,N_19827,N_19841);
xor U20199 (N_20199,N_19864,N_19832);
or U20200 (N_20200,N_20102,N_20131);
or U20201 (N_20201,N_20192,N_20035);
nand U20202 (N_20202,N_20175,N_20138);
and U20203 (N_20203,N_20031,N_20080);
nor U20204 (N_20204,N_20158,N_20045);
and U20205 (N_20205,N_20195,N_20147);
and U20206 (N_20206,N_20066,N_20086);
nor U20207 (N_20207,N_20083,N_20159);
nand U20208 (N_20208,N_20003,N_20129);
nand U20209 (N_20209,N_20120,N_20198);
nor U20210 (N_20210,N_20132,N_20028);
xnor U20211 (N_20211,N_20111,N_20104);
nor U20212 (N_20212,N_20133,N_20010);
and U20213 (N_20213,N_20013,N_20172);
and U20214 (N_20214,N_20163,N_20098);
and U20215 (N_20215,N_20089,N_20077);
xor U20216 (N_20216,N_20007,N_20157);
xor U20217 (N_20217,N_20014,N_20166);
and U20218 (N_20218,N_20069,N_20062);
or U20219 (N_20219,N_20092,N_20151);
and U20220 (N_20220,N_20054,N_20182);
and U20221 (N_20221,N_20115,N_20008);
xor U20222 (N_20222,N_20180,N_20162);
nand U20223 (N_20223,N_20072,N_20100);
nand U20224 (N_20224,N_20191,N_20029);
and U20225 (N_20225,N_20018,N_20169);
xor U20226 (N_20226,N_20012,N_20134);
or U20227 (N_20227,N_20020,N_20135);
xnor U20228 (N_20228,N_20081,N_20053);
or U20229 (N_20229,N_20095,N_20040);
or U20230 (N_20230,N_20124,N_20178);
nor U20231 (N_20231,N_20002,N_20064);
nor U20232 (N_20232,N_20137,N_20179);
xor U20233 (N_20233,N_20148,N_20041);
and U20234 (N_20234,N_20128,N_20055);
or U20235 (N_20235,N_20079,N_20156);
xnor U20236 (N_20236,N_20122,N_20042);
and U20237 (N_20237,N_20037,N_20052);
nand U20238 (N_20238,N_20142,N_20190);
nor U20239 (N_20239,N_20068,N_20170);
nand U20240 (N_20240,N_20161,N_20057);
nor U20241 (N_20241,N_20006,N_20094);
or U20242 (N_20242,N_20073,N_20181);
or U20243 (N_20243,N_20036,N_20183);
nor U20244 (N_20244,N_20032,N_20019);
nor U20245 (N_20245,N_20107,N_20177);
xnor U20246 (N_20246,N_20164,N_20034);
or U20247 (N_20247,N_20196,N_20143);
or U20248 (N_20248,N_20171,N_20165);
and U20249 (N_20249,N_20021,N_20011);
nand U20250 (N_20250,N_20155,N_20022);
or U20251 (N_20251,N_20103,N_20154);
xor U20252 (N_20252,N_20105,N_20121);
nor U20253 (N_20253,N_20000,N_20005);
and U20254 (N_20254,N_20146,N_20071);
and U20255 (N_20255,N_20091,N_20149);
nor U20256 (N_20256,N_20189,N_20194);
and U20257 (N_20257,N_20141,N_20173);
and U20258 (N_20258,N_20130,N_20090);
xnor U20259 (N_20259,N_20023,N_20174);
xnor U20260 (N_20260,N_20176,N_20009);
or U20261 (N_20261,N_20185,N_20075);
and U20262 (N_20262,N_20061,N_20015);
and U20263 (N_20263,N_20168,N_20106);
and U20264 (N_20264,N_20197,N_20160);
or U20265 (N_20265,N_20067,N_20026);
or U20266 (N_20266,N_20101,N_20060);
nand U20267 (N_20267,N_20199,N_20112);
or U20268 (N_20268,N_20016,N_20088);
nand U20269 (N_20269,N_20145,N_20150);
xnor U20270 (N_20270,N_20058,N_20187);
xor U20271 (N_20271,N_20044,N_20082);
xor U20272 (N_20272,N_20047,N_20184);
nand U20273 (N_20273,N_20004,N_20114);
or U20274 (N_20274,N_20096,N_20017);
xor U20275 (N_20275,N_20051,N_20118);
or U20276 (N_20276,N_20078,N_20070);
nand U20277 (N_20277,N_20125,N_20076);
or U20278 (N_20278,N_20050,N_20084);
nor U20279 (N_20279,N_20025,N_20065);
and U20280 (N_20280,N_20001,N_20074);
xor U20281 (N_20281,N_20108,N_20027);
nor U20282 (N_20282,N_20046,N_20043);
nand U20283 (N_20283,N_20099,N_20093);
or U20284 (N_20284,N_20063,N_20140);
or U20285 (N_20285,N_20024,N_20059);
xnor U20286 (N_20286,N_20116,N_20097);
xor U20287 (N_20287,N_20136,N_20186);
nor U20288 (N_20288,N_20153,N_20113);
nor U20289 (N_20289,N_20119,N_20049);
and U20290 (N_20290,N_20193,N_20056);
nand U20291 (N_20291,N_20085,N_20167);
or U20292 (N_20292,N_20139,N_20110);
or U20293 (N_20293,N_20030,N_20152);
xnor U20294 (N_20294,N_20117,N_20127);
or U20295 (N_20295,N_20126,N_20144);
or U20296 (N_20296,N_20048,N_20109);
nand U20297 (N_20297,N_20038,N_20123);
and U20298 (N_20298,N_20033,N_20188);
nand U20299 (N_20299,N_20087,N_20039);
xor U20300 (N_20300,N_20026,N_20190);
or U20301 (N_20301,N_20056,N_20194);
nand U20302 (N_20302,N_20096,N_20177);
nand U20303 (N_20303,N_20122,N_20081);
nor U20304 (N_20304,N_20069,N_20183);
xnor U20305 (N_20305,N_20197,N_20030);
nor U20306 (N_20306,N_20101,N_20194);
nor U20307 (N_20307,N_20166,N_20008);
nor U20308 (N_20308,N_20074,N_20089);
or U20309 (N_20309,N_20015,N_20141);
nor U20310 (N_20310,N_20057,N_20104);
or U20311 (N_20311,N_20143,N_20152);
nand U20312 (N_20312,N_20090,N_20029);
and U20313 (N_20313,N_20179,N_20011);
or U20314 (N_20314,N_20183,N_20051);
or U20315 (N_20315,N_20176,N_20041);
xnor U20316 (N_20316,N_20007,N_20142);
and U20317 (N_20317,N_20029,N_20186);
nor U20318 (N_20318,N_20049,N_20010);
xnor U20319 (N_20319,N_20196,N_20082);
nand U20320 (N_20320,N_20060,N_20047);
nor U20321 (N_20321,N_20160,N_20067);
nor U20322 (N_20322,N_20045,N_20103);
nor U20323 (N_20323,N_20107,N_20025);
or U20324 (N_20324,N_20188,N_20181);
nor U20325 (N_20325,N_20046,N_20127);
and U20326 (N_20326,N_20189,N_20036);
xnor U20327 (N_20327,N_20109,N_20030);
or U20328 (N_20328,N_20022,N_20105);
and U20329 (N_20329,N_20102,N_20142);
nor U20330 (N_20330,N_20145,N_20021);
and U20331 (N_20331,N_20144,N_20063);
and U20332 (N_20332,N_20006,N_20126);
xnor U20333 (N_20333,N_20192,N_20050);
or U20334 (N_20334,N_20105,N_20023);
and U20335 (N_20335,N_20094,N_20014);
and U20336 (N_20336,N_20006,N_20091);
xor U20337 (N_20337,N_20015,N_20093);
xor U20338 (N_20338,N_20194,N_20118);
nand U20339 (N_20339,N_20120,N_20117);
nand U20340 (N_20340,N_20093,N_20167);
nand U20341 (N_20341,N_20189,N_20042);
nand U20342 (N_20342,N_20156,N_20196);
nor U20343 (N_20343,N_20194,N_20043);
or U20344 (N_20344,N_20010,N_20101);
xor U20345 (N_20345,N_20087,N_20001);
xor U20346 (N_20346,N_20186,N_20067);
nand U20347 (N_20347,N_20154,N_20149);
or U20348 (N_20348,N_20069,N_20118);
xor U20349 (N_20349,N_20048,N_20097);
or U20350 (N_20350,N_20093,N_20116);
xor U20351 (N_20351,N_20053,N_20079);
nor U20352 (N_20352,N_20127,N_20087);
xor U20353 (N_20353,N_20032,N_20110);
xor U20354 (N_20354,N_20110,N_20197);
xor U20355 (N_20355,N_20197,N_20055);
xor U20356 (N_20356,N_20176,N_20025);
nor U20357 (N_20357,N_20156,N_20088);
xnor U20358 (N_20358,N_20003,N_20165);
or U20359 (N_20359,N_20197,N_20063);
nand U20360 (N_20360,N_20101,N_20190);
or U20361 (N_20361,N_20034,N_20184);
and U20362 (N_20362,N_20145,N_20175);
or U20363 (N_20363,N_20061,N_20093);
nand U20364 (N_20364,N_20103,N_20176);
nor U20365 (N_20365,N_20195,N_20039);
or U20366 (N_20366,N_20176,N_20106);
or U20367 (N_20367,N_20043,N_20081);
or U20368 (N_20368,N_20020,N_20115);
or U20369 (N_20369,N_20127,N_20097);
nor U20370 (N_20370,N_20189,N_20047);
xnor U20371 (N_20371,N_20170,N_20116);
nor U20372 (N_20372,N_20145,N_20193);
nand U20373 (N_20373,N_20176,N_20067);
xnor U20374 (N_20374,N_20190,N_20036);
nor U20375 (N_20375,N_20093,N_20071);
or U20376 (N_20376,N_20126,N_20073);
xnor U20377 (N_20377,N_20039,N_20151);
nand U20378 (N_20378,N_20022,N_20138);
xor U20379 (N_20379,N_20105,N_20077);
nor U20380 (N_20380,N_20113,N_20108);
nand U20381 (N_20381,N_20122,N_20058);
nand U20382 (N_20382,N_20092,N_20115);
or U20383 (N_20383,N_20074,N_20005);
nor U20384 (N_20384,N_20161,N_20104);
or U20385 (N_20385,N_20178,N_20029);
nor U20386 (N_20386,N_20132,N_20098);
nand U20387 (N_20387,N_20030,N_20171);
or U20388 (N_20388,N_20147,N_20132);
or U20389 (N_20389,N_20159,N_20038);
xor U20390 (N_20390,N_20191,N_20196);
xor U20391 (N_20391,N_20174,N_20048);
nor U20392 (N_20392,N_20032,N_20071);
nand U20393 (N_20393,N_20037,N_20050);
nor U20394 (N_20394,N_20199,N_20121);
or U20395 (N_20395,N_20076,N_20183);
or U20396 (N_20396,N_20009,N_20091);
nand U20397 (N_20397,N_20113,N_20107);
xor U20398 (N_20398,N_20112,N_20151);
nor U20399 (N_20399,N_20073,N_20132);
xnor U20400 (N_20400,N_20335,N_20290);
xor U20401 (N_20401,N_20285,N_20209);
nor U20402 (N_20402,N_20354,N_20389);
nor U20403 (N_20403,N_20367,N_20309);
and U20404 (N_20404,N_20321,N_20296);
nor U20405 (N_20405,N_20260,N_20327);
nor U20406 (N_20406,N_20228,N_20240);
nand U20407 (N_20407,N_20220,N_20250);
xnor U20408 (N_20408,N_20256,N_20274);
or U20409 (N_20409,N_20387,N_20230);
nor U20410 (N_20410,N_20324,N_20223);
nand U20411 (N_20411,N_20395,N_20392);
or U20412 (N_20412,N_20291,N_20337);
nand U20413 (N_20413,N_20259,N_20348);
nand U20414 (N_20414,N_20361,N_20264);
nand U20415 (N_20415,N_20272,N_20380);
nor U20416 (N_20416,N_20360,N_20333);
xnor U20417 (N_20417,N_20287,N_20301);
nor U20418 (N_20418,N_20233,N_20266);
nor U20419 (N_20419,N_20219,N_20334);
and U20420 (N_20420,N_20263,N_20307);
nand U20421 (N_20421,N_20273,N_20214);
and U20422 (N_20422,N_20341,N_20353);
xor U20423 (N_20423,N_20316,N_20247);
or U20424 (N_20424,N_20232,N_20339);
or U20425 (N_20425,N_20304,N_20236);
or U20426 (N_20426,N_20203,N_20217);
xor U20427 (N_20427,N_20234,N_20363);
xnor U20428 (N_20428,N_20325,N_20308);
and U20429 (N_20429,N_20295,N_20330);
nand U20430 (N_20430,N_20373,N_20237);
and U20431 (N_20431,N_20208,N_20344);
nand U20432 (N_20432,N_20218,N_20347);
and U20433 (N_20433,N_20311,N_20362);
or U20434 (N_20434,N_20338,N_20298);
and U20435 (N_20435,N_20229,N_20222);
nand U20436 (N_20436,N_20394,N_20286);
nand U20437 (N_20437,N_20224,N_20319);
and U20438 (N_20438,N_20352,N_20397);
nor U20439 (N_20439,N_20366,N_20281);
or U20440 (N_20440,N_20244,N_20215);
nand U20441 (N_20441,N_20378,N_20267);
nand U20442 (N_20442,N_20293,N_20205);
nor U20443 (N_20443,N_20204,N_20312);
nor U20444 (N_20444,N_20221,N_20386);
nor U20445 (N_20445,N_20279,N_20358);
and U20446 (N_20446,N_20270,N_20289);
xnor U20447 (N_20447,N_20235,N_20251);
or U20448 (N_20448,N_20346,N_20343);
and U20449 (N_20449,N_20246,N_20323);
or U20450 (N_20450,N_20328,N_20216);
or U20451 (N_20451,N_20258,N_20342);
or U20452 (N_20452,N_20269,N_20374);
nand U20453 (N_20453,N_20303,N_20288);
nand U20454 (N_20454,N_20369,N_20255);
or U20455 (N_20455,N_20261,N_20384);
or U20456 (N_20456,N_20372,N_20396);
nand U20457 (N_20457,N_20284,N_20315);
and U20458 (N_20458,N_20283,N_20375);
xor U20459 (N_20459,N_20207,N_20383);
nor U20460 (N_20460,N_20340,N_20359);
or U20461 (N_20461,N_20276,N_20271);
and U20462 (N_20462,N_20239,N_20297);
nand U20463 (N_20463,N_20379,N_20368);
and U20464 (N_20464,N_20249,N_20371);
nor U20465 (N_20465,N_20213,N_20331);
and U20466 (N_20466,N_20201,N_20355);
and U20467 (N_20467,N_20318,N_20227);
nor U20468 (N_20468,N_20243,N_20310);
nor U20469 (N_20469,N_20282,N_20351);
and U20470 (N_20470,N_20370,N_20275);
nand U20471 (N_20471,N_20305,N_20225);
xnor U20472 (N_20472,N_20390,N_20382);
xor U20473 (N_20473,N_20226,N_20320);
nand U20474 (N_20474,N_20211,N_20299);
nor U20475 (N_20475,N_20280,N_20391);
or U20476 (N_20476,N_20202,N_20306);
and U20477 (N_20477,N_20356,N_20254);
nand U20478 (N_20478,N_20399,N_20349);
and U20479 (N_20479,N_20268,N_20265);
or U20480 (N_20480,N_20350,N_20377);
nand U20481 (N_20481,N_20313,N_20252);
xor U20482 (N_20482,N_20257,N_20314);
and U20483 (N_20483,N_20238,N_20262);
nor U20484 (N_20484,N_20242,N_20388);
xor U20485 (N_20485,N_20277,N_20200);
nand U20486 (N_20486,N_20231,N_20253);
xor U20487 (N_20487,N_20248,N_20326);
and U20488 (N_20488,N_20365,N_20336);
nor U20489 (N_20489,N_20398,N_20376);
xor U20490 (N_20490,N_20381,N_20278);
nor U20491 (N_20491,N_20393,N_20210);
and U20492 (N_20492,N_20292,N_20212);
xnor U20493 (N_20493,N_20322,N_20357);
nor U20494 (N_20494,N_20241,N_20329);
and U20495 (N_20495,N_20332,N_20317);
or U20496 (N_20496,N_20364,N_20245);
xor U20497 (N_20497,N_20206,N_20302);
or U20498 (N_20498,N_20385,N_20294);
nand U20499 (N_20499,N_20300,N_20345);
and U20500 (N_20500,N_20287,N_20398);
and U20501 (N_20501,N_20365,N_20202);
xnor U20502 (N_20502,N_20209,N_20270);
or U20503 (N_20503,N_20259,N_20307);
and U20504 (N_20504,N_20355,N_20307);
and U20505 (N_20505,N_20244,N_20371);
nor U20506 (N_20506,N_20246,N_20325);
nand U20507 (N_20507,N_20255,N_20363);
xor U20508 (N_20508,N_20365,N_20269);
xor U20509 (N_20509,N_20231,N_20234);
and U20510 (N_20510,N_20215,N_20232);
and U20511 (N_20511,N_20398,N_20378);
nor U20512 (N_20512,N_20346,N_20288);
and U20513 (N_20513,N_20288,N_20255);
and U20514 (N_20514,N_20371,N_20383);
nor U20515 (N_20515,N_20343,N_20290);
xnor U20516 (N_20516,N_20329,N_20293);
and U20517 (N_20517,N_20248,N_20266);
nand U20518 (N_20518,N_20326,N_20370);
xor U20519 (N_20519,N_20354,N_20353);
nor U20520 (N_20520,N_20367,N_20232);
xor U20521 (N_20521,N_20288,N_20219);
nand U20522 (N_20522,N_20235,N_20386);
and U20523 (N_20523,N_20303,N_20260);
nor U20524 (N_20524,N_20318,N_20338);
nor U20525 (N_20525,N_20249,N_20266);
and U20526 (N_20526,N_20268,N_20294);
xor U20527 (N_20527,N_20256,N_20305);
or U20528 (N_20528,N_20287,N_20255);
or U20529 (N_20529,N_20253,N_20289);
nor U20530 (N_20530,N_20211,N_20284);
nand U20531 (N_20531,N_20257,N_20340);
or U20532 (N_20532,N_20293,N_20335);
and U20533 (N_20533,N_20318,N_20294);
or U20534 (N_20534,N_20261,N_20214);
or U20535 (N_20535,N_20244,N_20265);
xnor U20536 (N_20536,N_20265,N_20229);
xor U20537 (N_20537,N_20395,N_20222);
nand U20538 (N_20538,N_20296,N_20357);
or U20539 (N_20539,N_20277,N_20327);
nand U20540 (N_20540,N_20283,N_20365);
xor U20541 (N_20541,N_20295,N_20297);
and U20542 (N_20542,N_20265,N_20389);
xnor U20543 (N_20543,N_20226,N_20275);
and U20544 (N_20544,N_20330,N_20341);
or U20545 (N_20545,N_20271,N_20278);
nand U20546 (N_20546,N_20217,N_20319);
xnor U20547 (N_20547,N_20218,N_20390);
and U20548 (N_20548,N_20223,N_20278);
xnor U20549 (N_20549,N_20362,N_20379);
and U20550 (N_20550,N_20331,N_20208);
xor U20551 (N_20551,N_20316,N_20265);
xor U20552 (N_20552,N_20323,N_20362);
or U20553 (N_20553,N_20335,N_20232);
or U20554 (N_20554,N_20376,N_20287);
nor U20555 (N_20555,N_20318,N_20384);
or U20556 (N_20556,N_20349,N_20350);
nand U20557 (N_20557,N_20267,N_20225);
nor U20558 (N_20558,N_20296,N_20398);
and U20559 (N_20559,N_20263,N_20260);
nand U20560 (N_20560,N_20308,N_20372);
and U20561 (N_20561,N_20296,N_20378);
nor U20562 (N_20562,N_20282,N_20324);
or U20563 (N_20563,N_20294,N_20210);
nand U20564 (N_20564,N_20212,N_20388);
xor U20565 (N_20565,N_20247,N_20293);
and U20566 (N_20566,N_20395,N_20284);
xnor U20567 (N_20567,N_20257,N_20253);
xnor U20568 (N_20568,N_20313,N_20347);
nand U20569 (N_20569,N_20395,N_20378);
nand U20570 (N_20570,N_20304,N_20271);
nand U20571 (N_20571,N_20237,N_20208);
xnor U20572 (N_20572,N_20362,N_20394);
nor U20573 (N_20573,N_20280,N_20325);
xor U20574 (N_20574,N_20261,N_20288);
and U20575 (N_20575,N_20259,N_20295);
nor U20576 (N_20576,N_20333,N_20348);
and U20577 (N_20577,N_20332,N_20243);
nand U20578 (N_20578,N_20369,N_20286);
xnor U20579 (N_20579,N_20224,N_20337);
and U20580 (N_20580,N_20374,N_20260);
or U20581 (N_20581,N_20235,N_20281);
nor U20582 (N_20582,N_20346,N_20355);
xor U20583 (N_20583,N_20213,N_20383);
nand U20584 (N_20584,N_20369,N_20278);
and U20585 (N_20585,N_20207,N_20336);
or U20586 (N_20586,N_20397,N_20212);
and U20587 (N_20587,N_20281,N_20218);
nor U20588 (N_20588,N_20360,N_20305);
nand U20589 (N_20589,N_20390,N_20372);
nor U20590 (N_20590,N_20332,N_20212);
nor U20591 (N_20591,N_20215,N_20294);
nor U20592 (N_20592,N_20386,N_20307);
xnor U20593 (N_20593,N_20307,N_20237);
or U20594 (N_20594,N_20320,N_20281);
or U20595 (N_20595,N_20209,N_20263);
and U20596 (N_20596,N_20222,N_20340);
xnor U20597 (N_20597,N_20308,N_20262);
xnor U20598 (N_20598,N_20391,N_20213);
nor U20599 (N_20599,N_20391,N_20350);
and U20600 (N_20600,N_20549,N_20516);
nand U20601 (N_20601,N_20456,N_20567);
nor U20602 (N_20602,N_20490,N_20540);
xnor U20603 (N_20603,N_20588,N_20541);
xor U20604 (N_20604,N_20491,N_20446);
or U20605 (N_20605,N_20436,N_20468);
or U20606 (N_20606,N_20577,N_20508);
nand U20607 (N_20607,N_20521,N_20578);
nand U20608 (N_20608,N_20463,N_20496);
and U20609 (N_20609,N_20466,N_20592);
nand U20610 (N_20610,N_20504,N_20531);
xnor U20611 (N_20611,N_20507,N_20447);
or U20612 (N_20612,N_20492,N_20558);
and U20613 (N_20613,N_20520,N_20569);
nand U20614 (N_20614,N_20537,N_20429);
nand U20615 (N_20615,N_20559,N_20568);
xor U20616 (N_20616,N_20488,N_20554);
and U20617 (N_20617,N_20506,N_20511);
nor U20618 (N_20618,N_20421,N_20501);
xnor U20619 (N_20619,N_20406,N_20465);
xnor U20620 (N_20620,N_20582,N_20473);
nor U20621 (N_20621,N_20505,N_20597);
nand U20622 (N_20622,N_20533,N_20563);
or U20623 (N_20623,N_20530,N_20514);
and U20624 (N_20624,N_20437,N_20596);
or U20625 (N_20625,N_20418,N_20560);
and U20626 (N_20626,N_20518,N_20550);
xor U20627 (N_20627,N_20510,N_20551);
or U20628 (N_20628,N_20420,N_20599);
nand U20629 (N_20629,N_20556,N_20402);
and U20630 (N_20630,N_20425,N_20415);
or U20631 (N_20631,N_20509,N_20548);
or U20632 (N_20632,N_20442,N_20574);
nor U20633 (N_20633,N_20502,N_20528);
nand U20634 (N_20634,N_20562,N_20409);
nand U20635 (N_20635,N_20542,N_20566);
nand U20636 (N_20636,N_20552,N_20519);
xnor U20637 (N_20637,N_20433,N_20443);
or U20638 (N_20638,N_20479,N_20523);
and U20639 (N_20639,N_20480,N_20476);
or U20640 (N_20640,N_20590,N_20407);
and U20641 (N_20641,N_20464,N_20576);
or U20642 (N_20642,N_20401,N_20478);
xor U20643 (N_20643,N_20484,N_20474);
xor U20644 (N_20644,N_20424,N_20428);
nor U20645 (N_20645,N_20461,N_20595);
and U20646 (N_20646,N_20539,N_20494);
and U20647 (N_20647,N_20515,N_20543);
xnor U20648 (N_20648,N_20454,N_20585);
xnor U20649 (N_20649,N_20522,N_20482);
or U20650 (N_20650,N_20439,N_20512);
or U20651 (N_20651,N_20457,N_20580);
xnor U20652 (N_20652,N_20583,N_20513);
nor U20653 (N_20653,N_20547,N_20452);
nor U20654 (N_20654,N_20586,N_20544);
nand U20655 (N_20655,N_20458,N_20444);
nor U20656 (N_20656,N_20419,N_20411);
nor U20657 (N_20657,N_20410,N_20589);
and U20658 (N_20658,N_20427,N_20561);
or U20659 (N_20659,N_20404,N_20538);
and U20660 (N_20660,N_20405,N_20434);
nand U20661 (N_20661,N_20571,N_20467);
nand U20662 (N_20662,N_20498,N_20477);
or U20663 (N_20663,N_20573,N_20449);
nor U20664 (N_20664,N_20593,N_20412);
xnor U20665 (N_20665,N_20432,N_20536);
or U20666 (N_20666,N_20584,N_20471);
nand U20667 (N_20667,N_20435,N_20400);
xnor U20668 (N_20668,N_20553,N_20489);
and U20669 (N_20669,N_20526,N_20459);
xor U20670 (N_20670,N_20416,N_20546);
xor U20671 (N_20671,N_20534,N_20450);
and U20672 (N_20672,N_20564,N_20451);
and U20673 (N_20673,N_20487,N_20426);
nand U20674 (N_20674,N_20441,N_20598);
nand U20675 (N_20675,N_20493,N_20485);
or U20676 (N_20676,N_20403,N_20503);
nand U20677 (N_20677,N_20565,N_20408);
nand U20678 (N_20678,N_20413,N_20579);
xor U20679 (N_20679,N_20470,N_20499);
nand U20680 (N_20680,N_20453,N_20587);
nor U20681 (N_20681,N_20570,N_20472);
xor U20682 (N_20682,N_20438,N_20423);
and U20683 (N_20683,N_20555,N_20414);
or U20684 (N_20684,N_20529,N_20455);
nand U20685 (N_20685,N_20497,N_20445);
and U20686 (N_20686,N_20532,N_20431);
nand U20687 (N_20687,N_20481,N_20524);
nand U20688 (N_20688,N_20591,N_20517);
and U20689 (N_20689,N_20575,N_20495);
or U20690 (N_20690,N_20500,N_20545);
nor U20691 (N_20691,N_20422,N_20572);
nor U20692 (N_20692,N_20527,N_20462);
xnor U20693 (N_20693,N_20594,N_20486);
nand U20694 (N_20694,N_20417,N_20557);
or U20695 (N_20695,N_20525,N_20448);
nor U20696 (N_20696,N_20581,N_20430);
or U20697 (N_20697,N_20440,N_20460);
nand U20698 (N_20698,N_20483,N_20475);
and U20699 (N_20699,N_20469,N_20535);
and U20700 (N_20700,N_20445,N_20570);
nor U20701 (N_20701,N_20463,N_20448);
and U20702 (N_20702,N_20423,N_20552);
xor U20703 (N_20703,N_20490,N_20511);
nand U20704 (N_20704,N_20522,N_20523);
xnor U20705 (N_20705,N_20426,N_20509);
and U20706 (N_20706,N_20477,N_20443);
and U20707 (N_20707,N_20568,N_20470);
or U20708 (N_20708,N_20579,N_20586);
xnor U20709 (N_20709,N_20445,N_20486);
or U20710 (N_20710,N_20493,N_20556);
xor U20711 (N_20711,N_20584,N_20596);
nand U20712 (N_20712,N_20583,N_20481);
xor U20713 (N_20713,N_20531,N_20572);
xor U20714 (N_20714,N_20465,N_20538);
xor U20715 (N_20715,N_20417,N_20443);
nor U20716 (N_20716,N_20598,N_20565);
nor U20717 (N_20717,N_20451,N_20492);
xnor U20718 (N_20718,N_20446,N_20476);
nor U20719 (N_20719,N_20507,N_20413);
xor U20720 (N_20720,N_20571,N_20522);
nor U20721 (N_20721,N_20416,N_20539);
or U20722 (N_20722,N_20576,N_20557);
nand U20723 (N_20723,N_20478,N_20417);
nand U20724 (N_20724,N_20580,N_20514);
or U20725 (N_20725,N_20527,N_20497);
nand U20726 (N_20726,N_20514,N_20479);
or U20727 (N_20727,N_20420,N_20556);
or U20728 (N_20728,N_20472,N_20589);
nand U20729 (N_20729,N_20451,N_20580);
nand U20730 (N_20730,N_20569,N_20580);
or U20731 (N_20731,N_20415,N_20408);
xnor U20732 (N_20732,N_20530,N_20532);
or U20733 (N_20733,N_20520,N_20588);
nand U20734 (N_20734,N_20467,N_20426);
xnor U20735 (N_20735,N_20508,N_20521);
nand U20736 (N_20736,N_20483,N_20468);
or U20737 (N_20737,N_20527,N_20455);
or U20738 (N_20738,N_20493,N_20512);
xor U20739 (N_20739,N_20549,N_20566);
nor U20740 (N_20740,N_20560,N_20431);
or U20741 (N_20741,N_20529,N_20467);
nor U20742 (N_20742,N_20564,N_20486);
xor U20743 (N_20743,N_20594,N_20589);
or U20744 (N_20744,N_20519,N_20539);
nand U20745 (N_20745,N_20492,N_20546);
and U20746 (N_20746,N_20538,N_20578);
nor U20747 (N_20747,N_20517,N_20530);
nand U20748 (N_20748,N_20403,N_20449);
nor U20749 (N_20749,N_20474,N_20458);
and U20750 (N_20750,N_20501,N_20592);
nor U20751 (N_20751,N_20531,N_20474);
or U20752 (N_20752,N_20409,N_20596);
and U20753 (N_20753,N_20452,N_20448);
nand U20754 (N_20754,N_20554,N_20514);
or U20755 (N_20755,N_20506,N_20555);
nand U20756 (N_20756,N_20579,N_20518);
nor U20757 (N_20757,N_20579,N_20508);
xnor U20758 (N_20758,N_20426,N_20558);
nor U20759 (N_20759,N_20473,N_20455);
and U20760 (N_20760,N_20567,N_20436);
and U20761 (N_20761,N_20525,N_20450);
and U20762 (N_20762,N_20403,N_20571);
and U20763 (N_20763,N_20447,N_20432);
or U20764 (N_20764,N_20551,N_20429);
nand U20765 (N_20765,N_20478,N_20432);
or U20766 (N_20766,N_20466,N_20516);
and U20767 (N_20767,N_20548,N_20531);
or U20768 (N_20768,N_20457,N_20573);
nor U20769 (N_20769,N_20436,N_20426);
nand U20770 (N_20770,N_20518,N_20412);
nand U20771 (N_20771,N_20407,N_20431);
xnor U20772 (N_20772,N_20431,N_20505);
nand U20773 (N_20773,N_20440,N_20469);
xnor U20774 (N_20774,N_20597,N_20595);
xnor U20775 (N_20775,N_20420,N_20525);
or U20776 (N_20776,N_20442,N_20570);
nand U20777 (N_20777,N_20580,N_20564);
xnor U20778 (N_20778,N_20567,N_20574);
xor U20779 (N_20779,N_20496,N_20567);
or U20780 (N_20780,N_20596,N_20400);
or U20781 (N_20781,N_20476,N_20441);
and U20782 (N_20782,N_20586,N_20472);
and U20783 (N_20783,N_20466,N_20402);
nor U20784 (N_20784,N_20451,N_20568);
xnor U20785 (N_20785,N_20569,N_20404);
or U20786 (N_20786,N_20406,N_20573);
xnor U20787 (N_20787,N_20574,N_20400);
xor U20788 (N_20788,N_20582,N_20513);
nor U20789 (N_20789,N_20584,N_20489);
xor U20790 (N_20790,N_20489,N_20438);
xnor U20791 (N_20791,N_20451,N_20478);
or U20792 (N_20792,N_20519,N_20498);
nand U20793 (N_20793,N_20556,N_20592);
or U20794 (N_20794,N_20483,N_20423);
nor U20795 (N_20795,N_20430,N_20548);
or U20796 (N_20796,N_20407,N_20443);
nor U20797 (N_20797,N_20474,N_20425);
nand U20798 (N_20798,N_20570,N_20540);
and U20799 (N_20799,N_20526,N_20445);
nand U20800 (N_20800,N_20774,N_20630);
and U20801 (N_20801,N_20738,N_20748);
or U20802 (N_20802,N_20778,N_20792);
nor U20803 (N_20803,N_20698,N_20780);
or U20804 (N_20804,N_20604,N_20790);
nor U20805 (N_20805,N_20660,N_20740);
xnor U20806 (N_20806,N_20721,N_20672);
xnor U20807 (N_20807,N_20713,N_20677);
nor U20808 (N_20808,N_20763,N_20719);
xnor U20809 (N_20809,N_20741,N_20603);
or U20810 (N_20810,N_20701,N_20600);
and U20811 (N_20811,N_20707,N_20723);
nand U20812 (N_20812,N_20631,N_20728);
nand U20813 (N_20813,N_20687,N_20753);
and U20814 (N_20814,N_20773,N_20720);
and U20815 (N_20815,N_20644,N_20769);
xor U20816 (N_20816,N_20680,N_20796);
or U20817 (N_20817,N_20612,N_20781);
or U20818 (N_20818,N_20654,N_20619);
nor U20819 (N_20819,N_20626,N_20706);
nand U20820 (N_20820,N_20651,N_20730);
or U20821 (N_20821,N_20791,N_20695);
and U20822 (N_20822,N_20662,N_20611);
nand U20823 (N_20823,N_20647,N_20655);
and U20824 (N_20824,N_20751,N_20643);
or U20825 (N_20825,N_20637,N_20742);
or U20826 (N_20826,N_20733,N_20605);
or U20827 (N_20827,N_20788,N_20711);
nor U20828 (N_20828,N_20722,N_20666);
xor U20829 (N_20829,N_20640,N_20779);
nor U20830 (N_20830,N_20623,N_20610);
and U20831 (N_20831,N_20745,N_20732);
or U20832 (N_20832,N_20658,N_20767);
nor U20833 (N_20833,N_20601,N_20754);
nor U20834 (N_20834,N_20682,N_20777);
nor U20835 (N_20835,N_20709,N_20782);
nor U20836 (N_20836,N_20755,N_20608);
nand U20837 (N_20837,N_20775,N_20737);
xnor U20838 (N_20838,N_20629,N_20684);
nand U20839 (N_20839,N_20793,N_20614);
nor U20840 (N_20840,N_20727,N_20712);
or U20841 (N_20841,N_20699,N_20691);
nor U20842 (N_20842,N_20648,N_20636);
xnor U20843 (N_20843,N_20690,N_20679);
xnor U20844 (N_20844,N_20606,N_20764);
nor U20845 (N_20845,N_20661,N_20708);
and U20846 (N_20846,N_20659,N_20736);
or U20847 (N_20847,N_20752,N_20770);
nor U20848 (N_20848,N_20704,N_20726);
nor U20849 (N_20849,N_20671,N_20750);
or U20850 (N_20850,N_20725,N_20642);
nand U20851 (N_20851,N_20784,N_20797);
or U20852 (N_20852,N_20795,N_20625);
xor U20853 (N_20853,N_20632,N_20613);
and U20854 (N_20854,N_20670,N_20789);
and U20855 (N_20855,N_20760,N_20786);
nor U20856 (N_20856,N_20735,N_20743);
xor U20857 (N_20857,N_20765,N_20674);
xnor U20858 (N_20858,N_20710,N_20627);
xor U20859 (N_20859,N_20649,N_20676);
or U20860 (N_20860,N_20693,N_20705);
and U20861 (N_20861,N_20694,N_20634);
or U20862 (N_20862,N_20734,N_20729);
nand U20863 (N_20863,N_20717,N_20768);
or U20864 (N_20864,N_20602,N_20757);
and U20865 (N_20865,N_20669,N_20652);
or U20866 (N_20866,N_20697,N_20702);
xor U20867 (N_20867,N_20620,N_20696);
or U20868 (N_20868,N_20639,N_20618);
xnor U20869 (N_20869,N_20746,N_20749);
or U20870 (N_20870,N_20689,N_20656);
nand U20871 (N_20871,N_20759,N_20724);
or U20872 (N_20872,N_20714,N_20799);
xnor U20873 (N_20873,N_20641,N_20715);
nand U20874 (N_20874,N_20673,N_20664);
nand U20875 (N_20875,N_20667,N_20756);
and U20876 (N_20876,N_20758,N_20683);
or U20877 (N_20877,N_20615,N_20646);
and U20878 (N_20878,N_20616,N_20624);
nand U20879 (N_20879,N_20794,N_20787);
nor U20880 (N_20880,N_20650,N_20692);
xnor U20881 (N_20881,N_20703,N_20663);
xnor U20882 (N_20882,N_20716,N_20653);
or U20883 (N_20883,N_20783,N_20747);
nor U20884 (N_20884,N_20771,N_20686);
and U20885 (N_20885,N_20617,N_20668);
xor U20886 (N_20886,N_20638,N_20766);
or U20887 (N_20887,N_20622,N_20772);
and U20888 (N_20888,N_20681,N_20665);
xnor U20889 (N_20889,N_20762,N_20700);
nand U20890 (N_20890,N_20628,N_20609);
or U20891 (N_20891,N_20657,N_20675);
or U20892 (N_20892,N_20678,N_20798);
nor U20893 (N_20893,N_20635,N_20607);
and U20894 (N_20894,N_20645,N_20776);
or U20895 (N_20895,N_20739,N_20761);
or U20896 (N_20896,N_20688,N_20744);
nand U20897 (N_20897,N_20621,N_20718);
or U20898 (N_20898,N_20731,N_20785);
xor U20899 (N_20899,N_20633,N_20685);
nor U20900 (N_20900,N_20680,N_20631);
and U20901 (N_20901,N_20656,N_20729);
or U20902 (N_20902,N_20602,N_20660);
xor U20903 (N_20903,N_20665,N_20621);
nand U20904 (N_20904,N_20797,N_20667);
and U20905 (N_20905,N_20668,N_20670);
and U20906 (N_20906,N_20716,N_20678);
and U20907 (N_20907,N_20614,N_20739);
or U20908 (N_20908,N_20715,N_20658);
xor U20909 (N_20909,N_20756,N_20790);
nor U20910 (N_20910,N_20716,N_20715);
xor U20911 (N_20911,N_20708,N_20693);
or U20912 (N_20912,N_20753,N_20773);
xor U20913 (N_20913,N_20613,N_20628);
xor U20914 (N_20914,N_20711,N_20678);
or U20915 (N_20915,N_20779,N_20766);
or U20916 (N_20916,N_20768,N_20690);
and U20917 (N_20917,N_20705,N_20709);
and U20918 (N_20918,N_20720,N_20788);
and U20919 (N_20919,N_20682,N_20739);
nand U20920 (N_20920,N_20734,N_20794);
xnor U20921 (N_20921,N_20610,N_20725);
xnor U20922 (N_20922,N_20658,N_20769);
xnor U20923 (N_20923,N_20743,N_20611);
or U20924 (N_20924,N_20703,N_20769);
and U20925 (N_20925,N_20719,N_20620);
nor U20926 (N_20926,N_20744,N_20723);
or U20927 (N_20927,N_20697,N_20651);
nor U20928 (N_20928,N_20761,N_20693);
nand U20929 (N_20929,N_20645,N_20669);
nor U20930 (N_20930,N_20645,N_20770);
and U20931 (N_20931,N_20730,N_20727);
or U20932 (N_20932,N_20745,N_20663);
nand U20933 (N_20933,N_20748,N_20700);
or U20934 (N_20934,N_20622,N_20610);
nand U20935 (N_20935,N_20699,N_20636);
and U20936 (N_20936,N_20674,N_20685);
nor U20937 (N_20937,N_20679,N_20736);
xnor U20938 (N_20938,N_20757,N_20742);
nand U20939 (N_20939,N_20727,N_20626);
nor U20940 (N_20940,N_20747,N_20719);
nand U20941 (N_20941,N_20781,N_20652);
nor U20942 (N_20942,N_20710,N_20696);
and U20943 (N_20943,N_20792,N_20690);
nor U20944 (N_20944,N_20627,N_20743);
nand U20945 (N_20945,N_20796,N_20777);
xor U20946 (N_20946,N_20746,N_20600);
and U20947 (N_20947,N_20751,N_20634);
and U20948 (N_20948,N_20601,N_20771);
nand U20949 (N_20949,N_20693,N_20772);
nor U20950 (N_20950,N_20676,N_20710);
xor U20951 (N_20951,N_20668,N_20710);
nand U20952 (N_20952,N_20699,N_20733);
xor U20953 (N_20953,N_20671,N_20607);
and U20954 (N_20954,N_20750,N_20631);
and U20955 (N_20955,N_20733,N_20764);
xor U20956 (N_20956,N_20753,N_20617);
nand U20957 (N_20957,N_20607,N_20638);
or U20958 (N_20958,N_20773,N_20676);
nor U20959 (N_20959,N_20758,N_20749);
xnor U20960 (N_20960,N_20621,N_20722);
or U20961 (N_20961,N_20738,N_20756);
or U20962 (N_20962,N_20763,N_20693);
nor U20963 (N_20963,N_20791,N_20644);
and U20964 (N_20964,N_20766,N_20681);
and U20965 (N_20965,N_20744,N_20639);
nor U20966 (N_20966,N_20704,N_20619);
nand U20967 (N_20967,N_20649,N_20613);
xor U20968 (N_20968,N_20608,N_20708);
nand U20969 (N_20969,N_20657,N_20658);
nand U20970 (N_20970,N_20771,N_20626);
or U20971 (N_20971,N_20657,N_20622);
nand U20972 (N_20972,N_20779,N_20736);
or U20973 (N_20973,N_20684,N_20738);
or U20974 (N_20974,N_20694,N_20764);
or U20975 (N_20975,N_20761,N_20724);
or U20976 (N_20976,N_20787,N_20759);
or U20977 (N_20977,N_20772,N_20743);
xnor U20978 (N_20978,N_20602,N_20750);
and U20979 (N_20979,N_20724,N_20648);
nand U20980 (N_20980,N_20612,N_20777);
nand U20981 (N_20981,N_20777,N_20787);
and U20982 (N_20982,N_20702,N_20634);
or U20983 (N_20983,N_20746,N_20753);
and U20984 (N_20984,N_20727,N_20782);
nand U20985 (N_20985,N_20654,N_20739);
nor U20986 (N_20986,N_20630,N_20634);
nor U20987 (N_20987,N_20719,N_20706);
nor U20988 (N_20988,N_20743,N_20781);
xnor U20989 (N_20989,N_20611,N_20715);
and U20990 (N_20990,N_20771,N_20652);
nand U20991 (N_20991,N_20691,N_20632);
and U20992 (N_20992,N_20670,N_20722);
and U20993 (N_20993,N_20682,N_20625);
nand U20994 (N_20994,N_20655,N_20645);
nand U20995 (N_20995,N_20734,N_20755);
nand U20996 (N_20996,N_20705,N_20634);
and U20997 (N_20997,N_20727,N_20777);
or U20998 (N_20998,N_20649,N_20787);
xnor U20999 (N_20999,N_20768,N_20609);
nand U21000 (N_21000,N_20813,N_20965);
or U21001 (N_21001,N_20856,N_20968);
nand U21002 (N_21002,N_20928,N_20932);
nand U21003 (N_21003,N_20877,N_20936);
and U21004 (N_21004,N_20855,N_20830);
xor U21005 (N_21005,N_20970,N_20861);
xor U21006 (N_21006,N_20822,N_20801);
xor U21007 (N_21007,N_20890,N_20918);
nor U21008 (N_21008,N_20800,N_20922);
nand U21009 (N_21009,N_20899,N_20979);
nand U21010 (N_21010,N_20914,N_20852);
nand U21011 (N_21011,N_20943,N_20886);
or U21012 (N_21012,N_20872,N_20818);
or U21013 (N_21013,N_20986,N_20871);
nor U21014 (N_21014,N_20854,N_20876);
nand U21015 (N_21015,N_20901,N_20962);
or U21016 (N_21016,N_20878,N_20804);
nand U21017 (N_21017,N_20907,N_20860);
nand U21018 (N_21018,N_20926,N_20897);
xnor U21019 (N_21019,N_20933,N_20808);
nor U21020 (N_21020,N_20963,N_20823);
or U21021 (N_21021,N_20868,N_20863);
nor U21022 (N_21022,N_20880,N_20974);
nor U21023 (N_21023,N_20846,N_20882);
nor U21024 (N_21024,N_20848,N_20879);
nor U21025 (N_21025,N_20817,N_20973);
and U21026 (N_21026,N_20991,N_20840);
nor U21027 (N_21027,N_20850,N_20853);
xnor U21028 (N_21028,N_20833,N_20893);
or U21029 (N_21029,N_20838,N_20858);
or U21030 (N_21030,N_20917,N_20810);
and U21031 (N_21031,N_20946,N_20889);
nand U21032 (N_21032,N_20990,N_20807);
xor U21033 (N_21033,N_20997,N_20969);
xor U21034 (N_21034,N_20814,N_20908);
and U21035 (N_21035,N_20957,N_20951);
nor U21036 (N_21036,N_20919,N_20955);
and U21037 (N_21037,N_20819,N_20975);
xnor U21038 (N_21038,N_20966,N_20815);
xnor U21039 (N_21039,N_20865,N_20915);
nor U21040 (N_21040,N_20867,N_20942);
nand U21041 (N_21041,N_20811,N_20906);
and U21042 (N_21042,N_20869,N_20891);
nor U21043 (N_21043,N_20839,N_20836);
and U21044 (N_21044,N_20993,N_20845);
xor U21045 (N_21045,N_20925,N_20904);
nor U21046 (N_21046,N_20894,N_20842);
or U21047 (N_21047,N_20913,N_20900);
or U21048 (N_21048,N_20960,N_20859);
xnor U21049 (N_21049,N_20945,N_20809);
nand U21050 (N_21050,N_20950,N_20857);
and U21051 (N_21051,N_20977,N_20929);
nand U21052 (N_21052,N_20985,N_20939);
nand U21053 (N_21053,N_20829,N_20980);
xor U21054 (N_21054,N_20866,N_20989);
xnor U21055 (N_21055,N_20952,N_20982);
nor U21056 (N_21056,N_20949,N_20826);
nand U21057 (N_21057,N_20851,N_20916);
nor U21058 (N_21058,N_20972,N_20884);
and U21059 (N_21059,N_20964,N_20883);
and U21060 (N_21060,N_20837,N_20896);
and U21061 (N_21061,N_20930,N_20995);
and U21062 (N_21062,N_20983,N_20956);
nor U21063 (N_21063,N_20844,N_20958);
and U21064 (N_21064,N_20825,N_20988);
and U21065 (N_21065,N_20987,N_20940);
xor U21066 (N_21066,N_20967,N_20992);
nor U21067 (N_21067,N_20921,N_20862);
and U21068 (N_21068,N_20816,N_20948);
nand U21069 (N_21069,N_20805,N_20978);
or U21070 (N_21070,N_20938,N_20902);
or U21071 (N_21071,N_20953,N_20888);
or U21072 (N_21072,N_20976,N_20803);
xnor U21073 (N_21073,N_20887,N_20927);
nor U21074 (N_21074,N_20996,N_20944);
or U21075 (N_21075,N_20821,N_20935);
xnor U21076 (N_21076,N_20981,N_20834);
or U21077 (N_21077,N_20961,N_20920);
and U21078 (N_21078,N_20873,N_20831);
xnor U21079 (N_21079,N_20984,N_20954);
and U21080 (N_21080,N_20827,N_20937);
nor U21081 (N_21081,N_20895,N_20905);
and U21082 (N_21082,N_20998,N_20841);
and U21083 (N_21083,N_20832,N_20806);
or U21084 (N_21084,N_20849,N_20847);
xor U21085 (N_21085,N_20923,N_20885);
or U21086 (N_21086,N_20881,N_20874);
nor U21087 (N_21087,N_20802,N_20947);
and U21088 (N_21088,N_20843,N_20835);
and U21089 (N_21089,N_20934,N_20812);
nand U21090 (N_21090,N_20870,N_20910);
nand U21091 (N_21091,N_20903,N_20864);
or U21092 (N_21092,N_20999,N_20971);
xor U21093 (N_21093,N_20912,N_20959);
nand U21094 (N_21094,N_20898,N_20994);
nand U21095 (N_21095,N_20909,N_20820);
and U21096 (N_21096,N_20828,N_20931);
or U21097 (N_21097,N_20875,N_20941);
xnor U21098 (N_21098,N_20824,N_20892);
nand U21099 (N_21099,N_20911,N_20924);
and U21100 (N_21100,N_20906,N_20922);
or U21101 (N_21101,N_20973,N_20991);
nor U21102 (N_21102,N_20924,N_20898);
or U21103 (N_21103,N_20834,N_20986);
nand U21104 (N_21104,N_20975,N_20964);
xnor U21105 (N_21105,N_20820,N_20845);
nand U21106 (N_21106,N_20993,N_20913);
nor U21107 (N_21107,N_20922,N_20947);
and U21108 (N_21108,N_20971,N_20813);
nor U21109 (N_21109,N_20930,N_20981);
nor U21110 (N_21110,N_20853,N_20825);
nand U21111 (N_21111,N_20943,N_20983);
nor U21112 (N_21112,N_20930,N_20864);
and U21113 (N_21113,N_20976,N_20899);
or U21114 (N_21114,N_20853,N_20823);
nor U21115 (N_21115,N_20920,N_20986);
nand U21116 (N_21116,N_20801,N_20879);
xnor U21117 (N_21117,N_20807,N_20801);
and U21118 (N_21118,N_20893,N_20877);
nor U21119 (N_21119,N_20808,N_20968);
or U21120 (N_21120,N_20968,N_20938);
nor U21121 (N_21121,N_20956,N_20912);
nor U21122 (N_21122,N_20945,N_20991);
and U21123 (N_21123,N_20814,N_20823);
and U21124 (N_21124,N_20953,N_20962);
nor U21125 (N_21125,N_20936,N_20811);
xnor U21126 (N_21126,N_20835,N_20817);
xnor U21127 (N_21127,N_20894,N_20933);
and U21128 (N_21128,N_20902,N_20983);
or U21129 (N_21129,N_20990,N_20821);
or U21130 (N_21130,N_20982,N_20940);
nand U21131 (N_21131,N_20899,N_20804);
or U21132 (N_21132,N_20846,N_20913);
nor U21133 (N_21133,N_20955,N_20858);
xor U21134 (N_21134,N_20843,N_20943);
xor U21135 (N_21135,N_20898,N_20871);
nor U21136 (N_21136,N_20844,N_20977);
nor U21137 (N_21137,N_20874,N_20978);
or U21138 (N_21138,N_20973,N_20976);
or U21139 (N_21139,N_20807,N_20940);
and U21140 (N_21140,N_20885,N_20852);
nor U21141 (N_21141,N_20923,N_20994);
or U21142 (N_21142,N_20906,N_20920);
and U21143 (N_21143,N_20852,N_20825);
xnor U21144 (N_21144,N_20973,N_20895);
nor U21145 (N_21145,N_20907,N_20827);
nand U21146 (N_21146,N_20947,N_20941);
nor U21147 (N_21147,N_20987,N_20829);
nor U21148 (N_21148,N_20973,N_20864);
xnor U21149 (N_21149,N_20845,N_20858);
nand U21150 (N_21150,N_20920,N_20968);
nand U21151 (N_21151,N_20895,N_20814);
xnor U21152 (N_21152,N_20942,N_20906);
nand U21153 (N_21153,N_20909,N_20999);
or U21154 (N_21154,N_20859,N_20836);
xor U21155 (N_21155,N_20913,N_20825);
or U21156 (N_21156,N_20923,N_20997);
and U21157 (N_21157,N_20907,N_20868);
nand U21158 (N_21158,N_20867,N_20965);
and U21159 (N_21159,N_20869,N_20830);
and U21160 (N_21160,N_20939,N_20868);
nand U21161 (N_21161,N_20852,N_20906);
xor U21162 (N_21162,N_20918,N_20937);
xor U21163 (N_21163,N_20926,N_20841);
xor U21164 (N_21164,N_20955,N_20918);
and U21165 (N_21165,N_20869,N_20851);
nand U21166 (N_21166,N_20880,N_20857);
nand U21167 (N_21167,N_20851,N_20873);
nand U21168 (N_21168,N_20993,N_20958);
nor U21169 (N_21169,N_20892,N_20885);
nor U21170 (N_21170,N_20976,N_20883);
and U21171 (N_21171,N_20910,N_20936);
nor U21172 (N_21172,N_20862,N_20966);
nor U21173 (N_21173,N_20980,N_20867);
or U21174 (N_21174,N_20936,N_20849);
nand U21175 (N_21175,N_20870,N_20988);
nand U21176 (N_21176,N_20895,N_20949);
and U21177 (N_21177,N_20905,N_20827);
xnor U21178 (N_21178,N_20872,N_20912);
and U21179 (N_21179,N_20815,N_20804);
or U21180 (N_21180,N_20884,N_20881);
and U21181 (N_21181,N_20869,N_20957);
or U21182 (N_21182,N_20821,N_20844);
or U21183 (N_21183,N_20864,N_20871);
or U21184 (N_21184,N_20919,N_20802);
and U21185 (N_21185,N_20851,N_20806);
or U21186 (N_21186,N_20901,N_20879);
nor U21187 (N_21187,N_20932,N_20802);
nand U21188 (N_21188,N_20883,N_20867);
or U21189 (N_21189,N_20883,N_20960);
nor U21190 (N_21190,N_20816,N_20812);
nor U21191 (N_21191,N_20971,N_20926);
nor U21192 (N_21192,N_20889,N_20917);
nand U21193 (N_21193,N_20953,N_20845);
and U21194 (N_21194,N_20865,N_20972);
xor U21195 (N_21195,N_20909,N_20893);
xor U21196 (N_21196,N_20955,N_20887);
xnor U21197 (N_21197,N_20869,N_20801);
xor U21198 (N_21198,N_20954,N_20847);
and U21199 (N_21199,N_20861,N_20869);
or U21200 (N_21200,N_21007,N_21101);
nor U21201 (N_21201,N_21077,N_21061);
nand U21202 (N_21202,N_21185,N_21087);
and U21203 (N_21203,N_21191,N_21036);
and U21204 (N_21204,N_21066,N_21016);
or U21205 (N_21205,N_21162,N_21004);
nor U21206 (N_21206,N_21054,N_21058);
or U21207 (N_21207,N_21116,N_21002);
and U21208 (N_21208,N_21167,N_21117);
nand U21209 (N_21209,N_21031,N_21135);
xor U21210 (N_21210,N_21013,N_21043);
nand U21211 (N_21211,N_21086,N_21027);
and U21212 (N_21212,N_21063,N_21093);
nand U21213 (N_21213,N_21178,N_21045);
xnor U21214 (N_21214,N_21192,N_21049);
nor U21215 (N_21215,N_21080,N_21074);
nor U21216 (N_21216,N_21136,N_21060);
xnor U21217 (N_21217,N_21001,N_21173);
xnor U21218 (N_21218,N_21131,N_21181);
nor U21219 (N_21219,N_21003,N_21121);
and U21220 (N_21220,N_21120,N_21047);
nand U21221 (N_21221,N_21175,N_21000);
nand U21222 (N_21222,N_21183,N_21041);
xor U21223 (N_21223,N_21111,N_21008);
xor U21224 (N_21224,N_21194,N_21071);
nor U21225 (N_21225,N_21124,N_21062);
xnor U21226 (N_21226,N_21021,N_21102);
nor U21227 (N_21227,N_21127,N_21156);
xnor U21228 (N_21228,N_21046,N_21020);
nor U21229 (N_21229,N_21025,N_21174);
xnor U21230 (N_21230,N_21095,N_21105);
nor U21231 (N_21231,N_21139,N_21104);
xor U21232 (N_21232,N_21072,N_21079);
nor U21233 (N_21233,N_21017,N_21155);
and U21234 (N_21234,N_21166,N_21188);
nand U21235 (N_21235,N_21040,N_21195);
nand U21236 (N_21236,N_21033,N_21038);
and U21237 (N_21237,N_21048,N_21141);
and U21238 (N_21238,N_21164,N_21186);
and U21239 (N_21239,N_21085,N_21010);
xnor U21240 (N_21240,N_21112,N_21078);
nor U21241 (N_21241,N_21076,N_21106);
xor U21242 (N_21242,N_21052,N_21125);
nand U21243 (N_21243,N_21115,N_21152);
nand U21244 (N_21244,N_21184,N_21199);
nor U21245 (N_21245,N_21144,N_21159);
nand U21246 (N_21246,N_21015,N_21098);
xor U21247 (N_21247,N_21119,N_21196);
and U21248 (N_21248,N_21108,N_21073);
nand U21249 (N_21249,N_21107,N_21090);
xnor U21250 (N_21250,N_21147,N_21100);
nor U21251 (N_21251,N_21011,N_21037);
and U21252 (N_21252,N_21064,N_21146);
and U21253 (N_21253,N_21067,N_21172);
nor U21254 (N_21254,N_21158,N_21130);
or U21255 (N_21255,N_21182,N_21140);
or U21256 (N_21256,N_21059,N_21030);
or U21257 (N_21257,N_21154,N_21161);
nand U21258 (N_21258,N_21169,N_21193);
or U21259 (N_21259,N_21103,N_21143);
nand U21260 (N_21260,N_21133,N_21171);
or U21261 (N_21261,N_21065,N_21018);
or U21262 (N_21262,N_21042,N_21122);
xor U21263 (N_21263,N_21142,N_21006);
or U21264 (N_21264,N_21023,N_21170);
xor U21265 (N_21265,N_21082,N_21097);
or U21266 (N_21266,N_21089,N_21019);
xnor U21267 (N_21267,N_21138,N_21032);
nand U21268 (N_21268,N_21075,N_21110);
xnor U21269 (N_21269,N_21190,N_21150);
nand U21270 (N_21270,N_21134,N_21005);
and U21271 (N_21271,N_21092,N_21081);
or U21272 (N_21272,N_21024,N_21053);
nor U21273 (N_21273,N_21198,N_21176);
xor U21274 (N_21274,N_21022,N_21118);
nor U21275 (N_21275,N_21180,N_21070);
xor U21276 (N_21276,N_21114,N_21113);
and U21277 (N_21277,N_21160,N_21187);
nand U21278 (N_21278,N_21035,N_21109);
nor U21279 (N_21279,N_21157,N_21028);
and U21280 (N_21280,N_21039,N_21069);
nand U21281 (N_21281,N_21068,N_21163);
xor U21282 (N_21282,N_21148,N_21197);
and U21283 (N_21283,N_21050,N_21153);
and U21284 (N_21284,N_21132,N_21096);
xnor U21285 (N_21285,N_21034,N_21129);
nand U21286 (N_21286,N_21084,N_21137);
xor U21287 (N_21287,N_21128,N_21165);
xor U21288 (N_21288,N_21177,N_21055);
or U21289 (N_21289,N_21083,N_21051);
nand U21290 (N_21290,N_21014,N_21189);
or U21291 (N_21291,N_21009,N_21056);
nand U21292 (N_21292,N_21151,N_21012);
nand U21293 (N_21293,N_21099,N_21094);
xnor U21294 (N_21294,N_21179,N_21057);
and U21295 (N_21295,N_21091,N_21149);
nor U21296 (N_21296,N_21123,N_21088);
and U21297 (N_21297,N_21126,N_21044);
xor U21298 (N_21298,N_21168,N_21029);
xor U21299 (N_21299,N_21026,N_21145);
xor U21300 (N_21300,N_21122,N_21079);
nand U21301 (N_21301,N_21073,N_21179);
xnor U21302 (N_21302,N_21079,N_21041);
or U21303 (N_21303,N_21062,N_21147);
and U21304 (N_21304,N_21163,N_21034);
or U21305 (N_21305,N_21114,N_21025);
xnor U21306 (N_21306,N_21148,N_21150);
xor U21307 (N_21307,N_21124,N_21100);
xnor U21308 (N_21308,N_21080,N_21099);
nor U21309 (N_21309,N_21017,N_21149);
and U21310 (N_21310,N_21083,N_21187);
nor U21311 (N_21311,N_21078,N_21140);
and U21312 (N_21312,N_21075,N_21170);
nand U21313 (N_21313,N_21134,N_21060);
and U21314 (N_21314,N_21045,N_21153);
or U21315 (N_21315,N_21147,N_21178);
and U21316 (N_21316,N_21041,N_21086);
xnor U21317 (N_21317,N_21125,N_21162);
and U21318 (N_21318,N_21019,N_21152);
nand U21319 (N_21319,N_21021,N_21042);
xor U21320 (N_21320,N_21184,N_21123);
xnor U21321 (N_21321,N_21131,N_21064);
or U21322 (N_21322,N_21019,N_21106);
xnor U21323 (N_21323,N_21189,N_21061);
nand U21324 (N_21324,N_21161,N_21188);
nor U21325 (N_21325,N_21092,N_21190);
nor U21326 (N_21326,N_21191,N_21146);
and U21327 (N_21327,N_21094,N_21053);
xnor U21328 (N_21328,N_21076,N_21163);
and U21329 (N_21329,N_21151,N_21001);
and U21330 (N_21330,N_21159,N_21148);
xnor U21331 (N_21331,N_21138,N_21175);
and U21332 (N_21332,N_21045,N_21172);
or U21333 (N_21333,N_21161,N_21086);
or U21334 (N_21334,N_21090,N_21081);
or U21335 (N_21335,N_21199,N_21062);
or U21336 (N_21336,N_21131,N_21183);
xnor U21337 (N_21337,N_21163,N_21198);
nor U21338 (N_21338,N_21092,N_21083);
or U21339 (N_21339,N_21036,N_21182);
xnor U21340 (N_21340,N_21153,N_21106);
nand U21341 (N_21341,N_21161,N_21082);
and U21342 (N_21342,N_21177,N_21137);
nor U21343 (N_21343,N_21157,N_21036);
nor U21344 (N_21344,N_21155,N_21092);
nor U21345 (N_21345,N_21196,N_21013);
nand U21346 (N_21346,N_21125,N_21110);
and U21347 (N_21347,N_21147,N_21043);
xor U21348 (N_21348,N_21125,N_21146);
xor U21349 (N_21349,N_21132,N_21191);
or U21350 (N_21350,N_21130,N_21195);
xnor U21351 (N_21351,N_21068,N_21012);
or U21352 (N_21352,N_21049,N_21093);
nor U21353 (N_21353,N_21032,N_21149);
nand U21354 (N_21354,N_21031,N_21066);
or U21355 (N_21355,N_21113,N_21198);
or U21356 (N_21356,N_21102,N_21053);
and U21357 (N_21357,N_21140,N_21131);
nor U21358 (N_21358,N_21011,N_21149);
and U21359 (N_21359,N_21058,N_21070);
and U21360 (N_21360,N_21142,N_21183);
nand U21361 (N_21361,N_21174,N_21141);
nor U21362 (N_21362,N_21095,N_21052);
nand U21363 (N_21363,N_21057,N_21027);
nor U21364 (N_21364,N_21059,N_21099);
and U21365 (N_21365,N_21163,N_21061);
or U21366 (N_21366,N_21060,N_21180);
nor U21367 (N_21367,N_21171,N_21028);
and U21368 (N_21368,N_21074,N_21096);
and U21369 (N_21369,N_21031,N_21130);
xnor U21370 (N_21370,N_21032,N_21020);
and U21371 (N_21371,N_21006,N_21175);
xnor U21372 (N_21372,N_21063,N_21149);
xnor U21373 (N_21373,N_21003,N_21089);
xnor U21374 (N_21374,N_21024,N_21031);
nor U21375 (N_21375,N_21032,N_21037);
nand U21376 (N_21376,N_21042,N_21032);
nor U21377 (N_21377,N_21181,N_21029);
and U21378 (N_21378,N_21059,N_21027);
xor U21379 (N_21379,N_21192,N_21020);
and U21380 (N_21380,N_21066,N_21024);
nor U21381 (N_21381,N_21147,N_21086);
nor U21382 (N_21382,N_21009,N_21174);
nor U21383 (N_21383,N_21168,N_21103);
xor U21384 (N_21384,N_21062,N_21028);
nand U21385 (N_21385,N_21092,N_21116);
nand U21386 (N_21386,N_21041,N_21092);
and U21387 (N_21387,N_21006,N_21113);
nor U21388 (N_21388,N_21040,N_21143);
xor U21389 (N_21389,N_21018,N_21048);
xnor U21390 (N_21390,N_21146,N_21037);
or U21391 (N_21391,N_21197,N_21010);
and U21392 (N_21392,N_21079,N_21196);
nand U21393 (N_21393,N_21010,N_21189);
or U21394 (N_21394,N_21151,N_21106);
xor U21395 (N_21395,N_21010,N_21138);
xnor U21396 (N_21396,N_21177,N_21101);
or U21397 (N_21397,N_21155,N_21142);
or U21398 (N_21398,N_21129,N_21148);
or U21399 (N_21399,N_21180,N_21192);
nor U21400 (N_21400,N_21230,N_21357);
and U21401 (N_21401,N_21302,N_21385);
nand U21402 (N_21402,N_21296,N_21340);
xor U21403 (N_21403,N_21256,N_21352);
nand U21404 (N_21404,N_21323,N_21247);
nand U21405 (N_21405,N_21358,N_21396);
nor U21406 (N_21406,N_21374,N_21345);
nand U21407 (N_21407,N_21209,N_21367);
or U21408 (N_21408,N_21262,N_21238);
nand U21409 (N_21409,N_21382,N_21306);
and U21410 (N_21410,N_21378,N_21221);
and U21411 (N_21411,N_21332,N_21217);
nand U21412 (N_21412,N_21308,N_21285);
or U21413 (N_21413,N_21274,N_21204);
xor U21414 (N_21414,N_21369,N_21252);
and U21415 (N_21415,N_21389,N_21336);
or U21416 (N_21416,N_21213,N_21348);
xor U21417 (N_21417,N_21260,N_21318);
nand U21418 (N_21418,N_21282,N_21280);
nand U21419 (N_21419,N_21223,N_21360);
xnor U21420 (N_21420,N_21248,N_21351);
and U21421 (N_21421,N_21341,N_21354);
and U21422 (N_21422,N_21203,N_21328);
nand U21423 (N_21423,N_21355,N_21338);
or U21424 (N_21424,N_21244,N_21218);
or U21425 (N_21425,N_21215,N_21379);
nand U21426 (N_21426,N_21236,N_21245);
or U21427 (N_21427,N_21372,N_21392);
or U21428 (N_21428,N_21290,N_21224);
and U21429 (N_21429,N_21383,N_21258);
nand U21430 (N_21430,N_21210,N_21387);
nor U21431 (N_21431,N_21324,N_21349);
nor U21432 (N_21432,N_21225,N_21271);
nand U21433 (N_21433,N_21366,N_21362);
xor U21434 (N_21434,N_21309,N_21377);
xnor U21435 (N_21435,N_21370,N_21257);
or U21436 (N_21436,N_21263,N_21399);
nand U21437 (N_21437,N_21212,N_21319);
nor U21438 (N_21438,N_21266,N_21335);
nor U21439 (N_21439,N_21316,N_21286);
xnor U21440 (N_21440,N_21331,N_21222);
and U21441 (N_21441,N_21311,N_21297);
xnor U21442 (N_21442,N_21344,N_21391);
nand U21443 (N_21443,N_21314,N_21317);
or U21444 (N_21444,N_21350,N_21315);
xor U21445 (N_21445,N_21241,N_21291);
nand U21446 (N_21446,N_21220,N_21239);
and U21447 (N_21447,N_21246,N_21284);
and U21448 (N_21448,N_21243,N_21232);
and U21449 (N_21449,N_21205,N_21395);
xnor U21450 (N_21450,N_21333,N_21289);
nor U21451 (N_21451,N_21361,N_21254);
xnor U21452 (N_21452,N_21303,N_21216);
xnor U21453 (N_21453,N_21249,N_21278);
or U21454 (N_21454,N_21281,N_21277);
xnor U21455 (N_21455,N_21259,N_21321);
and U21456 (N_21456,N_21253,N_21270);
and U21457 (N_21457,N_21255,N_21330);
or U21458 (N_21458,N_21273,N_21214);
and U21459 (N_21459,N_21310,N_21265);
or U21460 (N_21460,N_21307,N_21343);
nand U21461 (N_21461,N_21211,N_21368);
nor U21462 (N_21462,N_21339,N_21279);
or U21463 (N_21463,N_21337,N_21287);
and U21464 (N_21464,N_21234,N_21342);
and U21465 (N_21465,N_21375,N_21272);
nand U21466 (N_21466,N_21201,N_21334);
nor U21467 (N_21467,N_21386,N_21398);
and U21468 (N_21468,N_21347,N_21276);
nand U21469 (N_21469,N_21329,N_21363);
and U21470 (N_21470,N_21295,N_21293);
or U21471 (N_21471,N_21288,N_21275);
or U21472 (N_21472,N_21390,N_21356);
nand U21473 (N_21473,N_21320,N_21300);
and U21474 (N_21474,N_21380,N_21219);
nand U21475 (N_21475,N_21235,N_21327);
or U21476 (N_21476,N_21207,N_21228);
nor U21477 (N_21477,N_21229,N_21283);
or U21478 (N_21478,N_21200,N_21299);
and U21479 (N_21479,N_21325,N_21226);
nand U21480 (N_21480,N_21326,N_21268);
and U21481 (N_21481,N_21346,N_21298);
nand U21482 (N_21482,N_21294,N_21364);
xor U21483 (N_21483,N_21371,N_21359);
nor U21484 (N_21484,N_21384,N_21381);
nor U21485 (N_21485,N_21240,N_21261);
nor U21486 (N_21486,N_21264,N_21242);
xnor U21487 (N_21487,N_21227,N_21304);
nand U21488 (N_21488,N_21388,N_21269);
or U21489 (N_21489,N_21208,N_21267);
nor U21490 (N_21490,N_21365,N_21231);
nand U21491 (N_21491,N_21376,N_21373);
xor U21492 (N_21492,N_21393,N_21394);
nor U21493 (N_21493,N_21305,N_21233);
nor U21494 (N_21494,N_21312,N_21313);
nor U21495 (N_21495,N_21251,N_21292);
nand U21496 (N_21496,N_21322,N_21237);
or U21497 (N_21497,N_21202,N_21250);
and U21498 (N_21498,N_21397,N_21206);
and U21499 (N_21499,N_21301,N_21353);
nor U21500 (N_21500,N_21294,N_21250);
or U21501 (N_21501,N_21395,N_21218);
xor U21502 (N_21502,N_21370,N_21296);
and U21503 (N_21503,N_21221,N_21298);
or U21504 (N_21504,N_21386,N_21263);
or U21505 (N_21505,N_21293,N_21344);
xnor U21506 (N_21506,N_21314,N_21217);
nand U21507 (N_21507,N_21255,N_21244);
nor U21508 (N_21508,N_21357,N_21343);
or U21509 (N_21509,N_21250,N_21314);
nor U21510 (N_21510,N_21258,N_21344);
xnor U21511 (N_21511,N_21209,N_21277);
xor U21512 (N_21512,N_21319,N_21362);
or U21513 (N_21513,N_21265,N_21228);
or U21514 (N_21514,N_21336,N_21343);
or U21515 (N_21515,N_21306,N_21295);
nor U21516 (N_21516,N_21265,N_21256);
nand U21517 (N_21517,N_21323,N_21244);
and U21518 (N_21518,N_21301,N_21317);
nor U21519 (N_21519,N_21361,N_21277);
and U21520 (N_21520,N_21346,N_21266);
xor U21521 (N_21521,N_21344,N_21353);
or U21522 (N_21522,N_21325,N_21383);
xnor U21523 (N_21523,N_21328,N_21229);
nor U21524 (N_21524,N_21304,N_21296);
nor U21525 (N_21525,N_21255,N_21316);
nand U21526 (N_21526,N_21394,N_21237);
or U21527 (N_21527,N_21381,N_21363);
nand U21528 (N_21528,N_21338,N_21330);
or U21529 (N_21529,N_21291,N_21250);
nand U21530 (N_21530,N_21299,N_21392);
or U21531 (N_21531,N_21263,N_21286);
nor U21532 (N_21532,N_21340,N_21294);
or U21533 (N_21533,N_21204,N_21363);
nor U21534 (N_21534,N_21214,N_21281);
or U21535 (N_21535,N_21273,N_21345);
and U21536 (N_21536,N_21341,N_21326);
nor U21537 (N_21537,N_21273,N_21283);
or U21538 (N_21538,N_21322,N_21228);
and U21539 (N_21539,N_21314,N_21340);
and U21540 (N_21540,N_21329,N_21299);
nand U21541 (N_21541,N_21258,N_21247);
nor U21542 (N_21542,N_21284,N_21268);
nor U21543 (N_21543,N_21206,N_21332);
nor U21544 (N_21544,N_21316,N_21370);
or U21545 (N_21545,N_21328,N_21339);
nand U21546 (N_21546,N_21218,N_21249);
or U21547 (N_21547,N_21206,N_21365);
xor U21548 (N_21548,N_21315,N_21326);
nor U21549 (N_21549,N_21278,N_21234);
nand U21550 (N_21550,N_21290,N_21365);
xor U21551 (N_21551,N_21374,N_21211);
nand U21552 (N_21552,N_21310,N_21359);
and U21553 (N_21553,N_21339,N_21316);
nand U21554 (N_21554,N_21231,N_21354);
nand U21555 (N_21555,N_21385,N_21206);
or U21556 (N_21556,N_21338,N_21249);
nor U21557 (N_21557,N_21259,N_21253);
nand U21558 (N_21558,N_21313,N_21249);
nand U21559 (N_21559,N_21235,N_21206);
nor U21560 (N_21560,N_21234,N_21275);
nor U21561 (N_21561,N_21271,N_21393);
nand U21562 (N_21562,N_21309,N_21275);
nand U21563 (N_21563,N_21205,N_21278);
nor U21564 (N_21564,N_21316,N_21384);
xor U21565 (N_21565,N_21285,N_21268);
and U21566 (N_21566,N_21263,N_21255);
nor U21567 (N_21567,N_21327,N_21304);
xor U21568 (N_21568,N_21271,N_21226);
and U21569 (N_21569,N_21339,N_21302);
nand U21570 (N_21570,N_21250,N_21345);
nand U21571 (N_21571,N_21391,N_21374);
and U21572 (N_21572,N_21324,N_21279);
nor U21573 (N_21573,N_21243,N_21220);
xnor U21574 (N_21574,N_21310,N_21309);
xor U21575 (N_21575,N_21343,N_21393);
nor U21576 (N_21576,N_21213,N_21229);
nand U21577 (N_21577,N_21357,N_21262);
xnor U21578 (N_21578,N_21394,N_21211);
nor U21579 (N_21579,N_21226,N_21322);
xnor U21580 (N_21580,N_21328,N_21288);
nor U21581 (N_21581,N_21331,N_21276);
xor U21582 (N_21582,N_21259,N_21390);
xor U21583 (N_21583,N_21367,N_21327);
xnor U21584 (N_21584,N_21348,N_21372);
xnor U21585 (N_21585,N_21340,N_21247);
xnor U21586 (N_21586,N_21281,N_21315);
nor U21587 (N_21587,N_21360,N_21378);
xor U21588 (N_21588,N_21217,N_21303);
nor U21589 (N_21589,N_21274,N_21224);
nor U21590 (N_21590,N_21228,N_21387);
nand U21591 (N_21591,N_21275,N_21266);
nand U21592 (N_21592,N_21298,N_21206);
nor U21593 (N_21593,N_21323,N_21274);
nand U21594 (N_21594,N_21371,N_21376);
and U21595 (N_21595,N_21241,N_21372);
and U21596 (N_21596,N_21329,N_21312);
nor U21597 (N_21597,N_21378,N_21384);
or U21598 (N_21598,N_21296,N_21242);
nor U21599 (N_21599,N_21279,N_21271);
or U21600 (N_21600,N_21487,N_21590);
or U21601 (N_21601,N_21557,N_21580);
and U21602 (N_21602,N_21473,N_21589);
or U21603 (N_21603,N_21509,N_21505);
nor U21604 (N_21604,N_21432,N_21442);
and U21605 (N_21605,N_21477,N_21591);
or U21606 (N_21606,N_21500,N_21458);
and U21607 (N_21607,N_21460,N_21485);
and U21608 (N_21608,N_21554,N_21585);
and U21609 (N_21609,N_21405,N_21549);
nor U21610 (N_21610,N_21437,N_21436);
nor U21611 (N_21611,N_21519,N_21444);
or U21612 (N_21612,N_21406,N_21561);
xnor U21613 (N_21613,N_21420,N_21467);
and U21614 (N_21614,N_21596,N_21546);
or U21615 (N_21615,N_21447,N_21451);
xor U21616 (N_21616,N_21572,N_21465);
or U21617 (N_21617,N_21412,N_21493);
nand U21618 (N_21618,N_21598,N_21403);
xor U21619 (N_21619,N_21512,N_21408);
xnor U21620 (N_21620,N_21494,N_21541);
nor U21621 (N_21621,N_21527,N_21441);
xor U21622 (N_21622,N_21479,N_21440);
nor U21623 (N_21623,N_21423,N_21491);
and U21624 (N_21624,N_21478,N_21503);
or U21625 (N_21625,N_21414,N_21461);
xor U21626 (N_21626,N_21559,N_21521);
xor U21627 (N_21627,N_21492,N_21449);
xnor U21628 (N_21628,N_21453,N_21525);
or U21629 (N_21629,N_21599,N_21537);
and U21630 (N_21630,N_21466,N_21552);
nand U21631 (N_21631,N_21535,N_21555);
and U21632 (N_21632,N_21484,N_21563);
nor U21633 (N_21633,N_21486,N_21568);
or U21634 (N_21634,N_21501,N_21578);
nand U21635 (N_21635,N_21518,N_21565);
nand U21636 (N_21636,N_21579,N_21566);
xnor U21637 (N_21637,N_21413,N_21513);
or U21638 (N_21638,N_21400,N_21439);
and U21639 (N_21639,N_21416,N_21488);
nand U21640 (N_21640,N_21564,N_21569);
and U21641 (N_21641,N_21475,N_21548);
nand U21642 (N_21642,N_21502,N_21480);
nor U21643 (N_21643,N_21415,N_21520);
nand U21644 (N_21644,N_21510,N_21404);
nand U21645 (N_21645,N_21407,N_21528);
and U21646 (N_21646,N_21504,N_21586);
or U21647 (N_21647,N_21529,N_21411);
or U21648 (N_21648,N_21402,N_21531);
nor U21649 (N_21649,N_21542,N_21551);
xnor U21650 (N_21650,N_21536,N_21417);
and U21651 (N_21651,N_21496,N_21524);
nor U21652 (N_21652,N_21592,N_21576);
and U21653 (N_21653,N_21421,N_21570);
nand U21654 (N_21654,N_21574,N_21553);
nor U21655 (N_21655,N_21545,N_21457);
nor U21656 (N_21656,N_21426,N_21588);
and U21657 (N_21657,N_21543,N_21489);
nand U21658 (N_21658,N_21560,N_21474);
or U21659 (N_21659,N_21468,N_21443);
and U21660 (N_21660,N_21435,N_21556);
nor U21661 (N_21661,N_21418,N_21401);
nor U21662 (N_21662,N_21470,N_21431);
or U21663 (N_21663,N_21446,N_21597);
or U21664 (N_21664,N_21425,N_21472);
nor U21665 (N_21665,N_21532,N_21511);
nor U21666 (N_21666,N_21539,N_21594);
nor U21667 (N_21667,N_21515,N_21595);
nand U21668 (N_21668,N_21583,N_21538);
or U21669 (N_21669,N_21409,N_21419);
and U21670 (N_21670,N_21498,N_21454);
or U21671 (N_21671,N_21448,N_21482);
xor U21672 (N_21672,N_21450,N_21438);
or U21673 (N_21673,N_21434,N_21582);
xor U21674 (N_21674,N_21464,N_21533);
xor U21675 (N_21675,N_21445,N_21573);
xor U21676 (N_21676,N_21540,N_21429);
or U21677 (N_21677,N_21483,N_21558);
and U21678 (N_21678,N_21490,N_21497);
nand U21679 (N_21679,N_21534,N_21526);
or U21680 (N_21680,N_21469,N_21508);
xnor U21681 (N_21681,N_21567,N_21463);
or U21682 (N_21682,N_21433,N_21581);
nor U21683 (N_21683,N_21517,N_21471);
nand U21684 (N_21684,N_21481,N_21495);
nor U21685 (N_21685,N_21452,N_21593);
nand U21686 (N_21686,N_21476,N_21427);
and U21687 (N_21687,N_21547,N_21530);
and U21688 (N_21688,N_21428,N_21455);
or U21689 (N_21689,N_21430,N_21575);
xnor U21690 (N_21690,N_21507,N_21584);
and U21691 (N_21691,N_21562,N_21577);
or U21692 (N_21692,N_21516,N_21459);
or U21693 (N_21693,N_21410,N_21424);
or U21694 (N_21694,N_21571,N_21550);
nand U21695 (N_21695,N_21587,N_21522);
nor U21696 (N_21696,N_21499,N_21456);
nor U21697 (N_21697,N_21422,N_21462);
xor U21698 (N_21698,N_21514,N_21544);
and U21699 (N_21699,N_21523,N_21506);
nand U21700 (N_21700,N_21401,N_21479);
xnor U21701 (N_21701,N_21487,N_21544);
xor U21702 (N_21702,N_21577,N_21440);
xor U21703 (N_21703,N_21451,N_21429);
or U21704 (N_21704,N_21594,N_21581);
nand U21705 (N_21705,N_21419,N_21564);
nor U21706 (N_21706,N_21585,N_21569);
and U21707 (N_21707,N_21547,N_21409);
nand U21708 (N_21708,N_21572,N_21540);
and U21709 (N_21709,N_21598,N_21507);
nand U21710 (N_21710,N_21426,N_21568);
nor U21711 (N_21711,N_21580,N_21523);
and U21712 (N_21712,N_21478,N_21406);
nand U21713 (N_21713,N_21500,N_21576);
nand U21714 (N_21714,N_21567,N_21556);
or U21715 (N_21715,N_21409,N_21453);
and U21716 (N_21716,N_21530,N_21569);
or U21717 (N_21717,N_21420,N_21502);
or U21718 (N_21718,N_21466,N_21589);
nand U21719 (N_21719,N_21443,N_21512);
xor U21720 (N_21720,N_21446,N_21423);
and U21721 (N_21721,N_21547,N_21485);
nor U21722 (N_21722,N_21551,N_21526);
nand U21723 (N_21723,N_21580,N_21463);
or U21724 (N_21724,N_21558,N_21515);
or U21725 (N_21725,N_21451,N_21521);
nand U21726 (N_21726,N_21543,N_21540);
nand U21727 (N_21727,N_21566,N_21580);
nand U21728 (N_21728,N_21404,N_21595);
nor U21729 (N_21729,N_21505,N_21515);
nand U21730 (N_21730,N_21575,N_21434);
nand U21731 (N_21731,N_21515,N_21589);
nor U21732 (N_21732,N_21477,N_21429);
or U21733 (N_21733,N_21458,N_21547);
or U21734 (N_21734,N_21596,N_21496);
xor U21735 (N_21735,N_21549,N_21439);
or U21736 (N_21736,N_21436,N_21475);
nor U21737 (N_21737,N_21427,N_21460);
xor U21738 (N_21738,N_21418,N_21554);
nand U21739 (N_21739,N_21507,N_21427);
nor U21740 (N_21740,N_21555,N_21442);
and U21741 (N_21741,N_21414,N_21469);
nand U21742 (N_21742,N_21581,N_21459);
and U21743 (N_21743,N_21590,N_21434);
nand U21744 (N_21744,N_21415,N_21411);
and U21745 (N_21745,N_21405,N_21406);
and U21746 (N_21746,N_21538,N_21400);
nand U21747 (N_21747,N_21459,N_21523);
xnor U21748 (N_21748,N_21542,N_21407);
or U21749 (N_21749,N_21445,N_21408);
nor U21750 (N_21750,N_21598,N_21556);
nor U21751 (N_21751,N_21500,N_21565);
and U21752 (N_21752,N_21402,N_21486);
nand U21753 (N_21753,N_21554,N_21529);
nor U21754 (N_21754,N_21526,N_21523);
xnor U21755 (N_21755,N_21441,N_21560);
and U21756 (N_21756,N_21455,N_21563);
and U21757 (N_21757,N_21532,N_21550);
nor U21758 (N_21758,N_21583,N_21410);
nand U21759 (N_21759,N_21487,N_21497);
nor U21760 (N_21760,N_21441,N_21422);
nor U21761 (N_21761,N_21471,N_21413);
nand U21762 (N_21762,N_21565,N_21507);
and U21763 (N_21763,N_21411,N_21461);
xnor U21764 (N_21764,N_21417,N_21457);
nand U21765 (N_21765,N_21507,N_21533);
nand U21766 (N_21766,N_21471,N_21511);
nand U21767 (N_21767,N_21465,N_21504);
or U21768 (N_21768,N_21578,N_21503);
xnor U21769 (N_21769,N_21470,N_21561);
xnor U21770 (N_21770,N_21486,N_21552);
and U21771 (N_21771,N_21523,N_21496);
or U21772 (N_21772,N_21553,N_21480);
xnor U21773 (N_21773,N_21496,N_21443);
and U21774 (N_21774,N_21565,N_21424);
nor U21775 (N_21775,N_21433,N_21424);
nor U21776 (N_21776,N_21599,N_21554);
nand U21777 (N_21777,N_21424,N_21507);
nor U21778 (N_21778,N_21577,N_21430);
or U21779 (N_21779,N_21472,N_21516);
xor U21780 (N_21780,N_21593,N_21472);
nand U21781 (N_21781,N_21415,N_21526);
or U21782 (N_21782,N_21564,N_21563);
xnor U21783 (N_21783,N_21529,N_21593);
or U21784 (N_21784,N_21493,N_21419);
nor U21785 (N_21785,N_21499,N_21536);
nand U21786 (N_21786,N_21578,N_21506);
and U21787 (N_21787,N_21593,N_21446);
nand U21788 (N_21788,N_21416,N_21452);
or U21789 (N_21789,N_21546,N_21526);
nor U21790 (N_21790,N_21416,N_21493);
xor U21791 (N_21791,N_21414,N_21596);
nor U21792 (N_21792,N_21578,N_21518);
xnor U21793 (N_21793,N_21428,N_21555);
and U21794 (N_21794,N_21517,N_21453);
xnor U21795 (N_21795,N_21513,N_21477);
nor U21796 (N_21796,N_21553,N_21587);
nor U21797 (N_21797,N_21485,N_21499);
xor U21798 (N_21798,N_21554,N_21504);
nor U21799 (N_21799,N_21456,N_21574);
nand U21800 (N_21800,N_21703,N_21671);
or U21801 (N_21801,N_21634,N_21739);
nor U21802 (N_21802,N_21669,N_21787);
nand U21803 (N_21803,N_21720,N_21636);
or U21804 (N_21804,N_21611,N_21777);
and U21805 (N_21805,N_21701,N_21735);
nor U21806 (N_21806,N_21738,N_21609);
nand U21807 (N_21807,N_21748,N_21689);
nand U21808 (N_21808,N_21608,N_21708);
xor U21809 (N_21809,N_21675,N_21640);
nand U21810 (N_21810,N_21688,N_21758);
nand U21811 (N_21811,N_21788,N_21616);
and U21812 (N_21812,N_21767,N_21681);
nor U21813 (N_21813,N_21657,N_21664);
nor U21814 (N_21814,N_21783,N_21755);
nor U21815 (N_21815,N_21638,N_21759);
or U21816 (N_21816,N_21668,N_21600);
and U21817 (N_21817,N_21679,N_21656);
xnor U21818 (N_21818,N_21621,N_21658);
nor U21819 (N_21819,N_21781,N_21606);
and U21820 (N_21820,N_21778,N_21713);
or U21821 (N_21821,N_21741,N_21762);
or U21822 (N_21822,N_21674,N_21729);
xnor U21823 (N_21823,N_21740,N_21722);
nand U21824 (N_21824,N_21717,N_21673);
xor U21825 (N_21825,N_21776,N_21624);
and U21826 (N_21826,N_21761,N_21644);
nand U21827 (N_21827,N_21628,N_21769);
and U21828 (N_21828,N_21766,N_21650);
nand U21829 (N_21829,N_21629,N_21682);
xor U21830 (N_21830,N_21604,N_21772);
or U21831 (N_21831,N_21775,N_21627);
xnor U21832 (N_21832,N_21709,N_21760);
and U21833 (N_21833,N_21715,N_21757);
and U21834 (N_21834,N_21641,N_21618);
and U21835 (N_21835,N_21710,N_21661);
and U21836 (N_21836,N_21645,N_21693);
nor U21837 (N_21837,N_21680,N_21737);
or U21838 (N_21838,N_21652,N_21770);
or U21839 (N_21839,N_21662,N_21605);
or U21840 (N_21840,N_21746,N_21793);
or U21841 (N_21841,N_21651,N_21718);
nand U21842 (N_21842,N_21734,N_21747);
or U21843 (N_21843,N_21780,N_21768);
nand U21844 (N_21844,N_21789,N_21716);
nand U21845 (N_21845,N_21602,N_21721);
nand U21846 (N_21846,N_21784,N_21691);
or U21847 (N_21847,N_21614,N_21617);
xor U21848 (N_21848,N_21779,N_21736);
and U21849 (N_21849,N_21782,N_21684);
nor U21850 (N_21850,N_21727,N_21712);
or U21851 (N_21851,N_21696,N_21786);
and U21852 (N_21852,N_21750,N_21795);
xor U21853 (N_21853,N_21765,N_21654);
xor U21854 (N_21854,N_21647,N_21764);
nand U21855 (N_21855,N_21763,N_21615);
nand U21856 (N_21856,N_21745,N_21714);
nand U21857 (N_21857,N_21601,N_21612);
nor U21858 (N_21858,N_21625,N_21702);
nand U21859 (N_21859,N_21631,N_21695);
xor U21860 (N_21860,N_21756,N_21633);
or U21861 (N_21861,N_21677,N_21791);
or U21862 (N_21862,N_21626,N_21683);
nor U21863 (N_21863,N_21620,N_21700);
nor U21864 (N_21864,N_21665,N_21667);
nand U21865 (N_21865,N_21676,N_21642);
nand U21866 (N_21866,N_21799,N_21666);
nand U21867 (N_21867,N_21610,N_21685);
nor U21868 (N_21868,N_21774,N_21706);
and U21869 (N_21869,N_21663,N_21632);
nor U21870 (N_21870,N_21649,N_21790);
xnor U21871 (N_21871,N_21711,N_21732);
nand U21872 (N_21872,N_21698,N_21607);
and U21873 (N_21873,N_21686,N_21687);
and U21874 (N_21874,N_21730,N_21655);
and U21875 (N_21875,N_21622,N_21692);
xnor U21876 (N_21876,N_21794,N_21660);
nand U21877 (N_21877,N_21653,N_21726);
and U21878 (N_21878,N_21613,N_21704);
or U21879 (N_21879,N_21743,N_21751);
and U21880 (N_21880,N_21672,N_21733);
or U21881 (N_21881,N_21643,N_21637);
nand U21882 (N_21882,N_21744,N_21773);
or U21883 (N_21883,N_21742,N_21719);
nand U21884 (N_21884,N_21731,N_21670);
xor U21885 (N_21885,N_21792,N_21648);
and U21886 (N_21886,N_21785,N_21771);
and U21887 (N_21887,N_21630,N_21725);
nor U21888 (N_21888,N_21646,N_21659);
or U21889 (N_21889,N_21723,N_21635);
nand U21890 (N_21890,N_21749,N_21690);
nor U21891 (N_21891,N_21796,N_21697);
xor U21892 (N_21892,N_21639,N_21678);
and U21893 (N_21893,N_21798,N_21724);
nand U21894 (N_21894,N_21754,N_21707);
or U21895 (N_21895,N_21619,N_21603);
xor U21896 (N_21896,N_21694,N_21797);
xnor U21897 (N_21897,N_21705,N_21623);
nand U21898 (N_21898,N_21752,N_21753);
nand U21899 (N_21899,N_21699,N_21728);
or U21900 (N_21900,N_21760,N_21665);
nand U21901 (N_21901,N_21684,N_21626);
xnor U21902 (N_21902,N_21667,N_21687);
and U21903 (N_21903,N_21668,N_21656);
xor U21904 (N_21904,N_21621,N_21635);
and U21905 (N_21905,N_21701,N_21676);
and U21906 (N_21906,N_21674,N_21771);
xnor U21907 (N_21907,N_21712,N_21759);
nor U21908 (N_21908,N_21608,N_21754);
nand U21909 (N_21909,N_21713,N_21643);
xor U21910 (N_21910,N_21669,N_21754);
and U21911 (N_21911,N_21603,N_21729);
nand U21912 (N_21912,N_21616,N_21623);
nor U21913 (N_21913,N_21724,N_21685);
or U21914 (N_21914,N_21602,N_21770);
nor U21915 (N_21915,N_21636,N_21614);
or U21916 (N_21916,N_21674,N_21645);
and U21917 (N_21917,N_21788,N_21766);
nand U21918 (N_21918,N_21772,N_21755);
xor U21919 (N_21919,N_21672,N_21649);
nand U21920 (N_21920,N_21733,N_21706);
nand U21921 (N_21921,N_21674,N_21735);
nand U21922 (N_21922,N_21705,N_21707);
nand U21923 (N_21923,N_21646,N_21685);
or U21924 (N_21924,N_21687,N_21704);
and U21925 (N_21925,N_21653,N_21797);
nand U21926 (N_21926,N_21642,N_21713);
or U21927 (N_21927,N_21778,N_21633);
xnor U21928 (N_21928,N_21629,N_21611);
nor U21929 (N_21929,N_21725,N_21758);
nor U21930 (N_21930,N_21729,N_21689);
nor U21931 (N_21931,N_21658,N_21646);
nor U21932 (N_21932,N_21636,N_21732);
or U21933 (N_21933,N_21701,N_21753);
and U21934 (N_21934,N_21693,N_21652);
nand U21935 (N_21935,N_21744,N_21619);
or U21936 (N_21936,N_21766,N_21742);
xor U21937 (N_21937,N_21601,N_21691);
or U21938 (N_21938,N_21789,N_21685);
or U21939 (N_21939,N_21712,N_21711);
xnor U21940 (N_21940,N_21648,N_21615);
nor U21941 (N_21941,N_21623,N_21663);
and U21942 (N_21942,N_21743,N_21740);
and U21943 (N_21943,N_21636,N_21792);
and U21944 (N_21944,N_21634,N_21732);
nor U21945 (N_21945,N_21624,N_21651);
or U21946 (N_21946,N_21690,N_21712);
or U21947 (N_21947,N_21681,N_21744);
or U21948 (N_21948,N_21747,N_21636);
xor U21949 (N_21949,N_21752,N_21778);
and U21950 (N_21950,N_21700,N_21793);
xnor U21951 (N_21951,N_21650,N_21667);
nor U21952 (N_21952,N_21758,N_21799);
nand U21953 (N_21953,N_21618,N_21736);
xor U21954 (N_21954,N_21667,N_21790);
nand U21955 (N_21955,N_21608,N_21630);
and U21956 (N_21956,N_21646,N_21757);
or U21957 (N_21957,N_21731,N_21782);
nand U21958 (N_21958,N_21754,N_21625);
nor U21959 (N_21959,N_21713,N_21727);
or U21960 (N_21960,N_21726,N_21640);
nand U21961 (N_21961,N_21603,N_21654);
nand U21962 (N_21962,N_21649,N_21674);
and U21963 (N_21963,N_21615,N_21613);
and U21964 (N_21964,N_21663,N_21620);
xor U21965 (N_21965,N_21781,N_21636);
and U21966 (N_21966,N_21644,N_21636);
xnor U21967 (N_21967,N_21631,N_21636);
nand U21968 (N_21968,N_21639,N_21660);
nand U21969 (N_21969,N_21724,N_21734);
nor U21970 (N_21970,N_21783,N_21732);
and U21971 (N_21971,N_21687,N_21614);
xor U21972 (N_21972,N_21726,N_21765);
or U21973 (N_21973,N_21692,N_21714);
nand U21974 (N_21974,N_21631,N_21646);
nor U21975 (N_21975,N_21781,N_21600);
nor U21976 (N_21976,N_21618,N_21749);
or U21977 (N_21977,N_21670,N_21684);
and U21978 (N_21978,N_21689,N_21780);
and U21979 (N_21979,N_21654,N_21633);
nor U21980 (N_21980,N_21799,N_21623);
xor U21981 (N_21981,N_21797,N_21758);
and U21982 (N_21982,N_21621,N_21796);
nor U21983 (N_21983,N_21755,N_21745);
or U21984 (N_21984,N_21739,N_21759);
or U21985 (N_21985,N_21782,N_21708);
nor U21986 (N_21986,N_21651,N_21748);
nand U21987 (N_21987,N_21684,N_21793);
xnor U21988 (N_21988,N_21791,N_21761);
or U21989 (N_21989,N_21703,N_21619);
or U21990 (N_21990,N_21632,N_21770);
xor U21991 (N_21991,N_21681,N_21615);
nand U21992 (N_21992,N_21644,N_21695);
or U21993 (N_21993,N_21667,N_21698);
xnor U21994 (N_21994,N_21655,N_21746);
or U21995 (N_21995,N_21651,N_21749);
nand U21996 (N_21996,N_21768,N_21690);
or U21997 (N_21997,N_21768,N_21702);
and U21998 (N_21998,N_21686,N_21742);
nand U21999 (N_21999,N_21667,N_21660);
nor U22000 (N_22000,N_21846,N_21867);
or U22001 (N_22001,N_21905,N_21976);
or U22002 (N_22002,N_21861,N_21904);
xnor U22003 (N_22003,N_21862,N_21851);
nand U22004 (N_22004,N_21860,N_21901);
nor U22005 (N_22005,N_21809,N_21962);
nor U22006 (N_22006,N_21898,N_21990);
and U22007 (N_22007,N_21813,N_21938);
xnor U22008 (N_22008,N_21810,N_21829);
and U22009 (N_22009,N_21893,N_21815);
nor U22010 (N_22010,N_21966,N_21805);
nand U22011 (N_22011,N_21839,N_21924);
nand U22012 (N_22012,N_21854,N_21800);
nand U22013 (N_22013,N_21832,N_21921);
nor U22014 (N_22014,N_21998,N_21896);
nand U22015 (N_22015,N_21947,N_21910);
nor U22016 (N_22016,N_21928,N_21926);
nand U22017 (N_22017,N_21817,N_21930);
and U22018 (N_22018,N_21961,N_21915);
xnor U22019 (N_22019,N_21963,N_21886);
nor U22020 (N_22020,N_21837,N_21881);
xnor U22021 (N_22021,N_21819,N_21918);
nand U22022 (N_22022,N_21876,N_21989);
and U22023 (N_22023,N_21820,N_21865);
or U22024 (N_22024,N_21909,N_21873);
and U22025 (N_22025,N_21841,N_21965);
nand U22026 (N_22026,N_21833,N_21954);
nand U22027 (N_22027,N_21945,N_21994);
nor U22028 (N_22028,N_21870,N_21834);
or U22029 (N_22029,N_21948,N_21955);
nand U22030 (N_22030,N_21978,N_21824);
nor U22031 (N_22031,N_21823,N_21911);
nand U22032 (N_22032,N_21987,N_21914);
or U22033 (N_22033,N_21892,N_21985);
xor U22034 (N_22034,N_21912,N_21874);
and U22035 (N_22035,N_21877,N_21825);
nor U22036 (N_22036,N_21887,N_21808);
and U22037 (N_22037,N_21864,N_21958);
nor U22038 (N_22038,N_21866,N_21888);
nor U22039 (N_22039,N_21925,N_21889);
xnor U22040 (N_22040,N_21803,N_21814);
and U22041 (N_22041,N_21879,N_21895);
nor U22042 (N_22042,N_21818,N_21953);
nand U22043 (N_22043,N_21806,N_21950);
nand U22044 (N_22044,N_21929,N_21845);
and U22045 (N_22045,N_21848,N_21807);
and U22046 (N_22046,N_21944,N_21986);
nand U22047 (N_22047,N_21849,N_21996);
nand U22048 (N_22048,N_21973,N_21847);
and U22049 (N_22049,N_21890,N_21974);
and U22050 (N_22050,N_21812,N_21967);
nor U22051 (N_22051,N_21875,N_21826);
and U22052 (N_22052,N_21844,N_21899);
xnor U22053 (N_22053,N_21964,N_21968);
nor U22054 (N_22054,N_21984,N_21852);
xnor U22055 (N_22055,N_21835,N_21997);
nor U22056 (N_22056,N_21941,N_21913);
nor U22057 (N_22057,N_21932,N_21983);
xnor U22058 (N_22058,N_21816,N_21802);
or U22059 (N_22059,N_21900,N_21894);
xnor U22060 (N_22060,N_21917,N_21882);
and U22061 (N_22061,N_21811,N_21871);
or U22062 (N_22062,N_21884,N_21858);
nor U22063 (N_22063,N_21916,N_21843);
xnor U22064 (N_22064,N_21878,N_21999);
nor U22065 (N_22065,N_21856,N_21920);
nor U22066 (N_22066,N_21949,N_21927);
and U22067 (N_22067,N_21972,N_21850);
xnor U22068 (N_22068,N_21922,N_21863);
xnor U22069 (N_22069,N_21934,N_21891);
xor U22070 (N_22070,N_21902,N_21946);
or U22071 (N_22071,N_21971,N_21988);
or U22072 (N_22072,N_21907,N_21933);
nand U22073 (N_22073,N_21992,N_21957);
or U22074 (N_22074,N_21956,N_21977);
nor U22075 (N_22075,N_21830,N_21980);
and U22076 (N_22076,N_21855,N_21991);
xor U22077 (N_22077,N_21943,N_21857);
nor U22078 (N_22078,N_21821,N_21936);
or U22079 (N_22079,N_21981,N_21801);
xnor U22080 (N_22080,N_21923,N_21868);
xor U22081 (N_22081,N_21908,N_21842);
nor U22082 (N_22082,N_21919,N_21869);
or U22083 (N_22083,N_21906,N_21838);
nand U22084 (N_22084,N_21880,N_21939);
or U22085 (N_22085,N_21804,N_21952);
and U22086 (N_22086,N_21897,N_21959);
xor U22087 (N_22087,N_21885,N_21995);
and U22088 (N_22088,N_21827,N_21883);
or U22089 (N_22089,N_21960,N_21872);
xnor U22090 (N_22090,N_21840,N_21853);
or U22091 (N_22091,N_21940,N_21951);
or U22092 (N_22092,N_21903,N_21831);
or U22093 (N_22093,N_21969,N_21937);
nor U22094 (N_22094,N_21982,N_21975);
or U22095 (N_22095,N_21931,N_21993);
xor U22096 (N_22096,N_21970,N_21859);
xor U22097 (N_22097,N_21979,N_21822);
nand U22098 (N_22098,N_21942,N_21935);
or U22099 (N_22099,N_21836,N_21828);
or U22100 (N_22100,N_21847,N_21980);
nor U22101 (N_22101,N_21997,N_21847);
xnor U22102 (N_22102,N_21939,N_21971);
nand U22103 (N_22103,N_21883,N_21860);
nor U22104 (N_22104,N_21946,N_21986);
and U22105 (N_22105,N_21857,N_21884);
nor U22106 (N_22106,N_21885,N_21836);
and U22107 (N_22107,N_21979,N_21836);
or U22108 (N_22108,N_21807,N_21953);
and U22109 (N_22109,N_21969,N_21872);
or U22110 (N_22110,N_21907,N_21949);
and U22111 (N_22111,N_21939,N_21817);
xnor U22112 (N_22112,N_21804,N_21852);
xnor U22113 (N_22113,N_21845,N_21994);
or U22114 (N_22114,N_21939,N_21864);
nand U22115 (N_22115,N_21829,N_21814);
nand U22116 (N_22116,N_21951,N_21962);
nand U22117 (N_22117,N_21906,N_21941);
nor U22118 (N_22118,N_21824,N_21947);
or U22119 (N_22119,N_21991,N_21826);
and U22120 (N_22120,N_21963,N_21991);
xor U22121 (N_22121,N_21928,N_21958);
xor U22122 (N_22122,N_21945,N_21923);
and U22123 (N_22123,N_21967,N_21992);
nor U22124 (N_22124,N_21804,N_21862);
xnor U22125 (N_22125,N_21933,N_21967);
xnor U22126 (N_22126,N_21832,N_21882);
nand U22127 (N_22127,N_21805,N_21819);
or U22128 (N_22128,N_21903,N_21917);
nand U22129 (N_22129,N_21879,N_21848);
or U22130 (N_22130,N_21983,N_21966);
nand U22131 (N_22131,N_21954,N_21848);
nand U22132 (N_22132,N_21908,N_21871);
nor U22133 (N_22133,N_21806,N_21931);
nand U22134 (N_22134,N_21838,N_21818);
xnor U22135 (N_22135,N_21883,N_21905);
nor U22136 (N_22136,N_21904,N_21913);
or U22137 (N_22137,N_21996,N_21824);
xnor U22138 (N_22138,N_21897,N_21812);
or U22139 (N_22139,N_21914,N_21842);
nand U22140 (N_22140,N_21925,N_21835);
or U22141 (N_22141,N_21930,N_21855);
and U22142 (N_22142,N_21831,N_21816);
nor U22143 (N_22143,N_21949,N_21818);
xnor U22144 (N_22144,N_21904,N_21821);
nor U22145 (N_22145,N_21973,N_21882);
nor U22146 (N_22146,N_21912,N_21826);
and U22147 (N_22147,N_21996,N_21884);
nor U22148 (N_22148,N_21971,N_21981);
nor U22149 (N_22149,N_21935,N_21831);
xor U22150 (N_22150,N_21915,N_21825);
or U22151 (N_22151,N_21842,N_21863);
and U22152 (N_22152,N_21889,N_21953);
and U22153 (N_22153,N_21962,N_21936);
or U22154 (N_22154,N_21826,N_21982);
nor U22155 (N_22155,N_21913,N_21922);
nand U22156 (N_22156,N_21837,N_21894);
or U22157 (N_22157,N_21829,N_21945);
or U22158 (N_22158,N_21976,N_21850);
and U22159 (N_22159,N_21885,N_21908);
or U22160 (N_22160,N_21835,N_21829);
xor U22161 (N_22161,N_21804,N_21939);
nand U22162 (N_22162,N_21904,N_21813);
xor U22163 (N_22163,N_21990,N_21876);
and U22164 (N_22164,N_21892,N_21925);
xor U22165 (N_22165,N_21802,N_21929);
xnor U22166 (N_22166,N_21860,N_21826);
and U22167 (N_22167,N_21892,N_21849);
or U22168 (N_22168,N_21887,N_21836);
or U22169 (N_22169,N_21833,N_21944);
xnor U22170 (N_22170,N_21911,N_21925);
and U22171 (N_22171,N_21989,N_21898);
nand U22172 (N_22172,N_21942,N_21939);
and U22173 (N_22173,N_21944,N_21822);
nor U22174 (N_22174,N_21902,N_21861);
nand U22175 (N_22175,N_21924,N_21905);
xnor U22176 (N_22176,N_21877,N_21925);
or U22177 (N_22177,N_21823,N_21832);
and U22178 (N_22178,N_21978,N_21829);
nand U22179 (N_22179,N_21892,N_21822);
nor U22180 (N_22180,N_21900,N_21860);
and U22181 (N_22181,N_21922,N_21931);
xnor U22182 (N_22182,N_21894,N_21893);
nor U22183 (N_22183,N_21995,N_21877);
nand U22184 (N_22184,N_21813,N_21817);
xor U22185 (N_22185,N_21953,N_21816);
or U22186 (N_22186,N_21926,N_21957);
and U22187 (N_22187,N_21884,N_21992);
nor U22188 (N_22188,N_21998,N_21959);
or U22189 (N_22189,N_21984,N_21897);
and U22190 (N_22190,N_21817,N_21982);
xor U22191 (N_22191,N_21810,N_21953);
nand U22192 (N_22192,N_21897,N_21886);
xor U22193 (N_22193,N_21871,N_21901);
or U22194 (N_22194,N_21808,N_21810);
xor U22195 (N_22195,N_21967,N_21883);
xor U22196 (N_22196,N_21903,N_21814);
or U22197 (N_22197,N_21952,N_21884);
or U22198 (N_22198,N_21801,N_21909);
or U22199 (N_22199,N_21813,N_21972);
or U22200 (N_22200,N_22198,N_22064);
nand U22201 (N_22201,N_22100,N_22154);
or U22202 (N_22202,N_22138,N_22150);
nor U22203 (N_22203,N_22188,N_22008);
or U22204 (N_22204,N_22136,N_22159);
nor U22205 (N_22205,N_22025,N_22019);
nand U22206 (N_22206,N_22003,N_22163);
xor U22207 (N_22207,N_22114,N_22185);
or U22208 (N_22208,N_22140,N_22023);
nand U22209 (N_22209,N_22101,N_22117);
nor U22210 (N_22210,N_22178,N_22009);
nand U22211 (N_22211,N_22021,N_22046);
xnor U22212 (N_22212,N_22134,N_22020);
and U22213 (N_22213,N_22062,N_22034);
nor U22214 (N_22214,N_22146,N_22190);
or U22215 (N_22215,N_22094,N_22036);
xor U22216 (N_22216,N_22093,N_22084);
and U22217 (N_22217,N_22180,N_22041);
or U22218 (N_22218,N_22016,N_22037);
nand U22219 (N_22219,N_22077,N_22014);
or U22220 (N_22220,N_22083,N_22080);
nor U22221 (N_22221,N_22032,N_22054);
nand U22222 (N_22222,N_22107,N_22106);
or U22223 (N_22223,N_22103,N_22112);
nor U22224 (N_22224,N_22119,N_22005);
and U22225 (N_22225,N_22113,N_22027);
nand U22226 (N_22226,N_22065,N_22174);
xor U22227 (N_22227,N_22011,N_22124);
or U22228 (N_22228,N_22142,N_22092);
and U22229 (N_22229,N_22081,N_22164);
xnor U22230 (N_22230,N_22066,N_22004);
xor U22231 (N_22231,N_22022,N_22177);
or U22232 (N_22232,N_22196,N_22049);
and U22233 (N_22233,N_22144,N_22076);
nor U22234 (N_22234,N_22038,N_22052);
and U22235 (N_22235,N_22125,N_22109);
and U22236 (N_22236,N_22123,N_22026);
or U22237 (N_22237,N_22090,N_22176);
nand U22238 (N_22238,N_22001,N_22017);
and U22239 (N_22239,N_22085,N_22051);
and U22240 (N_22240,N_22120,N_22089);
nor U22241 (N_22241,N_22193,N_22039);
or U22242 (N_22242,N_22153,N_22068);
or U22243 (N_22243,N_22195,N_22015);
and U22244 (N_22244,N_22096,N_22069);
xnor U22245 (N_22245,N_22116,N_22070);
nand U22246 (N_22246,N_22099,N_22098);
and U22247 (N_22247,N_22082,N_22168);
or U22248 (N_22248,N_22060,N_22013);
or U22249 (N_22249,N_22151,N_22104);
or U22250 (N_22250,N_22133,N_22149);
xnor U22251 (N_22251,N_22167,N_22139);
or U22252 (N_22252,N_22043,N_22007);
and U22253 (N_22253,N_22197,N_22157);
and U22254 (N_22254,N_22102,N_22111);
nand U22255 (N_22255,N_22179,N_22121);
xnor U22256 (N_22256,N_22187,N_22095);
nand U22257 (N_22257,N_22131,N_22061);
xor U22258 (N_22258,N_22192,N_22024);
or U22259 (N_22259,N_22172,N_22182);
nand U22260 (N_22260,N_22087,N_22028);
xnor U22261 (N_22261,N_22018,N_22000);
nor U22262 (N_22262,N_22170,N_22072);
and U22263 (N_22263,N_22067,N_22199);
xor U22264 (N_22264,N_22152,N_22128);
xnor U22265 (N_22265,N_22181,N_22126);
nor U22266 (N_22266,N_22002,N_22162);
nand U22267 (N_22267,N_22122,N_22115);
or U22268 (N_22268,N_22166,N_22097);
nor U22269 (N_22269,N_22074,N_22156);
xnor U22270 (N_22270,N_22044,N_22059);
or U22271 (N_22271,N_22029,N_22160);
xor U22272 (N_22272,N_22047,N_22141);
and U22273 (N_22273,N_22189,N_22183);
or U22274 (N_22274,N_22105,N_22048);
nor U22275 (N_22275,N_22071,N_22161);
nand U22276 (N_22276,N_22147,N_22035);
nor U22277 (N_22277,N_22063,N_22031);
or U22278 (N_22278,N_22173,N_22055);
nor U22279 (N_22279,N_22169,N_22135);
xnor U22280 (N_22280,N_22186,N_22132);
xor U22281 (N_22281,N_22030,N_22012);
and U22282 (N_22282,N_22108,N_22088);
xnor U22283 (N_22283,N_22075,N_22042);
nor U22284 (N_22284,N_22040,N_22086);
xor U22285 (N_22285,N_22078,N_22194);
and U22286 (N_22286,N_22184,N_22118);
nand U22287 (N_22287,N_22079,N_22053);
nor U22288 (N_22288,N_22127,N_22191);
nor U22289 (N_22289,N_22006,N_22175);
xor U22290 (N_22290,N_22137,N_22091);
or U22291 (N_22291,N_22045,N_22155);
and U22292 (N_22292,N_22148,N_22033);
or U22293 (N_22293,N_22130,N_22145);
xnor U22294 (N_22294,N_22143,N_22110);
xor U22295 (N_22295,N_22010,N_22050);
nand U22296 (N_22296,N_22158,N_22171);
xor U22297 (N_22297,N_22073,N_22057);
nand U22298 (N_22298,N_22056,N_22165);
nand U22299 (N_22299,N_22129,N_22058);
and U22300 (N_22300,N_22195,N_22131);
nand U22301 (N_22301,N_22034,N_22126);
nand U22302 (N_22302,N_22176,N_22140);
nand U22303 (N_22303,N_22187,N_22140);
xnor U22304 (N_22304,N_22040,N_22129);
or U22305 (N_22305,N_22180,N_22009);
or U22306 (N_22306,N_22156,N_22172);
xor U22307 (N_22307,N_22043,N_22175);
and U22308 (N_22308,N_22195,N_22170);
and U22309 (N_22309,N_22085,N_22168);
and U22310 (N_22310,N_22122,N_22153);
and U22311 (N_22311,N_22041,N_22003);
nor U22312 (N_22312,N_22062,N_22020);
or U22313 (N_22313,N_22158,N_22116);
nor U22314 (N_22314,N_22037,N_22143);
nand U22315 (N_22315,N_22097,N_22073);
and U22316 (N_22316,N_22134,N_22017);
nor U22317 (N_22317,N_22030,N_22144);
nand U22318 (N_22318,N_22192,N_22184);
nand U22319 (N_22319,N_22076,N_22048);
nor U22320 (N_22320,N_22177,N_22071);
and U22321 (N_22321,N_22092,N_22116);
nor U22322 (N_22322,N_22181,N_22044);
and U22323 (N_22323,N_22062,N_22124);
and U22324 (N_22324,N_22157,N_22101);
nand U22325 (N_22325,N_22158,N_22072);
xor U22326 (N_22326,N_22107,N_22145);
or U22327 (N_22327,N_22063,N_22078);
or U22328 (N_22328,N_22034,N_22050);
or U22329 (N_22329,N_22133,N_22004);
nor U22330 (N_22330,N_22099,N_22195);
nor U22331 (N_22331,N_22140,N_22035);
or U22332 (N_22332,N_22136,N_22199);
or U22333 (N_22333,N_22127,N_22181);
or U22334 (N_22334,N_22185,N_22095);
nor U22335 (N_22335,N_22194,N_22051);
xnor U22336 (N_22336,N_22009,N_22131);
xor U22337 (N_22337,N_22073,N_22159);
nor U22338 (N_22338,N_22032,N_22026);
nand U22339 (N_22339,N_22109,N_22011);
xor U22340 (N_22340,N_22120,N_22107);
and U22341 (N_22341,N_22151,N_22045);
xor U22342 (N_22342,N_22189,N_22065);
nand U22343 (N_22343,N_22187,N_22039);
and U22344 (N_22344,N_22188,N_22134);
nor U22345 (N_22345,N_22162,N_22122);
xor U22346 (N_22346,N_22123,N_22012);
and U22347 (N_22347,N_22177,N_22090);
nor U22348 (N_22348,N_22132,N_22011);
or U22349 (N_22349,N_22150,N_22099);
nand U22350 (N_22350,N_22106,N_22087);
or U22351 (N_22351,N_22173,N_22054);
and U22352 (N_22352,N_22009,N_22089);
nand U22353 (N_22353,N_22039,N_22006);
nor U22354 (N_22354,N_22177,N_22067);
or U22355 (N_22355,N_22129,N_22045);
or U22356 (N_22356,N_22031,N_22169);
and U22357 (N_22357,N_22060,N_22064);
or U22358 (N_22358,N_22179,N_22112);
xor U22359 (N_22359,N_22193,N_22057);
or U22360 (N_22360,N_22114,N_22165);
or U22361 (N_22361,N_22194,N_22186);
xor U22362 (N_22362,N_22171,N_22152);
xor U22363 (N_22363,N_22133,N_22090);
and U22364 (N_22364,N_22041,N_22191);
or U22365 (N_22365,N_22124,N_22146);
or U22366 (N_22366,N_22173,N_22019);
or U22367 (N_22367,N_22008,N_22030);
nand U22368 (N_22368,N_22099,N_22096);
nand U22369 (N_22369,N_22025,N_22038);
or U22370 (N_22370,N_22097,N_22107);
xor U22371 (N_22371,N_22059,N_22090);
xor U22372 (N_22372,N_22164,N_22177);
or U22373 (N_22373,N_22043,N_22160);
or U22374 (N_22374,N_22097,N_22164);
nor U22375 (N_22375,N_22149,N_22126);
nand U22376 (N_22376,N_22013,N_22108);
or U22377 (N_22377,N_22191,N_22182);
and U22378 (N_22378,N_22028,N_22098);
nand U22379 (N_22379,N_22174,N_22151);
and U22380 (N_22380,N_22188,N_22129);
or U22381 (N_22381,N_22126,N_22169);
and U22382 (N_22382,N_22149,N_22127);
nor U22383 (N_22383,N_22029,N_22164);
and U22384 (N_22384,N_22019,N_22002);
and U22385 (N_22385,N_22168,N_22170);
xor U22386 (N_22386,N_22002,N_22023);
xnor U22387 (N_22387,N_22051,N_22163);
and U22388 (N_22388,N_22133,N_22068);
and U22389 (N_22389,N_22038,N_22015);
and U22390 (N_22390,N_22089,N_22131);
nand U22391 (N_22391,N_22076,N_22107);
nor U22392 (N_22392,N_22070,N_22055);
xnor U22393 (N_22393,N_22039,N_22023);
nor U22394 (N_22394,N_22136,N_22055);
or U22395 (N_22395,N_22133,N_22143);
or U22396 (N_22396,N_22117,N_22066);
nand U22397 (N_22397,N_22008,N_22173);
and U22398 (N_22398,N_22017,N_22142);
and U22399 (N_22399,N_22103,N_22079);
nand U22400 (N_22400,N_22322,N_22229);
nand U22401 (N_22401,N_22397,N_22273);
or U22402 (N_22402,N_22280,N_22227);
nand U22403 (N_22403,N_22374,N_22344);
or U22404 (N_22404,N_22303,N_22350);
nand U22405 (N_22405,N_22380,N_22204);
or U22406 (N_22406,N_22217,N_22315);
xor U22407 (N_22407,N_22275,N_22352);
nand U22408 (N_22408,N_22267,N_22333);
nor U22409 (N_22409,N_22294,N_22336);
nor U22410 (N_22410,N_22258,N_22393);
nand U22411 (N_22411,N_22238,N_22289);
xor U22412 (N_22412,N_22246,N_22292);
nor U22413 (N_22413,N_22335,N_22376);
and U22414 (N_22414,N_22203,N_22327);
nor U22415 (N_22415,N_22243,N_22394);
or U22416 (N_22416,N_22291,N_22373);
nor U22417 (N_22417,N_22363,N_22339);
or U22418 (N_22418,N_22228,N_22210);
and U22419 (N_22419,N_22237,N_22240);
or U22420 (N_22420,N_22247,N_22316);
xnor U22421 (N_22421,N_22221,N_22390);
or U22422 (N_22422,N_22392,N_22357);
nand U22423 (N_22423,N_22331,N_22297);
or U22424 (N_22424,N_22284,N_22313);
and U22425 (N_22425,N_22306,N_22272);
nand U22426 (N_22426,N_22356,N_22268);
and U22427 (N_22427,N_22220,N_22319);
nand U22428 (N_22428,N_22251,N_22388);
nor U22429 (N_22429,N_22330,N_22399);
xnor U22430 (N_22430,N_22208,N_22296);
or U22431 (N_22431,N_22353,N_22219);
nand U22432 (N_22432,N_22355,N_22385);
nand U22433 (N_22433,N_22255,N_22269);
or U22434 (N_22434,N_22307,N_22354);
nor U22435 (N_22435,N_22371,N_22233);
xnor U22436 (N_22436,N_22293,N_22326);
or U22437 (N_22437,N_22288,N_22398);
nor U22438 (N_22438,N_22245,N_22285);
xnor U22439 (N_22439,N_22351,N_22372);
xnor U22440 (N_22440,N_22301,N_22278);
or U22441 (N_22441,N_22231,N_22370);
nand U22442 (N_22442,N_22279,N_22264);
and U22443 (N_22443,N_22320,N_22378);
xor U22444 (N_22444,N_22348,N_22349);
nand U22445 (N_22445,N_22311,N_22260);
and U22446 (N_22446,N_22256,N_22235);
nand U22447 (N_22447,N_22242,N_22310);
or U22448 (N_22448,N_22299,N_22214);
nor U22449 (N_22449,N_22290,N_22334);
and U22450 (N_22450,N_22286,N_22274);
xor U22451 (N_22451,N_22263,N_22276);
nor U22452 (N_22452,N_22257,N_22324);
nand U22453 (N_22453,N_22250,N_22224);
and U22454 (N_22454,N_22328,N_22211);
or U22455 (N_22455,N_22207,N_22265);
xnor U22456 (N_22456,N_22359,N_22200);
and U22457 (N_22457,N_22241,N_22384);
and U22458 (N_22458,N_22360,N_22343);
nor U22459 (N_22459,N_22345,N_22283);
nand U22460 (N_22460,N_22261,N_22342);
nand U22461 (N_22461,N_22216,N_22318);
or U22462 (N_22462,N_22239,N_22358);
or U22463 (N_22463,N_22387,N_22340);
or U22464 (N_22464,N_22361,N_22201);
or U22465 (N_22465,N_22332,N_22300);
and U22466 (N_22466,N_22212,N_22375);
nand U22467 (N_22467,N_22341,N_22386);
xor U22468 (N_22468,N_22308,N_22329);
nand U22469 (N_22469,N_22277,N_22314);
or U22470 (N_22470,N_22254,N_22321);
nor U22471 (N_22471,N_22266,N_22362);
nand U22472 (N_22472,N_22298,N_22395);
nor U22473 (N_22473,N_22396,N_22312);
xnor U22474 (N_22474,N_22337,N_22262);
or U22475 (N_22475,N_22236,N_22367);
or U22476 (N_22476,N_22215,N_22249);
nor U22477 (N_22477,N_22305,N_22347);
or U22478 (N_22478,N_22377,N_22205);
nor U22479 (N_22479,N_22381,N_22202);
nand U22480 (N_22480,N_22244,N_22209);
and U22481 (N_22481,N_22281,N_22234);
nand U22482 (N_22482,N_22223,N_22287);
xor U22483 (N_22483,N_22325,N_22225);
xnor U22484 (N_22484,N_22304,N_22346);
nor U22485 (N_22485,N_22338,N_22379);
nand U22486 (N_22486,N_22232,N_22368);
nand U22487 (N_22487,N_22248,N_22366);
and U22488 (N_22488,N_22213,N_22230);
or U22489 (N_22489,N_22364,N_22252);
nor U22490 (N_22490,N_22222,N_22218);
or U22491 (N_22491,N_22365,N_22389);
and U22492 (N_22492,N_22295,N_22271);
or U22493 (N_22493,N_22382,N_22253);
or U22494 (N_22494,N_22309,N_22323);
xnor U22495 (N_22495,N_22259,N_22270);
and U22496 (N_22496,N_22369,N_22282);
xor U22497 (N_22497,N_22317,N_22302);
or U22498 (N_22498,N_22226,N_22383);
nor U22499 (N_22499,N_22206,N_22391);
or U22500 (N_22500,N_22251,N_22296);
nor U22501 (N_22501,N_22363,N_22253);
xnor U22502 (N_22502,N_22329,N_22324);
nor U22503 (N_22503,N_22395,N_22396);
nor U22504 (N_22504,N_22251,N_22249);
nand U22505 (N_22505,N_22311,N_22343);
or U22506 (N_22506,N_22391,N_22280);
xor U22507 (N_22507,N_22298,N_22246);
nor U22508 (N_22508,N_22283,N_22355);
nor U22509 (N_22509,N_22308,N_22305);
nor U22510 (N_22510,N_22254,N_22226);
nor U22511 (N_22511,N_22384,N_22274);
or U22512 (N_22512,N_22276,N_22248);
xnor U22513 (N_22513,N_22216,N_22204);
or U22514 (N_22514,N_22350,N_22309);
or U22515 (N_22515,N_22245,N_22291);
xor U22516 (N_22516,N_22379,N_22252);
nand U22517 (N_22517,N_22399,N_22398);
xor U22518 (N_22518,N_22292,N_22384);
nor U22519 (N_22519,N_22261,N_22330);
or U22520 (N_22520,N_22333,N_22266);
xor U22521 (N_22521,N_22223,N_22234);
and U22522 (N_22522,N_22242,N_22318);
and U22523 (N_22523,N_22339,N_22224);
and U22524 (N_22524,N_22254,N_22340);
nor U22525 (N_22525,N_22387,N_22373);
and U22526 (N_22526,N_22226,N_22347);
and U22527 (N_22527,N_22223,N_22264);
and U22528 (N_22528,N_22267,N_22202);
nor U22529 (N_22529,N_22244,N_22223);
and U22530 (N_22530,N_22357,N_22263);
or U22531 (N_22531,N_22222,N_22344);
and U22532 (N_22532,N_22268,N_22335);
nor U22533 (N_22533,N_22386,N_22397);
and U22534 (N_22534,N_22278,N_22281);
and U22535 (N_22535,N_22215,N_22273);
or U22536 (N_22536,N_22362,N_22228);
nand U22537 (N_22537,N_22302,N_22375);
nor U22538 (N_22538,N_22361,N_22378);
or U22539 (N_22539,N_22370,N_22279);
nor U22540 (N_22540,N_22330,N_22300);
xor U22541 (N_22541,N_22245,N_22326);
nor U22542 (N_22542,N_22375,N_22360);
nor U22543 (N_22543,N_22232,N_22303);
or U22544 (N_22544,N_22397,N_22389);
nor U22545 (N_22545,N_22336,N_22295);
nand U22546 (N_22546,N_22336,N_22219);
nand U22547 (N_22547,N_22363,N_22278);
and U22548 (N_22548,N_22316,N_22351);
xnor U22549 (N_22549,N_22309,N_22291);
nor U22550 (N_22550,N_22365,N_22210);
and U22551 (N_22551,N_22375,N_22210);
xnor U22552 (N_22552,N_22210,N_22231);
and U22553 (N_22553,N_22343,N_22348);
nor U22554 (N_22554,N_22358,N_22352);
or U22555 (N_22555,N_22250,N_22256);
or U22556 (N_22556,N_22289,N_22210);
nor U22557 (N_22557,N_22304,N_22317);
or U22558 (N_22558,N_22325,N_22290);
nand U22559 (N_22559,N_22344,N_22303);
and U22560 (N_22560,N_22386,N_22339);
and U22561 (N_22561,N_22227,N_22391);
nand U22562 (N_22562,N_22356,N_22254);
xor U22563 (N_22563,N_22207,N_22244);
or U22564 (N_22564,N_22315,N_22386);
nand U22565 (N_22565,N_22204,N_22359);
xor U22566 (N_22566,N_22375,N_22259);
nand U22567 (N_22567,N_22273,N_22292);
or U22568 (N_22568,N_22267,N_22343);
and U22569 (N_22569,N_22338,N_22335);
and U22570 (N_22570,N_22382,N_22293);
xnor U22571 (N_22571,N_22246,N_22252);
nand U22572 (N_22572,N_22353,N_22252);
and U22573 (N_22573,N_22298,N_22214);
nand U22574 (N_22574,N_22309,N_22318);
nor U22575 (N_22575,N_22286,N_22334);
xnor U22576 (N_22576,N_22273,N_22256);
nand U22577 (N_22577,N_22277,N_22378);
or U22578 (N_22578,N_22326,N_22307);
xor U22579 (N_22579,N_22357,N_22376);
xor U22580 (N_22580,N_22264,N_22306);
and U22581 (N_22581,N_22233,N_22243);
nor U22582 (N_22582,N_22239,N_22359);
and U22583 (N_22583,N_22251,N_22373);
or U22584 (N_22584,N_22359,N_22365);
nor U22585 (N_22585,N_22374,N_22305);
nor U22586 (N_22586,N_22288,N_22324);
or U22587 (N_22587,N_22226,N_22202);
or U22588 (N_22588,N_22384,N_22297);
nor U22589 (N_22589,N_22257,N_22329);
nand U22590 (N_22590,N_22252,N_22291);
xnor U22591 (N_22591,N_22288,N_22370);
nand U22592 (N_22592,N_22343,N_22320);
or U22593 (N_22593,N_22344,N_22279);
xor U22594 (N_22594,N_22259,N_22248);
and U22595 (N_22595,N_22298,N_22230);
or U22596 (N_22596,N_22270,N_22380);
and U22597 (N_22597,N_22217,N_22292);
or U22598 (N_22598,N_22231,N_22394);
nand U22599 (N_22599,N_22395,N_22227);
or U22600 (N_22600,N_22597,N_22552);
nor U22601 (N_22601,N_22540,N_22558);
nor U22602 (N_22602,N_22588,N_22577);
and U22603 (N_22603,N_22579,N_22551);
or U22604 (N_22604,N_22440,N_22562);
nand U22605 (N_22605,N_22449,N_22481);
nand U22606 (N_22606,N_22477,N_22598);
and U22607 (N_22607,N_22575,N_22414);
xor U22608 (N_22608,N_22549,N_22409);
nor U22609 (N_22609,N_22569,N_22479);
xnor U22610 (N_22610,N_22595,N_22469);
or U22611 (N_22611,N_22430,N_22590);
xor U22612 (N_22612,N_22524,N_22559);
or U22613 (N_22613,N_22416,N_22423);
xor U22614 (N_22614,N_22410,N_22435);
xor U22615 (N_22615,N_22487,N_22442);
nor U22616 (N_22616,N_22534,N_22537);
and U22617 (N_22617,N_22528,N_22420);
xnor U22618 (N_22618,N_22408,N_22424);
nand U22619 (N_22619,N_22523,N_22581);
xnor U22620 (N_22620,N_22454,N_22494);
and U22621 (N_22621,N_22436,N_22403);
nor U22622 (N_22622,N_22421,N_22531);
nand U22623 (N_22623,N_22473,N_22448);
and U22624 (N_22624,N_22413,N_22464);
nor U22625 (N_22625,N_22571,N_22517);
xnor U22626 (N_22626,N_22536,N_22434);
nand U22627 (N_22627,N_22483,N_22596);
nand U22628 (N_22628,N_22428,N_22505);
or U22629 (N_22629,N_22492,N_22520);
xor U22630 (N_22630,N_22583,N_22554);
nand U22631 (N_22631,N_22488,N_22411);
nor U22632 (N_22632,N_22507,N_22500);
or U22633 (N_22633,N_22498,N_22418);
and U22634 (N_22634,N_22580,N_22548);
or U22635 (N_22635,N_22412,N_22450);
nand U22636 (N_22636,N_22446,N_22496);
xnor U22637 (N_22637,N_22422,N_22586);
xor U22638 (N_22638,N_22429,N_22576);
or U22639 (N_22639,N_22566,N_22453);
xor U22640 (N_22640,N_22400,N_22417);
and U22641 (N_22641,N_22478,N_22447);
nand U22642 (N_22642,N_22485,N_22555);
nor U22643 (N_22643,N_22510,N_22427);
nor U22644 (N_22644,N_22516,N_22437);
nand U22645 (N_22645,N_22545,N_22574);
xor U22646 (N_22646,N_22565,N_22511);
or U22647 (N_22647,N_22512,N_22521);
nor U22648 (N_22648,N_22425,N_22539);
and U22649 (N_22649,N_22508,N_22543);
xnor U22650 (N_22650,N_22438,N_22444);
and U22651 (N_22651,N_22570,N_22567);
and U22652 (N_22652,N_22402,N_22513);
xor U22653 (N_22653,N_22405,N_22572);
and U22654 (N_22654,N_22461,N_22544);
nor U22655 (N_22655,N_22530,N_22529);
or U22656 (N_22656,N_22443,N_22484);
nand U22657 (N_22657,N_22406,N_22546);
xor U22658 (N_22658,N_22470,N_22527);
and U22659 (N_22659,N_22573,N_22568);
nor U22660 (N_22660,N_22467,N_22538);
xnor U22661 (N_22661,N_22495,N_22578);
nand U22662 (N_22662,N_22491,N_22457);
xnor U22663 (N_22663,N_22587,N_22582);
or U22664 (N_22664,N_22564,N_22493);
or U22665 (N_22665,N_22504,N_22415);
and U22666 (N_22666,N_22592,N_22466);
and U22667 (N_22667,N_22455,N_22525);
or U22668 (N_22668,N_22419,N_22499);
nor U22669 (N_22669,N_22584,N_22541);
nor U22670 (N_22670,N_22433,N_22475);
and U22671 (N_22671,N_22452,N_22471);
and U22672 (N_22672,N_22533,N_22490);
and U22673 (N_22673,N_22593,N_22515);
and U22674 (N_22674,N_22439,N_22514);
and U22675 (N_22675,N_22456,N_22476);
and U22676 (N_22676,N_22480,N_22441);
and U22677 (N_22677,N_22458,N_22426);
and U22678 (N_22678,N_22503,N_22445);
nor U22679 (N_22679,N_22553,N_22465);
nor U22680 (N_22680,N_22459,N_22519);
nor U22681 (N_22681,N_22451,N_22472);
nand U22682 (N_22682,N_22526,N_22557);
and U22683 (N_22683,N_22497,N_22506);
xor U22684 (N_22684,N_22486,N_22509);
or U22685 (N_22685,N_22502,N_22585);
nand U22686 (N_22686,N_22463,N_22431);
and U22687 (N_22687,N_22401,N_22594);
nor U22688 (N_22688,N_22560,N_22563);
or U22689 (N_22689,N_22589,N_22535);
or U22690 (N_22690,N_22561,N_22432);
nand U22691 (N_22691,N_22550,N_22591);
nor U22692 (N_22692,N_22462,N_22482);
xnor U22693 (N_22693,N_22532,N_22501);
and U22694 (N_22694,N_22468,N_22522);
or U22695 (N_22695,N_22460,N_22556);
and U22696 (N_22696,N_22542,N_22547);
nor U22697 (N_22697,N_22404,N_22474);
nor U22698 (N_22698,N_22518,N_22489);
xor U22699 (N_22699,N_22599,N_22407);
nor U22700 (N_22700,N_22467,N_22409);
nand U22701 (N_22701,N_22551,N_22545);
and U22702 (N_22702,N_22551,N_22412);
xor U22703 (N_22703,N_22495,N_22512);
xnor U22704 (N_22704,N_22438,N_22548);
or U22705 (N_22705,N_22404,N_22448);
or U22706 (N_22706,N_22515,N_22548);
nand U22707 (N_22707,N_22455,N_22417);
xnor U22708 (N_22708,N_22536,N_22545);
nor U22709 (N_22709,N_22529,N_22558);
xnor U22710 (N_22710,N_22465,N_22474);
xor U22711 (N_22711,N_22415,N_22400);
xor U22712 (N_22712,N_22435,N_22427);
or U22713 (N_22713,N_22433,N_22502);
and U22714 (N_22714,N_22542,N_22465);
nor U22715 (N_22715,N_22496,N_22495);
and U22716 (N_22716,N_22443,N_22532);
and U22717 (N_22717,N_22582,N_22522);
and U22718 (N_22718,N_22454,N_22511);
or U22719 (N_22719,N_22437,N_22513);
nand U22720 (N_22720,N_22581,N_22445);
xor U22721 (N_22721,N_22462,N_22518);
or U22722 (N_22722,N_22565,N_22424);
nor U22723 (N_22723,N_22575,N_22526);
and U22724 (N_22724,N_22430,N_22526);
xor U22725 (N_22725,N_22567,N_22589);
or U22726 (N_22726,N_22506,N_22450);
nand U22727 (N_22727,N_22485,N_22508);
nand U22728 (N_22728,N_22540,N_22440);
or U22729 (N_22729,N_22473,N_22465);
nor U22730 (N_22730,N_22541,N_22525);
and U22731 (N_22731,N_22487,N_22457);
nand U22732 (N_22732,N_22508,N_22476);
and U22733 (N_22733,N_22456,N_22440);
or U22734 (N_22734,N_22539,N_22418);
and U22735 (N_22735,N_22453,N_22549);
or U22736 (N_22736,N_22504,N_22575);
or U22737 (N_22737,N_22536,N_22476);
nand U22738 (N_22738,N_22409,N_22559);
nor U22739 (N_22739,N_22407,N_22531);
or U22740 (N_22740,N_22552,N_22464);
nor U22741 (N_22741,N_22523,N_22566);
nor U22742 (N_22742,N_22557,N_22451);
and U22743 (N_22743,N_22493,N_22561);
and U22744 (N_22744,N_22589,N_22592);
xnor U22745 (N_22745,N_22425,N_22583);
or U22746 (N_22746,N_22515,N_22465);
xor U22747 (N_22747,N_22555,N_22508);
nor U22748 (N_22748,N_22471,N_22570);
nand U22749 (N_22749,N_22566,N_22559);
nand U22750 (N_22750,N_22599,N_22538);
xnor U22751 (N_22751,N_22449,N_22466);
nand U22752 (N_22752,N_22582,N_22527);
nand U22753 (N_22753,N_22531,N_22525);
nor U22754 (N_22754,N_22515,N_22504);
and U22755 (N_22755,N_22558,N_22582);
xnor U22756 (N_22756,N_22402,N_22563);
or U22757 (N_22757,N_22571,N_22531);
or U22758 (N_22758,N_22463,N_22454);
nor U22759 (N_22759,N_22507,N_22542);
and U22760 (N_22760,N_22442,N_22432);
or U22761 (N_22761,N_22483,N_22528);
nor U22762 (N_22762,N_22432,N_22466);
nor U22763 (N_22763,N_22459,N_22480);
nor U22764 (N_22764,N_22469,N_22496);
or U22765 (N_22765,N_22585,N_22433);
nand U22766 (N_22766,N_22494,N_22469);
nor U22767 (N_22767,N_22538,N_22539);
nor U22768 (N_22768,N_22450,N_22474);
or U22769 (N_22769,N_22428,N_22450);
xnor U22770 (N_22770,N_22479,N_22561);
or U22771 (N_22771,N_22564,N_22413);
nor U22772 (N_22772,N_22472,N_22573);
nand U22773 (N_22773,N_22558,N_22481);
and U22774 (N_22774,N_22539,N_22567);
or U22775 (N_22775,N_22416,N_22528);
nor U22776 (N_22776,N_22556,N_22458);
and U22777 (N_22777,N_22507,N_22414);
or U22778 (N_22778,N_22538,N_22508);
nand U22779 (N_22779,N_22589,N_22517);
xor U22780 (N_22780,N_22576,N_22475);
xor U22781 (N_22781,N_22527,N_22528);
or U22782 (N_22782,N_22406,N_22505);
and U22783 (N_22783,N_22576,N_22526);
or U22784 (N_22784,N_22576,N_22556);
nand U22785 (N_22785,N_22547,N_22411);
or U22786 (N_22786,N_22401,N_22557);
xor U22787 (N_22787,N_22513,N_22450);
nor U22788 (N_22788,N_22501,N_22426);
nor U22789 (N_22789,N_22474,N_22487);
and U22790 (N_22790,N_22434,N_22484);
nand U22791 (N_22791,N_22583,N_22586);
xor U22792 (N_22792,N_22479,N_22566);
or U22793 (N_22793,N_22487,N_22435);
xnor U22794 (N_22794,N_22545,N_22582);
xor U22795 (N_22795,N_22462,N_22411);
and U22796 (N_22796,N_22553,N_22560);
nand U22797 (N_22797,N_22433,N_22529);
xnor U22798 (N_22798,N_22479,N_22439);
and U22799 (N_22799,N_22437,N_22404);
nor U22800 (N_22800,N_22688,N_22627);
nor U22801 (N_22801,N_22685,N_22790);
and U22802 (N_22802,N_22705,N_22743);
or U22803 (N_22803,N_22799,N_22714);
or U22804 (N_22804,N_22777,N_22640);
and U22805 (N_22805,N_22711,N_22626);
nand U22806 (N_22806,N_22652,N_22762);
and U22807 (N_22807,N_22655,N_22718);
and U22808 (N_22808,N_22701,N_22794);
nor U22809 (N_22809,N_22796,N_22621);
or U22810 (N_22810,N_22614,N_22611);
nand U22811 (N_22811,N_22648,N_22600);
nor U22812 (N_22812,N_22618,N_22740);
or U22813 (N_22813,N_22749,N_22689);
or U22814 (N_22814,N_22663,N_22695);
xnor U22815 (N_22815,N_22662,N_22677);
nor U22816 (N_22816,N_22620,N_22769);
or U22817 (N_22817,N_22725,N_22671);
nor U22818 (N_22818,N_22742,N_22696);
or U22819 (N_22819,N_22724,N_22673);
or U22820 (N_22820,N_22754,N_22690);
and U22821 (N_22821,N_22780,N_22734);
nand U22822 (N_22822,N_22751,N_22793);
or U22823 (N_22823,N_22782,N_22722);
xnor U22824 (N_22824,N_22646,N_22676);
nor U22825 (N_22825,N_22656,N_22721);
xor U22826 (N_22826,N_22694,N_22739);
nand U22827 (N_22827,N_22612,N_22710);
nand U22828 (N_22828,N_22736,N_22700);
and U22829 (N_22829,N_22792,N_22798);
and U22830 (N_22830,N_22659,N_22608);
or U22831 (N_22831,N_22687,N_22767);
and U22832 (N_22832,N_22791,N_22766);
xor U22833 (N_22833,N_22670,N_22678);
and U22834 (N_22834,N_22669,N_22660);
and U22835 (N_22835,N_22649,N_22738);
nand U22836 (N_22836,N_22747,N_22619);
nor U22837 (N_22837,N_22760,N_22604);
nand U22838 (N_22838,N_22682,N_22729);
xnor U22839 (N_22839,N_22759,N_22771);
xnor U22840 (N_22840,N_22756,N_22753);
or U22841 (N_22841,N_22787,N_22757);
xor U22842 (N_22842,N_22651,N_22784);
or U22843 (N_22843,N_22776,N_22768);
nor U22844 (N_22844,N_22664,N_22707);
nand U22845 (N_22845,N_22622,N_22709);
xor U22846 (N_22846,N_22720,N_22698);
or U22847 (N_22847,N_22786,N_22723);
nand U22848 (N_22848,N_22672,N_22746);
and U22849 (N_22849,N_22726,N_22617);
and U22850 (N_22850,N_22629,N_22775);
nand U22851 (N_22851,N_22772,N_22602);
or U22852 (N_22852,N_22650,N_22623);
nor U22853 (N_22853,N_22636,N_22732);
xor U22854 (N_22854,N_22624,N_22630);
nor U22855 (N_22855,N_22758,N_22713);
xor U22856 (N_22856,N_22783,N_22763);
nand U22857 (N_22857,N_22642,N_22702);
or U22858 (N_22858,N_22715,N_22765);
or U22859 (N_22859,N_22633,N_22730);
nand U22860 (N_22860,N_22657,N_22727);
or U22861 (N_22861,N_22628,N_22631);
nor U22862 (N_22862,N_22748,N_22741);
or U22863 (N_22863,N_22615,N_22643);
nor U22864 (N_22864,N_22789,N_22750);
nor U22865 (N_22865,N_22733,N_22691);
nand U22866 (N_22866,N_22745,N_22717);
xnor U22867 (N_22867,N_22609,N_22667);
nor U22868 (N_22868,N_22781,N_22704);
nand U22869 (N_22869,N_22675,N_22634);
nand U22870 (N_22870,N_22605,N_22697);
nor U22871 (N_22871,N_22637,N_22606);
nand U22872 (N_22872,N_22641,N_22683);
nor U22873 (N_22873,N_22744,N_22668);
xnor U22874 (N_22874,N_22778,N_22795);
nand U22875 (N_22875,N_22603,N_22692);
nand U22876 (N_22876,N_22658,N_22610);
and U22877 (N_22877,N_22647,N_22773);
and U22878 (N_22878,N_22706,N_22632);
nand U22879 (N_22879,N_22613,N_22712);
nand U22880 (N_22880,N_22797,N_22774);
or U22881 (N_22881,N_22674,N_22719);
or U22882 (N_22882,N_22703,N_22779);
xnor U22883 (N_22883,N_22737,N_22785);
nand U22884 (N_22884,N_22638,N_22770);
or U22885 (N_22885,N_22653,N_22693);
or U22886 (N_22886,N_22679,N_22699);
xnor U22887 (N_22887,N_22644,N_22731);
or U22888 (N_22888,N_22716,N_22616);
and U22889 (N_22889,N_22728,N_22684);
nor U22890 (N_22890,N_22601,N_22752);
nand U22891 (N_22891,N_22761,N_22680);
and U22892 (N_22892,N_22607,N_22708);
nor U22893 (N_22893,N_22654,N_22665);
xor U22894 (N_22894,N_22639,N_22686);
nand U22895 (N_22895,N_22661,N_22635);
and U22896 (N_22896,N_22625,N_22645);
and U22897 (N_22897,N_22735,N_22788);
xnor U22898 (N_22898,N_22666,N_22755);
nor U22899 (N_22899,N_22681,N_22764);
xor U22900 (N_22900,N_22678,N_22671);
or U22901 (N_22901,N_22727,N_22718);
or U22902 (N_22902,N_22732,N_22761);
xor U22903 (N_22903,N_22622,N_22637);
xnor U22904 (N_22904,N_22799,N_22697);
or U22905 (N_22905,N_22748,N_22742);
nor U22906 (N_22906,N_22712,N_22798);
nand U22907 (N_22907,N_22703,N_22748);
or U22908 (N_22908,N_22728,N_22776);
nand U22909 (N_22909,N_22624,N_22633);
and U22910 (N_22910,N_22778,N_22665);
nand U22911 (N_22911,N_22706,N_22677);
and U22912 (N_22912,N_22707,N_22708);
xor U22913 (N_22913,N_22791,N_22702);
nor U22914 (N_22914,N_22784,N_22701);
nor U22915 (N_22915,N_22624,N_22774);
nor U22916 (N_22916,N_22653,N_22661);
nor U22917 (N_22917,N_22781,N_22764);
xor U22918 (N_22918,N_22609,N_22748);
nor U22919 (N_22919,N_22675,N_22637);
nor U22920 (N_22920,N_22692,N_22600);
xnor U22921 (N_22921,N_22726,N_22629);
nand U22922 (N_22922,N_22634,N_22716);
xnor U22923 (N_22923,N_22657,N_22674);
or U22924 (N_22924,N_22684,N_22655);
and U22925 (N_22925,N_22622,N_22737);
xnor U22926 (N_22926,N_22748,N_22795);
and U22927 (N_22927,N_22688,N_22764);
nor U22928 (N_22928,N_22717,N_22780);
nand U22929 (N_22929,N_22745,N_22782);
and U22930 (N_22930,N_22724,N_22674);
or U22931 (N_22931,N_22671,N_22617);
nand U22932 (N_22932,N_22661,N_22668);
xor U22933 (N_22933,N_22700,N_22752);
nor U22934 (N_22934,N_22646,N_22727);
and U22935 (N_22935,N_22677,N_22609);
and U22936 (N_22936,N_22783,N_22705);
nor U22937 (N_22937,N_22745,N_22792);
or U22938 (N_22938,N_22608,N_22747);
or U22939 (N_22939,N_22740,N_22745);
or U22940 (N_22940,N_22653,N_22764);
xnor U22941 (N_22941,N_22600,N_22653);
and U22942 (N_22942,N_22753,N_22713);
and U22943 (N_22943,N_22746,N_22723);
xnor U22944 (N_22944,N_22790,N_22799);
and U22945 (N_22945,N_22742,N_22787);
or U22946 (N_22946,N_22789,N_22752);
and U22947 (N_22947,N_22778,N_22742);
nor U22948 (N_22948,N_22748,N_22790);
nand U22949 (N_22949,N_22797,N_22698);
or U22950 (N_22950,N_22799,N_22682);
and U22951 (N_22951,N_22684,N_22796);
xor U22952 (N_22952,N_22636,N_22769);
or U22953 (N_22953,N_22725,N_22704);
or U22954 (N_22954,N_22682,N_22716);
nor U22955 (N_22955,N_22760,N_22729);
xnor U22956 (N_22956,N_22782,N_22741);
xor U22957 (N_22957,N_22697,N_22626);
or U22958 (N_22958,N_22692,N_22712);
nand U22959 (N_22959,N_22604,N_22691);
nor U22960 (N_22960,N_22648,N_22636);
or U22961 (N_22961,N_22674,N_22702);
or U22962 (N_22962,N_22641,N_22790);
or U22963 (N_22963,N_22759,N_22790);
or U22964 (N_22964,N_22688,N_22758);
nand U22965 (N_22965,N_22743,N_22719);
nor U22966 (N_22966,N_22627,N_22695);
xnor U22967 (N_22967,N_22772,N_22797);
nand U22968 (N_22968,N_22793,N_22705);
and U22969 (N_22969,N_22786,N_22788);
xor U22970 (N_22970,N_22691,N_22609);
nand U22971 (N_22971,N_22734,N_22711);
xnor U22972 (N_22972,N_22703,N_22732);
nor U22973 (N_22973,N_22645,N_22656);
and U22974 (N_22974,N_22715,N_22760);
and U22975 (N_22975,N_22625,N_22769);
and U22976 (N_22976,N_22604,N_22752);
or U22977 (N_22977,N_22621,N_22606);
nor U22978 (N_22978,N_22760,N_22711);
and U22979 (N_22979,N_22768,N_22699);
nand U22980 (N_22980,N_22703,N_22608);
or U22981 (N_22981,N_22734,N_22769);
nor U22982 (N_22982,N_22780,N_22798);
nand U22983 (N_22983,N_22675,N_22712);
xor U22984 (N_22984,N_22743,N_22779);
xnor U22985 (N_22985,N_22786,N_22712);
xor U22986 (N_22986,N_22717,N_22731);
xor U22987 (N_22987,N_22610,N_22643);
or U22988 (N_22988,N_22745,N_22747);
and U22989 (N_22989,N_22645,N_22751);
or U22990 (N_22990,N_22761,N_22787);
or U22991 (N_22991,N_22600,N_22783);
and U22992 (N_22992,N_22624,N_22729);
nand U22993 (N_22993,N_22762,N_22645);
xnor U22994 (N_22994,N_22634,N_22607);
or U22995 (N_22995,N_22739,N_22745);
and U22996 (N_22996,N_22601,N_22788);
xnor U22997 (N_22997,N_22637,N_22703);
nand U22998 (N_22998,N_22619,N_22733);
xor U22999 (N_22999,N_22602,N_22673);
xnor U23000 (N_23000,N_22878,N_22898);
and U23001 (N_23001,N_22812,N_22939);
nand U23002 (N_23002,N_22849,N_22868);
and U23003 (N_23003,N_22991,N_22866);
and U23004 (N_23004,N_22988,N_22805);
and U23005 (N_23005,N_22938,N_22990);
nand U23006 (N_23006,N_22949,N_22968);
nor U23007 (N_23007,N_22915,N_22856);
xnor U23008 (N_23008,N_22891,N_22855);
xnor U23009 (N_23009,N_22916,N_22808);
xor U23010 (N_23010,N_22961,N_22934);
or U23011 (N_23011,N_22958,N_22972);
or U23012 (N_23012,N_22930,N_22974);
and U23013 (N_23013,N_22885,N_22962);
xor U23014 (N_23014,N_22980,N_22872);
and U23015 (N_23015,N_22945,N_22998);
nor U23016 (N_23016,N_22918,N_22865);
nand U23017 (N_23017,N_22895,N_22935);
or U23018 (N_23018,N_22937,N_22944);
nand U23019 (N_23019,N_22859,N_22952);
nor U23020 (N_23020,N_22862,N_22870);
or U23021 (N_23021,N_22888,N_22904);
or U23022 (N_23022,N_22928,N_22971);
and U23023 (N_23023,N_22841,N_22853);
nand U23024 (N_23024,N_22890,N_22903);
nor U23025 (N_23025,N_22943,N_22911);
xor U23026 (N_23026,N_22925,N_22927);
and U23027 (N_23027,N_22905,N_22992);
and U23028 (N_23028,N_22803,N_22882);
and U23029 (N_23029,N_22909,N_22947);
nand U23030 (N_23030,N_22850,N_22986);
nor U23031 (N_23031,N_22838,N_22957);
nor U23032 (N_23032,N_22807,N_22953);
or U23033 (N_23033,N_22910,N_22979);
or U23034 (N_23034,N_22831,N_22987);
nor U23035 (N_23035,N_22973,N_22846);
xnor U23036 (N_23036,N_22842,N_22902);
or U23037 (N_23037,N_22860,N_22861);
nor U23038 (N_23038,N_22880,N_22879);
xor U23039 (N_23039,N_22951,N_22875);
or U23040 (N_23040,N_22995,N_22919);
xor U23041 (N_23041,N_22920,N_22914);
nor U23042 (N_23042,N_22816,N_22897);
and U23043 (N_23043,N_22960,N_22815);
and U23044 (N_23044,N_22811,N_22852);
xor U23045 (N_23045,N_22829,N_22877);
nand U23046 (N_23046,N_22926,N_22956);
nor U23047 (N_23047,N_22825,N_22997);
nor U23048 (N_23048,N_22887,N_22906);
or U23049 (N_23049,N_22837,N_22821);
xnor U23050 (N_23050,N_22940,N_22889);
nand U23051 (N_23051,N_22933,N_22976);
and U23052 (N_23052,N_22839,N_22819);
and U23053 (N_23053,N_22854,N_22892);
or U23054 (N_23054,N_22802,N_22923);
or U23055 (N_23055,N_22843,N_22941);
xor U23056 (N_23056,N_22814,N_22848);
or U23057 (N_23057,N_22901,N_22834);
xor U23058 (N_23058,N_22827,N_22857);
or U23059 (N_23059,N_22921,N_22966);
nor U23060 (N_23060,N_22828,N_22820);
and U23061 (N_23061,N_22963,N_22886);
xor U23062 (N_23062,N_22948,N_22840);
nor U23063 (N_23063,N_22817,N_22893);
or U23064 (N_23064,N_22823,N_22864);
xor U23065 (N_23065,N_22884,N_22946);
nor U23066 (N_23066,N_22800,N_22806);
xor U23067 (N_23067,N_22871,N_22975);
and U23068 (N_23068,N_22874,N_22810);
nor U23069 (N_23069,N_22908,N_22954);
nor U23070 (N_23070,N_22822,N_22867);
and U23071 (N_23071,N_22896,N_22809);
nor U23072 (N_23072,N_22931,N_22801);
xor U23073 (N_23073,N_22936,N_22832);
or U23074 (N_23074,N_22985,N_22894);
nor U23075 (N_23075,N_22845,N_22869);
xor U23076 (N_23076,N_22950,N_22826);
nor U23077 (N_23077,N_22863,N_22981);
nand U23078 (N_23078,N_22907,N_22824);
nor U23079 (N_23079,N_22876,N_22996);
or U23080 (N_23080,N_22982,N_22970);
and U23081 (N_23081,N_22858,N_22873);
and U23082 (N_23082,N_22964,N_22978);
or U23083 (N_23083,N_22965,N_22917);
nor U23084 (N_23084,N_22818,N_22881);
or U23085 (N_23085,N_22942,N_22836);
nor U23086 (N_23086,N_22984,N_22913);
and U23087 (N_23087,N_22899,N_22932);
xor U23088 (N_23088,N_22804,N_22847);
and U23089 (N_23089,N_22967,N_22900);
xor U23090 (N_23090,N_22912,N_22999);
xor U23091 (N_23091,N_22813,N_22993);
xor U23092 (N_23092,N_22959,N_22929);
nand U23093 (N_23093,N_22969,N_22989);
nor U23094 (N_23094,N_22833,N_22994);
xor U23095 (N_23095,N_22883,N_22977);
and U23096 (N_23096,N_22851,N_22924);
and U23097 (N_23097,N_22955,N_22922);
nor U23098 (N_23098,N_22835,N_22983);
nor U23099 (N_23099,N_22844,N_22830);
or U23100 (N_23100,N_22933,N_22812);
nand U23101 (N_23101,N_22827,N_22880);
xnor U23102 (N_23102,N_22905,N_22904);
xor U23103 (N_23103,N_22829,N_22896);
and U23104 (N_23104,N_22932,N_22942);
or U23105 (N_23105,N_22855,N_22968);
or U23106 (N_23106,N_22954,N_22997);
or U23107 (N_23107,N_22982,N_22869);
nand U23108 (N_23108,N_22937,N_22930);
nand U23109 (N_23109,N_22815,N_22824);
xnor U23110 (N_23110,N_22963,N_22892);
nor U23111 (N_23111,N_22984,N_22894);
nor U23112 (N_23112,N_22943,N_22893);
nand U23113 (N_23113,N_22931,N_22852);
xor U23114 (N_23114,N_22920,N_22892);
or U23115 (N_23115,N_22883,N_22917);
or U23116 (N_23116,N_22994,N_22892);
nand U23117 (N_23117,N_22951,N_22979);
and U23118 (N_23118,N_22974,N_22832);
and U23119 (N_23119,N_22986,N_22875);
and U23120 (N_23120,N_22843,N_22997);
and U23121 (N_23121,N_22985,N_22920);
nor U23122 (N_23122,N_22824,N_22956);
xor U23123 (N_23123,N_22871,N_22873);
nand U23124 (N_23124,N_22902,N_22801);
and U23125 (N_23125,N_22941,N_22881);
xnor U23126 (N_23126,N_22955,N_22809);
nand U23127 (N_23127,N_22944,N_22987);
or U23128 (N_23128,N_22889,N_22906);
nand U23129 (N_23129,N_22926,N_22904);
or U23130 (N_23130,N_22816,N_22818);
and U23131 (N_23131,N_22934,N_22805);
and U23132 (N_23132,N_22989,N_22839);
or U23133 (N_23133,N_22861,N_22840);
xnor U23134 (N_23134,N_22960,N_22847);
nand U23135 (N_23135,N_22943,N_22882);
nand U23136 (N_23136,N_22830,N_22976);
nor U23137 (N_23137,N_22824,N_22989);
nand U23138 (N_23138,N_22957,N_22996);
nand U23139 (N_23139,N_22854,N_22852);
xor U23140 (N_23140,N_22879,N_22889);
xnor U23141 (N_23141,N_22960,N_22818);
xor U23142 (N_23142,N_22994,N_22930);
nand U23143 (N_23143,N_22997,N_22897);
xor U23144 (N_23144,N_22950,N_22959);
nand U23145 (N_23145,N_22955,N_22983);
nor U23146 (N_23146,N_22900,N_22882);
nor U23147 (N_23147,N_22860,N_22824);
nor U23148 (N_23148,N_22979,N_22801);
nor U23149 (N_23149,N_22839,N_22927);
or U23150 (N_23150,N_22968,N_22950);
or U23151 (N_23151,N_22910,N_22921);
or U23152 (N_23152,N_22952,N_22863);
nand U23153 (N_23153,N_22884,N_22961);
nand U23154 (N_23154,N_22946,N_22842);
nor U23155 (N_23155,N_22900,N_22974);
or U23156 (N_23156,N_22978,N_22940);
nand U23157 (N_23157,N_22965,N_22851);
xnor U23158 (N_23158,N_22904,N_22917);
nor U23159 (N_23159,N_22992,N_22952);
and U23160 (N_23160,N_22990,N_22930);
or U23161 (N_23161,N_22955,N_22835);
nand U23162 (N_23162,N_22994,N_22952);
and U23163 (N_23163,N_22845,N_22963);
and U23164 (N_23164,N_22988,N_22864);
nand U23165 (N_23165,N_22809,N_22977);
nor U23166 (N_23166,N_22804,N_22937);
xnor U23167 (N_23167,N_22959,N_22932);
and U23168 (N_23168,N_22847,N_22922);
or U23169 (N_23169,N_22830,N_22800);
nor U23170 (N_23170,N_22974,N_22834);
and U23171 (N_23171,N_22859,N_22851);
xnor U23172 (N_23172,N_22906,N_22954);
nand U23173 (N_23173,N_22921,N_22964);
and U23174 (N_23174,N_22892,N_22933);
and U23175 (N_23175,N_22868,N_22956);
and U23176 (N_23176,N_22819,N_22951);
and U23177 (N_23177,N_22838,N_22905);
and U23178 (N_23178,N_22834,N_22855);
xnor U23179 (N_23179,N_22878,N_22899);
and U23180 (N_23180,N_22897,N_22984);
or U23181 (N_23181,N_22942,N_22834);
xor U23182 (N_23182,N_22946,N_22852);
nand U23183 (N_23183,N_22861,N_22905);
xor U23184 (N_23184,N_22924,N_22976);
nand U23185 (N_23185,N_22804,N_22972);
or U23186 (N_23186,N_22971,N_22883);
nor U23187 (N_23187,N_22857,N_22822);
or U23188 (N_23188,N_22902,N_22896);
nor U23189 (N_23189,N_22804,N_22986);
or U23190 (N_23190,N_22824,N_22978);
and U23191 (N_23191,N_22886,N_22871);
or U23192 (N_23192,N_22852,N_22871);
or U23193 (N_23193,N_22806,N_22964);
nand U23194 (N_23194,N_22836,N_22975);
xnor U23195 (N_23195,N_22893,N_22950);
xnor U23196 (N_23196,N_22928,N_22953);
nand U23197 (N_23197,N_22812,N_22991);
xnor U23198 (N_23198,N_22876,N_22904);
nand U23199 (N_23199,N_22828,N_22944);
nand U23200 (N_23200,N_23084,N_23061);
or U23201 (N_23201,N_23153,N_23194);
or U23202 (N_23202,N_23196,N_23013);
and U23203 (N_23203,N_23046,N_23011);
nor U23204 (N_23204,N_23078,N_23089);
nor U23205 (N_23205,N_23192,N_23191);
xor U23206 (N_23206,N_23002,N_23132);
xnor U23207 (N_23207,N_23164,N_23081);
nand U23208 (N_23208,N_23105,N_23107);
xor U23209 (N_23209,N_23140,N_23008);
xnor U23210 (N_23210,N_23096,N_23059);
xnor U23211 (N_23211,N_23082,N_23016);
nor U23212 (N_23212,N_23039,N_23133);
xnor U23213 (N_23213,N_23136,N_23185);
xor U23214 (N_23214,N_23029,N_23079);
or U23215 (N_23215,N_23012,N_23049);
nand U23216 (N_23216,N_23111,N_23106);
nand U23217 (N_23217,N_23052,N_23175);
nor U23218 (N_23218,N_23118,N_23033);
and U23219 (N_23219,N_23053,N_23158);
xnor U23220 (N_23220,N_23067,N_23162);
or U23221 (N_23221,N_23117,N_23120);
xnor U23222 (N_23222,N_23143,N_23064);
and U23223 (N_23223,N_23065,N_23157);
and U23224 (N_23224,N_23027,N_23155);
nor U23225 (N_23225,N_23176,N_23086);
and U23226 (N_23226,N_23001,N_23083);
and U23227 (N_23227,N_23179,N_23068);
nor U23228 (N_23228,N_23050,N_23051);
nor U23229 (N_23229,N_23110,N_23161);
or U23230 (N_23230,N_23087,N_23057);
nand U23231 (N_23231,N_23072,N_23182);
nor U23232 (N_23232,N_23152,N_23165);
nand U23233 (N_23233,N_23129,N_23075);
or U23234 (N_23234,N_23149,N_23094);
xor U23235 (N_23235,N_23198,N_23028);
nor U23236 (N_23236,N_23101,N_23095);
or U23237 (N_23237,N_23180,N_23160);
xnor U23238 (N_23238,N_23115,N_23151);
or U23239 (N_23239,N_23036,N_23171);
and U23240 (N_23240,N_23116,N_23042);
nand U23241 (N_23241,N_23063,N_23174);
nand U23242 (N_23242,N_23097,N_23128);
xnor U23243 (N_23243,N_23170,N_23184);
and U23244 (N_23244,N_23187,N_23199);
and U23245 (N_23245,N_23043,N_23023);
or U23246 (N_23246,N_23092,N_23000);
or U23247 (N_23247,N_23124,N_23126);
xnor U23248 (N_23248,N_23005,N_23195);
nor U23249 (N_23249,N_23113,N_23159);
nor U23250 (N_23250,N_23030,N_23080);
or U23251 (N_23251,N_23148,N_23026);
xnor U23252 (N_23252,N_23031,N_23193);
xnor U23253 (N_23253,N_23037,N_23134);
nand U23254 (N_23254,N_23168,N_23085);
nand U23255 (N_23255,N_23104,N_23071);
nand U23256 (N_23256,N_23041,N_23019);
xor U23257 (N_23257,N_23090,N_23098);
and U23258 (N_23258,N_23144,N_23123);
nand U23259 (N_23259,N_23006,N_23137);
and U23260 (N_23260,N_23125,N_23054);
nand U23261 (N_23261,N_23074,N_23121);
and U23262 (N_23262,N_23055,N_23135);
nand U23263 (N_23263,N_23166,N_23142);
xor U23264 (N_23264,N_23021,N_23130);
nor U23265 (N_23265,N_23169,N_23156);
xnor U23266 (N_23266,N_23062,N_23178);
and U23267 (N_23267,N_23045,N_23127);
xnor U23268 (N_23268,N_23108,N_23044);
nand U23269 (N_23269,N_23099,N_23103);
nand U23270 (N_23270,N_23017,N_23189);
nor U23271 (N_23271,N_23093,N_23139);
xor U23272 (N_23272,N_23114,N_23009);
xor U23273 (N_23273,N_23004,N_23177);
or U23274 (N_23274,N_23183,N_23003);
nor U23275 (N_23275,N_23069,N_23109);
nand U23276 (N_23276,N_23038,N_23167);
or U23277 (N_23277,N_23073,N_23014);
and U23278 (N_23278,N_23173,N_23112);
or U23279 (N_23279,N_23060,N_23186);
nor U23280 (N_23280,N_23163,N_23015);
and U23281 (N_23281,N_23007,N_23091);
and U23282 (N_23282,N_23048,N_23147);
nand U23283 (N_23283,N_23150,N_23188);
nand U23284 (N_23284,N_23032,N_23035);
nand U23285 (N_23285,N_23131,N_23066);
or U23286 (N_23286,N_23154,N_23141);
nor U23287 (N_23287,N_23056,N_23146);
nand U23288 (N_23288,N_23190,N_23047);
nor U23289 (N_23289,N_23070,N_23020);
xor U23290 (N_23290,N_23022,N_23076);
nand U23291 (N_23291,N_23138,N_23122);
nor U23292 (N_23292,N_23102,N_23024);
and U23293 (N_23293,N_23077,N_23181);
nand U23294 (N_23294,N_23018,N_23197);
nor U23295 (N_23295,N_23145,N_23040);
and U23296 (N_23296,N_23172,N_23010);
xnor U23297 (N_23297,N_23058,N_23088);
nor U23298 (N_23298,N_23119,N_23025);
xor U23299 (N_23299,N_23034,N_23100);
nor U23300 (N_23300,N_23064,N_23181);
and U23301 (N_23301,N_23023,N_23168);
and U23302 (N_23302,N_23174,N_23142);
nor U23303 (N_23303,N_23032,N_23085);
nor U23304 (N_23304,N_23175,N_23103);
xnor U23305 (N_23305,N_23079,N_23077);
nor U23306 (N_23306,N_23087,N_23055);
xor U23307 (N_23307,N_23000,N_23007);
nor U23308 (N_23308,N_23034,N_23055);
or U23309 (N_23309,N_23107,N_23163);
xor U23310 (N_23310,N_23003,N_23143);
nor U23311 (N_23311,N_23179,N_23059);
nor U23312 (N_23312,N_23028,N_23003);
and U23313 (N_23313,N_23089,N_23184);
or U23314 (N_23314,N_23022,N_23176);
and U23315 (N_23315,N_23011,N_23121);
xnor U23316 (N_23316,N_23000,N_23022);
nand U23317 (N_23317,N_23107,N_23094);
xor U23318 (N_23318,N_23098,N_23152);
xnor U23319 (N_23319,N_23092,N_23162);
or U23320 (N_23320,N_23191,N_23078);
nor U23321 (N_23321,N_23025,N_23162);
xnor U23322 (N_23322,N_23132,N_23061);
nor U23323 (N_23323,N_23017,N_23179);
nand U23324 (N_23324,N_23082,N_23138);
nand U23325 (N_23325,N_23156,N_23002);
nand U23326 (N_23326,N_23023,N_23050);
or U23327 (N_23327,N_23180,N_23015);
nor U23328 (N_23328,N_23108,N_23034);
xnor U23329 (N_23329,N_23096,N_23112);
xor U23330 (N_23330,N_23163,N_23184);
xor U23331 (N_23331,N_23104,N_23137);
nor U23332 (N_23332,N_23196,N_23018);
nor U23333 (N_23333,N_23164,N_23013);
nand U23334 (N_23334,N_23023,N_23117);
xnor U23335 (N_23335,N_23085,N_23185);
nor U23336 (N_23336,N_23099,N_23141);
and U23337 (N_23337,N_23063,N_23149);
and U23338 (N_23338,N_23153,N_23109);
nand U23339 (N_23339,N_23155,N_23071);
and U23340 (N_23340,N_23008,N_23136);
or U23341 (N_23341,N_23110,N_23160);
xor U23342 (N_23342,N_23096,N_23166);
xnor U23343 (N_23343,N_23161,N_23186);
xnor U23344 (N_23344,N_23086,N_23140);
and U23345 (N_23345,N_23097,N_23049);
nor U23346 (N_23346,N_23148,N_23049);
xnor U23347 (N_23347,N_23039,N_23045);
nor U23348 (N_23348,N_23195,N_23176);
nand U23349 (N_23349,N_23016,N_23170);
xnor U23350 (N_23350,N_23123,N_23185);
nor U23351 (N_23351,N_23003,N_23034);
xnor U23352 (N_23352,N_23127,N_23131);
nand U23353 (N_23353,N_23110,N_23091);
or U23354 (N_23354,N_23025,N_23128);
xnor U23355 (N_23355,N_23109,N_23029);
xnor U23356 (N_23356,N_23198,N_23085);
xor U23357 (N_23357,N_23139,N_23143);
or U23358 (N_23358,N_23009,N_23110);
nand U23359 (N_23359,N_23169,N_23064);
nor U23360 (N_23360,N_23073,N_23135);
xor U23361 (N_23361,N_23087,N_23007);
nor U23362 (N_23362,N_23112,N_23106);
nor U23363 (N_23363,N_23029,N_23171);
and U23364 (N_23364,N_23186,N_23047);
nand U23365 (N_23365,N_23085,N_23148);
or U23366 (N_23366,N_23195,N_23030);
xnor U23367 (N_23367,N_23148,N_23136);
nor U23368 (N_23368,N_23048,N_23175);
xnor U23369 (N_23369,N_23044,N_23127);
or U23370 (N_23370,N_23030,N_23187);
nand U23371 (N_23371,N_23164,N_23127);
nand U23372 (N_23372,N_23053,N_23122);
xor U23373 (N_23373,N_23000,N_23192);
and U23374 (N_23374,N_23076,N_23063);
nand U23375 (N_23375,N_23154,N_23084);
and U23376 (N_23376,N_23062,N_23034);
nand U23377 (N_23377,N_23049,N_23151);
and U23378 (N_23378,N_23099,N_23194);
or U23379 (N_23379,N_23112,N_23083);
and U23380 (N_23380,N_23005,N_23178);
nand U23381 (N_23381,N_23047,N_23083);
nor U23382 (N_23382,N_23180,N_23032);
and U23383 (N_23383,N_23102,N_23134);
xor U23384 (N_23384,N_23006,N_23063);
nand U23385 (N_23385,N_23011,N_23019);
and U23386 (N_23386,N_23078,N_23057);
xnor U23387 (N_23387,N_23165,N_23092);
nor U23388 (N_23388,N_23020,N_23081);
or U23389 (N_23389,N_23108,N_23060);
xor U23390 (N_23390,N_23164,N_23005);
and U23391 (N_23391,N_23041,N_23187);
nor U23392 (N_23392,N_23186,N_23032);
and U23393 (N_23393,N_23074,N_23065);
and U23394 (N_23394,N_23125,N_23159);
nand U23395 (N_23395,N_23064,N_23093);
xnor U23396 (N_23396,N_23073,N_23084);
or U23397 (N_23397,N_23060,N_23055);
nand U23398 (N_23398,N_23032,N_23024);
nor U23399 (N_23399,N_23179,N_23109);
nand U23400 (N_23400,N_23398,N_23364);
and U23401 (N_23401,N_23316,N_23282);
nor U23402 (N_23402,N_23328,N_23231);
nand U23403 (N_23403,N_23389,N_23355);
and U23404 (N_23404,N_23343,N_23256);
nand U23405 (N_23405,N_23358,N_23253);
nor U23406 (N_23406,N_23326,N_23220);
or U23407 (N_23407,N_23266,N_23327);
nand U23408 (N_23408,N_23319,N_23271);
nor U23409 (N_23409,N_23232,N_23320);
nand U23410 (N_23410,N_23290,N_23393);
nand U23411 (N_23411,N_23242,N_23207);
or U23412 (N_23412,N_23276,N_23341);
or U23413 (N_23413,N_23272,N_23308);
nor U23414 (N_23414,N_23375,N_23273);
xnor U23415 (N_23415,N_23336,N_23222);
and U23416 (N_23416,N_23251,N_23299);
or U23417 (N_23417,N_23309,N_23218);
nor U23418 (N_23418,N_23278,N_23295);
xnor U23419 (N_23419,N_23270,N_23318);
xnor U23420 (N_23420,N_23324,N_23380);
or U23421 (N_23421,N_23313,N_23209);
nand U23422 (N_23422,N_23368,N_23377);
nor U23423 (N_23423,N_23345,N_23314);
nand U23424 (N_23424,N_23214,N_23296);
nor U23425 (N_23425,N_23286,N_23219);
nor U23426 (N_23426,N_23373,N_23221);
or U23427 (N_23427,N_23330,N_23352);
nor U23428 (N_23428,N_23339,N_23204);
xnor U23429 (N_23429,N_23386,N_23321);
nor U23430 (N_23430,N_23356,N_23285);
nor U23431 (N_23431,N_23293,N_23239);
xor U23432 (N_23432,N_23234,N_23268);
or U23433 (N_23433,N_23381,N_23390);
or U23434 (N_23434,N_23379,N_23280);
nand U23435 (N_23435,N_23211,N_23240);
nand U23436 (N_23436,N_23396,N_23365);
xor U23437 (N_23437,N_23310,N_23274);
nand U23438 (N_23438,N_23227,N_23262);
and U23439 (N_23439,N_23243,N_23241);
nor U23440 (N_23440,N_23325,N_23384);
and U23441 (N_23441,N_23264,N_23250);
nand U23442 (N_23442,N_23287,N_23357);
nor U23443 (N_23443,N_23298,N_23340);
nand U23444 (N_23444,N_23237,N_23351);
nor U23445 (N_23445,N_23317,N_23279);
nor U23446 (N_23446,N_23203,N_23329);
nor U23447 (N_23447,N_23344,N_23323);
nor U23448 (N_23448,N_23304,N_23247);
nand U23449 (N_23449,N_23283,N_23382);
and U23450 (N_23450,N_23391,N_23322);
nor U23451 (N_23451,N_23225,N_23347);
or U23452 (N_23452,N_23301,N_23236);
and U23453 (N_23453,N_23294,N_23223);
nand U23454 (N_23454,N_23258,N_23371);
nand U23455 (N_23455,N_23353,N_23230);
or U23456 (N_23456,N_23255,N_23210);
or U23457 (N_23457,N_23284,N_23315);
and U23458 (N_23458,N_23363,N_23332);
nand U23459 (N_23459,N_23254,N_23392);
nand U23460 (N_23460,N_23361,N_23267);
nor U23461 (N_23461,N_23263,N_23201);
xnor U23462 (N_23462,N_23307,N_23269);
xnor U23463 (N_23463,N_23248,N_23349);
nor U23464 (N_23464,N_23235,N_23338);
xor U23465 (N_23465,N_23394,N_23369);
and U23466 (N_23466,N_23215,N_23244);
and U23467 (N_23467,N_23229,N_23306);
nand U23468 (N_23468,N_23224,N_23261);
xor U23469 (N_23469,N_23228,N_23331);
xnor U23470 (N_23470,N_23300,N_23387);
or U23471 (N_23471,N_23399,N_23372);
or U23472 (N_23472,N_23370,N_23397);
nand U23473 (N_23473,N_23367,N_23205);
nand U23474 (N_23474,N_23202,N_23312);
or U23475 (N_23475,N_23291,N_23388);
nor U23476 (N_23476,N_23217,N_23311);
nor U23477 (N_23477,N_23305,N_23337);
nor U23478 (N_23478,N_23212,N_23259);
or U23479 (N_23479,N_23249,N_23360);
nand U23480 (N_23480,N_23208,N_23302);
nand U23481 (N_23481,N_23333,N_23385);
nor U23482 (N_23482,N_23200,N_23245);
nor U23483 (N_23483,N_23395,N_23275);
or U23484 (N_23484,N_23233,N_23383);
nor U23485 (N_23485,N_23292,N_23265);
nor U23486 (N_23486,N_23238,N_23346);
or U23487 (N_23487,N_23289,N_23354);
nand U23488 (N_23488,N_23378,N_23213);
and U23489 (N_23489,N_23252,N_23226);
nor U23490 (N_23490,N_23350,N_23374);
xnor U23491 (N_23491,N_23376,N_23303);
and U23492 (N_23492,N_23288,N_23359);
nand U23493 (N_23493,N_23348,N_23216);
nand U23494 (N_23494,N_23257,N_23246);
or U23495 (N_23495,N_23342,N_23335);
and U23496 (N_23496,N_23206,N_23297);
nand U23497 (N_23497,N_23366,N_23362);
nand U23498 (N_23498,N_23260,N_23281);
nor U23499 (N_23499,N_23334,N_23277);
nor U23500 (N_23500,N_23224,N_23318);
and U23501 (N_23501,N_23275,N_23311);
nand U23502 (N_23502,N_23230,N_23265);
nor U23503 (N_23503,N_23321,N_23360);
or U23504 (N_23504,N_23285,N_23213);
nand U23505 (N_23505,N_23229,N_23273);
and U23506 (N_23506,N_23366,N_23266);
or U23507 (N_23507,N_23209,N_23214);
nor U23508 (N_23508,N_23313,N_23330);
xnor U23509 (N_23509,N_23382,N_23271);
nand U23510 (N_23510,N_23331,N_23381);
xor U23511 (N_23511,N_23243,N_23364);
or U23512 (N_23512,N_23350,N_23353);
xor U23513 (N_23513,N_23361,N_23313);
nand U23514 (N_23514,N_23263,N_23329);
xor U23515 (N_23515,N_23320,N_23207);
or U23516 (N_23516,N_23260,N_23337);
nor U23517 (N_23517,N_23342,N_23259);
nand U23518 (N_23518,N_23343,N_23325);
or U23519 (N_23519,N_23267,N_23235);
and U23520 (N_23520,N_23388,N_23222);
or U23521 (N_23521,N_23287,N_23332);
nand U23522 (N_23522,N_23232,N_23207);
nor U23523 (N_23523,N_23236,N_23268);
nand U23524 (N_23524,N_23329,N_23369);
nor U23525 (N_23525,N_23369,N_23382);
xor U23526 (N_23526,N_23352,N_23389);
or U23527 (N_23527,N_23316,N_23383);
xor U23528 (N_23528,N_23219,N_23217);
and U23529 (N_23529,N_23391,N_23334);
and U23530 (N_23530,N_23220,N_23313);
or U23531 (N_23531,N_23233,N_23290);
nand U23532 (N_23532,N_23339,N_23313);
or U23533 (N_23533,N_23204,N_23258);
nor U23534 (N_23534,N_23366,N_23326);
nand U23535 (N_23535,N_23346,N_23297);
or U23536 (N_23536,N_23235,N_23369);
or U23537 (N_23537,N_23344,N_23396);
nor U23538 (N_23538,N_23258,N_23379);
nor U23539 (N_23539,N_23320,N_23343);
xor U23540 (N_23540,N_23368,N_23222);
nand U23541 (N_23541,N_23327,N_23354);
xor U23542 (N_23542,N_23282,N_23312);
nand U23543 (N_23543,N_23209,N_23247);
and U23544 (N_23544,N_23319,N_23363);
and U23545 (N_23545,N_23202,N_23260);
nor U23546 (N_23546,N_23380,N_23396);
nand U23547 (N_23547,N_23390,N_23312);
nand U23548 (N_23548,N_23399,N_23213);
xor U23549 (N_23549,N_23385,N_23209);
xor U23550 (N_23550,N_23213,N_23214);
nor U23551 (N_23551,N_23385,N_23323);
nor U23552 (N_23552,N_23339,N_23327);
and U23553 (N_23553,N_23346,N_23357);
nor U23554 (N_23554,N_23228,N_23330);
and U23555 (N_23555,N_23290,N_23202);
xnor U23556 (N_23556,N_23310,N_23220);
nor U23557 (N_23557,N_23328,N_23340);
xnor U23558 (N_23558,N_23247,N_23363);
or U23559 (N_23559,N_23337,N_23324);
and U23560 (N_23560,N_23326,N_23383);
or U23561 (N_23561,N_23326,N_23362);
or U23562 (N_23562,N_23205,N_23212);
and U23563 (N_23563,N_23306,N_23327);
xor U23564 (N_23564,N_23249,N_23333);
xnor U23565 (N_23565,N_23242,N_23263);
nand U23566 (N_23566,N_23224,N_23246);
or U23567 (N_23567,N_23322,N_23222);
nand U23568 (N_23568,N_23314,N_23334);
and U23569 (N_23569,N_23251,N_23369);
or U23570 (N_23570,N_23239,N_23370);
xor U23571 (N_23571,N_23317,N_23245);
or U23572 (N_23572,N_23224,N_23288);
xor U23573 (N_23573,N_23330,N_23310);
xor U23574 (N_23574,N_23325,N_23230);
nand U23575 (N_23575,N_23361,N_23286);
nor U23576 (N_23576,N_23239,N_23398);
nand U23577 (N_23577,N_23269,N_23280);
nor U23578 (N_23578,N_23238,N_23264);
xor U23579 (N_23579,N_23284,N_23242);
xor U23580 (N_23580,N_23286,N_23355);
nand U23581 (N_23581,N_23309,N_23239);
nand U23582 (N_23582,N_23217,N_23331);
or U23583 (N_23583,N_23373,N_23283);
xnor U23584 (N_23584,N_23313,N_23380);
or U23585 (N_23585,N_23244,N_23398);
xnor U23586 (N_23586,N_23259,N_23307);
nor U23587 (N_23587,N_23336,N_23334);
xnor U23588 (N_23588,N_23263,N_23209);
nor U23589 (N_23589,N_23389,N_23338);
and U23590 (N_23590,N_23310,N_23209);
or U23591 (N_23591,N_23280,N_23340);
nand U23592 (N_23592,N_23294,N_23286);
or U23593 (N_23593,N_23297,N_23359);
nand U23594 (N_23594,N_23280,N_23299);
nand U23595 (N_23595,N_23277,N_23260);
or U23596 (N_23596,N_23322,N_23304);
or U23597 (N_23597,N_23349,N_23207);
or U23598 (N_23598,N_23398,N_23345);
and U23599 (N_23599,N_23279,N_23269);
and U23600 (N_23600,N_23524,N_23410);
or U23601 (N_23601,N_23436,N_23448);
or U23602 (N_23602,N_23592,N_23591);
xnor U23603 (N_23603,N_23541,N_23508);
or U23604 (N_23604,N_23469,N_23593);
and U23605 (N_23605,N_23573,N_23523);
or U23606 (N_23606,N_23504,N_23493);
nor U23607 (N_23607,N_23483,N_23444);
xnor U23608 (N_23608,N_23519,N_23528);
and U23609 (N_23609,N_23516,N_23569);
and U23610 (N_23610,N_23470,N_23467);
and U23611 (N_23611,N_23513,N_23533);
and U23612 (N_23612,N_23505,N_23407);
and U23613 (N_23613,N_23438,N_23471);
and U23614 (N_23614,N_23501,N_23472);
nor U23615 (N_23615,N_23453,N_23535);
or U23616 (N_23616,N_23587,N_23478);
and U23617 (N_23617,N_23537,N_23550);
nor U23618 (N_23618,N_23595,N_23427);
or U23619 (N_23619,N_23416,N_23545);
nor U23620 (N_23620,N_23579,N_23589);
nor U23621 (N_23621,N_23577,N_23538);
and U23622 (N_23622,N_23485,N_23433);
nand U23623 (N_23623,N_23542,N_23449);
and U23624 (N_23624,N_23571,N_23582);
and U23625 (N_23625,N_23580,N_23463);
and U23626 (N_23626,N_23455,N_23498);
nand U23627 (N_23627,N_23583,N_23534);
nor U23628 (N_23628,N_23451,N_23423);
nor U23629 (N_23629,N_23584,N_23430);
and U23630 (N_23630,N_23531,N_23565);
nand U23631 (N_23631,N_23417,N_23500);
xnor U23632 (N_23632,N_23559,N_23495);
nand U23633 (N_23633,N_23465,N_23487);
xnor U23634 (N_23634,N_23494,N_23567);
nand U23635 (N_23635,N_23517,N_23461);
or U23636 (N_23636,N_23415,N_23484);
xor U23637 (N_23637,N_23553,N_23434);
nand U23638 (N_23638,N_23568,N_23409);
nor U23639 (N_23639,N_23489,N_23539);
and U23640 (N_23640,N_23413,N_23400);
nand U23641 (N_23641,N_23540,N_23402);
xnor U23642 (N_23642,N_23473,N_23464);
or U23643 (N_23643,N_23462,N_23514);
xnor U23644 (N_23644,N_23425,N_23586);
and U23645 (N_23645,N_23554,N_23570);
nand U23646 (N_23646,N_23441,N_23522);
nor U23647 (N_23647,N_23560,N_23401);
or U23648 (N_23648,N_23414,N_23428);
nor U23649 (N_23649,N_23403,N_23459);
xnor U23650 (N_23650,N_23581,N_23419);
xnor U23651 (N_23651,N_23510,N_23437);
xor U23652 (N_23652,N_23549,N_23511);
xor U23653 (N_23653,N_23450,N_23447);
or U23654 (N_23654,N_23561,N_23594);
nand U23655 (N_23655,N_23479,N_23555);
and U23656 (N_23656,N_23576,N_23599);
nor U23657 (N_23657,N_23548,N_23532);
or U23658 (N_23658,N_23527,N_23497);
nor U23659 (N_23659,N_23468,N_23481);
nor U23660 (N_23660,N_23518,N_23486);
xor U23661 (N_23661,N_23597,N_23544);
nor U23662 (N_23662,N_23488,N_23475);
xnor U23663 (N_23663,N_23543,N_23422);
nand U23664 (N_23664,N_23490,N_23454);
xnor U23665 (N_23665,N_23418,N_23426);
and U23666 (N_23666,N_23529,N_23482);
nand U23667 (N_23667,N_23598,N_23421);
or U23668 (N_23668,N_23578,N_23491);
xor U23669 (N_23669,N_23526,N_23445);
or U23670 (N_23670,N_23474,N_23408);
nand U23671 (N_23671,N_23557,N_23562);
nand U23672 (N_23672,N_23460,N_23457);
xor U23673 (N_23673,N_23536,N_23546);
nor U23674 (N_23674,N_23492,N_23520);
xnor U23675 (N_23675,N_23456,N_23440);
or U23676 (N_23676,N_23435,N_23439);
or U23677 (N_23677,N_23412,N_23525);
or U23678 (N_23678,N_23551,N_23507);
xnor U23679 (N_23679,N_23420,N_23575);
nor U23680 (N_23680,N_23443,N_23574);
nor U23681 (N_23681,N_23566,N_23590);
and U23682 (N_23682,N_23564,N_23411);
or U23683 (N_23683,N_23477,N_23552);
nor U23684 (N_23684,N_23432,N_23530);
nand U23685 (N_23685,N_23496,N_23404);
or U23686 (N_23686,N_23502,N_23556);
nand U23687 (N_23687,N_23405,N_23521);
or U23688 (N_23688,N_23458,N_23431);
nand U23689 (N_23689,N_23406,N_23446);
and U23690 (N_23690,N_23503,N_23563);
or U23691 (N_23691,N_23572,N_23466);
and U23692 (N_23692,N_23424,N_23515);
nand U23693 (N_23693,N_23547,N_23480);
xnor U23694 (N_23694,N_23585,N_23558);
xnor U23695 (N_23695,N_23429,N_23509);
nor U23696 (N_23696,N_23442,N_23499);
nor U23697 (N_23697,N_23588,N_23452);
xnor U23698 (N_23698,N_23506,N_23596);
or U23699 (N_23699,N_23512,N_23476);
and U23700 (N_23700,N_23584,N_23428);
or U23701 (N_23701,N_23485,N_23419);
and U23702 (N_23702,N_23517,N_23403);
xor U23703 (N_23703,N_23471,N_23485);
nand U23704 (N_23704,N_23562,N_23594);
or U23705 (N_23705,N_23428,N_23579);
or U23706 (N_23706,N_23593,N_23468);
and U23707 (N_23707,N_23429,N_23405);
nand U23708 (N_23708,N_23579,N_23509);
xor U23709 (N_23709,N_23478,N_23513);
xnor U23710 (N_23710,N_23533,N_23559);
or U23711 (N_23711,N_23526,N_23505);
nor U23712 (N_23712,N_23552,N_23457);
nor U23713 (N_23713,N_23412,N_23406);
or U23714 (N_23714,N_23401,N_23501);
or U23715 (N_23715,N_23458,N_23468);
nor U23716 (N_23716,N_23591,N_23560);
xnor U23717 (N_23717,N_23543,N_23533);
or U23718 (N_23718,N_23590,N_23531);
or U23719 (N_23719,N_23432,N_23587);
and U23720 (N_23720,N_23504,N_23485);
and U23721 (N_23721,N_23416,N_23406);
or U23722 (N_23722,N_23446,N_23514);
and U23723 (N_23723,N_23492,N_23514);
nand U23724 (N_23724,N_23430,N_23446);
nand U23725 (N_23725,N_23470,N_23504);
or U23726 (N_23726,N_23507,N_23460);
nand U23727 (N_23727,N_23481,N_23529);
or U23728 (N_23728,N_23565,N_23576);
and U23729 (N_23729,N_23524,N_23404);
or U23730 (N_23730,N_23560,N_23448);
nand U23731 (N_23731,N_23515,N_23416);
or U23732 (N_23732,N_23537,N_23586);
and U23733 (N_23733,N_23554,N_23427);
xnor U23734 (N_23734,N_23477,N_23554);
or U23735 (N_23735,N_23586,N_23463);
nand U23736 (N_23736,N_23457,N_23593);
nand U23737 (N_23737,N_23499,N_23489);
nor U23738 (N_23738,N_23417,N_23504);
xnor U23739 (N_23739,N_23473,N_23443);
and U23740 (N_23740,N_23523,N_23480);
xnor U23741 (N_23741,N_23504,N_23557);
and U23742 (N_23742,N_23537,N_23569);
or U23743 (N_23743,N_23587,N_23562);
xor U23744 (N_23744,N_23465,N_23454);
and U23745 (N_23745,N_23421,N_23575);
nor U23746 (N_23746,N_23542,N_23492);
xnor U23747 (N_23747,N_23480,N_23568);
xor U23748 (N_23748,N_23508,N_23445);
nor U23749 (N_23749,N_23590,N_23495);
or U23750 (N_23750,N_23553,N_23483);
and U23751 (N_23751,N_23514,N_23459);
nor U23752 (N_23752,N_23591,N_23556);
xor U23753 (N_23753,N_23415,N_23560);
nand U23754 (N_23754,N_23448,N_23539);
nand U23755 (N_23755,N_23487,N_23583);
or U23756 (N_23756,N_23558,N_23416);
nand U23757 (N_23757,N_23462,N_23591);
and U23758 (N_23758,N_23536,N_23575);
nand U23759 (N_23759,N_23551,N_23488);
and U23760 (N_23760,N_23536,N_23435);
and U23761 (N_23761,N_23475,N_23437);
or U23762 (N_23762,N_23442,N_23469);
nor U23763 (N_23763,N_23498,N_23585);
or U23764 (N_23764,N_23545,N_23451);
nor U23765 (N_23765,N_23432,N_23518);
nor U23766 (N_23766,N_23471,N_23540);
nor U23767 (N_23767,N_23553,N_23469);
xor U23768 (N_23768,N_23578,N_23501);
nor U23769 (N_23769,N_23507,N_23415);
xnor U23770 (N_23770,N_23410,N_23458);
and U23771 (N_23771,N_23405,N_23461);
or U23772 (N_23772,N_23474,N_23428);
nor U23773 (N_23773,N_23508,N_23436);
nand U23774 (N_23774,N_23495,N_23478);
and U23775 (N_23775,N_23461,N_23557);
and U23776 (N_23776,N_23570,N_23472);
xnor U23777 (N_23777,N_23518,N_23448);
and U23778 (N_23778,N_23585,N_23590);
nor U23779 (N_23779,N_23519,N_23514);
or U23780 (N_23780,N_23587,N_23475);
nor U23781 (N_23781,N_23520,N_23590);
xor U23782 (N_23782,N_23507,N_23466);
nor U23783 (N_23783,N_23541,N_23425);
or U23784 (N_23784,N_23458,N_23485);
nor U23785 (N_23785,N_23513,N_23588);
or U23786 (N_23786,N_23488,N_23502);
xnor U23787 (N_23787,N_23445,N_23405);
nand U23788 (N_23788,N_23426,N_23472);
or U23789 (N_23789,N_23490,N_23427);
or U23790 (N_23790,N_23582,N_23458);
nor U23791 (N_23791,N_23533,N_23506);
and U23792 (N_23792,N_23452,N_23583);
nor U23793 (N_23793,N_23570,N_23428);
xnor U23794 (N_23794,N_23474,N_23509);
nand U23795 (N_23795,N_23476,N_23477);
nor U23796 (N_23796,N_23447,N_23585);
and U23797 (N_23797,N_23585,N_23418);
or U23798 (N_23798,N_23440,N_23542);
and U23799 (N_23799,N_23504,N_23571);
xnor U23800 (N_23800,N_23761,N_23721);
nor U23801 (N_23801,N_23760,N_23649);
nor U23802 (N_23802,N_23778,N_23781);
nand U23803 (N_23803,N_23793,N_23794);
nor U23804 (N_23804,N_23777,N_23742);
or U23805 (N_23805,N_23653,N_23767);
or U23806 (N_23806,N_23636,N_23634);
and U23807 (N_23807,N_23678,N_23696);
xnor U23808 (N_23808,N_23662,N_23773);
nor U23809 (N_23809,N_23618,N_23744);
xnor U23810 (N_23810,N_23709,N_23762);
nand U23811 (N_23811,N_23642,N_23716);
or U23812 (N_23812,N_23681,N_23726);
xnor U23813 (N_23813,N_23701,N_23713);
nand U23814 (N_23814,N_23771,N_23787);
xnor U23815 (N_23815,N_23729,N_23748);
nor U23816 (N_23816,N_23743,N_23775);
nand U23817 (N_23817,N_23757,N_23699);
nor U23818 (N_23818,N_23605,N_23647);
xnor U23819 (N_23819,N_23658,N_23671);
nor U23820 (N_23820,N_23703,N_23786);
and U23821 (N_23821,N_23629,N_23625);
xor U23822 (N_23822,N_23666,N_23619);
nand U23823 (N_23823,N_23611,N_23790);
and U23824 (N_23824,N_23646,N_23604);
and U23825 (N_23825,N_23644,N_23704);
nand U23826 (N_23826,N_23684,N_23667);
nor U23827 (N_23827,N_23797,N_23745);
and U23828 (N_23828,N_23631,N_23645);
nand U23829 (N_23829,N_23774,N_23732);
or U23830 (N_23830,N_23680,N_23659);
nor U23831 (N_23831,N_23620,N_23609);
nand U23832 (N_23832,N_23627,N_23788);
and U23833 (N_23833,N_23792,N_23676);
nor U23834 (N_23834,N_23692,N_23612);
or U23835 (N_23835,N_23798,N_23746);
nor U23836 (N_23836,N_23769,N_23621);
or U23837 (N_23837,N_23683,N_23628);
or U23838 (N_23838,N_23724,N_23617);
nor U23839 (N_23839,N_23613,N_23750);
or U23840 (N_23840,N_23755,N_23664);
or U23841 (N_23841,N_23641,N_23686);
nand U23842 (N_23842,N_23710,N_23648);
xor U23843 (N_23843,N_23633,N_23722);
and U23844 (N_23844,N_23640,N_23727);
or U23845 (N_23845,N_23690,N_23725);
nor U23846 (N_23846,N_23615,N_23776);
or U23847 (N_23847,N_23623,N_23740);
or U23848 (N_23848,N_23702,N_23707);
or U23849 (N_23849,N_23624,N_23736);
xnor U23850 (N_23850,N_23655,N_23718);
nand U23851 (N_23851,N_23697,N_23749);
nor U23852 (N_23852,N_23714,N_23772);
nor U23853 (N_23853,N_23685,N_23679);
or U23854 (N_23854,N_23734,N_23657);
nand U23855 (N_23855,N_23616,N_23795);
and U23856 (N_23856,N_23688,N_23728);
xnor U23857 (N_23857,N_23751,N_23675);
nand U23858 (N_23858,N_23747,N_23601);
nand U23859 (N_23859,N_23717,N_23614);
nand U23860 (N_23860,N_23763,N_23695);
xor U23861 (N_23861,N_23731,N_23674);
xnor U23862 (N_23862,N_23715,N_23737);
nor U23863 (N_23863,N_23630,N_23708);
xor U23864 (N_23864,N_23610,N_23723);
nand U23865 (N_23865,N_23639,N_23651);
and U23866 (N_23866,N_23687,N_23677);
and U23867 (N_23867,N_23637,N_23741);
or U23868 (N_23868,N_23785,N_23770);
nand U23869 (N_23869,N_23600,N_23622);
xnor U23870 (N_23870,N_23643,N_23753);
nor U23871 (N_23871,N_23602,N_23668);
or U23872 (N_23872,N_23660,N_23756);
or U23873 (N_23873,N_23656,N_23733);
nand U23874 (N_23874,N_23796,N_23661);
or U23875 (N_23875,N_23780,N_23608);
and U23876 (N_23876,N_23673,N_23759);
nor U23877 (N_23877,N_23730,N_23752);
or U23878 (N_23878,N_23694,N_23765);
nor U23879 (N_23879,N_23783,N_23712);
nand U23880 (N_23880,N_23635,N_23738);
nor U23881 (N_23881,N_23663,N_23789);
xor U23882 (N_23882,N_23669,N_23768);
nor U23883 (N_23883,N_23766,N_23689);
and U23884 (N_23884,N_23739,N_23799);
nor U23885 (N_23885,N_23654,N_23652);
and U23886 (N_23886,N_23711,N_23698);
or U23887 (N_23887,N_23638,N_23626);
nand U23888 (N_23888,N_23720,N_23693);
or U23889 (N_23889,N_23735,N_23607);
and U23890 (N_23890,N_23706,N_23700);
xnor U23891 (N_23891,N_23606,N_23705);
or U23892 (N_23892,N_23632,N_23784);
xor U23893 (N_23893,N_23782,N_23791);
and U23894 (N_23894,N_23758,N_23603);
nand U23895 (N_23895,N_23670,N_23665);
xor U23896 (N_23896,N_23650,N_23682);
nand U23897 (N_23897,N_23672,N_23754);
nand U23898 (N_23898,N_23719,N_23691);
xnor U23899 (N_23899,N_23779,N_23764);
or U23900 (N_23900,N_23662,N_23784);
xnor U23901 (N_23901,N_23700,N_23619);
nand U23902 (N_23902,N_23768,N_23672);
nor U23903 (N_23903,N_23625,N_23718);
nand U23904 (N_23904,N_23658,N_23752);
nor U23905 (N_23905,N_23779,N_23669);
nand U23906 (N_23906,N_23793,N_23767);
or U23907 (N_23907,N_23761,N_23641);
nand U23908 (N_23908,N_23665,N_23721);
or U23909 (N_23909,N_23722,N_23680);
nand U23910 (N_23910,N_23766,N_23636);
nand U23911 (N_23911,N_23728,N_23605);
xnor U23912 (N_23912,N_23790,N_23604);
and U23913 (N_23913,N_23612,N_23636);
nor U23914 (N_23914,N_23694,N_23622);
nand U23915 (N_23915,N_23731,N_23727);
nand U23916 (N_23916,N_23722,N_23690);
nor U23917 (N_23917,N_23759,N_23679);
or U23918 (N_23918,N_23719,N_23752);
xor U23919 (N_23919,N_23722,N_23658);
nand U23920 (N_23920,N_23666,N_23656);
nand U23921 (N_23921,N_23625,N_23791);
and U23922 (N_23922,N_23799,N_23745);
nand U23923 (N_23923,N_23735,N_23790);
nor U23924 (N_23924,N_23706,N_23790);
and U23925 (N_23925,N_23657,N_23725);
nor U23926 (N_23926,N_23679,N_23699);
and U23927 (N_23927,N_23760,N_23626);
and U23928 (N_23928,N_23736,N_23621);
nand U23929 (N_23929,N_23731,N_23695);
and U23930 (N_23930,N_23716,N_23686);
or U23931 (N_23931,N_23640,N_23793);
xnor U23932 (N_23932,N_23785,N_23750);
nand U23933 (N_23933,N_23786,N_23733);
and U23934 (N_23934,N_23647,N_23769);
nor U23935 (N_23935,N_23751,N_23714);
xor U23936 (N_23936,N_23746,N_23649);
or U23937 (N_23937,N_23633,N_23789);
nand U23938 (N_23938,N_23641,N_23638);
nand U23939 (N_23939,N_23707,N_23611);
or U23940 (N_23940,N_23639,N_23770);
xnor U23941 (N_23941,N_23751,N_23637);
nand U23942 (N_23942,N_23768,N_23687);
nand U23943 (N_23943,N_23678,N_23627);
nand U23944 (N_23944,N_23767,N_23750);
nand U23945 (N_23945,N_23777,N_23636);
nor U23946 (N_23946,N_23617,N_23794);
and U23947 (N_23947,N_23698,N_23724);
nand U23948 (N_23948,N_23669,N_23715);
nor U23949 (N_23949,N_23776,N_23719);
or U23950 (N_23950,N_23679,N_23735);
nand U23951 (N_23951,N_23641,N_23706);
nor U23952 (N_23952,N_23735,N_23759);
nand U23953 (N_23953,N_23799,N_23701);
or U23954 (N_23954,N_23722,N_23613);
or U23955 (N_23955,N_23712,N_23701);
and U23956 (N_23956,N_23730,N_23630);
nand U23957 (N_23957,N_23669,N_23656);
xnor U23958 (N_23958,N_23620,N_23716);
and U23959 (N_23959,N_23759,N_23705);
or U23960 (N_23960,N_23692,N_23634);
nor U23961 (N_23961,N_23732,N_23736);
nor U23962 (N_23962,N_23690,N_23689);
nor U23963 (N_23963,N_23655,N_23742);
and U23964 (N_23964,N_23787,N_23768);
nand U23965 (N_23965,N_23616,N_23757);
nand U23966 (N_23966,N_23680,N_23601);
nand U23967 (N_23967,N_23638,N_23773);
and U23968 (N_23968,N_23715,N_23625);
nor U23969 (N_23969,N_23654,N_23776);
xnor U23970 (N_23970,N_23606,N_23628);
nand U23971 (N_23971,N_23719,N_23664);
xor U23972 (N_23972,N_23666,N_23764);
and U23973 (N_23973,N_23771,N_23657);
xnor U23974 (N_23974,N_23691,N_23779);
nand U23975 (N_23975,N_23779,N_23636);
nor U23976 (N_23976,N_23712,N_23796);
or U23977 (N_23977,N_23678,N_23616);
xor U23978 (N_23978,N_23605,N_23755);
nor U23979 (N_23979,N_23729,N_23792);
nor U23980 (N_23980,N_23783,N_23761);
nand U23981 (N_23981,N_23739,N_23646);
xor U23982 (N_23982,N_23771,N_23645);
or U23983 (N_23983,N_23714,N_23780);
nand U23984 (N_23984,N_23728,N_23630);
and U23985 (N_23985,N_23784,N_23648);
nor U23986 (N_23986,N_23607,N_23733);
and U23987 (N_23987,N_23794,N_23606);
nor U23988 (N_23988,N_23777,N_23717);
or U23989 (N_23989,N_23640,N_23782);
or U23990 (N_23990,N_23791,N_23728);
nor U23991 (N_23991,N_23668,N_23795);
and U23992 (N_23992,N_23606,N_23630);
or U23993 (N_23993,N_23750,N_23783);
and U23994 (N_23994,N_23746,N_23710);
nand U23995 (N_23995,N_23729,N_23740);
and U23996 (N_23996,N_23781,N_23634);
nor U23997 (N_23997,N_23612,N_23606);
or U23998 (N_23998,N_23705,N_23749);
nor U23999 (N_23999,N_23738,N_23766);
xnor U24000 (N_24000,N_23845,N_23867);
or U24001 (N_24001,N_23838,N_23913);
nand U24002 (N_24002,N_23939,N_23860);
and U24003 (N_24003,N_23878,N_23820);
or U24004 (N_24004,N_23974,N_23825);
nand U24005 (N_24005,N_23839,N_23888);
or U24006 (N_24006,N_23855,N_23812);
or U24007 (N_24007,N_23854,N_23964);
nor U24008 (N_24008,N_23973,N_23962);
nor U24009 (N_24009,N_23940,N_23995);
nor U24010 (N_24010,N_23906,N_23886);
or U24011 (N_24011,N_23941,N_23903);
xor U24012 (N_24012,N_23925,N_23975);
xnor U24013 (N_24013,N_23834,N_23880);
xor U24014 (N_24014,N_23923,N_23947);
and U24015 (N_24015,N_23905,N_23840);
nor U24016 (N_24016,N_23817,N_23891);
and U24017 (N_24017,N_23909,N_23896);
and U24018 (N_24018,N_23898,N_23857);
xnor U24019 (N_24019,N_23811,N_23800);
nand U24020 (N_24020,N_23980,N_23966);
nor U24021 (N_24021,N_23881,N_23833);
xnor U24022 (N_24022,N_23977,N_23885);
or U24023 (N_24023,N_23927,N_23872);
and U24024 (N_24024,N_23986,N_23951);
nand U24025 (N_24025,N_23979,N_23907);
nor U24026 (N_24026,N_23814,N_23876);
nand U24027 (N_24027,N_23931,N_23852);
or U24028 (N_24028,N_23937,N_23959);
xor U24029 (N_24029,N_23849,N_23868);
and U24030 (N_24030,N_23989,N_23978);
nand U24031 (N_24031,N_23908,N_23967);
xnor U24032 (N_24032,N_23809,N_23869);
and U24033 (N_24033,N_23998,N_23954);
xor U24034 (N_24034,N_23884,N_23853);
or U24035 (N_24035,N_23870,N_23938);
nor U24036 (N_24036,N_23890,N_23803);
nor U24037 (N_24037,N_23836,N_23922);
and U24038 (N_24038,N_23851,N_23960);
xnor U24039 (N_24039,N_23976,N_23987);
nand U24040 (N_24040,N_23879,N_23985);
or U24041 (N_24041,N_23994,N_23988);
nor U24042 (N_24042,N_23883,N_23900);
nand U24043 (N_24043,N_23972,N_23917);
xor U24044 (N_24044,N_23984,N_23861);
or U24045 (N_24045,N_23970,N_23807);
or U24046 (N_24046,N_23919,N_23821);
and U24047 (N_24047,N_23958,N_23929);
nand U24048 (N_24048,N_23841,N_23859);
and U24049 (N_24049,N_23918,N_23802);
or U24050 (N_24050,N_23950,N_23945);
or U24051 (N_24051,N_23952,N_23862);
or U24052 (N_24052,N_23949,N_23850);
nor U24053 (N_24053,N_23948,N_23889);
xnor U24054 (N_24054,N_23819,N_23961);
and U24055 (N_24055,N_23875,N_23921);
or U24056 (N_24056,N_23813,N_23893);
xnor U24057 (N_24057,N_23865,N_23806);
xor U24058 (N_24058,N_23955,N_23932);
or U24059 (N_24059,N_23804,N_23944);
nand U24060 (N_24060,N_23946,N_23963);
and U24061 (N_24061,N_23904,N_23933);
and U24062 (N_24062,N_23990,N_23887);
nor U24063 (N_24063,N_23824,N_23801);
nor U24064 (N_24064,N_23926,N_23936);
xnor U24065 (N_24065,N_23842,N_23835);
and U24066 (N_24066,N_23829,N_23895);
nand U24067 (N_24067,N_23816,N_23902);
and U24068 (N_24068,N_23928,N_23826);
nand U24069 (N_24069,N_23956,N_23877);
or U24070 (N_24070,N_23848,N_23957);
nor U24071 (N_24071,N_23847,N_23912);
nand U24072 (N_24072,N_23874,N_23943);
or U24073 (N_24073,N_23996,N_23942);
and U24074 (N_24074,N_23914,N_23846);
or U24075 (N_24075,N_23882,N_23993);
nand U24076 (N_24076,N_23856,N_23843);
nand U24077 (N_24077,N_23873,N_23915);
nor U24078 (N_24078,N_23828,N_23892);
and U24079 (N_24079,N_23832,N_23837);
xnor U24080 (N_24080,N_23911,N_23805);
and U24081 (N_24081,N_23991,N_23864);
or U24082 (N_24082,N_23858,N_23815);
nand U24083 (N_24083,N_23901,N_23844);
xnor U24084 (N_24084,N_23999,N_23823);
and U24085 (N_24085,N_23808,N_23982);
or U24086 (N_24086,N_23866,N_23924);
xnor U24087 (N_24087,N_23863,N_23810);
or U24088 (N_24088,N_23934,N_23968);
or U24089 (N_24089,N_23871,N_23822);
or U24090 (N_24090,N_23916,N_23935);
xor U24091 (N_24091,N_23953,N_23981);
or U24092 (N_24092,N_23830,N_23965);
or U24093 (N_24093,N_23894,N_23818);
nand U24094 (N_24094,N_23899,N_23897);
and U24095 (N_24095,N_23910,N_23971);
xor U24096 (N_24096,N_23983,N_23831);
and U24097 (N_24097,N_23930,N_23920);
nor U24098 (N_24098,N_23827,N_23997);
xor U24099 (N_24099,N_23992,N_23969);
or U24100 (N_24100,N_23953,N_23894);
or U24101 (N_24101,N_23961,N_23905);
nand U24102 (N_24102,N_23998,N_23973);
or U24103 (N_24103,N_23945,N_23944);
nor U24104 (N_24104,N_23926,N_23881);
and U24105 (N_24105,N_23818,N_23865);
nand U24106 (N_24106,N_23886,N_23833);
xor U24107 (N_24107,N_23977,N_23836);
nand U24108 (N_24108,N_23948,N_23907);
nor U24109 (N_24109,N_23819,N_23805);
and U24110 (N_24110,N_23909,N_23875);
nand U24111 (N_24111,N_23839,N_23950);
xor U24112 (N_24112,N_23914,N_23986);
nor U24113 (N_24113,N_23863,N_23803);
nor U24114 (N_24114,N_23990,N_23876);
nor U24115 (N_24115,N_23932,N_23919);
or U24116 (N_24116,N_23863,N_23927);
nor U24117 (N_24117,N_23824,N_23888);
nor U24118 (N_24118,N_23991,N_23931);
xnor U24119 (N_24119,N_23915,N_23800);
or U24120 (N_24120,N_23938,N_23906);
and U24121 (N_24121,N_23816,N_23945);
or U24122 (N_24122,N_23821,N_23909);
nor U24123 (N_24123,N_23857,N_23831);
nor U24124 (N_24124,N_23803,N_23848);
nor U24125 (N_24125,N_23992,N_23821);
nor U24126 (N_24126,N_23837,N_23812);
nor U24127 (N_24127,N_23835,N_23826);
nor U24128 (N_24128,N_23877,N_23804);
xor U24129 (N_24129,N_23881,N_23945);
or U24130 (N_24130,N_23982,N_23936);
nand U24131 (N_24131,N_23990,N_23890);
nor U24132 (N_24132,N_23885,N_23924);
and U24133 (N_24133,N_23828,N_23849);
xor U24134 (N_24134,N_23856,N_23944);
nand U24135 (N_24135,N_23862,N_23993);
xor U24136 (N_24136,N_23801,N_23996);
nor U24137 (N_24137,N_23851,N_23878);
xnor U24138 (N_24138,N_23963,N_23879);
xnor U24139 (N_24139,N_23884,N_23831);
nor U24140 (N_24140,N_23884,N_23843);
or U24141 (N_24141,N_23861,N_23934);
and U24142 (N_24142,N_23850,N_23800);
xnor U24143 (N_24143,N_23975,N_23893);
nor U24144 (N_24144,N_23979,N_23919);
xnor U24145 (N_24145,N_23982,N_23938);
and U24146 (N_24146,N_23820,N_23814);
nand U24147 (N_24147,N_23986,N_23963);
and U24148 (N_24148,N_23803,N_23943);
and U24149 (N_24149,N_23977,N_23894);
nor U24150 (N_24150,N_23989,N_23955);
or U24151 (N_24151,N_23843,N_23828);
or U24152 (N_24152,N_23849,N_23809);
and U24153 (N_24153,N_23969,N_23837);
or U24154 (N_24154,N_23888,N_23925);
nand U24155 (N_24155,N_23852,N_23929);
nand U24156 (N_24156,N_23825,N_23887);
or U24157 (N_24157,N_23866,N_23877);
nand U24158 (N_24158,N_23931,N_23975);
nor U24159 (N_24159,N_23984,N_23835);
nor U24160 (N_24160,N_23904,N_23932);
or U24161 (N_24161,N_23960,N_23886);
and U24162 (N_24162,N_23848,N_23903);
nor U24163 (N_24163,N_23995,N_23968);
and U24164 (N_24164,N_23939,N_23952);
nand U24165 (N_24165,N_23857,N_23963);
or U24166 (N_24166,N_23914,N_23826);
nand U24167 (N_24167,N_23906,N_23860);
xnor U24168 (N_24168,N_23943,N_23994);
nor U24169 (N_24169,N_23806,N_23842);
and U24170 (N_24170,N_23803,N_23947);
and U24171 (N_24171,N_23972,N_23944);
nand U24172 (N_24172,N_23830,N_23906);
and U24173 (N_24173,N_23804,N_23808);
nor U24174 (N_24174,N_23802,N_23904);
or U24175 (N_24175,N_23996,N_23848);
xor U24176 (N_24176,N_23880,N_23809);
xor U24177 (N_24177,N_23857,N_23813);
or U24178 (N_24178,N_23875,N_23920);
nand U24179 (N_24179,N_23869,N_23995);
nor U24180 (N_24180,N_23949,N_23892);
nor U24181 (N_24181,N_23942,N_23801);
or U24182 (N_24182,N_23864,N_23993);
or U24183 (N_24183,N_23949,N_23958);
or U24184 (N_24184,N_23826,N_23801);
nand U24185 (N_24185,N_23947,N_23936);
and U24186 (N_24186,N_23819,N_23946);
or U24187 (N_24187,N_23835,N_23992);
nor U24188 (N_24188,N_23966,N_23951);
xor U24189 (N_24189,N_23863,N_23838);
xor U24190 (N_24190,N_23831,N_23937);
xor U24191 (N_24191,N_23858,N_23940);
or U24192 (N_24192,N_23848,N_23994);
nand U24193 (N_24193,N_23855,N_23960);
or U24194 (N_24194,N_23932,N_23949);
nand U24195 (N_24195,N_23852,N_23937);
xor U24196 (N_24196,N_23920,N_23941);
nor U24197 (N_24197,N_23859,N_23915);
and U24198 (N_24198,N_23895,N_23907);
nor U24199 (N_24199,N_23949,N_23838);
nand U24200 (N_24200,N_24011,N_24074);
and U24201 (N_24201,N_24004,N_24164);
and U24202 (N_24202,N_24145,N_24064);
or U24203 (N_24203,N_24080,N_24195);
or U24204 (N_24204,N_24075,N_24028);
and U24205 (N_24205,N_24069,N_24143);
or U24206 (N_24206,N_24078,N_24012);
xor U24207 (N_24207,N_24108,N_24016);
and U24208 (N_24208,N_24156,N_24155);
xnor U24209 (N_24209,N_24100,N_24039);
or U24210 (N_24210,N_24045,N_24049);
and U24211 (N_24211,N_24068,N_24112);
or U24212 (N_24212,N_24190,N_24029);
xnor U24213 (N_24213,N_24042,N_24082);
and U24214 (N_24214,N_24087,N_24144);
nor U24215 (N_24215,N_24017,N_24110);
and U24216 (N_24216,N_24172,N_24111);
or U24217 (N_24217,N_24187,N_24133);
or U24218 (N_24218,N_24181,N_24173);
nand U24219 (N_24219,N_24095,N_24124);
nor U24220 (N_24220,N_24003,N_24109);
and U24221 (N_24221,N_24128,N_24114);
nand U24222 (N_24222,N_24047,N_24053);
and U24223 (N_24223,N_24138,N_24198);
xnor U24224 (N_24224,N_24113,N_24127);
nor U24225 (N_24225,N_24035,N_24005);
xor U24226 (N_24226,N_24159,N_24121);
nor U24227 (N_24227,N_24062,N_24022);
xnor U24228 (N_24228,N_24169,N_24158);
nand U24229 (N_24229,N_24160,N_24120);
xor U24230 (N_24230,N_24186,N_24140);
nand U24231 (N_24231,N_24076,N_24085);
nor U24232 (N_24232,N_24021,N_24048);
nor U24233 (N_24233,N_24034,N_24088);
or U24234 (N_24234,N_24197,N_24177);
xor U24235 (N_24235,N_24031,N_24125);
xnor U24236 (N_24236,N_24036,N_24052);
nor U24237 (N_24237,N_24098,N_24107);
xor U24238 (N_24238,N_24189,N_24072);
xor U24239 (N_24239,N_24063,N_24084);
and U24240 (N_24240,N_24077,N_24009);
or U24241 (N_24241,N_24055,N_24086);
nand U24242 (N_24242,N_24105,N_24101);
or U24243 (N_24243,N_24050,N_24083);
nor U24244 (N_24244,N_24175,N_24115);
and U24245 (N_24245,N_24196,N_24043);
xnor U24246 (N_24246,N_24081,N_24103);
nor U24247 (N_24247,N_24058,N_24135);
nor U24248 (N_24248,N_24019,N_24157);
xnor U24249 (N_24249,N_24153,N_24185);
xnor U24250 (N_24250,N_24129,N_24010);
xor U24251 (N_24251,N_24079,N_24091);
xor U24252 (N_24252,N_24023,N_24054);
and U24253 (N_24253,N_24027,N_24066);
xor U24254 (N_24254,N_24191,N_24166);
nor U24255 (N_24255,N_24161,N_24178);
xnor U24256 (N_24256,N_24122,N_24030);
or U24257 (N_24257,N_24170,N_24094);
nand U24258 (N_24258,N_24018,N_24152);
or U24259 (N_24259,N_24089,N_24180);
nand U24260 (N_24260,N_24056,N_24041);
and U24261 (N_24261,N_24148,N_24182);
nand U24262 (N_24262,N_24093,N_24174);
and U24263 (N_24263,N_24000,N_24102);
nor U24264 (N_24264,N_24119,N_24193);
nand U24265 (N_24265,N_24199,N_24044);
or U24266 (N_24266,N_24001,N_24131);
and U24267 (N_24267,N_24006,N_24057);
and U24268 (N_24268,N_24014,N_24176);
or U24269 (N_24269,N_24126,N_24188);
nor U24270 (N_24270,N_24020,N_24099);
and U24271 (N_24271,N_24059,N_24130);
and U24272 (N_24272,N_24123,N_24046);
nor U24273 (N_24273,N_24134,N_24008);
nor U24274 (N_24274,N_24092,N_24040);
nor U24275 (N_24275,N_24132,N_24067);
nor U24276 (N_24276,N_24024,N_24179);
nor U24277 (N_24277,N_24032,N_24106);
xor U24278 (N_24278,N_24136,N_24162);
or U24279 (N_24279,N_24071,N_24002);
or U24280 (N_24280,N_24184,N_24147);
or U24281 (N_24281,N_24192,N_24168);
or U24282 (N_24282,N_24150,N_24116);
and U24283 (N_24283,N_24151,N_24167);
nor U24284 (N_24284,N_24154,N_24026);
or U24285 (N_24285,N_24097,N_24015);
xnor U24286 (N_24286,N_24194,N_24013);
xor U24287 (N_24287,N_24137,N_24060);
xor U24288 (N_24288,N_24171,N_24070);
nor U24289 (N_24289,N_24061,N_24037);
xor U24290 (N_24290,N_24104,N_24146);
xor U24291 (N_24291,N_24007,N_24163);
or U24292 (N_24292,N_24051,N_24025);
or U24293 (N_24293,N_24141,N_24033);
xnor U24294 (N_24294,N_24073,N_24065);
or U24295 (N_24295,N_24117,N_24096);
nor U24296 (N_24296,N_24165,N_24183);
xor U24297 (N_24297,N_24142,N_24149);
xor U24298 (N_24298,N_24090,N_24038);
nand U24299 (N_24299,N_24139,N_24118);
xor U24300 (N_24300,N_24024,N_24102);
and U24301 (N_24301,N_24109,N_24111);
or U24302 (N_24302,N_24061,N_24087);
nor U24303 (N_24303,N_24186,N_24091);
nand U24304 (N_24304,N_24197,N_24110);
or U24305 (N_24305,N_24013,N_24169);
or U24306 (N_24306,N_24007,N_24067);
nand U24307 (N_24307,N_24018,N_24000);
or U24308 (N_24308,N_24013,N_24030);
xor U24309 (N_24309,N_24037,N_24136);
nor U24310 (N_24310,N_24030,N_24195);
nand U24311 (N_24311,N_24116,N_24074);
and U24312 (N_24312,N_24131,N_24023);
nand U24313 (N_24313,N_24082,N_24096);
and U24314 (N_24314,N_24063,N_24029);
nand U24315 (N_24315,N_24008,N_24121);
nor U24316 (N_24316,N_24055,N_24187);
or U24317 (N_24317,N_24031,N_24027);
and U24318 (N_24318,N_24115,N_24126);
or U24319 (N_24319,N_24188,N_24147);
or U24320 (N_24320,N_24011,N_24066);
nand U24321 (N_24321,N_24042,N_24079);
nand U24322 (N_24322,N_24128,N_24096);
xor U24323 (N_24323,N_24174,N_24037);
nand U24324 (N_24324,N_24129,N_24044);
nor U24325 (N_24325,N_24107,N_24189);
and U24326 (N_24326,N_24182,N_24082);
or U24327 (N_24327,N_24158,N_24009);
nand U24328 (N_24328,N_24180,N_24183);
xnor U24329 (N_24329,N_24018,N_24144);
xnor U24330 (N_24330,N_24027,N_24132);
xnor U24331 (N_24331,N_24002,N_24073);
nand U24332 (N_24332,N_24105,N_24137);
nor U24333 (N_24333,N_24134,N_24193);
or U24334 (N_24334,N_24114,N_24133);
or U24335 (N_24335,N_24111,N_24170);
or U24336 (N_24336,N_24040,N_24008);
or U24337 (N_24337,N_24104,N_24026);
or U24338 (N_24338,N_24006,N_24196);
and U24339 (N_24339,N_24017,N_24010);
or U24340 (N_24340,N_24030,N_24164);
nor U24341 (N_24341,N_24136,N_24093);
xnor U24342 (N_24342,N_24070,N_24196);
xnor U24343 (N_24343,N_24031,N_24047);
and U24344 (N_24344,N_24010,N_24171);
nand U24345 (N_24345,N_24104,N_24140);
xor U24346 (N_24346,N_24191,N_24164);
xor U24347 (N_24347,N_24157,N_24052);
nand U24348 (N_24348,N_24110,N_24014);
nor U24349 (N_24349,N_24080,N_24167);
nand U24350 (N_24350,N_24111,N_24168);
nor U24351 (N_24351,N_24119,N_24105);
xor U24352 (N_24352,N_24149,N_24196);
nand U24353 (N_24353,N_24121,N_24184);
nand U24354 (N_24354,N_24079,N_24098);
and U24355 (N_24355,N_24060,N_24005);
or U24356 (N_24356,N_24144,N_24106);
nor U24357 (N_24357,N_24013,N_24016);
nand U24358 (N_24358,N_24193,N_24049);
nand U24359 (N_24359,N_24087,N_24082);
nand U24360 (N_24360,N_24125,N_24032);
or U24361 (N_24361,N_24097,N_24144);
or U24362 (N_24362,N_24154,N_24072);
nand U24363 (N_24363,N_24198,N_24066);
and U24364 (N_24364,N_24073,N_24192);
nor U24365 (N_24365,N_24187,N_24099);
and U24366 (N_24366,N_24072,N_24089);
and U24367 (N_24367,N_24037,N_24097);
or U24368 (N_24368,N_24036,N_24079);
nand U24369 (N_24369,N_24115,N_24103);
and U24370 (N_24370,N_24155,N_24191);
nor U24371 (N_24371,N_24142,N_24117);
and U24372 (N_24372,N_24102,N_24172);
xor U24373 (N_24373,N_24195,N_24174);
or U24374 (N_24374,N_24145,N_24163);
nand U24375 (N_24375,N_24063,N_24082);
and U24376 (N_24376,N_24163,N_24159);
and U24377 (N_24377,N_24022,N_24150);
xor U24378 (N_24378,N_24031,N_24169);
nand U24379 (N_24379,N_24127,N_24028);
nand U24380 (N_24380,N_24182,N_24146);
xnor U24381 (N_24381,N_24107,N_24012);
nor U24382 (N_24382,N_24161,N_24114);
and U24383 (N_24383,N_24020,N_24045);
nor U24384 (N_24384,N_24104,N_24115);
and U24385 (N_24385,N_24000,N_24136);
or U24386 (N_24386,N_24064,N_24125);
or U24387 (N_24387,N_24028,N_24125);
or U24388 (N_24388,N_24117,N_24055);
nor U24389 (N_24389,N_24155,N_24053);
nand U24390 (N_24390,N_24132,N_24009);
nor U24391 (N_24391,N_24079,N_24109);
xnor U24392 (N_24392,N_24108,N_24074);
nand U24393 (N_24393,N_24040,N_24025);
xnor U24394 (N_24394,N_24014,N_24012);
nand U24395 (N_24395,N_24132,N_24151);
and U24396 (N_24396,N_24168,N_24191);
nor U24397 (N_24397,N_24181,N_24048);
and U24398 (N_24398,N_24050,N_24094);
nor U24399 (N_24399,N_24131,N_24109);
nor U24400 (N_24400,N_24235,N_24339);
nand U24401 (N_24401,N_24383,N_24232);
or U24402 (N_24402,N_24393,N_24336);
xnor U24403 (N_24403,N_24255,N_24386);
and U24404 (N_24404,N_24369,N_24337);
nand U24405 (N_24405,N_24233,N_24372);
and U24406 (N_24406,N_24251,N_24320);
xnor U24407 (N_24407,N_24399,N_24267);
nand U24408 (N_24408,N_24354,N_24273);
xor U24409 (N_24409,N_24329,N_24384);
or U24410 (N_24410,N_24264,N_24396);
nand U24411 (N_24411,N_24395,N_24229);
nand U24412 (N_24412,N_24268,N_24248);
nor U24413 (N_24413,N_24353,N_24388);
or U24414 (N_24414,N_24377,N_24200);
xor U24415 (N_24415,N_24299,N_24340);
or U24416 (N_24416,N_24281,N_24271);
xor U24417 (N_24417,N_24303,N_24231);
or U24418 (N_24418,N_24300,N_24343);
nand U24419 (N_24419,N_24293,N_24208);
xor U24420 (N_24420,N_24269,N_24335);
or U24421 (N_24421,N_24250,N_24366);
nor U24422 (N_24422,N_24297,N_24211);
nand U24423 (N_24423,N_24214,N_24258);
and U24424 (N_24424,N_24280,N_24302);
nor U24425 (N_24425,N_24311,N_24218);
nand U24426 (N_24426,N_24362,N_24202);
nand U24427 (N_24427,N_24242,N_24379);
and U24428 (N_24428,N_24294,N_24350);
and U24429 (N_24429,N_24387,N_24365);
nand U24430 (N_24430,N_24207,N_24334);
and U24431 (N_24431,N_24236,N_24282);
nand U24432 (N_24432,N_24237,N_24381);
or U24433 (N_24433,N_24244,N_24222);
nor U24434 (N_24434,N_24216,N_24241);
nor U24435 (N_24435,N_24260,N_24276);
nor U24436 (N_24436,N_24360,N_24219);
nand U24437 (N_24437,N_24325,N_24278);
or U24438 (N_24438,N_24358,N_24392);
xor U24439 (N_24439,N_24347,N_24368);
xor U24440 (N_24440,N_24304,N_24270);
or U24441 (N_24441,N_24287,N_24367);
or U24442 (N_24442,N_24301,N_24330);
or U24443 (N_24443,N_24221,N_24203);
nand U24444 (N_24444,N_24210,N_24263);
nor U24445 (N_24445,N_24382,N_24246);
or U24446 (N_24446,N_24385,N_24249);
nor U24447 (N_24447,N_24205,N_24213);
or U24448 (N_24448,N_24328,N_24274);
or U24449 (N_24449,N_24341,N_24319);
or U24450 (N_24450,N_24317,N_24361);
or U24451 (N_24451,N_24286,N_24209);
nand U24452 (N_24452,N_24227,N_24228);
xor U24453 (N_24453,N_24310,N_24277);
nand U24454 (N_24454,N_24225,N_24257);
xor U24455 (N_24455,N_24290,N_24363);
and U24456 (N_24456,N_24238,N_24373);
nor U24457 (N_24457,N_24344,N_24220);
nor U24458 (N_24458,N_24226,N_24288);
and U24459 (N_24459,N_24215,N_24322);
nor U24460 (N_24460,N_24289,N_24394);
nand U24461 (N_24461,N_24307,N_24239);
nand U24462 (N_24462,N_24259,N_24323);
nand U24463 (N_24463,N_24292,N_24389);
nor U24464 (N_24464,N_24357,N_24275);
or U24465 (N_24465,N_24342,N_24374);
and U24466 (N_24466,N_24245,N_24284);
and U24467 (N_24467,N_24305,N_24291);
xor U24468 (N_24468,N_24391,N_24398);
and U24469 (N_24469,N_24327,N_24397);
and U24470 (N_24470,N_24224,N_24308);
xnor U24471 (N_24471,N_24306,N_24223);
xor U24472 (N_24472,N_24333,N_24313);
and U24473 (N_24473,N_24318,N_24252);
nand U24474 (N_24474,N_24234,N_24378);
nand U24475 (N_24475,N_24262,N_24298);
and U24476 (N_24476,N_24364,N_24261);
nor U24477 (N_24477,N_24375,N_24331);
and U24478 (N_24478,N_24204,N_24326);
or U24479 (N_24479,N_24230,N_24352);
and U24480 (N_24480,N_24266,N_24206);
and U24481 (N_24481,N_24212,N_24295);
nor U24482 (N_24482,N_24283,N_24253);
and U24483 (N_24483,N_24345,N_24324);
xnor U24484 (N_24484,N_24371,N_24321);
nor U24485 (N_24485,N_24316,N_24359);
nand U24486 (N_24486,N_24315,N_24254);
and U24487 (N_24487,N_24351,N_24285);
nor U24488 (N_24488,N_24217,N_24370);
and U24489 (N_24489,N_24332,N_24240);
nand U24490 (N_24490,N_24338,N_24309);
nand U24491 (N_24491,N_24201,N_24256);
nor U24492 (N_24492,N_24348,N_24265);
or U24493 (N_24493,N_24346,N_24376);
or U24494 (N_24494,N_24356,N_24243);
nor U24495 (N_24495,N_24279,N_24314);
nor U24496 (N_24496,N_24312,N_24247);
nor U24497 (N_24497,N_24349,N_24355);
nor U24498 (N_24498,N_24296,N_24380);
nor U24499 (N_24499,N_24390,N_24272);
nor U24500 (N_24500,N_24231,N_24233);
or U24501 (N_24501,N_24224,N_24270);
xnor U24502 (N_24502,N_24396,N_24268);
and U24503 (N_24503,N_24353,N_24227);
nor U24504 (N_24504,N_24322,N_24286);
xor U24505 (N_24505,N_24376,N_24394);
xnor U24506 (N_24506,N_24354,N_24366);
and U24507 (N_24507,N_24301,N_24262);
xnor U24508 (N_24508,N_24230,N_24399);
xnor U24509 (N_24509,N_24374,N_24399);
nand U24510 (N_24510,N_24288,N_24246);
or U24511 (N_24511,N_24322,N_24241);
nand U24512 (N_24512,N_24363,N_24387);
nor U24513 (N_24513,N_24346,N_24210);
nor U24514 (N_24514,N_24376,N_24348);
nand U24515 (N_24515,N_24374,N_24322);
and U24516 (N_24516,N_24362,N_24381);
or U24517 (N_24517,N_24247,N_24278);
or U24518 (N_24518,N_24316,N_24272);
or U24519 (N_24519,N_24256,N_24261);
or U24520 (N_24520,N_24270,N_24234);
nand U24521 (N_24521,N_24376,N_24207);
or U24522 (N_24522,N_24378,N_24359);
and U24523 (N_24523,N_24382,N_24381);
xnor U24524 (N_24524,N_24273,N_24299);
nor U24525 (N_24525,N_24301,N_24343);
xor U24526 (N_24526,N_24355,N_24338);
nand U24527 (N_24527,N_24318,N_24339);
xnor U24528 (N_24528,N_24316,N_24391);
nor U24529 (N_24529,N_24322,N_24356);
xnor U24530 (N_24530,N_24238,N_24330);
nor U24531 (N_24531,N_24246,N_24323);
xor U24532 (N_24532,N_24372,N_24255);
nand U24533 (N_24533,N_24231,N_24274);
nor U24534 (N_24534,N_24235,N_24225);
nand U24535 (N_24535,N_24231,N_24339);
xnor U24536 (N_24536,N_24340,N_24338);
or U24537 (N_24537,N_24317,N_24299);
nor U24538 (N_24538,N_24336,N_24252);
nor U24539 (N_24539,N_24225,N_24332);
and U24540 (N_24540,N_24366,N_24389);
xor U24541 (N_24541,N_24205,N_24208);
nor U24542 (N_24542,N_24311,N_24277);
nor U24543 (N_24543,N_24372,N_24278);
or U24544 (N_24544,N_24254,N_24318);
and U24545 (N_24545,N_24227,N_24375);
or U24546 (N_24546,N_24326,N_24286);
nor U24547 (N_24547,N_24381,N_24260);
or U24548 (N_24548,N_24347,N_24321);
xnor U24549 (N_24549,N_24218,N_24373);
or U24550 (N_24550,N_24345,N_24249);
nand U24551 (N_24551,N_24266,N_24241);
nor U24552 (N_24552,N_24299,N_24211);
or U24553 (N_24553,N_24315,N_24360);
xor U24554 (N_24554,N_24376,N_24379);
and U24555 (N_24555,N_24317,N_24337);
xor U24556 (N_24556,N_24296,N_24223);
xor U24557 (N_24557,N_24374,N_24358);
nor U24558 (N_24558,N_24243,N_24295);
nor U24559 (N_24559,N_24323,N_24265);
nor U24560 (N_24560,N_24338,N_24335);
nand U24561 (N_24561,N_24290,N_24259);
nor U24562 (N_24562,N_24399,N_24389);
nor U24563 (N_24563,N_24346,N_24204);
or U24564 (N_24564,N_24354,N_24381);
xnor U24565 (N_24565,N_24387,N_24347);
nor U24566 (N_24566,N_24203,N_24298);
and U24567 (N_24567,N_24318,N_24298);
or U24568 (N_24568,N_24375,N_24337);
xnor U24569 (N_24569,N_24315,N_24380);
nor U24570 (N_24570,N_24352,N_24281);
and U24571 (N_24571,N_24240,N_24323);
and U24572 (N_24572,N_24338,N_24351);
nor U24573 (N_24573,N_24312,N_24397);
and U24574 (N_24574,N_24218,N_24274);
or U24575 (N_24575,N_24216,N_24208);
nor U24576 (N_24576,N_24350,N_24257);
or U24577 (N_24577,N_24252,N_24257);
nor U24578 (N_24578,N_24339,N_24264);
xnor U24579 (N_24579,N_24299,N_24246);
xor U24580 (N_24580,N_24296,N_24314);
nand U24581 (N_24581,N_24251,N_24369);
and U24582 (N_24582,N_24200,N_24244);
or U24583 (N_24583,N_24217,N_24203);
nor U24584 (N_24584,N_24228,N_24373);
or U24585 (N_24585,N_24206,N_24369);
xnor U24586 (N_24586,N_24245,N_24307);
nand U24587 (N_24587,N_24311,N_24370);
xor U24588 (N_24588,N_24311,N_24238);
and U24589 (N_24589,N_24385,N_24393);
and U24590 (N_24590,N_24236,N_24235);
nand U24591 (N_24591,N_24379,N_24240);
xnor U24592 (N_24592,N_24251,N_24312);
nor U24593 (N_24593,N_24251,N_24374);
nand U24594 (N_24594,N_24328,N_24252);
nor U24595 (N_24595,N_24253,N_24233);
or U24596 (N_24596,N_24263,N_24358);
nor U24597 (N_24597,N_24242,N_24274);
and U24598 (N_24598,N_24209,N_24229);
nand U24599 (N_24599,N_24371,N_24211);
nor U24600 (N_24600,N_24454,N_24522);
nor U24601 (N_24601,N_24588,N_24483);
nor U24602 (N_24602,N_24582,N_24578);
and U24603 (N_24603,N_24518,N_24587);
or U24604 (N_24604,N_24509,N_24583);
nand U24605 (N_24605,N_24408,N_24428);
or U24606 (N_24606,N_24597,N_24576);
and U24607 (N_24607,N_24598,N_24436);
or U24608 (N_24608,N_24554,N_24534);
nand U24609 (N_24609,N_24555,N_24417);
nor U24610 (N_24610,N_24403,N_24427);
nor U24611 (N_24611,N_24498,N_24482);
xnor U24612 (N_24612,N_24535,N_24574);
or U24613 (N_24613,N_24487,N_24416);
nand U24614 (N_24614,N_24586,N_24438);
and U24615 (N_24615,N_24523,N_24460);
nand U24616 (N_24616,N_24412,N_24435);
and U24617 (N_24617,N_24528,N_24500);
nor U24618 (N_24618,N_24453,N_24508);
nor U24619 (N_24619,N_24567,N_24504);
nand U24620 (N_24620,N_24432,N_24573);
nor U24621 (N_24621,N_24486,N_24451);
nand U24622 (N_24622,N_24414,N_24433);
or U24623 (N_24623,N_24543,N_24514);
or U24624 (N_24624,N_24422,N_24538);
xnor U24625 (N_24625,N_24485,N_24479);
and U24626 (N_24626,N_24564,N_24488);
nand U24627 (N_24627,N_24429,N_24410);
xnor U24628 (N_24628,N_24575,N_24547);
xnor U24629 (N_24629,N_24446,N_24517);
or U24630 (N_24630,N_24584,N_24515);
nor U24631 (N_24631,N_24579,N_24524);
nor U24632 (N_24632,N_24516,N_24476);
nand U24633 (N_24633,N_24466,N_24471);
nor U24634 (N_24634,N_24470,N_24491);
nor U24635 (N_24635,N_24541,N_24565);
nor U24636 (N_24636,N_24566,N_24507);
and U24637 (N_24637,N_24520,N_24420);
xnor U24638 (N_24638,N_24411,N_24569);
or U24639 (N_24639,N_24457,N_24477);
and U24640 (N_24640,N_24594,N_24546);
and U24641 (N_24641,N_24542,N_24404);
or U24642 (N_24642,N_24443,N_24592);
and U24643 (N_24643,N_24513,N_24447);
nand U24644 (N_24644,N_24532,N_24539);
and U24645 (N_24645,N_24556,N_24445);
nor U24646 (N_24646,N_24468,N_24502);
xor U24647 (N_24647,N_24406,N_24440);
nor U24648 (N_24648,N_24490,N_24434);
xor U24649 (N_24649,N_24484,N_24585);
nand U24650 (N_24650,N_24549,N_24595);
nand U24651 (N_24651,N_24455,N_24557);
nand U24652 (N_24652,N_24437,N_24560);
nand U24653 (N_24653,N_24581,N_24444);
and U24654 (N_24654,N_24450,N_24464);
nor U24655 (N_24655,N_24405,N_24577);
or U24656 (N_24656,N_24495,N_24489);
and U24657 (N_24657,N_24596,N_24472);
nor U24658 (N_24658,N_24473,N_24494);
nor U24659 (N_24659,N_24562,N_24525);
xor U24660 (N_24660,N_24481,N_24570);
nor U24661 (N_24661,N_24497,N_24544);
or U24662 (N_24662,N_24469,N_24458);
or U24663 (N_24663,N_24409,N_24423);
nor U24664 (N_24664,N_24492,N_24419);
xor U24665 (N_24665,N_24537,N_24506);
and U24666 (N_24666,N_24529,N_24591);
or U24667 (N_24667,N_24465,N_24449);
nand U24668 (N_24668,N_24467,N_24441);
nand U24669 (N_24669,N_24559,N_24401);
nor U24670 (N_24670,N_24568,N_24563);
and U24671 (N_24671,N_24510,N_24527);
and U24672 (N_24672,N_24462,N_24589);
xnor U24673 (N_24673,N_24499,N_24463);
or U24674 (N_24674,N_24413,N_24421);
nor U24675 (N_24675,N_24580,N_24439);
or U24676 (N_24676,N_24521,N_24550);
or U24677 (N_24677,N_24459,N_24430);
or U24678 (N_24678,N_24526,N_24496);
nor U24679 (N_24679,N_24475,N_24478);
xor U24680 (N_24680,N_24561,N_24548);
nand U24681 (N_24681,N_24511,N_24530);
and U24682 (N_24682,N_24400,N_24402);
nand U24683 (N_24683,N_24558,N_24407);
xnor U24684 (N_24684,N_24426,N_24572);
or U24685 (N_24685,N_24474,N_24461);
or U24686 (N_24686,N_24571,N_24551);
or U24687 (N_24687,N_24590,N_24552);
nor U24688 (N_24688,N_24425,N_24599);
nand U24689 (N_24689,N_24456,N_24480);
and U24690 (N_24690,N_24505,N_24493);
or U24691 (N_24691,N_24424,N_24418);
or U24692 (N_24692,N_24415,N_24531);
and U24693 (N_24693,N_24553,N_24448);
and U24694 (N_24694,N_24452,N_24540);
nand U24695 (N_24695,N_24442,N_24512);
or U24696 (N_24696,N_24593,N_24503);
and U24697 (N_24697,N_24431,N_24536);
xor U24698 (N_24698,N_24501,N_24533);
or U24699 (N_24699,N_24519,N_24545);
or U24700 (N_24700,N_24487,N_24422);
nand U24701 (N_24701,N_24448,N_24420);
and U24702 (N_24702,N_24420,N_24500);
nand U24703 (N_24703,N_24439,N_24434);
or U24704 (N_24704,N_24519,N_24433);
xnor U24705 (N_24705,N_24435,N_24500);
nor U24706 (N_24706,N_24544,N_24549);
nand U24707 (N_24707,N_24410,N_24412);
xnor U24708 (N_24708,N_24529,N_24540);
xor U24709 (N_24709,N_24415,N_24450);
and U24710 (N_24710,N_24455,N_24539);
xor U24711 (N_24711,N_24468,N_24591);
xor U24712 (N_24712,N_24548,N_24545);
xnor U24713 (N_24713,N_24437,N_24413);
or U24714 (N_24714,N_24415,N_24547);
nand U24715 (N_24715,N_24410,N_24544);
nand U24716 (N_24716,N_24557,N_24454);
nor U24717 (N_24717,N_24497,N_24495);
nand U24718 (N_24718,N_24570,N_24437);
or U24719 (N_24719,N_24494,N_24579);
xnor U24720 (N_24720,N_24566,N_24517);
xnor U24721 (N_24721,N_24484,N_24413);
and U24722 (N_24722,N_24583,N_24421);
nor U24723 (N_24723,N_24457,N_24503);
nand U24724 (N_24724,N_24490,N_24431);
xor U24725 (N_24725,N_24468,N_24595);
or U24726 (N_24726,N_24413,N_24585);
nor U24727 (N_24727,N_24501,N_24518);
xnor U24728 (N_24728,N_24583,N_24452);
nand U24729 (N_24729,N_24415,N_24423);
xnor U24730 (N_24730,N_24514,N_24454);
xnor U24731 (N_24731,N_24467,N_24593);
nand U24732 (N_24732,N_24527,N_24456);
and U24733 (N_24733,N_24487,N_24490);
nand U24734 (N_24734,N_24470,N_24530);
xor U24735 (N_24735,N_24501,N_24492);
nand U24736 (N_24736,N_24409,N_24471);
nand U24737 (N_24737,N_24487,N_24409);
nor U24738 (N_24738,N_24566,N_24496);
nand U24739 (N_24739,N_24599,N_24513);
xnor U24740 (N_24740,N_24588,N_24503);
nand U24741 (N_24741,N_24463,N_24582);
or U24742 (N_24742,N_24486,N_24598);
xor U24743 (N_24743,N_24409,N_24528);
nand U24744 (N_24744,N_24435,N_24495);
xnor U24745 (N_24745,N_24496,N_24567);
or U24746 (N_24746,N_24528,N_24425);
nand U24747 (N_24747,N_24549,N_24498);
and U24748 (N_24748,N_24419,N_24489);
nor U24749 (N_24749,N_24544,N_24567);
and U24750 (N_24750,N_24415,N_24448);
and U24751 (N_24751,N_24412,N_24439);
nor U24752 (N_24752,N_24436,N_24565);
xor U24753 (N_24753,N_24527,N_24571);
nand U24754 (N_24754,N_24420,N_24414);
xnor U24755 (N_24755,N_24492,N_24438);
or U24756 (N_24756,N_24577,N_24423);
and U24757 (N_24757,N_24562,N_24456);
and U24758 (N_24758,N_24535,N_24487);
nor U24759 (N_24759,N_24408,N_24580);
nor U24760 (N_24760,N_24536,N_24492);
xnor U24761 (N_24761,N_24403,N_24469);
nor U24762 (N_24762,N_24415,N_24469);
and U24763 (N_24763,N_24471,N_24533);
nor U24764 (N_24764,N_24461,N_24501);
nor U24765 (N_24765,N_24487,N_24520);
and U24766 (N_24766,N_24515,N_24453);
nand U24767 (N_24767,N_24543,N_24562);
xnor U24768 (N_24768,N_24407,N_24483);
and U24769 (N_24769,N_24478,N_24412);
and U24770 (N_24770,N_24512,N_24474);
nor U24771 (N_24771,N_24476,N_24534);
nand U24772 (N_24772,N_24421,N_24471);
or U24773 (N_24773,N_24408,N_24406);
and U24774 (N_24774,N_24518,N_24450);
nand U24775 (N_24775,N_24530,N_24437);
xnor U24776 (N_24776,N_24578,N_24536);
or U24777 (N_24777,N_24444,N_24542);
nor U24778 (N_24778,N_24524,N_24420);
nor U24779 (N_24779,N_24423,N_24447);
nor U24780 (N_24780,N_24549,N_24539);
and U24781 (N_24781,N_24411,N_24509);
and U24782 (N_24782,N_24579,N_24594);
or U24783 (N_24783,N_24407,N_24417);
and U24784 (N_24784,N_24406,N_24407);
and U24785 (N_24785,N_24406,N_24448);
xor U24786 (N_24786,N_24599,N_24499);
or U24787 (N_24787,N_24453,N_24542);
or U24788 (N_24788,N_24539,N_24559);
or U24789 (N_24789,N_24496,N_24483);
nand U24790 (N_24790,N_24457,N_24464);
nand U24791 (N_24791,N_24573,N_24598);
nand U24792 (N_24792,N_24400,N_24511);
and U24793 (N_24793,N_24519,N_24422);
and U24794 (N_24794,N_24545,N_24523);
nand U24795 (N_24795,N_24410,N_24456);
nand U24796 (N_24796,N_24425,N_24435);
and U24797 (N_24797,N_24428,N_24463);
and U24798 (N_24798,N_24467,N_24527);
or U24799 (N_24799,N_24583,N_24515);
xnor U24800 (N_24800,N_24723,N_24706);
nand U24801 (N_24801,N_24780,N_24749);
xnor U24802 (N_24802,N_24781,N_24758);
nand U24803 (N_24803,N_24601,N_24739);
and U24804 (N_24804,N_24612,N_24641);
and U24805 (N_24805,N_24752,N_24707);
and U24806 (N_24806,N_24618,N_24667);
or U24807 (N_24807,N_24740,N_24684);
and U24808 (N_24808,N_24760,N_24661);
xnor U24809 (N_24809,N_24726,N_24708);
and U24810 (N_24810,N_24794,N_24750);
xnor U24811 (N_24811,N_24621,N_24729);
xor U24812 (N_24812,N_24650,N_24738);
and U24813 (N_24813,N_24763,N_24784);
nor U24814 (N_24814,N_24751,N_24659);
nor U24815 (N_24815,N_24744,N_24608);
nor U24816 (N_24816,N_24776,N_24685);
and U24817 (N_24817,N_24725,N_24690);
xor U24818 (N_24818,N_24732,N_24673);
and U24819 (N_24819,N_24769,N_24619);
nor U24820 (N_24820,N_24761,N_24640);
xnor U24821 (N_24821,N_24622,N_24778);
nand U24822 (N_24822,N_24644,N_24658);
nand U24823 (N_24823,N_24754,N_24671);
xnor U24824 (N_24824,N_24787,N_24742);
nor U24825 (N_24825,N_24745,N_24747);
and U24826 (N_24826,N_24623,N_24722);
and U24827 (N_24827,N_24678,N_24616);
or U24828 (N_24828,N_24755,N_24771);
or U24829 (N_24829,N_24788,N_24798);
and U24830 (N_24830,N_24773,N_24696);
or U24831 (N_24831,N_24736,N_24688);
or U24832 (N_24832,N_24721,N_24648);
nor U24833 (N_24833,N_24686,N_24605);
or U24834 (N_24834,N_24692,N_24613);
and U24835 (N_24835,N_24663,N_24624);
or U24836 (N_24836,N_24772,N_24765);
xnor U24837 (N_24837,N_24774,N_24600);
xor U24838 (N_24838,N_24674,N_24665);
nor U24839 (N_24839,N_24793,N_24630);
and U24840 (N_24840,N_24629,N_24697);
or U24841 (N_24841,N_24651,N_24681);
nand U24842 (N_24842,N_24711,N_24639);
nand U24843 (N_24843,N_24636,N_24702);
or U24844 (N_24844,N_24786,N_24727);
xor U24845 (N_24845,N_24757,N_24677);
or U24846 (N_24846,N_24767,N_24660);
xor U24847 (N_24847,N_24657,N_24716);
nor U24848 (N_24848,N_24625,N_24637);
nand U24849 (N_24849,N_24743,N_24766);
nand U24850 (N_24850,N_24632,N_24642);
and U24851 (N_24851,N_24705,N_24741);
nand U24852 (N_24852,N_24689,N_24714);
and U24853 (N_24853,N_24775,N_24628);
and U24854 (N_24854,N_24762,N_24730);
nand U24855 (N_24855,N_24675,N_24609);
nand U24856 (N_24856,N_24728,N_24734);
and U24857 (N_24857,N_24668,N_24679);
xnor U24858 (N_24858,N_24709,N_24790);
nor U24859 (N_24859,N_24614,N_24626);
xor U24860 (N_24860,N_24764,N_24654);
xor U24861 (N_24861,N_24649,N_24796);
xor U24862 (N_24862,N_24615,N_24627);
xnor U24863 (N_24863,N_24735,N_24759);
nor U24864 (N_24864,N_24791,N_24704);
nand U24865 (N_24865,N_24653,N_24672);
or U24866 (N_24866,N_24610,N_24724);
nor U24867 (N_24867,N_24617,N_24646);
nor U24868 (N_24868,N_24737,N_24701);
nor U24869 (N_24869,N_24797,N_24785);
nand U24870 (N_24870,N_24795,N_24713);
or U24871 (N_24871,N_24783,N_24703);
and U24872 (N_24872,N_24733,N_24638);
and U24873 (N_24873,N_24682,N_24603);
nor U24874 (N_24874,N_24756,N_24669);
xor U24875 (N_24875,N_24643,N_24606);
xnor U24876 (N_24876,N_24645,N_24695);
nor U24877 (N_24877,N_24731,N_24700);
nand U24878 (N_24878,N_24770,N_24698);
nor U24879 (N_24879,N_24715,N_24631);
or U24880 (N_24880,N_24604,N_24691);
nor U24881 (N_24881,N_24634,N_24693);
xor U24882 (N_24882,N_24717,N_24719);
and U24883 (N_24883,N_24718,N_24666);
xnor U24884 (N_24884,N_24712,N_24664);
or U24885 (N_24885,N_24792,N_24670);
xor U24886 (N_24886,N_24687,N_24782);
and U24887 (N_24887,N_24748,N_24720);
and U24888 (N_24888,N_24779,N_24676);
nor U24889 (N_24889,N_24607,N_24647);
and U24890 (N_24890,N_24635,N_24662);
and U24891 (N_24891,N_24789,N_24710);
xnor U24892 (N_24892,N_24777,N_24753);
xnor U24893 (N_24893,N_24611,N_24656);
and U24894 (N_24894,N_24768,N_24746);
nor U24895 (N_24895,N_24620,N_24683);
or U24896 (N_24896,N_24694,N_24633);
nor U24897 (N_24897,N_24799,N_24655);
nand U24898 (N_24898,N_24652,N_24680);
xor U24899 (N_24899,N_24602,N_24699);
or U24900 (N_24900,N_24622,N_24768);
nand U24901 (N_24901,N_24676,N_24729);
xnor U24902 (N_24902,N_24644,N_24674);
nor U24903 (N_24903,N_24724,N_24629);
xor U24904 (N_24904,N_24673,N_24759);
nand U24905 (N_24905,N_24650,N_24622);
nor U24906 (N_24906,N_24608,N_24633);
or U24907 (N_24907,N_24675,N_24746);
nor U24908 (N_24908,N_24752,N_24613);
nor U24909 (N_24909,N_24723,N_24729);
or U24910 (N_24910,N_24758,N_24668);
and U24911 (N_24911,N_24649,N_24680);
nor U24912 (N_24912,N_24764,N_24777);
nand U24913 (N_24913,N_24606,N_24620);
and U24914 (N_24914,N_24755,N_24734);
and U24915 (N_24915,N_24678,N_24629);
or U24916 (N_24916,N_24666,N_24631);
nand U24917 (N_24917,N_24788,N_24617);
xor U24918 (N_24918,N_24795,N_24694);
and U24919 (N_24919,N_24612,N_24780);
and U24920 (N_24920,N_24656,N_24690);
xor U24921 (N_24921,N_24765,N_24739);
nor U24922 (N_24922,N_24658,N_24673);
or U24923 (N_24923,N_24613,N_24705);
nand U24924 (N_24924,N_24749,N_24769);
xnor U24925 (N_24925,N_24742,N_24717);
xor U24926 (N_24926,N_24639,N_24758);
nor U24927 (N_24927,N_24771,N_24712);
and U24928 (N_24928,N_24696,N_24723);
and U24929 (N_24929,N_24701,N_24650);
nor U24930 (N_24930,N_24719,N_24657);
nor U24931 (N_24931,N_24666,N_24695);
xnor U24932 (N_24932,N_24654,N_24629);
nand U24933 (N_24933,N_24764,N_24705);
or U24934 (N_24934,N_24799,N_24724);
nor U24935 (N_24935,N_24758,N_24619);
or U24936 (N_24936,N_24742,N_24706);
nor U24937 (N_24937,N_24777,N_24639);
xnor U24938 (N_24938,N_24624,N_24644);
xnor U24939 (N_24939,N_24605,N_24609);
and U24940 (N_24940,N_24618,N_24615);
or U24941 (N_24941,N_24751,N_24799);
xor U24942 (N_24942,N_24679,N_24721);
xor U24943 (N_24943,N_24700,N_24728);
nor U24944 (N_24944,N_24602,N_24659);
and U24945 (N_24945,N_24725,N_24766);
xor U24946 (N_24946,N_24772,N_24761);
nor U24947 (N_24947,N_24768,N_24683);
nor U24948 (N_24948,N_24705,N_24666);
nand U24949 (N_24949,N_24655,N_24783);
nor U24950 (N_24950,N_24678,N_24675);
nor U24951 (N_24951,N_24649,N_24628);
or U24952 (N_24952,N_24640,N_24717);
nand U24953 (N_24953,N_24722,N_24645);
or U24954 (N_24954,N_24643,N_24642);
xor U24955 (N_24955,N_24661,N_24748);
nand U24956 (N_24956,N_24780,N_24766);
nand U24957 (N_24957,N_24644,N_24669);
nand U24958 (N_24958,N_24708,N_24675);
or U24959 (N_24959,N_24624,N_24761);
and U24960 (N_24960,N_24608,N_24792);
and U24961 (N_24961,N_24760,N_24701);
xnor U24962 (N_24962,N_24770,N_24732);
nand U24963 (N_24963,N_24627,N_24798);
or U24964 (N_24964,N_24680,N_24679);
and U24965 (N_24965,N_24609,N_24749);
nor U24966 (N_24966,N_24647,N_24633);
nand U24967 (N_24967,N_24778,N_24656);
xor U24968 (N_24968,N_24727,N_24749);
xnor U24969 (N_24969,N_24735,N_24752);
nand U24970 (N_24970,N_24724,N_24757);
and U24971 (N_24971,N_24645,N_24633);
or U24972 (N_24972,N_24617,N_24651);
nand U24973 (N_24973,N_24621,N_24740);
or U24974 (N_24974,N_24639,N_24642);
or U24975 (N_24975,N_24752,N_24665);
xnor U24976 (N_24976,N_24710,N_24650);
and U24977 (N_24977,N_24745,N_24641);
and U24978 (N_24978,N_24694,N_24651);
and U24979 (N_24979,N_24662,N_24661);
and U24980 (N_24980,N_24628,N_24778);
or U24981 (N_24981,N_24709,N_24655);
xnor U24982 (N_24982,N_24635,N_24719);
nor U24983 (N_24983,N_24640,N_24617);
nor U24984 (N_24984,N_24710,N_24777);
nor U24985 (N_24985,N_24671,N_24659);
nor U24986 (N_24986,N_24773,N_24754);
and U24987 (N_24987,N_24699,N_24658);
nor U24988 (N_24988,N_24682,N_24654);
or U24989 (N_24989,N_24622,N_24647);
nor U24990 (N_24990,N_24657,N_24647);
or U24991 (N_24991,N_24670,N_24759);
or U24992 (N_24992,N_24676,N_24636);
and U24993 (N_24993,N_24637,N_24670);
nand U24994 (N_24994,N_24741,N_24708);
nor U24995 (N_24995,N_24794,N_24753);
nor U24996 (N_24996,N_24617,N_24729);
or U24997 (N_24997,N_24715,N_24738);
and U24998 (N_24998,N_24637,N_24629);
xnor U24999 (N_24999,N_24655,N_24787);
or U25000 (N_25000,N_24878,N_24945);
or U25001 (N_25001,N_24994,N_24966);
xnor U25002 (N_25002,N_24956,N_24926);
nand U25003 (N_25003,N_24979,N_24839);
nand U25004 (N_25004,N_24897,N_24901);
nor U25005 (N_25005,N_24815,N_24861);
or U25006 (N_25006,N_24944,N_24971);
nor U25007 (N_25007,N_24936,N_24942);
nor U25008 (N_25008,N_24943,N_24987);
nand U25009 (N_25009,N_24932,N_24876);
or U25010 (N_25010,N_24921,N_24875);
nand U25011 (N_25011,N_24894,N_24992);
and U25012 (N_25012,N_24978,N_24833);
or U25013 (N_25013,N_24968,N_24852);
nand U25014 (N_25014,N_24845,N_24883);
xor U25015 (N_25015,N_24811,N_24920);
xnor U25016 (N_25016,N_24870,N_24804);
nand U25017 (N_25017,N_24985,N_24820);
xnor U25018 (N_25018,N_24827,N_24910);
xor U25019 (N_25019,N_24832,N_24931);
and U25020 (N_25020,N_24958,N_24892);
and U25021 (N_25021,N_24840,N_24850);
xnor U25022 (N_25022,N_24882,N_24948);
xnor U25023 (N_25023,N_24924,N_24906);
and U25024 (N_25024,N_24998,N_24893);
or U25025 (N_25025,N_24961,N_24904);
or U25026 (N_25026,N_24866,N_24805);
xor U25027 (N_25027,N_24939,N_24843);
or U25028 (N_25028,N_24813,N_24929);
and U25029 (N_25029,N_24928,N_24844);
and U25030 (N_25030,N_24808,N_24916);
nor U25031 (N_25031,N_24884,N_24889);
or U25032 (N_25032,N_24886,N_24809);
xnor U25033 (N_25033,N_24940,N_24849);
nand U25034 (N_25034,N_24988,N_24887);
nand U25035 (N_25035,N_24825,N_24934);
or U25036 (N_25036,N_24935,N_24829);
xor U25037 (N_25037,N_24902,N_24818);
xnor U25038 (N_25038,N_24907,N_24891);
nand U25039 (N_25039,N_24999,N_24888);
and U25040 (N_25040,N_24819,N_24930);
nand U25041 (N_25041,N_24895,N_24857);
xor U25042 (N_25042,N_24983,N_24947);
xor U25043 (N_25043,N_24989,N_24970);
xor U25044 (N_25044,N_24856,N_24927);
xnor U25045 (N_25045,N_24836,N_24933);
or U25046 (N_25046,N_24898,N_24802);
and U25047 (N_25047,N_24858,N_24880);
nor U25048 (N_25048,N_24853,N_24810);
nor U25049 (N_25049,N_24997,N_24967);
nand U25050 (N_25050,N_24976,N_24990);
nor U25051 (N_25051,N_24879,N_24848);
and U25052 (N_25052,N_24919,N_24846);
nor U25053 (N_25053,N_24982,N_24964);
nand U25054 (N_25054,N_24915,N_24925);
and U25055 (N_25055,N_24957,N_24823);
xnor U25056 (N_25056,N_24995,N_24841);
nor U25057 (N_25057,N_24900,N_24980);
nor U25058 (N_25058,N_24868,N_24965);
or U25059 (N_25059,N_24969,N_24862);
or U25060 (N_25060,N_24996,N_24834);
xor U25061 (N_25061,N_24885,N_24812);
nand U25062 (N_25062,N_24950,N_24975);
and U25063 (N_25063,N_24984,N_24896);
nor U25064 (N_25064,N_24923,N_24864);
nand U25065 (N_25065,N_24801,N_24960);
or U25066 (N_25066,N_24986,N_24822);
nand U25067 (N_25067,N_24993,N_24949);
xor U25068 (N_25068,N_24973,N_24831);
nand U25069 (N_25069,N_24828,N_24952);
xnor U25070 (N_25070,N_24817,N_24977);
nor U25071 (N_25071,N_24873,N_24821);
nor U25072 (N_25072,N_24838,N_24918);
or U25073 (N_25073,N_24826,N_24872);
nand U25074 (N_25074,N_24913,N_24869);
nor U25075 (N_25075,N_24814,N_24972);
nand U25076 (N_25076,N_24954,N_24855);
and U25077 (N_25077,N_24865,N_24800);
and U25078 (N_25078,N_24938,N_24991);
xor U25079 (N_25079,N_24816,N_24963);
nand U25080 (N_25080,N_24874,N_24867);
nor U25081 (N_25081,N_24903,N_24881);
xnor U25082 (N_25082,N_24951,N_24937);
xnor U25083 (N_25083,N_24922,N_24851);
xor U25084 (N_25084,N_24877,N_24837);
and U25085 (N_25085,N_24905,N_24863);
xor U25086 (N_25086,N_24974,N_24890);
nand U25087 (N_25087,N_24803,N_24912);
nand U25088 (N_25088,N_24941,N_24946);
or U25089 (N_25089,N_24835,N_24911);
nand U25090 (N_25090,N_24914,N_24962);
and U25091 (N_25091,N_24824,N_24959);
and U25092 (N_25092,N_24830,N_24807);
or U25093 (N_25093,N_24917,N_24871);
xnor U25094 (N_25094,N_24981,N_24806);
nand U25095 (N_25095,N_24953,N_24908);
and U25096 (N_25096,N_24847,N_24859);
or U25097 (N_25097,N_24899,N_24842);
xnor U25098 (N_25098,N_24860,N_24955);
nor U25099 (N_25099,N_24909,N_24854);
xor U25100 (N_25100,N_24862,N_24804);
and U25101 (N_25101,N_24801,N_24969);
xnor U25102 (N_25102,N_24810,N_24945);
nand U25103 (N_25103,N_24901,N_24979);
and U25104 (N_25104,N_24814,N_24832);
and U25105 (N_25105,N_24807,N_24826);
and U25106 (N_25106,N_24880,N_24865);
and U25107 (N_25107,N_24924,N_24871);
and U25108 (N_25108,N_24827,N_24898);
nor U25109 (N_25109,N_24949,N_24824);
nor U25110 (N_25110,N_24824,N_24804);
nand U25111 (N_25111,N_24885,N_24915);
and U25112 (N_25112,N_24993,N_24899);
or U25113 (N_25113,N_24836,N_24928);
nand U25114 (N_25114,N_24829,N_24807);
xor U25115 (N_25115,N_24978,N_24971);
xnor U25116 (N_25116,N_24808,N_24992);
nand U25117 (N_25117,N_24859,N_24901);
or U25118 (N_25118,N_24882,N_24842);
xnor U25119 (N_25119,N_24825,N_24832);
xor U25120 (N_25120,N_24816,N_24834);
nand U25121 (N_25121,N_24809,N_24808);
or U25122 (N_25122,N_24877,N_24938);
xnor U25123 (N_25123,N_24876,N_24863);
nor U25124 (N_25124,N_24852,N_24942);
nand U25125 (N_25125,N_24954,N_24812);
nand U25126 (N_25126,N_24946,N_24916);
nor U25127 (N_25127,N_24836,N_24842);
xor U25128 (N_25128,N_24828,N_24984);
xor U25129 (N_25129,N_24803,N_24800);
or U25130 (N_25130,N_24971,N_24886);
and U25131 (N_25131,N_24928,N_24975);
nor U25132 (N_25132,N_24941,N_24977);
and U25133 (N_25133,N_24871,N_24969);
nor U25134 (N_25134,N_24994,N_24935);
nor U25135 (N_25135,N_24836,N_24949);
xor U25136 (N_25136,N_24905,N_24921);
or U25137 (N_25137,N_24921,N_24867);
nand U25138 (N_25138,N_24934,N_24823);
xor U25139 (N_25139,N_24985,N_24900);
or U25140 (N_25140,N_24832,N_24975);
or U25141 (N_25141,N_24811,N_24857);
or U25142 (N_25142,N_24984,N_24972);
nand U25143 (N_25143,N_24858,N_24986);
or U25144 (N_25144,N_24914,N_24874);
nor U25145 (N_25145,N_24868,N_24873);
or U25146 (N_25146,N_24800,N_24980);
nor U25147 (N_25147,N_24967,N_24953);
and U25148 (N_25148,N_24872,N_24909);
xnor U25149 (N_25149,N_24851,N_24820);
nor U25150 (N_25150,N_24867,N_24956);
nand U25151 (N_25151,N_24878,N_24830);
or U25152 (N_25152,N_24840,N_24846);
xor U25153 (N_25153,N_24955,N_24893);
xor U25154 (N_25154,N_24838,N_24837);
or U25155 (N_25155,N_24832,N_24809);
nor U25156 (N_25156,N_24993,N_24925);
xnor U25157 (N_25157,N_24957,N_24911);
xor U25158 (N_25158,N_24874,N_24981);
xnor U25159 (N_25159,N_24808,N_24827);
xor U25160 (N_25160,N_24940,N_24920);
xor U25161 (N_25161,N_24947,N_24939);
and U25162 (N_25162,N_24827,N_24979);
nor U25163 (N_25163,N_24912,N_24956);
nand U25164 (N_25164,N_24989,N_24906);
and U25165 (N_25165,N_24825,N_24819);
xnor U25166 (N_25166,N_24967,N_24955);
or U25167 (N_25167,N_24845,N_24822);
nand U25168 (N_25168,N_24974,N_24904);
and U25169 (N_25169,N_24828,N_24962);
and U25170 (N_25170,N_24828,N_24926);
and U25171 (N_25171,N_24924,N_24808);
nand U25172 (N_25172,N_24826,N_24953);
nand U25173 (N_25173,N_24861,N_24953);
nor U25174 (N_25174,N_24809,N_24830);
nand U25175 (N_25175,N_24946,N_24896);
nor U25176 (N_25176,N_24863,N_24896);
xnor U25177 (N_25177,N_24865,N_24978);
nor U25178 (N_25178,N_24859,N_24898);
and U25179 (N_25179,N_24986,N_24992);
nor U25180 (N_25180,N_24971,N_24823);
or U25181 (N_25181,N_24988,N_24876);
xor U25182 (N_25182,N_24856,N_24866);
nor U25183 (N_25183,N_24806,N_24852);
xnor U25184 (N_25184,N_24862,N_24999);
nor U25185 (N_25185,N_24821,N_24958);
or U25186 (N_25186,N_24950,N_24926);
xor U25187 (N_25187,N_24880,N_24852);
nand U25188 (N_25188,N_24823,N_24861);
and U25189 (N_25189,N_24936,N_24846);
xnor U25190 (N_25190,N_24815,N_24824);
nor U25191 (N_25191,N_24918,N_24985);
nand U25192 (N_25192,N_24815,N_24923);
and U25193 (N_25193,N_24970,N_24997);
and U25194 (N_25194,N_24878,N_24973);
and U25195 (N_25195,N_24847,N_24863);
xnor U25196 (N_25196,N_24823,N_24856);
and U25197 (N_25197,N_24930,N_24990);
xnor U25198 (N_25198,N_24812,N_24961);
and U25199 (N_25199,N_24912,N_24909);
or U25200 (N_25200,N_25009,N_25019);
nor U25201 (N_25201,N_25060,N_25143);
nand U25202 (N_25202,N_25035,N_25124);
nor U25203 (N_25203,N_25102,N_25047);
or U25204 (N_25204,N_25054,N_25138);
nor U25205 (N_25205,N_25165,N_25137);
or U25206 (N_25206,N_25184,N_25159);
nand U25207 (N_25207,N_25155,N_25023);
nor U25208 (N_25208,N_25166,N_25075);
or U25209 (N_25209,N_25111,N_25116);
or U25210 (N_25210,N_25072,N_25170);
xor U25211 (N_25211,N_25162,N_25128);
xnor U25212 (N_25212,N_25169,N_25038);
nor U25213 (N_25213,N_25123,N_25108);
or U25214 (N_25214,N_25193,N_25092);
xor U25215 (N_25215,N_25069,N_25064);
nor U25216 (N_25216,N_25039,N_25059);
nor U25217 (N_25217,N_25010,N_25154);
xor U25218 (N_25218,N_25121,N_25145);
xnor U25219 (N_25219,N_25134,N_25070);
and U25220 (N_25220,N_25183,N_25040);
nor U25221 (N_25221,N_25104,N_25084);
nand U25222 (N_25222,N_25050,N_25174);
nand U25223 (N_25223,N_25119,N_25005);
and U25224 (N_25224,N_25034,N_25133);
nand U25225 (N_25225,N_25077,N_25164);
xnor U25226 (N_25226,N_25018,N_25061);
nand U25227 (N_25227,N_25052,N_25125);
xnor U25228 (N_25228,N_25026,N_25085);
xor U25229 (N_25229,N_25103,N_25089);
and U25230 (N_25230,N_25012,N_25041);
and U25231 (N_25231,N_25056,N_25044);
nor U25232 (N_25232,N_25100,N_25198);
xor U25233 (N_25233,N_25016,N_25036);
xor U25234 (N_25234,N_25114,N_25106);
and U25235 (N_25235,N_25113,N_25006);
or U25236 (N_25236,N_25175,N_25140);
nor U25237 (N_25237,N_25105,N_25139);
nor U25238 (N_25238,N_25015,N_25008);
or U25239 (N_25239,N_25112,N_25107);
and U25240 (N_25240,N_25147,N_25000);
or U25241 (N_25241,N_25027,N_25045);
and U25242 (N_25242,N_25029,N_25049);
and U25243 (N_25243,N_25117,N_25033);
xnor U25244 (N_25244,N_25076,N_25028);
or U25245 (N_25245,N_25109,N_25135);
or U25246 (N_25246,N_25007,N_25014);
nor U25247 (N_25247,N_25190,N_25158);
nand U25248 (N_25248,N_25189,N_25046);
and U25249 (N_25249,N_25073,N_25081);
nand U25250 (N_25250,N_25030,N_25058);
nor U25251 (N_25251,N_25129,N_25068);
nor U25252 (N_25252,N_25024,N_25067);
nor U25253 (N_25253,N_25195,N_25186);
xor U25254 (N_25254,N_25071,N_25115);
or U25255 (N_25255,N_25099,N_25087);
and U25256 (N_25256,N_25130,N_25017);
and U25257 (N_25257,N_25197,N_25181);
nor U25258 (N_25258,N_25131,N_25149);
and U25259 (N_25259,N_25142,N_25161);
or U25260 (N_25260,N_25156,N_25180);
or U25261 (N_25261,N_25022,N_25110);
and U25262 (N_25262,N_25093,N_25004);
or U25263 (N_25263,N_25003,N_25074);
nand U25264 (N_25264,N_25178,N_25013);
or U25265 (N_25265,N_25001,N_25042);
or U25266 (N_25266,N_25063,N_25098);
or U25267 (N_25267,N_25031,N_25150);
nor U25268 (N_25268,N_25120,N_25152);
xnor U25269 (N_25269,N_25171,N_25177);
or U25270 (N_25270,N_25020,N_25136);
xnor U25271 (N_25271,N_25096,N_25021);
or U25272 (N_25272,N_25043,N_25053);
xor U25273 (N_25273,N_25199,N_25182);
and U25274 (N_25274,N_25153,N_25157);
or U25275 (N_25275,N_25188,N_25179);
or U25276 (N_25276,N_25002,N_25146);
xnor U25277 (N_25277,N_25051,N_25091);
and U25278 (N_25278,N_25011,N_25194);
or U25279 (N_25279,N_25037,N_25192);
nand U25280 (N_25280,N_25168,N_25132);
nand U25281 (N_25281,N_25086,N_25097);
and U25282 (N_25282,N_25078,N_25065);
or U25283 (N_25283,N_25191,N_25080);
xor U25284 (N_25284,N_25160,N_25055);
nor U25285 (N_25285,N_25173,N_25151);
nand U25286 (N_25286,N_25163,N_25088);
or U25287 (N_25287,N_25127,N_25126);
and U25288 (N_25288,N_25025,N_25122);
nor U25289 (N_25289,N_25148,N_25176);
xnor U25290 (N_25290,N_25118,N_25083);
or U25291 (N_25291,N_25066,N_25032);
nand U25292 (N_25292,N_25196,N_25057);
nor U25293 (N_25293,N_25095,N_25090);
and U25294 (N_25294,N_25141,N_25185);
and U25295 (N_25295,N_25167,N_25101);
xnor U25296 (N_25296,N_25144,N_25048);
nand U25297 (N_25297,N_25187,N_25094);
nor U25298 (N_25298,N_25172,N_25062);
nor U25299 (N_25299,N_25079,N_25082);
nor U25300 (N_25300,N_25008,N_25070);
and U25301 (N_25301,N_25072,N_25191);
or U25302 (N_25302,N_25038,N_25027);
xnor U25303 (N_25303,N_25186,N_25084);
nor U25304 (N_25304,N_25123,N_25144);
nor U25305 (N_25305,N_25102,N_25065);
and U25306 (N_25306,N_25110,N_25187);
and U25307 (N_25307,N_25028,N_25154);
and U25308 (N_25308,N_25139,N_25028);
nand U25309 (N_25309,N_25143,N_25015);
and U25310 (N_25310,N_25013,N_25026);
and U25311 (N_25311,N_25059,N_25188);
xnor U25312 (N_25312,N_25021,N_25115);
nand U25313 (N_25313,N_25137,N_25038);
nand U25314 (N_25314,N_25098,N_25162);
nor U25315 (N_25315,N_25077,N_25175);
or U25316 (N_25316,N_25074,N_25050);
and U25317 (N_25317,N_25080,N_25027);
or U25318 (N_25318,N_25049,N_25023);
nor U25319 (N_25319,N_25189,N_25144);
nor U25320 (N_25320,N_25172,N_25196);
xor U25321 (N_25321,N_25122,N_25104);
xnor U25322 (N_25322,N_25003,N_25022);
or U25323 (N_25323,N_25056,N_25101);
nor U25324 (N_25324,N_25010,N_25016);
or U25325 (N_25325,N_25031,N_25082);
xnor U25326 (N_25326,N_25143,N_25168);
xnor U25327 (N_25327,N_25032,N_25146);
nand U25328 (N_25328,N_25149,N_25085);
nand U25329 (N_25329,N_25076,N_25150);
and U25330 (N_25330,N_25115,N_25128);
and U25331 (N_25331,N_25088,N_25118);
nor U25332 (N_25332,N_25123,N_25034);
or U25333 (N_25333,N_25191,N_25116);
xor U25334 (N_25334,N_25199,N_25187);
xor U25335 (N_25335,N_25192,N_25007);
nor U25336 (N_25336,N_25010,N_25020);
xnor U25337 (N_25337,N_25142,N_25165);
and U25338 (N_25338,N_25102,N_25160);
or U25339 (N_25339,N_25126,N_25071);
xnor U25340 (N_25340,N_25085,N_25146);
and U25341 (N_25341,N_25091,N_25068);
nand U25342 (N_25342,N_25107,N_25127);
or U25343 (N_25343,N_25125,N_25082);
nor U25344 (N_25344,N_25125,N_25083);
nor U25345 (N_25345,N_25101,N_25160);
and U25346 (N_25346,N_25066,N_25010);
xnor U25347 (N_25347,N_25023,N_25060);
xor U25348 (N_25348,N_25067,N_25036);
nor U25349 (N_25349,N_25177,N_25064);
nor U25350 (N_25350,N_25072,N_25071);
xor U25351 (N_25351,N_25096,N_25003);
or U25352 (N_25352,N_25118,N_25028);
nand U25353 (N_25353,N_25123,N_25169);
xor U25354 (N_25354,N_25172,N_25024);
and U25355 (N_25355,N_25198,N_25097);
nand U25356 (N_25356,N_25048,N_25138);
or U25357 (N_25357,N_25086,N_25131);
or U25358 (N_25358,N_25097,N_25054);
nor U25359 (N_25359,N_25198,N_25030);
and U25360 (N_25360,N_25041,N_25088);
and U25361 (N_25361,N_25113,N_25085);
nor U25362 (N_25362,N_25150,N_25170);
nor U25363 (N_25363,N_25174,N_25018);
or U25364 (N_25364,N_25119,N_25189);
xor U25365 (N_25365,N_25199,N_25004);
xnor U25366 (N_25366,N_25094,N_25029);
xnor U25367 (N_25367,N_25166,N_25040);
or U25368 (N_25368,N_25118,N_25193);
nand U25369 (N_25369,N_25090,N_25004);
nor U25370 (N_25370,N_25117,N_25063);
nor U25371 (N_25371,N_25092,N_25009);
xnor U25372 (N_25372,N_25191,N_25028);
xnor U25373 (N_25373,N_25093,N_25012);
nand U25374 (N_25374,N_25051,N_25117);
or U25375 (N_25375,N_25151,N_25106);
xnor U25376 (N_25376,N_25020,N_25104);
and U25377 (N_25377,N_25127,N_25149);
xor U25378 (N_25378,N_25156,N_25052);
xnor U25379 (N_25379,N_25060,N_25170);
nor U25380 (N_25380,N_25031,N_25024);
nor U25381 (N_25381,N_25189,N_25101);
xnor U25382 (N_25382,N_25019,N_25180);
nand U25383 (N_25383,N_25110,N_25175);
and U25384 (N_25384,N_25016,N_25130);
or U25385 (N_25385,N_25186,N_25032);
xor U25386 (N_25386,N_25064,N_25059);
nor U25387 (N_25387,N_25177,N_25092);
and U25388 (N_25388,N_25029,N_25104);
xnor U25389 (N_25389,N_25156,N_25011);
xnor U25390 (N_25390,N_25198,N_25145);
xnor U25391 (N_25391,N_25060,N_25024);
nor U25392 (N_25392,N_25186,N_25193);
or U25393 (N_25393,N_25168,N_25053);
nor U25394 (N_25394,N_25140,N_25162);
nand U25395 (N_25395,N_25065,N_25146);
nand U25396 (N_25396,N_25051,N_25045);
xnor U25397 (N_25397,N_25123,N_25018);
and U25398 (N_25398,N_25030,N_25049);
and U25399 (N_25399,N_25115,N_25164);
nor U25400 (N_25400,N_25317,N_25386);
nand U25401 (N_25401,N_25387,N_25232);
xor U25402 (N_25402,N_25261,N_25297);
nand U25403 (N_25403,N_25358,N_25349);
xnor U25404 (N_25404,N_25398,N_25208);
or U25405 (N_25405,N_25298,N_25376);
nand U25406 (N_25406,N_25211,N_25347);
nor U25407 (N_25407,N_25252,N_25291);
nand U25408 (N_25408,N_25237,N_25395);
nand U25409 (N_25409,N_25339,N_25352);
and U25410 (N_25410,N_25381,N_25219);
xor U25411 (N_25411,N_25316,N_25348);
and U25412 (N_25412,N_25325,N_25268);
xnor U25413 (N_25413,N_25356,N_25305);
and U25414 (N_25414,N_25227,N_25224);
xor U25415 (N_25415,N_25238,N_25337);
xor U25416 (N_25416,N_25295,N_25311);
nand U25417 (N_25417,N_25215,N_25258);
xor U25418 (N_25418,N_25217,N_25384);
nand U25419 (N_25419,N_25221,N_25366);
nor U25420 (N_25420,N_25353,N_25363);
xor U25421 (N_25421,N_25326,N_25245);
nand U25422 (N_25422,N_25253,N_25204);
nor U25423 (N_25423,N_25259,N_25234);
or U25424 (N_25424,N_25323,N_25236);
xor U25425 (N_25425,N_25273,N_25378);
nand U25426 (N_25426,N_25357,N_25374);
xor U25427 (N_25427,N_25292,N_25275);
xor U25428 (N_25428,N_25331,N_25389);
or U25429 (N_25429,N_25399,N_25226);
or U25430 (N_25430,N_25385,N_25248);
and U25431 (N_25431,N_25302,N_25344);
and U25432 (N_25432,N_25225,N_25355);
or U25433 (N_25433,N_25365,N_25370);
xor U25434 (N_25434,N_25321,N_25343);
nor U25435 (N_25435,N_25334,N_25255);
xor U25436 (N_25436,N_25369,N_25303);
xnor U25437 (N_25437,N_25266,N_25306);
nor U25438 (N_25438,N_25284,N_25377);
nor U25439 (N_25439,N_25318,N_25346);
or U25440 (N_25440,N_25324,N_25201);
nand U25441 (N_25441,N_25239,N_25397);
or U25442 (N_25442,N_25265,N_25379);
nand U25443 (N_25443,N_25264,N_25315);
nor U25444 (N_25444,N_25393,N_25294);
and U25445 (N_25445,N_25229,N_25241);
and U25446 (N_25446,N_25330,N_25333);
nand U25447 (N_25447,N_25279,N_25280);
and U25448 (N_25448,N_25380,N_25375);
nor U25449 (N_25449,N_25216,N_25274);
and U25450 (N_25450,N_25319,N_25367);
and U25451 (N_25451,N_25340,N_25285);
or U25452 (N_25452,N_25256,N_25212);
and U25453 (N_25453,N_25342,N_25246);
or U25454 (N_25454,N_25281,N_25220);
and U25455 (N_25455,N_25230,N_25368);
or U25456 (N_25456,N_25300,N_25202);
and U25457 (N_25457,N_25301,N_25296);
nor U25458 (N_25458,N_25350,N_25359);
or U25459 (N_25459,N_25299,N_25332);
or U25460 (N_25460,N_25341,N_25262);
nor U25461 (N_25461,N_25362,N_25200);
nand U25462 (N_25462,N_25250,N_25270);
nor U25463 (N_25463,N_25293,N_25269);
nor U25464 (N_25464,N_25313,N_25263);
xor U25465 (N_25465,N_25214,N_25307);
xor U25466 (N_25466,N_25304,N_25251);
or U25467 (N_25467,N_25257,N_25322);
or U25468 (N_25468,N_25335,N_25210);
nand U25469 (N_25469,N_25314,N_25286);
and U25470 (N_25470,N_25213,N_25203);
xnor U25471 (N_25471,N_25283,N_25254);
xnor U25472 (N_25472,N_25276,N_25364);
nor U25473 (N_25473,N_25278,N_25231);
nor U25474 (N_25474,N_25243,N_25329);
xor U25475 (N_25475,N_25338,N_25310);
or U25476 (N_25476,N_25392,N_25328);
nor U25477 (N_25477,N_25247,N_25336);
nor U25478 (N_25478,N_25351,N_25396);
or U25479 (N_25479,N_25354,N_25206);
or U25480 (N_25480,N_25242,N_25205);
and U25481 (N_25481,N_25327,N_25312);
or U25482 (N_25482,N_25394,N_25240);
or U25483 (N_25483,N_25228,N_25289);
nor U25484 (N_25484,N_25260,N_25277);
and U25485 (N_25485,N_25271,N_25209);
xor U25486 (N_25486,N_25233,N_25320);
nor U25487 (N_25487,N_25373,N_25288);
and U25488 (N_25488,N_25249,N_25207);
xor U25489 (N_25489,N_25223,N_25361);
and U25490 (N_25490,N_25287,N_25382);
and U25491 (N_25491,N_25371,N_25290);
or U25492 (N_25492,N_25372,N_25244);
or U25493 (N_25493,N_25390,N_25345);
nand U25494 (N_25494,N_25282,N_25272);
xnor U25495 (N_25495,N_25360,N_25218);
nand U25496 (N_25496,N_25383,N_25391);
or U25497 (N_25497,N_25309,N_25308);
or U25498 (N_25498,N_25235,N_25267);
and U25499 (N_25499,N_25222,N_25388);
nand U25500 (N_25500,N_25210,N_25323);
and U25501 (N_25501,N_25387,N_25226);
and U25502 (N_25502,N_25393,N_25399);
and U25503 (N_25503,N_25288,N_25318);
and U25504 (N_25504,N_25207,N_25272);
nand U25505 (N_25505,N_25285,N_25327);
or U25506 (N_25506,N_25221,N_25208);
nor U25507 (N_25507,N_25294,N_25340);
and U25508 (N_25508,N_25216,N_25281);
nand U25509 (N_25509,N_25251,N_25277);
and U25510 (N_25510,N_25252,N_25273);
and U25511 (N_25511,N_25313,N_25228);
and U25512 (N_25512,N_25215,N_25292);
xor U25513 (N_25513,N_25348,N_25386);
or U25514 (N_25514,N_25382,N_25293);
or U25515 (N_25515,N_25219,N_25330);
nand U25516 (N_25516,N_25399,N_25312);
nor U25517 (N_25517,N_25290,N_25296);
or U25518 (N_25518,N_25296,N_25246);
and U25519 (N_25519,N_25349,N_25250);
nor U25520 (N_25520,N_25280,N_25239);
xnor U25521 (N_25521,N_25202,N_25203);
or U25522 (N_25522,N_25285,N_25371);
or U25523 (N_25523,N_25230,N_25350);
nand U25524 (N_25524,N_25221,N_25361);
nor U25525 (N_25525,N_25304,N_25363);
xnor U25526 (N_25526,N_25262,N_25320);
xor U25527 (N_25527,N_25255,N_25330);
xor U25528 (N_25528,N_25266,N_25360);
or U25529 (N_25529,N_25245,N_25244);
or U25530 (N_25530,N_25350,N_25271);
or U25531 (N_25531,N_25254,N_25234);
nor U25532 (N_25532,N_25312,N_25250);
or U25533 (N_25533,N_25380,N_25324);
nor U25534 (N_25534,N_25294,N_25298);
or U25535 (N_25535,N_25225,N_25331);
or U25536 (N_25536,N_25316,N_25205);
nor U25537 (N_25537,N_25346,N_25215);
nor U25538 (N_25538,N_25227,N_25350);
nand U25539 (N_25539,N_25271,N_25290);
xnor U25540 (N_25540,N_25259,N_25268);
nor U25541 (N_25541,N_25362,N_25294);
xor U25542 (N_25542,N_25256,N_25232);
nor U25543 (N_25543,N_25292,N_25227);
nor U25544 (N_25544,N_25250,N_25356);
or U25545 (N_25545,N_25290,N_25387);
and U25546 (N_25546,N_25391,N_25269);
or U25547 (N_25547,N_25213,N_25273);
and U25548 (N_25548,N_25315,N_25271);
nand U25549 (N_25549,N_25280,N_25391);
nand U25550 (N_25550,N_25243,N_25380);
and U25551 (N_25551,N_25284,N_25279);
and U25552 (N_25552,N_25363,N_25265);
nand U25553 (N_25553,N_25221,N_25309);
or U25554 (N_25554,N_25351,N_25357);
and U25555 (N_25555,N_25299,N_25390);
or U25556 (N_25556,N_25250,N_25263);
or U25557 (N_25557,N_25344,N_25289);
nor U25558 (N_25558,N_25208,N_25356);
nor U25559 (N_25559,N_25315,N_25200);
and U25560 (N_25560,N_25373,N_25321);
nor U25561 (N_25561,N_25277,N_25296);
nor U25562 (N_25562,N_25391,N_25222);
or U25563 (N_25563,N_25224,N_25202);
and U25564 (N_25564,N_25338,N_25227);
nand U25565 (N_25565,N_25217,N_25383);
nor U25566 (N_25566,N_25310,N_25304);
and U25567 (N_25567,N_25274,N_25315);
and U25568 (N_25568,N_25230,N_25274);
nand U25569 (N_25569,N_25334,N_25309);
nor U25570 (N_25570,N_25200,N_25219);
xor U25571 (N_25571,N_25385,N_25320);
nor U25572 (N_25572,N_25262,N_25288);
nand U25573 (N_25573,N_25210,N_25339);
or U25574 (N_25574,N_25280,N_25312);
nor U25575 (N_25575,N_25299,N_25347);
nand U25576 (N_25576,N_25354,N_25334);
or U25577 (N_25577,N_25205,N_25206);
nand U25578 (N_25578,N_25338,N_25312);
and U25579 (N_25579,N_25283,N_25243);
nor U25580 (N_25580,N_25212,N_25241);
nor U25581 (N_25581,N_25253,N_25336);
and U25582 (N_25582,N_25330,N_25245);
and U25583 (N_25583,N_25322,N_25382);
or U25584 (N_25584,N_25328,N_25356);
xor U25585 (N_25585,N_25371,N_25247);
xnor U25586 (N_25586,N_25343,N_25392);
xor U25587 (N_25587,N_25377,N_25308);
nand U25588 (N_25588,N_25202,N_25251);
and U25589 (N_25589,N_25337,N_25301);
or U25590 (N_25590,N_25345,N_25218);
or U25591 (N_25591,N_25218,N_25348);
xor U25592 (N_25592,N_25267,N_25281);
or U25593 (N_25593,N_25238,N_25335);
and U25594 (N_25594,N_25295,N_25328);
or U25595 (N_25595,N_25325,N_25246);
xnor U25596 (N_25596,N_25379,N_25217);
nand U25597 (N_25597,N_25350,N_25278);
xnor U25598 (N_25598,N_25357,N_25365);
or U25599 (N_25599,N_25230,N_25280);
nand U25600 (N_25600,N_25481,N_25422);
and U25601 (N_25601,N_25480,N_25569);
nor U25602 (N_25602,N_25583,N_25501);
xor U25603 (N_25603,N_25490,N_25443);
xor U25604 (N_25604,N_25446,N_25416);
nor U25605 (N_25605,N_25522,N_25542);
xnor U25606 (N_25606,N_25467,N_25455);
or U25607 (N_25607,N_25458,N_25461);
or U25608 (N_25608,N_25534,N_25464);
and U25609 (N_25609,N_25597,N_25469);
and U25610 (N_25610,N_25548,N_25475);
and U25611 (N_25611,N_25566,N_25429);
or U25612 (N_25612,N_25592,N_25578);
nor U25613 (N_25613,N_25580,N_25436);
and U25614 (N_25614,N_25411,N_25573);
or U25615 (N_25615,N_25457,N_25451);
nand U25616 (N_25616,N_25581,N_25540);
nor U25617 (N_25617,N_25421,N_25528);
or U25618 (N_25618,N_25401,N_25599);
nor U25619 (N_25619,N_25570,N_25479);
or U25620 (N_25620,N_25444,N_25417);
nor U25621 (N_25621,N_25449,N_25439);
nand U25622 (N_25622,N_25508,N_25530);
nor U25623 (N_25623,N_25527,N_25518);
nand U25624 (N_25624,N_25477,N_25571);
xor U25625 (N_25625,N_25456,N_25520);
and U25626 (N_25626,N_25563,N_25591);
xor U25627 (N_25627,N_25561,N_25590);
and U25628 (N_25628,N_25468,N_25559);
and U25629 (N_25629,N_25400,N_25558);
xnor U25630 (N_25630,N_25478,N_25550);
xor U25631 (N_25631,N_25586,N_25503);
xnor U25632 (N_25632,N_25415,N_25406);
xnor U25633 (N_25633,N_25408,N_25463);
or U25634 (N_25634,N_25402,N_25423);
nand U25635 (N_25635,N_25459,N_25504);
nor U25636 (N_25636,N_25489,N_25433);
and U25637 (N_25637,N_25552,N_25442);
or U25638 (N_25638,N_25462,N_25512);
nand U25639 (N_25639,N_25447,N_25526);
xor U25640 (N_25640,N_25596,N_25448);
nand U25641 (N_25641,N_25574,N_25557);
nor U25642 (N_25642,N_25576,N_25587);
and U25643 (N_25643,N_25556,N_25484);
xor U25644 (N_25644,N_25440,N_25419);
or U25645 (N_25645,N_25441,N_25515);
nand U25646 (N_25646,N_25488,N_25472);
nor U25647 (N_25647,N_25428,N_25506);
nand U25648 (N_25648,N_25470,N_25567);
and U25649 (N_25649,N_25516,N_25544);
or U25650 (N_25650,N_25565,N_25553);
xor U25651 (N_25651,N_25499,N_25505);
nor U25652 (N_25652,N_25535,N_25510);
nand U25653 (N_25653,N_25498,N_25546);
xnor U25654 (N_25654,N_25476,N_25577);
or U25655 (N_25655,N_25537,N_25543);
nand U25656 (N_25656,N_25466,N_25551);
and U25657 (N_25657,N_25453,N_25555);
and U25658 (N_25658,N_25460,N_25432);
and U25659 (N_25659,N_25509,N_25431);
and U25660 (N_25660,N_25529,N_25413);
xnor U25661 (N_25661,N_25496,N_25424);
xnor U25662 (N_25662,N_25507,N_25547);
nand U25663 (N_25663,N_25405,N_25562);
xnor U25664 (N_25664,N_25579,N_25523);
nor U25665 (N_25665,N_25582,N_25427);
nor U25666 (N_25666,N_25549,N_25485);
and U25667 (N_25667,N_25502,N_25532);
and U25668 (N_25668,N_25495,N_25598);
and U25669 (N_25669,N_25575,N_25425);
nor U25670 (N_25670,N_25568,N_25545);
nand U25671 (N_25671,N_25410,N_25450);
nor U25672 (N_25672,N_25560,N_25454);
nand U25673 (N_25673,N_25538,N_25492);
nor U25674 (N_25674,N_25465,N_25403);
nand U25675 (N_25675,N_25554,N_25536);
or U25676 (N_25676,N_25412,N_25407);
and U25677 (N_25677,N_25491,N_25595);
nand U25678 (N_25678,N_25525,N_25589);
xor U25679 (N_25679,N_25519,N_25494);
xor U25680 (N_25680,N_25497,N_25430);
nand U25681 (N_25681,N_25517,N_25514);
nand U25682 (N_25682,N_25404,N_25541);
or U25683 (N_25683,N_25572,N_25409);
nand U25684 (N_25684,N_25564,N_25531);
nand U25685 (N_25685,N_25585,N_25593);
or U25686 (N_25686,N_25486,N_25438);
xnor U25687 (N_25687,N_25426,N_25420);
nand U25688 (N_25688,N_25435,N_25414);
xor U25689 (N_25689,N_25483,N_25437);
nand U25690 (N_25690,N_25482,N_25500);
nand U25691 (N_25691,N_25511,N_25434);
nor U25692 (N_25692,N_25539,N_25588);
xor U25693 (N_25693,N_25418,N_25473);
nor U25694 (N_25694,N_25524,N_25584);
and U25695 (N_25695,N_25474,N_25452);
nand U25696 (N_25696,N_25513,N_25471);
and U25697 (N_25697,N_25487,N_25533);
nand U25698 (N_25698,N_25594,N_25521);
and U25699 (N_25699,N_25445,N_25493);
or U25700 (N_25700,N_25598,N_25501);
xnor U25701 (N_25701,N_25523,N_25479);
or U25702 (N_25702,N_25539,N_25594);
xor U25703 (N_25703,N_25433,N_25598);
nor U25704 (N_25704,N_25532,N_25434);
xnor U25705 (N_25705,N_25592,N_25475);
nor U25706 (N_25706,N_25425,N_25413);
xor U25707 (N_25707,N_25447,N_25549);
nand U25708 (N_25708,N_25563,N_25480);
xnor U25709 (N_25709,N_25549,N_25585);
or U25710 (N_25710,N_25424,N_25573);
and U25711 (N_25711,N_25521,N_25575);
nand U25712 (N_25712,N_25510,N_25468);
xor U25713 (N_25713,N_25538,N_25542);
xor U25714 (N_25714,N_25515,N_25484);
nor U25715 (N_25715,N_25426,N_25498);
nand U25716 (N_25716,N_25466,N_25510);
or U25717 (N_25717,N_25484,N_25531);
nand U25718 (N_25718,N_25569,N_25590);
nor U25719 (N_25719,N_25583,N_25425);
nand U25720 (N_25720,N_25591,N_25521);
nand U25721 (N_25721,N_25401,N_25537);
nand U25722 (N_25722,N_25404,N_25555);
and U25723 (N_25723,N_25477,N_25484);
nand U25724 (N_25724,N_25543,N_25534);
or U25725 (N_25725,N_25416,N_25557);
nor U25726 (N_25726,N_25416,N_25423);
nor U25727 (N_25727,N_25410,N_25586);
or U25728 (N_25728,N_25471,N_25492);
nor U25729 (N_25729,N_25567,N_25555);
nand U25730 (N_25730,N_25592,N_25412);
nand U25731 (N_25731,N_25591,N_25577);
xor U25732 (N_25732,N_25421,N_25590);
xnor U25733 (N_25733,N_25429,N_25472);
or U25734 (N_25734,N_25446,N_25491);
or U25735 (N_25735,N_25450,N_25428);
nand U25736 (N_25736,N_25432,N_25451);
or U25737 (N_25737,N_25483,N_25585);
and U25738 (N_25738,N_25407,N_25581);
nand U25739 (N_25739,N_25521,N_25541);
xor U25740 (N_25740,N_25595,N_25596);
nor U25741 (N_25741,N_25541,N_25542);
xnor U25742 (N_25742,N_25574,N_25516);
xnor U25743 (N_25743,N_25413,N_25521);
and U25744 (N_25744,N_25513,N_25467);
and U25745 (N_25745,N_25552,N_25572);
nand U25746 (N_25746,N_25477,N_25493);
xor U25747 (N_25747,N_25410,N_25508);
nand U25748 (N_25748,N_25588,N_25436);
nor U25749 (N_25749,N_25566,N_25425);
or U25750 (N_25750,N_25558,N_25579);
nor U25751 (N_25751,N_25475,N_25433);
nand U25752 (N_25752,N_25408,N_25552);
nand U25753 (N_25753,N_25538,N_25454);
and U25754 (N_25754,N_25406,N_25537);
xor U25755 (N_25755,N_25553,N_25433);
and U25756 (N_25756,N_25553,N_25443);
and U25757 (N_25757,N_25402,N_25416);
xor U25758 (N_25758,N_25581,N_25435);
or U25759 (N_25759,N_25565,N_25554);
nand U25760 (N_25760,N_25427,N_25489);
nor U25761 (N_25761,N_25537,N_25470);
or U25762 (N_25762,N_25574,N_25590);
nand U25763 (N_25763,N_25481,N_25452);
or U25764 (N_25764,N_25461,N_25475);
nand U25765 (N_25765,N_25462,N_25567);
or U25766 (N_25766,N_25502,N_25515);
nand U25767 (N_25767,N_25552,N_25425);
nor U25768 (N_25768,N_25483,N_25559);
xor U25769 (N_25769,N_25454,N_25516);
and U25770 (N_25770,N_25572,N_25454);
nor U25771 (N_25771,N_25545,N_25570);
nand U25772 (N_25772,N_25561,N_25587);
nand U25773 (N_25773,N_25475,N_25424);
and U25774 (N_25774,N_25432,N_25505);
xor U25775 (N_25775,N_25574,N_25407);
and U25776 (N_25776,N_25494,N_25483);
nand U25777 (N_25777,N_25423,N_25530);
and U25778 (N_25778,N_25565,N_25418);
nor U25779 (N_25779,N_25484,N_25534);
nor U25780 (N_25780,N_25519,N_25527);
and U25781 (N_25781,N_25479,N_25471);
xor U25782 (N_25782,N_25475,N_25521);
nand U25783 (N_25783,N_25468,N_25401);
or U25784 (N_25784,N_25497,N_25480);
or U25785 (N_25785,N_25578,N_25576);
or U25786 (N_25786,N_25427,N_25548);
and U25787 (N_25787,N_25571,N_25441);
or U25788 (N_25788,N_25469,N_25547);
and U25789 (N_25789,N_25480,N_25527);
and U25790 (N_25790,N_25597,N_25593);
nor U25791 (N_25791,N_25405,N_25420);
xnor U25792 (N_25792,N_25420,N_25541);
or U25793 (N_25793,N_25461,N_25441);
xor U25794 (N_25794,N_25496,N_25557);
nor U25795 (N_25795,N_25523,N_25444);
nor U25796 (N_25796,N_25557,N_25583);
nor U25797 (N_25797,N_25572,N_25437);
nand U25798 (N_25798,N_25506,N_25447);
and U25799 (N_25799,N_25565,N_25519);
and U25800 (N_25800,N_25687,N_25696);
nand U25801 (N_25801,N_25742,N_25654);
nor U25802 (N_25802,N_25743,N_25795);
or U25803 (N_25803,N_25642,N_25652);
nand U25804 (N_25804,N_25622,N_25626);
or U25805 (N_25805,N_25740,N_25684);
xor U25806 (N_25806,N_25790,N_25776);
nand U25807 (N_25807,N_25739,N_25757);
and U25808 (N_25808,N_25601,N_25605);
and U25809 (N_25809,N_25699,N_25780);
nor U25810 (N_25810,N_25681,N_25784);
nand U25811 (N_25811,N_25621,N_25750);
nor U25812 (N_25812,N_25677,N_25786);
nand U25813 (N_25813,N_25744,N_25686);
and U25814 (N_25814,N_25771,N_25724);
nor U25815 (N_25815,N_25663,N_25640);
nand U25816 (N_25816,N_25615,N_25765);
or U25817 (N_25817,N_25644,N_25730);
or U25818 (N_25818,N_25702,N_25753);
or U25819 (N_25819,N_25665,N_25688);
xnor U25820 (N_25820,N_25606,N_25777);
nor U25821 (N_25821,N_25624,N_25729);
nand U25822 (N_25822,N_25643,N_25775);
and U25823 (N_25823,N_25719,N_25697);
xor U25824 (N_25824,N_25797,N_25761);
nor U25825 (N_25825,N_25655,N_25639);
and U25826 (N_25826,N_25610,N_25726);
nor U25827 (N_25827,N_25603,N_25732);
or U25828 (N_25828,N_25613,N_25628);
or U25829 (N_25829,N_25604,N_25645);
nor U25830 (N_25830,N_25612,N_25735);
xor U25831 (N_25831,N_25752,N_25781);
and U25832 (N_25832,N_25617,N_25782);
nand U25833 (N_25833,N_25635,N_25633);
or U25834 (N_25834,N_25798,N_25783);
xor U25835 (N_25835,N_25759,N_25658);
or U25836 (N_25836,N_25762,N_25703);
xnor U25837 (N_25837,N_25708,N_25768);
or U25838 (N_25838,N_25763,N_25794);
or U25839 (N_25839,N_25716,N_25737);
or U25840 (N_25840,N_25600,N_25650);
nor U25841 (N_25841,N_25689,N_25659);
nor U25842 (N_25842,N_25733,N_25669);
nor U25843 (N_25843,N_25602,N_25675);
nand U25844 (N_25844,N_25670,N_25676);
nor U25845 (N_25845,N_25636,N_25792);
and U25846 (N_25846,N_25711,N_25754);
and U25847 (N_25847,N_25700,N_25788);
xnor U25848 (N_25848,N_25727,N_25690);
xnor U25849 (N_25849,N_25647,N_25799);
nor U25850 (N_25850,N_25680,N_25692);
nor U25851 (N_25851,N_25651,N_25661);
nor U25852 (N_25852,N_25738,N_25704);
xnor U25853 (N_25853,N_25764,N_25769);
nor U25854 (N_25854,N_25674,N_25629);
nand U25855 (N_25855,N_25660,N_25685);
nor U25856 (N_25856,N_25646,N_25721);
xor U25857 (N_25857,N_25707,N_25749);
and U25858 (N_25858,N_25714,N_25793);
and U25859 (N_25859,N_25722,N_25666);
nor U25860 (N_25860,N_25789,N_25710);
nor U25861 (N_25861,N_25767,N_25634);
nor U25862 (N_25862,N_25630,N_25648);
and U25863 (N_25863,N_25760,N_25667);
and U25864 (N_25864,N_25785,N_25607);
nor U25865 (N_25865,N_25734,N_25672);
nor U25866 (N_25866,N_25627,N_25693);
nor U25867 (N_25867,N_25796,N_25747);
nand U25868 (N_25868,N_25691,N_25608);
xor U25869 (N_25869,N_25706,N_25656);
xor U25870 (N_25870,N_25683,N_25637);
xnor U25871 (N_25871,N_25791,N_25662);
nand U25872 (N_25872,N_25713,N_25701);
or U25873 (N_25873,N_25773,N_25787);
xnor U25874 (N_25874,N_25625,N_25649);
nand U25875 (N_25875,N_25657,N_25720);
and U25876 (N_25876,N_25609,N_25728);
xnor U25877 (N_25877,N_25736,N_25705);
nor U25878 (N_25878,N_25653,N_25694);
nand U25879 (N_25879,N_25755,N_25638);
xor U25880 (N_25880,N_25631,N_25751);
and U25881 (N_25881,N_25731,N_25758);
and U25882 (N_25882,N_25723,N_25671);
xnor U25883 (N_25883,N_25770,N_25682);
nand U25884 (N_25884,N_25679,N_25741);
nor U25885 (N_25885,N_25620,N_25632);
nor U25886 (N_25886,N_25756,N_25712);
nor U25887 (N_25887,N_25748,N_25766);
and U25888 (N_25888,N_25778,N_25614);
nor U25889 (N_25889,N_25664,N_25745);
nor U25890 (N_25890,N_25717,N_25709);
nor U25891 (N_25891,N_25725,N_25698);
nand U25892 (N_25892,N_25619,N_25772);
or U25893 (N_25893,N_25746,N_25774);
or U25894 (N_25894,N_25616,N_25715);
nor U25895 (N_25895,N_25678,N_25668);
nand U25896 (N_25896,N_25695,N_25718);
nand U25897 (N_25897,N_25779,N_25623);
nor U25898 (N_25898,N_25641,N_25618);
and U25899 (N_25899,N_25673,N_25611);
and U25900 (N_25900,N_25733,N_25687);
or U25901 (N_25901,N_25693,N_25648);
xnor U25902 (N_25902,N_25672,N_25663);
or U25903 (N_25903,N_25685,N_25611);
and U25904 (N_25904,N_25657,N_25711);
nor U25905 (N_25905,N_25729,N_25660);
and U25906 (N_25906,N_25769,N_25624);
and U25907 (N_25907,N_25618,N_25721);
nor U25908 (N_25908,N_25648,N_25623);
or U25909 (N_25909,N_25664,N_25704);
or U25910 (N_25910,N_25617,N_25710);
nor U25911 (N_25911,N_25703,N_25685);
xor U25912 (N_25912,N_25706,N_25714);
or U25913 (N_25913,N_25794,N_25635);
and U25914 (N_25914,N_25773,N_25683);
nor U25915 (N_25915,N_25604,N_25777);
and U25916 (N_25916,N_25641,N_25627);
nand U25917 (N_25917,N_25619,N_25642);
nand U25918 (N_25918,N_25676,N_25791);
and U25919 (N_25919,N_25650,N_25671);
nor U25920 (N_25920,N_25666,N_25714);
xor U25921 (N_25921,N_25726,N_25646);
xor U25922 (N_25922,N_25799,N_25631);
nand U25923 (N_25923,N_25607,N_25675);
and U25924 (N_25924,N_25621,N_25777);
nor U25925 (N_25925,N_25716,N_25711);
nor U25926 (N_25926,N_25698,N_25701);
or U25927 (N_25927,N_25662,N_25633);
nor U25928 (N_25928,N_25673,N_25772);
or U25929 (N_25929,N_25772,N_25786);
or U25930 (N_25930,N_25614,N_25728);
xnor U25931 (N_25931,N_25699,N_25797);
nor U25932 (N_25932,N_25744,N_25637);
nand U25933 (N_25933,N_25689,N_25755);
and U25934 (N_25934,N_25701,N_25664);
nor U25935 (N_25935,N_25691,N_25763);
xor U25936 (N_25936,N_25714,N_25687);
nor U25937 (N_25937,N_25625,N_25767);
nand U25938 (N_25938,N_25698,N_25659);
xor U25939 (N_25939,N_25612,N_25752);
nor U25940 (N_25940,N_25670,N_25741);
nor U25941 (N_25941,N_25715,N_25771);
and U25942 (N_25942,N_25650,N_25775);
nand U25943 (N_25943,N_25655,N_25742);
nand U25944 (N_25944,N_25616,N_25792);
and U25945 (N_25945,N_25694,N_25799);
nor U25946 (N_25946,N_25729,N_25701);
and U25947 (N_25947,N_25622,N_25650);
nand U25948 (N_25948,N_25603,N_25601);
or U25949 (N_25949,N_25707,N_25739);
nor U25950 (N_25950,N_25720,N_25683);
nand U25951 (N_25951,N_25693,N_25777);
or U25952 (N_25952,N_25721,N_25776);
or U25953 (N_25953,N_25726,N_25761);
or U25954 (N_25954,N_25626,N_25717);
nor U25955 (N_25955,N_25742,N_25630);
and U25956 (N_25956,N_25635,N_25697);
nand U25957 (N_25957,N_25718,N_25712);
xor U25958 (N_25958,N_25616,N_25671);
xor U25959 (N_25959,N_25705,N_25757);
and U25960 (N_25960,N_25740,N_25766);
xor U25961 (N_25961,N_25644,N_25745);
xor U25962 (N_25962,N_25679,N_25662);
nand U25963 (N_25963,N_25759,N_25679);
or U25964 (N_25964,N_25670,N_25730);
xor U25965 (N_25965,N_25768,N_25676);
xor U25966 (N_25966,N_25675,N_25719);
nor U25967 (N_25967,N_25705,N_25629);
xnor U25968 (N_25968,N_25717,N_25750);
or U25969 (N_25969,N_25744,N_25622);
nor U25970 (N_25970,N_25643,N_25716);
nor U25971 (N_25971,N_25670,N_25614);
or U25972 (N_25972,N_25736,N_25799);
xor U25973 (N_25973,N_25676,N_25654);
or U25974 (N_25974,N_25662,N_25600);
or U25975 (N_25975,N_25614,N_25790);
nor U25976 (N_25976,N_25760,N_25709);
and U25977 (N_25977,N_25660,N_25633);
and U25978 (N_25978,N_25640,N_25766);
xor U25979 (N_25979,N_25738,N_25640);
or U25980 (N_25980,N_25728,N_25791);
nand U25981 (N_25981,N_25608,N_25674);
nor U25982 (N_25982,N_25631,N_25613);
nor U25983 (N_25983,N_25781,N_25769);
and U25984 (N_25984,N_25614,N_25698);
and U25985 (N_25985,N_25708,N_25764);
or U25986 (N_25986,N_25697,N_25729);
nand U25987 (N_25987,N_25790,N_25671);
and U25988 (N_25988,N_25780,N_25746);
xnor U25989 (N_25989,N_25608,N_25737);
and U25990 (N_25990,N_25725,N_25736);
nand U25991 (N_25991,N_25793,N_25740);
and U25992 (N_25992,N_25690,N_25619);
and U25993 (N_25993,N_25654,N_25634);
nand U25994 (N_25994,N_25628,N_25641);
and U25995 (N_25995,N_25727,N_25781);
nor U25996 (N_25996,N_25605,N_25619);
or U25997 (N_25997,N_25719,N_25715);
and U25998 (N_25998,N_25692,N_25722);
xor U25999 (N_25999,N_25702,N_25783);
or U26000 (N_26000,N_25951,N_25974);
and U26001 (N_26001,N_25900,N_25965);
and U26002 (N_26002,N_25937,N_25925);
or U26003 (N_26003,N_25857,N_25835);
or U26004 (N_26004,N_25856,N_25822);
nand U26005 (N_26005,N_25927,N_25874);
and U26006 (N_26006,N_25980,N_25899);
nor U26007 (N_26007,N_25804,N_25904);
or U26008 (N_26008,N_25842,N_25948);
xnor U26009 (N_26009,N_25845,N_25991);
and U26010 (N_26010,N_25905,N_25946);
and U26011 (N_26011,N_25979,N_25893);
nor U26012 (N_26012,N_25993,N_25975);
or U26013 (N_26013,N_25877,N_25981);
xor U26014 (N_26014,N_25994,N_25918);
or U26015 (N_26015,N_25885,N_25929);
nand U26016 (N_26016,N_25935,N_25864);
or U26017 (N_26017,N_25992,N_25800);
nand U26018 (N_26018,N_25967,N_25880);
or U26019 (N_26019,N_25956,N_25851);
nand U26020 (N_26020,N_25843,N_25895);
or U26021 (N_26021,N_25821,N_25852);
nand U26022 (N_26022,N_25823,N_25999);
or U26023 (N_26023,N_25997,N_25969);
and U26024 (N_26024,N_25995,N_25832);
xnor U26025 (N_26025,N_25908,N_25962);
or U26026 (N_26026,N_25887,N_25973);
or U26027 (N_26027,N_25984,N_25878);
nand U26028 (N_26028,N_25959,N_25976);
xnor U26029 (N_26029,N_25872,N_25819);
and U26030 (N_26030,N_25901,N_25868);
nand U26031 (N_26031,N_25978,N_25849);
or U26032 (N_26032,N_25869,N_25854);
nor U26033 (N_26033,N_25910,N_25917);
or U26034 (N_26034,N_25846,N_25886);
nand U26035 (N_26035,N_25820,N_25943);
or U26036 (N_26036,N_25963,N_25862);
and U26037 (N_26037,N_25987,N_25894);
or U26038 (N_26038,N_25928,N_25989);
or U26039 (N_26039,N_25806,N_25924);
xor U26040 (N_26040,N_25824,N_25986);
nand U26041 (N_26041,N_25813,N_25801);
and U26042 (N_26042,N_25817,N_25947);
xor U26043 (N_26043,N_25884,N_25830);
and U26044 (N_26044,N_25903,N_25939);
nor U26045 (N_26045,N_25890,N_25985);
or U26046 (N_26046,N_25815,N_25998);
nand U26047 (N_26047,N_25811,N_25936);
or U26048 (N_26048,N_25915,N_25896);
nor U26049 (N_26049,N_25941,N_25838);
nand U26050 (N_26050,N_25945,N_25906);
xnor U26051 (N_26051,N_25810,N_25831);
nor U26052 (N_26052,N_25971,N_25911);
xor U26053 (N_26053,N_25802,N_25982);
xnor U26054 (N_26054,N_25960,N_25883);
nor U26055 (N_26055,N_25879,N_25934);
and U26056 (N_26056,N_25855,N_25818);
and U26057 (N_26057,N_25950,N_25921);
nand U26058 (N_26058,N_25949,N_25827);
nand U26059 (N_26059,N_25958,N_25844);
and U26060 (N_26060,N_25870,N_25876);
nor U26061 (N_26061,N_25840,N_25961);
and U26062 (N_26062,N_25940,N_25847);
xor U26063 (N_26063,N_25858,N_25836);
nor U26064 (N_26064,N_25996,N_25957);
xnor U26065 (N_26065,N_25865,N_25860);
and U26066 (N_26066,N_25912,N_25850);
nand U26067 (N_26067,N_25972,N_25988);
nand U26068 (N_26068,N_25873,N_25863);
nand U26069 (N_26069,N_25913,N_25931);
nor U26070 (N_26070,N_25933,N_25897);
and U26071 (N_26071,N_25861,N_25839);
xnor U26072 (N_26072,N_25859,N_25816);
or U26073 (N_26073,N_25983,N_25805);
nand U26074 (N_26074,N_25907,N_25825);
nand U26075 (N_26075,N_25814,N_25848);
xnor U26076 (N_26076,N_25942,N_25875);
and U26077 (N_26077,N_25966,N_25955);
xnor U26078 (N_26078,N_25834,N_25968);
or U26079 (N_26079,N_25871,N_25833);
nand U26080 (N_26080,N_25952,N_25954);
nor U26081 (N_26081,N_25889,N_25829);
and U26082 (N_26082,N_25809,N_25881);
xor U26083 (N_26083,N_25938,N_25828);
nor U26084 (N_26084,N_25867,N_25932);
or U26085 (N_26085,N_25898,N_25807);
or U26086 (N_26086,N_25826,N_25919);
nand U26087 (N_26087,N_25922,N_25953);
xor U26088 (N_26088,N_25892,N_25909);
or U26089 (N_26089,N_25970,N_25916);
and U26090 (N_26090,N_25977,N_25902);
and U26091 (N_26091,N_25891,N_25808);
nor U26092 (N_26092,N_25882,N_25837);
nand U26093 (N_26093,N_25866,N_25812);
xor U26094 (N_26094,N_25990,N_25841);
or U26095 (N_26095,N_25853,N_25930);
nor U26096 (N_26096,N_25914,N_25888);
xor U26097 (N_26097,N_25964,N_25923);
nor U26098 (N_26098,N_25920,N_25926);
or U26099 (N_26099,N_25944,N_25803);
or U26100 (N_26100,N_25809,N_25935);
or U26101 (N_26101,N_25805,N_25890);
and U26102 (N_26102,N_25959,N_25888);
or U26103 (N_26103,N_25877,N_25918);
nor U26104 (N_26104,N_25979,N_25884);
nor U26105 (N_26105,N_25812,N_25915);
xnor U26106 (N_26106,N_25985,N_25828);
nor U26107 (N_26107,N_25811,N_25902);
xnor U26108 (N_26108,N_25859,N_25911);
and U26109 (N_26109,N_25810,N_25996);
xor U26110 (N_26110,N_25984,N_25845);
or U26111 (N_26111,N_25953,N_25891);
and U26112 (N_26112,N_25915,N_25961);
nor U26113 (N_26113,N_25984,N_25930);
and U26114 (N_26114,N_25869,N_25945);
nor U26115 (N_26115,N_25898,N_25809);
nand U26116 (N_26116,N_25827,N_25823);
xnor U26117 (N_26117,N_25983,N_25936);
nand U26118 (N_26118,N_25959,N_25981);
nand U26119 (N_26119,N_25827,N_25845);
nand U26120 (N_26120,N_25894,N_25836);
or U26121 (N_26121,N_25982,N_25961);
or U26122 (N_26122,N_25890,N_25879);
or U26123 (N_26123,N_25877,N_25934);
nor U26124 (N_26124,N_25927,N_25899);
nand U26125 (N_26125,N_25873,N_25866);
or U26126 (N_26126,N_25941,N_25942);
nor U26127 (N_26127,N_25883,N_25909);
nor U26128 (N_26128,N_25877,N_25921);
nand U26129 (N_26129,N_25996,N_25815);
and U26130 (N_26130,N_25865,N_25924);
or U26131 (N_26131,N_25839,N_25924);
and U26132 (N_26132,N_25907,N_25977);
nor U26133 (N_26133,N_25964,N_25912);
nor U26134 (N_26134,N_25807,N_25980);
nand U26135 (N_26135,N_25823,N_25899);
nor U26136 (N_26136,N_25924,N_25802);
xor U26137 (N_26137,N_25891,N_25906);
or U26138 (N_26138,N_25914,N_25805);
or U26139 (N_26139,N_25829,N_25882);
nand U26140 (N_26140,N_25979,N_25803);
and U26141 (N_26141,N_25816,N_25911);
nand U26142 (N_26142,N_25817,N_25995);
nand U26143 (N_26143,N_25954,N_25901);
nand U26144 (N_26144,N_25969,N_25845);
or U26145 (N_26145,N_25841,N_25842);
and U26146 (N_26146,N_25956,N_25883);
xnor U26147 (N_26147,N_25947,N_25983);
and U26148 (N_26148,N_25891,N_25949);
or U26149 (N_26149,N_25984,N_25909);
or U26150 (N_26150,N_25886,N_25817);
nor U26151 (N_26151,N_25958,N_25852);
xor U26152 (N_26152,N_25966,N_25801);
nor U26153 (N_26153,N_25801,N_25834);
nor U26154 (N_26154,N_25959,N_25885);
or U26155 (N_26155,N_25985,N_25858);
nand U26156 (N_26156,N_25888,N_25942);
nand U26157 (N_26157,N_25896,N_25854);
nor U26158 (N_26158,N_25894,N_25964);
nor U26159 (N_26159,N_25879,N_25995);
or U26160 (N_26160,N_25852,N_25936);
xor U26161 (N_26161,N_25971,N_25846);
nand U26162 (N_26162,N_25853,N_25929);
or U26163 (N_26163,N_25906,N_25837);
nor U26164 (N_26164,N_25831,N_25847);
or U26165 (N_26165,N_25851,N_25818);
xor U26166 (N_26166,N_25996,N_25904);
or U26167 (N_26167,N_25812,N_25962);
nor U26168 (N_26168,N_25982,N_25914);
or U26169 (N_26169,N_25804,N_25921);
or U26170 (N_26170,N_25892,N_25805);
and U26171 (N_26171,N_25851,N_25945);
nand U26172 (N_26172,N_25958,N_25890);
nand U26173 (N_26173,N_25825,N_25966);
nand U26174 (N_26174,N_25911,N_25824);
nor U26175 (N_26175,N_25952,N_25820);
or U26176 (N_26176,N_25826,N_25872);
nor U26177 (N_26177,N_25823,N_25998);
nor U26178 (N_26178,N_25965,N_25902);
nand U26179 (N_26179,N_25871,N_25844);
nor U26180 (N_26180,N_25912,N_25833);
nor U26181 (N_26181,N_25874,N_25883);
or U26182 (N_26182,N_25961,N_25929);
nor U26183 (N_26183,N_25911,N_25960);
xor U26184 (N_26184,N_25974,N_25811);
nor U26185 (N_26185,N_25810,N_25867);
nand U26186 (N_26186,N_25817,N_25866);
or U26187 (N_26187,N_25975,N_25843);
nand U26188 (N_26188,N_25808,N_25820);
nand U26189 (N_26189,N_25957,N_25850);
nor U26190 (N_26190,N_25816,N_25836);
xnor U26191 (N_26191,N_25963,N_25900);
nand U26192 (N_26192,N_25841,N_25937);
and U26193 (N_26193,N_25985,N_25824);
xor U26194 (N_26194,N_25868,N_25823);
and U26195 (N_26195,N_25951,N_25988);
nor U26196 (N_26196,N_25932,N_25826);
xor U26197 (N_26197,N_25910,N_25923);
xnor U26198 (N_26198,N_25910,N_25993);
and U26199 (N_26199,N_25908,N_25905);
and U26200 (N_26200,N_26137,N_26193);
nor U26201 (N_26201,N_26073,N_26050);
nand U26202 (N_26202,N_26109,N_26185);
or U26203 (N_26203,N_26104,N_26140);
or U26204 (N_26204,N_26111,N_26002);
xnor U26205 (N_26205,N_26108,N_26102);
or U26206 (N_26206,N_26083,N_26196);
or U26207 (N_26207,N_26064,N_26165);
and U26208 (N_26208,N_26060,N_26003);
nand U26209 (N_26209,N_26084,N_26095);
xor U26210 (N_26210,N_26094,N_26045);
and U26211 (N_26211,N_26175,N_26163);
nor U26212 (N_26212,N_26098,N_26038);
and U26213 (N_26213,N_26047,N_26116);
xnor U26214 (N_26214,N_26029,N_26026);
nand U26215 (N_26215,N_26115,N_26033);
or U26216 (N_26216,N_26187,N_26182);
nand U26217 (N_26217,N_26001,N_26015);
xor U26218 (N_26218,N_26117,N_26171);
and U26219 (N_26219,N_26142,N_26020);
and U26220 (N_26220,N_26017,N_26123);
nor U26221 (N_26221,N_26048,N_26191);
or U26222 (N_26222,N_26063,N_26053);
and U26223 (N_26223,N_26099,N_26160);
xnor U26224 (N_26224,N_26180,N_26167);
xnor U26225 (N_26225,N_26061,N_26164);
or U26226 (N_26226,N_26176,N_26016);
xor U26227 (N_26227,N_26034,N_26028);
nor U26228 (N_26228,N_26105,N_26145);
nor U26229 (N_26229,N_26152,N_26172);
nand U26230 (N_26230,N_26122,N_26159);
nor U26231 (N_26231,N_26051,N_26067);
xor U26232 (N_26232,N_26069,N_26097);
or U26233 (N_26233,N_26025,N_26043);
and U26234 (N_26234,N_26155,N_26021);
or U26235 (N_26235,N_26081,N_26149);
nand U26236 (N_26236,N_26091,N_26089);
nor U26237 (N_26237,N_26046,N_26166);
nor U26238 (N_26238,N_26085,N_26019);
nand U26239 (N_26239,N_26106,N_26018);
nand U26240 (N_26240,N_26154,N_26134);
xnor U26241 (N_26241,N_26042,N_26030);
and U26242 (N_26242,N_26041,N_26143);
and U26243 (N_26243,N_26023,N_26103);
nand U26244 (N_26244,N_26027,N_26198);
xnor U26245 (N_26245,N_26192,N_26024);
and U26246 (N_26246,N_26054,N_26070);
xnor U26247 (N_26247,N_26161,N_26074);
nor U26248 (N_26248,N_26110,N_26199);
nand U26249 (N_26249,N_26181,N_26009);
nand U26250 (N_26250,N_26101,N_26133);
and U26251 (N_26251,N_26141,N_26135);
nor U26252 (N_26252,N_26014,N_26078);
xnor U26253 (N_26253,N_26113,N_26178);
nand U26254 (N_26254,N_26128,N_26184);
nor U26255 (N_26255,N_26077,N_26032);
nor U26256 (N_26256,N_26072,N_26000);
nor U26257 (N_26257,N_26082,N_26126);
nand U26258 (N_26258,N_26120,N_26153);
and U26259 (N_26259,N_26056,N_26156);
xor U26260 (N_26260,N_26066,N_26130);
xnor U26261 (N_26261,N_26146,N_26188);
nand U26262 (N_26262,N_26059,N_26186);
xnor U26263 (N_26263,N_26065,N_26151);
nand U26264 (N_26264,N_26131,N_26088);
nand U26265 (N_26265,N_26055,N_26007);
nand U26266 (N_26266,N_26010,N_26136);
nor U26267 (N_26267,N_26138,N_26093);
and U26268 (N_26268,N_26075,N_26006);
nand U26269 (N_26269,N_26079,N_26087);
or U26270 (N_26270,N_26036,N_26158);
nor U26271 (N_26271,N_26121,N_26129);
or U26272 (N_26272,N_26005,N_26035);
xnor U26273 (N_26273,N_26068,N_26144);
xor U26274 (N_26274,N_26058,N_26086);
xnor U26275 (N_26275,N_26183,N_26022);
or U26276 (N_26276,N_26076,N_26139);
nand U26277 (N_26277,N_26124,N_26011);
nor U26278 (N_26278,N_26062,N_26119);
and U26279 (N_26279,N_26150,N_26031);
and U26280 (N_26280,N_26148,N_26044);
nand U26281 (N_26281,N_26162,N_26013);
and U26282 (N_26282,N_26174,N_26157);
nor U26283 (N_26283,N_26039,N_26012);
nand U26284 (N_26284,N_26168,N_26173);
or U26285 (N_26285,N_26008,N_26037);
xnor U26286 (N_26286,N_26049,N_26052);
nand U26287 (N_26287,N_26177,N_26179);
or U26288 (N_26288,N_26090,N_26096);
xnor U26289 (N_26289,N_26169,N_26114);
nand U26290 (N_26290,N_26194,N_26092);
nand U26291 (N_26291,N_26118,N_26057);
nand U26292 (N_26292,N_26080,N_26197);
or U26293 (N_26293,N_26190,N_26147);
and U26294 (N_26294,N_26170,N_26195);
xnor U26295 (N_26295,N_26040,N_26112);
nand U26296 (N_26296,N_26125,N_26004);
xor U26297 (N_26297,N_26071,N_26132);
and U26298 (N_26298,N_26127,N_26189);
xor U26299 (N_26299,N_26107,N_26100);
and U26300 (N_26300,N_26061,N_26186);
nand U26301 (N_26301,N_26058,N_26015);
xnor U26302 (N_26302,N_26016,N_26096);
nand U26303 (N_26303,N_26070,N_26185);
nor U26304 (N_26304,N_26006,N_26012);
or U26305 (N_26305,N_26170,N_26151);
nor U26306 (N_26306,N_26054,N_26166);
xor U26307 (N_26307,N_26015,N_26074);
nor U26308 (N_26308,N_26029,N_26060);
xnor U26309 (N_26309,N_26009,N_26046);
xnor U26310 (N_26310,N_26029,N_26062);
nand U26311 (N_26311,N_26004,N_26010);
nor U26312 (N_26312,N_26044,N_26198);
or U26313 (N_26313,N_26028,N_26136);
nand U26314 (N_26314,N_26043,N_26181);
and U26315 (N_26315,N_26091,N_26037);
nor U26316 (N_26316,N_26194,N_26101);
or U26317 (N_26317,N_26079,N_26111);
nor U26318 (N_26318,N_26084,N_26149);
nand U26319 (N_26319,N_26043,N_26049);
xor U26320 (N_26320,N_26099,N_26101);
nand U26321 (N_26321,N_26073,N_26063);
and U26322 (N_26322,N_26044,N_26030);
nand U26323 (N_26323,N_26093,N_26032);
xor U26324 (N_26324,N_26128,N_26060);
or U26325 (N_26325,N_26170,N_26156);
or U26326 (N_26326,N_26025,N_26101);
nand U26327 (N_26327,N_26064,N_26185);
nand U26328 (N_26328,N_26035,N_26198);
nand U26329 (N_26329,N_26001,N_26183);
nor U26330 (N_26330,N_26080,N_26051);
nor U26331 (N_26331,N_26163,N_26145);
xor U26332 (N_26332,N_26177,N_26074);
nand U26333 (N_26333,N_26169,N_26112);
or U26334 (N_26334,N_26040,N_26144);
or U26335 (N_26335,N_26070,N_26179);
xor U26336 (N_26336,N_26158,N_26155);
or U26337 (N_26337,N_26071,N_26138);
xnor U26338 (N_26338,N_26175,N_26186);
and U26339 (N_26339,N_26085,N_26077);
and U26340 (N_26340,N_26077,N_26068);
xor U26341 (N_26341,N_26060,N_26082);
nand U26342 (N_26342,N_26107,N_26113);
or U26343 (N_26343,N_26051,N_26010);
nor U26344 (N_26344,N_26106,N_26048);
nand U26345 (N_26345,N_26112,N_26038);
xnor U26346 (N_26346,N_26073,N_26107);
or U26347 (N_26347,N_26034,N_26049);
or U26348 (N_26348,N_26175,N_26103);
or U26349 (N_26349,N_26196,N_26140);
xor U26350 (N_26350,N_26017,N_26109);
and U26351 (N_26351,N_26076,N_26131);
xor U26352 (N_26352,N_26171,N_26173);
nor U26353 (N_26353,N_26040,N_26077);
and U26354 (N_26354,N_26025,N_26012);
and U26355 (N_26355,N_26063,N_26182);
nand U26356 (N_26356,N_26035,N_26025);
and U26357 (N_26357,N_26094,N_26081);
nand U26358 (N_26358,N_26007,N_26121);
xor U26359 (N_26359,N_26186,N_26096);
nand U26360 (N_26360,N_26141,N_26142);
and U26361 (N_26361,N_26000,N_26004);
nand U26362 (N_26362,N_26094,N_26127);
nand U26363 (N_26363,N_26168,N_26190);
xnor U26364 (N_26364,N_26093,N_26021);
or U26365 (N_26365,N_26056,N_26069);
and U26366 (N_26366,N_26060,N_26057);
and U26367 (N_26367,N_26030,N_26008);
and U26368 (N_26368,N_26012,N_26076);
nand U26369 (N_26369,N_26095,N_26052);
or U26370 (N_26370,N_26082,N_26015);
or U26371 (N_26371,N_26195,N_26024);
or U26372 (N_26372,N_26039,N_26003);
nor U26373 (N_26373,N_26007,N_26069);
nand U26374 (N_26374,N_26131,N_26093);
nand U26375 (N_26375,N_26182,N_26163);
nor U26376 (N_26376,N_26076,N_26097);
nand U26377 (N_26377,N_26035,N_26027);
nand U26378 (N_26378,N_26144,N_26175);
xnor U26379 (N_26379,N_26144,N_26142);
xnor U26380 (N_26380,N_26015,N_26198);
or U26381 (N_26381,N_26192,N_26194);
and U26382 (N_26382,N_26009,N_26069);
xnor U26383 (N_26383,N_26124,N_26073);
and U26384 (N_26384,N_26034,N_26123);
and U26385 (N_26385,N_26012,N_26034);
nand U26386 (N_26386,N_26172,N_26162);
xnor U26387 (N_26387,N_26025,N_26019);
or U26388 (N_26388,N_26043,N_26169);
nor U26389 (N_26389,N_26006,N_26083);
nor U26390 (N_26390,N_26118,N_26058);
nor U26391 (N_26391,N_26043,N_26116);
xnor U26392 (N_26392,N_26185,N_26086);
or U26393 (N_26393,N_26160,N_26061);
nor U26394 (N_26394,N_26155,N_26144);
or U26395 (N_26395,N_26184,N_26180);
or U26396 (N_26396,N_26054,N_26090);
or U26397 (N_26397,N_26089,N_26186);
nor U26398 (N_26398,N_26104,N_26026);
and U26399 (N_26399,N_26155,N_26185);
xnor U26400 (N_26400,N_26313,N_26311);
xnor U26401 (N_26401,N_26260,N_26340);
xor U26402 (N_26402,N_26223,N_26300);
nand U26403 (N_26403,N_26322,N_26296);
or U26404 (N_26404,N_26297,N_26278);
xnor U26405 (N_26405,N_26203,N_26209);
and U26406 (N_26406,N_26335,N_26309);
and U26407 (N_26407,N_26253,N_26266);
and U26408 (N_26408,N_26380,N_26204);
nand U26409 (N_26409,N_26282,N_26274);
or U26410 (N_26410,N_26306,N_26333);
nand U26411 (N_26411,N_26331,N_26247);
or U26412 (N_26412,N_26254,N_26328);
and U26413 (N_26413,N_26276,N_26391);
nor U26414 (N_26414,N_26358,N_26373);
nor U26415 (N_26415,N_26366,N_26367);
or U26416 (N_26416,N_26320,N_26308);
or U26417 (N_26417,N_26210,N_26268);
or U26418 (N_26418,N_26377,N_26289);
and U26419 (N_26419,N_26299,N_26200);
nand U26420 (N_26420,N_26215,N_26239);
and U26421 (N_26421,N_26364,N_26399);
xor U26422 (N_26422,N_26393,N_26218);
or U26423 (N_26423,N_26387,N_26201);
and U26424 (N_26424,N_26235,N_26369);
xnor U26425 (N_26425,N_26326,N_26284);
or U26426 (N_26426,N_26305,N_26269);
nor U26427 (N_26427,N_26245,N_26376);
xnor U26428 (N_26428,N_26291,N_26265);
nor U26429 (N_26429,N_26233,N_26352);
nor U26430 (N_26430,N_26222,N_26270);
and U26431 (N_26431,N_26341,N_26386);
nor U26432 (N_26432,N_26287,N_26259);
nor U26433 (N_26433,N_26251,N_26250);
and U26434 (N_26434,N_26382,N_26318);
nand U26435 (N_26435,N_26319,N_26385);
nand U26436 (N_26436,N_26219,N_26396);
or U26437 (N_26437,N_26221,N_26310);
or U26438 (N_26438,N_26324,N_26304);
xnor U26439 (N_26439,N_26342,N_26224);
or U26440 (N_26440,N_26359,N_26280);
nor U26441 (N_26441,N_26336,N_26256);
xnor U26442 (N_26442,N_26220,N_26263);
or U26443 (N_26443,N_26240,N_26361);
and U26444 (N_26444,N_26234,N_26343);
xor U26445 (N_26445,N_26357,N_26321);
xor U26446 (N_26446,N_26271,N_26395);
nand U26447 (N_26447,N_26258,N_26248);
nand U26448 (N_26448,N_26273,N_26283);
nand U26449 (N_26449,N_26206,N_26261);
xor U26450 (N_26450,N_26211,N_26372);
and U26451 (N_26451,N_26232,N_26236);
or U26452 (N_26452,N_26327,N_26344);
and U26453 (N_26453,N_26348,N_26243);
and U26454 (N_26454,N_26293,N_26267);
and U26455 (N_26455,N_26317,N_26371);
nand U26456 (N_26456,N_26370,N_26337);
and U26457 (N_26457,N_26207,N_26355);
xor U26458 (N_26458,N_26356,N_26384);
and U26459 (N_26459,N_26338,N_26397);
nor U26460 (N_26460,N_26281,N_26398);
nor U26461 (N_26461,N_26330,N_26301);
nand U26462 (N_26462,N_26237,N_26388);
xor U26463 (N_26463,N_26242,N_26349);
nor U26464 (N_26464,N_26392,N_26363);
nor U26465 (N_26465,N_26362,N_26257);
xnor U26466 (N_26466,N_26231,N_26213);
nor U26467 (N_26467,N_26285,N_26228);
xor U26468 (N_26468,N_26378,N_26389);
xor U26469 (N_26469,N_26272,N_26286);
or U26470 (N_26470,N_26346,N_26262);
xnor U26471 (N_26471,N_26230,N_26303);
and U26472 (N_26472,N_26374,N_26394);
xnor U26473 (N_26473,N_26290,N_26315);
xor U26474 (N_26474,N_26390,N_26381);
nor U26475 (N_26475,N_26252,N_26312);
nand U26476 (N_26476,N_26302,N_26375);
xnor U26477 (N_26477,N_26353,N_26365);
or U26478 (N_26478,N_26277,N_26334);
and U26479 (N_26479,N_26379,N_26354);
xnor U26480 (N_26480,N_26227,N_26238);
nor U26481 (N_26481,N_26214,N_26217);
xor U26482 (N_26482,N_26288,N_26298);
xnor U26483 (N_26483,N_26339,N_26316);
nor U26484 (N_26484,N_26244,N_26264);
and U26485 (N_26485,N_26347,N_26368);
nor U26486 (N_26486,N_26216,N_26205);
nor U26487 (N_26487,N_26314,N_26332);
and U26488 (N_26488,N_26360,N_26202);
and U26489 (N_26489,N_26295,N_26226);
or U26490 (N_26490,N_26325,N_26229);
xnor U26491 (N_26491,N_26225,N_26294);
nand U26492 (N_26492,N_26208,N_26212);
or U26493 (N_26493,N_26241,N_26307);
xnor U26494 (N_26494,N_26292,N_26246);
xnor U26495 (N_26495,N_26383,N_26323);
xor U26496 (N_26496,N_26329,N_26350);
and U26497 (N_26497,N_26249,N_26255);
and U26498 (N_26498,N_26279,N_26351);
nor U26499 (N_26499,N_26275,N_26345);
and U26500 (N_26500,N_26359,N_26235);
or U26501 (N_26501,N_26291,N_26352);
xnor U26502 (N_26502,N_26264,N_26337);
nor U26503 (N_26503,N_26390,N_26335);
and U26504 (N_26504,N_26249,N_26202);
and U26505 (N_26505,N_26263,N_26326);
or U26506 (N_26506,N_26318,N_26324);
xnor U26507 (N_26507,N_26301,N_26243);
nand U26508 (N_26508,N_26291,N_26262);
and U26509 (N_26509,N_26348,N_26294);
or U26510 (N_26510,N_26342,N_26345);
or U26511 (N_26511,N_26365,N_26328);
nor U26512 (N_26512,N_26303,N_26360);
xor U26513 (N_26513,N_26310,N_26311);
and U26514 (N_26514,N_26211,N_26226);
nor U26515 (N_26515,N_26384,N_26332);
xnor U26516 (N_26516,N_26285,N_26372);
and U26517 (N_26517,N_26348,N_26255);
and U26518 (N_26518,N_26308,N_26278);
or U26519 (N_26519,N_26303,N_26330);
nor U26520 (N_26520,N_26316,N_26284);
nand U26521 (N_26521,N_26265,N_26314);
xor U26522 (N_26522,N_26201,N_26237);
and U26523 (N_26523,N_26255,N_26211);
or U26524 (N_26524,N_26391,N_26260);
and U26525 (N_26525,N_26320,N_26307);
or U26526 (N_26526,N_26378,N_26209);
nor U26527 (N_26527,N_26369,N_26233);
or U26528 (N_26528,N_26380,N_26302);
nand U26529 (N_26529,N_26270,N_26388);
or U26530 (N_26530,N_26216,N_26388);
xnor U26531 (N_26531,N_26325,N_26283);
nor U26532 (N_26532,N_26249,N_26325);
xor U26533 (N_26533,N_26395,N_26388);
and U26534 (N_26534,N_26323,N_26267);
xor U26535 (N_26535,N_26319,N_26221);
and U26536 (N_26536,N_26210,N_26349);
xnor U26537 (N_26537,N_26327,N_26348);
xnor U26538 (N_26538,N_26370,N_26219);
or U26539 (N_26539,N_26214,N_26286);
nor U26540 (N_26540,N_26243,N_26283);
and U26541 (N_26541,N_26267,N_26272);
nand U26542 (N_26542,N_26371,N_26339);
or U26543 (N_26543,N_26249,N_26286);
and U26544 (N_26544,N_26332,N_26329);
or U26545 (N_26545,N_26229,N_26322);
or U26546 (N_26546,N_26388,N_26202);
or U26547 (N_26547,N_26250,N_26206);
nand U26548 (N_26548,N_26283,N_26311);
or U26549 (N_26549,N_26347,N_26294);
nor U26550 (N_26550,N_26387,N_26239);
or U26551 (N_26551,N_26210,N_26360);
nand U26552 (N_26552,N_26353,N_26262);
xor U26553 (N_26553,N_26368,N_26352);
nor U26554 (N_26554,N_26258,N_26391);
or U26555 (N_26555,N_26323,N_26395);
xnor U26556 (N_26556,N_26228,N_26208);
nor U26557 (N_26557,N_26259,N_26223);
or U26558 (N_26558,N_26237,N_26319);
or U26559 (N_26559,N_26312,N_26327);
nor U26560 (N_26560,N_26342,N_26278);
nand U26561 (N_26561,N_26222,N_26263);
or U26562 (N_26562,N_26384,N_26347);
and U26563 (N_26563,N_26221,N_26343);
or U26564 (N_26564,N_26237,N_26205);
or U26565 (N_26565,N_26203,N_26234);
nor U26566 (N_26566,N_26389,N_26201);
xnor U26567 (N_26567,N_26364,N_26214);
nand U26568 (N_26568,N_26204,N_26314);
or U26569 (N_26569,N_26305,N_26209);
nor U26570 (N_26570,N_26238,N_26218);
nor U26571 (N_26571,N_26387,N_26236);
or U26572 (N_26572,N_26256,N_26326);
nand U26573 (N_26573,N_26257,N_26206);
nor U26574 (N_26574,N_26258,N_26340);
xor U26575 (N_26575,N_26213,N_26289);
nor U26576 (N_26576,N_26295,N_26248);
nand U26577 (N_26577,N_26286,N_26221);
or U26578 (N_26578,N_26360,N_26364);
and U26579 (N_26579,N_26255,N_26304);
nand U26580 (N_26580,N_26298,N_26360);
nand U26581 (N_26581,N_26379,N_26395);
or U26582 (N_26582,N_26277,N_26349);
nor U26583 (N_26583,N_26361,N_26335);
and U26584 (N_26584,N_26332,N_26399);
and U26585 (N_26585,N_26375,N_26292);
xnor U26586 (N_26586,N_26254,N_26360);
and U26587 (N_26587,N_26367,N_26282);
xor U26588 (N_26588,N_26273,N_26341);
and U26589 (N_26589,N_26296,N_26354);
and U26590 (N_26590,N_26307,N_26208);
nand U26591 (N_26591,N_26325,N_26344);
nor U26592 (N_26592,N_26368,N_26369);
xor U26593 (N_26593,N_26263,N_26378);
or U26594 (N_26594,N_26307,N_26334);
nor U26595 (N_26595,N_26331,N_26211);
nand U26596 (N_26596,N_26248,N_26301);
nand U26597 (N_26597,N_26312,N_26285);
xnor U26598 (N_26598,N_26295,N_26255);
nor U26599 (N_26599,N_26279,N_26330);
and U26600 (N_26600,N_26416,N_26511);
and U26601 (N_26601,N_26514,N_26467);
nand U26602 (N_26602,N_26487,N_26559);
xor U26603 (N_26603,N_26541,N_26579);
nor U26604 (N_26604,N_26540,N_26567);
xnor U26605 (N_26605,N_26476,N_26545);
and U26606 (N_26606,N_26455,N_26546);
and U26607 (N_26607,N_26493,N_26488);
nor U26608 (N_26608,N_26535,N_26562);
nand U26609 (N_26609,N_26417,N_26531);
or U26610 (N_26610,N_26402,N_26438);
or U26611 (N_26611,N_26563,N_26442);
nor U26612 (N_26612,N_26581,N_26549);
or U26613 (N_26613,N_26480,N_26586);
nor U26614 (N_26614,N_26453,N_26403);
nand U26615 (N_26615,N_26451,N_26406);
nor U26616 (N_26616,N_26461,N_26484);
and U26617 (N_26617,N_26483,N_26407);
or U26618 (N_26618,N_26552,N_26597);
xor U26619 (N_26619,N_26430,N_26570);
and U26620 (N_26620,N_26495,N_26459);
xnor U26621 (N_26621,N_26457,N_26526);
xor U26622 (N_26622,N_26513,N_26469);
or U26623 (N_26623,N_26536,N_26470);
and U26624 (N_26624,N_26528,N_26413);
or U26625 (N_26625,N_26422,N_26419);
and U26626 (N_26626,N_26569,N_26414);
nand U26627 (N_26627,N_26598,N_26582);
and U26628 (N_26628,N_26596,N_26449);
or U26629 (N_26629,N_26435,N_26491);
xor U26630 (N_26630,N_26557,N_26446);
or U26631 (N_26631,N_26599,N_26524);
or U26632 (N_26632,N_26441,N_26580);
xnor U26633 (N_26633,N_26590,N_26516);
nand U26634 (N_26634,N_26423,N_26592);
nor U26635 (N_26635,N_26421,N_26454);
or U26636 (N_26636,N_26431,N_26492);
nor U26637 (N_26637,N_26415,N_26497);
and U26638 (N_26638,N_26527,N_26517);
xor U26639 (N_26639,N_26444,N_26564);
or U26640 (N_26640,N_26412,N_26595);
nand U26641 (N_26641,N_26534,N_26588);
and U26642 (N_26642,N_26505,N_26466);
xor U26643 (N_26643,N_26477,N_26523);
nand U26644 (N_26644,N_26464,N_26481);
or U26645 (N_26645,N_26578,N_26479);
or U26646 (N_26646,N_26418,N_26452);
or U26647 (N_26647,N_26566,N_26560);
or U26648 (N_26648,N_26400,N_26472);
or U26649 (N_26649,N_26556,N_26542);
or U26650 (N_26650,N_26518,N_26428);
or U26651 (N_26651,N_26522,N_26551);
xor U26652 (N_26652,N_26494,N_26420);
or U26653 (N_26653,N_26520,N_26499);
or U26654 (N_26654,N_26489,N_26589);
and U26655 (N_26655,N_26445,N_26571);
nand U26656 (N_26656,N_26490,N_26515);
and U26657 (N_26657,N_26486,N_26425);
nor U26658 (N_26658,N_26574,N_26568);
nor U26659 (N_26659,N_26500,N_26573);
nor U26660 (N_26660,N_26496,N_26533);
nor U26661 (N_26661,N_26440,N_26553);
and U26662 (N_26662,N_26474,N_26507);
xnor U26663 (N_26663,N_26501,N_26432);
and U26664 (N_26664,N_26429,N_26539);
or U26665 (N_26665,N_26424,N_26555);
nand U26666 (N_26666,N_26405,N_26576);
nor U26667 (N_26667,N_26565,N_26434);
or U26668 (N_26668,N_26519,N_26550);
or U26669 (N_26669,N_26575,N_26538);
xnor U26670 (N_26670,N_26525,N_26506);
nor U26671 (N_26671,N_26585,N_26437);
xor U26672 (N_26672,N_26404,N_26594);
nand U26673 (N_26673,N_26577,N_26532);
nor U26674 (N_26674,N_26537,N_26561);
and U26675 (N_26675,N_26572,N_26458);
and U26676 (N_26676,N_26554,N_26544);
or U26677 (N_26677,N_26529,N_26471);
xor U26678 (N_26678,N_26460,N_26478);
and U26679 (N_26679,N_26468,N_26401);
nor U26680 (N_26680,N_26485,N_26548);
nor U26681 (N_26681,N_26512,N_26558);
xnor U26682 (N_26682,N_26593,N_26502);
nand U26683 (N_26683,N_26587,N_26427);
nor U26684 (N_26684,N_26436,N_26462);
xnor U26685 (N_26685,N_26473,N_26433);
nand U26686 (N_26686,N_26410,N_26503);
and U26687 (N_26687,N_26530,N_26508);
nand U26688 (N_26688,N_26463,N_26482);
nand U26689 (N_26689,N_26475,N_26504);
xnor U26690 (N_26690,N_26408,N_26426);
and U26691 (N_26691,N_26443,N_26584);
xnor U26692 (N_26692,N_26543,N_26509);
xnor U26693 (N_26693,N_26510,N_26465);
nor U26694 (N_26694,N_26547,N_26583);
and U26695 (N_26695,N_26521,N_26411);
and U26696 (N_26696,N_26450,N_26447);
nor U26697 (N_26697,N_26456,N_26448);
nand U26698 (N_26698,N_26498,N_26439);
or U26699 (N_26699,N_26409,N_26591);
nor U26700 (N_26700,N_26535,N_26581);
nor U26701 (N_26701,N_26565,N_26529);
and U26702 (N_26702,N_26574,N_26413);
xnor U26703 (N_26703,N_26455,N_26514);
or U26704 (N_26704,N_26427,N_26474);
or U26705 (N_26705,N_26549,N_26567);
xor U26706 (N_26706,N_26440,N_26522);
xor U26707 (N_26707,N_26406,N_26527);
nand U26708 (N_26708,N_26489,N_26407);
xor U26709 (N_26709,N_26424,N_26458);
xnor U26710 (N_26710,N_26424,N_26561);
and U26711 (N_26711,N_26479,N_26507);
nand U26712 (N_26712,N_26512,N_26590);
nor U26713 (N_26713,N_26465,N_26516);
xor U26714 (N_26714,N_26426,N_26578);
nand U26715 (N_26715,N_26506,N_26515);
and U26716 (N_26716,N_26532,N_26427);
nand U26717 (N_26717,N_26517,N_26538);
xor U26718 (N_26718,N_26511,N_26481);
and U26719 (N_26719,N_26478,N_26526);
and U26720 (N_26720,N_26422,N_26490);
xnor U26721 (N_26721,N_26463,N_26478);
nor U26722 (N_26722,N_26492,N_26421);
or U26723 (N_26723,N_26421,N_26530);
nand U26724 (N_26724,N_26466,N_26547);
xnor U26725 (N_26725,N_26474,N_26505);
xor U26726 (N_26726,N_26566,N_26575);
nor U26727 (N_26727,N_26521,N_26512);
or U26728 (N_26728,N_26572,N_26562);
xnor U26729 (N_26729,N_26494,N_26450);
or U26730 (N_26730,N_26506,N_26590);
and U26731 (N_26731,N_26492,N_26583);
and U26732 (N_26732,N_26483,N_26586);
nor U26733 (N_26733,N_26448,N_26595);
or U26734 (N_26734,N_26578,N_26533);
nand U26735 (N_26735,N_26444,N_26545);
xor U26736 (N_26736,N_26437,N_26422);
nor U26737 (N_26737,N_26462,N_26434);
nand U26738 (N_26738,N_26447,N_26489);
and U26739 (N_26739,N_26435,N_26544);
nand U26740 (N_26740,N_26590,N_26522);
nand U26741 (N_26741,N_26421,N_26550);
and U26742 (N_26742,N_26544,N_26456);
nand U26743 (N_26743,N_26560,N_26454);
nor U26744 (N_26744,N_26588,N_26552);
or U26745 (N_26745,N_26475,N_26454);
and U26746 (N_26746,N_26478,N_26501);
nor U26747 (N_26747,N_26484,N_26535);
xnor U26748 (N_26748,N_26441,N_26426);
xnor U26749 (N_26749,N_26458,N_26559);
or U26750 (N_26750,N_26518,N_26430);
xor U26751 (N_26751,N_26445,N_26564);
xor U26752 (N_26752,N_26563,N_26468);
xor U26753 (N_26753,N_26509,N_26588);
nor U26754 (N_26754,N_26427,N_26455);
and U26755 (N_26755,N_26552,N_26596);
nand U26756 (N_26756,N_26444,N_26414);
nand U26757 (N_26757,N_26432,N_26424);
or U26758 (N_26758,N_26521,N_26536);
or U26759 (N_26759,N_26575,N_26452);
nor U26760 (N_26760,N_26436,N_26468);
nand U26761 (N_26761,N_26576,N_26431);
or U26762 (N_26762,N_26576,N_26566);
xnor U26763 (N_26763,N_26469,N_26454);
xnor U26764 (N_26764,N_26538,N_26477);
xnor U26765 (N_26765,N_26481,N_26564);
xor U26766 (N_26766,N_26425,N_26570);
nand U26767 (N_26767,N_26595,N_26431);
nor U26768 (N_26768,N_26436,N_26402);
nor U26769 (N_26769,N_26477,N_26488);
xnor U26770 (N_26770,N_26493,N_26593);
nand U26771 (N_26771,N_26573,N_26513);
nand U26772 (N_26772,N_26505,N_26513);
nand U26773 (N_26773,N_26514,N_26585);
nor U26774 (N_26774,N_26598,N_26428);
nand U26775 (N_26775,N_26548,N_26420);
xor U26776 (N_26776,N_26489,N_26425);
xor U26777 (N_26777,N_26473,N_26534);
xor U26778 (N_26778,N_26472,N_26521);
nor U26779 (N_26779,N_26430,N_26464);
nand U26780 (N_26780,N_26427,N_26557);
or U26781 (N_26781,N_26558,N_26481);
xor U26782 (N_26782,N_26572,N_26411);
xor U26783 (N_26783,N_26530,N_26465);
nor U26784 (N_26784,N_26428,N_26586);
and U26785 (N_26785,N_26400,N_26578);
nor U26786 (N_26786,N_26530,N_26501);
and U26787 (N_26787,N_26465,N_26420);
nand U26788 (N_26788,N_26552,N_26469);
xnor U26789 (N_26789,N_26404,N_26486);
or U26790 (N_26790,N_26543,N_26584);
nand U26791 (N_26791,N_26572,N_26529);
xnor U26792 (N_26792,N_26408,N_26503);
nor U26793 (N_26793,N_26452,N_26584);
or U26794 (N_26794,N_26500,N_26555);
nor U26795 (N_26795,N_26488,N_26579);
and U26796 (N_26796,N_26504,N_26417);
nand U26797 (N_26797,N_26492,N_26406);
nor U26798 (N_26798,N_26442,N_26554);
nand U26799 (N_26799,N_26498,N_26479);
nor U26800 (N_26800,N_26670,N_26771);
and U26801 (N_26801,N_26604,N_26648);
nor U26802 (N_26802,N_26763,N_26664);
nor U26803 (N_26803,N_26762,N_26674);
and U26804 (N_26804,N_26779,N_26754);
xor U26805 (N_26805,N_26718,N_26743);
nand U26806 (N_26806,N_26736,N_26746);
and U26807 (N_26807,N_26642,N_26730);
nand U26808 (N_26808,N_26621,N_26678);
xnor U26809 (N_26809,N_26798,N_26715);
xnor U26810 (N_26810,N_26696,N_26645);
xor U26811 (N_26811,N_26729,N_26601);
xor U26812 (N_26812,N_26688,N_26697);
or U26813 (N_26813,N_26778,N_26727);
xnor U26814 (N_26814,N_26738,N_26704);
and U26815 (N_26815,N_26672,N_26711);
nand U26816 (N_26816,N_26745,N_26782);
xnor U26817 (N_26817,N_26628,N_26685);
xor U26818 (N_26818,N_26787,N_26695);
and U26819 (N_26819,N_26673,N_26653);
or U26820 (N_26820,N_26747,N_26796);
nand U26821 (N_26821,N_26629,N_26631);
or U26822 (N_26822,N_26622,N_26749);
xnor U26823 (N_26823,N_26777,N_26692);
nor U26824 (N_26824,N_26789,N_26658);
and U26825 (N_26825,N_26781,N_26624);
and U26826 (N_26826,N_26623,N_26775);
xor U26827 (N_26827,N_26660,N_26687);
and U26828 (N_26828,N_26752,N_26773);
nand U26829 (N_26829,N_26799,N_26740);
nor U26830 (N_26830,N_26683,N_26647);
xor U26831 (N_26831,N_26791,N_26641);
nor U26832 (N_26832,N_26659,N_26657);
or U26833 (N_26833,N_26735,N_26681);
and U26834 (N_26834,N_26783,N_26759);
nand U26835 (N_26835,N_26668,N_26793);
nand U26836 (N_26836,N_26689,N_26615);
nor U26837 (N_26837,N_26768,N_26691);
nor U26838 (N_26838,N_26760,N_26712);
or U26839 (N_26839,N_26675,N_26603);
nor U26840 (N_26840,N_26734,N_26679);
xnor U26841 (N_26841,N_26774,N_26717);
and U26842 (N_26842,N_26701,N_26721);
nand U26843 (N_26843,N_26635,N_26757);
nand U26844 (N_26844,N_26677,N_26665);
xnor U26845 (N_26845,N_26731,N_26723);
nand U26846 (N_26846,N_26707,N_26619);
nor U26847 (N_26847,N_26656,N_26710);
nor U26848 (N_26848,N_26652,N_26609);
and U26849 (N_26849,N_26766,N_26784);
xor U26850 (N_26850,N_26726,N_26769);
or U26851 (N_26851,N_26714,N_26719);
and U26852 (N_26852,N_26608,N_26680);
and U26853 (N_26853,N_26786,N_26669);
and U26854 (N_26854,N_26632,N_26755);
nand U26855 (N_26855,N_26698,N_26770);
xor U26856 (N_26856,N_26600,N_26722);
or U26857 (N_26857,N_26785,N_26612);
or U26858 (N_26858,N_26750,N_26613);
nand U26859 (N_26859,N_26767,N_26790);
or U26860 (N_26860,N_26666,N_26686);
or U26861 (N_26861,N_26741,N_26764);
nand U26862 (N_26862,N_26662,N_26617);
or U26863 (N_26863,N_26737,N_26667);
xnor U26864 (N_26864,N_26797,N_26765);
and U26865 (N_26865,N_26794,N_26690);
nand U26866 (N_26866,N_26616,N_26607);
nand U26867 (N_26867,N_26699,N_26702);
and U26868 (N_26868,N_26682,N_26788);
or U26869 (N_26869,N_26630,N_26761);
nand U26870 (N_26870,N_26606,N_26654);
nor U26871 (N_26871,N_26627,N_26694);
nor U26872 (N_26872,N_26728,N_26753);
xnor U26873 (N_26873,N_26716,N_26684);
nand U26874 (N_26874,N_26739,N_26639);
xor U26875 (N_26875,N_26671,N_26733);
nor U26876 (N_26876,N_26638,N_26643);
nor U26877 (N_26877,N_26725,N_26618);
xor U26878 (N_26878,N_26602,N_26661);
and U26879 (N_26879,N_26742,N_26676);
or U26880 (N_26880,N_26700,N_26634);
nand U26881 (N_26881,N_26795,N_26644);
nor U26882 (N_26882,N_26614,N_26703);
nor U26883 (N_26883,N_26776,N_26772);
and U26884 (N_26884,N_26625,N_26708);
or U26885 (N_26885,N_26792,N_26751);
xor U26886 (N_26886,N_26637,N_26705);
xnor U26887 (N_26887,N_26756,N_26605);
or U26888 (N_26888,N_26732,N_26713);
or U26889 (N_26889,N_26626,N_26748);
or U26890 (N_26890,N_26650,N_26693);
xnor U26891 (N_26891,N_26651,N_26724);
nor U26892 (N_26892,N_26709,N_26620);
nand U26893 (N_26893,N_26720,N_26758);
nand U26894 (N_26894,N_26611,N_26780);
xor U26895 (N_26895,N_26610,N_26663);
nor U26896 (N_26896,N_26636,N_26655);
nand U26897 (N_26897,N_26744,N_26649);
or U26898 (N_26898,N_26706,N_26646);
or U26899 (N_26899,N_26633,N_26640);
nand U26900 (N_26900,N_26655,N_26617);
or U26901 (N_26901,N_26754,N_26706);
or U26902 (N_26902,N_26749,N_26695);
nand U26903 (N_26903,N_26612,N_26768);
nor U26904 (N_26904,N_26729,N_26722);
and U26905 (N_26905,N_26674,N_26625);
xnor U26906 (N_26906,N_26726,N_26657);
nand U26907 (N_26907,N_26747,N_26678);
xnor U26908 (N_26908,N_26711,N_26740);
nor U26909 (N_26909,N_26603,N_26799);
nand U26910 (N_26910,N_26770,N_26694);
xor U26911 (N_26911,N_26629,N_26792);
nand U26912 (N_26912,N_26763,N_26792);
and U26913 (N_26913,N_26797,N_26618);
nand U26914 (N_26914,N_26756,N_26664);
nand U26915 (N_26915,N_26787,N_26630);
and U26916 (N_26916,N_26722,N_26701);
nand U26917 (N_26917,N_26617,N_26752);
nand U26918 (N_26918,N_26672,N_26638);
and U26919 (N_26919,N_26698,N_26739);
and U26920 (N_26920,N_26671,N_26633);
xor U26921 (N_26921,N_26777,N_26624);
and U26922 (N_26922,N_26672,N_26780);
nor U26923 (N_26923,N_26671,N_26706);
and U26924 (N_26924,N_26651,N_26796);
xor U26925 (N_26925,N_26734,N_26711);
nand U26926 (N_26926,N_26605,N_26749);
nor U26927 (N_26927,N_26697,N_26752);
or U26928 (N_26928,N_26689,N_26639);
nor U26929 (N_26929,N_26626,N_26751);
xnor U26930 (N_26930,N_26748,N_26744);
xor U26931 (N_26931,N_26669,N_26628);
and U26932 (N_26932,N_26638,N_26695);
and U26933 (N_26933,N_26787,N_26716);
or U26934 (N_26934,N_26670,N_26705);
nor U26935 (N_26935,N_26760,N_26762);
nand U26936 (N_26936,N_26748,N_26722);
nor U26937 (N_26937,N_26713,N_26723);
nor U26938 (N_26938,N_26607,N_26780);
xor U26939 (N_26939,N_26664,N_26674);
nand U26940 (N_26940,N_26736,N_26687);
or U26941 (N_26941,N_26651,N_26646);
nor U26942 (N_26942,N_26775,N_26688);
nand U26943 (N_26943,N_26721,N_26637);
nor U26944 (N_26944,N_26629,N_26640);
or U26945 (N_26945,N_26709,N_26675);
xor U26946 (N_26946,N_26778,N_26646);
nor U26947 (N_26947,N_26766,N_26643);
or U26948 (N_26948,N_26622,N_26670);
nor U26949 (N_26949,N_26656,N_26707);
and U26950 (N_26950,N_26678,N_26656);
and U26951 (N_26951,N_26642,N_26685);
nand U26952 (N_26952,N_26642,N_26672);
and U26953 (N_26953,N_26667,N_26751);
nor U26954 (N_26954,N_26629,N_26762);
xor U26955 (N_26955,N_26701,N_26668);
nand U26956 (N_26956,N_26621,N_26635);
xnor U26957 (N_26957,N_26643,N_26654);
or U26958 (N_26958,N_26761,N_26691);
nor U26959 (N_26959,N_26630,N_26611);
xnor U26960 (N_26960,N_26715,N_26686);
xnor U26961 (N_26961,N_26770,N_26616);
nor U26962 (N_26962,N_26692,N_26653);
nor U26963 (N_26963,N_26643,N_26709);
nor U26964 (N_26964,N_26778,N_26724);
nand U26965 (N_26965,N_26647,N_26780);
nand U26966 (N_26966,N_26708,N_26742);
xnor U26967 (N_26967,N_26705,N_26612);
xor U26968 (N_26968,N_26711,N_26664);
and U26969 (N_26969,N_26708,N_26775);
or U26970 (N_26970,N_26627,N_26664);
or U26971 (N_26971,N_26750,N_26788);
and U26972 (N_26972,N_26620,N_26760);
nand U26973 (N_26973,N_26712,N_26763);
nor U26974 (N_26974,N_26777,N_26740);
or U26975 (N_26975,N_26686,N_26725);
or U26976 (N_26976,N_26757,N_26797);
nand U26977 (N_26977,N_26701,N_26646);
and U26978 (N_26978,N_26782,N_26789);
nand U26979 (N_26979,N_26737,N_26726);
nor U26980 (N_26980,N_26770,N_26738);
nor U26981 (N_26981,N_26750,N_26657);
nor U26982 (N_26982,N_26749,N_26672);
and U26983 (N_26983,N_26755,N_26605);
or U26984 (N_26984,N_26679,N_26725);
xnor U26985 (N_26985,N_26664,N_26677);
nand U26986 (N_26986,N_26661,N_26689);
nor U26987 (N_26987,N_26773,N_26738);
xor U26988 (N_26988,N_26693,N_26655);
xnor U26989 (N_26989,N_26705,N_26617);
xor U26990 (N_26990,N_26699,N_26677);
nor U26991 (N_26991,N_26787,N_26613);
or U26992 (N_26992,N_26634,N_26746);
nand U26993 (N_26993,N_26784,N_26672);
nor U26994 (N_26994,N_26648,N_26734);
and U26995 (N_26995,N_26773,N_26663);
nor U26996 (N_26996,N_26656,N_26780);
nand U26997 (N_26997,N_26668,N_26652);
xor U26998 (N_26998,N_26728,N_26719);
xor U26999 (N_26999,N_26639,N_26766);
nor U27000 (N_27000,N_26962,N_26837);
and U27001 (N_27001,N_26839,N_26868);
and U27002 (N_27002,N_26831,N_26984);
nor U27003 (N_27003,N_26976,N_26825);
xnor U27004 (N_27004,N_26854,N_26987);
xnor U27005 (N_27005,N_26930,N_26895);
nand U27006 (N_27006,N_26832,N_26817);
nor U27007 (N_27007,N_26820,N_26904);
nand U27008 (N_27008,N_26999,N_26886);
or U27009 (N_27009,N_26857,N_26993);
nand U27010 (N_27010,N_26897,N_26815);
and U27011 (N_27011,N_26804,N_26823);
xnor U27012 (N_27012,N_26898,N_26903);
nand U27013 (N_27013,N_26953,N_26992);
nor U27014 (N_27014,N_26950,N_26920);
or U27015 (N_27015,N_26890,N_26805);
xor U27016 (N_27016,N_26935,N_26860);
and U27017 (N_27017,N_26906,N_26977);
nor U27018 (N_27018,N_26961,N_26916);
nand U27019 (N_27019,N_26814,N_26969);
nor U27020 (N_27020,N_26972,N_26866);
nor U27021 (N_27021,N_26818,N_26952);
nor U27022 (N_27022,N_26913,N_26970);
and U27023 (N_27023,N_26840,N_26864);
nand U27024 (N_27024,N_26939,N_26994);
nor U27025 (N_27025,N_26981,N_26990);
nand U27026 (N_27026,N_26967,N_26912);
nand U27027 (N_27027,N_26947,N_26809);
nand U27028 (N_27028,N_26963,N_26883);
xor U27029 (N_27029,N_26841,N_26836);
nor U27030 (N_27030,N_26980,N_26813);
and U27031 (N_27031,N_26936,N_26915);
or U27032 (N_27032,N_26975,N_26870);
nor U27033 (N_27033,N_26941,N_26811);
or U27034 (N_27034,N_26905,N_26964);
and U27035 (N_27035,N_26945,N_26900);
and U27036 (N_27036,N_26826,N_26867);
nor U27037 (N_27037,N_26810,N_26989);
xor U27038 (N_27038,N_26803,N_26958);
nor U27039 (N_27039,N_26991,N_26982);
and U27040 (N_27040,N_26908,N_26957);
or U27041 (N_27041,N_26948,N_26933);
xor U27042 (N_27042,N_26901,N_26943);
and U27043 (N_27043,N_26808,N_26812);
nand U27044 (N_27044,N_26855,N_26914);
and U27045 (N_27045,N_26858,N_26853);
nand U27046 (N_27046,N_26917,N_26835);
and U27047 (N_27047,N_26891,N_26986);
and U27048 (N_27048,N_26838,N_26876);
and U27049 (N_27049,N_26918,N_26988);
or U27050 (N_27050,N_26848,N_26956);
and U27051 (N_27051,N_26931,N_26910);
xnor U27052 (N_27052,N_26927,N_26872);
nor U27053 (N_27053,N_26965,N_26851);
xnor U27054 (N_27054,N_26859,N_26802);
nand U27055 (N_27055,N_26877,N_26925);
nand U27056 (N_27056,N_26911,N_26819);
or U27057 (N_27057,N_26899,N_26959);
and U27058 (N_27058,N_26827,N_26842);
or U27059 (N_27059,N_26955,N_26896);
or U27060 (N_27060,N_26806,N_26954);
and U27061 (N_27061,N_26882,N_26816);
xnor U27062 (N_27062,N_26881,N_26928);
and U27063 (N_27063,N_26834,N_26924);
nor U27064 (N_27064,N_26873,N_26887);
nor U27065 (N_27065,N_26833,N_26919);
nor U27066 (N_27066,N_26829,N_26862);
xnor U27067 (N_27067,N_26878,N_26879);
and U27068 (N_27068,N_26949,N_26934);
nand U27069 (N_27069,N_26971,N_26937);
xnor U27070 (N_27070,N_26946,N_26863);
and U27071 (N_27071,N_26940,N_26995);
nand U27072 (N_27072,N_26907,N_26997);
and U27073 (N_27073,N_26944,N_26996);
nor U27074 (N_27074,N_26824,N_26885);
or U27075 (N_27075,N_26998,N_26978);
nor U27076 (N_27076,N_26843,N_26921);
or U27077 (N_27077,N_26846,N_26894);
or U27078 (N_27078,N_26974,N_26985);
xor U27079 (N_27079,N_26902,N_26801);
and U27080 (N_27080,N_26888,N_26884);
and U27081 (N_27081,N_26929,N_26830);
nor U27082 (N_27082,N_26951,N_26923);
or U27083 (N_27083,N_26807,N_26821);
and U27084 (N_27084,N_26880,N_26889);
or U27085 (N_27085,N_26800,N_26850);
nand U27086 (N_27086,N_26844,N_26874);
and U27087 (N_27087,N_26828,N_26852);
nor U27088 (N_27088,N_26871,N_26942);
and U27089 (N_27089,N_26875,N_26893);
nand U27090 (N_27090,N_26960,N_26845);
and U27091 (N_27091,N_26822,N_26847);
xnor U27092 (N_27092,N_26865,N_26892);
and U27093 (N_27093,N_26922,N_26983);
xnor U27094 (N_27094,N_26966,N_26968);
or U27095 (N_27095,N_26973,N_26849);
nand U27096 (N_27096,N_26926,N_26856);
and U27097 (N_27097,N_26979,N_26932);
and U27098 (N_27098,N_26861,N_26909);
nand U27099 (N_27099,N_26938,N_26869);
nor U27100 (N_27100,N_26848,N_26933);
nand U27101 (N_27101,N_26811,N_26945);
xor U27102 (N_27102,N_26835,N_26908);
nor U27103 (N_27103,N_26892,N_26826);
nand U27104 (N_27104,N_26958,N_26921);
or U27105 (N_27105,N_26956,N_26960);
xor U27106 (N_27106,N_26852,N_26873);
or U27107 (N_27107,N_26951,N_26809);
and U27108 (N_27108,N_26810,N_26942);
and U27109 (N_27109,N_26974,N_26833);
xnor U27110 (N_27110,N_26990,N_26950);
nand U27111 (N_27111,N_26884,N_26885);
nand U27112 (N_27112,N_26955,N_26870);
nand U27113 (N_27113,N_26802,N_26882);
nor U27114 (N_27114,N_26832,N_26914);
nor U27115 (N_27115,N_26849,N_26834);
nor U27116 (N_27116,N_26825,N_26845);
or U27117 (N_27117,N_26922,N_26837);
and U27118 (N_27118,N_26864,N_26848);
nor U27119 (N_27119,N_26827,N_26917);
xor U27120 (N_27120,N_26853,N_26966);
or U27121 (N_27121,N_26856,N_26999);
xor U27122 (N_27122,N_26997,N_26843);
nor U27123 (N_27123,N_26857,N_26949);
nor U27124 (N_27124,N_26986,N_26960);
nand U27125 (N_27125,N_26889,N_26975);
nand U27126 (N_27126,N_26836,N_26984);
or U27127 (N_27127,N_26880,N_26954);
and U27128 (N_27128,N_26844,N_26918);
xor U27129 (N_27129,N_26954,N_26967);
nor U27130 (N_27130,N_26941,N_26845);
nor U27131 (N_27131,N_26975,N_26955);
nand U27132 (N_27132,N_26905,N_26822);
nand U27133 (N_27133,N_26892,N_26882);
and U27134 (N_27134,N_26927,N_26960);
and U27135 (N_27135,N_26995,N_26941);
xnor U27136 (N_27136,N_26928,N_26927);
nor U27137 (N_27137,N_26858,N_26857);
and U27138 (N_27138,N_26898,N_26927);
or U27139 (N_27139,N_26948,N_26945);
xnor U27140 (N_27140,N_26938,N_26918);
nand U27141 (N_27141,N_26816,N_26962);
nand U27142 (N_27142,N_26875,N_26892);
xnor U27143 (N_27143,N_26983,N_26945);
nor U27144 (N_27144,N_26958,N_26848);
nand U27145 (N_27145,N_26895,N_26928);
and U27146 (N_27146,N_26915,N_26902);
xnor U27147 (N_27147,N_26969,N_26825);
or U27148 (N_27148,N_26824,N_26931);
or U27149 (N_27149,N_26971,N_26889);
nand U27150 (N_27150,N_26868,N_26840);
and U27151 (N_27151,N_26888,N_26942);
nor U27152 (N_27152,N_26927,N_26931);
nor U27153 (N_27153,N_26898,N_26834);
and U27154 (N_27154,N_26881,N_26919);
and U27155 (N_27155,N_26899,N_26923);
nor U27156 (N_27156,N_26837,N_26949);
nor U27157 (N_27157,N_26998,N_26908);
nand U27158 (N_27158,N_26982,N_26865);
or U27159 (N_27159,N_26894,N_26984);
or U27160 (N_27160,N_26897,N_26868);
nor U27161 (N_27161,N_26998,N_26892);
or U27162 (N_27162,N_26889,N_26808);
nand U27163 (N_27163,N_26980,N_26814);
xor U27164 (N_27164,N_26864,N_26905);
nor U27165 (N_27165,N_26927,N_26946);
or U27166 (N_27166,N_26974,N_26802);
nand U27167 (N_27167,N_26935,N_26991);
nand U27168 (N_27168,N_26827,N_26993);
nor U27169 (N_27169,N_26975,N_26985);
and U27170 (N_27170,N_26840,N_26947);
nor U27171 (N_27171,N_26855,N_26987);
nand U27172 (N_27172,N_26846,N_26866);
nand U27173 (N_27173,N_26978,N_26861);
xnor U27174 (N_27174,N_26972,N_26838);
or U27175 (N_27175,N_26803,N_26908);
xor U27176 (N_27176,N_26929,N_26907);
and U27177 (N_27177,N_26895,N_26919);
xnor U27178 (N_27178,N_26884,N_26995);
nand U27179 (N_27179,N_26852,N_26832);
nor U27180 (N_27180,N_26851,N_26836);
or U27181 (N_27181,N_26958,N_26820);
nand U27182 (N_27182,N_26832,N_26980);
xnor U27183 (N_27183,N_26953,N_26933);
and U27184 (N_27184,N_26831,N_26878);
nor U27185 (N_27185,N_26990,N_26905);
xnor U27186 (N_27186,N_26913,N_26827);
and U27187 (N_27187,N_26830,N_26906);
xnor U27188 (N_27188,N_26914,N_26955);
xor U27189 (N_27189,N_26961,N_26962);
nand U27190 (N_27190,N_26867,N_26914);
and U27191 (N_27191,N_26976,N_26803);
and U27192 (N_27192,N_26966,N_26889);
and U27193 (N_27193,N_26805,N_26904);
nor U27194 (N_27194,N_26937,N_26984);
nand U27195 (N_27195,N_26853,N_26814);
nor U27196 (N_27196,N_26914,N_26848);
or U27197 (N_27197,N_26926,N_26838);
and U27198 (N_27198,N_26895,N_26986);
nand U27199 (N_27199,N_26887,N_26946);
xnor U27200 (N_27200,N_27051,N_27167);
or U27201 (N_27201,N_27139,N_27042);
nand U27202 (N_27202,N_27125,N_27128);
and U27203 (N_27203,N_27100,N_27124);
and U27204 (N_27204,N_27151,N_27183);
or U27205 (N_27205,N_27014,N_27045);
nor U27206 (N_27206,N_27115,N_27095);
and U27207 (N_27207,N_27121,N_27054);
and U27208 (N_27208,N_27010,N_27111);
xor U27209 (N_27209,N_27182,N_27047);
and U27210 (N_27210,N_27005,N_27065);
or U27211 (N_27211,N_27110,N_27107);
and U27212 (N_27212,N_27052,N_27187);
nand U27213 (N_27213,N_27062,N_27039);
nor U27214 (N_27214,N_27163,N_27033);
nand U27215 (N_27215,N_27082,N_27023);
and U27216 (N_27216,N_27037,N_27024);
or U27217 (N_27217,N_27074,N_27123);
xor U27218 (N_27218,N_27008,N_27188);
or U27219 (N_27219,N_27034,N_27175);
and U27220 (N_27220,N_27056,N_27155);
nand U27221 (N_27221,N_27018,N_27021);
xnor U27222 (N_27222,N_27050,N_27126);
and U27223 (N_27223,N_27043,N_27105);
nor U27224 (N_27224,N_27081,N_27067);
nor U27225 (N_27225,N_27179,N_27011);
xor U27226 (N_27226,N_27150,N_27057);
xnor U27227 (N_27227,N_27009,N_27135);
nand U27228 (N_27228,N_27093,N_27104);
or U27229 (N_27229,N_27154,N_27132);
or U27230 (N_27230,N_27092,N_27156);
xnor U27231 (N_27231,N_27068,N_27177);
or U27232 (N_27232,N_27157,N_27075);
and U27233 (N_27233,N_27070,N_27015);
xnor U27234 (N_27234,N_27060,N_27036);
xnor U27235 (N_27235,N_27174,N_27134);
and U27236 (N_27236,N_27038,N_27198);
nand U27237 (N_27237,N_27020,N_27089);
nand U27238 (N_27238,N_27130,N_27149);
and U27239 (N_27239,N_27152,N_27181);
nand U27240 (N_27240,N_27066,N_27117);
and U27241 (N_27241,N_27145,N_27087);
xnor U27242 (N_27242,N_27098,N_27173);
xor U27243 (N_27243,N_27116,N_27186);
xor U27244 (N_27244,N_27129,N_27000);
nor U27245 (N_27245,N_27076,N_27166);
or U27246 (N_27246,N_27184,N_27073);
nor U27247 (N_27247,N_27178,N_27103);
nand U27248 (N_27248,N_27164,N_27078);
xnor U27249 (N_27249,N_27133,N_27171);
nor U27250 (N_27250,N_27180,N_27048);
xnor U27251 (N_27251,N_27141,N_27168);
or U27252 (N_27252,N_27106,N_27003);
nand U27253 (N_27253,N_27099,N_27119);
and U27254 (N_27254,N_27137,N_27025);
and U27255 (N_27255,N_27035,N_27153);
and U27256 (N_27256,N_27108,N_27120);
and U27257 (N_27257,N_27122,N_27061);
xnor U27258 (N_27258,N_27096,N_27160);
nor U27259 (N_27259,N_27088,N_27097);
or U27260 (N_27260,N_27138,N_27114);
or U27261 (N_27261,N_27113,N_27090);
xor U27262 (N_27262,N_27063,N_27165);
and U27263 (N_27263,N_27016,N_27118);
nand U27264 (N_27264,N_27053,N_27191);
and U27265 (N_27265,N_27029,N_27112);
xor U27266 (N_27266,N_27190,N_27072);
and U27267 (N_27267,N_27077,N_27169);
and U27268 (N_27268,N_27071,N_27196);
and U27269 (N_27269,N_27146,N_27109);
or U27270 (N_27270,N_27162,N_27026);
and U27271 (N_27271,N_27194,N_27199);
or U27272 (N_27272,N_27193,N_27147);
and U27273 (N_27273,N_27197,N_27161);
nor U27274 (N_27274,N_27004,N_27032);
nor U27275 (N_27275,N_27148,N_27158);
xnor U27276 (N_27276,N_27002,N_27086);
or U27277 (N_27277,N_27044,N_27080);
nor U27278 (N_27278,N_27136,N_27170);
and U27279 (N_27279,N_27144,N_27159);
and U27280 (N_27280,N_27085,N_27195);
or U27281 (N_27281,N_27028,N_27049);
nand U27282 (N_27282,N_27030,N_27006);
or U27283 (N_27283,N_27041,N_27046);
xor U27284 (N_27284,N_27007,N_27131);
or U27285 (N_27285,N_27185,N_27022);
xor U27286 (N_27286,N_27172,N_27140);
nand U27287 (N_27287,N_27013,N_27091);
nor U27288 (N_27288,N_27055,N_27102);
nor U27289 (N_27289,N_27127,N_27083);
and U27290 (N_27290,N_27012,N_27079);
xor U27291 (N_27291,N_27019,N_27192);
nand U27292 (N_27292,N_27142,N_27101);
xor U27293 (N_27293,N_27189,N_27064);
xnor U27294 (N_27294,N_27001,N_27143);
and U27295 (N_27295,N_27027,N_27031);
xor U27296 (N_27296,N_27069,N_27040);
and U27297 (N_27297,N_27017,N_27084);
or U27298 (N_27298,N_27176,N_27059);
xnor U27299 (N_27299,N_27094,N_27058);
xnor U27300 (N_27300,N_27124,N_27106);
xor U27301 (N_27301,N_27033,N_27095);
or U27302 (N_27302,N_27162,N_27092);
nor U27303 (N_27303,N_27012,N_27125);
and U27304 (N_27304,N_27063,N_27187);
nor U27305 (N_27305,N_27153,N_27069);
or U27306 (N_27306,N_27113,N_27051);
and U27307 (N_27307,N_27171,N_27195);
and U27308 (N_27308,N_27182,N_27078);
nand U27309 (N_27309,N_27176,N_27049);
or U27310 (N_27310,N_27197,N_27015);
and U27311 (N_27311,N_27165,N_27190);
or U27312 (N_27312,N_27131,N_27003);
or U27313 (N_27313,N_27050,N_27125);
and U27314 (N_27314,N_27157,N_27026);
or U27315 (N_27315,N_27108,N_27049);
or U27316 (N_27316,N_27101,N_27131);
and U27317 (N_27317,N_27158,N_27062);
and U27318 (N_27318,N_27117,N_27135);
and U27319 (N_27319,N_27144,N_27006);
or U27320 (N_27320,N_27028,N_27038);
nor U27321 (N_27321,N_27020,N_27101);
and U27322 (N_27322,N_27077,N_27112);
or U27323 (N_27323,N_27125,N_27027);
xor U27324 (N_27324,N_27036,N_27042);
xnor U27325 (N_27325,N_27088,N_27179);
xor U27326 (N_27326,N_27171,N_27153);
and U27327 (N_27327,N_27187,N_27199);
nor U27328 (N_27328,N_27006,N_27054);
nand U27329 (N_27329,N_27022,N_27196);
nor U27330 (N_27330,N_27198,N_27170);
and U27331 (N_27331,N_27129,N_27117);
nand U27332 (N_27332,N_27020,N_27033);
nand U27333 (N_27333,N_27157,N_27125);
or U27334 (N_27334,N_27123,N_27092);
nand U27335 (N_27335,N_27174,N_27116);
or U27336 (N_27336,N_27148,N_27193);
xnor U27337 (N_27337,N_27090,N_27148);
xor U27338 (N_27338,N_27012,N_27073);
xor U27339 (N_27339,N_27136,N_27196);
nor U27340 (N_27340,N_27142,N_27121);
nor U27341 (N_27341,N_27151,N_27121);
nor U27342 (N_27342,N_27126,N_27084);
nor U27343 (N_27343,N_27102,N_27128);
or U27344 (N_27344,N_27023,N_27053);
and U27345 (N_27345,N_27074,N_27189);
nand U27346 (N_27346,N_27128,N_27093);
nand U27347 (N_27347,N_27021,N_27034);
nand U27348 (N_27348,N_27099,N_27118);
xnor U27349 (N_27349,N_27043,N_27136);
xnor U27350 (N_27350,N_27166,N_27199);
or U27351 (N_27351,N_27074,N_27168);
and U27352 (N_27352,N_27066,N_27050);
nand U27353 (N_27353,N_27096,N_27149);
or U27354 (N_27354,N_27139,N_27070);
xor U27355 (N_27355,N_27115,N_27162);
nand U27356 (N_27356,N_27172,N_27068);
xor U27357 (N_27357,N_27145,N_27132);
nor U27358 (N_27358,N_27118,N_27158);
xnor U27359 (N_27359,N_27086,N_27187);
xnor U27360 (N_27360,N_27145,N_27072);
or U27361 (N_27361,N_27043,N_27157);
and U27362 (N_27362,N_27146,N_27183);
nand U27363 (N_27363,N_27022,N_27036);
and U27364 (N_27364,N_27007,N_27012);
and U27365 (N_27365,N_27097,N_27050);
xnor U27366 (N_27366,N_27174,N_27129);
nand U27367 (N_27367,N_27119,N_27130);
nor U27368 (N_27368,N_27144,N_27170);
nor U27369 (N_27369,N_27146,N_27101);
nand U27370 (N_27370,N_27123,N_27164);
nor U27371 (N_27371,N_27002,N_27097);
and U27372 (N_27372,N_27177,N_27133);
xor U27373 (N_27373,N_27046,N_27107);
nand U27374 (N_27374,N_27074,N_27102);
and U27375 (N_27375,N_27028,N_27060);
nand U27376 (N_27376,N_27002,N_27019);
or U27377 (N_27377,N_27185,N_27093);
and U27378 (N_27378,N_27155,N_27016);
xor U27379 (N_27379,N_27008,N_27121);
nand U27380 (N_27380,N_27125,N_27069);
nor U27381 (N_27381,N_27193,N_27199);
or U27382 (N_27382,N_27022,N_27124);
nor U27383 (N_27383,N_27026,N_27194);
xor U27384 (N_27384,N_27090,N_27025);
nand U27385 (N_27385,N_27026,N_27058);
nor U27386 (N_27386,N_27092,N_27197);
or U27387 (N_27387,N_27126,N_27014);
nor U27388 (N_27388,N_27166,N_27158);
nand U27389 (N_27389,N_27076,N_27015);
nor U27390 (N_27390,N_27194,N_27135);
nor U27391 (N_27391,N_27021,N_27138);
nor U27392 (N_27392,N_27004,N_27126);
and U27393 (N_27393,N_27055,N_27198);
or U27394 (N_27394,N_27162,N_27069);
and U27395 (N_27395,N_27115,N_27091);
xor U27396 (N_27396,N_27083,N_27167);
xor U27397 (N_27397,N_27014,N_27040);
nor U27398 (N_27398,N_27117,N_27178);
or U27399 (N_27399,N_27106,N_27095);
nor U27400 (N_27400,N_27351,N_27333);
or U27401 (N_27401,N_27372,N_27271);
or U27402 (N_27402,N_27380,N_27382);
xnor U27403 (N_27403,N_27209,N_27324);
nand U27404 (N_27404,N_27326,N_27303);
nand U27405 (N_27405,N_27389,N_27267);
and U27406 (N_27406,N_27205,N_27361);
and U27407 (N_27407,N_27338,N_27280);
nand U27408 (N_27408,N_27343,N_27386);
xnor U27409 (N_27409,N_27387,N_27376);
or U27410 (N_27410,N_27286,N_27366);
or U27411 (N_27411,N_27224,N_27287);
or U27412 (N_27412,N_27296,N_27260);
nand U27413 (N_27413,N_27395,N_27290);
nor U27414 (N_27414,N_27394,N_27342);
nor U27415 (N_27415,N_27231,N_27336);
and U27416 (N_27416,N_27306,N_27255);
xor U27417 (N_27417,N_27369,N_27327);
or U27418 (N_27418,N_27264,N_27308);
or U27419 (N_27419,N_27298,N_27200);
nor U27420 (N_27420,N_27302,N_27216);
nor U27421 (N_27421,N_27341,N_27232);
and U27422 (N_27422,N_27370,N_27230);
xor U27423 (N_27423,N_27334,N_27259);
nor U27424 (N_27424,N_27226,N_27360);
or U27425 (N_27425,N_27270,N_27277);
nor U27426 (N_27426,N_27385,N_27335);
nand U27427 (N_27427,N_27238,N_27330);
and U27428 (N_27428,N_27265,N_27381);
xor U27429 (N_27429,N_27348,N_27236);
nand U27430 (N_27430,N_27261,N_27268);
nand U27431 (N_27431,N_27263,N_27354);
nand U27432 (N_27432,N_27279,N_27337);
and U27433 (N_27433,N_27283,N_27397);
nor U27434 (N_27434,N_27352,N_27235);
nor U27435 (N_27435,N_27258,N_27241);
nor U27436 (N_27436,N_27344,N_27347);
and U27437 (N_27437,N_27392,N_27234);
nand U27438 (N_27438,N_27225,N_27318);
and U27439 (N_27439,N_27221,N_27213);
nor U27440 (N_27440,N_27291,N_27295);
and U27441 (N_27441,N_27275,N_27207);
nor U27442 (N_27442,N_27276,N_27349);
nand U27443 (N_27443,N_27304,N_27239);
and U27444 (N_27444,N_27251,N_27305);
nand U27445 (N_27445,N_27229,N_27374);
xnor U27446 (N_27446,N_27219,N_27293);
xnor U27447 (N_27447,N_27253,N_27204);
and U27448 (N_27448,N_27388,N_27383);
nand U27449 (N_27449,N_27240,N_27285);
or U27450 (N_27450,N_27294,N_27345);
and U27451 (N_27451,N_27399,N_27320);
and U27452 (N_27452,N_27365,N_27249);
nand U27453 (N_27453,N_27310,N_27362);
nor U27454 (N_27454,N_27307,N_27379);
nand U27455 (N_27455,N_27266,N_27273);
and U27456 (N_27456,N_27214,N_27319);
and U27457 (N_27457,N_27329,N_27206);
or U27458 (N_27458,N_27315,N_27218);
and U27459 (N_27459,N_27384,N_27247);
nand U27460 (N_27460,N_27313,N_27359);
nand U27461 (N_27461,N_27311,N_27377);
nor U27462 (N_27462,N_27299,N_27212);
nor U27463 (N_27463,N_27346,N_27201);
and U27464 (N_27464,N_27367,N_27284);
and U27465 (N_27465,N_27203,N_27242);
and U27466 (N_27466,N_27355,N_27391);
or U27467 (N_27467,N_27227,N_27222);
xnor U27468 (N_27468,N_27332,N_27350);
or U27469 (N_27469,N_27278,N_27254);
nand U27470 (N_27470,N_27373,N_27371);
or U27471 (N_27471,N_27390,N_27353);
xor U27472 (N_27472,N_27243,N_27237);
xor U27473 (N_27473,N_27357,N_27339);
or U27474 (N_27474,N_27257,N_27244);
xor U27475 (N_27475,N_27228,N_27262);
or U27476 (N_27476,N_27208,N_27398);
nand U27477 (N_27477,N_27250,N_27363);
and U27478 (N_27478,N_27328,N_27288);
xnor U27479 (N_27479,N_27245,N_27269);
nor U27480 (N_27480,N_27215,N_27309);
nor U27481 (N_27481,N_27211,N_27282);
xnor U27482 (N_27482,N_27246,N_27274);
or U27483 (N_27483,N_27340,N_27248);
and U27484 (N_27484,N_27223,N_27289);
xnor U27485 (N_27485,N_27321,N_27202);
or U27486 (N_27486,N_27233,N_27331);
nor U27487 (N_27487,N_27364,N_27317);
xnor U27488 (N_27488,N_27396,N_27316);
nor U27489 (N_27489,N_27272,N_27312);
or U27490 (N_27490,N_27356,N_27252);
or U27491 (N_27491,N_27292,N_27393);
xnor U27492 (N_27492,N_27375,N_27325);
and U27493 (N_27493,N_27297,N_27323);
xor U27494 (N_27494,N_27368,N_27314);
and U27495 (N_27495,N_27322,N_27301);
nand U27496 (N_27496,N_27300,N_27220);
xor U27497 (N_27497,N_27281,N_27256);
and U27498 (N_27498,N_27210,N_27378);
xnor U27499 (N_27499,N_27358,N_27217);
and U27500 (N_27500,N_27386,N_27341);
and U27501 (N_27501,N_27389,N_27231);
xor U27502 (N_27502,N_27357,N_27322);
nor U27503 (N_27503,N_27310,N_27351);
and U27504 (N_27504,N_27261,N_27391);
nand U27505 (N_27505,N_27359,N_27202);
or U27506 (N_27506,N_27211,N_27268);
xnor U27507 (N_27507,N_27303,N_27317);
or U27508 (N_27508,N_27390,N_27315);
or U27509 (N_27509,N_27333,N_27364);
and U27510 (N_27510,N_27330,N_27302);
nand U27511 (N_27511,N_27269,N_27379);
and U27512 (N_27512,N_27236,N_27305);
and U27513 (N_27513,N_27244,N_27206);
and U27514 (N_27514,N_27307,N_27384);
or U27515 (N_27515,N_27278,N_27382);
and U27516 (N_27516,N_27200,N_27206);
nor U27517 (N_27517,N_27348,N_27245);
nor U27518 (N_27518,N_27283,N_27336);
and U27519 (N_27519,N_27245,N_27305);
xor U27520 (N_27520,N_27328,N_27269);
nand U27521 (N_27521,N_27296,N_27325);
or U27522 (N_27522,N_27248,N_27306);
and U27523 (N_27523,N_27230,N_27226);
and U27524 (N_27524,N_27257,N_27307);
or U27525 (N_27525,N_27262,N_27243);
xnor U27526 (N_27526,N_27238,N_27387);
nor U27527 (N_27527,N_27337,N_27241);
or U27528 (N_27528,N_27205,N_27348);
nand U27529 (N_27529,N_27306,N_27204);
nand U27530 (N_27530,N_27316,N_27397);
nor U27531 (N_27531,N_27388,N_27305);
xor U27532 (N_27532,N_27303,N_27269);
or U27533 (N_27533,N_27259,N_27350);
and U27534 (N_27534,N_27225,N_27326);
xor U27535 (N_27535,N_27240,N_27219);
and U27536 (N_27536,N_27272,N_27328);
nand U27537 (N_27537,N_27351,N_27253);
nand U27538 (N_27538,N_27347,N_27204);
nand U27539 (N_27539,N_27352,N_27200);
nor U27540 (N_27540,N_27335,N_27377);
nor U27541 (N_27541,N_27373,N_27352);
xor U27542 (N_27542,N_27205,N_27208);
xnor U27543 (N_27543,N_27236,N_27242);
and U27544 (N_27544,N_27278,N_27277);
xnor U27545 (N_27545,N_27283,N_27310);
and U27546 (N_27546,N_27223,N_27269);
nand U27547 (N_27547,N_27388,N_27380);
or U27548 (N_27548,N_27378,N_27386);
xor U27549 (N_27549,N_27383,N_27396);
nor U27550 (N_27550,N_27292,N_27283);
or U27551 (N_27551,N_27301,N_27225);
xor U27552 (N_27552,N_27277,N_27276);
and U27553 (N_27553,N_27267,N_27290);
nand U27554 (N_27554,N_27284,N_27309);
or U27555 (N_27555,N_27288,N_27255);
and U27556 (N_27556,N_27258,N_27243);
xor U27557 (N_27557,N_27240,N_27333);
or U27558 (N_27558,N_27303,N_27367);
or U27559 (N_27559,N_27280,N_27298);
nor U27560 (N_27560,N_27366,N_27341);
nand U27561 (N_27561,N_27382,N_27300);
xor U27562 (N_27562,N_27317,N_27295);
nor U27563 (N_27563,N_27244,N_27393);
xor U27564 (N_27564,N_27224,N_27302);
xor U27565 (N_27565,N_27388,N_27234);
or U27566 (N_27566,N_27377,N_27366);
or U27567 (N_27567,N_27351,N_27256);
nor U27568 (N_27568,N_27303,N_27345);
xnor U27569 (N_27569,N_27225,N_27291);
nand U27570 (N_27570,N_27213,N_27291);
nor U27571 (N_27571,N_27389,N_27234);
and U27572 (N_27572,N_27208,N_27348);
and U27573 (N_27573,N_27379,N_27249);
xor U27574 (N_27574,N_27386,N_27364);
and U27575 (N_27575,N_27252,N_27365);
xor U27576 (N_27576,N_27212,N_27389);
nor U27577 (N_27577,N_27396,N_27255);
or U27578 (N_27578,N_27280,N_27320);
xor U27579 (N_27579,N_27355,N_27250);
or U27580 (N_27580,N_27290,N_27237);
nand U27581 (N_27581,N_27273,N_27377);
or U27582 (N_27582,N_27369,N_27371);
nand U27583 (N_27583,N_27340,N_27339);
nand U27584 (N_27584,N_27318,N_27381);
nor U27585 (N_27585,N_27305,N_27372);
or U27586 (N_27586,N_27391,N_27202);
or U27587 (N_27587,N_27280,N_27285);
and U27588 (N_27588,N_27200,N_27306);
nand U27589 (N_27589,N_27262,N_27362);
xor U27590 (N_27590,N_27298,N_27390);
xnor U27591 (N_27591,N_27390,N_27272);
nor U27592 (N_27592,N_27305,N_27366);
xnor U27593 (N_27593,N_27292,N_27371);
nand U27594 (N_27594,N_27279,N_27208);
nor U27595 (N_27595,N_27282,N_27245);
nor U27596 (N_27596,N_27225,N_27281);
and U27597 (N_27597,N_27349,N_27278);
or U27598 (N_27598,N_27340,N_27389);
or U27599 (N_27599,N_27293,N_27225);
nor U27600 (N_27600,N_27567,N_27455);
nand U27601 (N_27601,N_27500,N_27502);
nor U27602 (N_27602,N_27573,N_27411);
or U27603 (N_27603,N_27418,N_27590);
xor U27604 (N_27604,N_27592,N_27430);
nand U27605 (N_27605,N_27540,N_27516);
nor U27606 (N_27606,N_27484,N_27523);
or U27607 (N_27607,N_27426,N_27550);
nor U27608 (N_27608,N_27504,N_27447);
or U27609 (N_27609,N_27412,N_27553);
nand U27610 (N_27610,N_27469,N_27467);
xnor U27611 (N_27611,N_27531,N_27422);
xnor U27612 (N_27612,N_27485,N_27511);
nand U27613 (N_27613,N_27558,N_27457);
and U27614 (N_27614,N_27581,N_27555);
nor U27615 (N_27615,N_27423,N_27518);
or U27616 (N_27616,N_27463,N_27443);
nor U27617 (N_27617,N_27537,N_27591);
or U27618 (N_27618,N_27454,N_27416);
xnor U27619 (N_27619,N_27508,N_27559);
nor U27620 (N_27620,N_27509,N_27431);
or U27621 (N_27621,N_27476,N_27488);
nor U27622 (N_27622,N_27572,N_27528);
and U27623 (N_27623,N_27565,N_27519);
and U27624 (N_27624,N_27425,N_27486);
nor U27625 (N_27625,N_27522,N_27532);
and U27626 (N_27626,N_27541,N_27595);
and U27627 (N_27627,N_27507,N_27492);
or U27628 (N_27628,N_27474,N_27438);
xnor U27629 (N_27629,N_27433,N_27582);
or U27630 (N_27630,N_27599,N_27493);
nor U27631 (N_27631,N_27529,N_27446);
and U27632 (N_27632,N_27452,N_27549);
nor U27633 (N_27633,N_27598,N_27527);
and U27634 (N_27634,N_27501,N_27442);
or U27635 (N_27635,N_27556,N_27506);
nor U27636 (N_27636,N_27533,N_27561);
or U27637 (N_27637,N_27409,N_27427);
nor U27638 (N_27638,N_27417,N_27594);
and U27639 (N_27639,N_27499,N_27441);
or U27640 (N_27640,N_27473,N_27576);
xnor U27641 (N_27641,N_27419,N_27539);
and U27642 (N_27642,N_27520,N_27514);
nand U27643 (N_27643,N_27468,N_27543);
and U27644 (N_27644,N_27566,N_27597);
xor U27645 (N_27645,N_27453,N_27428);
and U27646 (N_27646,N_27421,N_27478);
nand U27647 (N_27647,N_27521,N_27524);
and U27648 (N_27648,N_27587,N_27577);
xnor U27649 (N_27649,N_27448,N_27563);
and U27650 (N_27650,N_27451,N_27585);
xnor U27651 (N_27651,N_27546,N_27415);
nand U27652 (N_27652,N_27481,N_27593);
and U27653 (N_27653,N_27407,N_27480);
nand U27654 (N_27654,N_27545,N_27471);
and U27655 (N_27655,N_27403,N_27487);
nor U27656 (N_27656,N_27510,N_27408);
xor U27657 (N_27657,N_27482,N_27475);
nor U27658 (N_27658,N_27580,N_27569);
and U27659 (N_27659,N_27477,N_27483);
nand U27660 (N_27660,N_27459,N_27432);
or U27661 (N_27661,N_27579,N_27445);
and U27662 (N_27662,N_27460,N_27542);
xor U27663 (N_27663,N_27536,N_27497);
or U27664 (N_27664,N_27495,N_27464);
or U27665 (N_27665,N_27535,N_27584);
or U27666 (N_27666,N_27401,N_27413);
nor U27667 (N_27667,N_27560,N_27513);
and U27668 (N_27668,N_27470,N_27517);
and U27669 (N_27669,N_27498,N_27583);
nand U27670 (N_27670,N_27458,N_27515);
nor U27671 (N_27671,N_27491,N_27414);
or U27672 (N_27672,N_27547,N_27494);
nor U27673 (N_27673,N_27406,N_27554);
nor U27674 (N_27674,N_27596,N_27404);
nand U27675 (N_27675,N_27400,N_27461);
or U27676 (N_27676,N_27424,N_27525);
nor U27677 (N_27677,N_27534,N_27465);
xnor U27678 (N_27678,N_27512,N_27405);
or U27679 (N_27679,N_27429,N_27439);
xor U27680 (N_27680,N_27496,N_27402);
nor U27681 (N_27681,N_27489,N_27440);
or U27682 (N_27682,N_27437,N_27548);
nand U27683 (N_27683,N_27434,N_27530);
nor U27684 (N_27684,N_27551,N_27589);
or U27685 (N_27685,N_27570,N_27436);
and U27686 (N_27686,N_27571,N_27450);
nor U27687 (N_27687,N_27526,N_27505);
nor U27688 (N_27688,N_27435,N_27538);
and U27689 (N_27689,N_27456,N_27410);
nand U27690 (N_27690,N_27466,N_27578);
or U27691 (N_27691,N_27472,N_27479);
nor U27692 (N_27692,N_27586,N_27462);
and U27693 (N_27693,N_27490,N_27574);
and U27694 (N_27694,N_27557,N_27552);
and U27695 (N_27695,N_27544,N_27588);
and U27696 (N_27696,N_27575,N_27503);
xor U27697 (N_27697,N_27444,N_27564);
xnor U27698 (N_27698,N_27562,N_27568);
and U27699 (N_27699,N_27420,N_27449);
nand U27700 (N_27700,N_27581,N_27469);
nand U27701 (N_27701,N_27415,N_27457);
and U27702 (N_27702,N_27457,N_27447);
xor U27703 (N_27703,N_27536,N_27422);
nor U27704 (N_27704,N_27462,N_27505);
xor U27705 (N_27705,N_27487,N_27451);
nor U27706 (N_27706,N_27585,N_27406);
xor U27707 (N_27707,N_27439,N_27573);
xor U27708 (N_27708,N_27481,N_27436);
xor U27709 (N_27709,N_27570,N_27480);
nor U27710 (N_27710,N_27431,N_27541);
and U27711 (N_27711,N_27578,N_27492);
xnor U27712 (N_27712,N_27546,N_27446);
or U27713 (N_27713,N_27578,N_27469);
nor U27714 (N_27714,N_27489,N_27576);
xnor U27715 (N_27715,N_27449,N_27555);
or U27716 (N_27716,N_27508,N_27512);
and U27717 (N_27717,N_27411,N_27439);
nand U27718 (N_27718,N_27566,N_27586);
nor U27719 (N_27719,N_27482,N_27438);
xnor U27720 (N_27720,N_27508,N_27537);
or U27721 (N_27721,N_27533,N_27558);
xor U27722 (N_27722,N_27472,N_27574);
or U27723 (N_27723,N_27431,N_27442);
or U27724 (N_27724,N_27422,N_27529);
xnor U27725 (N_27725,N_27586,N_27473);
nand U27726 (N_27726,N_27426,N_27487);
nand U27727 (N_27727,N_27485,N_27524);
nor U27728 (N_27728,N_27573,N_27431);
nor U27729 (N_27729,N_27465,N_27504);
nor U27730 (N_27730,N_27560,N_27501);
xor U27731 (N_27731,N_27597,N_27544);
or U27732 (N_27732,N_27422,N_27530);
nor U27733 (N_27733,N_27586,N_27477);
nand U27734 (N_27734,N_27458,N_27522);
nor U27735 (N_27735,N_27493,N_27547);
or U27736 (N_27736,N_27578,N_27427);
nand U27737 (N_27737,N_27503,N_27426);
nor U27738 (N_27738,N_27598,N_27566);
and U27739 (N_27739,N_27438,N_27541);
or U27740 (N_27740,N_27496,N_27565);
or U27741 (N_27741,N_27520,N_27480);
or U27742 (N_27742,N_27456,N_27575);
nand U27743 (N_27743,N_27527,N_27542);
or U27744 (N_27744,N_27484,N_27427);
xnor U27745 (N_27745,N_27464,N_27453);
and U27746 (N_27746,N_27558,N_27408);
and U27747 (N_27747,N_27530,N_27443);
and U27748 (N_27748,N_27510,N_27581);
and U27749 (N_27749,N_27535,N_27426);
xor U27750 (N_27750,N_27483,N_27552);
and U27751 (N_27751,N_27531,N_27485);
nand U27752 (N_27752,N_27492,N_27427);
or U27753 (N_27753,N_27488,N_27413);
nand U27754 (N_27754,N_27575,N_27490);
nor U27755 (N_27755,N_27479,N_27532);
nand U27756 (N_27756,N_27552,N_27412);
and U27757 (N_27757,N_27404,N_27565);
or U27758 (N_27758,N_27532,N_27456);
and U27759 (N_27759,N_27547,N_27469);
nor U27760 (N_27760,N_27546,N_27549);
or U27761 (N_27761,N_27423,N_27528);
and U27762 (N_27762,N_27589,N_27473);
nand U27763 (N_27763,N_27448,N_27510);
nor U27764 (N_27764,N_27499,N_27439);
xor U27765 (N_27765,N_27505,N_27417);
nor U27766 (N_27766,N_27473,N_27475);
nand U27767 (N_27767,N_27476,N_27559);
xor U27768 (N_27768,N_27482,N_27462);
xor U27769 (N_27769,N_27587,N_27406);
nand U27770 (N_27770,N_27592,N_27549);
xnor U27771 (N_27771,N_27445,N_27551);
or U27772 (N_27772,N_27419,N_27446);
and U27773 (N_27773,N_27557,N_27591);
and U27774 (N_27774,N_27572,N_27582);
or U27775 (N_27775,N_27555,N_27431);
and U27776 (N_27776,N_27492,N_27482);
nand U27777 (N_27777,N_27509,N_27410);
nor U27778 (N_27778,N_27453,N_27546);
nand U27779 (N_27779,N_27563,N_27406);
xor U27780 (N_27780,N_27522,N_27548);
nand U27781 (N_27781,N_27571,N_27520);
nand U27782 (N_27782,N_27529,N_27427);
nand U27783 (N_27783,N_27594,N_27447);
xnor U27784 (N_27784,N_27437,N_27435);
or U27785 (N_27785,N_27509,N_27444);
or U27786 (N_27786,N_27589,N_27599);
xor U27787 (N_27787,N_27592,N_27515);
or U27788 (N_27788,N_27439,N_27408);
nor U27789 (N_27789,N_27405,N_27431);
or U27790 (N_27790,N_27461,N_27525);
and U27791 (N_27791,N_27542,N_27557);
or U27792 (N_27792,N_27496,N_27436);
or U27793 (N_27793,N_27580,N_27502);
or U27794 (N_27794,N_27444,N_27485);
or U27795 (N_27795,N_27435,N_27490);
and U27796 (N_27796,N_27455,N_27427);
or U27797 (N_27797,N_27411,N_27559);
nor U27798 (N_27798,N_27582,N_27550);
and U27799 (N_27799,N_27507,N_27411);
xnor U27800 (N_27800,N_27741,N_27659);
nor U27801 (N_27801,N_27699,N_27765);
xor U27802 (N_27802,N_27678,N_27616);
xnor U27803 (N_27803,N_27649,N_27688);
xnor U27804 (N_27804,N_27748,N_27762);
and U27805 (N_27805,N_27786,N_27719);
and U27806 (N_27806,N_27754,N_27770);
nor U27807 (N_27807,N_27687,N_27607);
xor U27808 (N_27808,N_27734,N_27796);
nand U27809 (N_27809,N_27689,N_27705);
or U27810 (N_27810,N_27655,N_27698);
or U27811 (N_27811,N_27738,N_27769);
nor U27812 (N_27812,N_27675,N_27685);
or U27813 (N_27813,N_27600,N_27642);
nor U27814 (N_27814,N_27610,N_27761);
nand U27815 (N_27815,N_27608,N_27601);
and U27816 (N_27816,N_27668,N_27701);
or U27817 (N_27817,N_27626,N_27684);
or U27818 (N_27818,N_27782,N_27708);
or U27819 (N_27819,N_27788,N_27760);
or U27820 (N_27820,N_27612,N_27713);
xor U27821 (N_27821,N_27722,N_27679);
or U27822 (N_27822,N_27707,N_27714);
or U27823 (N_27823,N_27620,N_27625);
nor U27824 (N_27824,N_27619,N_27650);
xor U27825 (N_27825,N_27697,N_27645);
nand U27826 (N_27826,N_27749,N_27778);
nand U27827 (N_27827,N_27797,N_27773);
nor U27828 (N_27828,N_27696,N_27723);
and U27829 (N_27829,N_27753,N_27634);
and U27830 (N_27830,N_27794,N_27643);
or U27831 (N_27831,N_27781,N_27720);
and U27832 (N_27832,N_27690,N_27744);
nand U27833 (N_27833,N_27758,N_27768);
or U27834 (N_27834,N_27694,N_27751);
or U27835 (N_27835,N_27793,N_27680);
and U27836 (N_27836,N_27629,N_27672);
nand U27837 (N_27837,N_27644,N_27767);
and U27838 (N_27838,N_27779,N_27771);
nor U27839 (N_27839,N_27654,N_27683);
and U27840 (N_27840,N_27739,N_27665);
and U27841 (N_27841,N_27799,N_27666);
xnor U27842 (N_27842,N_27740,N_27732);
nor U27843 (N_27843,N_27658,N_27641);
and U27844 (N_27844,N_27712,N_27736);
xor U27845 (N_27845,N_27671,N_27693);
nor U27846 (N_27846,N_27648,N_27664);
nor U27847 (N_27847,N_27727,N_27766);
and U27848 (N_27848,N_27710,N_27783);
and U27849 (N_27849,N_27622,N_27759);
nand U27850 (N_27850,N_27700,N_27681);
nand U27851 (N_27851,N_27624,N_27611);
nand U27852 (N_27852,N_27728,N_27764);
and U27853 (N_27853,N_27798,N_27795);
and U27854 (N_27854,N_27730,N_27669);
nand U27855 (N_27855,N_27657,N_27718);
xnor U27856 (N_27856,N_27731,N_27628);
xnor U27857 (N_27857,N_27606,N_27691);
and U27858 (N_27858,N_27784,N_27603);
xnor U27859 (N_27859,N_27682,N_27735);
xor U27860 (N_27860,N_27776,N_27677);
or U27861 (N_27861,N_27711,N_27737);
nand U27862 (N_27862,N_27617,N_27633);
xor U27863 (N_27863,N_27777,N_27717);
nor U27864 (N_27864,N_27638,N_27792);
nor U27865 (N_27865,N_27618,N_27651);
nor U27866 (N_27866,N_27652,N_27686);
and U27867 (N_27867,N_27615,N_27757);
or U27868 (N_27868,N_27673,N_27660);
nand U27869 (N_27869,N_27695,N_27621);
xor U27870 (N_27870,N_27656,N_27750);
or U27871 (N_27871,N_27789,N_27637);
and U27872 (N_27872,N_27646,N_27787);
and U27873 (N_27873,N_27623,N_27632);
nand U27874 (N_27874,N_27670,N_27791);
xor U27875 (N_27875,N_27640,N_27692);
nor U27876 (N_27876,N_27630,N_27733);
or U27877 (N_27877,N_27613,N_27663);
and U27878 (N_27878,N_27790,N_27631);
and U27879 (N_27879,N_27676,N_27756);
and U27880 (N_27880,N_27775,N_27674);
nand U27881 (N_27881,N_27725,N_27627);
or U27882 (N_27882,N_27667,N_27780);
or U27883 (N_27883,N_27772,N_27774);
nor U27884 (N_27884,N_27716,N_27635);
nor U27885 (N_27885,N_27752,N_27742);
xnor U27886 (N_27886,N_27721,N_27661);
and U27887 (N_27887,N_27746,N_27745);
nor U27888 (N_27888,N_27703,N_27614);
xor U27889 (N_27889,N_27763,N_27604);
nor U27890 (N_27890,N_27639,N_27647);
nor U27891 (N_27891,N_27702,N_27706);
nand U27892 (N_27892,N_27709,N_27729);
nand U27893 (N_27893,N_27747,N_27609);
and U27894 (N_27894,N_27662,N_27605);
or U27895 (N_27895,N_27785,N_27755);
or U27896 (N_27896,N_27726,N_27704);
and U27897 (N_27897,N_27715,N_27636);
nor U27898 (N_27898,N_27653,N_27724);
nand U27899 (N_27899,N_27743,N_27602);
and U27900 (N_27900,N_27707,N_27612);
nor U27901 (N_27901,N_27735,N_27789);
or U27902 (N_27902,N_27737,N_27644);
and U27903 (N_27903,N_27626,N_27782);
and U27904 (N_27904,N_27672,N_27709);
xor U27905 (N_27905,N_27601,N_27688);
nor U27906 (N_27906,N_27737,N_27604);
xor U27907 (N_27907,N_27601,N_27674);
nor U27908 (N_27908,N_27678,N_27635);
xnor U27909 (N_27909,N_27707,N_27796);
nor U27910 (N_27910,N_27761,N_27652);
nor U27911 (N_27911,N_27760,N_27699);
xor U27912 (N_27912,N_27751,N_27614);
or U27913 (N_27913,N_27665,N_27697);
and U27914 (N_27914,N_27728,N_27676);
nor U27915 (N_27915,N_27629,N_27794);
nand U27916 (N_27916,N_27794,N_27604);
nand U27917 (N_27917,N_27791,N_27689);
or U27918 (N_27918,N_27648,N_27768);
xor U27919 (N_27919,N_27763,N_27635);
nor U27920 (N_27920,N_27611,N_27795);
and U27921 (N_27921,N_27610,N_27771);
nand U27922 (N_27922,N_27773,N_27609);
nand U27923 (N_27923,N_27656,N_27758);
nor U27924 (N_27924,N_27623,N_27784);
nand U27925 (N_27925,N_27629,N_27760);
xor U27926 (N_27926,N_27661,N_27728);
xor U27927 (N_27927,N_27706,N_27602);
nor U27928 (N_27928,N_27709,N_27750);
nor U27929 (N_27929,N_27793,N_27722);
or U27930 (N_27930,N_27778,N_27753);
or U27931 (N_27931,N_27696,N_27642);
and U27932 (N_27932,N_27614,N_27760);
or U27933 (N_27933,N_27641,N_27617);
nand U27934 (N_27934,N_27789,N_27762);
xnor U27935 (N_27935,N_27685,N_27784);
xnor U27936 (N_27936,N_27740,N_27650);
nand U27937 (N_27937,N_27631,N_27752);
nand U27938 (N_27938,N_27711,N_27636);
nor U27939 (N_27939,N_27751,N_27662);
and U27940 (N_27940,N_27790,N_27721);
nor U27941 (N_27941,N_27636,N_27654);
nor U27942 (N_27942,N_27714,N_27794);
or U27943 (N_27943,N_27777,N_27677);
xnor U27944 (N_27944,N_27736,N_27628);
and U27945 (N_27945,N_27624,N_27660);
nor U27946 (N_27946,N_27646,N_27732);
nor U27947 (N_27947,N_27742,N_27772);
nand U27948 (N_27948,N_27663,N_27693);
nor U27949 (N_27949,N_27707,N_27709);
and U27950 (N_27950,N_27736,N_27734);
xor U27951 (N_27951,N_27688,N_27617);
nor U27952 (N_27952,N_27759,N_27678);
nor U27953 (N_27953,N_27714,N_27655);
nand U27954 (N_27954,N_27658,N_27765);
and U27955 (N_27955,N_27652,N_27619);
xnor U27956 (N_27956,N_27658,N_27771);
nor U27957 (N_27957,N_27704,N_27780);
nand U27958 (N_27958,N_27726,N_27610);
or U27959 (N_27959,N_27609,N_27642);
nand U27960 (N_27960,N_27765,N_27637);
or U27961 (N_27961,N_27751,N_27654);
xor U27962 (N_27962,N_27686,N_27691);
and U27963 (N_27963,N_27727,N_27763);
xnor U27964 (N_27964,N_27798,N_27698);
or U27965 (N_27965,N_27669,N_27744);
nor U27966 (N_27966,N_27620,N_27729);
or U27967 (N_27967,N_27779,N_27742);
nand U27968 (N_27968,N_27765,N_27639);
xnor U27969 (N_27969,N_27703,N_27784);
or U27970 (N_27970,N_27686,N_27626);
xor U27971 (N_27971,N_27778,N_27642);
nor U27972 (N_27972,N_27709,N_27702);
and U27973 (N_27973,N_27703,N_27742);
or U27974 (N_27974,N_27751,N_27691);
xnor U27975 (N_27975,N_27647,N_27721);
nor U27976 (N_27976,N_27784,N_27622);
or U27977 (N_27977,N_27717,N_27631);
and U27978 (N_27978,N_27623,N_27673);
nand U27979 (N_27979,N_27661,N_27621);
nand U27980 (N_27980,N_27754,N_27776);
or U27981 (N_27981,N_27774,N_27612);
nor U27982 (N_27982,N_27798,N_27664);
xnor U27983 (N_27983,N_27761,N_27632);
nor U27984 (N_27984,N_27747,N_27618);
nand U27985 (N_27985,N_27769,N_27675);
xor U27986 (N_27986,N_27629,N_27757);
and U27987 (N_27987,N_27683,N_27618);
and U27988 (N_27988,N_27758,N_27769);
and U27989 (N_27989,N_27637,N_27739);
nand U27990 (N_27990,N_27731,N_27730);
xor U27991 (N_27991,N_27778,N_27760);
nand U27992 (N_27992,N_27684,N_27672);
and U27993 (N_27993,N_27700,N_27787);
nor U27994 (N_27994,N_27629,N_27714);
nand U27995 (N_27995,N_27794,N_27614);
or U27996 (N_27996,N_27763,N_27790);
and U27997 (N_27997,N_27773,N_27619);
xor U27998 (N_27998,N_27695,N_27763);
nor U27999 (N_27999,N_27798,N_27644);
nand U28000 (N_28000,N_27814,N_27816);
and U28001 (N_28001,N_27981,N_27969);
xor U28002 (N_28002,N_27920,N_27892);
xnor U28003 (N_28003,N_27871,N_27877);
nor U28004 (N_28004,N_27849,N_27974);
nor U28005 (N_28005,N_27885,N_27954);
and U28006 (N_28006,N_27917,N_27983);
and U28007 (N_28007,N_27838,N_27870);
nand U28008 (N_28008,N_27991,N_27821);
or U28009 (N_28009,N_27873,N_27956);
and U28010 (N_28010,N_27947,N_27908);
nor U28011 (N_28011,N_27957,N_27979);
nand U28012 (N_28012,N_27907,N_27913);
or U28013 (N_28013,N_27990,N_27976);
and U28014 (N_28014,N_27832,N_27972);
or U28015 (N_28015,N_27881,N_27841);
and U28016 (N_28016,N_27867,N_27930);
xor U28017 (N_28017,N_27928,N_27804);
nand U28018 (N_28018,N_27802,N_27915);
nor U28019 (N_28019,N_27936,N_27940);
or U28020 (N_28020,N_27805,N_27800);
or U28021 (N_28021,N_27888,N_27831);
and U28022 (N_28022,N_27883,N_27842);
nor U28023 (N_28023,N_27891,N_27989);
and U28024 (N_28024,N_27852,N_27894);
xnor U28025 (N_28025,N_27929,N_27955);
or U28026 (N_28026,N_27809,N_27828);
or U28027 (N_28027,N_27997,N_27878);
and U28028 (N_28028,N_27911,N_27824);
nor U28029 (N_28029,N_27925,N_27910);
or U28030 (N_28030,N_27810,N_27906);
xor U28031 (N_28031,N_27876,N_27951);
nand U28032 (N_28032,N_27855,N_27909);
and U28033 (N_28033,N_27840,N_27811);
xnor U28034 (N_28034,N_27865,N_27825);
nor U28035 (N_28035,N_27939,N_27985);
nor U28036 (N_28036,N_27986,N_27851);
or U28037 (N_28037,N_27836,N_27900);
nor U28038 (N_28038,N_27998,N_27950);
nand U28039 (N_28039,N_27975,N_27833);
or U28040 (N_28040,N_27971,N_27826);
or U28041 (N_28041,N_27854,N_27932);
and U28042 (N_28042,N_27837,N_27890);
nand U28043 (N_28043,N_27801,N_27984);
nor U28044 (N_28044,N_27903,N_27964);
xor U28045 (N_28045,N_27944,N_27866);
and U28046 (N_28046,N_27819,N_27970);
nor U28047 (N_28047,N_27818,N_27962);
and U28048 (N_28048,N_27921,N_27963);
nand U28049 (N_28049,N_27961,N_27923);
xor U28050 (N_28050,N_27834,N_27848);
xnor U28051 (N_28051,N_27864,N_27914);
nand U28052 (N_28052,N_27872,N_27935);
xor U28053 (N_28053,N_27806,N_27982);
and U28054 (N_28054,N_27808,N_27999);
nand U28055 (N_28055,N_27978,N_27996);
nor U28056 (N_28056,N_27843,N_27893);
or U28057 (N_28057,N_27958,N_27992);
nor U28058 (N_28058,N_27846,N_27904);
xnor U28059 (N_28059,N_27880,N_27959);
nor U28060 (N_28060,N_27980,N_27902);
and U28061 (N_28061,N_27835,N_27862);
xor U28062 (N_28062,N_27977,N_27889);
xor U28063 (N_28063,N_27931,N_27820);
and U28064 (N_28064,N_27937,N_27847);
nand U28065 (N_28065,N_27812,N_27945);
xor U28066 (N_28066,N_27987,N_27941);
xor U28067 (N_28067,N_27857,N_27919);
xor U28068 (N_28068,N_27844,N_27829);
and U28069 (N_28069,N_27813,N_27868);
nand U28070 (N_28070,N_27922,N_27927);
xnor U28071 (N_28071,N_27817,N_27898);
nor U28072 (N_28072,N_27901,N_27918);
and U28073 (N_28073,N_27861,N_27887);
or U28074 (N_28074,N_27839,N_27994);
or U28075 (N_28075,N_27973,N_27905);
xnor U28076 (N_28076,N_27899,N_27875);
and U28077 (N_28077,N_27860,N_27938);
nor U28078 (N_28078,N_27933,N_27807);
nor U28079 (N_28079,N_27993,N_27858);
and U28080 (N_28080,N_27966,N_27897);
xor U28081 (N_28081,N_27845,N_27988);
nand U28082 (N_28082,N_27823,N_27853);
or U28083 (N_28083,N_27896,N_27953);
nand U28084 (N_28084,N_27912,N_27859);
or U28085 (N_28085,N_27916,N_27943);
and U28086 (N_28086,N_27960,N_27949);
nand U28087 (N_28087,N_27924,N_27803);
nor U28088 (N_28088,N_27827,N_27830);
nand U28089 (N_28089,N_27869,N_27879);
xor U28090 (N_28090,N_27948,N_27822);
and U28091 (N_28091,N_27968,N_27946);
and U28092 (N_28092,N_27995,N_27942);
or U28093 (N_28093,N_27882,N_27874);
nand U28094 (N_28094,N_27967,N_27884);
and U28095 (N_28095,N_27952,N_27926);
or U28096 (N_28096,N_27856,N_27850);
xnor U28097 (N_28097,N_27863,N_27965);
nand U28098 (N_28098,N_27815,N_27895);
or U28099 (N_28099,N_27934,N_27886);
nand U28100 (N_28100,N_27814,N_27993);
or U28101 (N_28101,N_27867,N_27982);
nand U28102 (N_28102,N_27814,N_27824);
xnor U28103 (N_28103,N_27975,N_27876);
and U28104 (N_28104,N_27860,N_27858);
or U28105 (N_28105,N_27925,N_27955);
xnor U28106 (N_28106,N_27937,N_27969);
xor U28107 (N_28107,N_27955,N_27918);
nand U28108 (N_28108,N_27882,N_27986);
xnor U28109 (N_28109,N_27996,N_27886);
nand U28110 (N_28110,N_27999,N_27950);
and U28111 (N_28111,N_27983,N_27814);
nand U28112 (N_28112,N_27900,N_27928);
nand U28113 (N_28113,N_27931,N_27949);
xor U28114 (N_28114,N_27935,N_27878);
nand U28115 (N_28115,N_27868,N_27833);
and U28116 (N_28116,N_27943,N_27996);
nand U28117 (N_28117,N_27935,N_27819);
nand U28118 (N_28118,N_27884,N_27993);
nor U28119 (N_28119,N_27911,N_27896);
nor U28120 (N_28120,N_27846,N_27872);
and U28121 (N_28121,N_27869,N_27976);
or U28122 (N_28122,N_27812,N_27846);
nor U28123 (N_28123,N_27844,N_27800);
nand U28124 (N_28124,N_27883,N_27964);
or U28125 (N_28125,N_27964,N_27845);
or U28126 (N_28126,N_27969,N_27940);
xor U28127 (N_28127,N_27909,N_27913);
xnor U28128 (N_28128,N_27897,N_27928);
and U28129 (N_28129,N_27926,N_27982);
xor U28130 (N_28130,N_27978,N_27954);
and U28131 (N_28131,N_27927,N_27914);
and U28132 (N_28132,N_27886,N_27878);
and U28133 (N_28133,N_27998,N_27940);
nor U28134 (N_28134,N_27846,N_27980);
nand U28135 (N_28135,N_27929,N_27835);
nand U28136 (N_28136,N_27936,N_27865);
xor U28137 (N_28137,N_27914,N_27930);
xnor U28138 (N_28138,N_27845,N_27941);
nand U28139 (N_28139,N_27872,N_27946);
nor U28140 (N_28140,N_27883,N_27860);
xor U28141 (N_28141,N_27971,N_27913);
or U28142 (N_28142,N_27887,N_27951);
or U28143 (N_28143,N_27914,N_27978);
xor U28144 (N_28144,N_27830,N_27951);
nand U28145 (N_28145,N_27856,N_27955);
xor U28146 (N_28146,N_27980,N_27972);
nor U28147 (N_28147,N_27858,N_27922);
or U28148 (N_28148,N_27977,N_27983);
nand U28149 (N_28149,N_27920,N_27933);
or U28150 (N_28150,N_27859,N_27848);
nand U28151 (N_28151,N_27826,N_27806);
nor U28152 (N_28152,N_27819,N_27802);
nand U28153 (N_28153,N_27899,N_27918);
or U28154 (N_28154,N_27856,N_27917);
nor U28155 (N_28155,N_27976,N_27993);
xnor U28156 (N_28156,N_27834,N_27947);
and U28157 (N_28157,N_27800,N_27920);
or U28158 (N_28158,N_27842,N_27847);
or U28159 (N_28159,N_27816,N_27835);
nand U28160 (N_28160,N_27951,N_27938);
and U28161 (N_28161,N_27835,N_27916);
and U28162 (N_28162,N_27807,N_27895);
nor U28163 (N_28163,N_27923,N_27942);
or U28164 (N_28164,N_27903,N_27884);
nor U28165 (N_28165,N_27938,N_27864);
nand U28166 (N_28166,N_27895,N_27967);
nor U28167 (N_28167,N_27941,N_27817);
and U28168 (N_28168,N_27910,N_27847);
nor U28169 (N_28169,N_27864,N_27892);
nand U28170 (N_28170,N_27913,N_27834);
and U28171 (N_28171,N_27964,N_27834);
or U28172 (N_28172,N_27846,N_27924);
nand U28173 (N_28173,N_27810,N_27915);
nand U28174 (N_28174,N_27999,N_27929);
nor U28175 (N_28175,N_27909,N_27976);
xor U28176 (N_28176,N_27825,N_27896);
and U28177 (N_28177,N_27871,N_27836);
nand U28178 (N_28178,N_27955,N_27902);
xnor U28179 (N_28179,N_27965,N_27959);
or U28180 (N_28180,N_27835,N_27868);
or U28181 (N_28181,N_27960,N_27866);
and U28182 (N_28182,N_27813,N_27959);
nor U28183 (N_28183,N_27968,N_27828);
nor U28184 (N_28184,N_27842,N_27990);
xnor U28185 (N_28185,N_27919,N_27943);
and U28186 (N_28186,N_27929,N_27800);
xor U28187 (N_28187,N_27902,N_27969);
nand U28188 (N_28188,N_27907,N_27945);
nor U28189 (N_28189,N_27912,N_27842);
xnor U28190 (N_28190,N_27828,N_27948);
or U28191 (N_28191,N_27857,N_27804);
and U28192 (N_28192,N_27914,N_27951);
and U28193 (N_28193,N_27908,N_27845);
xnor U28194 (N_28194,N_27889,N_27896);
nand U28195 (N_28195,N_27860,N_27863);
nand U28196 (N_28196,N_27979,N_27924);
and U28197 (N_28197,N_27937,N_27849);
or U28198 (N_28198,N_27856,N_27832);
xor U28199 (N_28199,N_27854,N_27911);
nor U28200 (N_28200,N_28137,N_28042);
and U28201 (N_28201,N_28005,N_28100);
or U28202 (N_28202,N_28165,N_28022);
and U28203 (N_28203,N_28103,N_28036);
nand U28204 (N_28204,N_28021,N_28027);
xnor U28205 (N_28205,N_28032,N_28112);
nor U28206 (N_28206,N_28195,N_28080);
nand U28207 (N_28207,N_28006,N_28128);
xnor U28208 (N_28208,N_28064,N_28188);
xor U28209 (N_28209,N_28016,N_28065);
nor U28210 (N_28210,N_28074,N_28040);
nor U28211 (N_28211,N_28157,N_28122);
and U28212 (N_28212,N_28182,N_28124);
xor U28213 (N_28213,N_28172,N_28133);
xnor U28214 (N_28214,N_28190,N_28175);
and U28215 (N_28215,N_28098,N_28177);
nand U28216 (N_28216,N_28046,N_28097);
xor U28217 (N_28217,N_28012,N_28115);
xnor U28218 (N_28218,N_28028,N_28158);
nor U28219 (N_28219,N_28143,N_28018);
and U28220 (N_28220,N_28029,N_28164);
nand U28221 (N_28221,N_28031,N_28118);
and U28222 (N_28222,N_28166,N_28070);
nand U28223 (N_28223,N_28107,N_28192);
and U28224 (N_28224,N_28058,N_28108);
nor U28225 (N_28225,N_28049,N_28059);
xnor U28226 (N_28226,N_28136,N_28000);
nor U28227 (N_28227,N_28198,N_28011);
nand U28228 (N_28228,N_28078,N_28130);
xnor U28229 (N_28229,N_28194,N_28057);
nor U28230 (N_28230,N_28077,N_28176);
xor U28231 (N_28231,N_28147,N_28092);
nor U28232 (N_28232,N_28174,N_28020);
nand U28233 (N_28233,N_28045,N_28185);
xnor U28234 (N_28234,N_28087,N_28061);
nand U28235 (N_28235,N_28019,N_28180);
nor U28236 (N_28236,N_28110,N_28134);
nor U28237 (N_28237,N_28041,N_28150);
nor U28238 (N_28238,N_28141,N_28106);
and U28239 (N_28239,N_28086,N_28037);
nor U28240 (N_28240,N_28125,N_28144);
xnor U28241 (N_28241,N_28052,N_28063);
nor U28242 (N_28242,N_28024,N_28127);
nor U28243 (N_28243,N_28187,N_28056);
nand U28244 (N_28244,N_28048,N_28197);
or U28245 (N_28245,N_28113,N_28169);
nand U28246 (N_28246,N_28116,N_28093);
and U28247 (N_28247,N_28178,N_28142);
and U28248 (N_28248,N_28009,N_28154);
nand U28249 (N_28249,N_28160,N_28094);
xor U28250 (N_28250,N_28167,N_28162);
and U28251 (N_28251,N_28196,N_28026);
xor U28252 (N_28252,N_28114,N_28193);
nand U28253 (N_28253,N_28084,N_28034);
or U28254 (N_28254,N_28007,N_28129);
and U28255 (N_28255,N_28126,N_28123);
or U28256 (N_28256,N_28138,N_28173);
or U28257 (N_28257,N_28153,N_28109);
nor U28258 (N_28258,N_28035,N_28139);
nor U28259 (N_28259,N_28067,N_28102);
nor U28260 (N_28260,N_28183,N_28184);
nor U28261 (N_28261,N_28071,N_28003);
nand U28262 (N_28262,N_28117,N_28179);
xor U28263 (N_28263,N_28051,N_28072);
and U28264 (N_28264,N_28025,N_28199);
xnor U28265 (N_28265,N_28145,N_28146);
xor U28266 (N_28266,N_28053,N_28002);
nand U28267 (N_28267,N_28168,N_28076);
xor U28268 (N_28268,N_28105,N_28159);
and U28269 (N_28269,N_28068,N_28140);
and U28270 (N_28270,N_28161,N_28008);
xnor U28271 (N_28271,N_28014,N_28131);
nand U28272 (N_28272,N_28151,N_28060);
nor U28273 (N_28273,N_28135,N_28069);
nor U28274 (N_28274,N_28132,N_28081);
xor U28275 (N_28275,N_28083,N_28050);
xor U28276 (N_28276,N_28010,N_28099);
or U28277 (N_28277,N_28030,N_28170);
xor U28278 (N_28278,N_28189,N_28149);
nor U28279 (N_28279,N_28039,N_28090);
nand U28280 (N_28280,N_28004,N_28075);
or U28281 (N_28281,N_28054,N_28186);
nor U28282 (N_28282,N_28101,N_28038);
nand U28283 (N_28283,N_28095,N_28148);
and U28284 (N_28284,N_28088,N_28073);
nand U28285 (N_28285,N_28047,N_28163);
and U28286 (N_28286,N_28017,N_28062);
nor U28287 (N_28287,N_28066,N_28091);
nand U28288 (N_28288,N_28120,N_28171);
nor U28289 (N_28289,N_28013,N_28152);
or U28290 (N_28290,N_28191,N_28096);
and U28291 (N_28291,N_28121,N_28033);
and U28292 (N_28292,N_28156,N_28015);
nor U28293 (N_28293,N_28089,N_28111);
xor U28294 (N_28294,N_28119,N_28079);
nand U28295 (N_28295,N_28055,N_28023);
and U28296 (N_28296,N_28082,N_28043);
nor U28297 (N_28297,N_28104,N_28155);
xor U28298 (N_28298,N_28181,N_28001);
nor U28299 (N_28299,N_28085,N_28044);
or U28300 (N_28300,N_28196,N_28091);
xnor U28301 (N_28301,N_28006,N_28096);
nor U28302 (N_28302,N_28113,N_28127);
nor U28303 (N_28303,N_28177,N_28143);
and U28304 (N_28304,N_28072,N_28062);
nor U28305 (N_28305,N_28109,N_28154);
nand U28306 (N_28306,N_28111,N_28076);
nor U28307 (N_28307,N_28134,N_28181);
or U28308 (N_28308,N_28102,N_28100);
or U28309 (N_28309,N_28185,N_28150);
xnor U28310 (N_28310,N_28081,N_28048);
and U28311 (N_28311,N_28083,N_28199);
or U28312 (N_28312,N_28101,N_28143);
nor U28313 (N_28313,N_28108,N_28024);
xnor U28314 (N_28314,N_28030,N_28083);
nand U28315 (N_28315,N_28030,N_28189);
xnor U28316 (N_28316,N_28119,N_28142);
xnor U28317 (N_28317,N_28198,N_28185);
or U28318 (N_28318,N_28151,N_28016);
nand U28319 (N_28319,N_28023,N_28173);
xnor U28320 (N_28320,N_28191,N_28161);
xor U28321 (N_28321,N_28098,N_28029);
xor U28322 (N_28322,N_28052,N_28185);
xor U28323 (N_28323,N_28056,N_28042);
or U28324 (N_28324,N_28136,N_28100);
and U28325 (N_28325,N_28034,N_28059);
nor U28326 (N_28326,N_28183,N_28174);
nor U28327 (N_28327,N_28129,N_28193);
and U28328 (N_28328,N_28102,N_28154);
or U28329 (N_28329,N_28190,N_28082);
and U28330 (N_28330,N_28139,N_28104);
xor U28331 (N_28331,N_28118,N_28173);
xor U28332 (N_28332,N_28093,N_28135);
nand U28333 (N_28333,N_28106,N_28167);
and U28334 (N_28334,N_28031,N_28192);
xnor U28335 (N_28335,N_28088,N_28173);
nor U28336 (N_28336,N_28087,N_28142);
and U28337 (N_28337,N_28032,N_28189);
nor U28338 (N_28338,N_28003,N_28007);
nor U28339 (N_28339,N_28111,N_28197);
and U28340 (N_28340,N_28194,N_28036);
xnor U28341 (N_28341,N_28134,N_28096);
nor U28342 (N_28342,N_28079,N_28098);
xnor U28343 (N_28343,N_28106,N_28003);
nor U28344 (N_28344,N_28152,N_28080);
xor U28345 (N_28345,N_28033,N_28124);
nor U28346 (N_28346,N_28016,N_28024);
xnor U28347 (N_28347,N_28003,N_28197);
xor U28348 (N_28348,N_28034,N_28014);
and U28349 (N_28349,N_28186,N_28135);
or U28350 (N_28350,N_28058,N_28148);
xor U28351 (N_28351,N_28129,N_28188);
nor U28352 (N_28352,N_28195,N_28151);
nand U28353 (N_28353,N_28170,N_28147);
or U28354 (N_28354,N_28100,N_28093);
nor U28355 (N_28355,N_28153,N_28118);
nor U28356 (N_28356,N_28000,N_28025);
nor U28357 (N_28357,N_28047,N_28196);
or U28358 (N_28358,N_28136,N_28184);
nor U28359 (N_28359,N_28142,N_28064);
xnor U28360 (N_28360,N_28061,N_28010);
nand U28361 (N_28361,N_28020,N_28054);
nor U28362 (N_28362,N_28079,N_28108);
nor U28363 (N_28363,N_28190,N_28171);
and U28364 (N_28364,N_28006,N_28097);
or U28365 (N_28365,N_28183,N_28145);
or U28366 (N_28366,N_28062,N_28198);
xnor U28367 (N_28367,N_28042,N_28169);
or U28368 (N_28368,N_28056,N_28154);
nor U28369 (N_28369,N_28152,N_28025);
nor U28370 (N_28370,N_28162,N_28154);
xnor U28371 (N_28371,N_28142,N_28095);
xnor U28372 (N_28372,N_28108,N_28155);
and U28373 (N_28373,N_28103,N_28102);
xor U28374 (N_28374,N_28018,N_28129);
xor U28375 (N_28375,N_28074,N_28002);
nor U28376 (N_28376,N_28119,N_28108);
nor U28377 (N_28377,N_28199,N_28096);
xnor U28378 (N_28378,N_28119,N_28048);
or U28379 (N_28379,N_28007,N_28036);
nand U28380 (N_28380,N_28077,N_28150);
xnor U28381 (N_28381,N_28125,N_28074);
nand U28382 (N_28382,N_28067,N_28145);
xnor U28383 (N_28383,N_28096,N_28018);
or U28384 (N_28384,N_28071,N_28149);
xnor U28385 (N_28385,N_28021,N_28071);
and U28386 (N_28386,N_28183,N_28080);
or U28387 (N_28387,N_28082,N_28008);
and U28388 (N_28388,N_28113,N_28034);
xor U28389 (N_28389,N_28104,N_28092);
nor U28390 (N_28390,N_28190,N_28113);
nand U28391 (N_28391,N_28193,N_28157);
and U28392 (N_28392,N_28043,N_28048);
nand U28393 (N_28393,N_28093,N_28101);
nor U28394 (N_28394,N_28126,N_28150);
or U28395 (N_28395,N_28170,N_28004);
nand U28396 (N_28396,N_28099,N_28031);
xnor U28397 (N_28397,N_28142,N_28177);
and U28398 (N_28398,N_28085,N_28042);
nand U28399 (N_28399,N_28021,N_28123);
nand U28400 (N_28400,N_28208,N_28218);
and U28401 (N_28401,N_28320,N_28382);
and U28402 (N_28402,N_28252,N_28302);
or U28403 (N_28403,N_28286,N_28383);
nand U28404 (N_28404,N_28344,N_28305);
nor U28405 (N_28405,N_28367,N_28328);
and U28406 (N_28406,N_28349,N_28378);
xnor U28407 (N_28407,N_28225,N_28317);
nor U28408 (N_28408,N_28211,N_28290);
nand U28409 (N_28409,N_28205,N_28299);
or U28410 (N_28410,N_28303,N_28337);
nor U28411 (N_28411,N_28363,N_28352);
xnor U28412 (N_28412,N_28316,N_28330);
xnor U28413 (N_28413,N_28321,N_28256);
xor U28414 (N_28414,N_28276,N_28325);
nor U28415 (N_28415,N_28206,N_28280);
xnor U28416 (N_28416,N_28377,N_28322);
nand U28417 (N_28417,N_28358,N_28255);
and U28418 (N_28418,N_28222,N_28233);
nand U28419 (N_28419,N_28306,N_28271);
nand U28420 (N_28420,N_28294,N_28257);
xnor U28421 (N_28421,N_28370,N_28212);
or U28422 (N_28422,N_28369,N_28304);
and U28423 (N_28423,N_28270,N_28292);
and U28424 (N_28424,N_28339,N_28341);
nand U28425 (N_28425,N_28266,N_28334);
xnor U28426 (N_28426,N_28376,N_28249);
or U28427 (N_28427,N_28393,N_28269);
nand U28428 (N_28428,N_28210,N_28283);
or U28429 (N_28429,N_28373,N_28391);
nand U28430 (N_28430,N_28204,N_28336);
nor U28431 (N_28431,N_28372,N_28386);
or U28432 (N_28432,N_28223,N_28265);
nor U28433 (N_28433,N_28356,N_28282);
or U28434 (N_28434,N_28277,N_28389);
or U28435 (N_28435,N_28278,N_28384);
xnor U28436 (N_28436,N_28251,N_28227);
xor U28437 (N_28437,N_28236,N_28293);
nor U28438 (N_28438,N_28247,N_28207);
xor U28439 (N_28439,N_28357,N_28381);
nand U28440 (N_28440,N_28245,N_28388);
or U28441 (N_28441,N_28229,N_28331);
and U28442 (N_28442,N_28274,N_28361);
or U28443 (N_28443,N_28326,N_28260);
nor U28444 (N_28444,N_28379,N_28279);
nand U28445 (N_28445,N_28281,N_28392);
or U28446 (N_28446,N_28237,N_28309);
or U28447 (N_28447,N_28209,N_28345);
xor U28448 (N_28448,N_28355,N_28217);
nor U28449 (N_28449,N_28390,N_28284);
or U28450 (N_28450,N_28200,N_28387);
xnor U28451 (N_28451,N_28259,N_28288);
xnor U28452 (N_28452,N_28346,N_28243);
nand U28453 (N_28453,N_28323,N_28380);
or U28454 (N_28454,N_28267,N_28220);
nand U28455 (N_28455,N_28241,N_28365);
and U28456 (N_28456,N_28248,N_28254);
nor U28457 (N_28457,N_28301,N_28335);
xor U28458 (N_28458,N_28359,N_28333);
and U28459 (N_28459,N_28395,N_28246);
nor U28460 (N_28460,N_28224,N_28332);
and U28461 (N_28461,N_28287,N_28351);
nand U28462 (N_28462,N_28340,N_28347);
or U28463 (N_28463,N_28258,N_28315);
nand U28464 (N_28464,N_28275,N_28368);
nand U28465 (N_28465,N_28295,N_28231);
xnor U28466 (N_28466,N_28364,N_28362);
and U28467 (N_28467,N_28250,N_28371);
or U28468 (N_28468,N_28268,N_28289);
xnor U28469 (N_28469,N_28348,N_28308);
nor U28470 (N_28470,N_28313,N_28385);
nor U28471 (N_28471,N_28375,N_28261);
and U28472 (N_28472,N_28226,N_28202);
xnor U28473 (N_28473,N_28285,N_28240);
or U28474 (N_28474,N_28262,N_28329);
xor U28475 (N_28475,N_28353,N_28307);
xnor U28476 (N_28476,N_28234,N_28235);
or U28477 (N_28477,N_28242,N_28215);
and U28478 (N_28478,N_28327,N_28264);
or U28479 (N_28479,N_28314,N_28213);
nand U28480 (N_28480,N_28272,N_28203);
nor U28481 (N_28481,N_28366,N_28298);
and U28482 (N_28482,N_28343,N_28310);
xnor U28483 (N_28483,N_28230,N_28350);
or U28484 (N_28484,N_28273,N_28201);
or U28485 (N_28485,N_28396,N_28354);
or U28486 (N_28486,N_28263,N_28219);
xor U28487 (N_28487,N_28214,N_28338);
and U28488 (N_28488,N_28399,N_28397);
or U28489 (N_28489,N_28311,N_28394);
or U28490 (N_28490,N_28360,N_28374);
nand U28491 (N_28491,N_28291,N_28318);
and U28492 (N_28492,N_28312,N_28238);
and U28493 (N_28493,N_28297,N_28216);
and U28494 (N_28494,N_28244,N_28296);
or U28495 (N_28495,N_28300,N_28342);
and U28496 (N_28496,N_28319,N_28253);
and U28497 (N_28497,N_28239,N_28221);
nand U28498 (N_28498,N_28232,N_28228);
nand U28499 (N_28499,N_28324,N_28398);
or U28500 (N_28500,N_28247,N_28320);
and U28501 (N_28501,N_28278,N_28373);
and U28502 (N_28502,N_28376,N_28222);
and U28503 (N_28503,N_28282,N_28347);
xnor U28504 (N_28504,N_28245,N_28221);
and U28505 (N_28505,N_28363,N_28213);
nand U28506 (N_28506,N_28263,N_28283);
or U28507 (N_28507,N_28341,N_28281);
nand U28508 (N_28508,N_28340,N_28391);
nor U28509 (N_28509,N_28368,N_28313);
xnor U28510 (N_28510,N_28248,N_28205);
xor U28511 (N_28511,N_28249,N_28331);
or U28512 (N_28512,N_28326,N_28319);
and U28513 (N_28513,N_28215,N_28235);
nor U28514 (N_28514,N_28210,N_28357);
and U28515 (N_28515,N_28295,N_28348);
and U28516 (N_28516,N_28275,N_28257);
or U28517 (N_28517,N_28301,N_28213);
xor U28518 (N_28518,N_28313,N_28265);
or U28519 (N_28519,N_28325,N_28220);
xnor U28520 (N_28520,N_28273,N_28245);
nor U28521 (N_28521,N_28364,N_28250);
nand U28522 (N_28522,N_28217,N_28335);
nor U28523 (N_28523,N_28364,N_28271);
nand U28524 (N_28524,N_28294,N_28371);
nor U28525 (N_28525,N_28384,N_28366);
xor U28526 (N_28526,N_28297,N_28224);
nand U28527 (N_28527,N_28377,N_28357);
xor U28528 (N_28528,N_28227,N_28234);
and U28529 (N_28529,N_28353,N_28320);
nand U28530 (N_28530,N_28246,N_28269);
and U28531 (N_28531,N_28367,N_28223);
and U28532 (N_28532,N_28376,N_28371);
and U28533 (N_28533,N_28395,N_28346);
nor U28534 (N_28534,N_28280,N_28388);
or U28535 (N_28535,N_28278,N_28392);
nor U28536 (N_28536,N_28300,N_28285);
and U28537 (N_28537,N_28347,N_28389);
nand U28538 (N_28538,N_28291,N_28264);
nor U28539 (N_28539,N_28349,N_28245);
or U28540 (N_28540,N_28354,N_28216);
nor U28541 (N_28541,N_28399,N_28234);
nand U28542 (N_28542,N_28248,N_28382);
and U28543 (N_28543,N_28347,N_28365);
or U28544 (N_28544,N_28395,N_28323);
nand U28545 (N_28545,N_28202,N_28300);
nor U28546 (N_28546,N_28344,N_28264);
nand U28547 (N_28547,N_28249,N_28267);
or U28548 (N_28548,N_28335,N_28356);
xor U28549 (N_28549,N_28208,N_28226);
nand U28550 (N_28550,N_28363,N_28367);
nor U28551 (N_28551,N_28362,N_28248);
or U28552 (N_28552,N_28226,N_28369);
or U28553 (N_28553,N_28215,N_28320);
and U28554 (N_28554,N_28362,N_28315);
or U28555 (N_28555,N_28330,N_28252);
or U28556 (N_28556,N_28253,N_28371);
nor U28557 (N_28557,N_28323,N_28265);
xnor U28558 (N_28558,N_28346,N_28399);
nand U28559 (N_28559,N_28246,N_28279);
and U28560 (N_28560,N_28327,N_28228);
and U28561 (N_28561,N_28370,N_28309);
nor U28562 (N_28562,N_28327,N_28300);
nand U28563 (N_28563,N_28359,N_28336);
or U28564 (N_28564,N_28231,N_28259);
or U28565 (N_28565,N_28241,N_28266);
and U28566 (N_28566,N_28373,N_28322);
xor U28567 (N_28567,N_28282,N_28352);
nor U28568 (N_28568,N_28242,N_28321);
xnor U28569 (N_28569,N_28336,N_28209);
nor U28570 (N_28570,N_28302,N_28271);
nand U28571 (N_28571,N_28350,N_28382);
and U28572 (N_28572,N_28298,N_28228);
or U28573 (N_28573,N_28338,N_28340);
nor U28574 (N_28574,N_28399,N_28334);
nor U28575 (N_28575,N_28214,N_28244);
and U28576 (N_28576,N_28329,N_28296);
nand U28577 (N_28577,N_28345,N_28266);
or U28578 (N_28578,N_28336,N_28248);
xnor U28579 (N_28579,N_28377,N_28254);
or U28580 (N_28580,N_28223,N_28345);
xnor U28581 (N_28581,N_28206,N_28212);
nor U28582 (N_28582,N_28280,N_28282);
or U28583 (N_28583,N_28300,N_28398);
and U28584 (N_28584,N_28348,N_28360);
nor U28585 (N_28585,N_28290,N_28268);
nand U28586 (N_28586,N_28346,N_28218);
and U28587 (N_28587,N_28206,N_28305);
and U28588 (N_28588,N_28265,N_28269);
nor U28589 (N_28589,N_28336,N_28387);
nor U28590 (N_28590,N_28269,N_28360);
nor U28591 (N_28591,N_28223,N_28377);
and U28592 (N_28592,N_28263,N_28361);
or U28593 (N_28593,N_28215,N_28205);
xor U28594 (N_28594,N_28231,N_28226);
or U28595 (N_28595,N_28398,N_28356);
nand U28596 (N_28596,N_28297,N_28335);
nand U28597 (N_28597,N_28253,N_28268);
nand U28598 (N_28598,N_28325,N_28266);
xnor U28599 (N_28599,N_28342,N_28239);
xor U28600 (N_28600,N_28426,N_28468);
or U28601 (N_28601,N_28408,N_28525);
or U28602 (N_28602,N_28479,N_28497);
nand U28603 (N_28603,N_28466,N_28577);
or U28604 (N_28604,N_28549,N_28597);
or U28605 (N_28605,N_28480,N_28578);
and U28606 (N_28606,N_28512,N_28505);
xor U28607 (N_28607,N_28588,N_28552);
or U28608 (N_28608,N_28403,N_28483);
xnor U28609 (N_28609,N_28493,N_28567);
nand U28610 (N_28610,N_28532,N_28438);
nor U28611 (N_28611,N_28470,N_28490);
nor U28612 (N_28612,N_28478,N_28410);
and U28613 (N_28613,N_28414,N_28432);
or U28614 (N_28614,N_28436,N_28526);
and U28615 (N_28615,N_28407,N_28443);
or U28616 (N_28616,N_28545,N_28553);
xnor U28617 (N_28617,N_28457,N_28402);
and U28618 (N_28618,N_28596,N_28535);
or U28619 (N_28619,N_28467,N_28430);
and U28620 (N_28620,N_28435,N_28458);
and U28621 (N_28621,N_28453,N_28562);
and U28622 (N_28622,N_28531,N_28476);
nand U28623 (N_28623,N_28534,N_28513);
and U28624 (N_28624,N_28474,N_28557);
nor U28625 (N_28625,N_28489,N_28570);
and U28626 (N_28626,N_28541,N_28548);
and U28627 (N_28627,N_28580,N_28439);
nand U28628 (N_28628,N_28496,N_28565);
xor U28629 (N_28629,N_28437,N_28592);
nand U28630 (N_28630,N_28550,N_28451);
xnor U28631 (N_28631,N_28584,N_28487);
and U28632 (N_28632,N_28423,N_28463);
and U28633 (N_28633,N_28576,N_28581);
xor U28634 (N_28634,N_28546,N_28415);
xor U28635 (N_28635,N_28412,N_28447);
and U28636 (N_28636,N_28507,N_28593);
or U28637 (N_28637,N_28573,N_28523);
and U28638 (N_28638,N_28564,N_28509);
or U28639 (N_28639,N_28568,N_28456);
xor U28640 (N_28640,N_28405,N_28522);
nor U28641 (N_28641,N_28400,N_28506);
or U28642 (N_28642,N_28599,N_28477);
xor U28643 (N_28643,N_28518,N_28559);
nor U28644 (N_28644,N_28589,N_28401);
xor U28645 (N_28645,N_28529,N_28419);
and U28646 (N_28646,N_28571,N_28475);
nand U28647 (N_28647,N_28533,N_28500);
xnor U28648 (N_28648,N_28462,N_28465);
or U28649 (N_28649,N_28498,N_28538);
nor U28650 (N_28650,N_28574,N_28417);
xor U28651 (N_28651,N_28520,N_28502);
nand U28652 (N_28652,N_28488,N_28404);
nand U28653 (N_28653,N_28544,N_28455);
and U28654 (N_28654,N_28411,N_28424);
or U28655 (N_28655,N_28555,N_28585);
or U28656 (N_28656,N_28537,N_28547);
xnor U28657 (N_28657,N_28421,N_28459);
or U28658 (N_28658,N_28495,N_28521);
nor U28659 (N_28659,N_28440,N_28485);
nor U28660 (N_28660,N_28563,N_28575);
and U28661 (N_28661,N_28418,N_28482);
or U28662 (N_28662,N_28527,N_28514);
nand U28663 (N_28663,N_28422,N_28413);
nor U28664 (N_28664,N_28528,N_28586);
nand U28665 (N_28665,N_28554,N_28539);
nand U28666 (N_28666,N_28484,N_28454);
and U28667 (N_28667,N_28591,N_28543);
and U28668 (N_28668,N_28446,N_28460);
or U28669 (N_28669,N_28595,N_28444);
and U28670 (N_28670,N_28569,N_28464);
xnor U28671 (N_28671,N_28556,N_28433);
or U28672 (N_28672,N_28420,N_28434);
xor U28673 (N_28673,N_28579,N_28510);
xor U28674 (N_28674,N_28486,N_28530);
xor U28675 (N_28675,N_28504,N_28516);
and U28676 (N_28676,N_28540,N_28425);
xnor U28677 (N_28677,N_28450,N_28469);
xnor U28678 (N_28678,N_28508,N_28501);
xor U28679 (N_28679,N_28448,N_28471);
nand U28680 (N_28680,N_28449,N_28481);
xnor U28681 (N_28681,N_28594,N_28566);
nand U28682 (N_28682,N_28572,N_28558);
nor U28683 (N_28683,N_28409,N_28511);
nand U28684 (N_28684,N_28517,N_28561);
and U28685 (N_28685,N_28429,N_28542);
or U28686 (N_28686,N_28445,N_28428);
nand U28687 (N_28687,N_28491,N_28431);
nor U28688 (N_28688,N_28452,N_28442);
or U28689 (N_28689,N_28472,N_28590);
nor U28690 (N_28690,N_28587,N_28427);
xor U28691 (N_28691,N_28461,N_28416);
nor U28692 (N_28692,N_28583,N_28598);
and U28693 (N_28693,N_28536,N_28503);
nor U28694 (N_28694,N_28551,N_28494);
or U28695 (N_28695,N_28582,N_28499);
xor U28696 (N_28696,N_28519,N_28515);
and U28697 (N_28697,N_28441,N_28473);
or U28698 (N_28698,N_28560,N_28406);
nand U28699 (N_28699,N_28492,N_28524);
nor U28700 (N_28700,N_28405,N_28403);
or U28701 (N_28701,N_28590,N_28402);
nor U28702 (N_28702,N_28497,N_28532);
xnor U28703 (N_28703,N_28465,N_28504);
xnor U28704 (N_28704,N_28461,N_28465);
nand U28705 (N_28705,N_28430,N_28568);
xor U28706 (N_28706,N_28413,N_28479);
xnor U28707 (N_28707,N_28566,N_28407);
and U28708 (N_28708,N_28431,N_28441);
xor U28709 (N_28709,N_28543,N_28538);
and U28710 (N_28710,N_28587,N_28540);
xor U28711 (N_28711,N_28463,N_28483);
or U28712 (N_28712,N_28487,N_28571);
nor U28713 (N_28713,N_28510,N_28598);
or U28714 (N_28714,N_28521,N_28523);
nor U28715 (N_28715,N_28586,N_28498);
and U28716 (N_28716,N_28507,N_28560);
xor U28717 (N_28717,N_28427,N_28496);
nand U28718 (N_28718,N_28484,N_28476);
nor U28719 (N_28719,N_28453,N_28454);
and U28720 (N_28720,N_28425,N_28576);
xor U28721 (N_28721,N_28573,N_28519);
nand U28722 (N_28722,N_28572,N_28498);
and U28723 (N_28723,N_28469,N_28574);
nor U28724 (N_28724,N_28475,N_28440);
nor U28725 (N_28725,N_28572,N_28434);
or U28726 (N_28726,N_28497,N_28425);
or U28727 (N_28727,N_28416,N_28410);
and U28728 (N_28728,N_28463,N_28487);
nand U28729 (N_28729,N_28514,N_28542);
xor U28730 (N_28730,N_28590,N_28535);
or U28731 (N_28731,N_28494,N_28516);
or U28732 (N_28732,N_28513,N_28565);
and U28733 (N_28733,N_28449,N_28580);
or U28734 (N_28734,N_28593,N_28408);
nand U28735 (N_28735,N_28450,N_28472);
nor U28736 (N_28736,N_28596,N_28548);
nand U28737 (N_28737,N_28407,N_28484);
xnor U28738 (N_28738,N_28588,N_28587);
and U28739 (N_28739,N_28541,N_28485);
nor U28740 (N_28740,N_28413,N_28585);
and U28741 (N_28741,N_28424,N_28534);
xor U28742 (N_28742,N_28432,N_28496);
xor U28743 (N_28743,N_28426,N_28412);
xor U28744 (N_28744,N_28568,N_28555);
or U28745 (N_28745,N_28573,N_28542);
nand U28746 (N_28746,N_28507,N_28540);
and U28747 (N_28747,N_28444,N_28522);
or U28748 (N_28748,N_28479,N_28434);
or U28749 (N_28749,N_28447,N_28516);
xnor U28750 (N_28750,N_28523,N_28486);
nor U28751 (N_28751,N_28567,N_28523);
nand U28752 (N_28752,N_28566,N_28562);
xnor U28753 (N_28753,N_28504,N_28474);
and U28754 (N_28754,N_28443,N_28461);
nand U28755 (N_28755,N_28597,N_28518);
nand U28756 (N_28756,N_28482,N_28511);
nand U28757 (N_28757,N_28416,N_28530);
or U28758 (N_28758,N_28494,N_28580);
xnor U28759 (N_28759,N_28557,N_28404);
nand U28760 (N_28760,N_28405,N_28597);
or U28761 (N_28761,N_28486,N_28448);
nand U28762 (N_28762,N_28547,N_28488);
nand U28763 (N_28763,N_28532,N_28404);
xnor U28764 (N_28764,N_28474,N_28488);
nand U28765 (N_28765,N_28525,N_28495);
nor U28766 (N_28766,N_28418,N_28479);
nand U28767 (N_28767,N_28599,N_28471);
nand U28768 (N_28768,N_28430,N_28567);
xnor U28769 (N_28769,N_28509,N_28574);
nand U28770 (N_28770,N_28404,N_28459);
nand U28771 (N_28771,N_28561,N_28466);
and U28772 (N_28772,N_28572,N_28587);
nor U28773 (N_28773,N_28544,N_28448);
xor U28774 (N_28774,N_28466,N_28410);
nand U28775 (N_28775,N_28455,N_28588);
xnor U28776 (N_28776,N_28593,N_28473);
nor U28777 (N_28777,N_28477,N_28484);
and U28778 (N_28778,N_28509,N_28594);
nand U28779 (N_28779,N_28472,N_28479);
or U28780 (N_28780,N_28525,N_28583);
nor U28781 (N_28781,N_28426,N_28475);
nand U28782 (N_28782,N_28597,N_28474);
xnor U28783 (N_28783,N_28572,N_28477);
and U28784 (N_28784,N_28421,N_28580);
and U28785 (N_28785,N_28456,N_28590);
nand U28786 (N_28786,N_28543,N_28438);
nand U28787 (N_28787,N_28525,N_28497);
nand U28788 (N_28788,N_28433,N_28412);
nor U28789 (N_28789,N_28411,N_28513);
nand U28790 (N_28790,N_28564,N_28552);
nand U28791 (N_28791,N_28433,N_28512);
nand U28792 (N_28792,N_28425,N_28599);
or U28793 (N_28793,N_28460,N_28558);
and U28794 (N_28794,N_28599,N_28443);
and U28795 (N_28795,N_28490,N_28408);
or U28796 (N_28796,N_28418,N_28422);
and U28797 (N_28797,N_28518,N_28400);
nand U28798 (N_28798,N_28433,N_28414);
xnor U28799 (N_28799,N_28521,N_28589);
xor U28800 (N_28800,N_28655,N_28686);
xor U28801 (N_28801,N_28799,N_28648);
and U28802 (N_28802,N_28727,N_28628);
and U28803 (N_28803,N_28735,N_28640);
xor U28804 (N_28804,N_28693,N_28695);
or U28805 (N_28805,N_28713,N_28688);
or U28806 (N_28806,N_28613,N_28672);
nand U28807 (N_28807,N_28758,N_28651);
xnor U28808 (N_28808,N_28793,N_28738);
nand U28809 (N_28809,N_28742,N_28615);
or U28810 (N_28810,N_28700,N_28631);
nand U28811 (N_28811,N_28662,N_28682);
nor U28812 (N_28812,N_28726,N_28683);
xor U28813 (N_28813,N_28756,N_28654);
nand U28814 (N_28814,N_28754,N_28685);
nand U28815 (N_28815,N_28603,N_28743);
nand U28816 (N_28816,N_28600,N_28678);
nor U28817 (N_28817,N_28666,N_28730);
xor U28818 (N_28818,N_28724,N_28676);
xnor U28819 (N_28819,N_28755,N_28767);
nand U28820 (N_28820,N_28771,N_28733);
xor U28821 (N_28821,N_28670,N_28636);
or U28822 (N_28822,N_28680,N_28750);
nor U28823 (N_28823,N_28798,N_28637);
nand U28824 (N_28824,N_28759,N_28617);
nor U28825 (N_28825,N_28790,N_28772);
nand U28826 (N_28826,N_28620,N_28657);
nand U28827 (N_28827,N_28792,N_28629);
or U28828 (N_28828,N_28737,N_28720);
or U28829 (N_28829,N_28736,N_28739);
nor U28830 (N_28830,N_28639,N_28766);
nand U28831 (N_28831,N_28622,N_28797);
nor U28832 (N_28832,N_28644,N_28709);
xor U28833 (N_28833,N_28770,N_28674);
and U28834 (N_28834,N_28669,N_28769);
or U28835 (N_28835,N_28635,N_28722);
and U28836 (N_28836,N_28747,N_28623);
xor U28837 (N_28837,N_28647,N_28675);
xnor U28838 (N_28838,N_28712,N_28661);
xnor U28839 (N_28839,N_28701,N_28783);
and U28840 (N_28840,N_28760,N_28786);
xor U28841 (N_28841,N_28723,N_28681);
and U28842 (N_28842,N_28717,N_28660);
and U28843 (N_28843,N_28784,N_28716);
nand U28844 (N_28844,N_28734,N_28610);
nand U28845 (N_28845,N_28665,N_28656);
or U28846 (N_28846,N_28638,N_28630);
nor U28847 (N_28847,N_28626,N_28751);
and U28848 (N_28848,N_28643,N_28663);
xor U28849 (N_28849,N_28763,N_28787);
nor U28850 (N_28850,N_28791,N_28746);
and U28851 (N_28851,N_28778,N_28621);
nand U28852 (N_28852,N_28782,N_28796);
xnor U28853 (N_28853,N_28697,N_28616);
nand U28854 (N_28854,N_28728,N_28602);
xnor U28855 (N_28855,N_28773,N_28689);
and U28856 (N_28856,N_28625,N_28671);
and U28857 (N_28857,N_28627,N_28764);
nand U28858 (N_28858,N_28677,N_28725);
nand U28859 (N_28859,N_28707,N_28776);
and U28860 (N_28860,N_28794,N_28761);
or U28861 (N_28861,N_28774,N_28719);
nand U28862 (N_28862,N_28609,N_28789);
nor U28863 (N_28863,N_28698,N_28729);
or U28864 (N_28864,N_28658,N_28641);
and U28865 (N_28865,N_28624,N_28748);
and U28866 (N_28866,N_28606,N_28731);
nand U28867 (N_28867,N_28684,N_28777);
and U28868 (N_28868,N_28646,N_28645);
xnor U28869 (N_28869,N_28668,N_28704);
xor U28870 (N_28870,N_28705,N_28718);
nand U28871 (N_28871,N_28633,N_28741);
xor U28872 (N_28872,N_28740,N_28673);
nand U28873 (N_28873,N_28604,N_28702);
nand U28874 (N_28874,N_28618,N_28692);
xnor U28875 (N_28875,N_28775,N_28752);
nand U28876 (N_28876,N_28788,N_28785);
nand U28877 (N_28877,N_28765,N_28614);
or U28878 (N_28878,N_28652,N_28650);
nor U28879 (N_28879,N_28649,N_28753);
nand U28880 (N_28880,N_28659,N_28781);
or U28881 (N_28881,N_28711,N_28653);
xnor U28882 (N_28882,N_28679,N_28696);
nand U28883 (N_28883,N_28642,N_28611);
nor U28884 (N_28884,N_28708,N_28703);
xnor U28885 (N_28885,N_28608,N_28632);
or U28886 (N_28886,N_28779,N_28710);
and U28887 (N_28887,N_28732,N_28768);
and U28888 (N_28888,N_28612,N_28667);
xor U28889 (N_28889,N_28721,N_28714);
xor U28890 (N_28890,N_28706,N_28757);
and U28891 (N_28891,N_28744,N_28601);
nand U28892 (N_28892,N_28687,N_28715);
and U28893 (N_28893,N_28691,N_28749);
or U28894 (N_28894,N_28699,N_28605);
xnor U28895 (N_28895,N_28619,N_28795);
xnor U28896 (N_28896,N_28745,N_28664);
and U28897 (N_28897,N_28690,N_28634);
and U28898 (N_28898,N_28694,N_28762);
or U28899 (N_28899,N_28780,N_28607);
or U28900 (N_28900,N_28696,N_28790);
xnor U28901 (N_28901,N_28640,N_28707);
xor U28902 (N_28902,N_28745,N_28737);
or U28903 (N_28903,N_28767,N_28693);
nand U28904 (N_28904,N_28690,N_28660);
nand U28905 (N_28905,N_28610,N_28673);
nand U28906 (N_28906,N_28755,N_28621);
and U28907 (N_28907,N_28772,N_28681);
nor U28908 (N_28908,N_28655,N_28767);
nand U28909 (N_28909,N_28696,N_28714);
nor U28910 (N_28910,N_28668,N_28638);
nand U28911 (N_28911,N_28601,N_28673);
and U28912 (N_28912,N_28779,N_28794);
xnor U28913 (N_28913,N_28677,N_28627);
or U28914 (N_28914,N_28647,N_28736);
xnor U28915 (N_28915,N_28709,N_28742);
nor U28916 (N_28916,N_28666,N_28705);
and U28917 (N_28917,N_28645,N_28719);
xor U28918 (N_28918,N_28794,N_28676);
nor U28919 (N_28919,N_28608,N_28770);
nor U28920 (N_28920,N_28611,N_28678);
nand U28921 (N_28921,N_28724,N_28704);
or U28922 (N_28922,N_28628,N_28720);
nor U28923 (N_28923,N_28757,N_28740);
nor U28924 (N_28924,N_28711,N_28683);
nand U28925 (N_28925,N_28726,N_28655);
nand U28926 (N_28926,N_28696,N_28663);
or U28927 (N_28927,N_28781,N_28600);
nor U28928 (N_28928,N_28601,N_28732);
and U28929 (N_28929,N_28785,N_28680);
and U28930 (N_28930,N_28608,N_28745);
nor U28931 (N_28931,N_28716,N_28674);
nand U28932 (N_28932,N_28681,N_28649);
and U28933 (N_28933,N_28785,N_28760);
nand U28934 (N_28934,N_28643,N_28661);
nor U28935 (N_28935,N_28677,N_28695);
and U28936 (N_28936,N_28614,N_28783);
nand U28937 (N_28937,N_28677,N_28607);
nor U28938 (N_28938,N_28795,N_28725);
xnor U28939 (N_28939,N_28675,N_28636);
nor U28940 (N_28940,N_28646,N_28794);
and U28941 (N_28941,N_28622,N_28657);
or U28942 (N_28942,N_28762,N_28676);
or U28943 (N_28943,N_28712,N_28721);
xnor U28944 (N_28944,N_28705,N_28622);
and U28945 (N_28945,N_28665,N_28664);
or U28946 (N_28946,N_28750,N_28755);
and U28947 (N_28947,N_28665,N_28796);
nor U28948 (N_28948,N_28649,N_28733);
or U28949 (N_28949,N_28681,N_28628);
and U28950 (N_28950,N_28761,N_28655);
nand U28951 (N_28951,N_28767,N_28716);
nand U28952 (N_28952,N_28672,N_28725);
and U28953 (N_28953,N_28791,N_28602);
nand U28954 (N_28954,N_28735,N_28683);
or U28955 (N_28955,N_28763,N_28690);
xor U28956 (N_28956,N_28741,N_28797);
or U28957 (N_28957,N_28747,N_28668);
and U28958 (N_28958,N_28620,N_28777);
nand U28959 (N_28959,N_28750,N_28738);
nand U28960 (N_28960,N_28621,N_28631);
nor U28961 (N_28961,N_28709,N_28659);
or U28962 (N_28962,N_28745,N_28727);
or U28963 (N_28963,N_28791,N_28629);
or U28964 (N_28964,N_28731,N_28667);
or U28965 (N_28965,N_28705,N_28667);
nand U28966 (N_28966,N_28719,N_28782);
nand U28967 (N_28967,N_28613,N_28637);
nand U28968 (N_28968,N_28710,N_28679);
or U28969 (N_28969,N_28722,N_28653);
nand U28970 (N_28970,N_28712,N_28713);
and U28971 (N_28971,N_28751,N_28745);
xnor U28972 (N_28972,N_28685,N_28647);
or U28973 (N_28973,N_28755,N_28717);
nor U28974 (N_28974,N_28723,N_28717);
nand U28975 (N_28975,N_28672,N_28683);
and U28976 (N_28976,N_28731,N_28703);
nor U28977 (N_28977,N_28614,N_28604);
and U28978 (N_28978,N_28679,N_28719);
nor U28979 (N_28979,N_28661,N_28744);
nand U28980 (N_28980,N_28739,N_28634);
or U28981 (N_28981,N_28784,N_28640);
nor U28982 (N_28982,N_28712,N_28761);
nor U28983 (N_28983,N_28773,N_28726);
or U28984 (N_28984,N_28773,N_28714);
nor U28985 (N_28985,N_28702,N_28607);
nor U28986 (N_28986,N_28607,N_28786);
nor U28987 (N_28987,N_28785,N_28648);
and U28988 (N_28988,N_28620,N_28714);
nor U28989 (N_28989,N_28795,N_28744);
nor U28990 (N_28990,N_28773,N_28684);
xnor U28991 (N_28991,N_28774,N_28664);
and U28992 (N_28992,N_28707,N_28761);
nor U28993 (N_28993,N_28697,N_28706);
xor U28994 (N_28994,N_28715,N_28672);
or U28995 (N_28995,N_28733,N_28792);
xor U28996 (N_28996,N_28729,N_28639);
or U28997 (N_28997,N_28613,N_28612);
and U28998 (N_28998,N_28647,N_28735);
xor U28999 (N_28999,N_28671,N_28650);
xor U29000 (N_29000,N_28890,N_28906);
nand U29001 (N_29001,N_28991,N_28836);
nor U29002 (N_29002,N_28850,N_28893);
nand U29003 (N_29003,N_28925,N_28889);
nor U29004 (N_29004,N_28897,N_28873);
xor U29005 (N_29005,N_28984,N_28804);
nor U29006 (N_29006,N_28802,N_28999);
and U29007 (N_29007,N_28884,N_28855);
nor U29008 (N_29008,N_28932,N_28911);
or U29009 (N_29009,N_28910,N_28950);
and U29010 (N_29010,N_28819,N_28908);
nor U29011 (N_29011,N_28875,N_28936);
xnor U29012 (N_29012,N_28805,N_28961);
nand U29013 (N_29013,N_28979,N_28913);
and U29014 (N_29014,N_28833,N_28982);
or U29015 (N_29015,N_28864,N_28993);
nand U29016 (N_29016,N_28807,N_28837);
and U29017 (N_29017,N_28972,N_28831);
xnor U29018 (N_29018,N_28958,N_28959);
or U29019 (N_29019,N_28813,N_28983);
and U29020 (N_29020,N_28944,N_28960);
xnor U29021 (N_29021,N_28929,N_28964);
or U29022 (N_29022,N_28834,N_28814);
nor U29023 (N_29023,N_28882,N_28947);
or U29024 (N_29024,N_28871,N_28969);
or U29025 (N_29025,N_28894,N_28899);
nor U29026 (N_29026,N_28803,N_28851);
xnor U29027 (N_29027,N_28902,N_28973);
xnor U29028 (N_29028,N_28967,N_28892);
or U29029 (N_29029,N_28918,N_28857);
and U29030 (N_29030,N_28885,N_28867);
and U29031 (N_29031,N_28863,N_28916);
or U29032 (N_29032,N_28801,N_28954);
or U29033 (N_29033,N_28841,N_28981);
or U29034 (N_29034,N_28974,N_28975);
nor U29035 (N_29035,N_28856,N_28905);
nor U29036 (N_29036,N_28806,N_28881);
or U29037 (N_29037,N_28956,N_28879);
nand U29038 (N_29038,N_28962,N_28827);
and U29039 (N_29039,N_28848,N_28996);
nand U29040 (N_29040,N_28858,N_28994);
nor U29041 (N_29041,N_28872,N_28939);
or U29042 (N_29042,N_28989,N_28970);
nand U29043 (N_29043,N_28933,N_28976);
nor U29044 (N_29044,N_28965,N_28883);
nor U29045 (N_29045,N_28809,N_28840);
nand U29046 (N_29046,N_28832,N_28852);
nand U29047 (N_29047,N_28868,N_28869);
xnor U29048 (N_29048,N_28912,N_28854);
nand U29049 (N_29049,N_28921,N_28937);
and U29050 (N_29050,N_28943,N_28919);
or U29051 (N_29051,N_28823,N_28824);
xor U29052 (N_29052,N_28971,N_28904);
nor U29053 (N_29053,N_28810,N_28862);
nor U29054 (N_29054,N_28920,N_28928);
nor U29055 (N_29055,N_28949,N_28845);
or U29056 (N_29056,N_28818,N_28930);
xnor U29057 (N_29057,N_28992,N_28865);
nand U29058 (N_29058,N_28825,N_28843);
and U29059 (N_29059,N_28900,N_28822);
or U29060 (N_29060,N_28842,N_28812);
and U29061 (N_29061,N_28927,N_28938);
nor U29062 (N_29062,N_28980,N_28820);
or U29063 (N_29063,N_28977,N_28859);
and U29064 (N_29064,N_28821,N_28838);
nand U29065 (N_29065,N_28826,N_28895);
nor U29066 (N_29066,N_28901,N_28876);
or U29067 (N_29067,N_28909,N_28934);
xnor U29068 (N_29068,N_28829,N_28839);
nand U29069 (N_29069,N_28877,N_28835);
nor U29070 (N_29070,N_28811,N_28953);
and U29071 (N_29071,N_28997,N_28963);
or U29072 (N_29072,N_28907,N_28887);
or U29073 (N_29073,N_28931,N_28870);
and U29074 (N_29074,N_28861,N_28800);
and U29075 (N_29075,N_28998,N_28874);
nor U29076 (N_29076,N_28952,N_28985);
nand U29077 (N_29077,N_28987,N_28828);
xnor U29078 (N_29078,N_28817,N_28955);
nand U29079 (N_29079,N_28966,N_28888);
and U29080 (N_29080,N_28986,N_28923);
and U29081 (N_29081,N_28896,N_28924);
and U29082 (N_29082,N_28880,N_28847);
nand U29083 (N_29083,N_28844,N_28951);
and U29084 (N_29084,N_28903,N_28915);
and U29085 (N_29085,N_28878,N_28808);
and U29086 (N_29086,N_28816,N_28957);
nand U29087 (N_29087,N_28891,N_28898);
nor U29088 (N_29088,N_28990,N_28830);
and U29089 (N_29089,N_28945,N_28860);
nor U29090 (N_29090,N_28846,N_28940);
nor U29091 (N_29091,N_28815,N_28914);
or U29092 (N_29092,N_28849,N_28941);
nor U29093 (N_29093,N_28988,N_28886);
or U29094 (N_29094,N_28948,N_28866);
nor U29095 (N_29095,N_28995,N_28917);
and U29096 (N_29096,N_28935,N_28946);
nor U29097 (N_29097,N_28978,N_28942);
or U29098 (N_29098,N_28853,N_28926);
nor U29099 (N_29099,N_28968,N_28922);
nor U29100 (N_29100,N_28893,N_28855);
xnor U29101 (N_29101,N_28830,N_28805);
and U29102 (N_29102,N_28964,N_28865);
xor U29103 (N_29103,N_28943,N_28932);
xnor U29104 (N_29104,N_28946,N_28821);
xnor U29105 (N_29105,N_28865,N_28968);
nor U29106 (N_29106,N_28999,N_28893);
nor U29107 (N_29107,N_28941,N_28997);
nand U29108 (N_29108,N_28972,N_28889);
xor U29109 (N_29109,N_28821,N_28904);
or U29110 (N_29110,N_28807,N_28968);
nand U29111 (N_29111,N_28985,N_28890);
or U29112 (N_29112,N_28873,N_28993);
nand U29113 (N_29113,N_28862,N_28912);
xor U29114 (N_29114,N_28835,N_28912);
and U29115 (N_29115,N_28942,N_28882);
xnor U29116 (N_29116,N_28864,N_28822);
and U29117 (N_29117,N_28918,N_28964);
nor U29118 (N_29118,N_28968,N_28941);
nand U29119 (N_29119,N_28976,N_28854);
nand U29120 (N_29120,N_28998,N_28841);
and U29121 (N_29121,N_28903,N_28871);
and U29122 (N_29122,N_28843,N_28830);
or U29123 (N_29123,N_28908,N_28941);
or U29124 (N_29124,N_28979,N_28859);
and U29125 (N_29125,N_28967,N_28801);
or U29126 (N_29126,N_28811,N_28848);
or U29127 (N_29127,N_28849,N_28817);
nand U29128 (N_29128,N_28905,N_28915);
nor U29129 (N_29129,N_28953,N_28871);
xnor U29130 (N_29130,N_28837,N_28925);
nor U29131 (N_29131,N_28841,N_28938);
or U29132 (N_29132,N_28929,N_28806);
or U29133 (N_29133,N_28929,N_28979);
and U29134 (N_29134,N_28871,N_28958);
nor U29135 (N_29135,N_28879,N_28853);
and U29136 (N_29136,N_28849,N_28968);
xor U29137 (N_29137,N_28803,N_28972);
xnor U29138 (N_29138,N_28994,N_28941);
xnor U29139 (N_29139,N_28906,N_28813);
xor U29140 (N_29140,N_28807,N_28953);
xnor U29141 (N_29141,N_28832,N_28887);
and U29142 (N_29142,N_28923,N_28942);
or U29143 (N_29143,N_28834,N_28916);
nand U29144 (N_29144,N_28875,N_28975);
and U29145 (N_29145,N_28816,N_28863);
nand U29146 (N_29146,N_28809,N_28802);
nor U29147 (N_29147,N_28809,N_28907);
and U29148 (N_29148,N_28982,N_28963);
or U29149 (N_29149,N_28962,N_28952);
nand U29150 (N_29150,N_28934,N_28802);
and U29151 (N_29151,N_28801,N_28883);
and U29152 (N_29152,N_28963,N_28999);
nand U29153 (N_29153,N_28857,N_28901);
and U29154 (N_29154,N_28802,N_28909);
nand U29155 (N_29155,N_28899,N_28904);
nor U29156 (N_29156,N_28965,N_28934);
and U29157 (N_29157,N_28910,N_28880);
nor U29158 (N_29158,N_28879,N_28833);
or U29159 (N_29159,N_28982,N_28991);
nand U29160 (N_29160,N_28952,N_28819);
nor U29161 (N_29161,N_28909,N_28974);
xnor U29162 (N_29162,N_28803,N_28839);
nor U29163 (N_29163,N_28832,N_28800);
nor U29164 (N_29164,N_28875,N_28911);
and U29165 (N_29165,N_28914,N_28871);
and U29166 (N_29166,N_28881,N_28938);
nand U29167 (N_29167,N_28847,N_28920);
or U29168 (N_29168,N_28925,N_28933);
nor U29169 (N_29169,N_28811,N_28919);
nor U29170 (N_29170,N_28847,N_28975);
xnor U29171 (N_29171,N_28997,N_28896);
and U29172 (N_29172,N_28946,N_28917);
and U29173 (N_29173,N_28824,N_28813);
nor U29174 (N_29174,N_28957,N_28873);
and U29175 (N_29175,N_28953,N_28892);
and U29176 (N_29176,N_28948,N_28832);
and U29177 (N_29177,N_28956,N_28934);
nand U29178 (N_29178,N_28927,N_28954);
or U29179 (N_29179,N_28807,N_28864);
nor U29180 (N_29180,N_28915,N_28934);
nand U29181 (N_29181,N_28871,N_28971);
nor U29182 (N_29182,N_28834,N_28860);
or U29183 (N_29183,N_28833,N_28929);
nor U29184 (N_29184,N_28919,N_28839);
nand U29185 (N_29185,N_28814,N_28804);
nor U29186 (N_29186,N_28966,N_28823);
and U29187 (N_29187,N_28828,N_28803);
xnor U29188 (N_29188,N_28809,N_28899);
nand U29189 (N_29189,N_28933,N_28877);
xor U29190 (N_29190,N_28841,N_28815);
xor U29191 (N_29191,N_28845,N_28864);
nor U29192 (N_29192,N_28959,N_28951);
or U29193 (N_29193,N_28977,N_28956);
nor U29194 (N_29194,N_28989,N_28935);
and U29195 (N_29195,N_28977,N_28964);
and U29196 (N_29196,N_28927,N_28803);
or U29197 (N_29197,N_28832,N_28938);
or U29198 (N_29198,N_28819,N_28938);
nor U29199 (N_29199,N_28897,N_28953);
and U29200 (N_29200,N_29161,N_29146);
xor U29201 (N_29201,N_29098,N_29102);
nand U29202 (N_29202,N_29068,N_29075);
and U29203 (N_29203,N_29114,N_29083);
and U29204 (N_29204,N_29108,N_29174);
and U29205 (N_29205,N_29086,N_29096);
xnor U29206 (N_29206,N_29077,N_29131);
and U29207 (N_29207,N_29142,N_29165);
and U29208 (N_29208,N_29121,N_29011);
nand U29209 (N_29209,N_29125,N_29040);
nor U29210 (N_29210,N_29107,N_29028);
nor U29211 (N_29211,N_29118,N_29063);
nand U29212 (N_29212,N_29160,N_29122);
xnor U29213 (N_29213,N_29032,N_29124);
nand U29214 (N_29214,N_29074,N_29018);
nor U29215 (N_29215,N_29056,N_29129);
and U29216 (N_29216,N_29171,N_29059);
xnor U29217 (N_29217,N_29187,N_29035);
and U29218 (N_29218,N_29128,N_29095);
and U29219 (N_29219,N_29081,N_29180);
xnor U29220 (N_29220,N_29072,N_29136);
nand U29221 (N_29221,N_29065,N_29120);
nand U29222 (N_29222,N_29179,N_29026);
xor U29223 (N_29223,N_29046,N_29042);
nand U29224 (N_29224,N_29104,N_29139);
nor U29225 (N_29225,N_29084,N_29027);
xor U29226 (N_29226,N_29001,N_29051);
or U29227 (N_29227,N_29033,N_29005);
nand U29228 (N_29228,N_29143,N_29111);
xnor U29229 (N_29229,N_29015,N_29182);
nand U29230 (N_29230,N_29024,N_29135);
and U29231 (N_29231,N_29163,N_29197);
and U29232 (N_29232,N_29186,N_29195);
nor U29233 (N_29233,N_29130,N_29004);
or U29234 (N_29234,N_29048,N_29127);
and U29235 (N_29235,N_29061,N_29181);
and U29236 (N_29236,N_29031,N_29184);
and U29237 (N_29237,N_29087,N_29100);
or U29238 (N_29238,N_29038,N_29183);
xnor U29239 (N_29239,N_29088,N_29052);
xor U29240 (N_29240,N_29002,N_29091);
and U29241 (N_29241,N_29144,N_29079);
or U29242 (N_29242,N_29037,N_29071);
xor U29243 (N_29243,N_29082,N_29199);
nand U29244 (N_29244,N_29117,N_29198);
nor U29245 (N_29245,N_29062,N_29113);
or U29246 (N_29246,N_29034,N_29140);
xor U29247 (N_29247,N_29092,N_29064);
nor U29248 (N_29248,N_29151,N_29022);
xor U29249 (N_29249,N_29194,N_29150);
xor U29250 (N_29250,N_29189,N_29073);
or U29251 (N_29251,N_29029,N_29112);
and U29252 (N_29252,N_29177,N_29191);
or U29253 (N_29253,N_29017,N_29185);
and U29254 (N_29254,N_29009,N_29093);
and U29255 (N_29255,N_29049,N_29154);
xnor U29256 (N_29256,N_29133,N_29134);
nor U29257 (N_29257,N_29045,N_29178);
nor U29258 (N_29258,N_29192,N_29020);
nor U29259 (N_29259,N_29090,N_29141);
nand U29260 (N_29260,N_29013,N_29021);
xnor U29261 (N_29261,N_29016,N_29053);
or U29262 (N_29262,N_29066,N_29054);
xnor U29263 (N_29263,N_29132,N_29010);
nand U29264 (N_29264,N_29176,N_29159);
nor U29265 (N_29265,N_29055,N_29157);
nor U29266 (N_29266,N_29025,N_29105);
nand U29267 (N_29267,N_29070,N_29023);
or U29268 (N_29268,N_29152,N_29039);
xor U29269 (N_29269,N_29030,N_29036);
or U29270 (N_29270,N_29050,N_29014);
nand U29271 (N_29271,N_29109,N_29097);
nor U29272 (N_29272,N_29115,N_29193);
xor U29273 (N_29273,N_29047,N_29137);
nor U29274 (N_29274,N_29123,N_29138);
nor U29275 (N_29275,N_29078,N_29101);
nor U29276 (N_29276,N_29076,N_29110);
nand U29277 (N_29277,N_29147,N_29188);
or U29278 (N_29278,N_29057,N_29106);
and U29279 (N_29279,N_29162,N_29169);
nand U29280 (N_29280,N_29044,N_29156);
and U29281 (N_29281,N_29099,N_29196);
nand U29282 (N_29282,N_29119,N_29173);
nand U29283 (N_29283,N_29190,N_29094);
nor U29284 (N_29284,N_29058,N_29019);
xnor U29285 (N_29285,N_29103,N_29168);
xnor U29286 (N_29286,N_29166,N_29175);
xor U29287 (N_29287,N_29067,N_29126);
xnor U29288 (N_29288,N_29043,N_29085);
or U29289 (N_29289,N_29003,N_29116);
or U29290 (N_29290,N_29158,N_29008);
nor U29291 (N_29291,N_29170,N_29148);
or U29292 (N_29292,N_29172,N_29000);
or U29293 (N_29293,N_29167,N_29069);
nor U29294 (N_29294,N_29060,N_29149);
or U29295 (N_29295,N_29155,N_29089);
or U29296 (N_29296,N_29080,N_29164);
or U29297 (N_29297,N_29041,N_29145);
xnor U29298 (N_29298,N_29007,N_29153);
and U29299 (N_29299,N_29012,N_29006);
nand U29300 (N_29300,N_29131,N_29038);
nor U29301 (N_29301,N_29197,N_29193);
or U29302 (N_29302,N_29142,N_29020);
or U29303 (N_29303,N_29166,N_29077);
or U29304 (N_29304,N_29055,N_29020);
nor U29305 (N_29305,N_29171,N_29120);
xnor U29306 (N_29306,N_29034,N_29151);
nor U29307 (N_29307,N_29187,N_29117);
nor U29308 (N_29308,N_29154,N_29040);
xnor U29309 (N_29309,N_29115,N_29042);
and U29310 (N_29310,N_29010,N_29083);
nor U29311 (N_29311,N_29101,N_29136);
or U29312 (N_29312,N_29137,N_29100);
and U29313 (N_29313,N_29197,N_29099);
and U29314 (N_29314,N_29025,N_29155);
and U29315 (N_29315,N_29129,N_29094);
nor U29316 (N_29316,N_29142,N_29041);
xnor U29317 (N_29317,N_29000,N_29135);
xnor U29318 (N_29318,N_29119,N_29074);
nor U29319 (N_29319,N_29195,N_29153);
or U29320 (N_29320,N_29013,N_29138);
or U29321 (N_29321,N_29032,N_29085);
nand U29322 (N_29322,N_29159,N_29014);
or U29323 (N_29323,N_29103,N_29004);
and U29324 (N_29324,N_29017,N_29074);
xor U29325 (N_29325,N_29189,N_29025);
or U29326 (N_29326,N_29171,N_29051);
or U29327 (N_29327,N_29187,N_29014);
or U29328 (N_29328,N_29137,N_29114);
and U29329 (N_29329,N_29197,N_29192);
and U29330 (N_29330,N_29116,N_29168);
nand U29331 (N_29331,N_29036,N_29047);
nand U29332 (N_29332,N_29112,N_29094);
xnor U29333 (N_29333,N_29192,N_29111);
or U29334 (N_29334,N_29023,N_29042);
nand U29335 (N_29335,N_29049,N_29100);
nor U29336 (N_29336,N_29139,N_29178);
or U29337 (N_29337,N_29077,N_29081);
or U29338 (N_29338,N_29144,N_29037);
and U29339 (N_29339,N_29084,N_29119);
nand U29340 (N_29340,N_29108,N_29103);
and U29341 (N_29341,N_29069,N_29010);
nand U29342 (N_29342,N_29192,N_29028);
and U29343 (N_29343,N_29120,N_29134);
and U29344 (N_29344,N_29141,N_29059);
nor U29345 (N_29345,N_29004,N_29115);
and U29346 (N_29346,N_29021,N_29082);
nor U29347 (N_29347,N_29033,N_29181);
or U29348 (N_29348,N_29166,N_29048);
nand U29349 (N_29349,N_29097,N_29082);
nand U29350 (N_29350,N_29012,N_29139);
or U29351 (N_29351,N_29197,N_29037);
nor U29352 (N_29352,N_29091,N_29086);
or U29353 (N_29353,N_29105,N_29052);
nor U29354 (N_29354,N_29116,N_29155);
and U29355 (N_29355,N_29082,N_29018);
or U29356 (N_29356,N_29021,N_29055);
xnor U29357 (N_29357,N_29158,N_29193);
nor U29358 (N_29358,N_29074,N_29031);
or U29359 (N_29359,N_29143,N_29068);
nand U29360 (N_29360,N_29193,N_29024);
nand U29361 (N_29361,N_29001,N_29161);
nor U29362 (N_29362,N_29156,N_29019);
xor U29363 (N_29363,N_29058,N_29142);
nand U29364 (N_29364,N_29196,N_29180);
or U29365 (N_29365,N_29199,N_29100);
xnor U29366 (N_29366,N_29006,N_29034);
and U29367 (N_29367,N_29131,N_29188);
or U29368 (N_29368,N_29112,N_29076);
nor U29369 (N_29369,N_29163,N_29011);
nor U29370 (N_29370,N_29009,N_29187);
and U29371 (N_29371,N_29116,N_29152);
xnor U29372 (N_29372,N_29066,N_29117);
or U29373 (N_29373,N_29058,N_29092);
nand U29374 (N_29374,N_29029,N_29103);
nor U29375 (N_29375,N_29123,N_29007);
or U29376 (N_29376,N_29161,N_29158);
xor U29377 (N_29377,N_29155,N_29017);
or U29378 (N_29378,N_29090,N_29020);
nor U29379 (N_29379,N_29053,N_29038);
xor U29380 (N_29380,N_29132,N_29085);
and U29381 (N_29381,N_29100,N_29017);
nand U29382 (N_29382,N_29049,N_29093);
and U29383 (N_29383,N_29043,N_29083);
nand U29384 (N_29384,N_29144,N_29182);
nand U29385 (N_29385,N_29138,N_29037);
xor U29386 (N_29386,N_29099,N_29146);
and U29387 (N_29387,N_29142,N_29088);
nor U29388 (N_29388,N_29004,N_29090);
xnor U29389 (N_29389,N_29175,N_29172);
nand U29390 (N_29390,N_29045,N_29157);
nor U29391 (N_29391,N_29126,N_29033);
nor U29392 (N_29392,N_29077,N_29046);
and U29393 (N_29393,N_29113,N_29027);
and U29394 (N_29394,N_29130,N_29072);
xor U29395 (N_29395,N_29197,N_29109);
nor U29396 (N_29396,N_29045,N_29148);
nand U29397 (N_29397,N_29179,N_29029);
xnor U29398 (N_29398,N_29199,N_29079);
or U29399 (N_29399,N_29163,N_29175);
nor U29400 (N_29400,N_29265,N_29302);
xor U29401 (N_29401,N_29370,N_29262);
xor U29402 (N_29402,N_29327,N_29398);
or U29403 (N_29403,N_29392,N_29359);
nor U29404 (N_29404,N_29349,N_29279);
xnor U29405 (N_29405,N_29323,N_29283);
and U29406 (N_29406,N_29223,N_29291);
nor U29407 (N_29407,N_29368,N_29271);
and U29408 (N_29408,N_29273,N_29364);
nor U29409 (N_29409,N_29236,N_29288);
nand U29410 (N_29410,N_29284,N_29313);
and U29411 (N_29411,N_29232,N_29237);
and U29412 (N_29412,N_29325,N_29391);
nand U29413 (N_29413,N_29310,N_29258);
and U29414 (N_29414,N_29299,N_29255);
xor U29415 (N_29415,N_29275,N_29251);
nand U29416 (N_29416,N_29296,N_29252);
and U29417 (N_29417,N_29340,N_29214);
xor U29418 (N_29418,N_29231,N_29375);
nand U29419 (N_29419,N_29385,N_29295);
nor U29420 (N_29420,N_29300,N_29307);
and U29421 (N_29421,N_29344,N_29361);
nor U29422 (N_29422,N_29347,N_29355);
and U29423 (N_29423,N_29297,N_29233);
xnor U29424 (N_29424,N_29358,N_29380);
xnor U29425 (N_29425,N_29376,N_29207);
and U29426 (N_29426,N_29204,N_29274);
or U29427 (N_29427,N_29248,N_29387);
or U29428 (N_29428,N_29206,N_29253);
and U29429 (N_29429,N_29256,N_29215);
nand U29430 (N_29430,N_29239,N_29245);
or U29431 (N_29431,N_29338,N_29238);
or U29432 (N_29432,N_29241,N_29303);
or U29433 (N_29433,N_29203,N_29377);
nor U29434 (N_29434,N_29286,N_29316);
or U29435 (N_29435,N_29229,N_29278);
and U29436 (N_29436,N_29335,N_29315);
nor U29437 (N_29437,N_29319,N_29244);
or U29438 (N_29438,N_29201,N_29314);
and U29439 (N_29439,N_29209,N_29343);
and U29440 (N_29440,N_29342,N_29285);
or U29441 (N_29441,N_29366,N_29381);
nor U29442 (N_29442,N_29269,N_29351);
nor U29443 (N_29443,N_29280,N_29333);
nor U29444 (N_29444,N_29304,N_29257);
xnor U29445 (N_29445,N_29369,N_29270);
or U29446 (N_29446,N_29200,N_29260);
or U29447 (N_29447,N_29308,N_29242);
xnor U29448 (N_29448,N_29261,N_29390);
nand U29449 (N_29449,N_29254,N_29220);
and U29450 (N_29450,N_29395,N_29217);
and U29451 (N_29451,N_29216,N_29287);
xor U29452 (N_29452,N_29332,N_29218);
xor U29453 (N_29453,N_29331,N_29305);
and U29454 (N_29454,N_29277,N_29240);
or U29455 (N_29455,N_29328,N_29399);
xor U29456 (N_29456,N_29379,N_29378);
nand U29457 (N_29457,N_29309,N_29234);
xnor U29458 (N_29458,N_29324,N_29329);
nand U29459 (N_29459,N_29290,N_29318);
nand U29460 (N_29460,N_29228,N_29371);
xnor U29461 (N_29461,N_29341,N_29263);
nand U29462 (N_29462,N_29357,N_29336);
nand U29463 (N_29463,N_29219,N_29330);
nand U29464 (N_29464,N_29334,N_29363);
nand U29465 (N_29465,N_29348,N_29243);
nand U29466 (N_29466,N_29282,N_29339);
xnor U29467 (N_29467,N_29235,N_29322);
nand U29468 (N_29468,N_29221,N_29373);
xor U29469 (N_29469,N_29227,N_29360);
xnor U29470 (N_29470,N_29394,N_29292);
and U29471 (N_29471,N_29320,N_29211);
xor U29472 (N_29472,N_29393,N_29312);
and U29473 (N_29473,N_29213,N_29202);
nor U29474 (N_29474,N_29362,N_29293);
and U29475 (N_29475,N_29208,N_29298);
nand U29476 (N_29476,N_29301,N_29225);
or U29477 (N_29477,N_29388,N_29326);
and U29478 (N_29478,N_29383,N_29281);
nand U29479 (N_29479,N_29397,N_29212);
and U29480 (N_29480,N_29345,N_29250);
or U29481 (N_29481,N_29382,N_29311);
and U29482 (N_29482,N_29294,N_29224);
nor U29483 (N_29483,N_29396,N_29365);
and U29484 (N_29484,N_29354,N_29367);
nand U29485 (N_29485,N_29317,N_29306);
xnor U29486 (N_29486,N_29353,N_29352);
xor U29487 (N_29487,N_29374,N_29350);
xnor U29488 (N_29488,N_29222,N_29346);
xnor U29489 (N_29489,N_29356,N_29372);
and U29490 (N_29490,N_29264,N_29321);
or U29491 (N_29491,N_29267,N_29266);
or U29492 (N_29492,N_29259,N_29276);
nand U29493 (N_29493,N_29210,N_29389);
nor U29494 (N_29494,N_29246,N_29289);
and U29495 (N_29495,N_29272,N_29205);
or U29496 (N_29496,N_29268,N_29386);
xnor U29497 (N_29497,N_29337,N_29226);
xor U29498 (N_29498,N_29384,N_29249);
or U29499 (N_29499,N_29247,N_29230);
or U29500 (N_29500,N_29259,N_29290);
or U29501 (N_29501,N_29393,N_29372);
nand U29502 (N_29502,N_29307,N_29250);
or U29503 (N_29503,N_29238,N_29208);
nor U29504 (N_29504,N_29212,N_29386);
nand U29505 (N_29505,N_29201,N_29329);
nor U29506 (N_29506,N_29379,N_29361);
nand U29507 (N_29507,N_29312,N_29293);
xor U29508 (N_29508,N_29279,N_29372);
or U29509 (N_29509,N_29339,N_29314);
xor U29510 (N_29510,N_29300,N_29382);
and U29511 (N_29511,N_29319,N_29206);
and U29512 (N_29512,N_29231,N_29346);
or U29513 (N_29513,N_29285,N_29205);
xnor U29514 (N_29514,N_29333,N_29249);
or U29515 (N_29515,N_29253,N_29378);
nor U29516 (N_29516,N_29301,N_29251);
nor U29517 (N_29517,N_29289,N_29298);
nor U29518 (N_29518,N_29387,N_29200);
and U29519 (N_29519,N_29316,N_29308);
and U29520 (N_29520,N_29357,N_29264);
xnor U29521 (N_29521,N_29290,N_29224);
nand U29522 (N_29522,N_29324,N_29214);
and U29523 (N_29523,N_29230,N_29246);
nand U29524 (N_29524,N_29251,N_29206);
or U29525 (N_29525,N_29391,N_29289);
nor U29526 (N_29526,N_29248,N_29212);
nand U29527 (N_29527,N_29229,N_29238);
or U29528 (N_29528,N_29291,N_29220);
xnor U29529 (N_29529,N_29207,N_29306);
xnor U29530 (N_29530,N_29337,N_29259);
nand U29531 (N_29531,N_29255,N_29327);
nor U29532 (N_29532,N_29272,N_29341);
xnor U29533 (N_29533,N_29360,N_29394);
nor U29534 (N_29534,N_29375,N_29309);
nor U29535 (N_29535,N_29223,N_29210);
xor U29536 (N_29536,N_29276,N_29201);
nor U29537 (N_29537,N_29261,N_29392);
nor U29538 (N_29538,N_29313,N_29211);
and U29539 (N_29539,N_29315,N_29361);
nand U29540 (N_29540,N_29276,N_29274);
and U29541 (N_29541,N_29342,N_29266);
or U29542 (N_29542,N_29226,N_29343);
xnor U29543 (N_29543,N_29359,N_29362);
or U29544 (N_29544,N_29217,N_29255);
nor U29545 (N_29545,N_29320,N_29398);
xor U29546 (N_29546,N_29328,N_29294);
nand U29547 (N_29547,N_29273,N_29258);
nand U29548 (N_29548,N_29370,N_29256);
nor U29549 (N_29549,N_29223,N_29251);
xor U29550 (N_29550,N_29319,N_29235);
and U29551 (N_29551,N_29316,N_29292);
xor U29552 (N_29552,N_29289,N_29373);
xnor U29553 (N_29553,N_29318,N_29257);
and U29554 (N_29554,N_29344,N_29302);
or U29555 (N_29555,N_29362,N_29308);
nor U29556 (N_29556,N_29232,N_29219);
nand U29557 (N_29557,N_29346,N_29294);
nor U29558 (N_29558,N_29227,N_29398);
nor U29559 (N_29559,N_29210,N_29305);
nor U29560 (N_29560,N_29216,N_29242);
nor U29561 (N_29561,N_29243,N_29324);
xor U29562 (N_29562,N_29204,N_29285);
and U29563 (N_29563,N_29289,N_29307);
nand U29564 (N_29564,N_29296,N_29289);
nand U29565 (N_29565,N_29339,N_29245);
xnor U29566 (N_29566,N_29388,N_29349);
xor U29567 (N_29567,N_29234,N_29397);
nor U29568 (N_29568,N_29286,N_29306);
xnor U29569 (N_29569,N_29361,N_29360);
and U29570 (N_29570,N_29383,N_29392);
nor U29571 (N_29571,N_29285,N_29220);
xnor U29572 (N_29572,N_29256,N_29280);
and U29573 (N_29573,N_29332,N_29304);
xnor U29574 (N_29574,N_29337,N_29294);
nor U29575 (N_29575,N_29208,N_29306);
or U29576 (N_29576,N_29358,N_29365);
or U29577 (N_29577,N_29368,N_29373);
nand U29578 (N_29578,N_29283,N_29388);
nand U29579 (N_29579,N_29230,N_29251);
nor U29580 (N_29580,N_29380,N_29363);
and U29581 (N_29581,N_29234,N_29271);
nor U29582 (N_29582,N_29333,N_29339);
xor U29583 (N_29583,N_29381,N_29382);
xor U29584 (N_29584,N_29202,N_29394);
nand U29585 (N_29585,N_29384,N_29382);
nor U29586 (N_29586,N_29339,N_29338);
nand U29587 (N_29587,N_29227,N_29201);
and U29588 (N_29588,N_29228,N_29314);
nor U29589 (N_29589,N_29396,N_29364);
or U29590 (N_29590,N_29206,N_29371);
or U29591 (N_29591,N_29299,N_29353);
or U29592 (N_29592,N_29366,N_29203);
nor U29593 (N_29593,N_29365,N_29341);
nor U29594 (N_29594,N_29309,N_29238);
nand U29595 (N_29595,N_29259,N_29346);
or U29596 (N_29596,N_29260,N_29214);
or U29597 (N_29597,N_29208,N_29258);
nor U29598 (N_29598,N_29265,N_29330);
nor U29599 (N_29599,N_29238,N_29397);
or U29600 (N_29600,N_29524,N_29407);
and U29601 (N_29601,N_29469,N_29413);
nand U29602 (N_29602,N_29426,N_29519);
or U29603 (N_29603,N_29548,N_29567);
nor U29604 (N_29604,N_29557,N_29569);
xor U29605 (N_29605,N_29513,N_29423);
and U29606 (N_29606,N_29565,N_29539);
and U29607 (N_29607,N_29492,N_29574);
xnor U29608 (N_29608,N_29401,N_29405);
nand U29609 (N_29609,N_29562,N_29590);
or U29610 (N_29610,N_29585,N_29502);
or U29611 (N_29611,N_29532,N_29444);
xor U29612 (N_29612,N_29463,N_29435);
and U29613 (N_29613,N_29579,N_29566);
nor U29614 (N_29614,N_29408,N_29589);
nor U29615 (N_29615,N_29410,N_29448);
xor U29616 (N_29616,N_29450,N_29593);
nor U29617 (N_29617,N_29558,N_29555);
nand U29618 (N_29618,N_29531,N_29545);
and U29619 (N_29619,N_29456,N_29577);
nor U29620 (N_29620,N_29588,N_29507);
or U29621 (N_29621,N_29442,N_29505);
nor U29622 (N_29622,N_29521,N_29454);
nand U29623 (N_29623,N_29535,N_29592);
nand U29624 (N_29624,N_29495,N_29510);
and U29625 (N_29625,N_29475,N_29420);
xnor U29626 (N_29626,N_29432,N_29561);
and U29627 (N_29627,N_29533,N_29525);
xnor U29628 (N_29628,N_29440,N_29549);
nand U29629 (N_29629,N_29596,N_29512);
nand U29630 (N_29630,N_29580,N_29459);
nor U29631 (N_29631,N_29404,N_29493);
and U29632 (N_29632,N_29526,N_29508);
or U29633 (N_29633,N_29418,N_29527);
xor U29634 (N_29634,N_29546,N_29416);
or U29635 (N_29635,N_29434,N_29570);
xor U29636 (N_29636,N_29449,N_29427);
and U29637 (N_29637,N_29455,N_29514);
xor U29638 (N_29638,N_29551,N_29537);
xnor U29639 (N_29639,N_29443,N_29554);
nor U29640 (N_29640,N_29458,N_29522);
and U29641 (N_29641,N_29598,N_29485);
or U29642 (N_29642,N_29576,N_29529);
and U29643 (N_29643,N_29412,N_29453);
xnor U29644 (N_29644,N_29451,N_29536);
nand U29645 (N_29645,N_29501,N_29544);
and U29646 (N_29646,N_29494,N_29528);
nor U29647 (N_29647,N_29564,N_29597);
xor U29648 (N_29648,N_29511,N_29452);
and U29649 (N_29649,N_29474,N_29419);
and U29650 (N_29650,N_29406,N_29473);
nor U29651 (N_29651,N_29484,N_29468);
nor U29652 (N_29652,N_29515,N_29403);
and U29653 (N_29653,N_29509,N_29472);
nand U29654 (N_29654,N_29461,N_29595);
or U29655 (N_29655,N_29490,N_29457);
and U29656 (N_29656,N_29563,N_29479);
xnor U29657 (N_29657,N_29431,N_29424);
nand U29658 (N_29658,N_29488,N_29542);
or U29659 (N_29659,N_29552,N_29486);
or U29660 (N_29660,N_29599,N_29568);
nor U29661 (N_29661,N_29543,N_29587);
or U29662 (N_29662,N_29430,N_29517);
and U29663 (N_29663,N_29584,N_29591);
nand U29664 (N_29664,N_29421,N_29433);
xor U29665 (N_29665,N_29460,N_29429);
nand U29666 (N_29666,N_29446,N_29439);
xnor U29667 (N_29667,N_29541,N_29578);
or U29668 (N_29668,N_29425,N_29445);
nand U29669 (N_29669,N_29491,N_29550);
and U29670 (N_29670,N_29471,N_29523);
nor U29671 (N_29671,N_29470,N_29506);
nand U29672 (N_29672,N_29573,N_29498);
or U29673 (N_29673,N_29441,N_29503);
nor U29674 (N_29674,N_29594,N_29547);
xor U29675 (N_29675,N_29560,N_29556);
nor U29676 (N_29676,N_29571,N_29559);
or U29677 (N_29677,N_29496,N_29583);
and U29678 (N_29678,N_29518,N_29582);
nand U29679 (N_29679,N_29417,N_29428);
nand U29680 (N_29680,N_29516,N_29520);
nand U29681 (N_29681,N_29500,N_29553);
or U29682 (N_29682,N_29447,N_29482);
or U29683 (N_29683,N_29415,N_29497);
or U29684 (N_29684,N_29422,N_29572);
and U29685 (N_29685,N_29478,N_29436);
xnor U29686 (N_29686,N_29462,N_29487);
xor U29687 (N_29687,N_29409,N_29530);
or U29688 (N_29688,N_29402,N_29534);
or U29689 (N_29689,N_29400,N_29489);
or U29690 (N_29690,N_29581,N_29476);
nand U29691 (N_29691,N_29540,N_29504);
nand U29692 (N_29692,N_29538,N_29477);
or U29693 (N_29693,N_29466,N_29480);
or U29694 (N_29694,N_29586,N_29483);
nor U29695 (N_29695,N_29437,N_29481);
nor U29696 (N_29696,N_29438,N_29499);
nand U29697 (N_29697,N_29464,N_29465);
or U29698 (N_29698,N_29411,N_29414);
or U29699 (N_29699,N_29467,N_29575);
xor U29700 (N_29700,N_29474,N_29412);
or U29701 (N_29701,N_29565,N_29400);
and U29702 (N_29702,N_29472,N_29427);
nor U29703 (N_29703,N_29499,N_29475);
nand U29704 (N_29704,N_29414,N_29454);
nand U29705 (N_29705,N_29548,N_29489);
nor U29706 (N_29706,N_29527,N_29589);
xor U29707 (N_29707,N_29416,N_29497);
nor U29708 (N_29708,N_29556,N_29506);
or U29709 (N_29709,N_29459,N_29432);
xnor U29710 (N_29710,N_29518,N_29451);
and U29711 (N_29711,N_29553,N_29538);
xor U29712 (N_29712,N_29487,N_29573);
nand U29713 (N_29713,N_29468,N_29531);
nand U29714 (N_29714,N_29404,N_29520);
or U29715 (N_29715,N_29485,N_29495);
and U29716 (N_29716,N_29597,N_29459);
or U29717 (N_29717,N_29476,N_29520);
nor U29718 (N_29718,N_29577,N_29400);
and U29719 (N_29719,N_29515,N_29461);
and U29720 (N_29720,N_29456,N_29581);
nand U29721 (N_29721,N_29486,N_29558);
and U29722 (N_29722,N_29507,N_29583);
nor U29723 (N_29723,N_29526,N_29473);
xnor U29724 (N_29724,N_29503,N_29571);
nand U29725 (N_29725,N_29496,N_29486);
xor U29726 (N_29726,N_29593,N_29423);
and U29727 (N_29727,N_29488,N_29529);
xnor U29728 (N_29728,N_29532,N_29433);
and U29729 (N_29729,N_29494,N_29573);
xnor U29730 (N_29730,N_29466,N_29405);
nor U29731 (N_29731,N_29416,N_29412);
nand U29732 (N_29732,N_29503,N_29582);
and U29733 (N_29733,N_29492,N_29420);
xor U29734 (N_29734,N_29484,N_29496);
xnor U29735 (N_29735,N_29483,N_29577);
xor U29736 (N_29736,N_29564,N_29470);
and U29737 (N_29737,N_29536,N_29590);
or U29738 (N_29738,N_29539,N_29543);
and U29739 (N_29739,N_29557,N_29407);
nor U29740 (N_29740,N_29557,N_29564);
nand U29741 (N_29741,N_29598,N_29592);
xnor U29742 (N_29742,N_29434,N_29514);
xnor U29743 (N_29743,N_29425,N_29484);
and U29744 (N_29744,N_29487,N_29437);
nor U29745 (N_29745,N_29468,N_29578);
xnor U29746 (N_29746,N_29477,N_29401);
nor U29747 (N_29747,N_29434,N_29492);
xor U29748 (N_29748,N_29443,N_29515);
nand U29749 (N_29749,N_29490,N_29472);
nand U29750 (N_29750,N_29486,N_29523);
or U29751 (N_29751,N_29513,N_29551);
and U29752 (N_29752,N_29581,N_29596);
nor U29753 (N_29753,N_29500,N_29512);
and U29754 (N_29754,N_29406,N_29420);
or U29755 (N_29755,N_29406,N_29408);
or U29756 (N_29756,N_29558,N_29525);
or U29757 (N_29757,N_29467,N_29481);
nor U29758 (N_29758,N_29402,N_29406);
nand U29759 (N_29759,N_29559,N_29580);
nor U29760 (N_29760,N_29470,N_29532);
xor U29761 (N_29761,N_29472,N_29453);
xor U29762 (N_29762,N_29466,N_29524);
nor U29763 (N_29763,N_29486,N_29505);
and U29764 (N_29764,N_29541,N_29576);
and U29765 (N_29765,N_29403,N_29542);
xor U29766 (N_29766,N_29558,N_29485);
nand U29767 (N_29767,N_29536,N_29492);
or U29768 (N_29768,N_29442,N_29509);
nor U29769 (N_29769,N_29550,N_29523);
or U29770 (N_29770,N_29449,N_29597);
nand U29771 (N_29771,N_29556,N_29554);
xor U29772 (N_29772,N_29554,N_29435);
nand U29773 (N_29773,N_29400,N_29551);
nand U29774 (N_29774,N_29474,N_29596);
xnor U29775 (N_29775,N_29426,N_29474);
nand U29776 (N_29776,N_29577,N_29448);
nor U29777 (N_29777,N_29596,N_29410);
xnor U29778 (N_29778,N_29485,N_29454);
or U29779 (N_29779,N_29459,N_29538);
nor U29780 (N_29780,N_29570,N_29522);
or U29781 (N_29781,N_29584,N_29462);
xnor U29782 (N_29782,N_29490,N_29598);
or U29783 (N_29783,N_29493,N_29424);
nand U29784 (N_29784,N_29583,N_29517);
xor U29785 (N_29785,N_29592,N_29434);
xor U29786 (N_29786,N_29473,N_29590);
or U29787 (N_29787,N_29489,N_29561);
xor U29788 (N_29788,N_29555,N_29412);
xnor U29789 (N_29789,N_29489,N_29533);
nand U29790 (N_29790,N_29423,N_29567);
xor U29791 (N_29791,N_29470,N_29553);
nor U29792 (N_29792,N_29577,N_29432);
or U29793 (N_29793,N_29597,N_29518);
or U29794 (N_29794,N_29480,N_29412);
xnor U29795 (N_29795,N_29567,N_29554);
nand U29796 (N_29796,N_29475,N_29450);
xor U29797 (N_29797,N_29413,N_29484);
and U29798 (N_29798,N_29479,N_29577);
or U29799 (N_29799,N_29453,N_29546);
and U29800 (N_29800,N_29690,N_29786);
xnor U29801 (N_29801,N_29671,N_29687);
nor U29802 (N_29802,N_29792,N_29732);
nor U29803 (N_29803,N_29753,N_29625);
nand U29804 (N_29804,N_29617,N_29610);
nand U29805 (N_29805,N_29787,N_29730);
or U29806 (N_29806,N_29710,N_29655);
xnor U29807 (N_29807,N_29632,N_29760);
xnor U29808 (N_29808,N_29627,N_29776);
and U29809 (N_29809,N_29676,N_29620);
and U29810 (N_29810,N_29759,N_29640);
nand U29811 (N_29811,N_29612,N_29737);
nand U29812 (N_29812,N_29649,N_29782);
or U29813 (N_29813,N_29635,N_29750);
xor U29814 (N_29814,N_29720,N_29734);
nor U29815 (N_29815,N_29684,N_29660);
nand U29816 (N_29816,N_29774,N_29773);
nor U29817 (N_29817,N_29794,N_29658);
and U29818 (N_29818,N_29719,N_29670);
and U29819 (N_29819,N_29765,N_29609);
nand U29820 (N_29820,N_29745,N_29700);
and U29821 (N_29821,N_29642,N_29704);
and U29822 (N_29822,N_29613,N_29699);
nor U29823 (N_29823,N_29761,N_29716);
or U29824 (N_29824,N_29736,N_29702);
or U29825 (N_29825,N_29769,N_29742);
xor U29826 (N_29826,N_29752,N_29672);
xnor U29827 (N_29827,N_29758,N_29789);
or U29828 (N_29828,N_29603,N_29638);
and U29829 (N_29829,N_29731,N_29729);
xnor U29830 (N_29830,N_29735,N_29641);
nor U29831 (N_29831,N_29784,N_29696);
or U29832 (N_29832,N_29673,N_29726);
nand U29833 (N_29833,N_29712,N_29659);
nor U29834 (N_29834,N_29739,N_29775);
and U29835 (N_29835,N_29706,N_29652);
xnor U29836 (N_29836,N_29683,N_29631);
nor U29837 (N_29837,N_29654,N_29755);
nand U29838 (N_29838,N_29777,N_29644);
nand U29839 (N_29839,N_29727,N_29779);
or U29840 (N_29840,N_29615,N_29692);
nor U29841 (N_29841,N_29778,N_29698);
nand U29842 (N_29842,N_29667,N_29767);
or U29843 (N_29843,N_29661,N_29682);
nand U29844 (N_29844,N_29703,N_29733);
nor U29845 (N_29845,N_29708,N_29633);
xor U29846 (N_29846,N_29677,N_29743);
nor U29847 (N_29847,N_29600,N_29653);
and U29848 (N_29848,N_29715,N_29711);
or U29849 (N_29849,N_29685,N_29645);
nor U29850 (N_29850,N_29689,N_29694);
nand U29851 (N_29851,N_29669,N_29668);
and U29852 (N_29852,N_29681,N_29747);
xnor U29853 (N_29853,N_29738,N_29717);
or U29854 (N_29854,N_29772,N_29788);
and U29855 (N_29855,N_29764,N_29662);
xnor U29856 (N_29856,N_29666,N_29763);
and U29857 (N_29857,N_29780,N_29626);
xnor U29858 (N_29858,N_29607,N_29746);
and U29859 (N_29859,N_29680,N_29608);
xor U29860 (N_29860,N_29714,N_29605);
nor U29861 (N_29861,N_29756,N_29639);
nor U29862 (N_29862,N_29770,N_29749);
nand U29863 (N_29863,N_29709,N_29618);
xnor U29864 (N_29864,N_29793,N_29637);
nor U29865 (N_29865,N_29674,N_29648);
and U29866 (N_29866,N_29604,N_29630);
nand U29867 (N_29867,N_29650,N_29705);
nand U29868 (N_29868,N_29728,N_29713);
and U29869 (N_29869,N_29724,N_29606);
and U29870 (N_29870,N_29790,N_29697);
or U29871 (N_29871,N_29781,N_29741);
and U29872 (N_29872,N_29688,N_29616);
xnor U29873 (N_29873,N_29665,N_29796);
and U29874 (N_29874,N_29799,N_29722);
nor U29875 (N_29875,N_29721,N_29622);
xor U29876 (N_29876,N_29766,N_29771);
and U29877 (N_29877,N_29646,N_29695);
or U29878 (N_29878,N_29701,N_29718);
nand U29879 (N_29879,N_29621,N_29611);
nand U29880 (N_29880,N_29628,N_29614);
and U29881 (N_29881,N_29623,N_29643);
and U29882 (N_29882,N_29744,N_29636);
and U29883 (N_29883,N_29785,N_29754);
nor U29884 (N_29884,N_29693,N_29691);
or U29885 (N_29885,N_29783,N_29678);
xnor U29886 (N_29886,N_29791,N_29725);
nand U29887 (N_29887,N_29634,N_29795);
xnor U29888 (N_29888,N_29762,N_29751);
xor U29889 (N_29889,N_29707,N_29602);
nand U29890 (N_29890,N_29601,N_29686);
xor U29891 (N_29891,N_29768,N_29651);
xor U29892 (N_29892,N_29748,N_29664);
xnor U29893 (N_29893,N_29757,N_29647);
xor U29894 (N_29894,N_29656,N_29619);
xor U29895 (N_29895,N_29797,N_29629);
nor U29896 (N_29896,N_29675,N_29663);
nand U29897 (N_29897,N_29740,N_29798);
nand U29898 (N_29898,N_29624,N_29679);
nand U29899 (N_29899,N_29657,N_29723);
and U29900 (N_29900,N_29784,N_29695);
and U29901 (N_29901,N_29685,N_29617);
xnor U29902 (N_29902,N_29733,N_29759);
or U29903 (N_29903,N_29633,N_29759);
xnor U29904 (N_29904,N_29687,N_29738);
or U29905 (N_29905,N_29729,N_29636);
xor U29906 (N_29906,N_29715,N_29624);
or U29907 (N_29907,N_29729,N_29609);
or U29908 (N_29908,N_29678,N_29701);
nand U29909 (N_29909,N_29662,N_29784);
and U29910 (N_29910,N_29783,N_29634);
or U29911 (N_29911,N_29796,N_29746);
or U29912 (N_29912,N_29692,N_29701);
xor U29913 (N_29913,N_29723,N_29663);
and U29914 (N_29914,N_29676,N_29648);
or U29915 (N_29915,N_29720,N_29782);
xnor U29916 (N_29916,N_29619,N_29760);
and U29917 (N_29917,N_29664,N_29726);
and U29918 (N_29918,N_29704,N_29760);
nand U29919 (N_29919,N_29672,N_29791);
nor U29920 (N_29920,N_29748,N_29770);
nand U29921 (N_29921,N_29721,N_29799);
nor U29922 (N_29922,N_29635,N_29606);
or U29923 (N_29923,N_29788,N_29769);
nand U29924 (N_29924,N_29630,N_29602);
xnor U29925 (N_29925,N_29706,N_29771);
or U29926 (N_29926,N_29659,N_29696);
xor U29927 (N_29927,N_29679,N_29628);
and U29928 (N_29928,N_29617,N_29604);
or U29929 (N_29929,N_29668,N_29731);
and U29930 (N_29930,N_29690,N_29612);
nor U29931 (N_29931,N_29682,N_29620);
and U29932 (N_29932,N_29639,N_29707);
xnor U29933 (N_29933,N_29666,N_29663);
nand U29934 (N_29934,N_29719,N_29612);
nor U29935 (N_29935,N_29773,N_29697);
or U29936 (N_29936,N_29612,N_29798);
xnor U29937 (N_29937,N_29786,N_29765);
or U29938 (N_29938,N_29724,N_29781);
xor U29939 (N_29939,N_29640,N_29620);
nand U29940 (N_29940,N_29693,N_29636);
or U29941 (N_29941,N_29764,N_29611);
xnor U29942 (N_29942,N_29633,N_29717);
nand U29943 (N_29943,N_29651,N_29790);
or U29944 (N_29944,N_29707,N_29664);
nand U29945 (N_29945,N_29622,N_29641);
xnor U29946 (N_29946,N_29707,N_29754);
and U29947 (N_29947,N_29646,N_29785);
and U29948 (N_29948,N_29767,N_29717);
nor U29949 (N_29949,N_29788,N_29694);
and U29950 (N_29950,N_29658,N_29696);
or U29951 (N_29951,N_29770,N_29703);
or U29952 (N_29952,N_29754,N_29602);
nor U29953 (N_29953,N_29704,N_29752);
nor U29954 (N_29954,N_29600,N_29640);
nor U29955 (N_29955,N_29704,N_29672);
or U29956 (N_29956,N_29732,N_29620);
nand U29957 (N_29957,N_29702,N_29796);
nor U29958 (N_29958,N_29682,N_29722);
and U29959 (N_29959,N_29701,N_29603);
nand U29960 (N_29960,N_29643,N_29609);
xor U29961 (N_29961,N_29666,N_29694);
nor U29962 (N_29962,N_29790,N_29721);
nand U29963 (N_29963,N_29772,N_29668);
xnor U29964 (N_29964,N_29778,N_29699);
or U29965 (N_29965,N_29607,N_29640);
or U29966 (N_29966,N_29732,N_29673);
nor U29967 (N_29967,N_29703,N_29767);
and U29968 (N_29968,N_29785,N_29799);
xor U29969 (N_29969,N_29642,N_29683);
nor U29970 (N_29970,N_29759,N_29637);
xnor U29971 (N_29971,N_29646,N_29735);
or U29972 (N_29972,N_29635,N_29794);
and U29973 (N_29973,N_29748,N_29734);
and U29974 (N_29974,N_29676,N_29763);
nand U29975 (N_29975,N_29637,N_29636);
and U29976 (N_29976,N_29700,N_29622);
or U29977 (N_29977,N_29656,N_29699);
nand U29978 (N_29978,N_29700,N_29786);
nor U29979 (N_29979,N_29650,N_29601);
and U29980 (N_29980,N_29650,N_29748);
and U29981 (N_29981,N_29624,N_29635);
xor U29982 (N_29982,N_29618,N_29799);
xor U29983 (N_29983,N_29783,N_29795);
nand U29984 (N_29984,N_29740,N_29674);
xnor U29985 (N_29985,N_29648,N_29754);
and U29986 (N_29986,N_29636,N_29767);
and U29987 (N_29987,N_29695,N_29715);
and U29988 (N_29988,N_29780,N_29695);
and U29989 (N_29989,N_29656,N_29705);
nor U29990 (N_29990,N_29645,N_29617);
xnor U29991 (N_29991,N_29794,N_29788);
and U29992 (N_29992,N_29644,N_29702);
and U29993 (N_29993,N_29772,N_29712);
and U29994 (N_29994,N_29630,N_29794);
nand U29995 (N_29995,N_29624,N_29746);
and U29996 (N_29996,N_29654,N_29723);
or U29997 (N_29997,N_29774,N_29640);
xor U29998 (N_29998,N_29776,N_29714);
xnor U29999 (N_29999,N_29604,N_29626);
xnor UO_0 (O_0,N_29967,N_29875);
nand UO_1 (O_1,N_29803,N_29914);
nand UO_2 (O_2,N_29992,N_29873);
and UO_3 (O_3,N_29852,N_29834);
and UO_4 (O_4,N_29923,N_29994);
nand UO_5 (O_5,N_29839,N_29940);
nand UO_6 (O_6,N_29897,N_29951);
or UO_7 (O_7,N_29856,N_29950);
or UO_8 (O_8,N_29814,N_29865);
nor UO_9 (O_9,N_29926,N_29809);
nand UO_10 (O_10,N_29905,N_29825);
xnor UO_11 (O_11,N_29882,N_29972);
nor UO_12 (O_12,N_29880,N_29954);
and UO_13 (O_13,N_29931,N_29981);
nand UO_14 (O_14,N_29812,N_29946);
nor UO_15 (O_15,N_29901,N_29878);
xnor UO_16 (O_16,N_29935,N_29840);
nor UO_17 (O_17,N_29986,N_29831);
nor UO_18 (O_18,N_29985,N_29947);
and UO_19 (O_19,N_29989,N_29820);
nand UO_20 (O_20,N_29888,N_29930);
xor UO_21 (O_21,N_29848,N_29917);
nand UO_22 (O_22,N_29970,N_29960);
nor UO_23 (O_23,N_29861,N_29958);
and UO_24 (O_24,N_29939,N_29998);
nor UO_25 (O_25,N_29889,N_29857);
xor UO_26 (O_26,N_29844,N_29904);
nor UO_27 (O_27,N_29934,N_29838);
and UO_28 (O_28,N_29973,N_29898);
xnor UO_29 (O_29,N_29872,N_29870);
and UO_30 (O_30,N_29948,N_29876);
nor UO_31 (O_31,N_29868,N_29822);
nor UO_32 (O_32,N_29910,N_29996);
or UO_33 (O_33,N_29842,N_29900);
and UO_34 (O_34,N_29828,N_29826);
and UO_35 (O_35,N_29936,N_29938);
and UO_36 (O_36,N_29881,N_29961);
or UO_37 (O_37,N_29995,N_29866);
or UO_38 (O_38,N_29885,N_29851);
xor UO_39 (O_39,N_29997,N_29903);
nor UO_40 (O_40,N_29832,N_29845);
and UO_41 (O_41,N_29999,N_29979);
or UO_42 (O_42,N_29993,N_29922);
xnor UO_43 (O_43,N_29815,N_29977);
and UO_44 (O_44,N_29827,N_29883);
nor UO_45 (O_45,N_29983,N_29806);
and UO_46 (O_46,N_29969,N_29855);
xnor UO_47 (O_47,N_29801,N_29821);
nor UO_48 (O_48,N_29974,N_29920);
or UO_49 (O_49,N_29982,N_29943);
and UO_50 (O_50,N_29886,N_29819);
nor UO_51 (O_51,N_29813,N_29836);
nor UO_52 (O_52,N_29800,N_29863);
xor UO_53 (O_53,N_29871,N_29833);
nand UO_54 (O_54,N_29975,N_29915);
and UO_55 (O_55,N_29906,N_29835);
or UO_56 (O_56,N_29879,N_29932);
nand UO_57 (O_57,N_29858,N_29808);
and UO_58 (O_58,N_29824,N_29908);
xnor UO_59 (O_59,N_29945,N_29823);
nand UO_60 (O_60,N_29916,N_29877);
nand UO_61 (O_61,N_29887,N_29942);
xnor UO_62 (O_62,N_29849,N_29850);
or UO_63 (O_63,N_29817,N_29918);
or UO_64 (O_64,N_29988,N_29971);
xnor UO_65 (O_65,N_29893,N_29937);
nor UO_66 (O_66,N_29927,N_29956);
and UO_67 (O_67,N_29978,N_29860);
nand UO_68 (O_68,N_29896,N_29909);
nor UO_69 (O_69,N_29966,N_29802);
nor UO_70 (O_70,N_29949,N_29955);
or UO_71 (O_71,N_29987,N_29843);
xnor UO_72 (O_72,N_29810,N_29874);
xnor UO_73 (O_73,N_29853,N_29913);
xnor UO_74 (O_74,N_29869,N_29990);
or UO_75 (O_75,N_29854,N_29864);
and UO_76 (O_76,N_29921,N_29894);
and UO_77 (O_77,N_29804,N_29964);
nand UO_78 (O_78,N_29980,N_29933);
nand UO_79 (O_79,N_29928,N_29907);
nor UO_80 (O_80,N_29902,N_29924);
or UO_81 (O_81,N_29811,N_29962);
or UO_82 (O_82,N_29968,N_29816);
nor UO_83 (O_83,N_29829,N_29859);
and UO_84 (O_84,N_29890,N_29884);
xor UO_85 (O_85,N_29965,N_29805);
xor UO_86 (O_86,N_29941,N_29867);
nor UO_87 (O_87,N_29976,N_29919);
xor UO_88 (O_88,N_29952,N_29841);
and UO_89 (O_89,N_29895,N_29912);
or UO_90 (O_90,N_29807,N_29984);
nand UO_91 (O_91,N_29891,N_29957);
and UO_92 (O_92,N_29991,N_29899);
nor UO_93 (O_93,N_29837,N_29892);
and UO_94 (O_94,N_29846,N_29911);
and UO_95 (O_95,N_29818,N_29929);
xnor UO_96 (O_96,N_29830,N_29862);
nor UO_97 (O_97,N_29953,N_29944);
and UO_98 (O_98,N_29959,N_29925);
nor UO_99 (O_99,N_29847,N_29963);
and UO_100 (O_100,N_29980,N_29898);
nand UO_101 (O_101,N_29823,N_29957);
nand UO_102 (O_102,N_29997,N_29801);
and UO_103 (O_103,N_29991,N_29828);
xnor UO_104 (O_104,N_29865,N_29902);
or UO_105 (O_105,N_29808,N_29826);
nor UO_106 (O_106,N_29836,N_29840);
xor UO_107 (O_107,N_29890,N_29926);
nand UO_108 (O_108,N_29845,N_29813);
nor UO_109 (O_109,N_29978,N_29843);
and UO_110 (O_110,N_29951,N_29914);
nor UO_111 (O_111,N_29908,N_29874);
nand UO_112 (O_112,N_29980,N_29882);
xnor UO_113 (O_113,N_29831,N_29881);
or UO_114 (O_114,N_29885,N_29998);
nor UO_115 (O_115,N_29838,N_29952);
nor UO_116 (O_116,N_29872,N_29809);
xnor UO_117 (O_117,N_29863,N_29873);
or UO_118 (O_118,N_29928,N_29834);
or UO_119 (O_119,N_29929,N_29985);
and UO_120 (O_120,N_29842,N_29836);
nand UO_121 (O_121,N_29818,N_29891);
nand UO_122 (O_122,N_29986,N_29828);
and UO_123 (O_123,N_29807,N_29879);
xnor UO_124 (O_124,N_29971,N_29806);
nor UO_125 (O_125,N_29886,N_29909);
xnor UO_126 (O_126,N_29918,N_29828);
and UO_127 (O_127,N_29888,N_29856);
nand UO_128 (O_128,N_29819,N_29989);
xnor UO_129 (O_129,N_29979,N_29900);
and UO_130 (O_130,N_29831,N_29930);
nor UO_131 (O_131,N_29973,N_29993);
or UO_132 (O_132,N_29848,N_29986);
xor UO_133 (O_133,N_29848,N_29915);
nand UO_134 (O_134,N_29871,N_29972);
nor UO_135 (O_135,N_29986,N_29990);
or UO_136 (O_136,N_29861,N_29825);
or UO_137 (O_137,N_29889,N_29887);
or UO_138 (O_138,N_29960,N_29988);
nor UO_139 (O_139,N_29819,N_29921);
xnor UO_140 (O_140,N_29967,N_29904);
and UO_141 (O_141,N_29822,N_29876);
or UO_142 (O_142,N_29911,N_29828);
xor UO_143 (O_143,N_29953,N_29843);
xnor UO_144 (O_144,N_29906,N_29981);
nor UO_145 (O_145,N_29847,N_29808);
and UO_146 (O_146,N_29898,N_29866);
xor UO_147 (O_147,N_29863,N_29807);
and UO_148 (O_148,N_29967,N_29930);
and UO_149 (O_149,N_29859,N_29825);
or UO_150 (O_150,N_29813,N_29881);
nor UO_151 (O_151,N_29840,N_29981);
nand UO_152 (O_152,N_29994,N_29801);
nand UO_153 (O_153,N_29865,N_29959);
xnor UO_154 (O_154,N_29917,N_29880);
and UO_155 (O_155,N_29936,N_29961);
nor UO_156 (O_156,N_29912,N_29801);
or UO_157 (O_157,N_29938,N_29859);
or UO_158 (O_158,N_29910,N_29887);
and UO_159 (O_159,N_29976,N_29986);
and UO_160 (O_160,N_29858,N_29883);
or UO_161 (O_161,N_29890,N_29879);
or UO_162 (O_162,N_29926,N_29994);
nand UO_163 (O_163,N_29885,N_29806);
nand UO_164 (O_164,N_29804,N_29963);
xnor UO_165 (O_165,N_29903,N_29885);
nor UO_166 (O_166,N_29980,N_29954);
and UO_167 (O_167,N_29931,N_29903);
or UO_168 (O_168,N_29811,N_29855);
and UO_169 (O_169,N_29915,N_29899);
xnor UO_170 (O_170,N_29995,N_29804);
nor UO_171 (O_171,N_29820,N_29972);
xor UO_172 (O_172,N_29905,N_29912);
nor UO_173 (O_173,N_29916,N_29899);
nor UO_174 (O_174,N_29991,N_29898);
xor UO_175 (O_175,N_29893,N_29998);
nand UO_176 (O_176,N_29964,N_29906);
nand UO_177 (O_177,N_29885,N_29926);
and UO_178 (O_178,N_29840,N_29933);
nor UO_179 (O_179,N_29819,N_29896);
xor UO_180 (O_180,N_29870,N_29975);
or UO_181 (O_181,N_29895,N_29968);
nand UO_182 (O_182,N_29986,N_29874);
xnor UO_183 (O_183,N_29962,N_29823);
and UO_184 (O_184,N_29859,N_29892);
and UO_185 (O_185,N_29938,N_29966);
and UO_186 (O_186,N_29915,N_29971);
nor UO_187 (O_187,N_29850,N_29938);
or UO_188 (O_188,N_29982,N_29889);
nor UO_189 (O_189,N_29830,N_29997);
nor UO_190 (O_190,N_29811,N_29810);
and UO_191 (O_191,N_29834,N_29917);
nor UO_192 (O_192,N_29890,N_29875);
and UO_193 (O_193,N_29832,N_29805);
xnor UO_194 (O_194,N_29892,N_29842);
or UO_195 (O_195,N_29893,N_29857);
xnor UO_196 (O_196,N_29914,N_29952);
and UO_197 (O_197,N_29978,N_29956);
xnor UO_198 (O_198,N_29984,N_29911);
xor UO_199 (O_199,N_29876,N_29907);
or UO_200 (O_200,N_29812,N_29973);
or UO_201 (O_201,N_29927,N_29970);
xnor UO_202 (O_202,N_29819,N_29982);
and UO_203 (O_203,N_29856,N_29969);
or UO_204 (O_204,N_29919,N_29865);
nand UO_205 (O_205,N_29806,N_29828);
nand UO_206 (O_206,N_29896,N_29820);
or UO_207 (O_207,N_29869,N_29960);
or UO_208 (O_208,N_29934,N_29826);
nand UO_209 (O_209,N_29841,N_29822);
or UO_210 (O_210,N_29802,N_29994);
or UO_211 (O_211,N_29823,N_29851);
xnor UO_212 (O_212,N_29822,N_29880);
nand UO_213 (O_213,N_29959,N_29863);
nor UO_214 (O_214,N_29993,N_29980);
nor UO_215 (O_215,N_29953,N_29972);
or UO_216 (O_216,N_29925,N_29947);
and UO_217 (O_217,N_29843,N_29921);
nor UO_218 (O_218,N_29910,N_29854);
nand UO_219 (O_219,N_29909,N_29999);
or UO_220 (O_220,N_29894,N_29915);
nand UO_221 (O_221,N_29984,N_29962);
nor UO_222 (O_222,N_29900,N_29895);
nand UO_223 (O_223,N_29854,N_29912);
xnor UO_224 (O_224,N_29800,N_29944);
and UO_225 (O_225,N_29890,N_29973);
or UO_226 (O_226,N_29895,N_29864);
nor UO_227 (O_227,N_29867,N_29980);
or UO_228 (O_228,N_29810,N_29894);
xor UO_229 (O_229,N_29919,N_29932);
nand UO_230 (O_230,N_29810,N_29890);
nor UO_231 (O_231,N_29829,N_29848);
or UO_232 (O_232,N_29968,N_29892);
nand UO_233 (O_233,N_29841,N_29854);
and UO_234 (O_234,N_29931,N_29995);
xor UO_235 (O_235,N_29817,N_29980);
or UO_236 (O_236,N_29946,N_29896);
and UO_237 (O_237,N_29968,N_29917);
nor UO_238 (O_238,N_29884,N_29985);
and UO_239 (O_239,N_29941,N_29936);
xnor UO_240 (O_240,N_29868,N_29998);
nor UO_241 (O_241,N_29930,N_29838);
or UO_242 (O_242,N_29818,N_29861);
nand UO_243 (O_243,N_29997,N_29979);
and UO_244 (O_244,N_29956,N_29822);
xnor UO_245 (O_245,N_29923,N_29984);
and UO_246 (O_246,N_29939,N_29970);
nand UO_247 (O_247,N_29974,N_29953);
xor UO_248 (O_248,N_29826,N_29916);
nand UO_249 (O_249,N_29953,N_29955);
nand UO_250 (O_250,N_29827,N_29834);
nor UO_251 (O_251,N_29826,N_29871);
nor UO_252 (O_252,N_29894,N_29852);
nor UO_253 (O_253,N_29867,N_29839);
xnor UO_254 (O_254,N_29872,N_29951);
or UO_255 (O_255,N_29808,N_29913);
xor UO_256 (O_256,N_29826,N_29820);
nor UO_257 (O_257,N_29903,N_29823);
nor UO_258 (O_258,N_29844,N_29865);
or UO_259 (O_259,N_29958,N_29923);
or UO_260 (O_260,N_29803,N_29993);
nand UO_261 (O_261,N_29992,N_29980);
and UO_262 (O_262,N_29897,N_29861);
nand UO_263 (O_263,N_29834,N_29832);
and UO_264 (O_264,N_29842,N_29884);
nand UO_265 (O_265,N_29876,N_29978);
nor UO_266 (O_266,N_29876,N_29847);
or UO_267 (O_267,N_29911,N_29915);
nor UO_268 (O_268,N_29806,N_29823);
nor UO_269 (O_269,N_29875,N_29956);
nor UO_270 (O_270,N_29828,N_29825);
nand UO_271 (O_271,N_29882,N_29928);
nand UO_272 (O_272,N_29956,N_29981);
or UO_273 (O_273,N_29954,N_29971);
nor UO_274 (O_274,N_29825,N_29952);
or UO_275 (O_275,N_29910,N_29982);
xor UO_276 (O_276,N_29998,N_29931);
or UO_277 (O_277,N_29884,N_29991);
or UO_278 (O_278,N_29993,N_29827);
xor UO_279 (O_279,N_29818,N_29944);
xor UO_280 (O_280,N_29999,N_29918);
xnor UO_281 (O_281,N_29905,N_29984);
and UO_282 (O_282,N_29825,N_29919);
xnor UO_283 (O_283,N_29830,N_29819);
nor UO_284 (O_284,N_29835,N_29880);
and UO_285 (O_285,N_29925,N_29831);
and UO_286 (O_286,N_29857,N_29954);
nor UO_287 (O_287,N_29906,N_29873);
or UO_288 (O_288,N_29845,N_29810);
xnor UO_289 (O_289,N_29813,N_29936);
and UO_290 (O_290,N_29947,N_29810);
and UO_291 (O_291,N_29875,N_29864);
and UO_292 (O_292,N_29855,N_29997);
or UO_293 (O_293,N_29803,N_29951);
nand UO_294 (O_294,N_29903,N_29859);
or UO_295 (O_295,N_29978,N_29981);
xor UO_296 (O_296,N_29839,N_29804);
and UO_297 (O_297,N_29912,N_29837);
xor UO_298 (O_298,N_29957,N_29837);
nor UO_299 (O_299,N_29926,N_29933);
xnor UO_300 (O_300,N_29973,N_29920);
or UO_301 (O_301,N_29846,N_29969);
or UO_302 (O_302,N_29964,N_29840);
or UO_303 (O_303,N_29981,N_29977);
or UO_304 (O_304,N_29832,N_29801);
nor UO_305 (O_305,N_29824,N_29801);
or UO_306 (O_306,N_29952,N_29966);
nor UO_307 (O_307,N_29966,N_29856);
or UO_308 (O_308,N_29881,N_29868);
xor UO_309 (O_309,N_29902,N_29960);
nand UO_310 (O_310,N_29939,N_29889);
nand UO_311 (O_311,N_29945,N_29842);
nor UO_312 (O_312,N_29943,N_29869);
or UO_313 (O_313,N_29902,N_29904);
nand UO_314 (O_314,N_29832,N_29907);
nand UO_315 (O_315,N_29966,N_29813);
xor UO_316 (O_316,N_29950,N_29979);
and UO_317 (O_317,N_29938,N_29838);
nor UO_318 (O_318,N_29856,N_29954);
or UO_319 (O_319,N_29885,N_29879);
xor UO_320 (O_320,N_29892,N_29929);
xor UO_321 (O_321,N_29911,N_29965);
nor UO_322 (O_322,N_29817,N_29882);
xor UO_323 (O_323,N_29988,N_29889);
nor UO_324 (O_324,N_29999,N_29833);
xnor UO_325 (O_325,N_29869,N_29812);
nand UO_326 (O_326,N_29864,N_29881);
and UO_327 (O_327,N_29875,N_29886);
nor UO_328 (O_328,N_29935,N_29814);
xnor UO_329 (O_329,N_29902,N_29919);
nor UO_330 (O_330,N_29807,N_29801);
nor UO_331 (O_331,N_29852,N_29893);
nor UO_332 (O_332,N_29806,N_29952);
nor UO_333 (O_333,N_29804,N_29865);
or UO_334 (O_334,N_29936,N_29893);
and UO_335 (O_335,N_29811,N_29803);
nor UO_336 (O_336,N_29974,N_29885);
or UO_337 (O_337,N_29824,N_29883);
and UO_338 (O_338,N_29957,N_29973);
nor UO_339 (O_339,N_29957,N_29869);
xnor UO_340 (O_340,N_29872,N_29894);
or UO_341 (O_341,N_29809,N_29942);
nand UO_342 (O_342,N_29977,N_29941);
nand UO_343 (O_343,N_29826,N_29991);
xnor UO_344 (O_344,N_29893,N_29959);
and UO_345 (O_345,N_29991,N_29929);
nor UO_346 (O_346,N_29822,N_29953);
xnor UO_347 (O_347,N_29810,N_29865);
and UO_348 (O_348,N_29916,N_29942);
xor UO_349 (O_349,N_29866,N_29984);
and UO_350 (O_350,N_29842,N_29830);
and UO_351 (O_351,N_29919,N_29889);
or UO_352 (O_352,N_29992,N_29868);
xor UO_353 (O_353,N_29958,N_29804);
nand UO_354 (O_354,N_29913,N_29844);
and UO_355 (O_355,N_29997,N_29815);
and UO_356 (O_356,N_29829,N_29850);
nor UO_357 (O_357,N_29951,N_29871);
nor UO_358 (O_358,N_29862,N_29963);
nor UO_359 (O_359,N_29987,N_29933);
nor UO_360 (O_360,N_29989,N_29900);
nand UO_361 (O_361,N_29810,N_29879);
xor UO_362 (O_362,N_29910,N_29884);
xnor UO_363 (O_363,N_29986,N_29800);
nor UO_364 (O_364,N_29850,N_29807);
nand UO_365 (O_365,N_29976,N_29973);
nand UO_366 (O_366,N_29925,N_29809);
nand UO_367 (O_367,N_29879,N_29878);
nor UO_368 (O_368,N_29872,N_29974);
nor UO_369 (O_369,N_29999,N_29845);
nand UO_370 (O_370,N_29931,N_29806);
nor UO_371 (O_371,N_29915,N_29918);
xor UO_372 (O_372,N_29899,N_29833);
nand UO_373 (O_373,N_29976,N_29956);
xnor UO_374 (O_374,N_29883,N_29951);
and UO_375 (O_375,N_29940,N_29958);
nor UO_376 (O_376,N_29955,N_29851);
nor UO_377 (O_377,N_29994,N_29837);
or UO_378 (O_378,N_29912,N_29906);
and UO_379 (O_379,N_29981,N_29874);
xnor UO_380 (O_380,N_29865,N_29884);
xnor UO_381 (O_381,N_29919,N_29893);
and UO_382 (O_382,N_29840,N_29998);
or UO_383 (O_383,N_29898,N_29917);
and UO_384 (O_384,N_29852,N_29970);
and UO_385 (O_385,N_29840,N_29816);
nand UO_386 (O_386,N_29805,N_29963);
or UO_387 (O_387,N_29984,N_29979);
nand UO_388 (O_388,N_29846,N_29881);
xnor UO_389 (O_389,N_29800,N_29843);
xor UO_390 (O_390,N_29858,N_29963);
nand UO_391 (O_391,N_29851,N_29990);
nand UO_392 (O_392,N_29986,N_29967);
nor UO_393 (O_393,N_29999,N_29830);
nand UO_394 (O_394,N_29815,N_29853);
nand UO_395 (O_395,N_29982,N_29926);
or UO_396 (O_396,N_29935,N_29803);
or UO_397 (O_397,N_29916,N_29844);
nor UO_398 (O_398,N_29828,N_29852);
and UO_399 (O_399,N_29877,N_29804);
nor UO_400 (O_400,N_29941,N_29875);
and UO_401 (O_401,N_29991,N_29961);
xnor UO_402 (O_402,N_29952,N_29824);
nand UO_403 (O_403,N_29857,N_29907);
nand UO_404 (O_404,N_29829,N_29979);
xor UO_405 (O_405,N_29925,N_29887);
or UO_406 (O_406,N_29849,N_29812);
xnor UO_407 (O_407,N_29892,N_29961);
nand UO_408 (O_408,N_29941,N_29911);
and UO_409 (O_409,N_29918,N_29802);
nor UO_410 (O_410,N_29892,N_29959);
nand UO_411 (O_411,N_29980,N_29878);
xor UO_412 (O_412,N_29875,N_29995);
and UO_413 (O_413,N_29981,N_29801);
and UO_414 (O_414,N_29823,N_29910);
nor UO_415 (O_415,N_29867,N_29905);
and UO_416 (O_416,N_29903,N_29871);
or UO_417 (O_417,N_29899,N_29862);
or UO_418 (O_418,N_29891,N_29999);
nand UO_419 (O_419,N_29900,N_29870);
xnor UO_420 (O_420,N_29970,N_29973);
and UO_421 (O_421,N_29819,N_29826);
nand UO_422 (O_422,N_29808,N_29958);
nand UO_423 (O_423,N_29988,N_29933);
xnor UO_424 (O_424,N_29986,N_29912);
or UO_425 (O_425,N_29879,N_29835);
nor UO_426 (O_426,N_29927,N_29972);
nand UO_427 (O_427,N_29852,N_29851);
or UO_428 (O_428,N_29948,N_29831);
or UO_429 (O_429,N_29961,N_29822);
xor UO_430 (O_430,N_29884,N_29914);
xor UO_431 (O_431,N_29967,N_29846);
nor UO_432 (O_432,N_29928,N_29973);
and UO_433 (O_433,N_29836,N_29909);
or UO_434 (O_434,N_29964,N_29905);
or UO_435 (O_435,N_29949,N_29919);
xor UO_436 (O_436,N_29950,N_29983);
and UO_437 (O_437,N_29816,N_29854);
xor UO_438 (O_438,N_29967,N_29803);
nor UO_439 (O_439,N_29815,N_29805);
xor UO_440 (O_440,N_29993,N_29862);
or UO_441 (O_441,N_29899,N_29998);
and UO_442 (O_442,N_29969,N_29895);
nor UO_443 (O_443,N_29888,N_29823);
and UO_444 (O_444,N_29860,N_29994);
xor UO_445 (O_445,N_29835,N_29842);
nor UO_446 (O_446,N_29972,N_29849);
xnor UO_447 (O_447,N_29979,N_29879);
or UO_448 (O_448,N_29992,N_29918);
nor UO_449 (O_449,N_29999,N_29857);
or UO_450 (O_450,N_29832,N_29896);
or UO_451 (O_451,N_29943,N_29992);
and UO_452 (O_452,N_29850,N_29852);
and UO_453 (O_453,N_29998,N_29985);
xnor UO_454 (O_454,N_29886,N_29931);
nor UO_455 (O_455,N_29971,N_29836);
or UO_456 (O_456,N_29858,N_29809);
nand UO_457 (O_457,N_29810,N_29833);
and UO_458 (O_458,N_29853,N_29891);
nor UO_459 (O_459,N_29880,N_29995);
or UO_460 (O_460,N_29933,N_29921);
nand UO_461 (O_461,N_29896,N_29877);
or UO_462 (O_462,N_29978,N_29820);
nor UO_463 (O_463,N_29883,N_29935);
nor UO_464 (O_464,N_29905,N_29859);
xor UO_465 (O_465,N_29917,N_29816);
xnor UO_466 (O_466,N_29902,N_29894);
nand UO_467 (O_467,N_29962,N_29899);
nor UO_468 (O_468,N_29983,N_29889);
nand UO_469 (O_469,N_29842,N_29972);
xor UO_470 (O_470,N_29988,N_29898);
nor UO_471 (O_471,N_29959,N_29838);
or UO_472 (O_472,N_29874,N_29887);
nand UO_473 (O_473,N_29945,N_29991);
or UO_474 (O_474,N_29869,N_29976);
nand UO_475 (O_475,N_29998,N_29916);
and UO_476 (O_476,N_29931,N_29883);
and UO_477 (O_477,N_29967,N_29801);
or UO_478 (O_478,N_29923,N_29824);
xor UO_479 (O_479,N_29956,N_29958);
xor UO_480 (O_480,N_29952,N_29849);
nand UO_481 (O_481,N_29813,N_29933);
nand UO_482 (O_482,N_29951,N_29900);
and UO_483 (O_483,N_29896,N_29928);
nor UO_484 (O_484,N_29992,N_29946);
or UO_485 (O_485,N_29974,N_29909);
nand UO_486 (O_486,N_29991,N_29859);
xor UO_487 (O_487,N_29837,N_29848);
or UO_488 (O_488,N_29959,N_29867);
or UO_489 (O_489,N_29949,N_29831);
nand UO_490 (O_490,N_29988,N_29811);
nor UO_491 (O_491,N_29905,N_29881);
nor UO_492 (O_492,N_29998,N_29805);
and UO_493 (O_493,N_29913,N_29921);
nand UO_494 (O_494,N_29813,N_29994);
nor UO_495 (O_495,N_29956,N_29849);
xnor UO_496 (O_496,N_29994,N_29976);
xnor UO_497 (O_497,N_29981,N_29962);
nand UO_498 (O_498,N_29922,N_29978);
nand UO_499 (O_499,N_29849,N_29953);
and UO_500 (O_500,N_29835,N_29869);
or UO_501 (O_501,N_29946,N_29986);
and UO_502 (O_502,N_29849,N_29872);
nand UO_503 (O_503,N_29813,N_29910);
or UO_504 (O_504,N_29929,N_29968);
xor UO_505 (O_505,N_29941,N_29939);
xnor UO_506 (O_506,N_29921,N_29885);
nor UO_507 (O_507,N_29988,N_29950);
nor UO_508 (O_508,N_29981,N_29892);
nand UO_509 (O_509,N_29974,N_29949);
xor UO_510 (O_510,N_29944,N_29909);
xor UO_511 (O_511,N_29924,N_29977);
and UO_512 (O_512,N_29849,N_29809);
and UO_513 (O_513,N_29904,N_29888);
nor UO_514 (O_514,N_29961,N_29981);
nand UO_515 (O_515,N_29870,N_29892);
and UO_516 (O_516,N_29843,N_29914);
and UO_517 (O_517,N_29894,N_29985);
nand UO_518 (O_518,N_29824,N_29928);
nand UO_519 (O_519,N_29912,N_29904);
xor UO_520 (O_520,N_29818,N_29852);
nor UO_521 (O_521,N_29999,N_29961);
or UO_522 (O_522,N_29983,N_29830);
nor UO_523 (O_523,N_29837,N_29820);
nor UO_524 (O_524,N_29987,N_29959);
nor UO_525 (O_525,N_29980,N_29810);
or UO_526 (O_526,N_29903,N_29881);
or UO_527 (O_527,N_29894,N_29980);
xnor UO_528 (O_528,N_29879,N_29928);
nor UO_529 (O_529,N_29848,N_29948);
xor UO_530 (O_530,N_29993,N_29984);
and UO_531 (O_531,N_29938,N_29920);
xor UO_532 (O_532,N_29856,N_29879);
xor UO_533 (O_533,N_29973,N_29810);
nand UO_534 (O_534,N_29940,N_29997);
xnor UO_535 (O_535,N_29906,N_29816);
or UO_536 (O_536,N_29920,N_29883);
xnor UO_537 (O_537,N_29801,N_29965);
xnor UO_538 (O_538,N_29989,N_29982);
and UO_539 (O_539,N_29939,N_29958);
xnor UO_540 (O_540,N_29993,N_29960);
nand UO_541 (O_541,N_29804,N_29921);
and UO_542 (O_542,N_29882,N_29850);
xor UO_543 (O_543,N_29903,N_29906);
xor UO_544 (O_544,N_29802,N_29903);
or UO_545 (O_545,N_29945,N_29811);
and UO_546 (O_546,N_29924,N_29872);
nor UO_547 (O_547,N_29871,N_29958);
or UO_548 (O_548,N_29899,N_29835);
nor UO_549 (O_549,N_29943,N_29882);
nor UO_550 (O_550,N_29805,N_29962);
xor UO_551 (O_551,N_29809,N_29802);
or UO_552 (O_552,N_29866,N_29862);
xor UO_553 (O_553,N_29817,N_29945);
xnor UO_554 (O_554,N_29804,N_29910);
nand UO_555 (O_555,N_29920,N_29862);
or UO_556 (O_556,N_29966,N_29880);
nand UO_557 (O_557,N_29803,N_29886);
nand UO_558 (O_558,N_29913,N_29987);
xor UO_559 (O_559,N_29879,N_29800);
and UO_560 (O_560,N_29897,N_29930);
or UO_561 (O_561,N_29857,N_29839);
or UO_562 (O_562,N_29937,N_29856);
nand UO_563 (O_563,N_29997,N_29849);
nand UO_564 (O_564,N_29924,N_29918);
and UO_565 (O_565,N_29823,N_29819);
xor UO_566 (O_566,N_29807,N_29985);
nor UO_567 (O_567,N_29892,N_29900);
xor UO_568 (O_568,N_29845,N_29877);
nand UO_569 (O_569,N_29938,N_29992);
and UO_570 (O_570,N_29832,N_29824);
and UO_571 (O_571,N_29951,N_29823);
or UO_572 (O_572,N_29838,N_29912);
xor UO_573 (O_573,N_29982,N_29915);
and UO_574 (O_574,N_29999,N_29882);
and UO_575 (O_575,N_29870,N_29933);
xnor UO_576 (O_576,N_29889,N_29934);
and UO_577 (O_577,N_29967,N_29804);
nor UO_578 (O_578,N_29851,N_29853);
and UO_579 (O_579,N_29954,N_29832);
xor UO_580 (O_580,N_29865,N_29872);
nor UO_581 (O_581,N_29972,N_29868);
xnor UO_582 (O_582,N_29857,N_29871);
nand UO_583 (O_583,N_29859,N_29841);
nand UO_584 (O_584,N_29839,N_29960);
xor UO_585 (O_585,N_29875,N_29858);
and UO_586 (O_586,N_29961,N_29984);
nor UO_587 (O_587,N_29821,N_29858);
or UO_588 (O_588,N_29997,N_29902);
nor UO_589 (O_589,N_29977,N_29979);
xnor UO_590 (O_590,N_29836,N_29997);
and UO_591 (O_591,N_29801,N_29820);
nor UO_592 (O_592,N_29961,N_29853);
xor UO_593 (O_593,N_29866,N_29805);
and UO_594 (O_594,N_29864,N_29932);
or UO_595 (O_595,N_29962,N_29806);
xor UO_596 (O_596,N_29802,N_29829);
and UO_597 (O_597,N_29966,N_29928);
or UO_598 (O_598,N_29955,N_29990);
xnor UO_599 (O_599,N_29965,N_29987);
and UO_600 (O_600,N_29980,N_29871);
nor UO_601 (O_601,N_29838,N_29899);
and UO_602 (O_602,N_29838,N_29980);
and UO_603 (O_603,N_29803,N_29827);
nor UO_604 (O_604,N_29831,N_29814);
and UO_605 (O_605,N_29981,N_29882);
nand UO_606 (O_606,N_29891,N_29821);
nand UO_607 (O_607,N_29942,N_29952);
or UO_608 (O_608,N_29900,N_29802);
or UO_609 (O_609,N_29860,N_29906);
or UO_610 (O_610,N_29949,N_29868);
or UO_611 (O_611,N_29954,N_29816);
and UO_612 (O_612,N_29951,N_29832);
nor UO_613 (O_613,N_29841,N_29876);
or UO_614 (O_614,N_29804,N_29812);
or UO_615 (O_615,N_29969,N_29825);
and UO_616 (O_616,N_29956,N_29994);
and UO_617 (O_617,N_29912,N_29994);
or UO_618 (O_618,N_29921,N_29844);
xor UO_619 (O_619,N_29976,N_29959);
and UO_620 (O_620,N_29859,N_29931);
and UO_621 (O_621,N_29894,N_29944);
nor UO_622 (O_622,N_29813,N_29876);
xnor UO_623 (O_623,N_29983,N_29967);
nor UO_624 (O_624,N_29978,N_29848);
nor UO_625 (O_625,N_29845,N_29939);
nand UO_626 (O_626,N_29970,N_29829);
nand UO_627 (O_627,N_29962,N_29968);
nand UO_628 (O_628,N_29975,N_29979);
xnor UO_629 (O_629,N_29959,N_29870);
xor UO_630 (O_630,N_29876,N_29949);
xor UO_631 (O_631,N_29994,N_29971);
nand UO_632 (O_632,N_29865,N_29873);
or UO_633 (O_633,N_29961,N_29873);
nand UO_634 (O_634,N_29874,N_29855);
xor UO_635 (O_635,N_29815,N_29897);
xnor UO_636 (O_636,N_29908,N_29923);
nand UO_637 (O_637,N_29831,N_29946);
or UO_638 (O_638,N_29919,N_29844);
nor UO_639 (O_639,N_29944,N_29819);
nor UO_640 (O_640,N_29896,N_29879);
nand UO_641 (O_641,N_29902,N_29833);
and UO_642 (O_642,N_29929,N_29896);
nand UO_643 (O_643,N_29920,N_29879);
nor UO_644 (O_644,N_29976,N_29882);
xor UO_645 (O_645,N_29912,N_29802);
nand UO_646 (O_646,N_29884,N_29879);
nor UO_647 (O_647,N_29950,N_29804);
and UO_648 (O_648,N_29947,N_29812);
or UO_649 (O_649,N_29902,N_29819);
nand UO_650 (O_650,N_29939,N_29954);
nor UO_651 (O_651,N_29846,N_29801);
xor UO_652 (O_652,N_29971,N_29904);
nand UO_653 (O_653,N_29914,N_29909);
xnor UO_654 (O_654,N_29904,N_29899);
and UO_655 (O_655,N_29995,N_29944);
nand UO_656 (O_656,N_29857,N_29811);
and UO_657 (O_657,N_29966,N_29923);
or UO_658 (O_658,N_29857,N_29814);
or UO_659 (O_659,N_29887,N_29957);
xnor UO_660 (O_660,N_29941,N_29889);
xor UO_661 (O_661,N_29842,N_29852);
xnor UO_662 (O_662,N_29959,N_29868);
nand UO_663 (O_663,N_29993,N_29896);
and UO_664 (O_664,N_29893,N_29882);
nand UO_665 (O_665,N_29884,N_29981);
xnor UO_666 (O_666,N_29860,N_29817);
nand UO_667 (O_667,N_29817,N_29983);
and UO_668 (O_668,N_29907,N_29810);
or UO_669 (O_669,N_29862,N_29840);
nor UO_670 (O_670,N_29886,N_29893);
xor UO_671 (O_671,N_29906,N_29895);
and UO_672 (O_672,N_29924,N_29954);
nand UO_673 (O_673,N_29824,N_29885);
nor UO_674 (O_674,N_29805,N_29981);
or UO_675 (O_675,N_29860,N_29949);
xor UO_676 (O_676,N_29815,N_29999);
or UO_677 (O_677,N_29947,N_29866);
nor UO_678 (O_678,N_29817,N_29813);
xnor UO_679 (O_679,N_29982,N_29817);
nor UO_680 (O_680,N_29919,N_29996);
nand UO_681 (O_681,N_29976,N_29970);
nand UO_682 (O_682,N_29895,N_29951);
or UO_683 (O_683,N_29956,N_29848);
nor UO_684 (O_684,N_29911,N_29887);
nand UO_685 (O_685,N_29890,N_29924);
nor UO_686 (O_686,N_29879,N_29985);
or UO_687 (O_687,N_29823,N_29993);
xnor UO_688 (O_688,N_29839,N_29825);
or UO_689 (O_689,N_29867,N_29860);
xnor UO_690 (O_690,N_29950,N_29964);
nor UO_691 (O_691,N_29939,N_29932);
nand UO_692 (O_692,N_29839,N_29929);
nand UO_693 (O_693,N_29989,N_29800);
or UO_694 (O_694,N_29974,N_29815);
xor UO_695 (O_695,N_29973,N_29992);
and UO_696 (O_696,N_29927,N_29969);
and UO_697 (O_697,N_29999,N_29967);
nand UO_698 (O_698,N_29838,N_29921);
or UO_699 (O_699,N_29825,N_29921);
nor UO_700 (O_700,N_29983,N_29839);
nor UO_701 (O_701,N_29993,N_29828);
and UO_702 (O_702,N_29914,N_29835);
nor UO_703 (O_703,N_29889,N_29880);
xor UO_704 (O_704,N_29871,N_29909);
xnor UO_705 (O_705,N_29979,N_29850);
or UO_706 (O_706,N_29822,N_29849);
nand UO_707 (O_707,N_29953,N_29960);
or UO_708 (O_708,N_29915,N_29926);
nor UO_709 (O_709,N_29877,N_29840);
nand UO_710 (O_710,N_29994,N_29946);
and UO_711 (O_711,N_29941,N_29833);
or UO_712 (O_712,N_29979,N_29803);
nand UO_713 (O_713,N_29956,N_29983);
and UO_714 (O_714,N_29855,N_29994);
and UO_715 (O_715,N_29894,N_29815);
nor UO_716 (O_716,N_29961,N_29884);
and UO_717 (O_717,N_29839,N_29809);
or UO_718 (O_718,N_29995,N_29801);
nand UO_719 (O_719,N_29842,N_29888);
xor UO_720 (O_720,N_29995,N_29884);
nand UO_721 (O_721,N_29890,N_29893);
nand UO_722 (O_722,N_29983,N_29973);
nor UO_723 (O_723,N_29959,N_29878);
or UO_724 (O_724,N_29841,N_29931);
or UO_725 (O_725,N_29859,N_29803);
and UO_726 (O_726,N_29980,N_29978);
or UO_727 (O_727,N_29966,N_29898);
xnor UO_728 (O_728,N_29940,N_29988);
nor UO_729 (O_729,N_29959,N_29982);
xnor UO_730 (O_730,N_29930,N_29914);
xor UO_731 (O_731,N_29996,N_29867);
and UO_732 (O_732,N_29951,N_29919);
xor UO_733 (O_733,N_29965,N_29921);
xor UO_734 (O_734,N_29990,N_29879);
and UO_735 (O_735,N_29938,N_29888);
nor UO_736 (O_736,N_29851,N_29892);
nand UO_737 (O_737,N_29985,N_29848);
nand UO_738 (O_738,N_29903,N_29979);
or UO_739 (O_739,N_29806,N_29914);
nor UO_740 (O_740,N_29828,N_29965);
xor UO_741 (O_741,N_29879,N_29828);
and UO_742 (O_742,N_29909,N_29837);
nor UO_743 (O_743,N_29933,N_29809);
xor UO_744 (O_744,N_29909,N_29888);
or UO_745 (O_745,N_29842,N_29856);
xor UO_746 (O_746,N_29803,N_29986);
and UO_747 (O_747,N_29816,N_29818);
xor UO_748 (O_748,N_29953,N_29905);
xor UO_749 (O_749,N_29947,N_29936);
nand UO_750 (O_750,N_29943,N_29962);
or UO_751 (O_751,N_29819,N_29909);
nand UO_752 (O_752,N_29954,N_29887);
xor UO_753 (O_753,N_29817,N_29908);
or UO_754 (O_754,N_29895,N_29822);
and UO_755 (O_755,N_29824,N_29960);
and UO_756 (O_756,N_29890,N_29960);
nand UO_757 (O_757,N_29884,N_29958);
xnor UO_758 (O_758,N_29829,N_29914);
or UO_759 (O_759,N_29965,N_29934);
nor UO_760 (O_760,N_29804,N_29901);
or UO_761 (O_761,N_29933,N_29819);
or UO_762 (O_762,N_29964,N_29800);
and UO_763 (O_763,N_29952,N_29878);
nand UO_764 (O_764,N_29843,N_29853);
nand UO_765 (O_765,N_29898,N_29865);
nor UO_766 (O_766,N_29965,N_29982);
nor UO_767 (O_767,N_29891,N_29822);
xor UO_768 (O_768,N_29889,N_29990);
and UO_769 (O_769,N_29923,N_29887);
xor UO_770 (O_770,N_29884,N_29805);
and UO_771 (O_771,N_29978,N_29987);
and UO_772 (O_772,N_29856,N_29902);
and UO_773 (O_773,N_29879,N_29917);
nand UO_774 (O_774,N_29904,N_29829);
and UO_775 (O_775,N_29874,N_29835);
nor UO_776 (O_776,N_29844,N_29970);
nor UO_777 (O_777,N_29898,N_29850);
xor UO_778 (O_778,N_29840,N_29838);
nand UO_779 (O_779,N_29901,N_29826);
nand UO_780 (O_780,N_29867,N_29813);
and UO_781 (O_781,N_29916,N_29971);
nor UO_782 (O_782,N_29888,N_29995);
xnor UO_783 (O_783,N_29978,N_29929);
nor UO_784 (O_784,N_29999,N_29920);
xnor UO_785 (O_785,N_29880,N_29989);
nand UO_786 (O_786,N_29839,N_29828);
and UO_787 (O_787,N_29856,N_29990);
xnor UO_788 (O_788,N_29825,N_29858);
nor UO_789 (O_789,N_29981,N_29938);
and UO_790 (O_790,N_29879,N_29910);
xor UO_791 (O_791,N_29843,N_29809);
xor UO_792 (O_792,N_29991,N_29912);
nor UO_793 (O_793,N_29976,N_29909);
nand UO_794 (O_794,N_29950,N_29873);
nand UO_795 (O_795,N_29957,N_29848);
and UO_796 (O_796,N_29848,N_29858);
nor UO_797 (O_797,N_29924,N_29875);
and UO_798 (O_798,N_29940,N_29850);
nor UO_799 (O_799,N_29975,N_29944);
xnor UO_800 (O_800,N_29977,N_29825);
or UO_801 (O_801,N_29844,N_29933);
nor UO_802 (O_802,N_29868,N_29821);
and UO_803 (O_803,N_29965,N_29883);
xor UO_804 (O_804,N_29913,N_29847);
or UO_805 (O_805,N_29911,N_29808);
nor UO_806 (O_806,N_29963,N_29961);
nor UO_807 (O_807,N_29879,N_29850);
nor UO_808 (O_808,N_29918,N_29842);
xor UO_809 (O_809,N_29977,N_29972);
and UO_810 (O_810,N_29965,N_29959);
and UO_811 (O_811,N_29850,N_29916);
nor UO_812 (O_812,N_29992,N_29999);
xor UO_813 (O_813,N_29898,N_29861);
and UO_814 (O_814,N_29976,N_29925);
nand UO_815 (O_815,N_29952,N_29940);
xor UO_816 (O_816,N_29817,N_29943);
and UO_817 (O_817,N_29846,N_29913);
or UO_818 (O_818,N_29903,N_29987);
or UO_819 (O_819,N_29905,N_29891);
nor UO_820 (O_820,N_29992,N_29833);
nor UO_821 (O_821,N_29902,N_29982);
and UO_822 (O_822,N_29994,N_29847);
or UO_823 (O_823,N_29872,N_29838);
nor UO_824 (O_824,N_29971,N_29853);
and UO_825 (O_825,N_29803,N_29955);
or UO_826 (O_826,N_29933,N_29886);
or UO_827 (O_827,N_29858,N_29934);
or UO_828 (O_828,N_29957,N_29809);
nor UO_829 (O_829,N_29912,N_29996);
xor UO_830 (O_830,N_29917,N_29888);
xnor UO_831 (O_831,N_29906,N_29957);
and UO_832 (O_832,N_29916,N_29888);
nor UO_833 (O_833,N_29864,N_29829);
nand UO_834 (O_834,N_29833,N_29933);
xor UO_835 (O_835,N_29813,N_29967);
or UO_836 (O_836,N_29981,N_29812);
and UO_837 (O_837,N_29801,N_29836);
xnor UO_838 (O_838,N_29928,N_29830);
or UO_839 (O_839,N_29956,N_29805);
nor UO_840 (O_840,N_29833,N_29865);
or UO_841 (O_841,N_29889,N_29914);
nand UO_842 (O_842,N_29807,N_29982);
xnor UO_843 (O_843,N_29823,N_29861);
xor UO_844 (O_844,N_29853,N_29935);
nor UO_845 (O_845,N_29920,N_29989);
nand UO_846 (O_846,N_29997,N_29867);
xnor UO_847 (O_847,N_29839,N_29802);
nor UO_848 (O_848,N_29807,N_29892);
and UO_849 (O_849,N_29820,N_29865);
nand UO_850 (O_850,N_29831,N_29939);
nand UO_851 (O_851,N_29833,N_29905);
xor UO_852 (O_852,N_29894,N_29949);
nor UO_853 (O_853,N_29969,N_29874);
nand UO_854 (O_854,N_29960,N_29985);
xnor UO_855 (O_855,N_29825,N_29901);
or UO_856 (O_856,N_29838,N_29935);
or UO_857 (O_857,N_29953,N_29947);
and UO_858 (O_858,N_29871,N_29867);
or UO_859 (O_859,N_29812,N_29922);
xor UO_860 (O_860,N_29876,N_29958);
nand UO_861 (O_861,N_29992,N_29803);
or UO_862 (O_862,N_29965,N_29806);
and UO_863 (O_863,N_29941,N_29800);
nand UO_864 (O_864,N_29825,N_29959);
or UO_865 (O_865,N_29802,N_29943);
nor UO_866 (O_866,N_29977,N_29999);
or UO_867 (O_867,N_29845,N_29826);
and UO_868 (O_868,N_29937,N_29812);
or UO_869 (O_869,N_29839,N_29805);
or UO_870 (O_870,N_29858,N_29873);
nor UO_871 (O_871,N_29960,N_29888);
or UO_872 (O_872,N_29943,N_29890);
xnor UO_873 (O_873,N_29962,N_29862);
nand UO_874 (O_874,N_29818,N_29882);
xor UO_875 (O_875,N_29822,N_29949);
and UO_876 (O_876,N_29834,N_29976);
or UO_877 (O_877,N_29948,N_29950);
or UO_878 (O_878,N_29813,N_29999);
xnor UO_879 (O_879,N_29895,N_29911);
or UO_880 (O_880,N_29892,N_29821);
or UO_881 (O_881,N_29927,N_29966);
and UO_882 (O_882,N_29881,N_29876);
and UO_883 (O_883,N_29846,N_29995);
nor UO_884 (O_884,N_29833,N_29820);
and UO_885 (O_885,N_29851,N_29986);
nand UO_886 (O_886,N_29937,N_29877);
and UO_887 (O_887,N_29917,N_29955);
nor UO_888 (O_888,N_29945,N_29861);
xor UO_889 (O_889,N_29921,N_29919);
and UO_890 (O_890,N_29924,N_29914);
nand UO_891 (O_891,N_29967,N_29976);
nor UO_892 (O_892,N_29845,N_29989);
xnor UO_893 (O_893,N_29921,N_29935);
nand UO_894 (O_894,N_29812,N_29976);
nor UO_895 (O_895,N_29933,N_29800);
xor UO_896 (O_896,N_29822,N_29814);
xnor UO_897 (O_897,N_29969,N_29814);
or UO_898 (O_898,N_29887,N_29881);
and UO_899 (O_899,N_29914,N_29871);
nor UO_900 (O_900,N_29844,N_29807);
xnor UO_901 (O_901,N_29851,N_29928);
xnor UO_902 (O_902,N_29867,N_29939);
nor UO_903 (O_903,N_29916,N_29977);
or UO_904 (O_904,N_29944,N_29922);
or UO_905 (O_905,N_29906,N_29856);
nor UO_906 (O_906,N_29853,N_29996);
and UO_907 (O_907,N_29802,N_29825);
or UO_908 (O_908,N_29950,N_29965);
nor UO_909 (O_909,N_29911,N_29850);
nand UO_910 (O_910,N_29903,N_29968);
nand UO_911 (O_911,N_29832,N_29902);
nand UO_912 (O_912,N_29942,N_29921);
or UO_913 (O_913,N_29936,N_29894);
or UO_914 (O_914,N_29966,N_29814);
and UO_915 (O_915,N_29966,N_29888);
and UO_916 (O_916,N_29844,N_29931);
and UO_917 (O_917,N_29946,N_29926);
nand UO_918 (O_918,N_29962,N_29802);
and UO_919 (O_919,N_29980,N_29862);
or UO_920 (O_920,N_29938,N_29890);
nor UO_921 (O_921,N_29875,N_29865);
and UO_922 (O_922,N_29919,N_29938);
nand UO_923 (O_923,N_29922,N_29983);
xor UO_924 (O_924,N_29876,N_29820);
and UO_925 (O_925,N_29894,N_29883);
xor UO_926 (O_926,N_29989,N_29978);
or UO_927 (O_927,N_29990,N_29877);
nor UO_928 (O_928,N_29908,N_29844);
and UO_929 (O_929,N_29952,N_29943);
or UO_930 (O_930,N_29836,N_29958);
nor UO_931 (O_931,N_29957,N_29893);
nor UO_932 (O_932,N_29866,N_29967);
nand UO_933 (O_933,N_29827,N_29829);
nor UO_934 (O_934,N_29926,N_29845);
or UO_935 (O_935,N_29862,N_29914);
nor UO_936 (O_936,N_29968,N_29819);
xnor UO_937 (O_937,N_29901,N_29934);
nand UO_938 (O_938,N_29905,N_29974);
or UO_939 (O_939,N_29972,N_29994);
and UO_940 (O_940,N_29914,N_29817);
nor UO_941 (O_941,N_29862,N_29911);
or UO_942 (O_942,N_29847,N_29956);
and UO_943 (O_943,N_29856,N_29953);
and UO_944 (O_944,N_29806,N_29847);
nor UO_945 (O_945,N_29890,N_29804);
xnor UO_946 (O_946,N_29866,N_29980);
nand UO_947 (O_947,N_29872,N_29933);
nor UO_948 (O_948,N_29954,N_29827);
xnor UO_949 (O_949,N_29942,N_29931);
nor UO_950 (O_950,N_29938,N_29997);
or UO_951 (O_951,N_29987,N_29941);
nand UO_952 (O_952,N_29867,N_29963);
or UO_953 (O_953,N_29911,N_29946);
xor UO_954 (O_954,N_29867,N_29987);
nor UO_955 (O_955,N_29934,N_29972);
or UO_956 (O_956,N_29940,N_29949);
or UO_957 (O_957,N_29816,N_29862);
and UO_958 (O_958,N_29961,N_29979);
or UO_959 (O_959,N_29833,N_29852);
or UO_960 (O_960,N_29993,N_29858);
nand UO_961 (O_961,N_29987,N_29989);
nor UO_962 (O_962,N_29947,N_29938);
nand UO_963 (O_963,N_29940,N_29893);
xnor UO_964 (O_964,N_29988,N_29856);
nor UO_965 (O_965,N_29829,N_29994);
and UO_966 (O_966,N_29860,N_29872);
or UO_967 (O_967,N_29849,N_29973);
nand UO_968 (O_968,N_29921,N_29823);
and UO_969 (O_969,N_29954,N_29985);
nand UO_970 (O_970,N_29826,N_29973);
nor UO_971 (O_971,N_29854,N_29921);
or UO_972 (O_972,N_29961,N_29867);
and UO_973 (O_973,N_29910,N_29924);
or UO_974 (O_974,N_29876,N_29863);
xnor UO_975 (O_975,N_29977,N_29973);
or UO_976 (O_976,N_29874,N_29816);
nand UO_977 (O_977,N_29967,N_29928);
nor UO_978 (O_978,N_29942,N_29812);
nor UO_979 (O_979,N_29945,N_29961);
nand UO_980 (O_980,N_29990,N_29874);
xor UO_981 (O_981,N_29909,N_29813);
nor UO_982 (O_982,N_29895,N_29910);
or UO_983 (O_983,N_29808,N_29979);
and UO_984 (O_984,N_29972,N_29866);
or UO_985 (O_985,N_29999,N_29841);
nand UO_986 (O_986,N_29973,N_29813);
and UO_987 (O_987,N_29901,N_29802);
and UO_988 (O_988,N_29919,N_29864);
nor UO_989 (O_989,N_29902,N_29933);
and UO_990 (O_990,N_29847,N_29993);
nand UO_991 (O_991,N_29909,N_29952);
nor UO_992 (O_992,N_29976,N_29907);
xor UO_993 (O_993,N_29834,N_29874);
and UO_994 (O_994,N_29930,N_29823);
nand UO_995 (O_995,N_29993,N_29956);
xor UO_996 (O_996,N_29809,N_29833);
or UO_997 (O_997,N_29933,N_29845);
or UO_998 (O_998,N_29824,N_29842);
or UO_999 (O_999,N_29917,N_29950);
or UO_1000 (O_1000,N_29956,N_29828);
nor UO_1001 (O_1001,N_29972,N_29976);
nand UO_1002 (O_1002,N_29921,N_29882);
xnor UO_1003 (O_1003,N_29940,N_29804);
nand UO_1004 (O_1004,N_29892,N_29848);
and UO_1005 (O_1005,N_29860,N_29955);
nand UO_1006 (O_1006,N_29985,N_29802);
or UO_1007 (O_1007,N_29922,N_29885);
and UO_1008 (O_1008,N_29937,N_29972);
xnor UO_1009 (O_1009,N_29838,N_29942);
xnor UO_1010 (O_1010,N_29807,N_29962);
and UO_1011 (O_1011,N_29920,N_29901);
and UO_1012 (O_1012,N_29986,N_29868);
or UO_1013 (O_1013,N_29809,N_29882);
and UO_1014 (O_1014,N_29917,N_29923);
xnor UO_1015 (O_1015,N_29894,N_29816);
nor UO_1016 (O_1016,N_29891,N_29850);
and UO_1017 (O_1017,N_29821,N_29980);
nand UO_1018 (O_1018,N_29971,N_29876);
nand UO_1019 (O_1019,N_29806,N_29942);
and UO_1020 (O_1020,N_29860,N_29971);
nand UO_1021 (O_1021,N_29974,N_29932);
xnor UO_1022 (O_1022,N_29935,N_29962);
nand UO_1023 (O_1023,N_29942,N_29951);
xnor UO_1024 (O_1024,N_29916,N_29929);
nor UO_1025 (O_1025,N_29884,N_29853);
nor UO_1026 (O_1026,N_29864,N_29943);
nand UO_1027 (O_1027,N_29878,N_29914);
xor UO_1028 (O_1028,N_29801,N_29883);
nand UO_1029 (O_1029,N_29846,N_29810);
xor UO_1030 (O_1030,N_29959,N_29889);
nand UO_1031 (O_1031,N_29976,N_29957);
nand UO_1032 (O_1032,N_29852,N_29983);
and UO_1033 (O_1033,N_29962,N_29941);
and UO_1034 (O_1034,N_29979,N_29896);
xor UO_1035 (O_1035,N_29907,N_29941);
xnor UO_1036 (O_1036,N_29814,N_29975);
and UO_1037 (O_1037,N_29938,N_29970);
or UO_1038 (O_1038,N_29927,N_29983);
and UO_1039 (O_1039,N_29807,N_29859);
nand UO_1040 (O_1040,N_29987,N_29935);
and UO_1041 (O_1041,N_29941,N_29815);
nor UO_1042 (O_1042,N_29976,N_29900);
xor UO_1043 (O_1043,N_29831,N_29920);
xor UO_1044 (O_1044,N_29901,N_29846);
xor UO_1045 (O_1045,N_29855,N_29901);
xor UO_1046 (O_1046,N_29958,N_29898);
nand UO_1047 (O_1047,N_29944,N_29831);
nand UO_1048 (O_1048,N_29802,N_29910);
and UO_1049 (O_1049,N_29855,N_29948);
nor UO_1050 (O_1050,N_29866,N_29826);
nand UO_1051 (O_1051,N_29909,N_29991);
nor UO_1052 (O_1052,N_29995,N_29892);
nor UO_1053 (O_1053,N_29835,N_29918);
nor UO_1054 (O_1054,N_29871,N_29838);
or UO_1055 (O_1055,N_29895,N_29838);
nand UO_1056 (O_1056,N_29913,N_29880);
and UO_1057 (O_1057,N_29865,N_29911);
or UO_1058 (O_1058,N_29874,N_29906);
and UO_1059 (O_1059,N_29893,N_29983);
nand UO_1060 (O_1060,N_29858,N_29942);
or UO_1061 (O_1061,N_29939,N_29948);
xnor UO_1062 (O_1062,N_29960,N_29907);
xor UO_1063 (O_1063,N_29889,N_29987);
and UO_1064 (O_1064,N_29993,N_29856);
nand UO_1065 (O_1065,N_29972,N_29827);
or UO_1066 (O_1066,N_29965,N_29825);
nor UO_1067 (O_1067,N_29902,N_29883);
nor UO_1068 (O_1068,N_29971,N_29975);
nor UO_1069 (O_1069,N_29836,N_29950);
nand UO_1070 (O_1070,N_29821,N_29823);
or UO_1071 (O_1071,N_29977,N_29875);
xor UO_1072 (O_1072,N_29963,N_29855);
and UO_1073 (O_1073,N_29922,N_29866);
nor UO_1074 (O_1074,N_29810,N_29841);
xnor UO_1075 (O_1075,N_29844,N_29863);
and UO_1076 (O_1076,N_29931,N_29971);
and UO_1077 (O_1077,N_29900,N_29820);
nor UO_1078 (O_1078,N_29848,N_29898);
xnor UO_1079 (O_1079,N_29834,N_29900);
nor UO_1080 (O_1080,N_29883,N_29856);
xnor UO_1081 (O_1081,N_29882,N_29827);
nand UO_1082 (O_1082,N_29819,N_29809);
nand UO_1083 (O_1083,N_29887,N_29839);
or UO_1084 (O_1084,N_29820,N_29945);
nor UO_1085 (O_1085,N_29844,N_29964);
or UO_1086 (O_1086,N_29952,N_29955);
xor UO_1087 (O_1087,N_29991,N_29969);
and UO_1088 (O_1088,N_29810,N_29948);
nor UO_1089 (O_1089,N_29894,N_29896);
xor UO_1090 (O_1090,N_29850,N_29844);
and UO_1091 (O_1091,N_29964,N_29843);
nand UO_1092 (O_1092,N_29958,N_29824);
xnor UO_1093 (O_1093,N_29850,N_29912);
nand UO_1094 (O_1094,N_29923,N_29937);
or UO_1095 (O_1095,N_29985,N_29895);
xnor UO_1096 (O_1096,N_29957,N_29921);
nand UO_1097 (O_1097,N_29979,N_29982);
and UO_1098 (O_1098,N_29870,N_29998);
nor UO_1099 (O_1099,N_29962,N_29828);
nor UO_1100 (O_1100,N_29989,N_29901);
nand UO_1101 (O_1101,N_29865,N_29972);
nor UO_1102 (O_1102,N_29812,N_29921);
nor UO_1103 (O_1103,N_29979,N_29949);
and UO_1104 (O_1104,N_29807,N_29967);
xor UO_1105 (O_1105,N_29955,N_29861);
or UO_1106 (O_1106,N_29845,N_29969);
xnor UO_1107 (O_1107,N_29809,N_29981);
nand UO_1108 (O_1108,N_29906,N_29931);
nor UO_1109 (O_1109,N_29807,N_29943);
or UO_1110 (O_1110,N_29953,N_29951);
xor UO_1111 (O_1111,N_29816,N_29950);
nor UO_1112 (O_1112,N_29869,N_29968);
and UO_1113 (O_1113,N_29856,N_29891);
or UO_1114 (O_1114,N_29939,N_29895);
nor UO_1115 (O_1115,N_29936,N_29913);
nand UO_1116 (O_1116,N_29902,N_29862);
nand UO_1117 (O_1117,N_29948,N_29816);
nor UO_1118 (O_1118,N_29938,N_29812);
nand UO_1119 (O_1119,N_29911,N_29967);
nor UO_1120 (O_1120,N_29808,N_29859);
xnor UO_1121 (O_1121,N_29976,N_29985);
nand UO_1122 (O_1122,N_29843,N_29878);
and UO_1123 (O_1123,N_29942,N_29833);
nor UO_1124 (O_1124,N_29948,N_29936);
and UO_1125 (O_1125,N_29914,N_29850);
xnor UO_1126 (O_1126,N_29938,N_29940);
nand UO_1127 (O_1127,N_29815,N_29902);
or UO_1128 (O_1128,N_29867,N_29840);
or UO_1129 (O_1129,N_29815,N_29868);
nor UO_1130 (O_1130,N_29849,N_29881);
and UO_1131 (O_1131,N_29978,N_29984);
or UO_1132 (O_1132,N_29985,N_29949);
nand UO_1133 (O_1133,N_29803,N_29896);
nor UO_1134 (O_1134,N_29814,N_29992);
or UO_1135 (O_1135,N_29976,N_29908);
or UO_1136 (O_1136,N_29920,N_29967);
nor UO_1137 (O_1137,N_29880,N_29990);
nand UO_1138 (O_1138,N_29969,N_29945);
xor UO_1139 (O_1139,N_29868,N_29895);
or UO_1140 (O_1140,N_29943,N_29939);
nor UO_1141 (O_1141,N_29834,N_29979);
nand UO_1142 (O_1142,N_29924,N_29830);
nor UO_1143 (O_1143,N_29923,N_29999);
nand UO_1144 (O_1144,N_29853,N_29933);
nor UO_1145 (O_1145,N_29801,N_29855);
or UO_1146 (O_1146,N_29838,N_29962);
xor UO_1147 (O_1147,N_29811,N_29869);
and UO_1148 (O_1148,N_29925,N_29906);
nor UO_1149 (O_1149,N_29827,N_29843);
or UO_1150 (O_1150,N_29938,N_29897);
xor UO_1151 (O_1151,N_29832,N_29813);
nor UO_1152 (O_1152,N_29894,N_29839);
or UO_1153 (O_1153,N_29863,N_29864);
nor UO_1154 (O_1154,N_29809,N_29949);
xnor UO_1155 (O_1155,N_29908,N_29902);
or UO_1156 (O_1156,N_29827,N_29872);
or UO_1157 (O_1157,N_29890,N_29956);
nand UO_1158 (O_1158,N_29836,N_29975);
nor UO_1159 (O_1159,N_29991,N_29995);
nor UO_1160 (O_1160,N_29897,N_29802);
nand UO_1161 (O_1161,N_29923,N_29804);
xor UO_1162 (O_1162,N_29852,N_29854);
and UO_1163 (O_1163,N_29954,N_29942);
or UO_1164 (O_1164,N_29839,N_29997);
xnor UO_1165 (O_1165,N_29980,N_29930);
and UO_1166 (O_1166,N_29830,N_29941);
or UO_1167 (O_1167,N_29826,N_29907);
nand UO_1168 (O_1168,N_29953,N_29896);
xor UO_1169 (O_1169,N_29899,N_29852);
or UO_1170 (O_1170,N_29876,N_29929);
nand UO_1171 (O_1171,N_29839,N_29998);
xnor UO_1172 (O_1172,N_29865,N_29840);
and UO_1173 (O_1173,N_29881,N_29939);
nor UO_1174 (O_1174,N_29861,N_29938);
and UO_1175 (O_1175,N_29969,N_29884);
and UO_1176 (O_1176,N_29885,N_29813);
nor UO_1177 (O_1177,N_29945,N_29800);
or UO_1178 (O_1178,N_29829,N_29992);
nor UO_1179 (O_1179,N_29974,N_29846);
or UO_1180 (O_1180,N_29831,N_29960);
nor UO_1181 (O_1181,N_29989,N_29825);
nor UO_1182 (O_1182,N_29997,N_29838);
xor UO_1183 (O_1183,N_29946,N_29944);
and UO_1184 (O_1184,N_29806,N_29877);
xnor UO_1185 (O_1185,N_29826,N_29986);
nor UO_1186 (O_1186,N_29870,N_29898);
nor UO_1187 (O_1187,N_29946,N_29818);
xnor UO_1188 (O_1188,N_29951,N_29983);
and UO_1189 (O_1189,N_29986,N_29904);
or UO_1190 (O_1190,N_29879,N_29816);
nor UO_1191 (O_1191,N_29812,N_29918);
nor UO_1192 (O_1192,N_29829,N_29845);
and UO_1193 (O_1193,N_29831,N_29978);
nor UO_1194 (O_1194,N_29946,N_29860);
xor UO_1195 (O_1195,N_29963,N_29845);
xnor UO_1196 (O_1196,N_29892,N_29947);
nand UO_1197 (O_1197,N_29823,N_29922);
nand UO_1198 (O_1198,N_29874,N_29938);
nor UO_1199 (O_1199,N_29826,N_29956);
xor UO_1200 (O_1200,N_29870,N_29991);
or UO_1201 (O_1201,N_29933,N_29975);
xnor UO_1202 (O_1202,N_29812,N_29882);
or UO_1203 (O_1203,N_29992,N_29879);
xor UO_1204 (O_1204,N_29996,N_29935);
nor UO_1205 (O_1205,N_29910,N_29929);
nand UO_1206 (O_1206,N_29885,N_29984);
nor UO_1207 (O_1207,N_29973,N_29969);
nor UO_1208 (O_1208,N_29881,N_29931);
or UO_1209 (O_1209,N_29947,N_29811);
and UO_1210 (O_1210,N_29960,N_29826);
nor UO_1211 (O_1211,N_29919,N_29959);
nand UO_1212 (O_1212,N_29994,N_29816);
nor UO_1213 (O_1213,N_29887,N_29985);
xor UO_1214 (O_1214,N_29889,N_29909);
and UO_1215 (O_1215,N_29835,N_29907);
xnor UO_1216 (O_1216,N_29890,N_29957);
xnor UO_1217 (O_1217,N_29946,N_29849);
xor UO_1218 (O_1218,N_29903,N_29930);
nand UO_1219 (O_1219,N_29875,N_29852);
and UO_1220 (O_1220,N_29802,N_29992);
or UO_1221 (O_1221,N_29950,N_29827);
nand UO_1222 (O_1222,N_29973,N_29857);
xor UO_1223 (O_1223,N_29939,N_29839);
xnor UO_1224 (O_1224,N_29856,N_29997);
nand UO_1225 (O_1225,N_29948,N_29990);
nor UO_1226 (O_1226,N_29852,N_29877);
or UO_1227 (O_1227,N_29849,N_29948);
and UO_1228 (O_1228,N_29875,N_29902);
or UO_1229 (O_1229,N_29920,N_29970);
nor UO_1230 (O_1230,N_29883,N_29849);
nand UO_1231 (O_1231,N_29833,N_29925);
or UO_1232 (O_1232,N_29839,N_29823);
xor UO_1233 (O_1233,N_29919,N_29805);
and UO_1234 (O_1234,N_29890,N_29840);
nand UO_1235 (O_1235,N_29869,N_29860);
or UO_1236 (O_1236,N_29811,N_29919);
and UO_1237 (O_1237,N_29821,N_29860);
nand UO_1238 (O_1238,N_29897,N_29972);
nor UO_1239 (O_1239,N_29861,N_29868);
and UO_1240 (O_1240,N_29807,N_29874);
nor UO_1241 (O_1241,N_29925,N_29826);
and UO_1242 (O_1242,N_29992,N_29871);
nor UO_1243 (O_1243,N_29911,N_29916);
xnor UO_1244 (O_1244,N_29986,N_29880);
nand UO_1245 (O_1245,N_29868,N_29874);
nand UO_1246 (O_1246,N_29913,N_29929);
and UO_1247 (O_1247,N_29890,N_29838);
nand UO_1248 (O_1248,N_29878,N_29810);
xnor UO_1249 (O_1249,N_29808,N_29987);
or UO_1250 (O_1250,N_29827,N_29814);
xnor UO_1251 (O_1251,N_29973,N_29948);
xnor UO_1252 (O_1252,N_29801,N_29928);
xor UO_1253 (O_1253,N_29841,N_29959);
nand UO_1254 (O_1254,N_29985,N_29840);
xor UO_1255 (O_1255,N_29908,N_29868);
nand UO_1256 (O_1256,N_29812,N_29980);
and UO_1257 (O_1257,N_29968,N_29947);
nand UO_1258 (O_1258,N_29989,N_29940);
nand UO_1259 (O_1259,N_29865,N_29963);
or UO_1260 (O_1260,N_29995,N_29878);
xnor UO_1261 (O_1261,N_29831,N_29804);
nor UO_1262 (O_1262,N_29958,N_29829);
or UO_1263 (O_1263,N_29804,N_29875);
xor UO_1264 (O_1264,N_29923,N_29901);
xnor UO_1265 (O_1265,N_29970,N_29952);
nor UO_1266 (O_1266,N_29864,N_29880);
xor UO_1267 (O_1267,N_29958,N_29942);
or UO_1268 (O_1268,N_29855,N_29941);
and UO_1269 (O_1269,N_29979,N_29832);
and UO_1270 (O_1270,N_29863,N_29821);
nand UO_1271 (O_1271,N_29923,N_29924);
xnor UO_1272 (O_1272,N_29982,N_29888);
xnor UO_1273 (O_1273,N_29876,N_29996);
nor UO_1274 (O_1274,N_29968,N_29840);
nor UO_1275 (O_1275,N_29856,N_29929);
or UO_1276 (O_1276,N_29940,N_29976);
or UO_1277 (O_1277,N_29884,N_29925);
and UO_1278 (O_1278,N_29824,N_29825);
nand UO_1279 (O_1279,N_29810,N_29827);
xor UO_1280 (O_1280,N_29853,N_29859);
xnor UO_1281 (O_1281,N_29812,N_29940);
and UO_1282 (O_1282,N_29924,N_29845);
and UO_1283 (O_1283,N_29830,N_29954);
nor UO_1284 (O_1284,N_29875,N_29842);
or UO_1285 (O_1285,N_29921,N_29977);
nand UO_1286 (O_1286,N_29904,N_29974);
and UO_1287 (O_1287,N_29874,N_29983);
nand UO_1288 (O_1288,N_29962,N_29931);
and UO_1289 (O_1289,N_29848,N_29847);
nor UO_1290 (O_1290,N_29828,N_29819);
nor UO_1291 (O_1291,N_29951,N_29898);
or UO_1292 (O_1292,N_29974,N_29811);
xor UO_1293 (O_1293,N_29921,N_29967);
or UO_1294 (O_1294,N_29993,N_29952);
and UO_1295 (O_1295,N_29954,N_29846);
nor UO_1296 (O_1296,N_29915,N_29863);
nand UO_1297 (O_1297,N_29902,N_29800);
xor UO_1298 (O_1298,N_29941,N_29919);
and UO_1299 (O_1299,N_29915,N_29902);
and UO_1300 (O_1300,N_29829,N_29800);
nor UO_1301 (O_1301,N_29905,N_29899);
nand UO_1302 (O_1302,N_29878,N_29935);
nor UO_1303 (O_1303,N_29944,N_29931);
xnor UO_1304 (O_1304,N_29864,N_29900);
and UO_1305 (O_1305,N_29814,N_29908);
nand UO_1306 (O_1306,N_29813,N_29805);
xor UO_1307 (O_1307,N_29863,N_29930);
nand UO_1308 (O_1308,N_29807,N_29992);
nand UO_1309 (O_1309,N_29838,N_29911);
and UO_1310 (O_1310,N_29821,N_29991);
or UO_1311 (O_1311,N_29939,N_29823);
xor UO_1312 (O_1312,N_29978,N_29822);
and UO_1313 (O_1313,N_29957,N_29914);
or UO_1314 (O_1314,N_29979,N_29831);
xnor UO_1315 (O_1315,N_29904,N_29962);
xnor UO_1316 (O_1316,N_29871,N_29856);
and UO_1317 (O_1317,N_29916,N_29997);
nor UO_1318 (O_1318,N_29870,N_29826);
nor UO_1319 (O_1319,N_29850,N_29857);
or UO_1320 (O_1320,N_29828,N_29866);
xor UO_1321 (O_1321,N_29919,N_29924);
nand UO_1322 (O_1322,N_29995,N_29963);
or UO_1323 (O_1323,N_29988,N_29870);
xnor UO_1324 (O_1324,N_29804,N_29858);
nor UO_1325 (O_1325,N_29954,N_29928);
nor UO_1326 (O_1326,N_29836,N_29951);
nand UO_1327 (O_1327,N_29820,N_29953);
nand UO_1328 (O_1328,N_29879,N_29829);
and UO_1329 (O_1329,N_29845,N_29921);
nor UO_1330 (O_1330,N_29853,N_29936);
nand UO_1331 (O_1331,N_29849,N_29874);
xnor UO_1332 (O_1332,N_29981,N_29974);
and UO_1333 (O_1333,N_29824,N_29851);
xnor UO_1334 (O_1334,N_29875,N_29968);
nor UO_1335 (O_1335,N_29998,N_29918);
nand UO_1336 (O_1336,N_29943,N_29812);
or UO_1337 (O_1337,N_29837,N_29915);
nor UO_1338 (O_1338,N_29826,N_29811);
xnor UO_1339 (O_1339,N_29910,N_29901);
nand UO_1340 (O_1340,N_29941,N_29884);
nand UO_1341 (O_1341,N_29800,N_29872);
xnor UO_1342 (O_1342,N_29883,N_29952);
xor UO_1343 (O_1343,N_29807,N_29926);
xnor UO_1344 (O_1344,N_29968,N_29997);
or UO_1345 (O_1345,N_29966,N_29973);
and UO_1346 (O_1346,N_29813,N_29934);
xor UO_1347 (O_1347,N_29996,N_29929);
nand UO_1348 (O_1348,N_29949,N_29934);
and UO_1349 (O_1349,N_29843,N_29898);
or UO_1350 (O_1350,N_29945,N_29814);
nand UO_1351 (O_1351,N_29864,N_29805);
nor UO_1352 (O_1352,N_29824,N_29927);
nor UO_1353 (O_1353,N_29832,N_29848);
nor UO_1354 (O_1354,N_29967,N_29869);
and UO_1355 (O_1355,N_29999,N_29956);
and UO_1356 (O_1356,N_29904,N_29884);
xnor UO_1357 (O_1357,N_29958,N_29842);
nand UO_1358 (O_1358,N_29801,N_29898);
xor UO_1359 (O_1359,N_29878,N_29900);
nand UO_1360 (O_1360,N_29841,N_29988);
xor UO_1361 (O_1361,N_29924,N_29922);
xnor UO_1362 (O_1362,N_29848,N_29840);
xnor UO_1363 (O_1363,N_29911,N_29827);
nand UO_1364 (O_1364,N_29959,N_29851);
nor UO_1365 (O_1365,N_29882,N_29857);
or UO_1366 (O_1366,N_29938,N_29815);
xnor UO_1367 (O_1367,N_29894,N_29994);
nand UO_1368 (O_1368,N_29926,N_29993);
nor UO_1369 (O_1369,N_29957,N_29986);
nor UO_1370 (O_1370,N_29992,N_29862);
nand UO_1371 (O_1371,N_29925,N_29993);
nor UO_1372 (O_1372,N_29883,N_29848);
and UO_1373 (O_1373,N_29845,N_29923);
and UO_1374 (O_1374,N_29865,N_29992);
xnor UO_1375 (O_1375,N_29861,N_29913);
and UO_1376 (O_1376,N_29809,N_29803);
xor UO_1377 (O_1377,N_29867,N_29988);
and UO_1378 (O_1378,N_29918,N_29959);
nand UO_1379 (O_1379,N_29816,N_29967);
nand UO_1380 (O_1380,N_29870,N_29999);
nand UO_1381 (O_1381,N_29923,N_29806);
or UO_1382 (O_1382,N_29830,N_29807);
nor UO_1383 (O_1383,N_29905,N_29925);
or UO_1384 (O_1384,N_29892,N_29931);
or UO_1385 (O_1385,N_29818,N_29890);
nand UO_1386 (O_1386,N_29835,N_29845);
nor UO_1387 (O_1387,N_29850,N_29889);
and UO_1388 (O_1388,N_29871,N_29848);
and UO_1389 (O_1389,N_29957,N_29950);
and UO_1390 (O_1390,N_29932,N_29985);
xor UO_1391 (O_1391,N_29944,N_29993);
nor UO_1392 (O_1392,N_29840,N_29921);
xor UO_1393 (O_1393,N_29974,N_29965);
or UO_1394 (O_1394,N_29831,N_29867);
nor UO_1395 (O_1395,N_29922,N_29863);
nor UO_1396 (O_1396,N_29997,N_29818);
xor UO_1397 (O_1397,N_29873,N_29804);
nor UO_1398 (O_1398,N_29819,N_29882);
nand UO_1399 (O_1399,N_29843,N_29952);
or UO_1400 (O_1400,N_29922,N_29860);
and UO_1401 (O_1401,N_29848,N_29949);
xor UO_1402 (O_1402,N_29961,N_29886);
nand UO_1403 (O_1403,N_29948,N_29863);
nand UO_1404 (O_1404,N_29904,N_29900);
nor UO_1405 (O_1405,N_29951,N_29815);
or UO_1406 (O_1406,N_29876,N_29830);
or UO_1407 (O_1407,N_29989,N_29924);
nor UO_1408 (O_1408,N_29953,N_29957);
xnor UO_1409 (O_1409,N_29974,N_29805);
or UO_1410 (O_1410,N_29922,N_29828);
or UO_1411 (O_1411,N_29838,N_29877);
nor UO_1412 (O_1412,N_29910,N_29889);
xnor UO_1413 (O_1413,N_29861,N_29851);
nor UO_1414 (O_1414,N_29978,N_29851);
or UO_1415 (O_1415,N_29877,N_29828);
nand UO_1416 (O_1416,N_29882,N_29988);
and UO_1417 (O_1417,N_29868,N_29988);
nand UO_1418 (O_1418,N_29822,N_29985);
xor UO_1419 (O_1419,N_29878,N_29894);
and UO_1420 (O_1420,N_29879,N_29898);
nor UO_1421 (O_1421,N_29923,N_29980);
nand UO_1422 (O_1422,N_29857,N_29972);
nand UO_1423 (O_1423,N_29815,N_29988);
and UO_1424 (O_1424,N_29992,N_29828);
xor UO_1425 (O_1425,N_29978,N_29898);
xnor UO_1426 (O_1426,N_29995,N_29900);
xnor UO_1427 (O_1427,N_29961,N_29982);
or UO_1428 (O_1428,N_29944,N_29865);
and UO_1429 (O_1429,N_29881,N_29973);
or UO_1430 (O_1430,N_29860,N_29839);
and UO_1431 (O_1431,N_29992,N_29872);
or UO_1432 (O_1432,N_29944,N_29941);
nand UO_1433 (O_1433,N_29925,N_29958);
and UO_1434 (O_1434,N_29845,N_29991);
or UO_1435 (O_1435,N_29917,N_29967);
nand UO_1436 (O_1436,N_29927,N_29986);
or UO_1437 (O_1437,N_29867,N_29872);
nand UO_1438 (O_1438,N_29868,N_29889);
or UO_1439 (O_1439,N_29882,N_29880);
or UO_1440 (O_1440,N_29876,N_29800);
and UO_1441 (O_1441,N_29912,N_29899);
xnor UO_1442 (O_1442,N_29879,N_29823);
or UO_1443 (O_1443,N_29810,N_29912);
and UO_1444 (O_1444,N_29844,N_29992);
and UO_1445 (O_1445,N_29919,N_29897);
nand UO_1446 (O_1446,N_29860,N_29890);
xor UO_1447 (O_1447,N_29882,N_29930);
xor UO_1448 (O_1448,N_29964,N_29839);
xor UO_1449 (O_1449,N_29905,N_29852);
nand UO_1450 (O_1450,N_29896,N_29836);
xnor UO_1451 (O_1451,N_29841,N_29901);
nor UO_1452 (O_1452,N_29854,N_29925);
xnor UO_1453 (O_1453,N_29927,N_29893);
xnor UO_1454 (O_1454,N_29872,N_29877);
and UO_1455 (O_1455,N_29823,N_29800);
nor UO_1456 (O_1456,N_29863,N_29816);
nand UO_1457 (O_1457,N_29859,N_29928);
and UO_1458 (O_1458,N_29812,N_29932);
or UO_1459 (O_1459,N_29871,N_29964);
and UO_1460 (O_1460,N_29849,N_29978);
xor UO_1461 (O_1461,N_29991,N_29928);
or UO_1462 (O_1462,N_29900,N_29812);
nand UO_1463 (O_1463,N_29874,N_29832);
xnor UO_1464 (O_1464,N_29857,N_29807);
nor UO_1465 (O_1465,N_29931,N_29835);
and UO_1466 (O_1466,N_29921,N_29958);
and UO_1467 (O_1467,N_29839,N_29803);
and UO_1468 (O_1468,N_29859,N_29975);
or UO_1469 (O_1469,N_29806,N_29980);
nand UO_1470 (O_1470,N_29935,N_29960);
nand UO_1471 (O_1471,N_29843,N_29989);
nor UO_1472 (O_1472,N_29959,N_29970);
and UO_1473 (O_1473,N_29968,N_29976);
nand UO_1474 (O_1474,N_29837,N_29863);
or UO_1475 (O_1475,N_29897,N_29850);
nor UO_1476 (O_1476,N_29819,N_29874);
and UO_1477 (O_1477,N_29977,N_29870);
or UO_1478 (O_1478,N_29952,N_29984);
or UO_1479 (O_1479,N_29800,N_29834);
nand UO_1480 (O_1480,N_29852,N_29967);
nor UO_1481 (O_1481,N_29935,N_29874);
nand UO_1482 (O_1482,N_29804,N_29980);
and UO_1483 (O_1483,N_29988,N_29902);
xor UO_1484 (O_1484,N_29811,N_29914);
nand UO_1485 (O_1485,N_29817,N_29802);
and UO_1486 (O_1486,N_29983,N_29870);
xnor UO_1487 (O_1487,N_29916,N_29953);
and UO_1488 (O_1488,N_29903,N_29926);
or UO_1489 (O_1489,N_29919,N_29994);
nand UO_1490 (O_1490,N_29878,N_29999);
nor UO_1491 (O_1491,N_29987,N_29859);
nand UO_1492 (O_1492,N_29910,N_29932);
xor UO_1493 (O_1493,N_29803,N_29825);
and UO_1494 (O_1494,N_29899,N_29956);
or UO_1495 (O_1495,N_29962,N_29910);
xnor UO_1496 (O_1496,N_29855,N_29907);
and UO_1497 (O_1497,N_29891,N_29920);
or UO_1498 (O_1498,N_29988,N_29906);
or UO_1499 (O_1499,N_29830,N_29889);
xnor UO_1500 (O_1500,N_29870,N_29804);
or UO_1501 (O_1501,N_29926,N_29944);
xnor UO_1502 (O_1502,N_29859,N_29961);
and UO_1503 (O_1503,N_29903,N_29838);
nand UO_1504 (O_1504,N_29984,N_29946);
nand UO_1505 (O_1505,N_29853,N_29800);
nand UO_1506 (O_1506,N_29865,N_29812);
or UO_1507 (O_1507,N_29816,N_29924);
xor UO_1508 (O_1508,N_29992,N_29981);
nand UO_1509 (O_1509,N_29905,N_29933);
nor UO_1510 (O_1510,N_29967,N_29964);
or UO_1511 (O_1511,N_29857,N_29996);
nand UO_1512 (O_1512,N_29950,N_29888);
nor UO_1513 (O_1513,N_29999,N_29983);
xnor UO_1514 (O_1514,N_29874,N_29985);
xor UO_1515 (O_1515,N_29824,N_29913);
and UO_1516 (O_1516,N_29916,N_29961);
nor UO_1517 (O_1517,N_29856,N_29973);
and UO_1518 (O_1518,N_29844,N_29988);
nand UO_1519 (O_1519,N_29842,N_29807);
xor UO_1520 (O_1520,N_29973,N_29906);
and UO_1521 (O_1521,N_29866,N_29847);
nand UO_1522 (O_1522,N_29811,N_29870);
xnor UO_1523 (O_1523,N_29925,N_29835);
or UO_1524 (O_1524,N_29829,N_29990);
or UO_1525 (O_1525,N_29964,N_29912);
or UO_1526 (O_1526,N_29840,N_29826);
or UO_1527 (O_1527,N_29876,N_29850);
nor UO_1528 (O_1528,N_29953,N_29959);
nand UO_1529 (O_1529,N_29817,N_29801);
xnor UO_1530 (O_1530,N_29851,N_29886);
xor UO_1531 (O_1531,N_29960,N_29963);
nand UO_1532 (O_1532,N_29947,N_29920);
xnor UO_1533 (O_1533,N_29954,N_29876);
nand UO_1534 (O_1534,N_29813,N_29811);
nand UO_1535 (O_1535,N_29883,N_29843);
nand UO_1536 (O_1536,N_29906,N_29852);
nor UO_1537 (O_1537,N_29885,N_29815);
or UO_1538 (O_1538,N_29854,N_29993);
or UO_1539 (O_1539,N_29945,N_29876);
xnor UO_1540 (O_1540,N_29938,N_29895);
and UO_1541 (O_1541,N_29923,N_29906);
nor UO_1542 (O_1542,N_29882,N_29884);
xnor UO_1543 (O_1543,N_29987,N_29945);
nor UO_1544 (O_1544,N_29832,N_29837);
and UO_1545 (O_1545,N_29839,N_29968);
or UO_1546 (O_1546,N_29936,N_29911);
and UO_1547 (O_1547,N_29869,N_29800);
and UO_1548 (O_1548,N_29959,N_29832);
and UO_1549 (O_1549,N_29868,N_29946);
nor UO_1550 (O_1550,N_29892,N_29990);
nor UO_1551 (O_1551,N_29855,N_29804);
nor UO_1552 (O_1552,N_29824,N_29978);
xnor UO_1553 (O_1553,N_29835,N_29864);
or UO_1554 (O_1554,N_29824,N_29896);
nor UO_1555 (O_1555,N_29981,N_29836);
or UO_1556 (O_1556,N_29968,N_29949);
nor UO_1557 (O_1557,N_29867,N_29924);
nor UO_1558 (O_1558,N_29844,N_29848);
xnor UO_1559 (O_1559,N_29935,N_29917);
nand UO_1560 (O_1560,N_29943,N_29913);
nor UO_1561 (O_1561,N_29803,N_29991);
or UO_1562 (O_1562,N_29950,N_29843);
xor UO_1563 (O_1563,N_29972,N_29910);
xnor UO_1564 (O_1564,N_29858,N_29861);
or UO_1565 (O_1565,N_29900,N_29849);
nand UO_1566 (O_1566,N_29986,N_29942);
or UO_1567 (O_1567,N_29965,N_29989);
xor UO_1568 (O_1568,N_29849,N_29878);
xnor UO_1569 (O_1569,N_29848,N_29946);
xnor UO_1570 (O_1570,N_29989,N_29973);
nor UO_1571 (O_1571,N_29985,N_29988);
xor UO_1572 (O_1572,N_29807,N_29825);
nor UO_1573 (O_1573,N_29988,N_29805);
and UO_1574 (O_1574,N_29967,N_29985);
and UO_1575 (O_1575,N_29868,N_29912);
nor UO_1576 (O_1576,N_29830,N_29946);
xor UO_1577 (O_1577,N_29922,N_29902);
and UO_1578 (O_1578,N_29860,N_29838);
nor UO_1579 (O_1579,N_29977,N_29990);
and UO_1580 (O_1580,N_29917,N_29997);
nor UO_1581 (O_1581,N_29889,N_29929);
xor UO_1582 (O_1582,N_29979,N_29940);
nand UO_1583 (O_1583,N_29979,N_29942);
nand UO_1584 (O_1584,N_29811,N_29829);
xor UO_1585 (O_1585,N_29947,N_29907);
xnor UO_1586 (O_1586,N_29858,N_29964);
nand UO_1587 (O_1587,N_29854,N_29836);
nand UO_1588 (O_1588,N_29808,N_29804);
nand UO_1589 (O_1589,N_29816,N_29940);
and UO_1590 (O_1590,N_29898,N_29857);
xnor UO_1591 (O_1591,N_29955,N_29908);
xor UO_1592 (O_1592,N_29986,N_29960);
xor UO_1593 (O_1593,N_29865,N_29805);
and UO_1594 (O_1594,N_29941,N_29864);
and UO_1595 (O_1595,N_29982,N_29810);
nand UO_1596 (O_1596,N_29806,N_29930);
nor UO_1597 (O_1597,N_29821,N_29950);
and UO_1598 (O_1598,N_29833,N_29823);
xnor UO_1599 (O_1599,N_29844,N_29810);
or UO_1600 (O_1600,N_29839,N_29971);
nor UO_1601 (O_1601,N_29886,N_29940);
nand UO_1602 (O_1602,N_29987,N_29920);
nor UO_1603 (O_1603,N_29924,N_29930);
nor UO_1604 (O_1604,N_29900,N_29907);
nor UO_1605 (O_1605,N_29954,N_29995);
nor UO_1606 (O_1606,N_29922,N_29862);
or UO_1607 (O_1607,N_29948,N_29926);
and UO_1608 (O_1608,N_29905,N_29913);
nand UO_1609 (O_1609,N_29842,N_29803);
nor UO_1610 (O_1610,N_29942,N_29946);
xnor UO_1611 (O_1611,N_29881,N_29974);
nand UO_1612 (O_1612,N_29863,N_29897);
or UO_1613 (O_1613,N_29974,N_29995);
nor UO_1614 (O_1614,N_29832,N_29833);
and UO_1615 (O_1615,N_29949,N_29836);
or UO_1616 (O_1616,N_29997,N_29871);
nand UO_1617 (O_1617,N_29840,N_29843);
and UO_1618 (O_1618,N_29820,N_29862);
and UO_1619 (O_1619,N_29827,N_29821);
nand UO_1620 (O_1620,N_29940,N_29871);
xor UO_1621 (O_1621,N_29813,N_29825);
nand UO_1622 (O_1622,N_29816,N_29878);
nand UO_1623 (O_1623,N_29819,N_29807);
or UO_1624 (O_1624,N_29873,N_29825);
and UO_1625 (O_1625,N_29947,N_29887);
xnor UO_1626 (O_1626,N_29918,N_29956);
nand UO_1627 (O_1627,N_29879,N_29947);
xor UO_1628 (O_1628,N_29863,N_29929);
xnor UO_1629 (O_1629,N_29857,N_29874);
and UO_1630 (O_1630,N_29907,N_29839);
nor UO_1631 (O_1631,N_29813,N_29904);
xnor UO_1632 (O_1632,N_29934,N_29935);
xor UO_1633 (O_1633,N_29905,N_29961);
and UO_1634 (O_1634,N_29928,N_29999);
or UO_1635 (O_1635,N_29847,N_29970);
xor UO_1636 (O_1636,N_29915,N_29849);
nand UO_1637 (O_1637,N_29874,N_29943);
and UO_1638 (O_1638,N_29823,N_29955);
nand UO_1639 (O_1639,N_29838,N_29981);
or UO_1640 (O_1640,N_29810,N_29954);
nor UO_1641 (O_1641,N_29869,N_29924);
xor UO_1642 (O_1642,N_29890,N_29904);
and UO_1643 (O_1643,N_29828,N_29964);
and UO_1644 (O_1644,N_29877,N_29880);
xor UO_1645 (O_1645,N_29889,N_29938);
nor UO_1646 (O_1646,N_29805,N_29984);
nand UO_1647 (O_1647,N_29882,N_29897);
nor UO_1648 (O_1648,N_29845,N_29851);
nor UO_1649 (O_1649,N_29937,N_29849);
nor UO_1650 (O_1650,N_29841,N_29911);
nand UO_1651 (O_1651,N_29981,N_29920);
and UO_1652 (O_1652,N_29869,N_29945);
nand UO_1653 (O_1653,N_29949,N_29869);
nand UO_1654 (O_1654,N_29995,N_29883);
nor UO_1655 (O_1655,N_29908,N_29818);
xor UO_1656 (O_1656,N_29986,N_29850);
or UO_1657 (O_1657,N_29975,N_29876);
and UO_1658 (O_1658,N_29951,N_29912);
and UO_1659 (O_1659,N_29927,N_29817);
xnor UO_1660 (O_1660,N_29959,N_29895);
nand UO_1661 (O_1661,N_29917,N_29982);
nor UO_1662 (O_1662,N_29887,N_29966);
and UO_1663 (O_1663,N_29921,N_29872);
nand UO_1664 (O_1664,N_29905,N_29907);
nand UO_1665 (O_1665,N_29906,N_29956);
xnor UO_1666 (O_1666,N_29824,N_29868);
and UO_1667 (O_1667,N_29907,N_29939);
xnor UO_1668 (O_1668,N_29956,N_29941);
or UO_1669 (O_1669,N_29864,N_29802);
xnor UO_1670 (O_1670,N_29895,N_29861);
nand UO_1671 (O_1671,N_29971,N_29912);
nand UO_1672 (O_1672,N_29835,N_29828);
xor UO_1673 (O_1673,N_29887,N_29878);
or UO_1674 (O_1674,N_29884,N_29986);
and UO_1675 (O_1675,N_29845,N_29908);
xnor UO_1676 (O_1676,N_29891,N_29931);
nand UO_1677 (O_1677,N_29983,N_29946);
and UO_1678 (O_1678,N_29825,N_29895);
or UO_1679 (O_1679,N_29803,N_29996);
nand UO_1680 (O_1680,N_29916,N_29856);
nand UO_1681 (O_1681,N_29938,N_29906);
xor UO_1682 (O_1682,N_29973,N_29985);
nand UO_1683 (O_1683,N_29901,N_29883);
nand UO_1684 (O_1684,N_29843,N_29894);
xor UO_1685 (O_1685,N_29814,N_29889);
xnor UO_1686 (O_1686,N_29952,N_29995);
and UO_1687 (O_1687,N_29845,N_29889);
nand UO_1688 (O_1688,N_29880,N_29922);
nand UO_1689 (O_1689,N_29926,N_29935);
xor UO_1690 (O_1690,N_29947,N_29994);
and UO_1691 (O_1691,N_29904,N_29987);
nor UO_1692 (O_1692,N_29917,N_29953);
nor UO_1693 (O_1693,N_29981,N_29907);
xnor UO_1694 (O_1694,N_29919,N_29815);
xor UO_1695 (O_1695,N_29836,N_29884);
and UO_1696 (O_1696,N_29927,N_29918);
or UO_1697 (O_1697,N_29880,N_29839);
nor UO_1698 (O_1698,N_29835,N_29962);
nand UO_1699 (O_1699,N_29808,N_29815);
nor UO_1700 (O_1700,N_29941,N_29955);
or UO_1701 (O_1701,N_29964,N_29902);
or UO_1702 (O_1702,N_29908,N_29854);
nor UO_1703 (O_1703,N_29961,N_29834);
nor UO_1704 (O_1704,N_29971,N_29960);
nand UO_1705 (O_1705,N_29855,N_29885);
xnor UO_1706 (O_1706,N_29953,N_29835);
or UO_1707 (O_1707,N_29835,N_29974);
or UO_1708 (O_1708,N_29894,N_29995);
or UO_1709 (O_1709,N_29962,N_29827);
or UO_1710 (O_1710,N_29963,N_29957);
and UO_1711 (O_1711,N_29980,N_29891);
nor UO_1712 (O_1712,N_29846,N_29922);
xor UO_1713 (O_1713,N_29830,N_29939);
nand UO_1714 (O_1714,N_29897,N_29878);
or UO_1715 (O_1715,N_29909,N_29977);
or UO_1716 (O_1716,N_29852,N_29968);
and UO_1717 (O_1717,N_29898,N_29811);
or UO_1718 (O_1718,N_29930,N_29932);
or UO_1719 (O_1719,N_29862,N_29974);
xnor UO_1720 (O_1720,N_29881,N_29860);
nor UO_1721 (O_1721,N_29822,N_29940);
or UO_1722 (O_1722,N_29979,N_29929);
nor UO_1723 (O_1723,N_29911,N_29842);
or UO_1724 (O_1724,N_29811,N_29955);
xnor UO_1725 (O_1725,N_29820,N_29872);
nand UO_1726 (O_1726,N_29942,N_29802);
or UO_1727 (O_1727,N_29890,N_29964);
nand UO_1728 (O_1728,N_29970,N_29882);
and UO_1729 (O_1729,N_29879,N_29959);
or UO_1730 (O_1730,N_29917,N_29965);
xnor UO_1731 (O_1731,N_29814,N_29811);
xor UO_1732 (O_1732,N_29951,N_29835);
nand UO_1733 (O_1733,N_29890,N_29968);
nand UO_1734 (O_1734,N_29833,N_29831);
or UO_1735 (O_1735,N_29822,N_29918);
nor UO_1736 (O_1736,N_29808,N_29966);
nand UO_1737 (O_1737,N_29825,N_29913);
nand UO_1738 (O_1738,N_29980,N_29925);
xnor UO_1739 (O_1739,N_29844,N_29873);
nor UO_1740 (O_1740,N_29807,N_29893);
xor UO_1741 (O_1741,N_29856,N_29915);
nand UO_1742 (O_1742,N_29805,N_29947);
xnor UO_1743 (O_1743,N_29927,N_29978);
nand UO_1744 (O_1744,N_29883,N_29831);
xor UO_1745 (O_1745,N_29831,N_29805);
or UO_1746 (O_1746,N_29891,N_29923);
nand UO_1747 (O_1747,N_29889,N_29864);
and UO_1748 (O_1748,N_29996,N_29861);
or UO_1749 (O_1749,N_29824,N_29990);
nor UO_1750 (O_1750,N_29814,N_29809);
xnor UO_1751 (O_1751,N_29942,N_29973);
and UO_1752 (O_1752,N_29968,N_29882);
or UO_1753 (O_1753,N_29829,N_29809);
nor UO_1754 (O_1754,N_29957,N_29933);
nor UO_1755 (O_1755,N_29994,N_29906);
xnor UO_1756 (O_1756,N_29962,N_29972);
xnor UO_1757 (O_1757,N_29973,N_29871);
xor UO_1758 (O_1758,N_29825,N_29988);
xnor UO_1759 (O_1759,N_29810,N_29963);
nor UO_1760 (O_1760,N_29824,N_29988);
nand UO_1761 (O_1761,N_29873,N_29942);
xnor UO_1762 (O_1762,N_29927,N_29816);
and UO_1763 (O_1763,N_29923,N_29913);
nand UO_1764 (O_1764,N_29955,N_29918);
and UO_1765 (O_1765,N_29948,N_29917);
and UO_1766 (O_1766,N_29927,N_29832);
and UO_1767 (O_1767,N_29993,N_29808);
xnor UO_1768 (O_1768,N_29839,N_29915);
xor UO_1769 (O_1769,N_29820,N_29850);
and UO_1770 (O_1770,N_29830,N_29922);
nand UO_1771 (O_1771,N_29912,N_29829);
xor UO_1772 (O_1772,N_29939,N_29926);
or UO_1773 (O_1773,N_29970,N_29928);
and UO_1774 (O_1774,N_29880,N_29861);
nand UO_1775 (O_1775,N_29848,N_29846);
nor UO_1776 (O_1776,N_29801,N_29937);
and UO_1777 (O_1777,N_29965,N_29841);
nand UO_1778 (O_1778,N_29956,N_29955);
and UO_1779 (O_1779,N_29886,N_29894);
xnor UO_1780 (O_1780,N_29800,N_29947);
nand UO_1781 (O_1781,N_29829,N_29836);
xor UO_1782 (O_1782,N_29862,N_29947);
and UO_1783 (O_1783,N_29832,N_29812);
or UO_1784 (O_1784,N_29888,N_29812);
xor UO_1785 (O_1785,N_29857,N_29956);
nor UO_1786 (O_1786,N_29918,N_29982);
and UO_1787 (O_1787,N_29847,N_29947);
and UO_1788 (O_1788,N_29992,N_29811);
xnor UO_1789 (O_1789,N_29916,N_29896);
and UO_1790 (O_1790,N_29911,N_29952);
xnor UO_1791 (O_1791,N_29858,N_29953);
nand UO_1792 (O_1792,N_29812,N_29846);
and UO_1793 (O_1793,N_29860,N_29974);
nand UO_1794 (O_1794,N_29999,N_29917);
and UO_1795 (O_1795,N_29888,N_29819);
xnor UO_1796 (O_1796,N_29853,N_29847);
or UO_1797 (O_1797,N_29801,N_29915);
or UO_1798 (O_1798,N_29936,N_29866);
xor UO_1799 (O_1799,N_29866,N_29938);
nand UO_1800 (O_1800,N_29985,N_29898);
nor UO_1801 (O_1801,N_29954,N_29975);
and UO_1802 (O_1802,N_29981,N_29814);
and UO_1803 (O_1803,N_29920,N_29849);
nor UO_1804 (O_1804,N_29843,N_29806);
xnor UO_1805 (O_1805,N_29980,N_29921);
or UO_1806 (O_1806,N_29921,N_29821);
nand UO_1807 (O_1807,N_29802,N_29851);
and UO_1808 (O_1808,N_29965,N_29901);
and UO_1809 (O_1809,N_29956,N_29868);
xor UO_1810 (O_1810,N_29853,N_29835);
and UO_1811 (O_1811,N_29929,N_29902);
or UO_1812 (O_1812,N_29816,N_29984);
xor UO_1813 (O_1813,N_29852,N_29885);
and UO_1814 (O_1814,N_29966,N_29843);
and UO_1815 (O_1815,N_29827,N_29959);
nor UO_1816 (O_1816,N_29937,N_29907);
and UO_1817 (O_1817,N_29878,N_29805);
xnor UO_1818 (O_1818,N_29944,N_29983);
or UO_1819 (O_1819,N_29990,N_29875);
nor UO_1820 (O_1820,N_29804,N_29900);
nor UO_1821 (O_1821,N_29862,N_29934);
nor UO_1822 (O_1822,N_29861,N_29889);
and UO_1823 (O_1823,N_29986,N_29894);
or UO_1824 (O_1824,N_29856,N_29896);
or UO_1825 (O_1825,N_29884,N_29928);
and UO_1826 (O_1826,N_29810,N_29997);
or UO_1827 (O_1827,N_29812,N_29850);
nand UO_1828 (O_1828,N_29835,N_29926);
xnor UO_1829 (O_1829,N_29881,N_29839);
xnor UO_1830 (O_1830,N_29837,N_29960);
nor UO_1831 (O_1831,N_29827,N_29930);
xor UO_1832 (O_1832,N_29831,N_29971);
xor UO_1833 (O_1833,N_29984,N_29865);
or UO_1834 (O_1834,N_29904,N_29852);
or UO_1835 (O_1835,N_29812,N_29843);
or UO_1836 (O_1836,N_29859,N_29994);
and UO_1837 (O_1837,N_29836,N_29902);
and UO_1838 (O_1838,N_29901,N_29865);
and UO_1839 (O_1839,N_29992,N_29913);
nand UO_1840 (O_1840,N_29897,N_29937);
nand UO_1841 (O_1841,N_29941,N_29902);
and UO_1842 (O_1842,N_29988,N_29921);
nor UO_1843 (O_1843,N_29881,N_29951);
nor UO_1844 (O_1844,N_29837,N_29903);
xor UO_1845 (O_1845,N_29901,N_29997);
nand UO_1846 (O_1846,N_29825,N_29821);
and UO_1847 (O_1847,N_29824,N_29878);
xor UO_1848 (O_1848,N_29835,N_29987);
nand UO_1849 (O_1849,N_29906,N_29987);
nand UO_1850 (O_1850,N_29867,N_29834);
and UO_1851 (O_1851,N_29861,N_29884);
and UO_1852 (O_1852,N_29939,N_29937);
nand UO_1853 (O_1853,N_29955,N_29817);
and UO_1854 (O_1854,N_29845,N_29834);
nor UO_1855 (O_1855,N_29873,N_29880);
xor UO_1856 (O_1856,N_29939,N_29874);
and UO_1857 (O_1857,N_29909,N_29920);
or UO_1858 (O_1858,N_29853,N_29975);
xor UO_1859 (O_1859,N_29896,N_29805);
and UO_1860 (O_1860,N_29817,N_29973);
xnor UO_1861 (O_1861,N_29892,N_29819);
and UO_1862 (O_1862,N_29919,N_29874);
nand UO_1863 (O_1863,N_29899,N_29887);
or UO_1864 (O_1864,N_29944,N_29852);
or UO_1865 (O_1865,N_29971,N_29925);
or UO_1866 (O_1866,N_29864,N_29877);
or UO_1867 (O_1867,N_29886,N_29960);
nor UO_1868 (O_1868,N_29916,N_29882);
and UO_1869 (O_1869,N_29932,N_29885);
nand UO_1870 (O_1870,N_29848,N_29996);
and UO_1871 (O_1871,N_29916,N_29854);
or UO_1872 (O_1872,N_29878,N_29866);
or UO_1873 (O_1873,N_29806,N_29902);
and UO_1874 (O_1874,N_29870,N_29858);
xor UO_1875 (O_1875,N_29817,N_29845);
and UO_1876 (O_1876,N_29806,N_29896);
xor UO_1877 (O_1877,N_29901,N_29999);
nor UO_1878 (O_1878,N_29994,N_29869);
or UO_1879 (O_1879,N_29827,N_29905);
or UO_1880 (O_1880,N_29956,N_29919);
xor UO_1881 (O_1881,N_29958,N_29928);
xor UO_1882 (O_1882,N_29995,N_29999);
nor UO_1883 (O_1883,N_29948,N_29975);
nand UO_1884 (O_1884,N_29994,N_29804);
or UO_1885 (O_1885,N_29858,N_29974);
nand UO_1886 (O_1886,N_29833,N_29882);
nor UO_1887 (O_1887,N_29888,N_29855);
or UO_1888 (O_1888,N_29874,N_29838);
or UO_1889 (O_1889,N_29986,N_29973);
nand UO_1890 (O_1890,N_29926,N_29999);
xnor UO_1891 (O_1891,N_29850,N_29841);
xor UO_1892 (O_1892,N_29944,N_29889);
and UO_1893 (O_1893,N_29828,N_29893);
nand UO_1894 (O_1894,N_29960,N_29889);
and UO_1895 (O_1895,N_29874,N_29806);
or UO_1896 (O_1896,N_29880,N_29870);
xnor UO_1897 (O_1897,N_29969,N_29894);
nand UO_1898 (O_1898,N_29990,N_29985);
or UO_1899 (O_1899,N_29983,N_29804);
or UO_1900 (O_1900,N_29877,N_29874);
nand UO_1901 (O_1901,N_29946,N_29884);
nor UO_1902 (O_1902,N_29890,N_29925);
nand UO_1903 (O_1903,N_29956,N_29995);
nor UO_1904 (O_1904,N_29826,N_29805);
nand UO_1905 (O_1905,N_29926,N_29945);
nor UO_1906 (O_1906,N_29986,N_29970);
and UO_1907 (O_1907,N_29935,N_29915);
nor UO_1908 (O_1908,N_29839,N_29942);
xnor UO_1909 (O_1909,N_29989,N_29863);
and UO_1910 (O_1910,N_29869,N_29881);
xnor UO_1911 (O_1911,N_29949,N_29975);
nand UO_1912 (O_1912,N_29879,N_29851);
xor UO_1913 (O_1913,N_29830,N_29877);
xnor UO_1914 (O_1914,N_29818,N_29927);
and UO_1915 (O_1915,N_29845,N_29806);
nor UO_1916 (O_1916,N_29828,N_29938);
or UO_1917 (O_1917,N_29866,N_29928);
nand UO_1918 (O_1918,N_29817,N_29949);
or UO_1919 (O_1919,N_29838,N_29982);
xnor UO_1920 (O_1920,N_29825,N_29800);
and UO_1921 (O_1921,N_29979,N_29811);
nor UO_1922 (O_1922,N_29850,N_29996);
xor UO_1923 (O_1923,N_29822,N_29977);
and UO_1924 (O_1924,N_29844,N_29981);
nor UO_1925 (O_1925,N_29842,N_29817);
nor UO_1926 (O_1926,N_29974,N_29882);
and UO_1927 (O_1927,N_29955,N_29979);
or UO_1928 (O_1928,N_29944,N_29959);
or UO_1929 (O_1929,N_29964,N_29812);
xnor UO_1930 (O_1930,N_29882,N_29932);
and UO_1931 (O_1931,N_29860,N_29943);
or UO_1932 (O_1932,N_29979,N_29853);
or UO_1933 (O_1933,N_29983,N_29995);
and UO_1934 (O_1934,N_29896,N_29817);
or UO_1935 (O_1935,N_29906,N_29883);
nand UO_1936 (O_1936,N_29968,N_29888);
and UO_1937 (O_1937,N_29872,N_29845);
or UO_1938 (O_1938,N_29892,N_29834);
nor UO_1939 (O_1939,N_29934,N_29967);
nor UO_1940 (O_1940,N_29961,N_29835);
nand UO_1941 (O_1941,N_29990,N_29929);
xnor UO_1942 (O_1942,N_29811,N_29980);
nand UO_1943 (O_1943,N_29827,N_29851);
and UO_1944 (O_1944,N_29937,N_29936);
and UO_1945 (O_1945,N_29853,N_29939);
xnor UO_1946 (O_1946,N_29870,N_29964);
and UO_1947 (O_1947,N_29969,N_29966);
nand UO_1948 (O_1948,N_29899,N_29936);
nor UO_1949 (O_1949,N_29846,N_29818);
nor UO_1950 (O_1950,N_29995,N_29912);
nand UO_1951 (O_1951,N_29891,N_29949);
xnor UO_1952 (O_1952,N_29991,N_29962);
nand UO_1953 (O_1953,N_29985,N_29837);
or UO_1954 (O_1954,N_29945,N_29805);
and UO_1955 (O_1955,N_29977,N_29802);
and UO_1956 (O_1956,N_29877,N_29868);
and UO_1957 (O_1957,N_29978,N_29917);
or UO_1958 (O_1958,N_29808,N_29948);
and UO_1959 (O_1959,N_29922,N_29890);
nand UO_1960 (O_1960,N_29851,N_29997);
nor UO_1961 (O_1961,N_29815,N_29968);
nand UO_1962 (O_1962,N_29972,N_29877);
nor UO_1963 (O_1963,N_29990,N_29891);
or UO_1964 (O_1964,N_29845,N_29850);
or UO_1965 (O_1965,N_29923,N_29939);
or UO_1966 (O_1966,N_29913,N_29960);
nor UO_1967 (O_1967,N_29942,N_29980);
nand UO_1968 (O_1968,N_29990,N_29976);
or UO_1969 (O_1969,N_29805,N_29927);
or UO_1970 (O_1970,N_29977,N_29804);
xor UO_1971 (O_1971,N_29939,N_29808);
xor UO_1972 (O_1972,N_29981,N_29935);
and UO_1973 (O_1973,N_29966,N_29801);
nand UO_1974 (O_1974,N_29855,N_29900);
or UO_1975 (O_1975,N_29993,N_29893);
nand UO_1976 (O_1976,N_29810,N_29934);
or UO_1977 (O_1977,N_29948,N_29901);
xnor UO_1978 (O_1978,N_29887,N_29814);
nor UO_1979 (O_1979,N_29891,N_29868);
nor UO_1980 (O_1980,N_29992,N_29805);
nand UO_1981 (O_1981,N_29996,N_29840);
xnor UO_1982 (O_1982,N_29955,N_29904);
nor UO_1983 (O_1983,N_29988,N_29849);
nor UO_1984 (O_1984,N_29931,N_29889);
nor UO_1985 (O_1985,N_29955,N_29837);
and UO_1986 (O_1986,N_29999,N_29863);
or UO_1987 (O_1987,N_29877,N_29876);
and UO_1988 (O_1988,N_29922,N_29999);
and UO_1989 (O_1989,N_29933,N_29885);
and UO_1990 (O_1990,N_29973,N_29967);
nand UO_1991 (O_1991,N_29984,N_29917);
or UO_1992 (O_1992,N_29944,N_29843);
xnor UO_1993 (O_1993,N_29922,N_29953);
and UO_1994 (O_1994,N_29856,N_29827);
or UO_1995 (O_1995,N_29904,N_29936);
or UO_1996 (O_1996,N_29925,N_29868);
or UO_1997 (O_1997,N_29891,N_29941);
and UO_1998 (O_1998,N_29874,N_29894);
xor UO_1999 (O_1999,N_29972,N_29973);
xnor UO_2000 (O_2000,N_29964,N_29931);
nor UO_2001 (O_2001,N_29827,N_29923);
or UO_2002 (O_2002,N_29943,N_29892);
or UO_2003 (O_2003,N_29876,N_29898);
or UO_2004 (O_2004,N_29803,N_29943);
and UO_2005 (O_2005,N_29883,N_29960);
nand UO_2006 (O_2006,N_29937,N_29986);
or UO_2007 (O_2007,N_29858,N_29958);
and UO_2008 (O_2008,N_29967,N_29843);
nor UO_2009 (O_2009,N_29998,N_29995);
and UO_2010 (O_2010,N_29929,N_29967);
xnor UO_2011 (O_2011,N_29993,N_29867);
or UO_2012 (O_2012,N_29837,N_29882);
xnor UO_2013 (O_2013,N_29960,N_29976);
and UO_2014 (O_2014,N_29913,N_29882);
xnor UO_2015 (O_2015,N_29893,N_29908);
and UO_2016 (O_2016,N_29897,N_29992);
and UO_2017 (O_2017,N_29957,N_29923);
and UO_2018 (O_2018,N_29882,N_29889);
xnor UO_2019 (O_2019,N_29825,N_29941);
nand UO_2020 (O_2020,N_29955,N_29986);
xnor UO_2021 (O_2021,N_29849,N_29911);
and UO_2022 (O_2022,N_29988,N_29934);
xnor UO_2023 (O_2023,N_29967,N_29931);
nand UO_2024 (O_2024,N_29812,N_29899);
and UO_2025 (O_2025,N_29820,N_29827);
and UO_2026 (O_2026,N_29958,N_29902);
nand UO_2027 (O_2027,N_29914,N_29815);
nor UO_2028 (O_2028,N_29843,N_29988);
or UO_2029 (O_2029,N_29995,N_29990);
and UO_2030 (O_2030,N_29918,N_29990);
nor UO_2031 (O_2031,N_29870,N_29965);
xor UO_2032 (O_2032,N_29986,N_29911);
and UO_2033 (O_2033,N_29822,N_29873);
and UO_2034 (O_2034,N_29905,N_29955);
nor UO_2035 (O_2035,N_29811,N_29965);
xor UO_2036 (O_2036,N_29823,N_29949);
nor UO_2037 (O_2037,N_29901,N_29835);
xor UO_2038 (O_2038,N_29992,N_29930);
xor UO_2039 (O_2039,N_29828,N_29882);
xnor UO_2040 (O_2040,N_29960,N_29875);
and UO_2041 (O_2041,N_29881,N_29809);
xor UO_2042 (O_2042,N_29924,N_29969);
xor UO_2043 (O_2043,N_29824,N_29889);
or UO_2044 (O_2044,N_29966,N_29955);
nor UO_2045 (O_2045,N_29887,N_29843);
or UO_2046 (O_2046,N_29973,N_29929);
nor UO_2047 (O_2047,N_29853,N_29836);
xor UO_2048 (O_2048,N_29958,N_29930);
nand UO_2049 (O_2049,N_29832,N_29807);
xor UO_2050 (O_2050,N_29998,N_29878);
or UO_2051 (O_2051,N_29977,N_29867);
nand UO_2052 (O_2052,N_29996,N_29869);
and UO_2053 (O_2053,N_29873,N_29955);
and UO_2054 (O_2054,N_29927,N_29994);
xor UO_2055 (O_2055,N_29842,N_29827);
xnor UO_2056 (O_2056,N_29971,N_29834);
and UO_2057 (O_2057,N_29976,N_29877);
or UO_2058 (O_2058,N_29883,N_29817);
or UO_2059 (O_2059,N_29836,N_29891);
nand UO_2060 (O_2060,N_29922,N_29894);
nand UO_2061 (O_2061,N_29803,N_29949);
nor UO_2062 (O_2062,N_29951,N_29993);
nor UO_2063 (O_2063,N_29845,N_29875);
or UO_2064 (O_2064,N_29972,N_29949);
or UO_2065 (O_2065,N_29959,N_29806);
nor UO_2066 (O_2066,N_29933,N_29857);
nor UO_2067 (O_2067,N_29903,N_29803);
nor UO_2068 (O_2068,N_29941,N_29863);
and UO_2069 (O_2069,N_29972,N_29902);
nor UO_2070 (O_2070,N_29836,N_29817);
xnor UO_2071 (O_2071,N_29842,N_29980);
and UO_2072 (O_2072,N_29858,N_29972);
and UO_2073 (O_2073,N_29869,N_29973);
nand UO_2074 (O_2074,N_29928,N_29943);
nor UO_2075 (O_2075,N_29810,N_29858);
and UO_2076 (O_2076,N_29849,N_29990);
nand UO_2077 (O_2077,N_29922,N_29979);
nor UO_2078 (O_2078,N_29877,N_29949);
nor UO_2079 (O_2079,N_29862,N_29875);
nand UO_2080 (O_2080,N_29867,N_29981);
or UO_2081 (O_2081,N_29839,N_29898);
and UO_2082 (O_2082,N_29873,N_29872);
nand UO_2083 (O_2083,N_29999,N_29895);
xnor UO_2084 (O_2084,N_29869,N_29891);
and UO_2085 (O_2085,N_29968,N_29836);
or UO_2086 (O_2086,N_29969,N_29907);
xnor UO_2087 (O_2087,N_29980,N_29999);
nor UO_2088 (O_2088,N_29856,N_29965);
or UO_2089 (O_2089,N_29908,N_29832);
and UO_2090 (O_2090,N_29807,N_29836);
nor UO_2091 (O_2091,N_29834,N_29878);
or UO_2092 (O_2092,N_29914,N_29992);
nand UO_2093 (O_2093,N_29990,N_29981);
xor UO_2094 (O_2094,N_29966,N_29904);
or UO_2095 (O_2095,N_29939,N_29885);
and UO_2096 (O_2096,N_29829,N_29884);
or UO_2097 (O_2097,N_29935,N_29966);
xor UO_2098 (O_2098,N_29957,N_29804);
xnor UO_2099 (O_2099,N_29840,N_29889);
nor UO_2100 (O_2100,N_29969,N_29800);
xor UO_2101 (O_2101,N_29812,N_29970);
xnor UO_2102 (O_2102,N_29965,N_29944);
nand UO_2103 (O_2103,N_29919,N_29837);
nand UO_2104 (O_2104,N_29838,N_29897);
nor UO_2105 (O_2105,N_29811,N_29833);
xnor UO_2106 (O_2106,N_29998,N_29978);
nand UO_2107 (O_2107,N_29944,N_29969);
and UO_2108 (O_2108,N_29989,N_29897);
and UO_2109 (O_2109,N_29897,N_29964);
or UO_2110 (O_2110,N_29946,N_29822);
nand UO_2111 (O_2111,N_29910,N_29846);
xor UO_2112 (O_2112,N_29965,N_29925);
and UO_2113 (O_2113,N_29928,N_29924);
xnor UO_2114 (O_2114,N_29800,N_29810);
nand UO_2115 (O_2115,N_29829,N_29922);
xor UO_2116 (O_2116,N_29992,N_29986);
and UO_2117 (O_2117,N_29914,N_29890);
nor UO_2118 (O_2118,N_29827,N_29836);
xor UO_2119 (O_2119,N_29816,N_29859);
nand UO_2120 (O_2120,N_29892,N_29813);
nand UO_2121 (O_2121,N_29981,N_29912);
and UO_2122 (O_2122,N_29996,N_29870);
and UO_2123 (O_2123,N_29858,N_29976);
xnor UO_2124 (O_2124,N_29958,N_29886);
nand UO_2125 (O_2125,N_29994,N_29885);
nand UO_2126 (O_2126,N_29890,N_29847);
nand UO_2127 (O_2127,N_29907,N_29919);
nand UO_2128 (O_2128,N_29962,N_29993);
nor UO_2129 (O_2129,N_29845,N_29802);
xor UO_2130 (O_2130,N_29956,N_29957);
nand UO_2131 (O_2131,N_29898,N_29902);
and UO_2132 (O_2132,N_29811,N_29946);
nand UO_2133 (O_2133,N_29809,N_29944);
or UO_2134 (O_2134,N_29969,N_29815);
and UO_2135 (O_2135,N_29890,N_29868);
xor UO_2136 (O_2136,N_29805,N_29871);
or UO_2137 (O_2137,N_29922,N_29856);
nand UO_2138 (O_2138,N_29999,N_29828);
or UO_2139 (O_2139,N_29961,N_29848);
nand UO_2140 (O_2140,N_29988,N_29853);
xor UO_2141 (O_2141,N_29988,N_29952);
nor UO_2142 (O_2142,N_29811,N_29858);
or UO_2143 (O_2143,N_29861,N_29967);
or UO_2144 (O_2144,N_29860,N_29868);
nand UO_2145 (O_2145,N_29931,N_29902);
xor UO_2146 (O_2146,N_29896,N_29844);
or UO_2147 (O_2147,N_29944,N_29987);
and UO_2148 (O_2148,N_29900,N_29977);
xnor UO_2149 (O_2149,N_29870,N_29883);
xnor UO_2150 (O_2150,N_29971,N_29810);
xnor UO_2151 (O_2151,N_29878,N_29825);
xor UO_2152 (O_2152,N_29813,N_29954);
xor UO_2153 (O_2153,N_29805,N_29898);
nor UO_2154 (O_2154,N_29889,N_29904);
nor UO_2155 (O_2155,N_29943,N_29946);
or UO_2156 (O_2156,N_29838,N_29998);
or UO_2157 (O_2157,N_29824,N_29869);
or UO_2158 (O_2158,N_29951,N_29827);
nand UO_2159 (O_2159,N_29844,N_29847);
xor UO_2160 (O_2160,N_29918,N_29839);
and UO_2161 (O_2161,N_29810,N_29885);
and UO_2162 (O_2162,N_29958,N_29856);
or UO_2163 (O_2163,N_29823,N_29987);
nand UO_2164 (O_2164,N_29823,N_29913);
nor UO_2165 (O_2165,N_29982,N_29894);
or UO_2166 (O_2166,N_29888,N_29817);
or UO_2167 (O_2167,N_29971,N_29981);
nor UO_2168 (O_2168,N_29895,N_29937);
or UO_2169 (O_2169,N_29974,N_29993);
or UO_2170 (O_2170,N_29848,N_29887);
xnor UO_2171 (O_2171,N_29918,N_29939);
nand UO_2172 (O_2172,N_29873,N_29897);
xnor UO_2173 (O_2173,N_29929,N_29888);
and UO_2174 (O_2174,N_29979,N_29877);
nor UO_2175 (O_2175,N_29965,N_29802);
and UO_2176 (O_2176,N_29970,N_29943);
and UO_2177 (O_2177,N_29819,N_29950);
xnor UO_2178 (O_2178,N_29870,N_29909);
nand UO_2179 (O_2179,N_29993,N_29938);
and UO_2180 (O_2180,N_29850,N_29872);
xor UO_2181 (O_2181,N_29837,N_29998);
nand UO_2182 (O_2182,N_29817,N_29965);
or UO_2183 (O_2183,N_29981,N_29959);
nand UO_2184 (O_2184,N_29993,N_29891);
and UO_2185 (O_2185,N_29909,N_29916);
nand UO_2186 (O_2186,N_29951,N_29901);
and UO_2187 (O_2187,N_29883,N_29963);
or UO_2188 (O_2188,N_29900,N_29867);
and UO_2189 (O_2189,N_29967,N_29887);
nor UO_2190 (O_2190,N_29884,N_29866);
nor UO_2191 (O_2191,N_29841,N_29900);
xnor UO_2192 (O_2192,N_29890,N_29978);
and UO_2193 (O_2193,N_29915,N_29817);
xnor UO_2194 (O_2194,N_29980,N_29931);
nor UO_2195 (O_2195,N_29924,N_29862);
xor UO_2196 (O_2196,N_29866,N_29909);
nor UO_2197 (O_2197,N_29861,N_29817);
nor UO_2198 (O_2198,N_29881,N_29878);
xor UO_2199 (O_2199,N_29927,N_29840);
nand UO_2200 (O_2200,N_29973,N_29863);
or UO_2201 (O_2201,N_29836,N_29869);
nor UO_2202 (O_2202,N_29934,N_29932);
nor UO_2203 (O_2203,N_29891,N_29813);
nor UO_2204 (O_2204,N_29918,N_29891);
nand UO_2205 (O_2205,N_29956,N_29912);
or UO_2206 (O_2206,N_29889,N_29807);
and UO_2207 (O_2207,N_29851,N_29953);
or UO_2208 (O_2208,N_29828,N_29850);
or UO_2209 (O_2209,N_29882,N_29911);
xor UO_2210 (O_2210,N_29887,N_29959);
nand UO_2211 (O_2211,N_29994,N_29807);
nand UO_2212 (O_2212,N_29940,N_29821);
nand UO_2213 (O_2213,N_29943,N_29924);
xor UO_2214 (O_2214,N_29945,N_29821);
xnor UO_2215 (O_2215,N_29958,N_29832);
nor UO_2216 (O_2216,N_29952,N_29956);
or UO_2217 (O_2217,N_29966,N_29906);
nand UO_2218 (O_2218,N_29804,N_29961);
or UO_2219 (O_2219,N_29915,N_29948);
and UO_2220 (O_2220,N_29892,N_29963);
or UO_2221 (O_2221,N_29861,N_29860);
xor UO_2222 (O_2222,N_29845,N_29827);
nand UO_2223 (O_2223,N_29813,N_29882);
xnor UO_2224 (O_2224,N_29847,N_29921);
nor UO_2225 (O_2225,N_29936,N_29844);
nor UO_2226 (O_2226,N_29929,N_29847);
or UO_2227 (O_2227,N_29966,N_29859);
nor UO_2228 (O_2228,N_29892,N_29812);
xor UO_2229 (O_2229,N_29804,N_29904);
or UO_2230 (O_2230,N_29867,N_29904);
nand UO_2231 (O_2231,N_29889,N_29809);
or UO_2232 (O_2232,N_29855,N_29996);
or UO_2233 (O_2233,N_29934,N_29816);
xor UO_2234 (O_2234,N_29837,N_29802);
or UO_2235 (O_2235,N_29896,N_29955);
and UO_2236 (O_2236,N_29854,N_29880);
and UO_2237 (O_2237,N_29971,N_29983);
and UO_2238 (O_2238,N_29993,N_29991);
or UO_2239 (O_2239,N_29911,N_29931);
nand UO_2240 (O_2240,N_29961,N_29805);
or UO_2241 (O_2241,N_29863,N_29814);
xnor UO_2242 (O_2242,N_29916,N_29867);
nor UO_2243 (O_2243,N_29932,N_29918);
xor UO_2244 (O_2244,N_29855,N_29999);
nor UO_2245 (O_2245,N_29921,N_29963);
or UO_2246 (O_2246,N_29951,N_29894);
nand UO_2247 (O_2247,N_29863,N_29842);
nand UO_2248 (O_2248,N_29931,N_29852);
xor UO_2249 (O_2249,N_29894,N_29829);
xor UO_2250 (O_2250,N_29860,N_29887);
nand UO_2251 (O_2251,N_29963,N_29871);
nand UO_2252 (O_2252,N_29922,N_29917);
nor UO_2253 (O_2253,N_29984,N_29875);
and UO_2254 (O_2254,N_29880,N_29914);
nand UO_2255 (O_2255,N_29957,N_29815);
nand UO_2256 (O_2256,N_29905,N_29979);
and UO_2257 (O_2257,N_29881,N_29816);
xnor UO_2258 (O_2258,N_29958,N_29879);
nor UO_2259 (O_2259,N_29874,N_29825);
nand UO_2260 (O_2260,N_29892,N_29852);
xnor UO_2261 (O_2261,N_29936,N_29952);
nor UO_2262 (O_2262,N_29974,N_29903);
xnor UO_2263 (O_2263,N_29850,N_29846);
or UO_2264 (O_2264,N_29949,N_29998);
or UO_2265 (O_2265,N_29800,N_29832);
nor UO_2266 (O_2266,N_29881,N_29982);
or UO_2267 (O_2267,N_29944,N_29836);
or UO_2268 (O_2268,N_29813,N_29938);
nand UO_2269 (O_2269,N_29982,N_29991);
or UO_2270 (O_2270,N_29898,N_29952);
nor UO_2271 (O_2271,N_29958,N_29844);
xor UO_2272 (O_2272,N_29929,N_29880);
nor UO_2273 (O_2273,N_29957,N_29936);
nand UO_2274 (O_2274,N_29901,N_29839);
nand UO_2275 (O_2275,N_29815,N_29983);
xor UO_2276 (O_2276,N_29826,N_29835);
nand UO_2277 (O_2277,N_29822,N_29844);
or UO_2278 (O_2278,N_29811,N_29836);
and UO_2279 (O_2279,N_29833,N_29962);
nor UO_2280 (O_2280,N_29988,N_29989);
and UO_2281 (O_2281,N_29936,N_29876);
nor UO_2282 (O_2282,N_29899,N_29825);
xor UO_2283 (O_2283,N_29857,N_29915);
and UO_2284 (O_2284,N_29978,N_29904);
or UO_2285 (O_2285,N_29815,N_29980);
or UO_2286 (O_2286,N_29938,N_29995);
and UO_2287 (O_2287,N_29930,N_29807);
nor UO_2288 (O_2288,N_29819,N_29914);
nand UO_2289 (O_2289,N_29807,N_29938);
nor UO_2290 (O_2290,N_29979,N_29802);
nor UO_2291 (O_2291,N_29976,N_29928);
xnor UO_2292 (O_2292,N_29947,N_29978);
and UO_2293 (O_2293,N_29950,N_29874);
nand UO_2294 (O_2294,N_29929,N_29947);
or UO_2295 (O_2295,N_29808,N_29937);
nor UO_2296 (O_2296,N_29894,N_29913);
nand UO_2297 (O_2297,N_29892,N_29853);
and UO_2298 (O_2298,N_29806,N_29857);
xnor UO_2299 (O_2299,N_29959,N_29811);
nor UO_2300 (O_2300,N_29941,N_29885);
nand UO_2301 (O_2301,N_29998,N_29993);
nor UO_2302 (O_2302,N_29814,N_29813);
and UO_2303 (O_2303,N_29899,N_29949);
nor UO_2304 (O_2304,N_29820,N_29841);
nor UO_2305 (O_2305,N_29875,N_29901);
and UO_2306 (O_2306,N_29811,N_29999);
nand UO_2307 (O_2307,N_29921,N_29858);
nor UO_2308 (O_2308,N_29962,N_29986);
and UO_2309 (O_2309,N_29939,N_29909);
xnor UO_2310 (O_2310,N_29802,N_29866);
and UO_2311 (O_2311,N_29866,N_29883);
nand UO_2312 (O_2312,N_29856,N_29828);
and UO_2313 (O_2313,N_29863,N_29843);
or UO_2314 (O_2314,N_29899,N_29813);
xor UO_2315 (O_2315,N_29922,N_29804);
nand UO_2316 (O_2316,N_29873,N_29933);
nand UO_2317 (O_2317,N_29876,N_29862);
and UO_2318 (O_2318,N_29824,N_29963);
xnor UO_2319 (O_2319,N_29914,N_29982);
and UO_2320 (O_2320,N_29891,N_29976);
nand UO_2321 (O_2321,N_29832,N_29849);
and UO_2322 (O_2322,N_29923,N_29914);
or UO_2323 (O_2323,N_29967,N_29885);
and UO_2324 (O_2324,N_29983,N_29992);
nand UO_2325 (O_2325,N_29946,N_29968);
xnor UO_2326 (O_2326,N_29873,N_29838);
nand UO_2327 (O_2327,N_29859,N_29963);
xnor UO_2328 (O_2328,N_29869,N_29935);
and UO_2329 (O_2329,N_29858,N_29815);
xor UO_2330 (O_2330,N_29896,N_29802);
nand UO_2331 (O_2331,N_29904,N_29960);
nor UO_2332 (O_2332,N_29828,N_29809);
and UO_2333 (O_2333,N_29910,N_29905);
xnor UO_2334 (O_2334,N_29818,N_29983);
xnor UO_2335 (O_2335,N_29998,N_29897);
nand UO_2336 (O_2336,N_29818,N_29815);
or UO_2337 (O_2337,N_29862,N_29971);
nand UO_2338 (O_2338,N_29839,N_29924);
nand UO_2339 (O_2339,N_29997,N_29886);
xnor UO_2340 (O_2340,N_29830,N_29958);
xnor UO_2341 (O_2341,N_29880,N_29802);
and UO_2342 (O_2342,N_29979,N_29993);
nand UO_2343 (O_2343,N_29915,N_29813);
or UO_2344 (O_2344,N_29985,N_29867);
and UO_2345 (O_2345,N_29885,N_29808);
xor UO_2346 (O_2346,N_29883,N_29948);
or UO_2347 (O_2347,N_29864,N_29801);
and UO_2348 (O_2348,N_29895,N_29965);
nor UO_2349 (O_2349,N_29898,N_29851);
xnor UO_2350 (O_2350,N_29863,N_29887);
xor UO_2351 (O_2351,N_29846,N_29865);
or UO_2352 (O_2352,N_29958,N_29909);
or UO_2353 (O_2353,N_29980,N_29964);
and UO_2354 (O_2354,N_29842,N_29853);
nor UO_2355 (O_2355,N_29820,N_29992);
and UO_2356 (O_2356,N_29935,N_29990);
nor UO_2357 (O_2357,N_29864,N_29817);
xnor UO_2358 (O_2358,N_29859,N_29933);
nor UO_2359 (O_2359,N_29806,N_29866);
nor UO_2360 (O_2360,N_29819,N_29984);
xor UO_2361 (O_2361,N_29866,N_29825);
nand UO_2362 (O_2362,N_29923,N_29839);
and UO_2363 (O_2363,N_29862,N_29828);
or UO_2364 (O_2364,N_29843,N_29818);
nor UO_2365 (O_2365,N_29895,N_29845);
nand UO_2366 (O_2366,N_29998,N_29946);
or UO_2367 (O_2367,N_29977,N_29850);
nor UO_2368 (O_2368,N_29854,N_29968);
xor UO_2369 (O_2369,N_29962,N_29932);
or UO_2370 (O_2370,N_29892,N_29863);
and UO_2371 (O_2371,N_29935,N_29832);
nor UO_2372 (O_2372,N_29850,N_29985);
nand UO_2373 (O_2373,N_29833,N_29959);
or UO_2374 (O_2374,N_29929,N_29930);
or UO_2375 (O_2375,N_29949,N_29818);
xor UO_2376 (O_2376,N_29965,N_29953);
xor UO_2377 (O_2377,N_29859,N_29840);
and UO_2378 (O_2378,N_29879,N_29956);
or UO_2379 (O_2379,N_29816,N_29889);
or UO_2380 (O_2380,N_29885,N_29908);
or UO_2381 (O_2381,N_29991,N_29927);
nor UO_2382 (O_2382,N_29945,N_29889);
nor UO_2383 (O_2383,N_29918,N_29905);
nor UO_2384 (O_2384,N_29879,N_29923);
and UO_2385 (O_2385,N_29878,N_29809);
and UO_2386 (O_2386,N_29943,N_29955);
nor UO_2387 (O_2387,N_29828,N_29847);
nor UO_2388 (O_2388,N_29951,N_29813);
nand UO_2389 (O_2389,N_29894,N_29826);
nor UO_2390 (O_2390,N_29836,N_29979);
or UO_2391 (O_2391,N_29803,N_29969);
xor UO_2392 (O_2392,N_29884,N_29899);
nand UO_2393 (O_2393,N_29993,N_29860);
nor UO_2394 (O_2394,N_29843,N_29819);
or UO_2395 (O_2395,N_29960,N_29989);
xnor UO_2396 (O_2396,N_29929,N_29807);
xor UO_2397 (O_2397,N_29868,N_29879);
xor UO_2398 (O_2398,N_29977,N_29922);
nand UO_2399 (O_2399,N_29831,N_29974);
xor UO_2400 (O_2400,N_29979,N_29934);
nor UO_2401 (O_2401,N_29863,N_29827);
nor UO_2402 (O_2402,N_29937,N_29924);
nor UO_2403 (O_2403,N_29870,N_29833);
or UO_2404 (O_2404,N_29926,N_29942);
and UO_2405 (O_2405,N_29801,N_29992);
and UO_2406 (O_2406,N_29866,N_29993);
or UO_2407 (O_2407,N_29961,N_29953);
nor UO_2408 (O_2408,N_29883,N_29966);
or UO_2409 (O_2409,N_29862,N_29965);
and UO_2410 (O_2410,N_29906,N_29930);
nand UO_2411 (O_2411,N_29896,N_29807);
nand UO_2412 (O_2412,N_29852,N_29864);
and UO_2413 (O_2413,N_29938,N_29911);
or UO_2414 (O_2414,N_29968,N_29919);
nor UO_2415 (O_2415,N_29853,N_29984);
nand UO_2416 (O_2416,N_29998,N_29922);
xnor UO_2417 (O_2417,N_29941,N_29843);
nor UO_2418 (O_2418,N_29895,N_29927);
xor UO_2419 (O_2419,N_29834,N_29916);
or UO_2420 (O_2420,N_29915,N_29835);
xor UO_2421 (O_2421,N_29809,N_29837);
and UO_2422 (O_2422,N_29936,N_29996);
and UO_2423 (O_2423,N_29887,N_29968);
and UO_2424 (O_2424,N_29885,N_29811);
nor UO_2425 (O_2425,N_29929,N_29877);
nand UO_2426 (O_2426,N_29936,N_29980);
nand UO_2427 (O_2427,N_29898,N_29969);
nor UO_2428 (O_2428,N_29954,N_29841);
xnor UO_2429 (O_2429,N_29950,N_29914);
and UO_2430 (O_2430,N_29995,N_29835);
nand UO_2431 (O_2431,N_29954,N_29994);
nor UO_2432 (O_2432,N_29813,N_29976);
or UO_2433 (O_2433,N_29841,N_29947);
nand UO_2434 (O_2434,N_29893,N_29939);
nor UO_2435 (O_2435,N_29938,N_29892);
or UO_2436 (O_2436,N_29916,N_29864);
and UO_2437 (O_2437,N_29855,N_29847);
nor UO_2438 (O_2438,N_29883,N_29905);
nand UO_2439 (O_2439,N_29910,N_29966);
and UO_2440 (O_2440,N_29988,N_29923);
xor UO_2441 (O_2441,N_29931,N_29803);
nand UO_2442 (O_2442,N_29972,N_29812);
nor UO_2443 (O_2443,N_29932,N_29851);
or UO_2444 (O_2444,N_29937,N_29820);
nand UO_2445 (O_2445,N_29932,N_29839);
or UO_2446 (O_2446,N_29934,N_29922);
and UO_2447 (O_2447,N_29961,N_29924);
or UO_2448 (O_2448,N_29877,N_29962);
nand UO_2449 (O_2449,N_29891,N_29939);
xor UO_2450 (O_2450,N_29800,N_29928);
xor UO_2451 (O_2451,N_29989,N_29865);
and UO_2452 (O_2452,N_29926,N_29803);
xor UO_2453 (O_2453,N_29944,N_29951);
and UO_2454 (O_2454,N_29859,N_29943);
xor UO_2455 (O_2455,N_29918,N_29832);
and UO_2456 (O_2456,N_29868,N_29892);
and UO_2457 (O_2457,N_29985,N_29911);
nor UO_2458 (O_2458,N_29992,N_29898);
nor UO_2459 (O_2459,N_29921,N_29948);
and UO_2460 (O_2460,N_29993,N_29834);
xnor UO_2461 (O_2461,N_29928,N_29960);
or UO_2462 (O_2462,N_29966,N_29860);
xnor UO_2463 (O_2463,N_29966,N_29980);
and UO_2464 (O_2464,N_29852,N_29916);
nand UO_2465 (O_2465,N_29952,N_29842);
nor UO_2466 (O_2466,N_29845,N_29825);
nor UO_2467 (O_2467,N_29992,N_29819);
nand UO_2468 (O_2468,N_29998,N_29914);
nor UO_2469 (O_2469,N_29833,N_29886);
or UO_2470 (O_2470,N_29914,N_29920);
xor UO_2471 (O_2471,N_29881,N_29940);
nor UO_2472 (O_2472,N_29886,N_29839);
or UO_2473 (O_2473,N_29975,N_29875);
and UO_2474 (O_2474,N_29977,N_29965);
or UO_2475 (O_2475,N_29949,N_29978);
xnor UO_2476 (O_2476,N_29899,N_29937);
nand UO_2477 (O_2477,N_29951,N_29885);
nor UO_2478 (O_2478,N_29972,N_29990);
nor UO_2479 (O_2479,N_29802,N_29873);
nand UO_2480 (O_2480,N_29869,N_29834);
xnor UO_2481 (O_2481,N_29801,N_29906);
nand UO_2482 (O_2482,N_29806,N_29949);
or UO_2483 (O_2483,N_29939,N_29922);
xnor UO_2484 (O_2484,N_29964,N_29827);
nand UO_2485 (O_2485,N_29884,N_29807);
nor UO_2486 (O_2486,N_29910,N_29936);
nand UO_2487 (O_2487,N_29914,N_29974);
and UO_2488 (O_2488,N_29954,N_29836);
nand UO_2489 (O_2489,N_29831,N_29993);
or UO_2490 (O_2490,N_29824,N_29857);
and UO_2491 (O_2491,N_29849,N_29924);
xor UO_2492 (O_2492,N_29941,N_29938);
nand UO_2493 (O_2493,N_29897,N_29933);
or UO_2494 (O_2494,N_29944,N_29974);
and UO_2495 (O_2495,N_29913,N_29989);
nor UO_2496 (O_2496,N_29857,N_29819);
xnor UO_2497 (O_2497,N_29983,N_29861);
or UO_2498 (O_2498,N_29952,N_29886);
and UO_2499 (O_2499,N_29852,N_29844);
nor UO_2500 (O_2500,N_29869,N_29980);
nor UO_2501 (O_2501,N_29911,N_29998);
nor UO_2502 (O_2502,N_29982,N_29867);
nor UO_2503 (O_2503,N_29867,N_29821);
nand UO_2504 (O_2504,N_29858,N_29893);
or UO_2505 (O_2505,N_29982,N_29925);
or UO_2506 (O_2506,N_29848,N_29835);
and UO_2507 (O_2507,N_29841,N_29835);
nand UO_2508 (O_2508,N_29998,N_29851);
nand UO_2509 (O_2509,N_29893,N_29898);
xor UO_2510 (O_2510,N_29928,N_29815);
or UO_2511 (O_2511,N_29802,N_29904);
nand UO_2512 (O_2512,N_29855,N_29957);
xnor UO_2513 (O_2513,N_29828,N_29899);
or UO_2514 (O_2514,N_29942,N_29857);
xnor UO_2515 (O_2515,N_29839,N_29948);
and UO_2516 (O_2516,N_29958,N_29937);
nand UO_2517 (O_2517,N_29914,N_29968);
nor UO_2518 (O_2518,N_29888,N_29934);
nand UO_2519 (O_2519,N_29954,N_29903);
or UO_2520 (O_2520,N_29892,N_29973);
xor UO_2521 (O_2521,N_29937,N_29967);
nand UO_2522 (O_2522,N_29932,N_29836);
or UO_2523 (O_2523,N_29954,N_29802);
nor UO_2524 (O_2524,N_29882,N_29984);
and UO_2525 (O_2525,N_29902,N_29977);
and UO_2526 (O_2526,N_29836,N_29834);
nand UO_2527 (O_2527,N_29923,N_29863);
and UO_2528 (O_2528,N_29980,N_29963);
and UO_2529 (O_2529,N_29929,N_29868);
or UO_2530 (O_2530,N_29925,N_29919);
and UO_2531 (O_2531,N_29934,N_29857);
nand UO_2532 (O_2532,N_29839,N_29909);
or UO_2533 (O_2533,N_29856,N_29986);
or UO_2534 (O_2534,N_29937,N_29963);
xnor UO_2535 (O_2535,N_29904,N_29983);
and UO_2536 (O_2536,N_29959,N_29937);
or UO_2537 (O_2537,N_29923,N_29893);
or UO_2538 (O_2538,N_29952,N_29945);
nor UO_2539 (O_2539,N_29857,N_29908);
nand UO_2540 (O_2540,N_29988,N_29864);
or UO_2541 (O_2541,N_29829,N_29913);
xnor UO_2542 (O_2542,N_29922,N_29936);
xnor UO_2543 (O_2543,N_29819,N_29898);
or UO_2544 (O_2544,N_29985,N_29927);
or UO_2545 (O_2545,N_29835,N_29958);
xnor UO_2546 (O_2546,N_29954,N_29935);
nand UO_2547 (O_2547,N_29878,N_29870);
and UO_2548 (O_2548,N_29955,N_29879);
xor UO_2549 (O_2549,N_29955,N_29977);
xor UO_2550 (O_2550,N_29953,N_29931);
xor UO_2551 (O_2551,N_29822,N_29865);
nand UO_2552 (O_2552,N_29957,N_29939);
nand UO_2553 (O_2553,N_29802,N_29949);
nand UO_2554 (O_2554,N_29873,N_29928);
and UO_2555 (O_2555,N_29886,N_29959);
and UO_2556 (O_2556,N_29823,N_29816);
or UO_2557 (O_2557,N_29884,N_29908);
nand UO_2558 (O_2558,N_29886,N_29823);
nor UO_2559 (O_2559,N_29842,N_29976);
or UO_2560 (O_2560,N_29970,N_29875);
or UO_2561 (O_2561,N_29931,N_29837);
nor UO_2562 (O_2562,N_29951,N_29923);
xnor UO_2563 (O_2563,N_29815,N_29890);
xor UO_2564 (O_2564,N_29853,N_29902);
or UO_2565 (O_2565,N_29953,N_29983);
nand UO_2566 (O_2566,N_29970,N_29801);
nand UO_2567 (O_2567,N_29946,N_29921);
or UO_2568 (O_2568,N_29958,N_29997);
nand UO_2569 (O_2569,N_29875,N_29982);
nand UO_2570 (O_2570,N_29891,N_29849);
or UO_2571 (O_2571,N_29962,N_29940);
xnor UO_2572 (O_2572,N_29992,N_29993);
nor UO_2573 (O_2573,N_29981,N_29888);
and UO_2574 (O_2574,N_29995,N_29966);
xnor UO_2575 (O_2575,N_29889,N_29981);
nor UO_2576 (O_2576,N_29876,N_29860);
xor UO_2577 (O_2577,N_29884,N_29922);
or UO_2578 (O_2578,N_29931,N_29975);
xnor UO_2579 (O_2579,N_29843,N_29956);
or UO_2580 (O_2580,N_29980,N_29989);
nor UO_2581 (O_2581,N_29821,N_29933);
nor UO_2582 (O_2582,N_29958,N_29838);
nand UO_2583 (O_2583,N_29867,N_29926);
or UO_2584 (O_2584,N_29940,N_29926);
xnor UO_2585 (O_2585,N_29880,N_29825);
xor UO_2586 (O_2586,N_29845,N_29961);
and UO_2587 (O_2587,N_29966,N_29806);
xnor UO_2588 (O_2588,N_29881,N_29817);
xor UO_2589 (O_2589,N_29977,N_29821);
or UO_2590 (O_2590,N_29803,N_29936);
xnor UO_2591 (O_2591,N_29842,N_29872);
nor UO_2592 (O_2592,N_29940,N_29849);
xor UO_2593 (O_2593,N_29987,N_29869);
or UO_2594 (O_2594,N_29915,N_29828);
xnor UO_2595 (O_2595,N_29984,N_29811);
nor UO_2596 (O_2596,N_29980,N_29875);
nor UO_2597 (O_2597,N_29896,N_29880);
and UO_2598 (O_2598,N_29903,N_29940);
xor UO_2599 (O_2599,N_29898,N_29826);
xor UO_2600 (O_2600,N_29928,N_29920);
or UO_2601 (O_2601,N_29837,N_29891);
nand UO_2602 (O_2602,N_29900,N_29801);
nand UO_2603 (O_2603,N_29899,N_29996);
or UO_2604 (O_2604,N_29990,N_29836);
or UO_2605 (O_2605,N_29942,N_29846);
xor UO_2606 (O_2606,N_29830,N_29893);
and UO_2607 (O_2607,N_29930,N_29859);
and UO_2608 (O_2608,N_29884,N_29938);
or UO_2609 (O_2609,N_29952,N_29820);
xnor UO_2610 (O_2610,N_29802,N_29920);
and UO_2611 (O_2611,N_29832,N_29929);
nand UO_2612 (O_2612,N_29897,N_29892);
nor UO_2613 (O_2613,N_29888,N_29922);
nor UO_2614 (O_2614,N_29905,N_29877);
nor UO_2615 (O_2615,N_29962,N_29866);
and UO_2616 (O_2616,N_29812,N_29851);
nand UO_2617 (O_2617,N_29848,N_29981);
xor UO_2618 (O_2618,N_29895,N_29905);
nor UO_2619 (O_2619,N_29998,N_29972);
or UO_2620 (O_2620,N_29965,N_29824);
nand UO_2621 (O_2621,N_29985,N_29924);
and UO_2622 (O_2622,N_29969,N_29810);
or UO_2623 (O_2623,N_29807,N_29959);
or UO_2624 (O_2624,N_29979,N_29923);
and UO_2625 (O_2625,N_29908,N_29907);
nand UO_2626 (O_2626,N_29896,N_29899);
xor UO_2627 (O_2627,N_29847,N_29999);
and UO_2628 (O_2628,N_29927,N_29947);
or UO_2629 (O_2629,N_29992,N_29835);
and UO_2630 (O_2630,N_29961,N_29988);
xnor UO_2631 (O_2631,N_29915,N_29961);
or UO_2632 (O_2632,N_29968,N_29820);
xor UO_2633 (O_2633,N_29976,N_29938);
or UO_2634 (O_2634,N_29827,N_29881);
xnor UO_2635 (O_2635,N_29901,N_29938);
or UO_2636 (O_2636,N_29995,N_29976);
nor UO_2637 (O_2637,N_29881,N_29837);
xnor UO_2638 (O_2638,N_29862,N_29883);
nand UO_2639 (O_2639,N_29817,N_29937);
or UO_2640 (O_2640,N_29874,N_29949);
xor UO_2641 (O_2641,N_29834,N_29973);
nor UO_2642 (O_2642,N_29901,N_29932);
nor UO_2643 (O_2643,N_29825,N_29981);
and UO_2644 (O_2644,N_29934,N_29814);
xor UO_2645 (O_2645,N_29908,N_29894);
xnor UO_2646 (O_2646,N_29823,N_29829);
nor UO_2647 (O_2647,N_29878,N_29898);
nor UO_2648 (O_2648,N_29868,N_29873);
and UO_2649 (O_2649,N_29959,N_29835);
nand UO_2650 (O_2650,N_29849,N_29983);
nor UO_2651 (O_2651,N_29856,N_29944);
and UO_2652 (O_2652,N_29974,N_29844);
nor UO_2653 (O_2653,N_29809,N_29918);
nor UO_2654 (O_2654,N_29996,N_29994);
and UO_2655 (O_2655,N_29829,N_29842);
and UO_2656 (O_2656,N_29975,N_29991);
xor UO_2657 (O_2657,N_29944,N_29844);
nor UO_2658 (O_2658,N_29824,N_29818);
nand UO_2659 (O_2659,N_29969,N_29873);
xnor UO_2660 (O_2660,N_29833,N_29923);
and UO_2661 (O_2661,N_29828,N_29822);
and UO_2662 (O_2662,N_29803,N_29965);
and UO_2663 (O_2663,N_29811,N_29861);
and UO_2664 (O_2664,N_29831,N_29861);
nor UO_2665 (O_2665,N_29968,N_29881);
xor UO_2666 (O_2666,N_29860,N_29813);
xnor UO_2667 (O_2667,N_29933,N_29932);
or UO_2668 (O_2668,N_29872,N_29813);
xor UO_2669 (O_2669,N_29800,N_29893);
and UO_2670 (O_2670,N_29845,N_29925);
nand UO_2671 (O_2671,N_29941,N_29916);
and UO_2672 (O_2672,N_29875,N_29908);
nor UO_2673 (O_2673,N_29807,N_29902);
and UO_2674 (O_2674,N_29887,N_29978);
nand UO_2675 (O_2675,N_29863,N_29927);
xor UO_2676 (O_2676,N_29877,N_29987);
xnor UO_2677 (O_2677,N_29805,N_29979);
or UO_2678 (O_2678,N_29800,N_29852);
nor UO_2679 (O_2679,N_29857,N_29975);
nand UO_2680 (O_2680,N_29891,N_29935);
or UO_2681 (O_2681,N_29952,N_29962);
nand UO_2682 (O_2682,N_29924,N_29815);
nor UO_2683 (O_2683,N_29982,N_29934);
nor UO_2684 (O_2684,N_29870,N_29934);
or UO_2685 (O_2685,N_29901,N_29968);
and UO_2686 (O_2686,N_29851,N_29837);
nand UO_2687 (O_2687,N_29813,N_29842);
nor UO_2688 (O_2688,N_29860,N_29907);
xor UO_2689 (O_2689,N_29999,N_29996);
or UO_2690 (O_2690,N_29948,N_29821);
nand UO_2691 (O_2691,N_29835,N_29940);
nor UO_2692 (O_2692,N_29916,N_29981);
nand UO_2693 (O_2693,N_29937,N_29842);
or UO_2694 (O_2694,N_29851,N_29940);
or UO_2695 (O_2695,N_29846,N_29892);
or UO_2696 (O_2696,N_29981,N_29919);
nand UO_2697 (O_2697,N_29949,N_29849);
and UO_2698 (O_2698,N_29944,N_29847);
and UO_2699 (O_2699,N_29975,N_29917);
or UO_2700 (O_2700,N_29926,N_29907);
xnor UO_2701 (O_2701,N_29971,N_29970);
and UO_2702 (O_2702,N_29825,N_29943);
and UO_2703 (O_2703,N_29804,N_29821);
nor UO_2704 (O_2704,N_29912,N_29856);
nand UO_2705 (O_2705,N_29990,N_29870);
or UO_2706 (O_2706,N_29984,N_29836);
and UO_2707 (O_2707,N_29956,N_29895);
xnor UO_2708 (O_2708,N_29953,N_29967);
nor UO_2709 (O_2709,N_29941,N_29856);
nor UO_2710 (O_2710,N_29850,N_29903);
nor UO_2711 (O_2711,N_29809,N_29928);
and UO_2712 (O_2712,N_29803,N_29941);
nand UO_2713 (O_2713,N_29823,N_29943);
nor UO_2714 (O_2714,N_29886,N_29854);
or UO_2715 (O_2715,N_29990,N_29873);
nand UO_2716 (O_2716,N_29932,N_29881);
nor UO_2717 (O_2717,N_29884,N_29858);
or UO_2718 (O_2718,N_29834,N_29868);
nand UO_2719 (O_2719,N_29868,N_29923);
and UO_2720 (O_2720,N_29849,N_29905);
xor UO_2721 (O_2721,N_29934,N_29951);
and UO_2722 (O_2722,N_29881,N_29934);
nor UO_2723 (O_2723,N_29830,N_29803);
or UO_2724 (O_2724,N_29996,N_29800);
or UO_2725 (O_2725,N_29863,N_29965);
and UO_2726 (O_2726,N_29894,N_29873);
nor UO_2727 (O_2727,N_29871,N_29999);
nor UO_2728 (O_2728,N_29926,N_29864);
and UO_2729 (O_2729,N_29981,N_29948);
and UO_2730 (O_2730,N_29838,N_29808);
and UO_2731 (O_2731,N_29978,N_29818);
xor UO_2732 (O_2732,N_29880,N_29931);
or UO_2733 (O_2733,N_29897,N_29875);
or UO_2734 (O_2734,N_29838,N_29977);
nor UO_2735 (O_2735,N_29823,N_29854);
nand UO_2736 (O_2736,N_29937,N_29944);
and UO_2737 (O_2737,N_29824,N_29957);
nand UO_2738 (O_2738,N_29933,N_29913);
xor UO_2739 (O_2739,N_29912,N_29870);
or UO_2740 (O_2740,N_29918,N_29843);
or UO_2741 (O_2741,N_29830,N_29899);
and UO_2742 (O_2742,N_29839,N_29966);
and UO_2743 (O_2743,N_29914,N_29851);
nand UO_2744 (O_2744,N_29819,N_29978);
nand UO_2745 (O_2745,N_29867,N_29960);
or UO_2746 (O_2746,N_29910,N_29814);
and UO_2747 (O_2747,N_29877,N_29950);
nor UO_2748 (O_2748,N_29910,N_29914);
xor UO_2749 (O_2749,N_29986,N_29936);
nand UO_2750 (O_2750,N_29927,N_29912);
or UO_2751 (O_2751,N_29812,N_29839);
nand UO_2752 (O_2752,N_29942,N_29842);
or UO_2753 (O_2753,N_29917,N_29946);
xnor UO_2754 (O_2754,N_29909,N_29891);
or UO_2755 (O_2755,N_29879,N_29924);
nor UO_2756 (O_2756,N_29882,N_29820);
nor UO_2757 (O_2757,N_29911,N_29856);
nor UO_2758 (O_2758,N_29900,N_29883);
or UO_2759 (O_2759,N_29896,N_29808);
nand UO_2760 (O_2760,N_29894,N_29891);
and UO_2761 (O_2761,N_29994,N_29904);
and UO_2762 (O_2762,N_29838,N_29994);
or UO_2763 (O_2763,N_29960,N_29969);
nor UO_2764 (O_2764,N_29966,N_29865);
xnor UO_2765 (O_2765,N_29991,N_29900);
xnor UO_2766 (O_2766,N_29817,N_29859);
and UO_2767 (O_2767,N_29828,N_29982);
and UO_2768 (O_2768,N_29890,N_29900);
nand UO_2769 (O_2769,N_29978,N_29990);
nand UO_2770 (O_2770,N_29892,N_29954);
nor UO_2771 (O_2771,N_29811,N_29837);
and UO_2772 (O_2772,N_29899,N_29890);
and UO_2773 (O_2773,N_29901,N_29914);
or UO_2774 (O_2774,N_29889,N_29993);
or UO_2775 (O_2775,N_29994,N_29963);
and UO_2776 (O_2776,N_29937,N_29881);
or UO_2777 (O_2777,N_29842,N_29840);
or UO_2778 (O_2778,N_29848,N_29959);
or UO_2779 (O_2779,N_29878,N_29851);
or UO_2780 (O_2780,N_29893,N_29892);
nand UO_2781 (O_2781,N_29934,N_29958);
and UO_2782 (O_2782,N_29938,N_29839);
and UO_2783 (O_2783,N_29966,N_29872);
or UO_2784 (O_2784,N_29961,N_29919);
nand UO_2785 (O_2785,N_29954,N_29870);
nor UO_2786 (O_2786,N_29830,N_29812);
and UO_2787 (O_2787,N_29879,N_29847);
and UO_2788 (O_2788,N_29973,N_29878);
nand UO_2789 (O_2789,N_29899,N_29947);
nand UO_2790 (O_2790,N_29945,N_29872);
or UO_2791 (O_2791,N_29930,N_29845);
nand UO_2792 (O_2792,N_29805,N_29829);
xor UO_2793 (O_2793,N_29822,N_29827);
nor UO_2794 (O_2794,N_29872,N_29905);
nand UO_2795 (O_2795,N_29970,N_29951);
nor UO_2796 (O_2796,N_29906,N_29846);
nor UO_2797 (O_2797,N_29969,N_29987);
nand UO_2798 (O_2798,N_29857,N_29812);
nand UO_2799 (O_2799,N_29861,N_29894);
and UO_2800 (O_2800,N_29964,N_29864);
and UO_2801 (O_2801,N_29805,N_29893);
nor UO_2802 (O_2802,N_29924,N_29998);
nand UO_2803 (O_2803,N_29838,N_29801);
xor UO_2804 (O_2804,N_29967,N_29962);
nand UO_2805 (O_2805,N_29811,N_29918);
xor UO_2806 (O_2806,N_29918,N_29951);
xor UO_2807 (O_2807,N_29882,N_29826);
and UO_2808 (O_2808,N_29924,N_29962);
nand UO_2809 (O_2809,N_29976,N_29979);
or UO_2810 (O_2810,N_29852,N_29912);
nor UO_2811 (O_2811,N_29848,N_29932);
nand UO_2812 (O_2812,N_29951,N_29960);
xnor UO_2813 (O_2813,N_29891,N_29828);
nand UO_2814 (O_2814,N_29985,N_29940);
xnor UO_2815 (O_2815,N_29996,N_29901);
and UO_2816 (O_2816,N_29884,N_29800);
or UO_2817 (O_2817,N_29878,N_29864);
or UO_2818 (O_2818,N_29807,N_29899);
or UO_2819 (O_2819,N_29877,N_29973);
and UO_2820 (O_2820,N_29853,N_29914);
xor UO_2821 (O_2821,N_29999,N_29805);
xor UO_2822 (O_2822,N_29969,N_29909);
nand UO_2823 (O_2823,N_29827,N_29875);
nor UO_2824 (O_2824,N_29884,N_29849);
xor UO_2825 (O_2825,N_29964,N_29856);
nor UO_2826 (O_2826,N_29918,N_29991);
nor UO_2827 (O_2827,N_29996,N_29842);
nor UO_2828 (O_2828,N_29857,N_29849);
nor UO_2829 (O_2829,N_29920,N_29825);
or UO_2830 (O_2830,N_29908,N_29994);
and UO_2831 (O_2831,N_29821,N_29897);
nor UO_2832 (O_2832,N_29866,N_29876);
or UO_2833 (O_2833,N_29936,N_29981);
nor UO_2834 (O_2834,N_29991,N_29840);
nand UO_2835 (O_2835,N_29816,N_29866);
xnor UO_2836 (O_2836,N_29893,N_29811);
nor UO_2837 (O_2837,N_29974,N_29947);
or UO_2838 (O_2838,N_29864,N_29872);
nand UO_2839 (O_2839,N_29859,N_29944);
nand UO_2840 (O_2840,N_29885,N_29990);
or UO_2841 (O_2841,N_29821,N_29970);
or UO_2842 (O_2842,N_29926,N_29863);
nor UO_2843 (O_2843,N_29951,N_29917);
or UO_2844 (O_2844,N_29962,N_29994);
nor UO_2845 (O_2845,N_29802,N_29999);
xor UO_2846 (O_2846,N_29997,N_29922);
nand UO_2847 (O_2847,N_29845,N_29915);
xor UO_2848 (O_2848,N_29825,N_29917);
xor UO_2849 (O_2849,N_29834,N_29966);
xor UO_2850 (O_2850,N_29924,N_29982);
or UO_2851 (O_2851,N_29966,N_29956);
nor UO_2852 (O_2852,N_29837,N_29917);
or UO_2853 (O_2853,N_29919,N_29998);
nor UO_2854 (O_2854,N_29841,N_29848);
and UO_2855 (O_2855,N_29890,N_29878);
nor UO_2856 (O_2856,N_29902,N_29987);
and UO_2857 (O_2857,N_29961,N_29877);
nand UO_2858 (O_2858,N_29945,N_29833);
nand UO_2859 (O_2859,N_29829,N_29801);
or UO_2860 (O_2860,N_29818,N_29838);
nand UO_2861 (O_2861,N_29964,N_29933);
or UO_2862 (O_2862,N_29985,N_29863);
nand UO_2863 (O_2863,N_29982,N_29832);
and UO_2864 (O_2864,N_29813,N_29801);
nand UO_2865 (O_2865,N_29953,N_29826);
xnor UO_2866 (O_2866,N_29975,N_29809);
xnor UO_2867 (O_2867,N_29867,N_29830);
nor UO_2868 (O_2868,N_29956,N_29905);
nand UO_2869 (O_2869,N_29880,N_29961);
or UO_2870 (O_2870,N_29825,N_29890);
nand UO_2871 (O_2871,N_29988,N_29994);
nor UO_2872 (O_2872,N_29934,N_29906);
xor UO_2873 (O_2873,N_29801,N_29952);
xor UO_2874 (O_2874,N_29887,N_29851);
nor UO_2875 (O_2875,N_29930,N_29862);
nor UO_2876 (O_2876,N_29874,N_29890);
nand UO_2877 (O_2877,N_29865,N_29954);
or UO_2878 (O_2878,N_29870,N_29821);
and UO_2879 (O_2879,N_29822,N_29931);
xor UO_2880 (O_2880,N_29926,N_29862);
and UO_2881 (O_2881,N_29874,N_29992);
xnor UO_2882 (O_2882,N_29814,N_29909);
and UO_2883 (O_2883,N_29987,N_29973);
nand UO_2884 (O_2884,N_29875,N_29800);
and UO_2885 (O_2885,N_29818,N_29954);
xnor UO_2886 (O_2886,N_29901,N_29908);
or UO_2887 (O_2887,N_29813,N_29901);
nor UO_2888 (O_2888,N_29934,N_29923);
or UO_2889 (O_2889,N_29815,N_29958);
xor UO_2890 (O_2890,N_29846,N_29898);
or UO_2891 (O_2891,N_29976,N_29876);
xor UO_2892 (O_2892,N_29913,N_29858);
xnor UO_2893 (O_2893,N_29981,N_29819);
xnor UO_2894 (O_2894,N_29966,N_29972);
nand UO_2895 (O_2895,N_29975,N_29833);
nor UO_2896 (O_2896,N_29858,N_29977);
nor UO_2897 (O_2897,N_29824,N_29968);
nor UO_2898 (O_2898,N_29831,N_29849);
nor UO_2899 (O_2899,N_29970,N_29879);
nor UO_2900 (O_2900,N_29882,N_29896);
xor UO_2901 (O_2901,N_29950,N_29834);
or UO_2902 (O_2902,N_29935,N_29955);
nand UO_2903 (O_2903,N_29850,N_29853);
or UO_2904 (O_2904,N_29911,N_29814);
or UO_2905 (O_2905,N_29929,N_29853);
nor UO_2906 (O_2906,N_29815,N_29908);
xor UO_2907 (O_2907,N_29841,N_29821);
or UO_2908 (O_2908,N_29826,N_29955);
and UO_2909 (O_2909,N_29954,N_29855);
and UO_2910 (O_2910,N_29979,N_29989);
nor UO_2911 (O_2911,N_29824,N_29905);
nand UO_2912 (O_2912,N_29900,N_29868);
nand UO_2913 (O_2913,N_29810,N_29951);
and UO_2914 (O_2914,N_29811,N_29967);
xor UO_2915 (O_2915,N_29921,N_29856);
xnor UO_2916 (O_2916,N_29959,N_29939);
nand UO_2917 (O_2917,N_29951,N_29820);
or UO_2918 (O_2918,N_29862,N_29932);
nor UO_2919 (O_2919,N_29844,N_29989);
or UO_2920 (O_2920,N_29832,N_29897);
or UO_2921 (O_2921,N_29976,N_29873);
xnor UO_2922 (O_2922,N_29865,N_29855);
nor UO_2923 (O_2923,N_29832,N_29816);
xor UO_2924 (O_2924,N_29998,N_29852);
or UO_2925 (O_2925,N_29811,N_29871);
nand UO_2926 (O_2926,N_29950,N_29929);
nor UO_2927 (O_2927,N_29958,N_29868);
and UO_2928 (O_2928,N_29882,N_29940);
nor UO_2929 (O_2929,N_29812,N_29988);
and UO_2930 (O_2930,N_29806,N_29947);
or UO_2931 (O_2931,N_29862,N_29898);
or UO_2932 (O_2932,N_29848,N_29875);
nand UO_2933 (O_2933,N_29801,N_29837);
xor UO_2934 (O_2934,N_29903,N_29985);
or UO_2935 (O_2935,N_29827,N_29975);
xor UO_2936 (O_2936,N_29829,N_29898);
and UO_2937 (O_2937,N_29924,N_29865);
nand UO_2938 (O_2938,N_29864,N_29884);
or UO_2939 (O_2939,N_29876,N_29886);
xnor UO_2940 (O_2940,N_29936,N_29977);
xnor UO_2941 (O_2941,N_29907,N_29875);
nand UO_2942 (O_2942,N_29995,N_29856);
nand UO_2943 (O_2943,N_29952,N_29890);
and UO_2944 (O_2944,N_29849,N_29922);
or UO_2945 (O_2945,N_29818,N_29837);
nor UO_2946 (O_2946,N_29804,N_29823);
and UO_2947 (O_2947,N_29921,N_29898);
xor UO_2948 (O_2948,N_29914,N_29958);
and UO_2949 (O_2949,N_29916,N_29873);
nand UO_2950 (O_2950,N_29806,N_29831);
or UO_2951 (O_2951,N_29873,N_29828);
or UO_2952 (O_2952,N_29969,N_29982);
or UO_2953 (O_2953,N_29807,N_29914);
xnor UO_2954 (O_2954,N_29863,N_29954);
and UO_2955 (O_2955,N_29824,N_29817);
nor UO_2956 (O_2956,N_29903,N_29833);
xor UO_2957 (O_2957,N_29881,N_29946);
xnor UO_2958 (O_2958,N_29912,N_29851);
nor UO_2959 (O_2959,N_29918,N_29923);
and UO_2960 (O_2960,N_29992,N_29902);
nand UO_2961 (O_2961,N_29818,N_29807);
xnor UO_2962 (O_2962,N_29833,N_29816);
or UO_2963 (O_2963,N_29930,N_29986);
and UO_2964 (O_2964,N_29908,N_29810);
nand UO_2965 (O_2965,N_29980,N_29805);
nor UO_2966 (O_2966,N_29931,N_29882);
xor UO_2967 (O_2967,N_29865,N_29958);
or UO_2968 (O_2968,N_29829,N_29946);
xor UO_2969 (O_2969,N_29922,N_29871);
xnor UO_2970 (O_2970,N_29904,N_29824);
xnor UO_2971 (O_2971,N_29861,N_29921);
or UO_2972 (O_2972,N_29931,N_29987);
and UO_2973 (O_2973,N_29841,N_29938);
and UO_2974 (O_2974,N_29826,N_29853);
nor UO_2975 (O_2975,N_29945,N_29854);
or UO_2976 (O_2976,N_29859,N_29976);
nor UO_2977 (O_2977,N_29810,N_29961);
nand UO_2978 (O_2978,N_29818,N_29809);
or UO_2979 (O_2979,N_29981,N_29903);
nand UO_2980 (O_2980,N_29910,N_29822);
nor UO_2981 (O_2981,N_29830,N_29931);
and UO_2982 (O_2982,N_29987,N_29998);
nand UO_2983 (O_2983,N_29933,N_29974);
nor UO_2984 (O_2984,N_29815,N_29835);
xnor UO_2985 (O_2985,N_29927,N_29987);
nand UO_2986 (O_2986,N_29977,N_29856);
nand UO_2987 (O_2987,N_29851,N_29922);
nor UO_2988 (O_2988,N_29904,N_29981);
nand UO_2989 (O_2989,N_29887,N_29815);
or UO_2990 (O_2990,N_29824,N_29844);
nor UO_2991 (O_2991,N_29822,N_29826);
nand UO_2992 (O_2992,N_29967,N_29925);
nor UO_2993 (O_2993,N_29904,N_29807);
or UO_2994 (O_2994,N_29835,N_29968);
xnor UO_2995 (O_2995,N_29861,N_29920);
nand UO_2996 (O_2996,N_29809,N_29983);
nand UO_2997 (O_2997,N_29992,N_29961);
nor UO_2998 (O_2998,N_29925,N_29988);
and UO_2999 (O_2999,N_29816,N_29995);
nor UO_3000 (O_3000,N_29980,N_29852);
xnor UO_3001 (O_3001,N_29998,N_29854);
and UO_3002 (O_3002,N_29854,N_29861);
xnor UO_3003 (O_3003,N_29829,N_29889);
nor UO_3004 (O_3004,N_29849,N_29859);
nor UO_3005 (O_3005,N_29921,N_29814);
nand UO_3006 (O_3006,N_29835,N_29970);
or UO_3007 (O_3007,N_29997,N_29848);
nor UO_3008 (O_3008,N_29946,N_29803);
nor UO_3009 (O_3009,N_29881,N_29863);
nor UO_3010 (O_3010,N_29875,N_29855);
or UO_3011 (O_3011,N_29880,N_29876);
or UO_3012 (O_3012,N_29993,N_29801);
and UO_3013 (O_3013,N_29965,N_29913);
and UO_3014 (O_3014,N_29936,N_29902);
xor UO_3015 (O_3015,N_29810,N_29861);
or UO_3016 (O_3016,N_29942,N_29879);
or UO_3017 (O_3017,N_29858,N_29947);
nand UO_3018 (O_3018,N_29807,N_29868);
and UO_3019 (O_3019,N_29930,N_29842);
and UO_3020 (O_3020,N_29900,N_29851);
nand UO_3021 (O_3021,N_29912,N_29831);
or UO_3022 (O_3022,N_29891,N_29952);
nand UO_3023 (O_3023,N_29933,N_29968);
and UO_3024 (O_3024,N_29821,N_29843);
or UO_3025 (O_3025,N_29996,N_29962);
and UO_3026 (O_3026,N_29976,N_29921);
and UO_3027 (O_3027,N_29957,N_29822);
xor UO_3028 (O_3028,N_29861,N_29907);
or UO_3029 (O_3029,N_29945,N_29847);
nor UO_3030 (O_3030,N_29815,N_29882);
nand UO_3031 (O_3031,N_29815,N_29912);
and UO_3032 (O_3032,N_29980,N_29826);
nand UO_3033 (O_3033,N_29928,N_29932);
or UO_3034 (O_3034,N_29995,N_29807);
nor UO_3035 (O_3035,N_29980,N_29996);
nor UO_3036 (O_3036,N_29807,N_29809);
nor UO_3037 (O_3037,N_29976,N_29863);
nor UO_3038 (O_3038,N_29815,N_29869);
nand UO_3039 (O_3039,N_29919,N_29948);
or UO_3040 (O_3040,N_29843,N_29913);
nand UO_3041 (O_3041,N_29879,N_29806);
or UO_3042 (O_3042,N_29841,N_29868);
nor UO_3043 (O_3043,N_29965,N_29956);
or UO_3044 (O_3044,N_29963,N_29885);
xor UO_3045 (O_3045,N_29957,N_29872);
xnor UO_3046 (O_3046,N_29900,N_29800);
xor UO_3047 (O_3047,N_29805,N_29993);
nand UO_3048 (O_3048,N_29984,N_29948);
nor UO_3049 (O_3049,N_29883,N_29826);
nand UO_3050 (O_3050,N_29893,N_29935);
nor UO_3051 (O_3051,N_29819,N_29965);
nor UO_3052 (O_3052,N_29814,N_29994);
nand UO_3053 (O_3053,N_29972,N_29997);
nor UO_3054 (O_3054,N_29820,N_29879);
xor UO_3055 (O_3055,N_29997,N_29800);
xor UO_3056 (O_3056,N_29800,N_29857);
nor UO_3057 (O_3057,N_29850,N_29936);
xor UO_3058 (O_3058,N_29945,N_29874);
nand UO_3059 (O_3059,N_29878,N_29802);
or UO_3060 (O_3060,N_29936,N_29825);
or UO_3061 (O_3061,N_29887,N_29813);
and UO_3062 (O_3062,N_29811,N_29975);
nand UO_3063 (O_3063,N_29952,N_29854);
xor UO_3064 (O_3064,N_29800,N_29842);
xor UO_3065 (O_3065,N_29879,N_29953);
nand UO_3066 (O_3066,N_29988,N_29975);
and UO_3067 (O_3067,N_29804,N_29889);
or UO_3068 (O_3068,N_29890,N_29881);
and UO_3069 (O_3069,N_29921,N_29936);
nand UO_3070 (O_3070,N_29882,N_29835);
and UO_3071 (O_3071,N_29956,N_29833);
and UO_3072 (O_3072,N_29975,N_29945);
xor UO_3073 (O_3073,N_29981,N_29846);
nand UO_3074 (O_3074,N_29835,N_29948);
xor UO_3075 (O_3075,N_29866,N_29895);
nand UO_3076 (O_3076,N_29961,N_29921);
nand UO_3077 (O_3077,N_29806,N_29814);
xnor UO_3078 (O_3078,N_29988,N_29990);
nor UO_3079 (O_3079,N_29895,N_29804);
xnor UO_3080 (O_3080,N_29945,N_29917);
and UO_3081 (O_3081,N_29871,N_29882);
or UO_3082 (O_3082,N_29981,N_29991);
or UO_3083 (O_3083,N_29953,N_29968);
and UO_3084 (O_3084,N_29983,N_29813);
or UO_3085 (O_3085,N_29935,N_29831);
nor UO_3086 (O_3086,N_29952,N_29857);
and UO_3087 (O_3087,N_29862,N_29958);
or UO_3088 (O_3088,N_29892,N_29839);
xor UO_3089 (O_3089,N_29982,N_29827);
or UO_3090 (O_3090,N_29805,N_29881);
xor UO_3091 (O_3091,N_29932,N_29945);
nor UO_3092 (O_3092,N_29805,N_29932);
nor UO_3093 (O_3093,N_29840,N_29839);
xor UO_3094 (O_3094,N_29985,N_29809);
and UO_3095 (O_3095,N_29934,N_29994);
and UO_3096 (O_3096,N_29892,N_29937);
nor UO_3097 (O_3097,N_29870,N_29890);
and UO_3098 (O_3098,N_29999,N_29822);
nor UO_3099 (O_3099,N_29883,N_29943);
nor UO_3100 (O_3100,N_29811,N_29966);
xnor UO_3101 (O_3101,N_29990,N_29806);
nor UO_3102 (O_3102,N_29871,N_29908);
xor UO_3103 (O_3103,N_29843,N_29902);
or UO_3104 (O_3104,N_29922,N_29802);
and UO_3105 (O_3105,N_29882,N_29953);
and UO_3106 (O_3106,N_29881,N_29818);
nand UO_3107 (O_3107,N_29965,N_29946);
or UO_3108 (O_3108,N_29915,N_29819);
nor UO_3109 (O_3109,N_29915,N_29846);
nand UO_3110 (O_3110,N_29870,N_29822);
xor UO_3111 (O_3111,N_29857,N_29902);
nor UO_3112 (O_3112,N_29999,N_29819);
nor UO_3113 (O_3113,N_29849,N_29985);
and UO_3114 (O_3114,N_29972,N_29933);
and UO_3115 (O_3115,N_29863,N_29825);
and UO_3116 (O_3116,N_29965,N_29845);
and UO_3117 (O_3117,N_29852,N_29883);
nor UO_3118 (O_3118,N_29963,N_29971);
and UO_3119 (O_3119,N_29834,N_29890);
nor UO_3120 (O_3120,N_29887,N_29811);
and UO_3121 (O_3121,N_29993,N_29997);
or UO_3122 (O_3122,N_29809,N_29886);
xnor UO_3123 (O_3123,N_29959,N_29936);
and UO_3124 (O_3124,N_29982,N_29895);
xnor UO_3125 (O_3125,N_29956,N_29987);
xnor UO_3126 (O_3126,N_29910,N_29890);
and UO_3127 (O_3127,N_29906,N_29932);
xnor UO_3128 (O_3128,N_29989,N_29936);
and UO_3129 (O_3129,N_29871,N_29987);
or UO_3130 (O_3130,N_29823,N_29960);
or UO_3131 (O_3131,N_29845,N_29977);
xor UO_3132 (O_3132,N_29959,N_29805);
nor UO_3133 (O_3133,N_29817,N_29999);
nor UO_3134 (O_3134,N_29826,N_29974);
nand UO_3135 (O_3135,N_29809,N_29938);
or UO_3136 (O_3136,N_29980,N_29979);
xnor UO_3137 (O_3137,N_29922,N_29906);
or UO_3138 (O_3138,N_29815,N_29907);
xnor UO_3139 (O_3139,N_29801,N_29975);
or UO_3140 (O_3140,N_29925,N_29817);
or UO_3141 (O_3141,N_29969,N_29954);
or UO_3142 (O_3142,N_29951,N_29896);
or UO_3143 (O_3143,N_29858,N_29949);
and UO_3144 (O_3144,N_29937,N_29867);
and UO_3145 (O_3145,N_29813,N_29998);
nor UO_3146 (O_3146,N_29950,N_29869);
or UO_3147 (O_3147,N_29816,N_29891);
xor UO_3148 (O_3148,N_29895,N_29993);
or UO_3149 (O_3149,N_29909,N_29846);
and UO_3150 (O_3150,N_29859,N_29945);
xor UO_3151 (O_3151,N_29849,N_29838);
xor UO_3152 (O_3152,N_29801,N_29800);
nand UO_3153 (O_3153,N_29972,N_29893);
nand UO_3154 (O_3154,N_29844,N_29980);
xor UO_3155 (O_3155,N_29887,N_29921);
xor UO_3156 (O_3156,N_29980,N_29950);
and UO_3157 (O_3157,N_29852,N_29832);
nor UO_3158 (O_3158,N_29943,N_29971);
nand UO_3159 (O_3159,N_29856,N_29967);
or UO_3160 (O_3160,N_29889,N_29923);
nand UO_3161 (O_3161,N_29999,N_29894);
or UO_3162 (O_3162,N_29930,N_29922);
xnor UO_3163 (O_3163,N_29894,N_29811);
and UO_3164 (O_3164,N_29947,N_29817);
or UO_3165 (O_3165,N_29801,N_29969);
nor UO_3166 (O_3166,N_29828,N_29933);
nor UO_3167 (O_3167,N_29851,N_29946);
nand UO_3168 (O_3168,N_29882,N_29946);
or UO_3169 (O_3169,N_29984,N_29928);
and UO_3170 (O_3170,N_29861,N_29916);
and UO_3171 (O_3171,N_29853,N_29965);
nand UO_3172 (O_3172,N_29826,N_29920);
nand UO_3173 (O_3173,N_29895,N_29898);
and UO_3174 (O_3174,N_29989,N_29891);
xnor UO_3175 (O_3175,N_29880,N_29819);
nand UO_3176 (O_3176,N_29983,N_29858);
nor UO_3177 (O_3177,N_29933,N_29801);
or UO_3178 (O_3178,N_29964,N_29830);
or UO_3179 (O_3179,N_29893,N_29835);
nor UO_3180 (O_3180,N_29914,N_29814);
nand UO_3181 (O_3181,N_29840,N_29934);
and UO_3182 (O_3182,N_29907,N_29980);
nand UO_3183 (O_3183,N_29822,N_29965);
and UO_3184 (O_3184,N_29845,N_29816);
nand UO_3185 (O_3185,N_29981,N_29873);
nor UO_3186 (O_3186,N_29990,N_29947);
nor UO_3187 (O_3187,N_29869,N_29965);
nor UO_3188 (O_3188,N_29848,N_29914);
nor UO_3189 (O_3189,N_29856,N_29813);
xnor UO_3190 (O_3190,N_29943,N_29929);
nand UO_3191 (O_3191,N_29962,N_29867);
or UO_3192 (O_3192,N_29851,N_29841);
xnor UO_3193 (O_3193,N_29808,N_29957);
xnor UO_3194 (O_3194,N_29909,N_29847);
nand UO_3195 (O_3195,N_29834,N_29817);
xor UO_3196 (O_3196,N_29898,N_29913);
xor UO_3197 (O_3197,N_29863,N_29891);
and UO_3198 (O_3198,N_29975,N_29864);
nand UO_3199 (O_3199,N_29963,N_29918);
xor UO_3200 (O_3200,N_29834,N_29906);
nand UO_3201 (O_3201,N_29980,N_29924);
or UO_3202 (O_3202,N_29987,N_29912);
nand UO_3203 (O_3203,N_29878,N_29958);
nor UO_3204 (O_3204,N_29920,N_29869);
xnor UO_3205 (O_3205,N_29999,N_29952);
and UO_3206 (O_3206,N_29951,N_29959);
and UO_3207 (O_3207,N_29996,N_29820);
nand UO_3208 (O_3208,N_29812,N_29923);
or UO_3209 (O_3209,N_29991,N_29843);
nor UO_3210 (O_3210,N_29804,N_29932);
nor UO_3211 (O_3211,N_29993,N_29868);
xor UO_3212 (O_3212,N_29862,N_29915);
nand UO_3213 (O_3213,N_29816,N_29985);
nand UO_3214 (O_3214,N_29958,N_29996);
nand UO_3215 (O_3215,N_29925,N_29801);
nand UO_3216 (O_3216,N_29892,N_29930);
and UO_3217 (O_3217,N_29841,N_29913);
and UO_3218 (O_3218,N_29916,N_29851);
nand UO_3219 (O_3219,N_29933,N_29904);
or UO_3220 (O_3220,N_29862,N_29931);
nor UO_3221 (O_3221,N_29958,N_29833);
or UO_3222 (O_3222,N_29888,N_29853);
or UO_3223 (O_3223,N_29810,N_29891);
and UO_3224 (O_3224,N_29934,N_29811);
or UO_3225 (O_3225,N_29844,N_29826);
or UO_3226 (O_3226,N_29872,N_29973);
xnor UO_3227 (O_3227,N_29899,N_29878);
or UO_3228 (O_3228,N_29904,N_29965);
and UO_3229 (O_3229,N_29955,N_29985);
or UO_3230 (O_3230,N_29951,N_29893);
nand UO_3231 (O_3231,N_29933,N_29825);
and UO_3232 (O_3232,N_29897,N_29935);
or UO_3233 (O_3233,N_29974,N_29918);
or UO_3234 (O_3234,N_29927,N_29940);
or UO_3235 (O_3235,N_29855,N_29982);
xor UO_3236 (O_3236,N_29971,N_29955);
and UO_3237 (O_3237,N_29843,N_29851);
and UO_3238 (O_3238,N_29833,N_29879);
nand UO_3239 (O_3239,N_29911,N_29949);
or UO_3240 (O_3240,N_29994,N_29917);
nand UO_3241 (O_3241,N_29977,N_29873);
or UO_3242 (O_3242,N_29932,N_29817);
nand UO_3243 (O_3243,N_29901,N_29823);
or UO_3244 (O_3244,N_29900,N_29829);
or UO_3245 (O_3245,N_29885,N_29946);
xor UO_3246 (O_3246,N_29913,N_29957);
or UO_3247 (O_3247,N_29883,N_29877);
nand UO_3248 (O_3248,N_29885,N_29924);
and UO_3249 (O_3249,N_29931,N_29801);
nor UO_3250 (O_3250,N_29884,N_29844);
xor UO_3251 (O_3251,N_29906,N_29963);
nor UO_3252 (O_3252,N_29825,N_29834);
nand UO_3253 (O_3253,N_29819,N_29918);
or UO_3254 (O_3254,N_29966,N_29863);
or UO_3255 (O_3255,N_29860,N_29851);
nor UO_3256 (O_3256,N_29802,N_29858);
nor UO_3257 (O_3257,N_29844,N_29819);
and UO_3258 (O_3258,N_29939,N_29962);
nor UO_3259 (O_3259,N_29909,N_29801);
nand UO_3260 (O_3260,N_29975,N_29919);
xnor UO_3261 (O_3261,N_29960,N_29884);
xnor UO_3262 (O_3262,N_29983,N_29987);
xor UO_3263 (O_3263,N_29959,N_29860);
nand UO_3264 (O_3264,N_29971,N_29863);
xnor UO_3265 (O_3265,N_29946,N_29985);
or UO_3266 (O_3266,N_29956,N_29880);
nand UO_3267 (O_3267,N_29896,N_29828);
or UO_3268 (O_3268,N_29860,N_29842);
xor UO_3269 (O_3269,N_29983,N_29974);
xnor UO_3270 (O_3270,N_29810,N_29814);
nand UO_3271 (O_3271,N_29825,N_29925);
and UO_3272 (O_3272,N_29903,N_29946);
nor UO_3273 (O_3273,N_29992,N_29841);
xor UO_3274 (O_3274,N_29948,N_29888);
nor UO_3275 (O_3275,N_29821,N_29903);
or UO_3276 (O_3276,N_29846,N_29962);
or UO_3277 (O_3277,N_29894,N_29867);
and UO_3278 (O_3278,N_29814,N_29870);
and UO_3279 (O_3279,N_29942,N_29996);
and UO_3280 (O_3280,N_29833,N_29963);
xnor UO_3281 (O_3281,N_29912,N_29980);
xnor UO_3282 (O_3282,N_29969,N_29965);
and UO_3283 (O_3283,N_29854,N_29866);
nor UO_3284 (O_3284,N_29814,N_29993);
xor UO_3285 (O_3285,N_29944,N_29830);
or UO_3286 (O_3286,N_29818,N_29848);
or UO_3287 (O_3287,N_29972,N_29816);
xor UO_3288 (O_3288,N_29834,N_29882);
or UO_3289 (O_3289,N_29956,N_29907);
nand UO_3290 (O_3290,N_29966,N_29817);
xor UO_3291 (O_3291,N_29936,N_29849);
and UO_3292 (O_3292,N_29850,N_29836);
xor UO_3293 (O_3293,N_29869,N_29883);
nor UO_3294 (O_3294,N_29895,N_29857);
and UO_3295 (O_3295,N_29956,N_29949);
and UO_3296 (O_3296,N_29996,N_29989);
nand UO_3297 (O_3297,N_29808,N_29879);
or UO_3298 (O_3298,N_29865,N_29803);
nor UO_3299 (O_3299,N_29985,N_29995);
or UO_3300 (O_3300,N_29980,N_29960);
xor UO_3301 (O_3301,N_29938,N_29972);
and UO_3302 (O_3302,N_29977,N_29852);
nor UO_3303 (O_3303,N_29811,N_29936);
or UO_3304 (O_3304,N_29963,N_29934);
xor UO_3305 (O_3305,N_29857,N_29986);
nand UO_3306 (O_3306,N_29894,N_29929);
xor UO_3307 (O_3307,N_29970,N_29832);
or UO_3308 (O_3308,N_29940,N_29933);
or UO_3309 (O_3309,N_29887,N_29994);
and UO_3310 (O_3310,N_29856,N_29945);
and UO_3311 (O_3311,N_29838,N_29817);
and UO_3312 (O_3312,N_29956,N_29867);
xor UO_3313 (O_3313,N_29976,N_29843);
or UO_3314 (O_3314,N_29886,N_29808);
nand UO_3315 (O_3315,N_29857,N_29901);
xor UO_3316 (O_3316,N_29849,N_29803);
nand UO_3317 (O_3317,N_29972,N_29983);
or UO_3318 (O_3318,N_29968,N_29818);
nand UO_3319 (O_3319,N_29886,N_29936);
nand UO_3320 (O_3320,N_29989,N_29860);
or UO_3321 (O_3321,N_29980,N_29983);
or UO_3322 (O_3322,N_29941,N_29960);
and UO_3323 (O_3323,N_29970,N_29980);
nand UO_3324 (O_3324,N_29955,N_29900);
and UO_3325 (O_3325,N_29949,N_29914);
and UO_3326 (O_3326,N_29916,N_29805);
nor UO_3327 (O_3327,N_29885,N_29880);
nand UO_3328 (O_3328,N_29852,N_29981);
and UO_3329 (O_3329,N_29815,N_29820);
nor UO_3330 (O_3330,N_29866,N_29872);
nand UO_3331 (O_3331,N_29971,N_29807);
or UO_3332 (O_3332,N_29872,N_29979);
nand UO_3333 (O_3333,N_29952,N_29881);
xor UO_3334 (O_3334,N_29871,N_29875);
or UO_3335 (O_3335,N_29942,N_29985);
xor UO_3336 (O_3336,N_29807,N_29878);
xor UO_3337 (O_3337,N_29941,N_29965);
or UO_3338 (O_3338,N_29904,N_29996);
nor UO_3339 (O_3339,N_29952,N_29965);
nand UO_3340 (O_3340,N_29833,N_29970);
nor UO_3341 (O_3341,N_29923,N_29943);
nand UO_3342 (O_3342,N_29981,N_29999);
nor UO_3343 (O_3343,N_29806,N_29889);
or UO_3344 (O_3344,N_29992,N_29962);
or UO_3345 (O_3345,N_29965,N_29831);
nand UO_3346 (O_3346,N_29943,N_29873);
nand UO_3347 (O_3347,N_29851,N_29954);
nor UO_3348 (O_3348,N_29886,N_29864);
xor UO_3349 (O_3349,N_29840,N_29918);
and UO_3350 (O_3350,N_29966,N_29845);
nand UO_3351 (O_3351,N_29886,N_29957);
nor UO_3352 (O_3352,N_29986,N_29847);
and UO_3353 (O_3353,N_29845,N_29922);
xnor UO_3354 (O_3354,N_29976,N_29880);
and UO_3355 (O_3355,N_29900,N_29908);
nor UO_3356 (O_3356,N_29928,N_29821);
xnor UO_3357 (O_3357,N_29954,N_29951);
xnor UO_3358 (O_3358,N_29806,N_29871);
or UO_3359 (O_3359,N_29817,N_29936);
or UO_3360 (O_3360,N_29831,N_29897);
xnor UO_3361 (O_3361,N_29887,N_29917);
and UO_3362 (O_3362,N_29931,N_29918);
or UO_3363 (O_3363,N_29841,N_29816);
and UO_3364 (O_3364,N_29992,N_29806);
xnor UO_3365 (O_3365,N_29895,N_29827);
or UO_3366 (O_3366,N_29882,N_29948);
nand UO_3367 (O_3367,N_29904,N_29956);
nand UO_3368 (O_3368,N_29894,N_29990);
nand UO_3369 (O_3369,N_29809,N_29895);
or UO_3370 (O_3370,N_29987,N_29856);
xnor UO_3371 (O_3371,N_29888,N_29857);
and UO_3372 (O_3372,N_29813,N_29923);
nor UO_3373 (O_3373,N_29887,N_29821);
nor UO_3374 (O_3374,N_29912,N_29959);
nand UO_3375 (O_3375,N_29870,N_29830);
or UO_3376 (O_3376,N_29922,N_29819);
nand UO_3377 (O_3377,N_29887,N_29934);
or UO_3378 (O_3378,N_29904,N_29837);
nor UO_3379 (O_3379,N_29856,N_29980);
and UO_3380 (O_3380,N_29891,N_29966);
or UO_3381 (O_3381,N_29892,N_29866);
or UO_3382 (O_3382,N_29982,N_29830);
and UO_3383 (O_3383,N_29904,N_29806);
nand UO_3384 (O_3384,N_29904,N_29901);
xnor UO_3385 (O_3385,N_29915,N_29942);
and UO_3386 (O_3386,N_29823,N_29908);
nor UO_3387 (O_3387,N_29919,N_29895);
and UO_3388 (O_3388,N_29827,N_29811);
and UO_3389 (O_3389,N_29992,N_29984);
nor UO_3390 (O_3390,N_29845,N_29863);
and UO_3391 (O_3391,N_29871,N_29812);
and UO_3392 (O_3392,N_29807,N_29925);
and UO_3393 (O_3393,N_29935,N_29907);
or UO_3394 (O_3394,N_29927,N_29931);
nor UO_3395 (O_3395,N_29848,N_29874);
nand UO_3396 (O_3396,N_29991,N_29998);
nand UO_3397 (O_3397,N_29889,N_29948);
xor UO_3398 (O_3398,N_29879,N_29870);
or UO_3399 (O_3399,N_29912,N_29962);
nor UO_3400 (O_3400,N_29859,N_29988);
or UO_3401 (O_3401,N_29915,N_29806);
xnor UO_3402 (O_3402,N_29910,N_29807);
xnor UO_3403 (O_3403,N_29972,N_29929);
nor UO_3404 (O_3404,N_29961,N_29976);
nor UO_3405 (O_3405,N_29979,N_29852);
nor UO_3406 (O_3406,N_29826,N_29838);
and UO_3407 (O_3407,N_29904,N_29841);
nor UO_3408 (O_3408,N_29953,N_29911);
xnor UO_3409 (O_3409,N_29888,N_29839);
and UO_3410 (O_3410,N_29842,N_29858);
nand UO_3411 (O_3411,N_29877,N_29977);
xor UO_3412 (O_3412,N_29962,N_29978);
xnor UO_3413 (O_3413,N_29976,N_29930);
xnor UO_3414 (O_3414,N_29935,N_29837);
nand UO_3415 (O_3415,N_29817,N_29871);
or UO_3416 (O_3416,N_29929,N_29964);
nand UO_3417 (O_3417,N_29953,N_29978);
and UO_3418 (O_3418,N_29906,N_29991);
and UO_3419 (O_3419,N_29817,N_29839);
or UO_3420 (O_3420,N_29802,N_29925);
nand UO_3421 (O_3421,N_29929,N_29942);
xor UO_3422 (O_3422,N_29921,N_29922);
or UO_3423 (O_3423,N_29820,N_29873);
nand UO_3424 (O_3424,N_29941,N_29946);
nand UO_3425 (O_3425,N_29866,N_29923);
or UO_3426 (O_3426,N_29970,N_29937);
and UO_3427 (O_3427,N_29864,N_29966);
or UO_3428 (O_3428,N_29995,N_29925);
and UO_3429 (O_3429,N_29835,N_29820);
or UO_3430 (O_3430,N_29842,N_29826);
xor UO_3431 (O_3431,N_29975,N_29978);
xnor UO_3432 (O_3432,N_29934,N_29846);
xor UO_3433 (O_3433,N_29990,N_29819);
xnor UO_3434 (O_3434,N_29931,N_29804);
or UO_3435 (O_3435,N_29884,N_29979);
xnor UO_3436 (O_3436,N_29844,N_29932);
xor UO_3437 (O_3437,N_29848,N_29901);
nand UO_3438 (O_3438,N_29824,N_29941);
xor UO_3439 (O_3439,N_29848,N_29954);
nor UO_3440 (O_3440,N_29966,N_29889);
nand UO_3441 (O_3441,N_29874,N_29885);
xnor UO_3442 (O_3442,N_29955,N_29981);
or UO_3443 (O_3443,N_29878,N_29907);
nor UO_3444 (O_3444,N_29802,N_29842);
nor UO_3445 (O_3445,N_29998,N_29943);
nor UO_3446 (O_3446,N_29892,N_29811);
xor UO_3447 (O_3447,N_29820,N_29949);
and UO_3448 (O_3448,N_29899,N_29817);
and UO_3449 (O_3449,N_29814,N_29893);
nor UO_3450 (O_3450,N_29988,N_29970);
and UO_3451 (O_3451,N_29969,N_29832);
or UO_3452 (O_3452,N_29835,N_29817);
or UO_3453 (O_3453,N_29946,N_29964);
nand UO_3454 (O_3454,N_29998,N_29965);
xnor UO_3455 (O_3455,N_29947,N_29992);
or UO_3456 (O_3456,N_29838,N_29864);
xor UO_3457 (O_3457,N_29960,N_29949);
and UO_3458 (O_3458,N_29866,N_29809);
xnor UO_3459 (O_3459,N_29862,N_29871);
nor UO_3460 (O_3460,N_29854,N_29924);
and UO_3461 (O_3461,N_29889,N_29999);
nand UO_3462 (O_3462,N_29996,N_29826);
xnor UO_3463 (O_3463,N_29827,N_29924);
and UO_3464 (O_3464,N_29885,N_29928);
xnor UO_3465 (O_3465,N_29984,N_29932);
nor UO_3466 (O_3466,N_29902,N_29820);
nor UO_3467 (O_3467,N_29986,N_29908);
nand UO_3468 (O_3468,N_29935,N_29823);
or UO_3469 (O_3469,N_29843,N_29836);
xnor UO_3470 (O_3470,N_29995,N_29964);
and UO_3471 (O_3471,N_29901,N_29805);
nand UO_3472 (O_3472,N_29932,N_29859);
or UO_3473 (O_3473,N_29978,N_29881);
xor UO_3474 (O_3474,N_29847,N_29824);
xor UO_3475 (O_3475,N_29994,N_29800);
nand UO_3476 (O_3476,N_29820,N_29971);
nand UO_3477 (O_3477,N_29935,N_29939);
xnor UO_3478 (O_3478,N_29853,N_29824);
nor UO_3479 (O_3479,N_29887,N_29844);
nor UO_3480 (O_3480,N_29910,N_29825);
xnor UO_3481 (O_3481,N_29904,N_29891);
xnor UO_3482 (O_3482,N_29814,N_29964);
and UO_3483 (O_3483,N_29890,N_29942);
and UO_3484 (O_3484,N_29854,N_29956);
or UO_3485 (O_3485,N_29879,N_29840);
or UO_3486 (O_3486,N_29859,N_29974);
nand UO_3487 (O_3487,N_29968,N_29817);
or UO_3488 (O_3488,N_29904,N_29989);
and UO_3489 (O_3489,N_29822,N_29941);
or UO_3490 (O_3490,N_29994,N_29979);
or UO_3491 (O_3491,N_29924,N_29820);
xor UO_3492 (O_3492,N_29935,N_29850);
or UO_3493 (O_3493,N_29908,N_29863);
nand UO_3494 (O_3494,N_29989,N_29868);
and UO_3495 (O_3495,N_29942,N_29877);
xnor UO_3496 (O_3496,N_29859,N_29821);
xor UO_3497 (O_3497,N_29826,N_29886);
xnor UO_3498 (O_3498,N_29839,N_29863);
or UO_3499 (O_3499,N_29842,N_29831);
endmodule