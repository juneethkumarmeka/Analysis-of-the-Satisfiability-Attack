module basic_750_5000_1000_2_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2525,N_2526,N_2527,N_2529,N_2530,N_2531,N_2532,N_2533,N_2535,N_2536,N_2537,N_2538,N_2539,N_2543,N_2546,N_2548,N_2549,N_2550,N_2552,N_2553,N_2554,N_2555,N_2557,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2573,N_2575,N_2576,N_2577,N_2578,N_2579,N_2581,N_2582,N_2583,N_2584,N_2585,N_2587,N_2588,N_2592,N_2593,N_2594,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2607,N_2608,N_2609,N_2610,N_2611,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2621,N_2623,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2657,N_2658,N_2659,N_2661,N_2662,N_2663,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2680,N_2682,N_2684,N_2685,N_2686,N_2687,N_2688,N_2690,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2716,N_2717,N_2719,N_2720,N_2721,N_2722,N_2723,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2743,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2755,N_2756,N_2758,N_2759,N_2760,N_2762,N_2764,N_2765,N_2766,N_2768,N_2769,N_2771,N_2772,N_2773,N_2776,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2797,N_2798,N_2799,N_2800,N_2801,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2814,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2833,N_2834,N_2835,N_2838,N_2839,N_2840,N_2841,N_2842,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2857,N_2858,N_2859,N_2860,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2879,N_2880,N_2881,N_2883,N_2885,N_2887,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2932,N_2933,N_2934,N_2935,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2946,N_2948,N_2949,N_2950,N_2951,N_2953,N_2955,N_2956,N_2958,N_2959,N_2960,N_2961,N_2962,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2973,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2983,N_2984,N_2985,N_2986,N_2987,N_2991,N_2993,N_2994,N_2995,N_2996,N_2997,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3011,N_3012,N_3013,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3046,N_3048,N_3049,N_3051,N_3052,N_3053,N_3054,N_3055,N_3057,N_3058,N_3059,N_3062,N_3063,N_3064,N_3067,N_3068,N_3069,N_3070,N_3071,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3082,N_3083,N_3084,N_3085,N_3087,N_3089,N_3091,N_3092,N_3093,N_3094,N_3096,N_3097,N_3101,N_3102,N_3103,N_3104,N_3105,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3122,N_3123,N_3124,N_3125,N_3127,N_3128,N_3129,N_3131,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3140,N_3142,N_3143,N_3144,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3176,N_3177,N_3178,N_3179,N_3180,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3189,N_3190,N_3192,N_3193,N_3194,N_3195,N_3196,N_3199,N_3201,N_3202,N_3203,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3223,N_3224,N_3225,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3263,N_3264,N_3265,N_3266,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3280,N_3282,N_3283,N_3284,N_3286,N_3287,N_3289,N_3290,N_3291,N_3292,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3310,N_3312,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3351,N_3352,N_3353,N_3355,N_3357,N_3358,N_3359,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3374,N_3375,N_3376,N_3377,N_3379,N_3381,N_3382,N_3383,N_3384,N_3385,N_3387,N_3388,N_3389,N_3390,N_3393,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3412,N_3413,N_3415,N_3416,N_3417,N_3419,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3433,N_3435,N_3436,N_3437,N_3438,N_3441,N_3442,N_3443,N_3444,N_3445,N_3447,N_3448,N_3449,N_3450,N_3453,N_3454,N_3455,N_3456,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3476,N_3477,N_3478,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3487,N_3488,N_3489,N_3492,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3501,N_3502,N_3504,N_3505,N_3508,N_3510,N_3511,N_3512,N_3513,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3527,N_3528,N_3529,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3540,N_3542,N_3543,N_3545,N_3546,N_3547,N_3548,N_3551,N_3552,N_3553,N_3554,N_3555,N_3557,N_3558,N_3559,N_3561,N_3562,N_3563,N_3564,N_3565,N_3567,N_3568,N_3570,N_3571,N_3573,N_3574,N_3576,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3591,N_3592,N_3594,N_3595,N_3596,N_3597,N_3598,N_3601,N_3602,N_3605,N_3607,N_3608,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3621,N_3622,N_3623,N_3624,N_3625,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3640,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3652,N_3653,N_3654,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3664,N_3668,N_3671,N_3673,N_3674,N_3676,N_3677,N_3678,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3711,N_3712,N_3714,N_3715,N_3717,N_3718,N_3719,N_3720,N_3722,N_3723,N_3725,N_3726,N_3727,N_3730,N_3731,N_3732,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3761,N_3762,N_3764,N_3765,N_3766,N_3767,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3777,N_3778,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3795,N_3796,N_3797,N_3798,N_3800,N_3801,N_3803,N_3804,N_3807,N_3808,N_3810,N_3811,N_3812,N_3813,N_3815,N_3816,N_3817,N_3818,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3838,N_3839,N_3840,N_3842,N_3843,N_3844,N_3845,N_3847,N_3848,N_3849,N_3850,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3884,N_3885,N_3886,N_3887,N_3888,N_3891,N_3892,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3940,N_3941,N_3942,N_3943,N_3944,N_3946,N_3947,N_3950,N_3951,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3962,N_3963,N_3967,N_3968,N_3970,N_3971,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3986,N_3987,N_3988,N_3990,N_3992,N_3993,N_3994,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4009,N_4010,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4022,N_4023,N_4028,N_4029,N_4031,N_4032,N_4033,N_4036,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4049,N_4050,N_4051,N_4052,N_4054,N_4058,N_4059,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4070,N_4072,N_4073,N_4074,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4086,N_4088,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4134,N_4136,N_4137,N_4138,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4159,N_4160,N_4162,N_4163,N_4164,N_4165,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4176,N_4180,N_4181,N_4182,N_4183,N_4185,N_4186,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4197,N_4198,N_4199,N_4201,N_4202,N_4204,N_4205,N_4206,N_4207,N_4208,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4220,N_4221,N_4222,N_4223,N_4225,N_4226,N_4229,N_4230,N_4231,N_4233,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4244,N_4245,N_4246,N_4247,N_4248,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4276,N_4277,N_4278,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4287,N_4288,N_4290,N_4291,N_4292,N_4293,N_4294,N_4297,N_4298,N_4299,N_4301,N_4303,N_4304,N_4305,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4328,N_4329,N_4331,N_4332,N_4334,N_4335,N_4336,N_4337,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4346,N_4347,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4361,N_4362,N_4363,N_4364,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4381,N_4382,N_4383,N_4384,N_4386,N_4387,N_4389,N_4390,N_4392,N_4393,N_4395,N_4396,N_4397,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4413,N_4414,N_4415,N_4416,N_4417,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4431,N_4433,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4449,N_4452,N_4453,N_4454,N_4455,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4465,N_4466,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4480,N_4481,N_4482,N_4484,N_4485,N_4486,N_4487,N_4489,N_4491,N_4493,N_4494,N_4496,N_4497,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4544,N_4546,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4562,N_4563,N_4565,N_4566,N_4567,N_4568,N_4570,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4582,N_4583,N_4585,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4598,N_4599,N_4601,N_4602,N_4603,N_4604,N_4605,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4622,N_4623,N_4624,N_4626,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4636,N_4637,N_4638,N_4639,N_4641,N_4642,N_4643,N_4644,N_4646,N_4648,N_4649,N_4651,N_4655,N_4656,N_4659,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4668,N_4669,N_4670,N_4671,N_4672,N_4674,N_4675,N_4676,N_4677,N_4680,N_4681,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4690,N_4691,N_4693,N_4694,N_4695,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4705,N_4707,N_4709,N_4710,N_4711,N_4713,N_4714,N_4715,N_4717,N_4718,N_4719,N_4720,N_4722,N_4724,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4741,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4753,N_4754,N_4756,N_4757,N_4759,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4769,N_4770,N_4771,N_4772,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4790,N_4791,N_4792,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4811,N_4812,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4825,N_4827,N_4828,N_4829,N_4830,N_4831,N_4833,N_4834,N_4835,N_4836,N_4837,N_4839,N_4840,N_4841,N_4842,N_4844,N_4845,N_4846,N_4849,N_4851,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4869,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4882,N_4884,N_4885,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4903,N_4904,N_4906,N_4908,N_4909,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4932,N_4933,N_4934,N_4935,N_4936,N_4938,N_4941,N_4942,N_4944,N_4945,N_4946,N_4948,N_4950,N_4951,N_4952,N_4954,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4964,N_4965,N_4966,N_4968,N_4969,N_4970,N_4972,N_4973,N_4974,N_4975,N_4978,N_4979,N_4980,N_4982,N_4985,N_4986,N_4987,N_4991,N_4992,N_4993,N_4994,N_4995,N_4997,N_4999;
nor U0 (N_0,In_42,In_480);
xnor U1 (N_1,In_152,In_313);
or U2 (N_2,In_438,In_600);
or U3 (N_3,In_723,In_120);
and U4 (N_4,In_401,In_614);
xor U5 (N_5,In_440,In_726);
nand U6 (N_6,In_674,In_301);
nand U7 (N_7,In_353,In_170);
nand U8 (N_8,In_62,In_681);
nor U9 (N_9,In_113,In_327);
or U10 (N_10,In_141,In_549);
and U11 (N_11,In_660,In_457);
nor U12 (N_12,In_2,In_181);
xor U13 (N_13,In_349,In_148);
and U14 (N_14,In_57,In_0);
or U15 (N_15,In_583,In_559);
nand U16 (N_16,In_630,In_306);
xnor U17 (N_17,In_274,In_482);
xor U18 (N_18,In_531,In_633);
and U19 (N_19,In_203,In_748);
and U20 (N_20,In_355,In_212);
xor U21 (N_21,In_267,In_333);
nand U22 (N_22,In_716,In_540);
nor U23 (N_23,In_618,In_523);
or U24 (N_24,In_613,In_568);
xor U25 (N_25,In_235,In_490);
nand U26 (N_26,In_577,In_462);
nor U27 (N_27,In_185,In_467);
or U28 (N_28,In_142,In_663);
xor U29 (N_29,In_393,In_485);
or U30 (N_30,In_563,In_180);
or U31 (N_31,In_29,In_702);
nand U32 (N_32,In_744,In_690);
and U33 (N_33,In_75,In_6);
xnor U34 (N_34,In_534,In_528);
or U35 (N_35,In_352,In_698);
nand U36 (N_36,In_677,In_10);
or U37 (N_37,In_426,In_383);
xnor U38 (N_38,In_562,In_169);
and U39 (N_39,In_703,In_552);
xor U40 (N_40,In_286,In_470);
and U41 (N_41,In_419,In_557);
nor U42 (N_42,In_146,In_429);
nor U43 (N_43,In_724,In_687);
xnor U44 (N_44,In_163,In_91);
or U45 (N_45,In_332,In_733);
nor U46 (N_46,In_387,In_138);
nor U47 (N_47,In_159,In_592);
nor U48 (N_48,In_239,In_437);
xnor U49 (N_49,In_32,In_292);
nand U50 (N_50,In_705,In_623);
xor U51 (N_51,In_245,In_588);
nand U52 (N_52,In_591,In_231);
or U53 (N_53,In_565,In_463);
and U54 (N_54,In_629,In_136);
nand U55 (N_55,In_68,In_701);
nand U56 (N_56,In_688,In_519);
or U57 (N_57,In_340,In_342);
xnor U58 (N_58,In_520,In_628);
or U59 (N_59,In_213,In_553);
nand U60 (N_60,In_73,In_415);
and U61 (N_61,In_529,In_537);
xor U62 (N_62,In_334,In_337);
and U63 (N_63,In_365,In_211);
nor U64 (N_64,In_28,In_464);
nand U65 (N_65,In_83,In_294);
nor U66 (N_66,In_248,In_555);
or U67 (N_67,In_601,In_648);
and U68 (N_68,In_522,In_36);
or U69 (N_69,In_643,In_476);
xor U70 (N_70,In_339,In_536);
nand U71 (N_71,In_511,In_134);
nor U72 (N_72,In_240,In_499);
nor U73 (N_73,In_725,In_608);
nand U74 (N_74,In_742,In_575);
and U75 (N_75,In_244,In_609);
and U76 (N_76,In_38,In_578);
and U77 (N_77,In_434,In_341);
nand U78 (N_78,In_101,In_111);
or U79 (N_79,In_201,In_18);
nor U80 (N_80,In_281,In_45);
nand U81 (N_81,In_634,In_56);
and U82 (N_82,In_736,In_518);
nor U83 (N_83,In_264,In_139);
or U84 (N_84,In_727,In_597);
nor U85 (N_85,In_638,In_79);
and U86 (N_86,In_713,In_247);
nor U87 (N_87,In_535,In_654);
and U88 (N_88,In_372,In_295);
or U89 (N_89,In_734,In_494);
nor U90 (N_90,In_3,In_607);
nand U91 (N_91,In_197,In_722);
nor U92 (N_92,In_172,In_659);
nand U93 (N_93,In_465,In_740);
xor U94 (N_94,In_406,In_399);
or U95 (N_95,In_53,In_602);
nand U96 (N_96,In_521,In_530);
and U97 (N_97,In_508,In_130);
or U98 (N_98,In_305,In_194);
or U99 (N_99,In_689,In_533);
or U100 (N_100,In_509,In_256);
and U101 (N_101,In_550,In_547);
xor U102 (N_102,In_151,In_362);
nand U103 (N_103,In_7,In_664);
xor U104 (N_104,In_729,In_675);
or U105 (N_105,In_544,In_98);
and U106 (N_106,In_30,In_404);
or U107 (N_107,In_110,In_114);
or U108 (N_108,In_644,In_361);
xor U109 (N_109,In_495,In_593);
nor U110 (N_110,In_243,In_685);
nand U111 (N_111,In_206,In_155);
or U112 (N_112,In_627,In_52);
and U113 (N_113,In_241,In_187);
nor U114 (N_114,In_596,In_599);
nand U115 (N_115,In_266,In_513);
nor U116 (N_116,In_432,In_95);
nor U117 (N_117,In_708,In_587);
nor U118 (N_118,In_610,In_672);
nor U119 (N_119,In_217,In_396);
nor U120 (N_120,In_478,In_283);
and U121 (N_121,In_204,In_491);
xnor U122 (N_122,In_147,In_143);
xor U123 (N_123,In_459,In_431);
xnor U124 (N_124,In_317,In_356);
xnor U125 (N_125,In_706,In_749);
or U126 (N_126,In_299,In_541);
nor U127 (N_127,In_268,In_135);
nand U128 (N_128,In_377,In_254);
xnor U129 (N_129,In_220,In_566);
or U130 (N_130,In_397,In_154);
xor U131 (N_131,In_506,In_741);
xnor U132 (N_132,In_272,In_696);
and U133 (N_133,In_145,In_405);
nand U134 (N_134,In_580,In_473);
nor U135 (N_135,In_493,In_14);
nand U136 (N_136,In_604,In_363);
or U137 (N_137,In_449,In_474);
or U138 (N_138,In_5,In_72);
or U139 (N_139,In_157,In_164);
xnor U140 (N_140,In_394,In_65);
nand U141 (N_141,In_489,In_258);
and U142 (N_142,In_156,In_461);
and U143 (N_143,In_611,In_739);
nand U144 (N_144,In_642,In_226);
and U145 (N_145,In_308,In_284);
xnor U146 (N_146,In_477,In_210);
and U147 (N_147,In_27,In_214);
or U148 (N_148,In_400,In_423);
and U149 (N_149,In_561,In_350);
nand U150 (N_150,In_22,In_17);
and U151 (N_151,In_430,In_124);
xnor U152 (N_152,In_96,In_162);
xor U153 (N_153,In_416,In_285);
or U154 (N_154,In_719,In_78);
xnor U155 (N_155,In_487,In_103);
xnor U156 (N_156,In_469,In_665);
xor U157 (N_157,In_237,In_265);
nor U158 (N_158,In_586,In_109);
xor U159 (N_159,In_46,In_402);
nor U160 (N_160,In_300,In_326);
nand U161 (N_161,In_238,In_390);
xnor U162 (N_162,In_100,In_656);
nor U163 (N_163,In_88,In_571);
nor U164 (N_164,In_173,In_691);
nor U165 (N_165,In_684,In_730);
or U166 (N_166,In_460,In_380);
and U167 (N_167,In_358,In_505);
or U168 (N_168,In_297,In_354);
nor U169 (N_169,In_425,In_525);
or U170 (N_170,In_411,In_617);
xnor U171 (N_171,In_107,In_323);
nand U172 (N_172,In_153,In_526);
or U173 (N_173,In_621,In_71);
and U174 (N_174,In_196,In_165);
nor U175 (N_175,In_376,In_551);
nand U176 (N_176,In_125,In_382);
and U177 (N_177,In_123,In_199);
xor U178 (N_178,In_312,In_598);
and U179 (N_179,In_514,In_347);
or U180 (N_180,In_357,In_200);
or U181 (N_181,In_585,In_589);
nand U182 (N_182,In_167,In_497);
xor U183 (N_183,In_496,In_11);
and U184 (N_184,In_441,In_466);
xor U185 (N_185,In_403,In_82);
nand U186 (N_186,In_502,In_524);
nor U187 (N_187,In_695,In_503);
nand U188 (N_188,In_58,In_676);
xor U189 (N_189,In_360,In_417);
and U190 (N_190,In_90,In_289);
and U191 (N_191,In_126,In_658);
and U192 (N_192,In_686,In_177);
nand U193 (N_193,In_661,In_545);
xnor U194 (N_194,In_261,In_158);
nor U195 (N_195,In_330,In_699);
nor U196 (N_196,In_581,In_373);
nand U197 (N_197,In_407,In_21);
nand U198 (N_198,In_683,In_31);
nor U199 (N_199,In_34,In_15);
and U200 (N_200,In_121,In_398);
or U201 (N_201,In_445,In_37);
and U202 (N_202,In_635,In_50);
nor U203 (N_203,In_242,In_603);
nand U204 (N_204,In_646,In_171);
nand U205 (N_205,In_647,In_279);
xnor U206 (N_206,In_391,In_374);
nor U207 (N_207,In_296,In_472);
xor U208 (N_208,In_262,In_251);
or U209 (N_209,In_651,In_325);
and U210 (N_210,In_447,In_290);
nand U211 (N_211,In_302,In_178);
nand U212 (N_212,In_278,In_558);
nor U213 (N_213,In_632,In_218);
xnor U214 (N_214,In_395,In_202);
nand U215 (N_215,In_694,In_287);
nor U216 (N_216,In_392,In_564);
xnor U217 (N_217,In_378,In_682);
nand U218 (N_218,In_606,In_40);
and U219 (N_219,In_453,In_35);
nor U220 (N_220,In_288,In_700);
nand U221 (N_221,In_626,In_452);
nor U222 (N_222,In_479,In_737);
nand U223 (N_223,In_590,In_260);
and U224 (N_224,In_51,In_208);
or U225 (N_225,In_412,In_150);
nor U226 (N_226,In_731,In_85);
nand U227 (N_227,In_567,In_324);
and U228 (N_228,In_693,In_44);
or U229 (N_229,In_166,In_189);
and U230 (N_230,In_576,In_714);
xnor U231 (N_231,In_657,In_174);
or U232 (N_232,In_668,In_418);
or U233 (N_233,In_222,In_616);
nor U234 (N_234,In_198,In_662);
nor U235 (N_235,In_743,In_223);
nand U236 (N_236,In_542,In_328);
xor U237 (N_237,In_455,In_182);
or U238 (N_238,In_582,In_692);
xnor U239 (N_239,In_560,In_624);
xor U240 (N_240,In_483,In_81);
and U241 (N_241,In_670,In_527);
nor U242 (N_242,In_717,In_129);
nand U243 (N_243,In_93,In_720);
and U244 (N_244,In_570,In_225);
nand U245 (N_245,In_436,In_615);
and U246 (N_246,In_321,In_669);
nor U247 (N_247,In_351,In_252);
nand U248 (N_248,In_512,In_572);
and U249 (N_249,In_246,In_667);
nor U250 (N_250,In_538,In_66);
or U251 (N_251,In_303,In_671);
and U252 (N_252,In_707,In_137);
nor U253 (N_253,In_712,In_546);
or U254 (N_254,In_64,In_515);
and U255 (N_255,In_422,In_112);
or U256 (N_256,In_679,In_276);
xnor U257 (N_257,In_554,In_140);
nand U258 (N_258,In_364,In_548);
nand U259 (N_259,In_205,In_486);
and U260 (N_260,In_270,In_543);
nand U261 (N_261,In_25,In_448);
nor U262 (N_262,In_381,In_257);
and U263 (N_263,In_442,In_273);
nor U264 (N_264,In_424,In_386);
nor U265 (N_265,In_188,In_230);
or U266 (N_266,In_504,In_718);
xnor U267 (N_267,In_507,In_179);
xor U268 (N_268,In_343,In_1);
and U269 (N_269,In_47,In_336);
nand U270 (N_270,In_331,In_620);
xnor U271 (N_271,In_738,In_193);
and U272 (N_272,In_408,In_456);
and U273 (N_273,In_69,In_652);
nand U274 (N_274,In_277,In_4);
and U275 (N_275,In_732,In_655);
and U276 (N_276,In_492,In_366);
xnor U277 (N_277,In_275,In_569);
xor U278 (N_278,In_304,In_99);
xnor U279 (N_279,In_12,In_747);
nand U280 (N_280,In_20,In_293);
xor U281 (N_281,In_344,In_131);
xor U282 (N_282,In_63,In_595);
nand U283 (N_283,In_420,In_318);
xnor U284 (N_284,In_271,In_454);
nand U285 (N_285,In_33,In_116);
xnor U286 (N_286,In_314,In_584);
and U287 (N_287,In_379,In_161);
or U288 (N_288,In_49,In_59);
xor U289 (N_289,In_458,In_269);
nand U290 (N_290,In_428,In_255);
and U291 (N_291,In_122,In_622);
xnor U292 (N_292,In_221,In_128);
or U293 (N_293,In_532,In_574);
and U294 (N_294,In_89,In_329);
nor U295 (N_295,In_335,In_105);
xor U296 (N_296,In_232,In_253);
or U297 (N_297,In_715,In_410);
nand U298 (N_298,In_67,In_371);
xnor U299 (N_299,In_227,In_315);
or U300 (N_300,In_573,In_39);
and U301 (N_301,In_612,In_501);
or U302 (N_302,In_639,In_229);
and U303 (N_303,In_16,In_55);
or U304 (N_304,In_233,In_645);
and U305 (N_305,In_195,In_250);
and U306 (N_306,In_510,In_77);
nor U307 (N_307,In_192,In_637);
nor U308 (N_308,In_435,In_307);
and U309 (N_309,In_369,In_673);
nand U310 (N_310,In_653,In_481);
xnor U311 (N_311,In_444,In_48);
xor U312 (N_312,In_471,In_348);
nand U313 (N_313,In_119,In_413);
nor U314 (N_314,In_191,In_309);
xnor U315 (N_315,In_468,In_54);
nor U316 (N_316,In_500,In_517);
nand U317 (N_317,In_389,In_176);
xor U318 (N_318,In_87,In_280);
nor U319 (N_319,In_94,In_678);
or U320 (N_320,In_384,In_215);
nor U321 (N_321,In_539,In_433);
or U322 (N_322,In_367,In_108);
xor U323 (N_323,In_224,In_168);
and U324 (N_324,In_117,In_282);
xor U325 (N_325,In_704,In_319);
and U326 (N_326,In_84,In_132);
and U327 (N_327,In_641,In_190);
xor U328 (N_328,In_209,In_127);
or U329 (N_329,In_636,In_414);
nand U330 (N_330,In_345,In_666);
nand U331 (N_331,In_443,In_375);
xnor U332 (N_332,In_13,In_298);
nand U333 (N_333,In_144,In_236);
xor U334 (N_334,In_219,In_579);
nand U335 (N_335,In_625,In_97);
nor U336 (N_336,In_338,In_409);
or U337 (N_337,In_234,In_8);
nor U338 (N_338,In_475,In_76);
xnor U339 (N_339,In_186,In_207);
or U340 (N_340,In_649,In_70);
nor U341 (N_341,In_594,In_484);
and U342 (N_342,In_359,In_184);
nor U343 (N_343,In_322,In_439);
xnor U344 (N_344,In_263,In_709);
nor U345 (N_345,In_216,In_745);
xor U346 (N_346,In_19,In_118);
or U347 (N_347,In_311,In_446);
xnor U348 (N_348,In_385,In_106);
and U349 (N_349,In_249,In_516);
nor U350 (N_350,In_697,In_735);
or U351 (N_351,In_228,In_498);
or U352 (N_352,In_388,In_43);
xor U353 (N_353,In_102,In_721);
and U354 (N_354,In_316,In_26);
and U355 (N_355,In_23,In_133);
and U356 (N_356,In_619,In_728);
nor U357 (N_357,In_291,In_259);
or U358 (N_358,In_149,In_160);
or U359 (N_359,In_451,In_746);
xnor U360 (N_360,In_640,In_370);
and U361 (N_361,In_74,In_605);
nor U362 (N_362,In_368,In_556);
nand U363 (N_363,In_60,In_183);
xnor U364 (N_364,In_488,In_346);
nor U365 (N_365,In_92,In_680);
nor U366 (N_366,In_175,In_427);
nor U367 (N_367,In_115,In_320);
xnor U368 (N_368,In_650,In_310);
nor U369 (N_369,In_631,In_711);
nand U370 (N_370,In_710,In_450);
nor U371 (N_371,In_86,In_24);
or U372 (N_372,In_421,In_104);
nor U373 (N_373,In_41,In_9);
and U374 (N_374,In_61,In_80);
or U375 (N_375,In_4,In_234);
nor U376 (N_376,In_487,In_671);
nor U377 (N_377,In_267,In_51);
or U378 (N_378,In_76,In_146);
xor U379 (N_379,In_643,In_114);
xor U380 (N_380,In_16,In_488);
nand U381 (N_381,In_709,In_312);
xnor U382 (N_382,In_533,In_187);
nor U383 (N_383,In_680,In_415);
and U384 (N_384,In_636,In_411);
nand U385 (N_385,In_220,In_476);
and U386 (N_386,In_213,In_483);
nor U387 (N_387,In_102,In_625);
nor U388 (N_388,In_53,In_548);
and U389 (N_389,In_150,In_708);
nand U390 (N_390,In_26,In_648);
or U391 (N_391,In_748,In_136);
or U392 (N_392,In_419,In_556);
or U393 (N_393,In_253,In_200);
nor U394 (N_394,In_76,In_222);
or U395 (N_395,In_320,In_248);
xor U396 (N_396,In_536,In_652);
nor U397 (N_397,In_567,In_743);
xnor U398 (N_398,In_167,In_496);
xnor U399 (N_399,In_246,In_50);
xnor U400 (N_400,In_706,In_722);
nor U401 (N_401,In_153,In_126);
xor U402 (N_402,In_667,In_360);
or U403 (N_403,In_445,In_666);
and U404 (N_404,In_732,In_422);
and U405 (N_405,In_389,In_419);
or U406 (N_406,In_565,In_549);
nor U407 (N_407,In_157,In_148);
nand U408 (N_408,In_570,In_401);
nor U409 (N_409,In_338,In_453);
and U410 (N_410,In_685,In_710);
and U411 (N_411,In_89,In_638);
nand U412 (N_412,In_494,In_501);
nor U413 (N_413,In_285,In_733);
or U414 (N_414,In_736,In_372);
xor U415 (N_415,In_590,In_482);
nor U416 (N_416,In_403,In_391);
nand U417 (N_417,In_655,In_148);
xor U418 (N_418,In_511,In_527);
or U419 (N_419,In_292,In_478);
xnor U420 (N_420,In_568,In_57);
xnor U421 (N_421,In_251,In_314);
nand U422 (N_422,In_581,In_3);
nor U423 (N_423,In_451,In_409);
xor U424 (N_424,In_619,In_656);
nand U425 (N_425,In_270,In_69);
or U426 (N_426,In_674,In_589);
nand U427 (N_427,In_553,In_62);
nor U428 (N_428,In_113,In_348);
or U429 (N_429,In_657,In_199);
nand U430 (N_430,In_475,In_211);
nor U431 (N_431,In_676,In_212);
nor U432 (N_432,In_686,In_62);
or U433 (N_433,In_203,In_43);
or U434 (N_434,In_690,In_356);
or U435 (N_435,In_746,In_502);
nand U436 (N_436,In_407,In_233);
and U437 (N_437,In_521,In_169);
nand U438 (N_438,In_748,In_363);
and U439 (N_439,In_151,In_491);
nand U440 (N_440,In_721,In_613);
and U441 (N_441,In_418,In_301);
nand U442 (N_442,In_553,In_459);
or U443 (N_443,In_434,In_648);
and U444 (N_444,In_399,In_552);
or U445 (N_445,In_629,In_308);
or U446 (N_446,In_57,In_623);
nand U447 (N_447,In_214,In_699);
nor U448 (N_448,In_353,In_731);
nor U449 (N_449,In_409,In_233);
xor U450 (N_450,In_343,In_139);
nand U451 (N_451,In_578,In_633);
or U452 (N_452,In_247,In_8);
nand U453 (N_453,In_670,In_222);
or U454 (N_454,In_247,In_424);
nor U455 (N_455,In_704,In_176);
nand U456 (N_456,In_602,In_4);
or U457 (N_457,In_330,In_439);
xnor U458 (N_458,In_28,In_719);
or U459 (N_459,In_170,In_146);
nand U460 (N_460,In_327,In_16);
xnor U461 (N_461,In_54,In_138);
nor U462 (N_462,In_473,In_588);
nor U463 (N_463,In_303,In_75);
nand U464 (N_464,In_745,In_532);
and U465 (N_465,In_449,In_255);
and U466 (N_466,In_93,In_165);
or U467 (N_467,In_446,In_455);
nand U468 (N_468,In_331,In_336);
xnor U469 (N_469,In_557,In_442);
or U470 (N_470,In_277,In_667);
nor U471 (N_471,In_450,In_22);
nor U472 (N_472,In_709,In_512);
nor U473 (N_473,In_742,In_543);
or U474 (N_474,In_478,In_339);
nor U475 (N_475,In_693,In_577);
or U476 (N_476,In_618,In_608);
nand U477 (N_477,In_364,In_300);
and U478 (N_478,In_286,In_631);
xnor U479 (N_479,In_22,In_381);
nor U480 (N_480,In_496,In_140);
and U481 (N_481,In_666,In_576);
or U482 (N_482,In_410,In_215);
or U483 (N_483,In_641,In_742);
or U484 (N_484,In_496,In_158);
nor U485 (N_485,In_408,In_186);
nor U486 (N_486,In_558,In_549);
or U487 (N_487,In_27,In_695);
xor U488 (N_488,In_288,In_725);
nand U489 (N_489,In_548,In_1);
xnor U490 (N_490,In_514,In_120);
xor U491 (N_491,In_319,In_78);
and U492 (N_492,In_160,In_363);
nand U493 (N_493,In_14,In_198);
nand U494 (N_494,In_342,In_111);
nand U495 (N_495,In_709,In_631);
nand U496 (N_496,In_180,In_300);
nand U497 (N_497,In_242,In_47);
nor U498 (N_498,In_403,In_396);
nor U499 (N_499,In_211,In_314);
nand U500 (N_500,In_419,In_471);
nand U501 (N_501,In_379,In_594);
or U502 (N_502,In_148,In_16);
xor U503 (N_503,In_37,In_263);
or U504 (N_504,In_302,In_366);
nor U505 (N_505,In_178,In_229);
nor U506 (N_506,In_220,In_541);
or U507 (N_507,In_129,In_372);
nand U508 (N_508,In_431,In_386);
nor U509 (N_509,In_142,In_168);
and U510 (N_510,In_147,In_258);
nor U511 (N_511,In_592,In_200);
nor U512 (N_512,In_40,In_720);
or U513 (N_513,In_453,In_358);
and U514 (N_514,In_705,In_203);
nor U515 (N_515,In_243,In_161);
or U516 (N_516,In_700,In_734);
nor U517 (N_517,In_130,In_78);
or U518 (N_518,In_205,In_227);
or U519 (N_519,In_410,In_335);
nor U520 (N_520,In_711,In_650);
and U521 (N_521,In_159,In_57);
xnor U522 (N_522,In_729,In_406);
xnor U523 (N_523,In_739,In_358);
xnor U524 (N_524,In_236,In_495);
or U525 (N_525,In_102,In_500);
nor U526 (N_526,In_474,In_360);
xnor U527 (N_527,In_470,In_278);
nor U528 (N_528,In_552,In_14);
nor U529 (N_529,In_347,In_206);
nand U530 (N_530,In_126,In_221);
and U531 (N_531,In_322,In_280);
or U532 (N_532,In_29,In_716);
and U533 (N_533,In_167,In_532);
nand U534 (N_534,In_677,In_482);
xnor U535 (N_535,In_696,In_157);
and U536 (N_536,In_85,In_177);
and U537 (N_537,In_453,In_346);
nand U538 (N_538,In_218,In_124);
nand U539 (N_539,In_175,In_729);
xnor U540 (N_540,In_454,In_124);
and U541 (N_541,In_654,In_691);
xnor U542 (N_542,In_203,In_181);
xnor U543 (N_543,In_404,In_528);
and U544 (N_544,In_544,In_707);
nand U545 (N_545,In_7,In_647);
and U546 (N_546,In_584,In_284);
nand U547 (N_547,In_296,In_364);
or U548 (N_548,In_4,In_135);
or U549 (N_549,In_614,In_304);
nand U550 (N_550,In_219,In_437);
or U551 (N_551,In_329,In_323);
or U552 (N_552,In_36,In_278);
or U553 (N_553,In_285,In_275);
nand U554 (N_554,In_117,In_52);
nor U555 (N_555,In_513,In_480);
xor U556 (N_556,In_54,In_273);
xor U557 (N_557,In_401,In_181);
xnor U558 (N_558,In_621,In_241);
or U559 (N_559,In_454,In_205);
xnor U560 (N_560,In_261,In_162);
or U561 (N_561,In_629,In_497);
nand U562 (N_562,In_542,In_325);
and U563 (N_563,In_469,In_133);
or U564 (N_564,In_87,In_220);
and U565 (N_565,In_355,In_353);
xor U566 (N_566,In_615,In_384);
or U567 (N_567,In_597,In_415);
and U568 (N_568,In_520,In_416);
and U569 (N_569,In_688,In_547);
nand U570 (N_570,In_210,In_729);
or U571 (N_571,In_673,In_449);
and U572 (N_572,In_173,In_229);
xor U573 (N_573,In_702,In_430);
or U574 (N_574,In_658,In_329);
and U575 (N_575,In_95,In_695);
xnor U576 (N_576,In_611,In_186);
nand U577 (N_577,In_535,In_447);
and U578 (N_578,In_159,In_445);
or U579 (N_579,In_257,In_587);
nand U580 (N_580,In_263,In_674);
nor U581 (N_581,In_730,In_495);
nand U582 (N_582,In_9,In_51);
nor U583 (N_583,In_183,In_349);
xor U584 (N_584,In_145,In_712);
or U585 (N_585,In_148,In_645);
xnor U586 (N_586,In_666,In_658);
nand U587 (N_587,In_392,In_409);
or U588 (N_588,In_481,In_129);
nor U589 (N_589,In_157,In_521);
nor U590 (N_590,In_163,In_343);
or U591 (N_591,In_497,In_663);
xnor U592 (N_592,In_330,In_724);
or U593 (N_593,In_244,In_434);
nor U594 (N_594,In_605,In_273);
nor U595 (N_595,In_623,In_452);
xor U596 (N_596,In_638,In_685);
or U597 (N_597,In_143,In_582);
xor U598 (N_598,In_177,In_117);
nand U599 (N_599,In_628,In_650);
or U600 (N_600,In_727,In_368);
nand U601 (N_601,In_141,In_381);
xor U602 (N_602,In_501,In_445);
or U603 (N_603,In_15,In_172);
nand U604 (N_604,In_719,In_680);
xor U605 (N_605,In_579,In_451);
xor U606 (N_606,In_407,In_370);
and U607 (N_607,In_2,In_635);
or U608 (N_608,In_651,In_567);
and U609 (N_609,In_205,In_54);
and U610 (N_610,In_70,In_305);
nand U611 (N_611,In_353,In_331);
and U612 (N_612,In_306,In_505);
and U613 (N_613,In_738,In_495);
or U614 (N_614,In_276,In_175);
or U615 (N_615,In_578,In_113);
nand U616 (N_616,In_581,In_186);
and U617 (N_617,In_483,In_655);
nor U618 (N_618,In_327,In_157);
and U619 (N_619,In_435,In_686);
or U620 (N_620,In_366,In_488);
or U621 (N_621,In_572,In_344);
nand U622 (N_622,In_636,In_476);
nand U623 (N_623,In_121,In_254);
nor U624 (N_624,In_638,In_368);
and U625 (N_625,In_358,In_161);
and U626 (N_626,In_155,In_662);
or U627 (N_627,In_288,In_529);
and U628 (N_628,In_169,In_82);
nand U629 (N_629,In_192,In_266);
nand U630 (N_630,In_102,In_679);
nor U631 (N_631,In_551,In_351);
and U632 (N_632,In_173,In_385);
xnor U633 (N_633,In_105,In_34);
nand U634 (N_634,In_148,In_570);
or U635 (N_635,In_733,In_411);
nor U636 (N_636,In_317,In_496);
and U637 (N_637,In_444,In_659);
xnor U638 (N_638,In_724,In_615);
nand U639 (N_639,In_377,In_356);
nor U640 (N_640,In_48,In_668);
nand U641 (N_641,In_591,In_71);
and U642 (N_642,In_63,In_54);
nand U643 (N_643,In_45,In_460);
and U644 (N_644,In_574,In_420);
nand U645 (N_645,In_94,In_232);
nand U646 (N_646,In_405,In_53);
nor U647 (N_647,In_201,In_647);
and U648 (N_648,In_403,In_277);
xor U649 (N_649,In_489,In_123);
nor U650 (N_650,In_153,In_586);
nand U651 (N_651,In_424,In_267);
nand U652 (N_652,In_686,In_396);
nor U653 (N_653,In_677,In_537);
or U654 (N_654,In_651,In_523);
nor U655 (N_655,In_124,In_120);
and U656 (N_656,In_655,In_658);
xnor U657 (N_657,In_96,In_435);
or U658 (N_658,In_705,In_541);
xnor U659 (N_659,In_723,In_171);
xor U660 (N_660,In_106,In_165);
xor U661 (N_661,In_591,In_431);
xnor U662 (N_662,In_471,In_106);
and U663 (N_663,In_74,In_367);
nor U664 (N_664,In_86,In_617);
or U665 (N_665,In_491,In_217);
and U666 (N_666,In_146,In_532);
nor U667 (N_667,In_10,In_531);
xor U668 (N_668,In_612,In_178);
nor U669 (N_669,In_584,In_259);
nand U670 (N_670,In_603,In_158);
nor U671 (N_671,In_501,In_687);
or U672 (N_672,In_174,In_627);
or U673 (N_673,In_288,In_48);
nand U674 (N_674,In_534,In_631);
and U675 (N_675,In_475,In_600);
and U676 (N_676,In_306,In_573);
nor U677 (N_677,In_15,In_666);
or U678 (N_678,In_63,In_25);
and U679 (N_679,In_554,In_696);
xnor U680 (N_680,In_544,In_337);
or U681 (N_681,In_11,In_251);
xnor U682 (N_682,In_724,In_134);
nand U683 (N_683,In_701,In_170);
or U684 (N_684,In_704,In_244);
nor U685 (N_685,In_612,In_115);
nand U686 (N_686,In_411,In_581);
xor U687 (N_687,In_191,In_390);
and U688 (N_688,In_552,In_596);
or U689 (N_689,In_100,In_319);
and U690 (N_690,In_258,In_45);
xor U691 (N_691,In_184,In_132);
xnor U692 (N_692,In_24,In_670);
or U693 (N_693,In_474,In_245);
xor U694 (N_694,In_651,In_228);
nand U695 (N_695,In_33,In_163);
nor U696 (N_696,In_669,In_635);
xnor U697 (N_697,In_43,In_696);
and U698 (N_698,In_355,In_737);
and U699 (N_699,In_482,In_582);
xnor U700 (N_700,In_419,In_627);
xnor U701 (N_701,In_116,In_437);
xnor U702 (N_702,In_338,In_23);
nand U703 (N_703,In_735,In_369);
xor U704 (N_704,In_255,In_55);
xor U705 (N_705,In_709,In_417);
or U706 (N_706,In_353,In_736);
xor U707 (N_707,In_418,In_288);
nand U708 (N_708,In_521,In_599);
nand U709 (N_709,In_428,In_37);
nor U710 (N_710,In_17,In_733);
xor U711 (N_711,In_50,In_476);
nand U712 (N_712,In_207,In_251);
nor U713 (N_713,In_524,In_217);
or U714 (N_714,In_370,In_591);
nor U715 (N_715,In_155,In_240);
or U716 (N_716,In_298,In_136);
or U717 (N_717,In_28,In_394);
nor U718 (N_718,In_477,In_87);
or U719 (N_719,In_689,In_48);
nor U720 (N_720,In_646,In_405);
and U721 (N_721,In_224,In_606);
or U722 (N_722,In_164,In_371);
nand U723 (N_723,In_58,In_126);
nand U724 (N_724,In_377,In_283);
nand U725 (N_725,In_268,In_159);
nand U726 (N_726,In_469,In_683);
nand U727 (N_727,In_88,In_202);
nor U728 (N_728,In_507,In_747);
xnor U729 (N_729,In_568,In_136);
xnor U730 (N_730,In_331,In_51);
xor U731 (N_731,In_665,In_573);
or U732 (N_732,In_279,In_560);
and U733 (N_733,In_587,In_165);
or U734 (N_734,In_35,In_415);
xnor U735 (N_735,In_503,In_227);
and U736 (N_736,In_259,In_585);
xnor U737 (N_737,In_246,In_141);
nor U738 (N_738,In_46,In_564);
nor U739 (N_739,In_468,In_295);
or U740 (N_740,In_358,In_747);
or U741 (N_741,In_120,In_193);
nand U742 (N_742,In_368,In_453);
xnor U743 (N_743,In_459,In_6);
xor U744 (N_744,In_235,In_533);
xor U745 (N_745,In_607,In_344);
nor U746 (N_746,In_80,In_444);
xor U747 (N_747,In_16,In_22);
xnor U748 (N_748,In_573,In_710);
nor U749 (N_749,In_122,In_247);
xnor U750 (N_750,In_583,In_353);
or U751 (N_751,In_276,In_702);
nand U752 (N_752,In_164,In_703);
nand U753 (N_753,In_591,In_178);
xor U754 (N_754,In_258,In_386);
or U755 (N_755,In_127,In_467);
and U756 (N_756,In_350,In_590);
xor U757 (N_757,In_406,In_618);
and U758 (N_758,In_45,In_659);
nor U759 (N_759,In_86,In_348);
nand U760 (N_760,In_12,In_444);
nand U761 (N_761,In_592,In_144);
nand U762 (N_762,In_554,In_524);
and U763 (N_763,In_157,In_40);
xor U764 (N_764,In_539,In_575);
nor U765 (N_765,In_717,In_684);
xor U766 (N_766,In_746,In_232);
and U767 (N_767,In_289,In_67);
nand U768 (N_768,In_376,In_116);
nand U769 (N_769,In_69,In_153);
nand U770 (N_770,In_585,In_202);
and U771 (N_771,In_660,In_62);
or U772 (N_772,In_160,In_247);
and U773 (N_773,In_44,In_561);
nand U774 (N_774,In_32,In_453);
nor U775 (N_775,In_734,In_462);
xor U776 (N_776,In_594,In_269);
and U777 (N_777,In_316,In_114);
nand U778 (N_778,In_484,In_95);
xnor U779 (N_779,In_530,In_568);
nor U780 (N_780,In_278,In_203);
or U781 (N_781,In_223,In_173);
nor U782 (N_782,In_570,In_447);
and U783 (N_783,In_278,In_427);
nor U784 (N_784,In_676,In_378);
nand U785 (N_785,In_39,In_53);
and U786 (N_786,In_357,In_358);
nand U787 (N_787,In_682,In_118);
and U788 (N_788,In_434,In_665);
or U789 (N_789,In_530,In_655);
nand U790 (N_790,In_61,In_21);
and U791 (N_791,In_363,In_92);
or U792 (N_792,In_21,In_129);
nand U793 (N_793,In_284,In_380);
xor U794 (N_794,In_122,In_72);
nor U795 (N_795,In_201,In_163);
and U796 (N_796,In_417,In_537);
and U797 (N_797,In_327,In_613);
xor U798 (N_798,In_200,In_490);
xor U799 (N_799,In_457,In_478);
or U800 (N_800,In_670,In_387);
or U801 (N_801,In_683,In_325);
xor U802 (N_802,In_542,In_235);
and U803 (N_803,In_653,In_490);
xor U804 (N_804,In_358,In_403);
nand U805 (N_805,In_564,In_346);
nand U806 (N_806,In_380,In_661);
or U807 (N_807,In_288,In_108);
xnor U808 (N_808,In_268,In_137);
nor U809 (N_809,In_226,In_316);
xor U810 (N_810,In_541,In_368);
or U811 (N_811,In_574,In_237);
nor U812 (N_812,In_714,In_498);
nor U813 (N_813,In_393,In_209);
and U814 (N_814,In_493,In_259);
or U815 (N_815,In_149,In_222);
and U816 (N_816,In_247,In_392);
and U817 (N_817,In_608,In_656);
or U818 (N_818,In_442,In_427);
or U819 (N_819,In_386,In_213);
and U820 (N_820,In_211,In_182);
nor U821 (N_821,In_85,In_147);
or U822 (N_822,In_652,In_27);
nor U823 (N_823,In_390,In_184);
or U824 (N_824,In_476,In_380);
nor U825 (N_825,In_156,In_691);
xor U826 (N_826,In_131,In_46);
nand U827 (N_827,In_559,In_704);
and U828 (N_828,In_339,In_198);
nor U829 (N_829,In_173,In_180);
xnor U830 (N_830,In_740,In_733);
nand U831 (N_831,In_660,In_343);
nor U832 (N_832,In_456,In_252);
or U833 (N_833,In_363,In_703);
nand U834 (N_834,In_418,In_227);
or U835 (N_835,In_675,In_471);
nand U836 (N_836,In_479,In_222);
or U837 (N_837,In_513,In_97);
or U838 (N_838,In_44,In_349);
nor U839 (N_839,In_86,In_508);
or U840 (N_840,In_638,In_302);
nand U841 (N_841,In_293,In_283);
nor U842 (N_842,In_511,In_51);
or U843 (N_843,In_686,In_72);
or U844 (N_844,In_343,In_378);
nor U845 (N_845,In_46,In_729);
nor U846 (N_846,In_279,In_355);
or U847 (N_847,In_266,In_718);
xor U848 (N_848,In_532,In_519);
nand U849 (N_849,In_343,In_636);
nor U850 (N_850,In_485,In_375);
and U851 (N_851,In_171,In_713);
xnor U852 (N_852,In_701,In_132);
or U853 (N_853,In_108,In_120);
xor U854 (N_854,In_571,In_90);
nand U855 (N_855,In_469,In_588);
nand U856 (N_856,In_352,In_119);
and U857 (N_857,In_237,In_534);
and U858 (N_858,In_257,In_749);
and U859 (N_859,In_219,In_134);
or U860 (N_860,In_549,In_689);
xor U861 (N_861,In_539,In_149);
xor U862 (N_862,In_693,In_272);
nand U863 (N_863,In_269,In_325);
nor U864 (N_864,In_634,In_292);
nand U865 (N_865,In_692,In_564);
nand U866 (N_866,In_237,In_32);
nand U867 (N_867,In_629,In_628);
and U868 (N_868,In_196,In_395);
nor U869 (N_869,In_147,In_430);
and U870 (N_870,In_410,In_285);
xnor U871 (N_871,In_517,In_705);
nand U872 (N_872,In_428,In_181);
or U873 (N_873,In_79,In_657);
xor U874 (N_874,In_572,In_402);
or U875 (N_875,In_144,In_588);
xor U876 (N_876,In_624,In_457);
nand U877 (N_877,In_301,In_320);
nand U878 (N_878,In_466,In_511);
or U879 (N_879,In_14,In_708);
and U880 (N_880,In_523,In_652);
and U881 (N_881,In_646,In_187);
xnor U882 (N_882,In_582,In_391);
xnor U883 (N_883,In_100,In_650);
nor U884 (N_884,In_277,In_742);
xnor U885 (N_885,In_437,In_392);
and U886 (N_886,In_276,In_409);
or U887 (N_887,In_593,In_746);
nand U888 (N_888,In_93,In_342);
nor U889 (N_889,In_474,In_0);
and U890 (N_890,In_745,In_680);
nand U891 (N_891,In_717,In_476);
or U892 (N_892,In_134,In_741);
nor U893 (N_893,In_721,In_163);
xnor U894 (N_894,In_119,In_186);
nand U895 (N_895,In_612,In_470);
nand U896 (N_896,In_522,In_625);
nor U897 (N_897,In_729,In_89);
or U898 (N_898,In_432,In_296);
nand U899 (N_899,In_210,In_438);
xor U900 (N_900,In_176,In_277);
or U901 (N_901,In_198,In_122);
or U902 (N_902,In_236,In_299);
nand U903 (N_903,In_3,In_450);
nor U904 (N_904,In_698,In_651);
nor U905 (N_905,In_357,In_58);
or U906 (N_906,In_435,In_370);
and U907 (N_907,In_367,In_68);
or U908 (N_908,In_673,In_439);
nor U909 (N_909,In_430,In_362);
nand U910 (N_910,In_249,In_39);
nor U911 (N_911,In_153,In_556);
or U912 (N_912,In_180,In_316);
nor U913 (N_913,In_69,In_289);
nor U914 (N_914,In_561,In_4);
or U915 (N_915,In_276,In_123);
or U916 (N_916,In_443,In_157);
and U917 (N_917,In_421,In_619);
or U918 (N_918,In_60,In_634);
and U919 (N_919,In_153,In_544);
xnor U920 (N_920,In_701,In_244);
and U921 (N_921,In_230,In_681);
nor U922 (N_922,In_170,In_174);
nand U923 (N_923,In_279,In_331);
nand U924 (N_924,In_647,In_116);
nor U925 (N_925,In_656,In_476);
and U926 (N_926,In_323,In_270);
nand U927 (N_927,In_262,In_358);
nor U928 (N_928,In_163,In_579);
nor U929 (N_929,In_725,In_263);
and U930 (N_930,In_176,In_450);
nand U931 (N_931,In_165,In_673);
or U932 (N_932,In_285,In_394);
or U933 (N_933,In_743,In_476);
and U934 (N_934,In_687,In_281);
nand U935 (N_935,In_350,In_228);
nor U936 (N_936,In_372,In_601);
xor U937 (N_937,In_282,In_68);
or U938 (N_938,In_557,In_696);
or U939 (N_939,In_647,In_543);
or U940 (N_940,In_267,In_164);
and U941 (N_941,In_199,In_224);
xor U942 (N_942,In_250,In_351);
and U943 (N_943,In_101,In_236);
nand U944 (N_944,In_276,In_461);
and U945 (N_945,In_625,In_439);
nand U946 (N_946,In_381,In_286);
xor U947 (N_947,In_268,In_476);
nor U948 (N_948,In_382,In_664);
and U949 (N_949,In_683,In_673);
nand U950 (N_950,In_34,In_299);
xnor U951 (N_951,In_207,In_453);
nand U952 (N_952,In_100,In_133);
and U953 (N_953,In_185,In_678);
nand U954 (N_954,In_273,In_245);
xor U955 (N_955,In_455,In_368);
nand U956 (N_956,In_359,In_126);
xor U957 (N_957,In_677,In_93);
or U958 (N_958,In_484,In_563);
or U959 (N_959,In_62,In_113);
nor U960 (N_960,In_34,In_438);
nor U961 (N_961,In_139,In_427);
or U962 (N_962,In_369,In_3);
nand U963 (N_963,In_213,In_2);
and U964 (N_964,In_75,In_397);
xor U965 (N_965,In_494,In_441);
nand U966 (N_966,In_309,In_591);
nor U967 (N_967,In_265,In_572);
nand U968 (N_968,In_632,In_702);
xnor U969 (N_969,In_457,In_22);
xor U970 (N_970,In_230,In_316);
nand U971 (N_971,In_185,In_230);
or U972 (N_972,In_381,In_432);
or U973 (N_973,In_440,In_743);
nand U974 (N_974,In_395,In_140);
nand U975 (N_975,In_479,In_469);
nand U976 (N_976,In_568,In_663);
or U977 (N_977,In_416,In_523);
nand U978 (N_978,In_219,In_497);
or U979 (N_979,In_601,In_2);
nor U980 (N_980,In_742,In_398);
or U981 (N_981,In_91,In_679);
and U982 (N_982,In_340,In_101);
or U983 (N_983,In_23,In_185);
nand U984 (N_984,In_55,In_480);
xnor U985 (N_985,In_634,In_748);
or U986 (N_986,In_285,In_452);
and U987 (N_987,In_305,In_515);
or U988 (N_988,In_599,In_283);
and U989 (N_989,In_367,In_350);
xor U990 (N_990,In_471,In_550);
nand U991 (N_991,In_3,In_599);
and U992 (N_992,In_342,In_675);
nor U993 (N_993,In_361,In_412);
or U994 (N_994,In_31,In_482);
and U995 (N_995,In_11,In_430);
nor U996 (N_996,In_40,In_148);
or U997 (N_997,In_109,In_101);
nand U998 (N_998,In_407,In_454);
xnor U999 (N_999,In_197,In_274);
and U1000 (N_1000,In_414,In_38);
and U1001 (N_1001,In_498,In_53);
xnor U1002 (N_1002,In_40,In_272);
and U1003 (N_1003,In_394,In_345);
or U1004 (N_1004,In_577,In_661);
xnor U1005 (N_1005,In_231,In_407);
nor U1006 (N_1006,In_438,In_271);
and U1007 (N_1007,In_412,In_473);
nand U1008 (N_1008,In_432,In_703);
and U1009 (N_1009,In_713,In_748);
and U1010 (N_1010,In_444,In_183);
xnor U1011 (N_1011,In_617,In_649);
nand U1012 (N_1012,In_719,In_357);
xor U1013 (N_1013,In_434,In_110);
and U1014 (N_1014,In_539,In_700);
or U1015 (N_1015,In_744,In_730);
nor U1016 (N_1016,In_2,In_595);
or U1017 (N_1017,In_424,In_622);
nor U1018 (N_1018,In_523,In_660);
xnor U1019 (N_1019,In_515,In_711);
xor U1020 (N_1020,In_736,In_430);
xor U1021 (N_1021,In_13,In_620);
nand U1022 (N_1022,In_381,In_546);
and U1023 (N_1023,In_77,In_342);
or U1024 (N_1024,In_536,In_14);
or U1025 (N_1025,In_646,In_616);
xor U1026 (N_1026,In_584,In_722);
nor U1027 (N_1027,In_373,In_657);
or U1028 (N_1028,In_167,In_465);
or U1029 (N_1029,In_676,In_338);
and U1030 (N_1030,In_373,In_122);
nor U1031 (N_1031,In_227,In_318);
nor U1032 (N_1032,In_258,In_92);
or U1033 (N_1033,In_590,In_721);
or U1034 (N_1034,In_331,In_147);
or U1035 (N_1035,In_505,In_523);
nor U1036 (N_1036,In_451,In_713);
nor U1037 (N_1037,In_584,In_206);
xor U1038 (N_1038,In_618,In_83);
or U1039 (N_1039,In_495,In_484);
or U1040 (N_1040,In_39,In_602);
or U1041 (N_1041,In_481,In_417);
and U1042 (N_1042,In_474,In_627);
or U1043 (N_1043,In_146,In_424);
or U1044 (N_1044,In_151,In_264);
and U1045 (N_1045,In_634,In_378);
nand U1046 (N_1046,In_521,In_129);
or U1047 (N_1047,In_157,In_352);
nor U1048 (N_1048,In_68,In_678);
nor U1049 (N_1049,In_272,In_261);
and U1050 (N_1050,In_231,In_382);
xnor U1051 (N_1051,In_114,In_297);
nand U1052 (N_1052,In_712,In_487);
and U1053 (N_1053,In_166,In_568);
and U1054 (N_1054,In_736,In_251);
nand U1055 (N_1055,In_490,In_308);
nor U1056 (N_1056,In_552,In_641);
and U1057 (N_1057,In_246,In_160);
xnor U1058 (N_1058,In_595,In_95);
nor U1059 (N_1059,In_316,In_697);
or U1060 (N_1060,In_404,In_11);
xnor U1061 (N_1061,In_665,In_44);
xnor U1062 (N_1062,In_460,In_181);
nand U1063 (N_1063,In_282,In_305);
nand U1064 (N_1064,In_385,In_577);
or U1065 (N_1065,In_487,In_321);
and U1066 (N_1066,In_587,In_39);
xnor U1067 (N_1067,In_470,In_100);
xnor U1068 (N_1068,In_699,In_620);
xor U1069 (N_1069,In_119,In_230);
xnor U1070 (N_1070,In_414,In_389);
xor U1071 (N_1071,In_480,In_612);
and U1072 (N_1072,In_515,In_470);
or U1073 (N_1073,In_482,In_265);
or U1074 (N_1074,In_223,In_717);
nor U1075 (N_1075,In_477,In_126);
and U1076 (N_1076,In_20,In_29);
nand U1077 (N_1077,In_668,In_164);
nand U1078 (N_1078,In_83,In_653);
and U1079 (N_1079,In_300,In_742);
xnor U1080 (N_1080,In_592,In_526);
or U1081 (N_1081,In_46,In_273);
nand U1082 (N_1082,In_719,In_717);
and U1083 (N_1083,In_298,In_295);
nand U1084 (N_1084,In_597,In_380);
or U1085 (N_1085,In_624,In_453);
xnor U1086 (N_1086,In_474,In_605);
nor U1087 (N_1087,In_343,In_52);
nor U1088 (N_1088,In_657,In_362);
nand U1089 (N_1089,In_359,In_105);
or U1090 (N_1090,In_250,In_643);
and U1091 (N_1091,In_366,In_326);
nor U1092 (N_1092,In_275,In_197);
or U1093 (N_1093,In_96,In_239);
xor U1094 (N_1094,In_519,In_148);
nand U1095 (N_1095,In_182,In_661);
and U1096 (N_1096,In_108,In_369);
nand U1097 (N_1097,In_231,In_401);
nand U1098 (N_1098,In_653,In_68);
and U1099 (N_1099,In_371,In_440);
nand U1100 (N_1100,In_362,In_460);
nor U1101 (N_1101,In_490,In_698);
and U1102 (N_1102,In_300,In_486);
and U1103 (N_1103,In_66,In_180);
or U1104 (N_1104,In_121,In_396);
nand U1105 (N_1105,In_198,In_208);
nor U1106 (N_1106,In_37,In_583);
or U1107 (N_1107,In_103,In_325);
nor U1108 (N_1108,In_107,In_219);
nand U1109 (N_1109,In_745,In_583);
nor U1110 (N_1110,In_128,In_255);
nand U1111 (N_1111,In_91,In_484);
xnor U1112 (N_1112,In_101,In_488);
nor U1113 (N_1113,In_403,In_233);
nand U1114 (N_1114,In_609,In_653);
or U1115 (N_1115,In_342,In_559);
nand U1116 (N_1116,In_665,In_525);
or U1117 (N_1117,In_57,In_516);
and U1118 (N_1118,In_434,In_210);
and U1119 (N_1119,In_739,In_306);
nand U1120 (N_1120,In_3,In_109);
nor U1121 (N_1121,In_339,In_354);
xnor U1122 (N_1122,In_298,In_484);
nor U1123 (N_1123,In_52,In_252);
nor U1124 (N_1124,In_379,In_429);
xor U1125 (N_1125,In_346,In_523);
nand U1126 (N_1126,In_81,In_125);
xor U1127 (N_1127,In_255,In_252);
and U1128 (N_1128,In_308,In_546);
nor U1129 (N_1129,In_62,In_53);
nand U1130 (N_1130,In_526,In_208);
nand U1131 (N_1131,In_214,In_349);
or U1132 (N_1132,In_214,In_509);
and U1133 (N_1133,In_699,In_487);
and U1134 (N_1134,In_553,In_112);
or U1135 (N_1135,In_747,In_586);
nor U1136 (N_1136,In_209,In_237);
nor U1137 (N_1137,In_733,In_117);
nor U1138 (N_1138,In_283,In_689);
nand U1139 (N_1139,In_445,In_177);
and U1140 (N_1140,In_53,In_252);
and U1141 (N_1141,In_657,In_505);
nand U1142 (N_1142,In_737,In_361);
nand U1143 (N_1143,In_259,In_266);
or U1144 (N_1144,In_391,In_407);
and U1145 (N_1145,In_737,In_279);
xnor U1146 (N_1146,In_527,In_107);
or U1147 (N_1147,In_503,In_197);
nor U1148 (N_1148,In_66,In_200);
nor U1149 (N_1149,In_383,In_13);
nor U1150 (N_1150,In_646,In_266);
xnor U1151 (N_1151,In_221,In_256);
nand U1152 (N_1152,In_201,In_562);
xnor U1153 (N_1153,In_153,In_638);
or U1154 (N_1154,In_712,In_309);
nor U1155 (N_1155,In_426,In_304);
xnor U1156 (N_1156,In_204,In_290);
or U1157 (N_1157,In_226,In_614);
nand U1158 (N_1158,In_646,In_285);
and U1159 (N_1159,In_586,In_363);
nor U1160 (N_1160,In_367,In_534);
nand U1161 (N_1161,In_184,In_180);
or U1162 (N_1162,In_472,In_271);
nand U1163 (N_1163,In_609,In_394);
nor U1164 (N_1164,In_383,In_495);
nor U1165 (N_1165,In_249,In_539);
nor U1166 (N_1166,In_84,In_21);
nand U1167 (N_1167,In_380,In_602);
xor U1168 (N_1168,In_358,In_408);
and U1169 (N_1169,In_513,In_453);
and U1170 (N_1170,In_248,In_227);
xnor U1171 (N_1171,In_365,In_171);
nor U1172 (N_1172,In_86,In_493);
and U1173 (N_1173,In_348,In_660);
nor U1174 (N_1174,In_205,In_27);
or U1175 (N_1175,In_679,In_588);
nand U1176 (N_1176,In_650,In_68);
and U1177 (N_1177,In_573,In_229);
nand U1178 (N_1178,In_258,In_632);
nand U1179 (N_1179,In_12,In_230);
nor U1180 (N_1180,In_645,In_482);
xor U1181 (N_1181,In_473,In_566);
nor U1182 (N_1182,In_22,In_679);
and U1183 (N_1183,In_284,In_533);
nand U1184 (N_1184,In_119,In_39);
nand U1185 (N_1185,In_226,In_215);
and U1186 (N_1186,In_368,In_664);
nor U1187 (N_1187,In_494,In_414);
and U1188 (N_1188,In_521,In_131);
and U1189 (N_1189,In_158,In_124);
nand U1190 (N_1190,In_677,In_91);
or U1191 (N_1191,In_312,In_353);
nand U1192 (N_1192,In_410,In_369);
and U1193 (N_1193,In_408,In_566);
nor U1194 (N_1194,In_40,In_457);
and U1195 (N_1195,In_402,In_494);
nor U1196 (N_1196,In_86,In_441);
nor U1197 (N_1197,In_388,In_124);
nand U1198 (N_1198,In_309,In_122);
nor U1199 (N_1199,In_336,In_443);
nand U1200 (N_1200,In_262,In_478);
and U1201 (N_1201,In_494,In_241);
and U1202 (N_1202,In_550,In_519);
nor U1203 (N_1203,In_660,In_429);
or U1204 (N_1204,In_322,In_567);
nand U1205 (N_1205,In_354,In_137);
xnor U1206 (N_1206,In_463,In_731);
nor U1207 (N_1207,In_334,In_482);
and U1208 (N_1208,In_554,In_185);
xnor U1209 (N_1209,In_4,In_636);
and U1210 (N_1210,In_213,In_695);
nor U1211 (N_1211,In_108,In_320);
nand U1212 (N_1212,In_158,In_95);
xor U1213 (N_1213,In_294,In_6);
and U1214 (N_1214,In_224,In_321);
and U1215 (N_1215,In_388,In_122);
nand U1216 (N_1216,In_725,In_316);
and U1217 (N_1217,In_450,In_166);
xor U1218 (N_1218,In_718,In_204);
xnor U1219 (N_1219,In_661,In_469);
and U1220 (N_1220,In_645,In_90);
or U1221 (N_1221,In_12,In_501);
or U1222 (N_1222,In_723,In_385);
nand U1223 (N_1223,In_465,In_477);
and U1224 (N_1224,In_350,In_168);
xor U1225 (N_1225,In_742,In_455);
and U1226 (N_1226,In_718,In_444);
nor U1227 (N_1227,In_229,In_616);
or U1228 (N_1228,In_135,In_245);
nor U1229 (N_1229,In_258,In_299);
nand U1230 (N_1230,In_627,In_646);
or U1231 (N_1231,In_445,In_564);
and U1232 (N_1232,In_737,In_471);
xnor U1233 (N_1233,In_609,In_117);
and U1234 (N_1234,In_289,In_707);
and U1235 (N_1235,In_208,In_563);
or U1236 (N_1236,In_63,In_510);
xnor U1237 (N_1237,In_135,In_292);
xnor U1238 (N_1238,In_79,In_546);
and U1239 (N_1239,In_350,In_104);
or U1240 (N_1240,In_183,In_328);
nand U1241 (N_1241,In_41,In_602);
nand U1242 (N_1242,In_656,In_129);
and U1243 (N_1243,In_679,In_600);
and U1244 (N_1244,In_618,In_172);
nor U1245 (N_1245,In_276,In_339);
nor U1246 (N_1246,In_743,In_254);
and U1247 (N_1247,In_579,In_457);
nor U1248 (N_1248,In_230,In_36);
or U1249 (N_1249,In_335,In_371);
xnor U1250 (N_1250,In_273,In_627);
nor U1251 (N_1251,In_554,In_660);
nor U1252 (N_1252,In_105,In_241);
xnor U1253 (N_1253,In_435,In_593);
or U1254 (N_1254,In_237,In_278);
nand U1255 (N_1255,In_13,In_262);
nor U1256 (N_1256,In_733,In_609);
and U1257 (N_1257,In_221,In_474);
nand U1258 (N_1258,In_27,In_298);
and U1259 (N_1259,In_117,In_596);
nor U1260 (N_1260,In_693,In_671);
or U1261 (N_1261,In_646,In_299);
and U1262 (N_1262,In_84,In_392);
and U1263 (N_1263,In_692,In_695);
and U1264 (N_1264,In_204,In_673);
and U1265 (N_1265,In_548,In_430);
and U1266 (N_1266,In_11,In_661);
or U1267 (N_1267,In_100,In_241);
or U1268 (N_1268,In_559,In_544);
or U1269 (N_1269,In_205,In_246);
nor U1270 (N_1270,In_715,In_366);
nor U1271 (N_1271,In_12,In_128);
and U1272 (N_1272,In_75,In_51);
and U1273 (N_1273,In_660,In_404);
xnor U1274 (N_1274,In_267,In_434);
and U1275 (N_1275,In_448,In_720);
xor U1276 (N_1276,In_466,In_695);
nor U1277 (N_1277,In_390,In_74);
and U1278 (N_1278,In_482,In_124);
nor U1279 (N_1279,In_605,In_539);
and U1280 (N_1280,In_427,In_547);
or U1281 (N_1281,In_524,In_400);
and U1282 (N_1282,In_503,In_378);
and U1283 (N_1283,In_471,In_588);
and U1284 (N_1284,In_546,In_159);
and U1285 (N_1285,In_499,In_484);
or U1286 (N_1286,In_393,In_694);
nand U1287 (N_1287,In_542,In_683);
nor U1288 (N_1288,In_310,In_400);
nor U1289 (N_1289,In_550,In_95);
xnor U1290 (N_1290,In_40,In_62);
or U1291 (N_1291,In_35,In_70);
nand U1292 (N_1292,In_73,In_125);
xor U1293 (N_1293,In_728,In_242);
nand U1294 (N_1294,In_484,In_121);
nor U1295 (N_1295,In_79,In_301);
nor U1296 (N_1296,In_593,In_709);
or U1297 (N_1297,In_139,In_591);
or U1298 (N_1298,In_568,In_681);
and U1299 (N_1299,In_94,In_390);
or U1300 (N_1300,In_645,In_146);
nor U1301 (N_1301,In_43,In_652);
nor U1302 (N_1302,In_665,In_589);
nor U1303 (N_1303,In_151,In_688);
nor U1304 (N_1304,In_40,In_60);
nor U1305 (N_1305,In_315,In_360);
and U1306 (N_1306,In_181,In_554);
nor U1307 (N_1307,In_712,In_373);
or U1308 (N_1308,In_123,In_440);
nand U1309 (N_1309,In_57,In_497);
xnor U1310 (N_1310,In_566,In_643);
or U1311 (N_1311,In_324,In_335);
and U1312 (N_1312,In_631,In_134);
and U1313 (N_1313,In_5,In_496);
nand U1314 (N_1314,In_368,In_439);
or U1315 (N_1315,In_524,In_249);
nor U1316 (N_1316,In_181,In_503);
xnor U1317 (N_1317,In_584,In_684);
nand U1318 (N_1318,In_640,In_0);
and U1319 (N_1319,In_624,In_294);
or U1320 (N_1320,In_685,In_471);
nor U1321 (N_1321,In_123,In_391);
xnor U1322 (N_1322,In_166,In_252);
nor U1323 (N_1323,In_261,In_29);
nor U1324 (N_1324,In_302,In_389);
or U1325 (N_1325,In_391,In_137);
nand U1326 (N_1326,In_242,In_105);
or U1327 (N_1327,In_683,In_234);
xor U1328 (N_1328,In_497,In_225);
or U1329 (N_1329,In_450,In_468);
nand U1330 (N_1330,In_1,In_43);
nand U1331 (N_1331,In_150,In_45);
or U1332 (N_1332,In_199,In_233);
nand U1333 (N_1333,In_344,In_369);
xor U1334 (N_1334,In_332,In_372);
and U1335 (N_1335,In_469,In_396);
or U1336 (N_1336,In_110,In_458);
xor U1337 (N_1337,In_612,In_425);
or U1338 (N_1338,In_635,In_418);
xnor U1339 (N_1339,In_315,In_290);
nor U1340 (N_1340,In_8,In_501);
nor U1341 (N_1341,In_607,In_589);
or U1342 (N_1342,In_330,In_66);
xnor U1343 (N_1343,In_23,In_244);
nor U1344 (N_1344,In_670,In_489);
and U1345 (N_1345,In_433,In_389);
or U1346 (N_1346,In_149,In_99);
or U1347 (N_1347,In_292,In_569);
or U1348 (N_1348,In_279,In_215);
nor U1349 (N_1349,In_482,In_495);
nand U1350 (N_1350,In_430,In_450);
or U1351 (N_1351,In_163,In_205);
nor U1352 (N_1352,In_672,In_172);
nand U1353 (N_1353,In_96,In_686);
and U1354 (N_1354,In_14,In_742);
nor U1355 (N_1355,In_298,In_555);
nand U1356 (N_1356,In_297,In_429);
or U1357 (N_1357,In_336,In_287);
xor U1358 (N_1358,In_312,In_132);
xnor U1359 (N_1359,In_687,In_47);
nand U1360 (N_1360,In_45,In_145);
xor U1361 (N_1361,In_386,In_342);
xnor U1362 (N_1362,In_310,In_567);
nor U1363 (N_1363,In_489,In_61);
and U1364 (N_1364,In_651,In_525);
nor U1365 (N_1365,In_564,In_292);
nor U1366 (N_1366,In_23,In_265);
and U1367 (N_1367,In_409,In_262);
nor U1368 (N_1368,In_271,In_489);
nor U1369 (N_1369,In_39,In_335);
and U1370 (N_1370,In_603,In_687);
nor U1371 (N_1371,In_69,In_632);
xor U1372 (N_1372,In_733,In_132);
or U1373 (N_1373,In_20,In_438);
xor U1374 (N_1374,In_599,In_330);
and U1375 (N_1375,In_638,In_482);
nand U1376 (N_1376,In_254,In_677);
xnor U1377 (N_1377,In_512,In_534);
and U1378 (N_1378,In_116,In_373);
and U1379 (N_1379,In_10,In_400);
or U1380 (N_1380,In_591,In_128);
xor U1381 (N_1381,In_163,In_451);
or U1382 (N_1382,In_321,In_570);
xnor U1383 (N_1383,In_653,In_516);
nor U1384 (N_1384,In_141,In_243);
nor U1385 (N_1385,In_596,In_291);
or U1386 (N_1386,In_640,In_516);
and U1387 (N_1387,In_709,In_499);
or U1388 (N_1388,In_7,In_79);
and U1389 (N_1389,In_331,In_641);
nor U1390 (N_1390,In_309,In_183);
xor U1391 (N_1391,In_550,In_50);
and U1392 (N_1392,In_722,In_605);
xor U1393 (N_1393,In_75,In_458);
nand U1394 (N_1394,In_65,In_390);
and U1395 (N_1395,In_705,In_303);
and U1396 (N_1396,In_569,In_543);
nor U1397 (N_1397,In_659,In_295);
or U1398 (N_1398,In_150,In_663);
and U1399 (N_1399,In_98,In_43);
xor U1400 (N_1400,In_571,In_621);
and U1401 (N_1401,In_650,In_70);
nand U1402 (N_1402,In_355,In_576);
or U1403 (N_1403,In_428,In_547);
nor U1404 (N_1404,In_507,In_294);
xor U1405 (N_1405,In_172,In_727);
nand U1406 (N_1406,In_569,In_503);
or U1407 (N_1407,In_444,In_213);
nand U1408 (N_1408,In_731,In_520);
nand U1409 (N_1409,In_218,In_445);
nor U1410 (N_1410,In_685,In_97);
or U1411 (N_1411,In_63,In_21);
nand U1412 (N_1412,In_542,In_454);
xnor U1413 (N_1413,In_288,In_568);
or U1414 (N_1414,In_721,In_579);
nand U1415 (N_1415,In_717,In_482);
and U1416 (N_1416,In_744,In_346);
and U1417 (N_1417,In_545,In_195);
xor U1418 (N_1418,In_418,In_487);
nor U1419 (N_1419,In_105,In_315);
nor U1420 (N_1420,In_317,In_438);
xnor U1421 (N_1421,In_25,In_285);
or U1422 (N_1422,In_251,In_721);
nor U1423 (N_1423,In_576,In_397);
nand U1424 (N_1424,In_137,In_218);
nor U1425 (N_1425,In_550,In_340);
nor U1426 (N_1426,In_742,In_677);
nor U1427 (N_1427,In_530,In_154);
nand U1428 (N_1428,In_375,In_451);
xnor U1429 (N_1429,In_573,In_685);
xnor U1430 (N_1430,In_717,In_201);
or U1431 (N_1431,In_523,In_586);
xor U1432 (N_1432,In_626,In_187);
or U1433 (N_1433,In_41,In_99);
nand U1434 (N_1434,In_75,In_401);
and U1435 (N_1435,In_678,In_271);
and U1436 (N_1436,In_642,In_56);
nand U1437 (N_1437,In_407,In_495);
nor U1438 (N_1438,In_366,In_562);
xnor U1439 (N_1439,In_533,In_255);
nand U1440 (N_1440,In_520,In_289);
or U1441 (N_1441,In_348,In_547);
or U1442 (N_1442,In_405,In_610);
nand U1443 (N_1443,In_591,In_545);
xor U1444 (N_1444,In_456,In_324);
and U1445 (N_1445,In_552,In_506);
xor U1446 (N_1446,In_120,In_101);
and U1447 (N_1447,In_726,In_352);
and U1448 (N_1448,In_190,In_96);
and U1449 (N_1449,In_645,In_287);
and U1450 (N_1450,In_360,In_77);
and U1451 (N_1451,In_590,In_638);
and U1452 (N_1452,In_55,In_417);
and U1453 (N_1453,In_472,In_681);
xor U1454 (N_1454,In_82,In_0);
xor U1455 (N_1455,In_252,In_248);
nand U1456 (N_1456,In_204,In_661);
or U1457 (N_1457,In_745,In_140);
nand U1458 (N_1458,In_693,In_257);
xnor U1459 (N_1459,In_272,In_106);
nand U1460 (N_1460,In_598,In_470);
nand U1461 (N_1461,In_186,In_469);
or U1462 (N_1462,In_19,In_413);
nor U1463 (N_1463,In_531,In_557);
nor U1464 (N_1464,In_138,In_722);
nor U1465 (N_1465,In_2,In_499);
nor U1466 (N_1466,In_703,In_295);
or U1467 (N_1467,In_609,In_521);
or U1468 (N_1468,In_393,In_685);
and U1469 (N_1469,In_42,In_472);
and U1470 (N_1470,In_293,In_116);
or U1471 (N_1471,In_188,In_209);
or U1472 (N_1472,In_58,In_538);
nand U1473 (N_1473,In_263,In_321);
nor U1474 (N_1474,In_98,In_597);
nor U1475 (N_1475,In_127,In_521);
nor U1476 (N_1476,In_715,In_400);
and U1477 (N_1477,In_71,In_9);
nor U1478 (N_1478,In_712,In_79);
or U1479 (N_1479,In_429,In_645);
and U1480 (N_1480,In_427,In_425);
nor U1481 (N_1481,In_707,In_552);
and U1482 (N_1482,In_697,In_589);
xnor U1483 (N_1483,In_492,In_159);
nand U1484 (N_1484,In_480,In_109);
nand U1485 (N_1485,In_110,In_3);
xor U1486 (N_1486,In_659,In_191);
xnor U1487 (N_1487,In_574,In_608);
nand U1488 (N_1488,In_52,In_710);
or U1489 (N_1489,In_625,In_544);
nand U1490 (N_1490,In_332,In_348);
nand U1491 (N_1491,In_615,In_450);
or U1492 (N_1492,In_505,In_296);
xor U1493 (N_1493,In_693,In_238);
xor U1494 (N_1494,In_577,In_55);
nand U1495 (N_1495,In_728,In_159);
nor U1496 (N_1496,In_22,In_741);
or U1497 (N_1497,In_311,In_362);
and U1498 (N_1498,In_144,In_298);
nand U1499 (N_1499,In_613,In_199);
xnor U1500 (N_1500,In_72,In_517);
and U1501 (N_1501,In_120,In_637);
and U1502 (N_1502,In_481,In_637);
and U1503 (N_1503,In_615,In_75);
xor U1504 (N_1504,In_111,In_137);
nand U1505 (N_1505,In_362,In_86);
xnor U1506 (N_1506,In_536,In_242);
nor U1507 (N_1507,In_638,In_370);
nor U1508 (N_1508,In_718,In_467);
or U1509 (N_1509,In_199,In_561);
nand U1510 (N_1510,In_122,In_205);
nor U1511 (N_1511,In_583,In_28);
or U1512 (N_1512,In_23,In_182);
xor U1513 (N_1513,In_385,In_156);
nor U1514 (N_1514,In_40,In_701);
and U1515 (N_1515,In_472,In_713);
xnor U1516 (N_1516,In_436,In_495);
xnor U1517 (N_1517,In_428,In_352);
nor U1518 (N_1518,In_45,In_11);
nand U1519 (N_1519,In_320,In_409);
nor U1520 (N_1520,In_247,In_43);
nand U1521 (N_1521,In_627,In_534);
nor U1522 (N_1522,In_132,In_107);
nor U1523 (N_1523,In_580,In_292);
or U1524 (N_1524,In_464,In_401);
xnor U1525 (N_1525,In_351,In_63);
nand U1526 (N_1526,In_487,In_184);
or U1527 (N_1527,In_747,In_409);
or U1528 (N_1528,In_517,In_124);
nor U1529 (N_1529,In_480,In_175);
nand U1530 (N_1530,In_344,In_82);
or U1531 (N_1531,In_550,In_32);
or U1532 (N_1532,In_228,In_205);
nand U1533 (N_1533,In_389,In_563);
and U1534 (N_1534,In_264,In_333);
nor U1535 (N_1535,In_292,In_121);
or U1536 (N_1536,In_510,In_290);
or U1537 (N_1537,In_606,In_251);
xor U1538 (N_1538,In_744,In_10);
nor U1539 (N_1539,In_716,In_277);
xnor U1540 (N_1540,In_369,In_248);
and U1541 (N_1541,In_673,In_429);
nor U1542 (N_1542,In_349,In_146);
and U1543 (N_1543,In_732,In_16);
xor U1544 (N_1544,In_105,In_166);
xor U1545 (N_1545,In_54,In_104);
nor U1546 (N_1546,In_217,In_175);
and U1547 (N_1547,In_313,In_228);
nand U1548 (N_1548,In_568,In_217);
nand U1549 (N_1549,In_405,In_311);
or U1550 (N_1550,In_478,In_85);
nand U1551 (N_1551,In_428,In_161);
nand U1552 (N_1552,In_149,In_235);
xnor U1553 (N_1553,In_415,In_54);
xnor U1554 (N_1554,In_708,In_18);
nand U1555 (N_1555,In_152,In_314);
and U1556 (N_1556,In_134,In_150);
xnor U1557 (N_1557,In_70,In_540);
and U1558 (N_1558,In_690,In_105);
nand U1559 (N_1559,In_152,In_700);
nor U1560 (N_1560,In_64,In_298);
xor U1561 (N_1561,In_106,In_688);
nor U1562 (N_1562,In_531,In_338);
xor U1563 (N_1563,In_551,In_361);
and U1564 (N_1564,In_489,In_535);
xor U1565 (N_1565,In_526,In_660);
xor U1566 (N_1566,In_229,In_453);
nor U1567 (N_1567,In_369,In_606);
nor U1568 (N_1568,In_280,In_313);
and U1569 (N_1569,In_188,In_156);
and U1570 (N_1570,In_708,In_592);
or U1571 (N_1571,In_348,In_255);
or U1572 (N_1572,In_603,In_659);
xnor U1573 (N_1573,In_594,In_12);
or U1574 (N_1574,In_441,In_637);
nand U1575 (N_1575,In_558,In_33);
or U1576 (N_1576,In_130,In_546);
nor U1577 (N_1577,In_693,In_303);
xor U1578 (N_1578,In_329,In_367);
or U1579 (N_1579,In_609,In_191);
xnor U1580 (N_1580,In_20,In_296);
xor U1581 (N_1581,In_649,In_628);
nand U1582 (N_1582,In_462,In_84);
and U1583 (N_1583,In_674,In_99);
and U1584 (N_1584,In_381,In_370);
xnor U1585 (N_1585,In_651,In_46);
xnor U1586 (N_1586,In_368,In_662);
nand U1587 (N_1587,In_245,In_144);
nand U1588 (N_1588,In_353,In_271);
nor U1589 (N_1589,In_352,In_305);
or U1590 (N_1590,In_335,In_708);
nand U1591 (N_1591,In_187,In_591);
and U1592 (N_1592,In_658,In_456);
and U1593 (N_1593,In_133,In_86);
or U1594 (N_1594,In_564,In_447);
xnor U1595 (N_1595,In_361,In_399);
nor U1596 (N_1596,In_541,In_100);
and U1597 (N_1597,In_527,In_51);
or U1598 (N_1598,In_183,In_629);
nand U1599 (N_1599,In_738,In_519);
nand U1600 (N_1600,In_706,In_235);
nor U1601 (N_1601,In_401,In_713);
nor U1602 (N_1602,In_416,In_162);
xor U1603 (N_1603,In_476,In_524);
nor U1604 (N_1604,In_65,In_98);
nor U1605 (N_1605,In_248,In_486);
or U1606 (N_1606,In_639,In_154);
nor U1607 (N_1607,In_324,In_613);
nand U1608 (N_1608,In_625,In_46);
nand U1609 (N_1609,In_99,In_711);
nand U1610 (N_1610,In_17,In_689);
or U1611 (N_1611,In_744,In_258);
nor U1612 (N_1612,In_183,In_21);
nand U1613 (N_1613,In_383,In_545);
nor U1614 (N_1614,In_522,In_107);
nor U1615 (N_1615,In_408,In_46);
and U1616 (N_1616,In_494,In_269);
nand U1617 (N_1617,In_620,In_623);
or U1618 (N_1618,In_358,In_119);
or U1619 (N_1619,In_690,In_747);
nor U1620 (N_1620,In_442,In_111);
nor U1621 (N_1621,In_569,In_20);
nand U1622 (N_1622,In_739,In_169);
nand U1623 (N_1623,In_732,In_357);
or U1624 (N_1624,In_400,In_613);
nor U1625 (N_1625,In_706,In_276);
and U1626 (N_1626,In_393,In_294);
or U1627 (N_1627,In_63,In_600);
and U1628 (N_1628,In_336,In_282);
and U1629 (N_1629,In_141,In_744);
or U1630 (N_1630,In_469,In_520);
and U1631 (N_1631,In_483,In_729);
or U1632 (N_1632,In_560,In_228);
nand U1633 (N_1633,In_580,In_255);
and U1634 (N_1634,In_706,In_594);
nor U1635 (N_1635,In_739,In_163);
xor U1636 (N_1636,In_112,In_62);
and U1637 (N_1637,In_418,In_598);
nor U1638 (N_1638,In_300,In_735);
xnor U1639 (N_1639,In_489,In_348);
xnor U1640 (N_1640,In_573,In_197);
xnor U1641 (N_1641,In_391,In_177);
nor U1642 (N_1642,In_131,In_535);
and U1643 (N_1643,In_43,In_169);
xnor U1644 (N_1644,In_479,In_3);
nand U1645 (N_1645,In_669,In_677);
nor U1646 (N_1646,In_628,In_389);
xnor U1647 (N_1647,In_78,In_560);
xor U1648 (N_1648,In_174,In_639);
and U1649 (N_1649,In_613,In_536);
and U1650 (N_1650,In_456,In_676);
xor U1651 (N_1651,In_251,In_735);
and U1652 (N_1652,In_77,In_80);
or U1653 (N_1653,In_176,In_309);
and U1654 (N_1654,In_14,In_601);
xnor U1655 (N_1655,In_553,In_9);
or U1656 (N_1656,In_524,In_611);
xnor U1657 (N_1657,In_373,In_625);
or U1658 (N_1658,In_406,In_144);
or U1659 (N_1659,In_723,In_58);
and U1660 (N_1660,In_297,In_534);
nand U1661 (N_1661,In_653,In_234);
nand U1662 (N_1662,In_156,In_197);
or U1663 (N_1663,In_396,In_163);
and U1664 (N_1664,In_68,In_183);
xnor U1665 (N_1665,In_587,In_334);
xnor U1666 (N_1666,In_695,In_197);
xor U1667 (N_1667,In_16,In_1);
nand U1668 (N_1668,In_558,In_648);
nand U1669 (N_1669,In_163,In_167);
nor U1670 (N_1670,In_91,In_649);
xor U1671 (N_1671,In_491,In_455);
nor U1672 (N_1672,In_18,In_236);
and U1673 (N_1673,In_723,In_663);
nand U1674 (N_1674,In_695,In_460);
nor U1675 (N_1675,In_647,In_66);
and U1676 (N_1676,In_685,In_167);
and U1677 (N_1677,In_510,In_618);
or U1678 (N_1678,In_548,In_550);
nor U1679 (N_1679,In_305,In_197);
nand U1680 (N_1680,In_435,In_67);
xor U1681 (N_1681,In_16,In_448);
or U1682 (N_1682,In_529,In_249);
nor U1683 (N_1683,In_635,In_657);
xor U1684 (N_1684,In_459,In_135);
nand U1685 (N_1685,In_465,In_617);
or U1686 (N_1686,In_22,In_622);
nor U1687 (N_1687,In_421,In_252);
nand U1688 (N_1688,In_313,In_713);
and U1689 (N_1689,In_384,In_608);
and U1690 (N_1690,In_152,In_48);
nand U1691 (N_1691,In_234,In_597);
nand U1692 (N_1692,In_252,In_144);
nand U1693 (N_1693,In_349,In_675);
and U1694 (N_1694,In_675,In_343);
xor U1695 (N_1695,In_243,In_11);
nor U1696 (N_1696,In_49,In_118);
nand U1697 (N_1697,In_447,In_343);
nand U1698 (N_1698,In_188,In_476);
and U1699 (N_1699,In_208,In_144);
or U1700 (N_1700,In_212,In_501);
and U1701 (N_1701,In_489,In_119);
nor U1702 (N_1702,In_386,In_129);
and U1703 (N_1703,In_527,In_649);
and U1704 (N_1704,In_259,In_114);
and U1705 (N_1705,In_691,In_526);
or U1706 (N_1706,In_136,In_167);
or U1707 (N_1707,In_724,In_325);
nand U1708 (N_1708,In_538,In_532);
and U1709 (N_1709,In_537,In_6);
xor U1710 (N_1710,In_650,In_273);
and U1711 (N_1711,In_696,In_95);
xor U1712 (N_1712,In_355,In_494);
or U1713 (N_1713,In_701,In_437);
or U1714 (N_1714,In_271,In_595);
nor U1715 (N_1715,In_437,In_472);
nor U1716 (N_1716,In_572,In_176);
nand U1717 (N_1717,In_506,In_597);
xor U1718 (N_1718,In_730,In_28);
and U1719 (N_1719,In_226,In_71);
and U1720 (N_1720,In_165,In_586);
nor U1721 (N_1721,In_90,In_720);
and U1722 (N_1722,In_84,In_685);
nor U1723 (N_1723,In_229,In_343);
and U1724 (N_1724,In_399,In_522);
xnor U1725 (N_1725,In_205,In_548);
nand U1726 (N_1726,In_413,In_657);
nor U1727 (N_1727,In_210,In_2);
nand U1728 (N_1728,In_166,In_402);
nor U1729 (N_1729,In_699,In_88);
and U1730 (N_1730,In_29,In_483);
or U1731 (N_1731,In_202,In_332);
nand U1732 (N_1732,In_576,In_366);
and U1733 (N_1733,In_735,In_698);
nor U1734 (N_1734,In_544,In_445);
xor U1735 (N_1735,In_375,In_552);
nand U1736 (N_1736,In_664,In_2);
nor U1737 (N_1737,In_721,In_210);
or U1738 (N_1738,In_682,In_730);
nor U1739 (N_1739,In_36,In_220);
xor U1740 (N_1740,In_561,In_480);
xnor U1741 (N_1741,In_303,In_493);
xnor U1742 (N_1742,In_233,In_381);
or U1743 (N_1743,In_687,In_365);
nand U1744 (N_1744,In_613,In_484);
and U1745 (N_1745,In_584,In_18);
nand U1746 (N_1746,In_252,In_228);
or U1747 (N_1747,In_720,In_583);
and U1748 (N_1748,In_644,In_271);
nor U1749 (N_1749,In_560,In_113);
xnor U1750 (N_1750,In_212,In_725);
and U1751 (N_1751,In_246,In_343);
xnor U1752 (N_1752,In_547,In_332);
nand U1753 (N_1753,In_343,In_45);
nand U1754 (N_1754,In_185,In_168);
xor U1755 (N_1755,In_726,In_404);
nand U1756 (N_1756,In_531,In_405);
xnor U1757 (N_1757,In_605,In_70);
nand U1758 (N_1758,In_360,In_324);
xnor U1759 (N_1759,In_400,In_538);
and U1760 (N_1760,In_661,In_161);
nor U1761 (N_1761,In_285,In_223);
and U1762 (N_1762,In_483,In_340);
xor U1763 (N_1763,In_579,In_569);
nand U1764 (N_1764,In_142,In_117);
or U1765 (N_1765,In_271,In_596);
nor U1766 (N_1766,In_46,In_660);
or U1767 (N_1767,In_87,In_518);
xor U1768 (N_1768,In_318,In_229);
or U1769 (N_1769,In_54,In_464);
and U1770 (N_1770,In_222,In_282);
and U1771 (N_1771,In_610,In_52);
xnor U1772 (N_1772,In_433,In_131);
xor U1773 (N_1773,In_180,In_686);
nor U1774 (N_1774,In_723,In_749);
and U1775 (N_1775,In_740,In_361);
or U1776 (N_1776,In_455,In_453);
and U1777 (N_1777,In_535,In_291);
nor U1778 (N_1778,In_133,In_737);
nor U1779 (N_1779,In_603,In_512);
xor U1780 (N_1780,In_161,In_336);
nand U1781 (N_1781,In_646,In_700);
and U1782 (N_1782,In_729,In_569);
nor U1783 (N_1783,In_438,In_623);
and U1784 (N_1784,In_719,In_103);
nand U1785 (N_1785,In_146,In_119);
or U1786 (N_1786,In_361,In_243);
nor U1787 (N_1787,In_568,In_80);
and U1788 (N_1788,In_44,In_9);
nand U1789 (N_1789,In_237,In_9);
nand U1790 (N_1790,In_460,In_541);
and U1791 (N_1791,In_491,In_115);
or U1792 (N_1792,In_649,In_437);
xnor U1793 (N_1793,In_59,In_117);
or U1794 (N_1794,In_397,In_18);
nand U1795 (N_1795,In_51,In_403);
nor U1796 (N_1796,In_585,In_429);
nand U1797 (N_1797,In_120,In_49);
nor U1798 (N_1798,In_394,In_521);
nand U1799 (N_1799,In_465,In_65);
nand U1800 (N_1800,In_127,In_255);
nor U1801 (N_1801,In_180,In_620);
xnor U1802 (N_1802,In_320,In_169);
or U1803 (N_1803,In_297,In_138);
xor U1804 (N_1804,In_324,In_214);
nand U1805 (N_1805,In_711,In_616);
xnor U1806 (N_1806,In_35,In_348);
or U1807 (N_1807,In_369,In_652);
or U1808 (N_1808,In_187,In_597);
nand U1809 (N_1809,In_626,In_597);
or U1810 (N_1810,In_553,In_317);
or U1811 (N_1811,In_362,In_342);
nor U1812 (N_1812,In_548,In_745);
and U1813 (N_1813,In_68,In_122);
nand U1814 (N_1814,In_425,In_104);
nor U1815 (N_1815,In_638,In_649);
and U1816 (N_1816,In_667,In_534);
or U1817 (N_1817,In_78,In_581);
nor U1818 (N_1818,In_40,In_144);
xnor U1819 (N_1819,In_614,In_79);
nand U1820 (N_1820,In_115,In_127);
nor U1821 (N_1821,In_206,In_640);
nand U1822 (N_1822,In_526,In_262);
nor U1823 (N_1823,In_474,In_179);
nor U1824 (N_1824,In_358,In_102);
xor U1825 (N_1825,In_533,In_701);
or U1826 (N_1826,In_110,In_385);
nand U1827 (N_1827,In_3,In_556);
nor U1828 (N_1828,In_164,In_663);
or U1829 (N_1829,In_449,In_733);
nand U1830 (N_1830,In_437,In_605);
nand U1831 (N_1831,In_676,In_65);
nor U1832 (N_1832,In_165,In_160);
nor U1833 (N_1833,In_392,In_633);
nand U1834 (N_1834,In_398,In_718);
nand U1835 (N_1835,In_447,In_519);
and U1836 (N_1836,In_254,In_568);
nand U1837 (N_1837,In_115,In_307);
or U1838 (N_1838,In_352,In_510);
or U1839 (N_1839,In_127,In_407);
xor U1840 (N_1840,In_186,In_743);
nand U1841 (N_1841,In_441,In_742);
nand U1842 (N_1842,In_465,In_524);
nor U1843 (N_1843,In_733,In_143);
nand U1844 (N_1844,In_55,In_268);
nand U1845 (N_1845,In_121,In_643);
or U1846 (N_1846,In_367,In_545);
nor U1847 (N_1847,In_81,In_174);
and U1848 (N_1848,In_80,In_416);
nor U1849 (N_1849,In_532,In_609);
nor U1850 (N_1850,In_379,In_748);
nor U1851 (N_1851,In_410,In_678);
and U1852 (N_1852,In_330,In_217);
xor U1853 (N_1853,In_309,In_178);
nand U1854 (N_1854,In_748,In_403);
and U1855 (N_1855,In_339,In_15);
nor U1856 (N_1856,In_241,In_582);
nand U1857 (N_1857,In_308,In_688);
and U1858 (N_1858,In_2,In_645);
nor U1859 (N_1859,In_4,In_266);
and U1860 (N_1860,In_723,In_273);
and U1861 (N_1861,In_161,In_52);
or U1862 (N_1862,In_355,In_45);
nand U1863 (N_1863,In_453,In_369);
and U1864 (N_1864,In_518,In_249);
xor U1865 (N_1865,In_196,In_325);
xnor U1866 (N_1866,In_644,In_98);
nand U1867 (N_1867,In_712,In_333);
or U1868 (N_1868,In_41,In_115);
nor U1869 (N_1869,In_373,In_343);
or U1870 (N_1870,In_79,In_502);
or U1871 (N_1871,In_475,In_8);
nand U1872 (N_1872,In_310,In_664);
nand U1873 (N_1873,In_702,In_462);
xor U1874 (N_1874,In_528,In_612);
nor U1875 (N_1875,In_290,In_549);
or U1876 (N_1876,In_285,In_575);
and U1877 (N_1877,In_127,In_294);
xor U1878 (N_1878,In_550,In_459);
nor U1879 (N_1879,In_353,In_575);
and U1880 (N_1880,In_718,In_225);
xor U1881 (N_1881,In_143,In_363);
and U1882 (N_1882,In_338,In_249);
and U1883 (N_1883,In_542,In_28);
and U1884 (N_1884,In_708,In_483);
or U1885 (N_1885,In_167,In_174);
nand U1886 (N_1886,In_413,In_597);
or U1887 (N_1887,In_169,In_108);
nand U1888 (N_1888,In_374,In_614);
and U1889 (N_1889,In_401,In_51);
nand U1890 (N_1890,In_127,In_424);
or U1891 (N_1891,In_250,In_388);
nor U1892 (N_1892,In_164,In_596);
nor U1893 (N_1893,In_591,In_81);
nor U1894 (N_1894,In_464,In_301);
or U1895 (N_1895,In_279,In_455);
nor U1896 (N_1896,In_482,In_599);
nand U1897 (N_1897,In_575,In_150);
xnor U1898 (N_1898,In_501,In_624);
and U1899 (N_1899,In_683,In_303);
or U1900 (N_1900,In_133,In_548);
and U1901 (N_1901,In_500,In_75);
or U1902 (N_1902,In_485,In_587);
or U1903 (N_1903,In_172,In_680);
xnor U1904 (N_1904,In_575,In_244);
xnor U1905 (N_1905,In_341,In_745);
xnor U1906 (N_1906,In_742,In_485);
or U1907 (N_1907,In_609,In_651);
and U1908 (N_1908,In_14,In_575);
nor U1909 (N_1909,In_473,In_3);
or U1910 (N_1910,In_236,In_559);
nor U1911 (N_1911,In_340,In_436);
or U1912 (N_1912,In_16,In_315);
or U1913 (N_1913,In_415,In_676);
nand U1914 (N_1914,In_156,In_720);
xor U1915 (N_1915,In_741,In_270);
nand U1916 (N_1916,In_540,In_73);
or U1917 (N_1917,In_287,In_679);
xor U1918 (N_1918,In_626,In_152);
or U1919 (N_1919,In_649,In_392);
nand U1920 (N_1920,In_73,In_340);
nand U1921 (N_1921,In_382,In_299);
nand U1922 (N_1922,In_235,In_343);
nand U1923 (N_1923,In_75,In_639);
nand U1924 (N_1924,In_246,In_302);
or U1925 (N_1925,In_90,In_561);
xor U1926 (N_1926,In_123,In_636);
nor U1927 (N_1927,In_218,In_490);
and U1928 (N_1928,In_538,In_246);
or U1929 (N_1929,In_561,In_98);
nor U1930 (N_1930,In_746,In_182);
or U1931 (N_1931,In_20,In_191);
nor U1932 (N_1932,In_429,In_683);
or U1933 (N_1933,In_544,In_505);
nand U1934 (N_1934,In_184,In_476);
and U1935 (N_1935,In_621,In_155);
xor U1936 (N_1936,In_305,In_435);
or U1937 (N_1937,In_38,In_242);
nand U1938 (N_1938,In_337,In_203);
or U1939 (N_1939,In_412,In_429);
or U1940 (N_1940,In_254,In_565);
nor U1941 (N_1941,In_528,In_53);
nand U1942 (N_1942,In_585,In_727);
and U1943 (N_1943,In_558,In_310);
or U1944 (N_1944,In_320,In_328);
or U1945 (N_1945,In_89,In_313);
nand U1946 (N_1946,In_299,In_657);
nor U1947 (N_1947,In_298,In_442);
nand U1948 (N_1948,In_248,In_533);
and U1949 (N_1949,In_366,In_204);
or U1950 (N_1950,In_609,In_62);
xor U1951 (N_1951,In_128,In_560);
nand U1952 (N_1952,In_594,In_677);
nand U1953 (N_1953,In_212,In_392);
xnor U1954 (N_1954,In_87,In_636);
and U1955 (N_1955,In_83,In_487);
xnor U1956 (N_1956,In_601,In_400);
nor U1957 (N_1957,In_205,In_463);
and U1958 (N_1958,In_591,In_335);
nand U1959 (N_1959,In_153,In_446);
nor U1960 (N_1960,In_675,In_44);
nand U1961 (N_1961,In_303,In_178);
nand U1962 (N_1962,In_547,In_721);
and U1963 (N_1963,In_675,In_168);
xnor U1964 (N_1964,In_301,In_607);
or U1965 (N_1965,In_494,In_608);
and U1966 (N_1966,In_442,In_408);
or U1967 (N_1967,In_434,In_656);
and U1968 (N_1968,In_431,In_736);
nand U1969 (N_1969,In_541,In_185);
nor U1970 (N_1970,In_486,In_610);
nor U1971 (N_1971,In_714,In_568);
nand U1972 (N_1972,In_392,In_165);
or U1973 (N_1973,In_648,In_70);
or U1974 (N_1974,In_440,In_162);
nor U1975 (N_1975,In_729,In_555);
and U1976 (N_1976,In_620,In_399);
nand U1977 (N_1977,In_191,In_599);
nor U1978 (N_1978,In_402,In_435);
nor U1979 (N_1979,In_239,In_162);
or U1980 (N_1980,In_527,In_691);
nand U1981 (N_1981,In_73,In_243);
xnor U1982 (N_1982,In_239,In_554);
nand U1983 (N_1983,In_692,In_310);
nor U1984 (N_1984,In_176,In_533);
nand U1985 (N_1985,In_673,In_347);
nand U1986 (N_1986,In_216,In_189);
nor U1987 (N_1987,In_388,In_365);
or U1988 (N_1988,In_461,In_682);
nand U1989 (N_1989,In_42,In_43);
xnor U1990 (N_1990,In_520,In_295);
and U1991 (N_1991,In_698,In_55);
nand U1992 (N_1992,In_337,In_186);
xor U1993 (N_1993,In_668,In_598);
and U1994 (N_1994,In_2,In_169);
nor U1995 (N_1995,In_21,In_156);
nor U1996 (N_1996,In_219,In_273);
or U1997 (N_1997,In_129,In_350);
nor U1998 (N_1998,In_746,In_578);
nand U1999 (N_1999,In_318,In_144);
xor U2000 (N_2000,In_190,In_405);
xnor U2001 (N_2001,In_745,In_454);
nand U2002 (N_2002,In_683,In_411);
nor U2003 (N_2003,In_450,In_551);
xor U2004 (N_2004,In_291,In_682);
xor U2005 (N_2005,In_88,In_47);
or U2006 (N_2006,In_68,In_54);
and U2007 (N_2007,In_350,In_397);
xnor U2008 (N_2008,In_369,In_235);
nor U2009 (N_2009,In_569,In_332);
and U2010 (N_2010,In_119,In_414);
nor U2011 (N_2011,In_573,In_498);
or U2012 (N_2012,In_510,In_674);
or U2013 (N_2013,In_492,In_17);
and U2014 (N_2014,In_463,In_505);
nor U2015 (N_2015,In_104,In_545);
or U2016 (N_2016,In_58,In_726);
nor U2017 (N_2017,In_629,In_331);
and U2018 (N_2018,In_482,In_370);
or U2019 (N_2019,In_668,In_337);
nand U2020 (N_2020,In_151,In_639);
nor U2021 (N_2021,In_412,In_189);
nor U2022 (N_2022,In_241,In_544);
nor U2023 (N_2023,In_570,In_693);
nand U2024 (N_2024,In_448,In_403);
nand U2025 (N_2025,In_597,In_60);
nor U2026 (N_2026,In_515,In_710);
nor U2027 (N_2027,In_46,In_634);
xor U2028 (N_2028,In_128,In_582);
or U2029 (N_2029,In_252,In_34);
nor U2030 (N_2030,In_486,In_413);
and U2031 (N_2031,In_175,In_68);
or U2032 (N_2032,In_178,In_331);
nand U2033 (N_2033,In_677,In_688);
xnor U2034 (N_2034,In_404,In_79);
nor U2035 (N_2035,In_165,In_493);
nor U2036 (N_2036,In_540,In_452);
nand U2037 (N_2037,In_389,In_633);
nand U2038 (N_2038,In_71,In_430);
and U2039 (N_2039,In_32,In_261);
and U2040 (N_2040,In_409,In_37);
nor U2041 (N_2041,In_445,In_613);
nor U2042 (N_2042,In_245,In_533);
xnor U2043 (N_2043,In_224,In_524);
nor U2044 (N_2044,In_467,In_348);
nand U2045 (N_2045,In_247,In_110);
nor U2046 (N_2046,In_478,In_480);
xor U2047 (N_2047,In_550,In_464);
xnor U2048 (N_2048,In_323,In_577);
or U2049 (N_2049,In_467,In_712);
nand U2050 (N_2050,In_232,In_278);
and U2051 (N_2051,In_661,In_525);
or U2052 (N_2052,In_672,In_1);
xnor U2053 (N_2053,In_224,In_421);
or U2054 (N_2054,In_536,In_576);
and U2055 (N_2055,In_440,In_185);
or U2056 (N_2056,In_734,In_151);
xnor U2057 (N_2057,In_305,In_693);
or U2058 (N_2058,In_252,In_402);
and U2059 (N_2059,In_13,In_134);
nand U2060 (N_2060,In_248,In_356);
xor U2061 (N_2061,In_124,In_446);
and U2062 (N_2062,In_405,In_282);
and U2063 (N_2063,In_271,In_710);
nand U2064 (N_2064,In_700,In_36);
or U2065 (N_2065,In_663,In_210);
or U2066 (N_2066,In_461,In_734);
nor U2067 (N_2067,In_376,In_583);
nor U2068 (N_2068,In_6,In_559);
nor U2069 (N_2069,In_34,In_318);
xor U2070 (N_2070,In_346,In_419);
xnor U2071 (N_2071,In_727,In_562);
nor U2072 (N_2072,In_401,In_382);
xnor U2073 (N_2073,In_700,In_732);
nor U2074 (N_2074,In_15,In_344);
nor U2075 (N_2075,In_630,In_133);
or U2076 (N_2076,In_221,In_226);
nand U2077 (N_2077,In_35,In_714);
nor U2078 (N_2078,In_34,In_256);
xor U2079 (N_2079,In_730,In_383);
nor U2080 (N_2080,In_541,In_101);
and U2081 (N_2081,In_307,In_598);
xnor U2082 (N_2082,In_474,In_305);
or U2083 (N_2083,In_143,In_122);
nand U2084 (N_2084,In_360,In_664);
and U2085 (N_2085,In_511,In_372);
xnor U2086 (N_2086,In_331,In_197);
nand U2087 (N_2087,In_258,In_481);
or U2088 (N_2088,In_336,In_682);
or U2089 (N_2089,In_509,In_326);
nor U2090 (N_2090,In_137,In_233);
or U2091 (N_2091,In_192,In_725);
nor U2092 (N_2092,In_142,In_597);
nand U2093 (N_2093,In_702,In_26);
or U2094 (N_2094,In_643,In_735);
xnor U2095 (N_2095,In_91,In_230);
nand U2096 (N_2096,In_550,In_511);
xor U2097 (N_2097,In_195,In_675);
nor U2098 (N_2098,In_336,In_589);
nor U2099 (N_2099,In_231,In_171);
and U2100 (N_2100,In_100,In_490);
nor U2101 (N_2101,In_226,In_286);
xnor U2102 (N_2102,In_131,In_461);
nand U2103 (N_2103,In_119,In_291);
nor U2104 (N_2104,In_230,In_284);
and U2105 (N_2105,In_195,In_698);
and U2106 (N_2106,In_672,In_162);
or U2107 (N_2107,In_598,In_132);
nor U2108 (N_2108,In_591,In_286);
xor U2109 (N_2109,In_265,In_735);
nor U2110 (N_2110,In_12,In_475);
and U2111 (N_2111,In_254,In_11);
and U2112 (N_2112,In_687,In_398);
xnor U2113 (N_2113,In_637,In_153);
and U2114 (N_2114,In_666,In_663);
nor U2115 (N_2115,In_85,In_293);
nor U2116 (N_2116,In_685,In_628);
or U2117 (N_2117,In_542,In_345);
xor U2118 (N_2118,In_363,In_200);
and U2119 (N_2119,In_190,In_226);
nand U2120 (N_2120,In_47,In_503);
nand U2121 (N_2121,In_713,In_488);
nand U2122 (N_2122,In_155,In_454);
nand U2123 (N_2123,In_171,In_70);
xor U2124 (N_2124,In_460,In_374);
nand U2125 (N_2125,In_45,In_616);
xnor U2126 (N_2126,In_522,In_687);
nand U2127 (N_2127,In_250,In_202);
and U2128 (N_2128,In_531,In_565);
and U2129 (N_2129,In_102,In_146);
and U2130 (N_2130,In_183,In_79);
and U2131 (N_2131,In_346,In_330);
nor U2132 (N_2132,In_70,In_680);
and U2133 (N_2133,In_199,In_615);
nor U2134 (N_2134,In_241,In_145);
xor U2135 (N_2135,In_283,In_404);
or U2136 (N_2136,In_166,In_102);
and U2137 (N_2137,In_215,In_101);
or U2138 (N_2138,In_402,In_234);
xor U2139 (N_2139,In_138,In_544);
nor U2140 (N_2140,In_137,In_180);
and U2141 (N_2141,In_734,In_308);
xnor U2142 (N_2142,In_126,In_637);
or U2143 (N_2143,In_137,In_406);
nand U2144 (N_2144,In_70,In_48);
xor U2145 (N_2145,In_34,In_115);
xnor U2146 (N_2146,In_715,In_425);
and U2147 (N_2147,In_683,In_736);
or U2148 (N_2148,In_124,In_274);
nor U2149 (N_2149,In_523,In_310);
or U2150 (N_2150,In_221,In_644);
nand U2151 (N_2151,In_699,In_413);
and U2152 (N_2152,In_533,In_75);
nand U2153 (N_2153,In_331,In_95);
or U2154 (N_2154,In_452,In_125);
and U2155 (N_2155,In_653,In_427);
and U2156 (N_2156,In_15,In_485);
nor U2157 (N_2157,In_609,In_365);
nor U2158 (N_2158,In_77,In_549);
nor U2159 (N_2159,In_229,In_395);
xor U2160 (N_2160,In_360,In_249);
nand U2161 (N_2161,In_666,In_684);
xor U2162 (N_2162,In_96,In_656);
or U2163 (N_2163,In_597,In_174);
or U2164 (N_2164,In_548,In_199);
nor U2165 (N_2165,In_145,In_202);
xor U2166 (N_2166,In_479,In_485);
xnor U2167 (N_2167,In_740,In_693);
or U2168 (N_2168,In_562,In_662);
or U2169 (N_2169,In_266,In_381);
xnor U2170 (N_2170,In_180,In_535);
and U2171 (N_2171,In_337,In_268);
nand U2172 (N_2172,In_528,In_388);
and U2173 (N_2173,In_352,In_272);
nand U2174 (N_2174,In_454,In_424);
and U2175 (N_2175,In_676,In_28);
nor U2176 (N_2176,In_231,In_19);
nand U2177 (N_2177,In_726,In_574);
and U2178 (N_2178,In_638,In_697);
and U2179 (N_2179,In_438,In_637);
and U2180 (N_2180,In_360,In_613);
nor U2181 (N_2181,In_23,In_649);
nand U2182 (N_2182,In_255,In_43);
nand U2183 (N_2183,In_66,In_504);
and U2184 (N_2184,In_151,In_162);
nand U2185 (N_2185,In_29,In_123);
xor U2186 (N_2186,In_368,In_120);
nand U2187 (N_2187,In_653,In_125);
or U2188 (N_2188,In_344,In_655);
xnor U2189 (N_2189,In_680,In_491);
nor U2190 (N_2190,In_213,In_490);
or U2191 (N_2191,In_214,In_609);
nand U2192 (N_2192,In_133,In_180);
nand U2193 (N_2193,In_616,In_304);
nor U2194 (N_2194,In_423,In_698);
xnor U2195 (N_2195,In_172,In_575);
nor U2196 (N_2196,In_330,In_447);
nand U2197 (N_2197,In_232,In_229);
and U2198 (N_2198,In_298,In_535);
and U2199 (N_2199,In_292,In_28);
nand U2200 (N_2200,In_744,In_130);
nor U2201 (N_2201,In_562,In_622);
xor U2202 (N_2202,In_155,In_729);
or U2203 (N_2203,In_716,In_694);
nand U2204 (N_2204,In_658,In_561);
or U2205 (N_2205,In_251,In_658);
or U2206 (N_2206,In_384,In_485);
xor U2207 (N_2207,In_726,In_337);
or U2208 (N_2208,In_477,In_548);
nand U2209 (N_2209,In_43,In_164);
or U2210 (N_2210,In_156,In_30);
nor U2211 (N_2211,In_369,In_639);
xnor U2212 (N_2212,In_10,In_378);
nand U2213 (N_2213,In_717,In_254);
and U2214 (N_2214,In_317,In_441);
and U2215 (N_2215,In_365,In_579);
and U2216 (N_2216,In_573,In_13);
or U2217 (N_2217,In_267,In_404);
nand U2218 (N_2218,In_584,In_66);
xnor U2219 (N_2219,In_729,In_13);
nor U2220 (N_2220,In_633,In_36);
and U2221 (N_2221,In_454,In_67);
xor U2222 (N_2222,In_365,In_416);
or U2223 (N_2223,In_44,In_135);
and U2224 (N_2224,In_145,In_195);
nor U2225 (N_2225,In_498,In_554);
xor U2226 (N_2226,In_230,In_747);
xnor U2227 (N_2227,In_587,In_211);
and U2228 (N_2228,In_597,In_374);
or U2229 (N_2229,In_223,In_124);
nand U2230 (N_2230,In_526,In_325);
xor U2231 (N_2231,In_681,In_309);
or U2232 (N_2232,In_253,In_106);
xor U2233 (N_2233,In_271,In_261);
or U2234 (N_2234,In_412,In_476);
and U2235 (N_2235,In_588,In_140);
xnor U2236 (N_2236,In_361,In_635);
nor U2237 (N_2237,In_737,In_259);
xnor U2238 (N_2238,In_209,In_606);
nor U2239 (N_2239,In_14,In_473);
nor U2240 (N_2240,In_649,In_420);
and U2241 (N_2241,In_540,In_675);
nand U2242 (N_2242,In_524,In_96);
nand U2243 (N_2243,In_651,In_648);
and U2244 (N_2244,In_26,In_333);
xnor U2245 (N_2245,In_130,In_692);
or U2246 (N_2246,In_447,In_338);
and U2247 (N_2247,In_99,In_274);
and U2248 (N_2248,In_191,In_97);
xnor U2249 (N_2249,In_74,In_735);
xor U2250 (N_2250,In_229,In_62);
nor U2251 (N_2251,In_183,In_370);
nand U2252 (N_2252,In_444,In_245);
nand U2253 (N_2253,In_367,In_374);
xor U2254 (N_2254,In_704,In_614);
and U2255 (N_2255,In_538,In_700);
nor U2256 (N_2256,In_593,In_546);
nor U2257 (N_2257,In_466,In_613);
xnor U2258 (N_2258,In_106,In_388);
and U2259 (N_2259,In_272,In_449);
nor U2260 (N_2260,In_93,In_712);
xnor U2261 (N_2261,In_42,In_221);
nand U2262 (N_2262,In_472,In_743);
nand U2263 (N_2263,In_77,In_488);
and U2264 (N_2264,In_221,In_133);
nand U2265 (N_2265,In_587,In_499);
and U2266 (N_2266,In_349,In_729);
xnor U2267 (N_2267,In_412,In_74);
or U2268 (N_2268,In_612,In_199);
or U2269 (N_2269,In_97,In_386);
or U2270 (N_2270,In_51,In_206);
nand U2271 (N_2271,In_566,In_448);
nand U2272 (N_2272,In_93,In_728);
nand U2273 (N_2273,In_223,In_456);
or U2274 (N_2274,In_77,In_55);
and U2275 (N_2275,In_65,In_516);
nor U2276 (N_2276,In_386,In_329);
or U2277 (N_2277,In_164,In_243);
nand U2278 (N_2278,In_580,In_543);
and U2279 (N_2279,In_31,In_150);
or U2280 (N_2280,In_283,In_34);
or U2281 (N_2281,In_177,In_313);
and U2282 (N_2282,In_485,In_338);
nor U2283 (N_2283,In_318,In_715);
nand U2284 (N_2284,In_85,In_294);
nand U2285 (N_2285,In_367,In_78);
and U2286 (N_2286,In_338,In_636);
xor U2287 (N_2287,In_504,In_587);
or U2288 (N_2288,In_220,In_82);
xor U2289 (N_2289,In_168,In_90);
or U2290 (N_2290,In_399,In_586);
nor U2291 (N_2291,In_434,In_63);
nor U2292 (N_2292,In_404,In_70);
nand U2293 (N_2293,In_364,In_95);
or U2294 (N_2294,In_204,In_208);
nor U2295 (N_2295,In_220,In_393);
and U2296 (N_2296,In_251,In_242);
or U2297 (N_2297,In_673,In_651);
nand U2298 (N_2298,In_344,In_109);
nand U2299 (N_2299,In_269,In_228);
nand U2300 (N_2300,In_386,In_372);
nand U2301 (N_2301,In_234,In_651);
xor U2302 (N_2302,In_519,In_542);
nand U2303 (N_2303,In_530,In_35);
and U2304 (N_2304,In_708,In_557);
nand U2305 (N_2305,In_695,In_636);
xor U2306 (N_2306,In_676,In_368);
and U2307 (N_2307,In_713,In_9);
nand U2308 (N_2308,In_529,In_77);
xnor U2309 (N_2309,In_285,In_586);
nor U2310 (N_2310,In_522,In_71);
or U2311 (N_2311,In_117,In_664);
or U2312 (N_2312,In_299,In_193);
and U2313 (N_2313,In_624,In_579);
xor U2314 (N_2314,In_198,In_99);
xnor U2315 (N_2315,In_427,In_510);
xor U2316 (N_2316,In_428,In_718);
nand U2317 (N_2317,In_387,In_726);
xnor U2318 (N_2318,In_728,In_268);
nand U2319 (N_2319,In_420,In_171);
nand U2320 (N_2320,In_611,In_336);
nand U2321 (N_2321,In_239,In_567);
nor U2322 (N_2322,In_494,In_586);
and U2323 (N_2323,In_58,In_696);
nand U2324 (N_2324,In_689,In_459);
or U2325 (N_2325,In_450,In_485);
and U2326 (N_2326,In_572,In_414);
nand U2327 (N_2327,In_560,In_527);
and U2328 (N_2328,In_658,In_155);
or U2329 (N_2329,In_100,In_167);
or U2330 (N_2330,In_109,In_270);
xor U2331 (N_2331,In_736,In_98);
nor U2332 (N_2332,In_528,In_689);
nand U2333 (N_2333,In_345,In_398);
xor U2334 (N_2334,In_16,In_571);
and U2335 (N_2335,In_346,In_397);
nor U2336 (N_2336,In_97,In_666);
nor U2337 (N_2337,In_506,In_132);
nor U2338 (N_2338,In_624,In_212);
nand U2339 (N_2339,In_370,In_285);
xor U2340 (N_2340,In_651,In_661);
nand U2341 (N_2341,In_147,In_432);
nor U2342 (N_2342,In_367,In_537);
or U2343 (N_2343,In_470,In_706);
xnor U2344 (N_2344,In_79,In_425);
or U2345 (N_2345,In_390,In_385);
and U2346 (N_2346,In_142,In_652);
or U2347 (N_2347,In_358,In_124);
and U2348 (N_2348,In_517,In_44);
and U2349 (N_2349,In_98,In_418);
xnor U2350 (N_2350,In_271,In_641);
xnor U2351 (N_2351,In_539,In_217);
nand U2352 (N_2352,In_473,In_677);
nor U2353 (N_2353,In_153,In_404);
xnor U2354 (N_2354,In_137,In_105);
nand U2355 (N_2355,In_542,In_686);
nand U2356 (N_2356,In_385,In_369);
xnor U2357 (N_2357,In_575,In_127);
or U2358 (N_2358,In_233,In_3);
or U2359 (N_2359,In_523,In_443);
nor U2360 (N_2360,In_102,In_632);
xor U2361 (N_2361,In_101,In_36);
nand U2362 (N_2362,In_674,In_340);
or U2363 (N_2363,In_601,In_623);
nand U2364 (N_2364,In_439,In_84);
nor U2365 (N_2365,In_111,In_486);
nand U2366 (N_2366,In_607,In_333);
and U2367 (N_2367,In_501,In_723);
xnor U2368 (N_2368,In_308,In_111);
and U2369 (N_2369,In_148,In_488);
nor U2370 (N_2370,In_575,In_351);
nor U2371 (N_2371,In_363,In_291);
xnor U2372 (N_2372,In_174,In_31);
nand U2373 (N_2373,In_231,In_371);
and U2374 (N_2374,In_220,In_404);
xor U2375 (N_2375,In_713,In_400);
and U2376 (N_2376,In_438,In_414);
or U2377 (N_2377,In_264,In_16);
nand U2378 (N_2378,In_410,In_205);
nor U2379 (N_2379,In_528,In_414);
or U2380 (N_2380,In_640,In_653);
or U2381 (N_2381,In_206,In_614);
or U2382 (N_2382,In_82,In_739);
or U2383 (N_2383,In_371,In_135);
xnor U2384 (N_2384,In_315,In_218);
nor U2385 (N_2385,In_53,In_650);
nand U2386 (N_2386,In_43,In_355);
nand U2387 (N_2387,In_43,In_645);
and U2388 (N_2388,In_340,In_264);
nor U2389 (N_2389,In_250,In_712);
xnor U2390 (N_2390,In_621,In_308);
and U2391 (N_2391,In_273,In_735);
or U2392 (N_2392,In_87,In_268);
and U2393 (N_2393,In_80,In_747);
nor U2394 (N_2394,In_722,In_160);
and U2395 (N_2395,In_352,In_553);
xor U2396 (N_2396,In_78,In_475);
nand U2397 (N_2397,In_340,In_601);
or U2398 (N_2398,In_522,In_396);
or U2399 (N_2399,In_634,In_94);
nor U2400 (N_2400,In_674,In_325);
and U2401 (N_2401,In_383,In_469);
nand U2402 (N_2402,In_391,In_189);
nor U2403 (N_2403,In_696,In_621);
and U2404 (N_2404,In_418,In_417);
or U2405 (N_2405,In_519,In_500);
nor U2406 (N_2406,In_176,In_508);
nor U2407 (N_2407,In_454,In_258);
nand U2408 (N_2408,In_424,In_232);
or U2409 (N_2409,In_115,In_107);
xor U2410 (N_2410,In_501,In_95);
and U2411 (N_2411,In_224,In_670);
xnor U2412 (N_2412,In_290,In_329);
nand U2413 (N_2413,In_665,In_567);
and U2414 (N_2414,In_276,In_143);
and U2415 (N_2415,In_690,In_392);
and U2416 (N_2416,In_462,In_594);
nor U2417 (N_2417,In_183,In_286);
and U2418 (N_2418,In_344,In_11);
nand U2419 (N_2419,In_609,In_264);
nor U2420 (N_2420,In_535,In_317);
nor U2421 (N_2421,In_409,In_203);
or U2422 (N_2422,In_412,In_141);
nand U2423 (N_2423,In_479,In_593);
xnor U2424 (N_2424,In_91,In_241);
and U2425 (N_2425,In_461,In_39);
and U2426 (N_2426,In_666,In_71);
or U2427 (N_2427,In_382,In_129);
or U2428 (N_2428,In_631,In_406);
nor U2429 (N_2429,In_285,In_603);
and U2430 (N_2430,In_740,In_354);
and U2431 (N_2431,In_552,In_66);
nor U2432 (N_2432,In_419,In_397);
xor U2433 (N_2433,In_401,In_560);
or U2434 (N_2434,In_387,In_524);
or U2435 (N_2435,In_666,In_166);
or U2436 (N_2436,In_118,In_248);
xnor U2437 (N_2437,In_400,In_328);
and U2438 (N_2438,In_240,In_704);
and U2439 (N_2439,In_399,In_357);
and U2440 (N_2440,In_249,In_461);
xnor U2441 (N_2441,In_715,In_550);
xor U2442 (N_2442,In_76,In_487);
nor U2443 (N_2443,In_476,In_293);
nand U2444 (N_2444,In_296,In_117);
nor U2445 (N_2445,In_210,In_244);
or U2446 (N_2446,In_601,In_510);
or U2447 (N_2447,In_468,In_588);
xnor U2448 (N_2448,In_32,In_48);
nand U2449 (N_2449,In_389,In_468);
or U2450 (N_2450,In_336,In_92);
or U2451 (N_2451,In_157,In_274);
or U2452 (N_2452,In_680,In_139);
nand U2453 (N_2453,In_262,In_475);
or U2454 (N_2454,In_554,In_365);
or U2455 (N_2455,In_276,In_37);
nand U2456 (N_2456,In_615,In_509);
and U2457 (N_2457,In_331,In_323);
or U2458 (N_2458,In_524,In_371);
or U2459 (N_2459,In_208,In_411);
and U2460 (N_2460,In_280,In_210);
or U2461 (N_2461,In_521,In_90);
and U2462 (N_2462,In_644,In_224);
nor U2463 (N_2463,In_54,In_61);
or U2464 (N_2464,In_467,In_137);
nor U2465 (N_2465,In_699,In_603);
xor U2466 (N_2466,In_602,In_265);
nor U2467 (N_2467,In_421,In_427);
or U2468 (N_2468,In_665,In_424);
or U2469 (N_2469,In_699,In_90);
nand U2470 (N_2470,In_368,In_274);
nor U2471 (N_2471,In_89,In_13);
nor U2472 (N_2472,In_83,In_212);
or U2473 (N_2473,In_677,In_492);
nor U2474 (N_2474,In_164,In_516);
xor U2475 (N_2475,In_379,In_723);
and U2476 (N_2476,In_122,In_631);
nor U2477 (N_2477,In_643,In_331);
xor U2478 (N_2478,In_524,In_15);
nor U2479 (N_2479,In_305,In_51);
and U2480 (N_2480,In_261,In_54);
and U2481 (N_2481,In_728,In_500);
xnor U2482 (N_2482,In_548,In_163);
nand U2483 (N_2483,In_391,In_209);
and U2484 (N_2484,In_85,In_736);
xor U2485 (N_2485,In_215,In_436);
nand U2486 (N_2486,In_42,In_281);
and U2487 (N_2487,In_660,In_48);
and U2488 (N_2488,In_80,In_521);
xnor U2489 (N_2489,In_224,In_350);
or U2490 (N_2490,In_338,In_479);
and U2491 (N_2491,In_382,In_516);
nor U2492 (N_2492,In_219,In_690);
nand U2493 (N_2493,In_673,In_693);
xnor U2494 (N_2494,In_326,In_127);
nand U2495 (N_2495,In_235,In_557);
and U2496 (N_2496,In_737,In_155);
nand U2497 (N_2497,In_333,In_596);
or U2498 (N_2498,In_403,In_616);
and U2499 (N_2499,In_623,In_460);
or U2500 (N_2500,N_2261,N_1243);
nand U2501 (N_2501,N_2462,N_2352);
nor U2502 (N_2502,N_1754,N_842);
nand U2503 (N_2503,N_557,N_1156);
and U2504 (N_2504,N_787,N_1647);
and U2505 (N_2505,N_2019,N_896);
xnor U2506 (N_2506,N_1929,N_1442);
or U2507 (N_2507,N_948,N_962);
nand U2508 (N_2508,N_2309,N_1963);
nand U2509 (N_2509,N_2439,N_2395);
xnor U2510 (N_2510,N_281,N_1446);
xor U2511 (N_2511,N_2018,N_1848);
and U2512 (N_2512,N_2414,N_1146);
or U2513 (N_2513,N_1276,N_2407);
nand U2514 (N_2514,N_180,N_80);
nor U2515 (N_2515,N_21,N_1436);
and U2516 (N_2516,N_701,N_171);
xor U2517 (N_2517,N_1427,N_2228);
xnor U2518 (N_2518,N_1939,N_2481);
or U2519 (N_2519,N_1447,N_1942);
or U2520 (N_2520,N_705,N_1624);
and U2521 (N_2521,N_381,N_1496);
or U2522 (N_2522,N_1542,N_1905);
nand U2523 (N_2523,N_455,N_1172);
or U2524 (N_2524,N_2037,N_1532);
and U2525 (N_2525,N_1482,N_114);
xnor U2526 (N_2526,N_497,N_472);
nand U2527 (N_2527,N_432,N_1777);
and U2528 (N_2528,N_920,N_897);
or U2529 (N_2529,N_1057,N_24);
and U2530 (N_2530,N_521,N_1060);
and U2531 (N_2531,N_260,N_270);
or U2532 (N_2532,N_887,N_1852);
nor U2533 (N_2533,N_591,N_2343);
nor U2534 (N_2534,N_1823,N_1577);
and U2535 (N_2535,N_786,N_1541);
and U2536 (N_2536,N_1299,N_1165);
nand U2537 (N_2537,N_318,N_1519);
nor U2538 (N_2538,N_211,N_1045);
nand U2539 (N_2539,N_879,N_2301);
nand U2540 (N_2540,N_1055,N_1552);
or U2541 (N_2541,N_1562,N_141);
and U2542 (N_2542,N_2255,N_1538);
and U2543 (N_2543,N_2123,N_2154);
nor U2544 (N_2544,N_837,N_950);
and U2545 (N_2545,N_2480,N_253);
xnor U2546 (N_2546,N_353,N_662);
and U2547 (N_2547,N_1404,N_95);
or U2548 (N_2548,N_93,N_1326);
nor U2549 (N_2549,N_1162,N_963);
or U2550 (N_2550,N_1341,N_1293);
or U2551 (N_2551,N_1031,N_1451);
nor U2552 (N_2552,N_2162,N_2431);
xnor U2553 (N_2553,N_1066,N_101);
nor U2554 (N_2554,N_2077,N_1033);
xnor U2555 (N_2555,N_1186,N_1915);
and U2556 (N_2556,N_1775,N_1888);
and U2557 (N_2557,N_1679,N_1516);
and U2558 (N_2558,N_156,N_2119);
or U2559 (N_2559,N_397,N_998);
or U2560 (N_2560,N_1312,N_2111);
and U2561 (N_2561,N_1381,N_133);
nor U2562 (N_2562,N_53,N_732);
nand U2563 (N_2563,N_1484,N_1564);
nand U2564 (N_2564,N_2105,N_1596);
or U2565 (N_2565,N_359,N_2323);
nand U2566 (N_2566,N_1599,N_172);
and U2567 (N_2567,N_2155,N_2279);
nand U2568 (N_2568,N_1999,N_2339);
nand U2569 (N_2569,N_1643,N_2282);
xnor U2570 (N_2570,N_323,N_250);
nor U2571 (N_2571,N_45,N_2177);
or U2572 (N_2572,N_127,N_2398);
xnor U2573 (N_2573,N_1798,N_537);
and U2574 (N_2574,N_618,N_338);
xor U2575 (N_2575,N_2060,N_1937);
xnor U2576 (N_2576,N_2266,N_1614);
xnor U2577 (N_2577,N_326,N_2463);
nor U2578 (N_2578,N_1474,N_996);
or U2579 (N_2579,N_321,N_1870);
and U2580 (N_2580,N_765,N_988);
xor U2581 (N_2581,N_2044,N_2422);
xnor U2582 (N_2582,N_2058,N_984);
xor U2583 (N_2583,N_566,N_1159);
nand U2584 (N_2584,N_240,N_1169);
xor U2585 (N_2585,N_574,N_1131);
xor U2586 (N_2586,N_1800,N_1865);
nand U2587 (N_2587,N_116,N_367);
or U2588 (N_2588,N_1002,N_873);
and U2589 (N_2589,N_1602,N_1583);
xor U2590 (N_2590,N_246,N_1531);
xor U2591 (N_2591,N_619,N_2106);
xnor U2592 (N_2592,N_872,N_1278);
nand U2593 (N_2593,N_1654,N_1214);
or U2594 (N_2594,N_2373,N_483);
and U2595 (N_2595,N_1473,N_304);
and U2596 (N_2596,N_2391,N_1476);
nand U2597 (N_2597,N_92,N_1697);
and U2598 (N_2598,N_1553,N_1986);
and U2599 (N_2599,N_360,N_1137);
xnor U2600 (N_2600,N_334,N_2171);
xor U2601 (N_2601,N_598,N_333);
nor U2602 (N_2602,N_1648,N_1361);
nor U2603 (N_2603,N_1626,N_188);
xor U2604 (N_2604,N_76,N_498);
nand U2605 (N_2605,N_1843,N_901);
and U2606 (N_2606,N_623,N_265);
xor U2607 (N_2607,N_1544,N_1829);
or U2608 (N_2608,N_1700,N_1093);
xnor U2609 (N_2609,N_1920,N_2188);
nor U2610 (N_2610,N_1916,N_974);
and U2611 (N_2611,N_1816,N_1193);
or U2612 (N_2612,N_684,N_1724);
and U2613 (N_2613,N_2167,N_505);
or U2614 (N_2614,N_2420,N_1734);
or U2615 (N_2615,N_2361,N_1091);
xnor U2616 (N_2616,N_392,N_1160);
nand U2617 (N_2617,N_2107,N_2499);
nor U2618 (N_2618,N_183,N_1272);
nand U2619 (N_2619,N_1011,N_2483);
or U2620 (N_2620,N_1575,N_1120);
or U2621 (N_2621,N_534,N_2307);
nand U2622 (N_2622,N_2363,N_1669);
xnor U2623 (N_2623,N_860,N_1197);
and U2624 (N_2624,N_94,N_2131);
nand U2625 (N_2625,N_47,N_1994);
nor U2626 (N_2626,N_1522,N_1743);
and U2627 (N_2627,N_324,N_1855);
or U2628 (N_2628,N_1938,N_1713);
nand U2629 (N_2629,N_1880,N_339);
or U2630 (N_2630,N_926,N_1667);
or U2631 (N_2631,N_630,N_710);
and U2632 (N_2632,N_332,N_1658);
or U2633 (N_2633,N_67,N_1535);
xnor U2634 (N_2634,N_1048,N_344);
xnor U2635 (N_2635,N_655,N_1527);
and U2636 (N_2636,N_1729,N_2292);
or U2637 (N_2637,N_160,N_1611);
nor U2638 (N_2638,N_2023,N_1895);
nand U2639 (N_2639,N_632,N_1857);
and U2640 (N_2640,N_1149,N_2194);
xnor U2641 (N_2641,N_1995,N_1681);
nor U2642 (N_2642,N_638,N_1489);
and U2643 (N_2643,N_2072,N_1933);
xnor U2644 (N_2644,N_1357,N_2078);
or U2645 (N_2645,N_2114,N_2425);
nor U2646 (N_2646,N_2325,N_2400);
nor U2647 (N_2647,N_1500,N_2467);
or U2648 (N_2648,N_1101,N_227);
nor U2649 (N_2649,N_1808,N_991);
nor U2650 (N_2650,N_2021,N_401);
and U2651 (N_2651,N_1116,N_1683);
and U2652 (N_2652,N_2328,N_199);
xor U2653 (N_2653,N_1819,N_910);
xor U2654 (N_2654,N_261,N_1374);
or U2655 (N_2655,N_192,N_1042);
or U2656 (N_2656,N_1108,N_1504);
xnor U2657 (N_2657,N_2182,N_1270);
nand U2658 (N_2658,N_1715,N_1179);
nand U2659 (N_2659,N_1050,N_1130);
and U2660 (N_2660,N_420,N_1369);
and U2661 (N_2661,N_118,N_1439);
xnor U2662 (N_2662,N_783,N_82);
nor U2663 (N_2663,N_393,N_1891);
or U2664 (N_2664,N_124,N_2032);
nand U2665 (N_2665,N_558,N_1229);
nor U2666 (N_2666,N_486,N_1764);
xnor U2667 (N_2667,N_206,N_162);
nand U2668 (N_2668,N_2364,N_1690);
and U2669 (N_2669,N_1641,N_1712);
or U2670 (N_2670,N_1782,N_840);
or U2671 (N_2671,N_2087,N_2412);
or U2672 (N_2672,N_689,N_2306);
and U2673 (N_2673,N_760,N_2020);
nand U2674 (N_2674,N_602,N_687);
xnor U2675 (N_2675,N_1265,N_919);
nand U2676 (N_2676,N_1806,N_1356);
and U2677 (N_2677,N_1392,N_1714);
nand U2678 (N_2678,N_947,N_310);
and U2679 (N_2679,N_77,N_891);
nand U2680 (N_2680,N_789,N_63);
nand U2681 (N_2681,N_888,N_1271);
nand U2682 (N_2682,N_1420,N_1492);
nand U2683 (N_2683,N_1046,N_2247);
nand U2684 (N_2684,N_2369,N_805);
xor U2685 (N_2685,N_194,N_2362);
nor U2686 (N_2686,N_201,N_1904);
nor U2687 (N_2687,N_26,N_1608);
xnor U2688 (N_2688,N_1597,N_165);
and U2689 (N_2689,N_489,N_563);
nor U2690 (N_2690,N_2444,N_316);
nand U2691 (N_2691,N_2490,N_2047);
or U2692 (N_2692,N_106,N_286);
nor U2693 (N_2693,N_2426,N_1878);
nor U2694 (N_2694,N_1603,N_935);
or U2695 (N_2695,N_992,N_1205);
xor U2696 (N_2696,N_354,N_1298);
xor U2697 (N_2697,N_257,N_113);
nor U2698 (N_2698,N_774,N_166);
or U2699 (N_2699,N_654,N_622);
and U2700 (N_2700,N_337,N_1340);
xnor U2701 (N_2701,N_1642,N_1805);
or U2702 (N_2702,N_1956,N_535);
nor U2703 (N_2703,N_1784,N_2101);
nand U2704 (N_2704,N_288,N_1029);
nor U2705 (N_2705,N_578,N_2216);
nand U2706 (N_2706,N_1794,N_627);
or U2707 (N_2707,N_880,N_362);
xnor U2708 (N_2708,N_461,N_377);
xor U2709 (N_2709,N_565,N_676);
nand U2710 (N_2710,N_918,N_749);
nand U2711 (N_2711,N_2122,N_1256);
xnor U2712 (N_2712,N_1483,N_494);
and U2713 (N_2713,N_303,N_617);
or U2714 (N_2714,N_23,N_990);
or U2715 (N_2715,N_2433,N_149);
and U2716 (N_2716,N_834,N_1721);
xnor U2717 (N_2717,N_1136,N_1232);
nor U2718 (N_2718,N_709,N_959);
and U2719 (N_2719,N_2298,N_282);
xor U2720 (N_2720,N_13,N_2001);
or U2721 (N_2721,N_1285,N_1145);
nand U2722 (N_2722,N_358,N_1978);
xor U2723 (N_2723,N_1217,N_2148);
or U2724 (N_2724,N_1581,N_981);
and U2725 (N_2725,N_331,N_1830);
nand U2726 (N_2726,N_798,N_641);
and U2727 (N_2727,N_651,N_823);
xnor U2728 (N_2728,N_1004,N_999);
xnor U2729 (N_2729,N_1788,N_1637);
nand U2730 (N_2730,N_1772,N_661);
or U2731 (N_2731,N_683,N_1871);
nand U2732 (N_2732,N_1399,N_2272);
nor U2733 (N_2733,N_755,N_84);
nand U2734 (N_2734,N_479,N_1412);
xor U2735 (N_2735,N_1490,N_75);
or U2736 (N_2736,N_852,N_2442);
and U2737 (N_2737,N_1242,N_464);
nor U2738 (N_2738,N_1443,N_625);
nand U2739 (N_2739,N_2384,N_145);
xnor U2740 (N_2740,N_1558,N_1152);
nor U2741 (N_2741,N_148,N_2168);
xnor U2742 (N_2742,N_2176,N_568);
nor U2743 (N_2743,N_422,N_186);
or U2744 (N_2744,N_1491,N_876);
or U2745 (N_2745,N_463,N_1409);
xnor U2746 (N_2746,N_439,N_838);
nor U2747 (N_2747,N_175,N_821);
nand U2748 (N_2748,N_1216,N_1150);
nor U2749 (N_2749,N_68,N_2461);
nand U2750 (N_2750,N_1335,N_645);
or U2751 (N_2751,N_1716,N_1090);
xor U2752 (N_2752,N_913,N_752);
or U2753 (N_2753,N_2121,N_154);
or U2754 (N_2754,N_2102,N_226);
and U2755 (N_2755,N_2326,N_1345);
nor U2756 (N_2756,N_777,N_1418);
and U2757 (N_2757,N_1249,N_1016);
nand U2758 (N_2758,N_273,N_2006);
or U2759 (N_2759,N_2479,N_1115);
or U2760 (N_2760,N_225,N_2127);
nor U2761 (N_2761,N_674,N_1215);
nor U2762 (N_2762,N_395,N_958);
nand U2763 (N_2763,N_1006,N_2220);
or U2764 (N_2764,N_1651,N_835);
xor U2765 (N_2765,N_1177,N_1428);
nand U2766 (N_2766,N_2221,N_605);
nand U2767 (N_2767,N_2241,N_878);
nand U2768 (N_2768,N_874,N_419);
and U2769 (N_2769,N_697,N_2181);
nor U2770 (N_2770,N_279,N_696);
nor U2771 (N_2771,N_877,N_524);
nor U2772 (N_2772,N_1157,N_375);
nor U2773 (N_2773,N_445,N_886);
and U2774 (N_2774,N_849,N_1653);
and U2775 (N_2775,N_2297,N_2475);
and U2776 (N_2776,N_1495,N_1854);
nor U2777 (N_2777,N_1087,N_1148);
and U2778 (N_2778,N_1096,N_551);
nand U2779 (N_2779,N_1924,N_839);
xor U2780 (N_2780,N_668,N_658);
xnor U2781 (N_2781,N_2113,N_1897);
nor U2782 (N_2782,N_1606,N_1013);
nor U2783 (N_2783,N_2271,N_1918);
or U2784 (N_2784,N_809,N_1837);
nor U2785 (N_2785,N_647,N_613);
nor U2786 (N_2786,N_1189,N_234);
xnor U2787 (N_2787,N_933,N_64);
and U2788 (N_2788,N_1459,N_1590);
xnor U2789 (N_2789,N_1621,N_1138);
nand U2790 (N_2790,N_1831,N_1199);
xor U2791 (N_2791,N_1509,N_2287);
nor U2792 (N_2792,N_1435,N_549);
or U2793 (N_2793,N_1364,N_2149);
and U2794 (N_2794,N_1314,N_1824);
and U2795 (N_2795,N_305,N_2076);
xnor U2796 (N_2796,N_1687,N_2453);
xor U2797 (N_2797,N_1258,N_2342);
xor U2798 (N_2798,N_1524,N_2160);
nor U2799 (N_2799,N_2109,N_1325);
xor U2800 (N_2800,N_1635,N_1799);
nor U2801 (N_2801,N_2137,N_586);
nand U2802 (N_2802,N_1846,N_2039);
or U2803 (N_2803,N_2002,N_1927);
nand U2804 (N_2804,N_1455,N_2207);
and U2805 (N_2805,N_1505,N_1228);
xnor U2806 (N_2806,N_889,N_564);
nor U2807 (N_2807,N_681,N_2175);
nand U2808 (N_2808,N_754,N_2252);
xnor U2809 (N_2809,N_856,N_2022);
nor U2810 (N_2810,N_1103,N_590);
and U2811 (N_2811,N_184,N_2374);
and U2812 (N_2812,N_1555,N_1140);
nor U2813 (N_2813,N_979,N_2385);
nor U2814 (N_2814,N_488,N_1998);
or U2815 (N_2815,N_1753,N_802);
nand U2816 (N_2816,N_1955,N_155);
nand U2817 (N_2817,N_2450,N_2334);
nor U2818 (N_2818,N_425,N_1561);
or U2819 (N_2819,N_693,N_207);
or U2820 (N_2820,N_1945,N_2126);
nor U2821 (N_2821,N_2212,N_473);
and U2822 (N_2822,N_1849,N_620);
nor U2823 (N_2823,N_1885,N_567);
and U2824 (N_2824,N_1224,N_579);
xor U2825 (N_2825,N_932,N_431);
xor U2826 (N_2826,N_1853,N_546);
xor U2827 (N_2827,N_851,N_1142);
xnor U2828 (N_2828,N_1833,N_921);
or U2829 (N_2829,N_807,N_1385);
and U2830 (N_2830,N_1235,N_1537);
nand U2831 (N_2831,N_105,N_1809);
xor U2832 (N_2832,N_1617,N_2143);
and U2833 (N_2833,N_2213,N_1370);
xor U2834 (N_2834,N_2435,N_2203);
and U2835 (N_2835,N_2319,N_1909);
or U2836 (N_2836,N_673,N_664);
and U2837 (N_2837,N_767,N_1291);
and U2838 (N_2838,N_929,N_892);
nand U2839 (N_2839,N_648,N_995);
nand U2840 (N_2840,N_2215,N_571);
xnor U2841 (N_2841,N_301,N_1457);
nor U2842 (N_2842,N_499,N_2239);
or U2843 (N_2843,N_437,N_850);
or U2844 (N_2844,N_728,N_125);
nor U2845 (N_2845,N_1841,N_386);
nor U2846 (N_2846,N_1386,N_2132);
xnor U2847 (N_2847,N_2100,N_548);
nor U2848 (N_2848,N_1458,N_509);
or U2849 (N_2849,N_1979,N_2231);
and U2850 (N_2850,N_139,N_468);
or U2851 (N_2851,N_1468,N_1722);
or U2852 (N_2852,N_2392,N_639);
and U2853 (N_2853,N_624,N_2495);
xor U2854 (N_2854,N_1882,N_1812);
nand U2855 (N_2855,N_1631,N_955);
and U2856 (N_2856,N_290,N_30);
and U2857 (N_2857,N_2432,N_161);
and U2858 (N_2858,N_2464,N_720);
nand U2859 (N_2859,N_1273,N_1925);
nor U2860 (N_2860,N_2192,N_1430);
xnor U2861 (N_2861,N_1960,N_978);
nor U2862 (N_2862,N_2178,N_511);
and U2863 (N_2863,N_1184,N_956);
nand U2864 (N_2864,N_2250,N_39);
nor U2865 (N_2865,N_2232,N_1811);
xor U2866 (N_2866,N_1665,N_738);
nor U2867 (N_2867,N_2049,N_2075);
nor U2868 (N_2868,N_1350,N_1294);
xnor U2869 (N_2869,N_1322,N_440);
or U2870 (N_2870,N_2059,N_297);
or U2871 (N_2871,N_1040,N_1230);
nand U2872 (N_2872,N_50,N_715);
and U2873 (N_2873,N_819,N_703);
and U2874 (N_2874,N_309,N_1164);
or U2875 (N_2875,N_2270,N_203);
nor U2876 (N_2876,N_424,N_435);
nor U2877 (N_2877,N_1233,N_717);
xnor U2878 (N_2878,N_2024,N_1887);
or U2879 (N_2879,N_1192,N_670);
and U2880 (N_2880,N_1203,N_1699);
or U2881 (N_2881,N_1952,N_523);
nor U2882 (N_2882,N_1467,N_516);
or U2883 (N_2883,N_320,N_1431);
xor U2884 (N_2884,N_1737,N_1573);
xor U2885 (N_2885,N_233,N_2269);
and U2886 (N_2886,N_770,N_2159);
or U2887 (N_2887,N_912,N_2088);
xor U2888 (N_2888,N_1124,N_2291);
nor U2889 (N_2889,N_1081,N_1349);
nand U2890 (N_2890,N_469,N_542);
and U2891 (N_2891,N_430,N_1062);
xor U2892 (N_2892,N_1604,N_806);
xor U2893 (N_2893,N_1334,N_1413);
nor U2894 (N_2894,N_1208,N_2230);
xor U2895 (N_2895,N_408,N_1676);
xnor U2896 (N_2896,N_923,N_649);
or U2897 (N_2897,N_351,N_1674);
and U2898 (N_2898,N_1950,N_1084);
nand U2899 (N_2899,N_1645,N_2393);
or U2900 (N_2900,N_1280,N_607);
nand U2901 (N_2901,N_2313,N_1423);
xor U2902 (N_2902,N_501,N_1989);
nand U2903 (N_2903,N_1861,N_2187);
or U2904 (N_2904,N_742,N_724);
xor U2905 (N_2905,N_1311,N_1983);
nand U2906 (N_2906,N_131,N_1038);
nor U2907 (N_2907,N_376,N_828);
nand U2908 (N_2908,N_2267,N_2062);
nor U2909 (N_2909,N_708,N_447);
and U2910 (N_2910,N_1826,N_731);
or U2911 (N_2911,N_2492,N_808);
or U2912 (N_2912,N_1903,N_1434);
and U2913 (N_2913,N_899,N_1691);
xor U2914 (N_2914,N_626,N_88);
xnor U2915 (N_2915,N_1035,N_2090);
nor U2916 (N_2916,N_1976,N_1814);
or U2917 (N_2917,N_1736,N_223);
or U2918 (N_2918,N_1570,N_692);
or U2919 (N_2919,N_1039,N_580);
and U2920 (N_2920,N_1372,N_1477);
nor U2921 (N_2921,N_1007,N_2346);
xnor U2922 (N_2922,N_5,N_2413);
or U2923 (N_2923,N_83,N_1874);
or U2924 (N_2924,N_477,N_2086);
xnor U2925 (N_2925,N_138,N_1211);
or U2926 (N_2926,N_952,N_1320);
nor U2927 (N_2927,N_1946,N_1968);
xnor U2928 (N_2928,N_1127,N_1747);
xor U2929 (N_2929,N_2429,N_927);
or U2930 (N_2930,N_1987,N_307);
xor U2931 (N_2931,N_1308,N_1321);
or U2932 (N_2932,N_1533,N_2330);
or U2933 (N_2933,N_1622,N_1748);
and U2934 (N_2934,N_2015,N_797);
nand U2935 (N_2935,N_163,N_1615);
nand U2936 (N_2936,N_1685,N_986);
xor U2937 (N_2937,N_1770,N_788);
nor U2938 (N_2938,N_467,N_1718);
nor U2939 (N_2939,N_762,N_1940);
nand U2940 (N_2940,N_2173,N_1092);
xnor U2941 (N_2941,N_444,N_1020);
nand U2942 (N_2942,N_216,N_729);
or U2943 (N_2943,N_1969,N_1132);
nor U2944 (N_2944,N_698,N_1445);
nand U2945 (N_2945,N_1569,N_1371);
and U2946 (N_2946,N_476,N_1290);
or U2947 (N_2947,N_2205,N_1037);
or U2948 (N_2948,N_1008,N_2304);
nor U2949 (N_2949,N_1796,N_249);
or U2950 (N_2950,N_2445,N_2094);
nand U2951 (N_2951,N_41,N_86);
xor U2952 (N_2952,N_938,N_2063);
and U2953 (N_2953,N_1082,N_1450);
nand U2954 (N_2954,N_1212,N_176);
nand U2955 (N_2955,N_750,N_16);
or U2956 (N_2956,N_242,N_2417);
nor U2957 (N_2957,N_1953,N_1910);
nor U2958 (N_2958,N_2224,N_2390);
or U2959 (N_2959,N_1070,N_383);
xor U2960 (N_2960,N_1400,N_1954);
nand U2961 (N_2961,N_863,N_1227);
nand U2962 (N_2962,N_1773,N_1498);
and U2963 (N_2963,N_2074,N_771);
nor U2964 (N_2964,N_903,N_1073);
xor U2965 (N_2965,N_702,N_1992);
nand U2966 (N_2966,N_1281,N_928);
nor U2967 (N_2967,N_2071,N_1429);
nor U2968 (N_2968,N_434,N_2321);
nor U2969 (N_2969,N_1822,N_480);
or U2970 (N_2970,N_1323,N_1478);
and U2971 (N_2971,N_484,N_256);
xor U2972 (N_2972,N_1348,N_1262);
nand U2973 (N_2973,N_1644,N_650);
and U2974 (N_2974,N_1973,N_1664);
and U2975 (N_2975,N_2386,N_881);
nand U2976 (N_2976,N_209,N_1710);
xnor U2977 (N_2977,N_2332,N_983);
nand U2978 (N_2978,N_855,N_1886);
xnor U2979 (N_2979,N_104,N_2112);
nor U2980 (N_2980,N_2163,N_1543);
xor U2981 (N_2981,N_2276,N_2223);
or U2982 (N_2982,N_785,N_1288);
xnor U2983 (N_2983,N_1497,N_1639);
and U2984 (N_2984,N_109,N_2091);
or U2985 (N_2985,N_764,N_1607);
nor U2986 (N_2986,N_941,N_2283);
and U2987 (N_2987,N_2337,N_384);
xnor U2988 (N_2988,N_757,N_2441);
or U2989 (N_2989,N_1847,N_1448);
or U2990 (N_2990,N_1425,N_1684);
nand U2991 (N_2991,N_1894,N_103);
nor U2992 (N_2992,N_2310,N_2338);
and U2993 (N_2993,N_1387,N_796);
nor U2994 (N_2994,N_1098,N_1000);
xor U2995 (N_2995,N_2195,N_2070);
xnor U2996 (N_2996,N_1579,N_677);
and U2997 (N_2997,N_1287,N_328);
or U2998 (N_2998,N_2489,N_1802);
and U2999 (N_2999,N_545,N_1390);
nor U3000 (N_3000,N_740,N_1723);
and U3001 (N_3001,N_1206,N_1275);
or U3002 (N_3002,N_417,N_429);
and U3003 (N_3003,N_1842,N_1209);
and U3004 (N_3004,N_1656,N_562);
or U3005 (N_3005,N_1594,N_1362);
and U3006 (N_3006,N_1128,N_1768);
and U3007 (N_3007,N_500,N_400);
xnor U3008 (N_3008,N_1785,N_1742);
xnor U3009 (N_3009,N_688,N_1110);
nand U3010 (N_3010,N_115,N_1122);
or U3011 (N_3011,N_252,N_2093);
nor U3012 (N_3012,N_2082,N_937);
nor U3013 (N_3013,N_278,N_1240);
or U3014 (N_3014,N_458,N_1510);
or U3015 (N_3015,N_1449,N_853);
or U3016 (N_3016,N_2057,N_1572);
xnor U3017 (N_3017,N_1257,N_1352);
and U3018 (N_3018,N_866,N_2424);
xnor U3019 (N_3019,N_2166,N_1545);
xor U3020 (N_3020,N_119,N_1052);
and U3021 (N_3021,N_1997,N_2084);
nand U3022 (N_3022,N_123,N_1763);
nand U3023 (N_3023,N_723,N_215);
xor U3024 (N_3024,N_1499,N_1274);
nor U3025 (N_3025,N_1009,N_845);
xnor U3026 (N_3026,N_1163,N_1521);
and U3027 (N_3027,N_1301,N_1540);
nor U3028 (N_3028,N_825,N_1706);
xor U3029 (N_3029,N_2030,N_2116);
and U3030 (N_3030,N_218,N_530);
or U3031 (N_3031,N_369,N_61);
xnor U3032 (N_3032,N_2183,N_1787);
or U3033 (N_3033,N_945,N_1760);
or U3034 (N_3034,N_766,N_1752);
xor U3035 (N_3035,N_128,N_2157);
nor U3036 (N_3036,N_826,N_365);
and U3037 (N_3037,N_1061,N_2144);
xnor U3038 (N_3038,N_1027,N_1917);
nand U3039 (N_3039,N_2219,N_142);
nand U3040 (N_3040,N_2238,N_1375);
nand U3041 (N_3041,N_504,N_2055);
xor U3042 (N_3042,N_481,N_1661);
and U3043 (N_3043,N_2488,N_258);
or U3044 (N_3044,N_2141,N_1844);
nor U3045 (N_3045,N_2294,N_448);
xor U3046 (N_3046,N_1379,N_269);
nand U3047 (N_3047,N_725,N_1633);
or U3048 (N_3048,N_2317,N_325);
nand U3049 (N_3049,N_2134,N_372);
and U3050 (N_3050,N_653,N_315);
and U3051 (N_3051,N_1548,N_1958);
nor U3052 (N_3052,N_769,N_1266);
nand U3053 (N_3053,N_943,N_656);
nand U3054 (N_3054,N_18,N_1072);
nor U3055 (N_3055,N_2067,N_1306);
and U3056 (N_3056,N_1158,N_583);
and U3057 (N_3057,N_748,N_1902);
or U3058 (N_3058,N_1102,N_283);
and U3059 (N_3059,N_657,N_1133);
or U3060 (N_3060,N_1557,N_87);
and U3061 (N_3061,N_1619,N_97);
and U3062 (N_3062,N_42,N_1175);
xnor U3063 (N_3063,N_930,N_713);
nand U3064 (N_3064,N_1180,N_413);
or U3065 (N_3065,N_1720,N_2303);
nor U3066 (N_3066,N_2460,N_1432);
nor U3067 (N_3067,N_843,N_298);
or U3068 (N_3068,N_2341,N_2026);
or U3069 (N_3069,N_554,N_1139);
nor U3070 (N_3070,N_1017,N_2246);
xnor U3071 (N_3071,N_1289,N_2434);
nor U3072 (N_3072,N_989,N_1109);
nor U3073 (N_3073,N_2482,N_1239);
xnor U3074 (N_3074,N_960,N_540);
or U3075 (N_3075,N_975,N_190);
nor U3076 (N_3076,N_239,N_517);
xnor U3077 (N_3077,N_707,N_2428);
or U3078 (N_3078,N_669,N_861);
xnor U3079 (N_3079,N_621,N_1305);
or U3080 (N_3080,N_1058,N_859);
and U3081 (N_3081,N_174,N_1324);
nand U3082 (N_3082,N_2371,N_198);
or U3083 (N_3083,N_1354,N_1793);
nor U3084 (N_3084,N_870,N_1892);
and U3085 (N_3085,N_1901,N_603);
and U3086 (N_3086,N_1328,N_966);
xnor U3087 (N_3087,N_415,N_411);
and U3088 (N_3088,N_2358,N_2351);
xnor U3089 (N_3089,N_2050,N_1076);
and U3090 (N_3090,N_308,N_1221);
and U3091 (N_3091,N_1393,N_405);
and U3092 (N_3092,N_1185,N_665);
nor U3093 (N_3093,N_780,N_716);
xor U3094 (N_3094,N_736,N_2401);
and U3095 (N_3095,N_555,N_2472);
or U3096 (N_3096,N_1820,N_152);
or U3097 (N_3097,N_1100,N_940);
or U3098 (N_3098,N_1536,N_741);
and U3099 (N_3099,N_1858,N_2290);
nand U3100 (N_3100,N_34,N_2056);
xnor U3101 (N_3101,N_2381,N_311);
nor U3102 (N_3102,N_734,N_399);
nor U3103 (N_3103,N_559,N_1993);
xnor U3104 (N_3104,N_343,N_2289);
or U3105 (N_3105,N_1337,N_686);
nand U3106 (N_3106,N_1248,N_2388);
or U3107 (N_3107,N_714,N_478);
xor U3108 (N_3108,N_181,N_2096);
nor U3109 (N_3109,N_2204,N_1389);
and U3110 (N_3110,N_100,N_784);
nand U3111 (N_3111,N_980,N_1059);
nor U3112 (N_3112,N_1708,N_1170);
xor U3113 (N_3113,N_1625,N_38);
xnor U3114 (N_3114,N_112,N_1975);
nor U3115 (N_3115,N_482,N_2184);
xor U3116 (N_3116,N_600,N_594);
and U3117 (N_3117,N_2477,N_135);
or U3118 (N_3118,N_1546,N_2370);
and U3119 (N_3119,N_371,N_2041);
xor U3120 (N_3120,N_1908,N_173);
xnor U3121 (N_3121,N_1182,N_210);
nand U3122 (N_3122,N_1815,N_1469);
nor U3123 (N_3123,N_2331,N_490);
nand U3124 (N_3124,N_102,N_1610);
and U3125 (N_3125,N_27,N_1640);
and U3126 (N_3126,N_380,N_2201);
and U3127 (N_3127,N_1053,N_2033);
or U3128 (N_3128,N_1049,N_168);
nor U3129 (N_3129,N_1260,N_730);
nand U3130 (N_3130,N_245,N_1336);
xnor U3131 (N_3131,N_612,N_964);
or U3132 (N_3132,N_491,N_1675);
xnor U3133 (N_3133,N_733,N_2377);
and U3134 (N_3134,N_2497,N_427);
xnor U3135 (N_3135,N_553,N_1421);
nand U3136 (N_3136,N_1598,N_2421);
nand U3137 (N_3137,N_2073,N_582);
nor U3138 (N_3138,N_2237,N_1932);
nand U3139 (N_3139,N_609,N_2318);
or U3140 (N_3140,N_1360,N_1580);
or U3141 (N_3141,N_719,N_220);
and U3142 (N_3142,N_1795,N_1327);
nand U3143 (N_3143,N_1750,N_10);
or U3144 (N_3144,N_1106,N_2120);
or U3145 (N_3145,N_2222,N_1261);
and U3146 (N_3146,N_522,N_972);
or U3147 (N_3147,N_200,N_965);
nor U3148 (N_3148,N_949,N_43);
or U3149 (N_3149,N_219,N_847);
and U3150 (N_3150,N_3,N_268);
or U3151 (N_3151,N_2375,N_636);
xnor U3152 (N_3152,N_1204,N_1251);
or U3153 (N_3153,N_1756,N_2347);
nor U3154 (N_3154,N_150,N_1695);
xnor U3155 (N_3155,N_1028,N_1731);
nand U3156 (N_3156,N_994,N_1329);
or U3157 (N_3157,N_520,N_2169);
nand U3158 (N_3158,N_1678,N_1313);
nor U3159 (N_3159,N_1934,N_1682);
and U3160 (N_3160,N_515,N_423);
xnor U3161 (N_3161,N_474,N_1304);
nor U3162 (N_3162,N_2253,N_1080);
nand U3163 (N_3163,N_1876,N_1692);
nand U3164 (N_3164,N_824,N_370);
and U3165 (N_3165,N_759,N_1366);
nor U3166 (N_3166,N_1024,N_1991);
nor U3167 (N_3167,N_2458,N_1632);
and U3168 (N_3168,N_2013,N_2418);
nand U3169 (N_3169,N_2300,N_2034);
or U3170 (N_3170,N_827,N_1980);
nor U3171 (N_3171,N_2245,N_776);
or U3172 (N_3172,N_844,N_944);
nor U3173 (N_3173,N_312,N_1253);
nand U3174 (N_3174,N_1884,N_2308);
or U3175 (N_3175,N_208,N_247);
nor U3176 (N_3176,N_525,N_1501);
and U3177 (N_3177,N_2359,N_726);
nor U3178 (N_3178,N_466,N_1426);
xnor U3179 (N_3179,N_35,N_589);
or U3180 (N_3180,N_2382,N_1056);
nor U3181 (N_3181,N_756,N_1518);
and U3182 (N_3182,N_801,N_1526);
and U3183 (N_3183,N_836,N_2383);
xor U3184 (N_3184,N_2190,N_2180);
or U3185 (N_3185,N_778,N_1628);
and U3186 (N_3186,N_1774,N_961);
nor U3187 (N_3187,N_556,N_1317);
nor U3188 (N_3188,N_1419,N_727);
xor U3189 (N_3189,N_1382,N_243);
or U3190 (N_3190,N_1440,N_1584);
and U3191 (N_3191,N_1041,N_1415);
and U3192 (N_3192,N_1514,N_711);
nand U3193 (N_3193,N_404,N_187);
nor U3194 (N_3194,N_2311,N_1949);
xor U3195 (N_3195,N_2129,N_1022);
xnor U3196 (N_3196,N_487,N_721);
xnor U3197 (N_3197,N_902,N_1279);
xnor U3198 (N_3198,N_1034,N_883);
and U3199 (N_3199,N_1126,N_1810);
nor U3200 (N_3200,N_588,N_1745);
nand U3201 (N_3201,N_346,N_1636);
nand U3202 (N_3202,N_2097,N_1585);
xor U3203 (N_3203,N_1094,N_1649);
nand U3204 (N_3204,N_1487,N_2288);
or U3205 (N_3205,N_319,N_2437);
nand U3206 (N_3206,N_1972,N_2465);
nor U3207 (N_3207,N_1176,N_382);
nand U3208 (N_3208,N_396,N_1589);
xor U3209 (N_3209,N_368,N_1089);
or U3210 (N_3210,N_503,N_44);
nor U3211 (N_3211,N_659,N_235);
xor U3212 (N_3212,N_2108,N_452);
and U3213 (N_3213,N_2257,N_1019);
nand U3214 (N_3214,N_2256,N_1);
or U3215 (N_3215,N_1693,N_1365);
or U3216 (N_3216,N_969,N_1394);
xnor U3217 (N_3217,N_69,N_1143);
or U3218 (N_3218,N_898,N_675);
nand U3219 (N_3219,N_1190,N_1378);
nor U3220 (N_3220,N_1074,N_121);
xor U3221 (N_3221,N_1502,N_1485);
xnor U3222 (N_3222,N_1151,N_799);
nand U3223 (N_3223,N_793,N_36);
nor U3224 (N_3224,N_643,N_2124);
nor U3225 (N_3225,N_1587,N_1453);
and U3226 (N_3226,N_2189,N_1023);
xor U3227 (N_3227,N_1183,N_1735);
xnor U3228 (N_3228,N_682,N_1838);
and U3229 (N_3229,N_864,N_2344);
or U3230 (N_3230,N_1757,N_280);
nor U3231 (N_3231,N_228,N_936);
or U3232 (N_3232,N_1863,N_1003);
and U3233 (N_3233,N_330,N_2027);
nor U3234 (N_3234,N_99,N_1155);
nor U3235 (N_3235,N_409,N_2004);
nand U3236 (N_3236,N_854,N_1241);
nand U3237 (N_3237,N_634,N_1310);
xnor U3238 (N_3238,N_1539,N_957);
or U3239 (N_3239,N_1659,N_284);
or U3240 (N_3240,N_205,N_1746);
nand U3241 (N_3241,N_71,N_1766);
nor U3242 (N_3242,N_1226,N_1921);
and U3243 (N_3243,N_1225,N_1663);
nand U3244 (N_3244,N_905,N_1680);
and U3245 (N_3245,N_459,N_1698);
nand U3246 (N_3246,N_1879,N_1529);
xnor U3247 (N_3247,N_2128,N_74);
or U3248 (N_3248,N_212,N_1549);
xnor U3249 (N_3249,N_1263,N_587);
xnor U3250 (N_3250,N_2262,N_829);
or U3251 (N_3251,N_1967,N_1479);
nand U3252 (N_3252,N_968,N_2202);
nand U3253 (N_3253,N_1906,N_2172);
nand U3254 (N_3254,N_2103,N_1528);
xnor U3255 (N_3255,N_1755,N_2217);
or U3256 (N_3256,N_126,N_475);
xor U3257 (N_3257,N_85,N_2474);
nand U3258 (N_3258,N_2243,N_2117);
xor U3259 (N_3259,N_506,N_2146);
and U3260 (N_3260,N_1694,N_342);
xor U3261 (N_3261,N_925,N_1913);
xor U3262 (N_3262,N_695,N_1244);
nor U3263 (N_3263,N_347,N_1779);
nor U3264 (N_3264,N_2396,N_433);
xnor U3265 (N_3265,N_1762,N_248);
xnor U3266 (N_3266,N_1801,N_514);
xor U3267 (N_3267,N_1971,N_841);
nor U3268 (N_3268,N_329,N_1234);
nor U3269 (N_3269,N_59,N_2045);
or U3270 (N_3270,N_426,N_2206);
xor U3271 (N_3271,N_1717,N_111);
and U3272 (N_3272,N_2263,N_1303);
nand U3273 (N_3273,N_277,N_387);
xor U3274 (N_3274,N_2476,N_890);
and U3275 (N_3275,N_1930,N_502);
xnor U3276 (N_3276,N_1286,N_2061);
nand U3277 (N_3277,N_691,N_366);
xnor U3278 (N_3278,N_1187,N_1601);
and U3279 (N_3279,N_1466,N_58);
nand U3280 (N_3280,N_1307,N_32);
nor U3281 (N_3281,N_914,N_2350);
xnor U3282 (N_3282,N_340,N_2051);
nor U3283 (N_3283,N_1099,N_0);
and U3284 (N_3284,N_644,N_96);
nand U3285 (N_3285,N_12,N_904);
xor U3286 (N_3286,N_1965,N_266);
or U3287 (N_3287,N_1351,N_1804);
nor U3288 (N_3288,N_895,N_1296);
nor U3289 (N_3289,N_1666,N_2009);
nor U3290 (N_3290,N_1568,N_1907);
nand U3291 (N_3291,N_953,N_1069);
nand U3292 (N_3292,N_1749,N_1015);
xor U3293 (N_3293,N_1900,N_158);
nor U3294 (N_3294,N_2379,N_1864);
nand U3295 (N_3295,N_1494,N_544);
xor U3296 (N_3296,N_364,N_418);
nor U3297 (N_3297,N_1511,N_1786);
and U3298 (N_3298,N_1403,N_272);
xnor U3299 (N_3299,N_1065,N_1178);
or U3300 (N_3300,N_2469,N_1711);
nor U3301 (N_3301,N_993,N_1161);
nand U3302 (N_3302,N_291,N_917);
xnor U3303 (N_3303,N_1417,N_2095);
nand U3304 (N_3304,N_2320,N_1769);
nand U3305 (N_3305,N_637,N_1411);
or U3306 (N_3306,N_1832,N_2277);
or U3307 (N_3307,N_1835,N_2242);
nand U3308 (N_3308,N_2268,N_2125);
or U3309 (N_3309,N_2248,N_2104);
nand U3310 (N_3310,N_2110,N_1936);
or U3311 (N_3311,N_2080,N_189);
and U3312 (N_3312,N_1465,N_660);
and U3313 (N_3313,N_560,N_2365);
and U3314 (N_3314,N_739,N_1154);
or U3315 (N_3315,N_977,N_924);
or U3316 (N_3316,N_615,N_485);
nor U3317 (N_3317,N_81,N_1368);
or U3318 (N_3318,N_1890,N_970);
and U3319 (N_3319,N_2274,N_2264);
or U3320 (N_3320,N_573,N_1097);
and U3321 (N_3321,N_454,N_2449);
or U3322 (N_3322,N_471,N_1565);
nor U3323 (N_3323,N_610,N_1250);
nor U3324 (N_3324,N_2038,N_1629);
nor U3325 (N_3325,N_1347,N_633);
nor U3326 (N_3326,N_295,N_663);
or U3327 (N_3327,N_1839,N_857);
and U3328 (N_3328,N_2196,N_1118);
or U3329 (N_3329,N_1480,N_1593);
and U3330 (N_3330,N_758,N_1237);
and U3331 (N_3331,N_865,N_2043);
and U3332 (N_3332,N_72,N_182);
and U3333 (N_3333,N_292,N_2440);
or U3334 (N_3334,N_581,N_1452);
nor U3335 (N_3335,N_685,N_1893);
and U3336 (N_3336,N_1202,N_1623);
or U3337 (N_3337,N_179,N_385);
nor U3338 (N_3338,N_666,N_1673);
xor U3339 (N_3339,N_1220,N_1269);
and U3340 (N_3340,N_1207,N_1559);
nand U3341 (N_3341,N_275,N_1405);
nand U3342 (N_3342,N_197,N_1363);
nor U3343 (N_3343,N_773,N_2236);
nand U3344 (N_3344,N_743,N_107);
and U3345 (N_3345,N_1957,N_575);
xor U3346 (N_3346,N_2372,N_1383);
xnor U3347 (N_3347,N_136,N_1704);
or U3348 (N_3348,N_65,N_846);
nor U3349 (N_3349,N_90,N_1117);
xnor U3350 (N_3350,N_222,N_1582);
xor U3351 (N_3351,N_2447,N_601);
nor U3352 (N_3352,N_1210,N_1859);
nand U3353 (N_3353,N_893,N_2209);
xnor U3354 (N_3354,N_699,N_706);
and U3355 (N_3355,N_132,N_73);
nor U3356 (N_3356,N_1218,N_570);
nor U3357 (N_3357,N_195,N_2403);
and U3358 (N_3358,N_11,N_496);
and U3359 (N_3359,N_185,N_1650);
or U3360 (N_3360,N_746,N_1188);
or U3361 (N_3361,N_2179,N_31);
xnor U3362 (N_3362,N_1719,N_2452);
or U3363 (N_3363,N_751,N_2040);
nand U3364 (N_3364,N_289,N_264);
nand U3365 (N_3365,N_812,N_1567);
nor U3366 (N_3366,N_2042,N_1881);
and U3367 (N_3367,N_1018,N_167);
nor U3368 (N_3368,N_20,N_436);
and U3369 (N_3369,N_510,N_237);
or U3370 (N_3370,N_259,N_818);
and U3371 (N_3371,N_25,N_1247);
nand U3372 (N_3372,N_1595,N_690);
and U3373 (N_3373,N_1866,N_274);
xnor U3374 (N_3374,N_1922,N_1818);
nor U3375 (N_3375,N_2145,N_300);
or U3376 (N_3376,N_2485,N_1948);
or U3377 (N_3377,N_1318,N_1627);
xnor U3378 (N_3378,N_833,N_29);
nor U3379 (N_3379,N_782,N_606);
and U3380 (N_3380,N_2329,N_1959);
or U3381 (N_3381,N_1083,N_1701);
nor U3382 (N_3382,N_327,N_1486);
and U3383 (N_3383,N_2008,N_1438);
xnor U3384 (N_3384,N_1646,N_2446);
or U3385 (N_3385,N_62,N_1471);
nor U3386 (N_3386,N_2017,N_2466);
nor U3387 (N_3387,N_287,N_1869);
nor U3388 (N_3388,N_1195,N_1219);
nor U3389 (N_3389,N_599,N_1085);
or U3390 (N_3390,N_2025,N_1384);
and U3391 (N_3391,N_414,N_1079);
nor U3392 (N_3392,N_130,N_1778);
or U3393 (N_3393,N_1461,N_916);
nand U3394 (N_3394,N_900,N_1530);
nand U3395 (N_3395,N_2007,N_1277);
or U3396 (N_3396,N_37,N_2185);
nor U3397 (N_3397,N_1252,N_232);
nand U3398 (N_3398,N_753,N_1660);
and U3399 (N_3399,N_2156,N_942);
or U3400 (N_3400,N_2199,N_2281);
xnor U3401 (N_3401,N_2416,N_1141);
or U3402 (N_3402,N_56,N_263);
nand U3403 (N_3403,N_911,N_1246);
nand U3404 (N_3404,N_2029,N_1761);
xnor U3405 (N_3405,N_1776,N_202);
and U3406 (N_3406,N_1574,N_2003);
nor U3407 (N_3407,N_584,N_1740);
and U3408 (N_3408,N_820,N_1001);
or U3409 (N_3409,N_231,N_224);
nor U3410 (N_3410,N_1078,N_1733);
xor U3411 (N_3411,N_465,N_1662);
nor U3412 (N_3412,N_1104,N_1377);
or U3413 (N_3413,N_1896,N_2415);
nor U3414 (N_3414,N_768,N_2389);
nand U3415 (N_3415,N_1071,N_2016);
nand U3416 (N_3416,N_832,N_539);
nor U3417 (N_3417,N_1630,N_2200);
nand U3418 (N_3418,N_66,N_631);
nor U3419 (N_3419,N_2079,N_196);
nand U3420 (N_3420,N_1333,N_1463);
nor U3421 (N_3421,N_1875,N_1129);
nand U3422 (N_3422,N_1889,N_2135);
or U3423 (N_3423,N_867,N_2470);
xnor U3424 (N_3424,N_2349,N_1620);
or U3425 (N_3425,N_763,N_1396);
nor U3426 (N_3426,N_54,N_744);
or U3427 (N_3427,N_2438,N_388);
or U3428 (N_3428,N_2011,N_1507);
or U3429 (N_3429,N_2251,N_2083);
or U3430 (N_3430,N_1047,N_973);
or U3431 (N_3431,N_1067,N_2353);
xnor U3432 (N_3432,N_2054,N_2265);
xnor U3433 (N_3433,N_267,N_1827);
or U3434 (N_3434,N_538,N_1935);
nor U3435 (N_3435,N_137,N_737);
or U3436 (N_3436,N_2031,N_170);
nor U3437 (N_3437,N_2406,N_1600);
xor U3438 (N_3438,N_49,N_1236);
and U3439 (N_3439,N_78,N_51);
xor U3440 (N_3440,N_2161,N_1872);
nand U3441 (N_3441,N_2229,N_2367);
xor U3442 (N_3442,N_694,N_98);
or U3443 (N_3443,N_153,N_1612);
nand U3444 (N_3444,N_379,N_1836);
nor U3445 (N_3445,N_1730,N_1943);
nand U3446 (N_3446,N_1851,N_241);
and U3447 (N_3447,N_2473,N_2068);
nand U3448 (N_3448,N_1339,N_70);
nand U3449 (N_3449,N_761,N_470);
xor U3450 (N_3450,N_1726,N_2028);
and U3451 (N_3451,N_1981,N_2436);
or U3452 (N_3452,N_1021,N_2456);
xnor U3453 (N_3453,N_2193,N_1044);
and U3454 (N_3454,N_1988,N_804);
nor U3455 (N_3455,N_2035,N_1591);
xor U3456 (N_3456,N_398,N_967);
and U3457 (N_3457,N_552,N_6);
or U3458 (N_3458,N_985,N_2360);
nor U3459 (N_3459,N_254,N_2430);
or U3460 (N_3460,N_2314,N_577);
or U3461 (N_3461,N_1054,N_91);
nand U3462 (N_3462,N_811,N_1850);
and U3463 (N_3463,N_1010,N_667);
nor U3464 (N_3464,N_52,N_1292);
xor U3465 (N_3465,N_1523,N_2227);
nand U3466 (N_3466,N_2000,N_4);
xnor U3467 (N_3467,N_229,N_1391);
or U3468 (N_3468,N_1025,N_336);
nor U3469 (N_3469,N_1898,N_1373);
nor U3470 (N_3470,N_1670,N_2471);
and U3471 (N_3471,N_1515,N_1410);
or U3472 (N_3472,N_1513,N_456);
and U3473 (N_3473,N_1868,N_2052);
or U3474 (N_3474,N_1319,N_611);
xor U3475 (N_3475,N_2234,N_1343);
nor U3476 (N_3476,N_2133,N_1970);
nand U3477 (N_3477,N_394,N_236);
or U3478 (N_3478,N_230,N_238);
nand U3479 (N_3479,N_529,N_355);
nand U3480 (N_3480,N_2244,N_817);
or U3481 (N_3481,N_2118,N_1422);
or U3482 (N_3482,N_2399,N_1503);
or U3483 (N_3483,N_1825,N_518);
nand U3484 (N_3484,N_1454,N_635);
nand U3485 (N_3485,N_1095,N_2394);
or U3486 (N_3486,N_2496,N_1616);
or U3487 (N_3487,N_2240,N_2404);
nor U3488 (N_3488,N_1344,N_906);
xor U3489 (N_3489,N_2211,N_561);
nand U3490 (N_3490,N_2366,N_1547);
nand U3491 (N_3491,N_89,N_2142);
nand U3492 (N_3492,N_416,N_2092);
nor U3493 (N_3493,N_772,N_2151);
and U3494 (N_3494,N_1605,N_1064);
nand U3495 (N_3495,N_2494,N_939);
or U3496 (N_3496,N_1135,N_2336);
and U3497 (N_3497,N_1771,N_2130);
and U3498 (N_3498,N_848,N_997);
nand U3499 (N_3499,N_1834,N_794);
and U3500 (N_3500,N_1911,N_1703);
or U3501 (N_3501,N_1282,N_1201);
or U3502 (N_3502,N_378,N_1688);
or U3503 (N_3503,N_60,N_1166);
xnor U3504 (N_3504,N_2380,N_1153);
or U3505 (N_3505,N_869,N_1380);
or U3506 (N_3506,N_1300,N_513);
and U3507 (N_3507,N_402,N_2316);
and U3508 (N_3508,N_214,N_2064);
nand U3509 (N_3509,N_678,N_244);
nand U3510 (N_3510,N_1475,N_2014);
nand U3511 (N_3511,N_1732,N_1828);
or U3512 (N_3512,N_2010,N_810);
nor U3513 (N_3513,N_276,N_1346);
nor U3514 (N_3514,N_1036,N_2408);
xor U3515 (N_3515,N_2225,N_1222);
and U3516 (N_3516,N_1525,N_512);
and U3517 (N_3517,N_1578,N_722);
nor U3518 (N_3518,N_348,N_629);
and U3519 (N_3519,N_363,N_2493);
and U3520 (N_3520,N_1268,N_2410);
nand U3521 (N_3521,N_2448,N_1689);
or U3522 (N_3522,N_1738,N_2147);
nand U3523 (N_3523,N_1472,N_2191);
and U3524 (N_3524,N_428,N_221);
xnor U3525 (N_3525,N_1686,N_1255);
and U3526 (N_3526,N_1982,N_550);
nand U3527 (N_3527,N_151,N_1488);
nand U3528 (N_3528,N_2459,N_608);
nor U3529 (N_3529,N_1576,N_830);
and U3530 (N_3530,N_2498,N_391);
xnor U3531 (N_3531,N_1571,N_1807);
xor U3532 (N_3532,N_1353,N_9);
and U3533 (N_3533,N_2315,N_1727);
nor U3534 (N_3534,N_2099,N_120);
nor U3535 (N_3535,N_1424,N_1563);
and U3536 (N_3536,N_204,N_1259);
nor U3537 (N_3537,N_1134,N_299);
nand U3538 (N_3538,N_453,N_875);
nand U3539 (N_3539,N_2085,N_40);
and U3540 (N_3540,N_987,N_2280);
nand U3541 (N_3541,N_262,N_931);
nor U3542 (N_3542,N_862,N_410);
nand U3543 (N_3543,N_946,N_147);
xor U3544 (N_3544,N_349,N_169);
nor U3545 (N_3545,N_1588,N_1551);
xnor U3546 (N_3546,N_2170,N_1512);
nand U3547 (N_3547,N_533,N_1780);
nand U3548 (N_3548,N_704,N_1996);
nand U3549 (N_3549,N_14,N_1506);
nor U3550 (N_3550,N_1961,N_457);
xnor U3551 (N_3551,N_519,N_1556);
nand U3552 (N_3552,N_1355,N_1406);
nand U3553 (N_3553,N_2005,N_585);
and U3554 (N_3554,N_614,N_1797);
xor U3555 (N_3555,N_1677,N_1926);
and U3556 (N_3556,N_2411,N_1964);
xnor U3557 (N_3557,N_1283,N_2066);
nor U3558 (N_3558,N_792,N_2198);
nand U3559 (N_3559,N_361,N_747);
nor U3560 (N_3560,N_1696,N_2165);
nand U3561 (N_3561,N_1944,N_2299);
nor U3562 (N_3562,N_443,N_1985);
and U3563 (N_3563,N_193,N_2355);
nand U3564 (N_3564,N_1586,N_915);
nor U3565 (N_3565,N_1444,N_296);
or U3566 (N_3566,N_2152,N_527);
and U3567 (N_3567,N_1877,N_616);
or U3568 (N_3568,N_1912,N_2098);
or U3569 (N_3569,N_1671,N_882);
or U3570 (N_3570,N_2197,N_33);
xor U3571 (N_3571,N_1112,N_1297);
nand U3572 (N_3572,N_628,N_2275);
or U3573 (N_3573,N_356,N_2286);
nand U3574 (N_3574,N_438,N_680);
nor U3575 (N_3575,N_460,N_164);
and U3576 (N_3576,N_791,N_712);
and U3577 (N_3577,N_1481,N_1974);
and U3578 (N_3578,N_177,N_1181);
xor U3579 (N_3579,N_934,N_951);
xnor U3580 (N_3580,N_592,N_907);
and U3581 (N_3581,N_1194,N_1088);
nor U3582 (N_3582,N_2284,N_2273);
and U3583 (N_3583,N_1919,N_536);
or U3584 (N_3584,N_531,N_1191);
or U3585 (N_3585,N_450,N_1792);
nor U3586 (N_3586,N_1075,N_446);
nor U3587 (N_3587,N_2443,N_1264);
xor U3588 (N_3588,N_1652,N_117);
and U3589 (N_3589,N_1121,N_1845);
xor U3590 (N_3590,N_1043,N_1618);
or U3591 (N_3591,N_2278,N_1408);
xnor U3592 (N_3592,N_2478,N_1168);
and U3593 (N_3593,N_1751,N_1398);
nor U3594 (N_3594,N_1707,N_1063);
or U3595 (N_3595,N_412,N_1990);
nor U3596 (N_3596,N_831,N_2150);
nor U3597 (N_3597,N_217,N_2423);
or U3598 (N_3598,N_822,N_144);
nand U3599 (N_3599,N_495,N_593);
and U3600 (N_3600,N_908,N_492);
nor U3601 (N_3601,N_178,N_2376);
and U3602 (N_3602,N_1493,N_954);
xnor U3603 (N_3603,N_1767,N_157);
and U3604 (N_3604,N_2348,N_1554);
nor U3605 (N_3605,N_672,N_2322);
nor U3606 (N_3606,N_1520,N_1947);
nor U3607 (N_3607,N_1803,N_2258);
nor U3608 (N_3608,N_1407,N_2235);
nand U3609 (N_3609,N_2295,N_2327);
and U3610 (N_3610,N_1113,N_1470);
nor U3611 (N_3611,N_2302,N_1012);
nor U3612 (N_3612,N_22,N_1725);
nor U3613 (N_3613,N_2259,N_1883);
and U3614 (N_3614,N_1331,N_2451);
and U3615 (N_3615,N_2454,N_2285);
and U3616 (N_3616,N_1316,N_1550);
nor U3617 (N_3617,N_885,N_390);
and U3618 (N_3618,N_1171,N_322);
xnor U3619 (N_3619,N_1781,N_1508);
nand U3620 (N_3620,N_28,N_2164);
and U3621 (N_3621,N_1817,N_1196);
nand U3622 (N_3622,N_407,N_1941);
xnor U3623 (N_3623,N_815,N_1123);
and U3624 (N_3624,N_1873,N_1174);
and U3625 (N_3625,N_2254,N_1358);
xnor U3626 (N_3626,N_1267,N_2208);
nand U3627 (N_3627,N_1560,N_2378);
nor U3628 (N_3628,N_46,N_1441);
and U3629 (N_3629,N_1914,N_122);
nor U3630 (N_3630,N_159,N_1609);
xor U3631 (N_3631,N_57,N_718);
or U3632 (N_3632,N_317,N_1759);
xor U3633 (N_3633,N_1295,N_1114);
xor U3634 (N_3634,N_1821,N_2293);
and U3635 (N_3635,N_2405,N_2218);
and U3636 (N_3636,N_1860,N_302);
nor U3637 (N_3637,N_1456,N_2419);
xnor U3638 (N_3638,N_2324,N_541);
xnor U3639 (N_3639,N_462,N_2357);
xor U3640 (N_3640,N_671,N_775);
xnor U3641 (N_3641,N_2333,N_2484);
nand U3642 (N_3642,N_1951,N_1223);
nor U3643 (N_3643,N_1655,N_140);
or U3644 (N_3644,N_2305,N_814);
nor U3645 (N_3645,N_1315,N_306);
nand U3646 (N_3646,N_971,N_642);
nand U3647 (N_3647,N_48,N_569);
xnor U3648 (N_3648,N_2065,N_1231);
and U3649 (N_3649,N_646,N_1867);
nor U3650 (N_3650,N_2174,N_1198);
nand U3651 (N_3651,N_2296,N_1173);
nor U3652 (N_3652,N_640,N_1984);
xor U3653 (N_3653,N_871,N_2136);
and U3654 (N_3654,N_1862,N_884);
and U3655 (N_3655,N_313,N_1338);
or U3656 (N_3656,N_1395,N_1789);
and U3657 (N_3657,N_2397,N_1309);
or U3658 (N_3658,N_1668,N_374);
xor U3659 (N_3659,N_1284,N_1030);
nor U3660 (N_3660,N_543,N_1462);
or U3661 (N_3661,N_1592,N_2089);
or U3662 (N_3662,N_110,N_2233);
nand U3663 (N_3663,N_1367,N_19);
xor U3664 (N_3664,N_526,N_1517);
and U3665 (N_3665,N_2491,N_735);
xor U3666 (N_3666,N_1359,N_1144);
and U3667 (N_3667,N_909,N_781);
and U3668 (N_3668,N_700,N_1923);
or U3669 (N_3669,N_572,N_1744);
xnor U3670 (N_3670,N_2186,N_1464);
and U3671 (N_3671,N_373,N_1977);
nand U3672 (N_3672,N_652,N_528);
nand U3673 (N_3673,N_1613,N_1302);
xor U3674 (N_3674,N_7,N_2);
nand U3675 (N_3675,N_2455,N_1702);
or U3676 (N_3676,N_2487,N_1813);
and U3677 (N_3677,N_55,N_2427);
xor U3678 (N_3678,N_1437,N_1111);
or U3679 (N_3679,N_790,N_449);
xnor U3680 (N_3680,N_251,N_143);
or U3681 (N_3681,N_1032,N_1119);
or U3682 (N_3682,N_1928,N_2335);
xnor U3683 (N_3683,N_389,N_2312);
and U3684 (N_3684,N_146,N_2402);
or U3685 (N_3685,N_1791,N_2457);
or U3686 (N_3686,N_2226,N_1402);
nor U3687 (N_3687,N_451,N_803);
and U3688 (N_3688,N_679,N_2486);
nand U3689 (N_3689,N_1105,N_1342);
nor U3690 (N_3690,N_596,N_868);
nor U3691 (N_3691,N_134,N_576);
or U3692 (N_3692,N_1107,N_1401);
nand U3693 (N_3693,N_2368,N_8);
nor U3694 (N_3694,N_345,N_108);
nand U3695 (N_3695,N_2260,N_2468);
or U3696 (N_3696,N_1238,N_604);
xor U3697 (N_3697,N_858,N_1213);
and U3698 (N_3698,N_1758,N_352);
and U3699 (N_3699,N_2046,N_421);
nor U3700 (N_3700,N_1086,N_15);
nand U3701 (N_3701,N_1739,N_779);
xor U3702 (N_3702,N_795,N_403);
nor U3703 (N_3703,N_191,N_1856);
xnor U3704 (N_3704,N_1657,N_1566);
and U3705 (N_3705,N_1765,N_1433);
or U3706 (N_3706,N_1068,N_507);
xor U3707 (N_3707,N_1245,N_1962);
and U3708 (N_3708,N_982,N_2249);
xor U3709 (N_3709,N_1840,N_800);
and U3710 (N_3710,N_442,N_2340);
nand U3711 (N_3711,N_1026,N_976);
or U3712 (N_3712,N_2210,N_129);
or U3713 (N_3713,N_1200,N_1672);
xor U3714 (N_3714,N_17,N_1728);
xor U3715 (N_3715,N_532,N_595);
or U3716 (N_3716,N_1899,N_1125);
or U3717 (N_3717,N_2387,N_213);
nand U3718 (N_3718,N_293,N_2158);
nand U3719 (N_3719,N_79,N_2036);
xor U3720 (N_3720,N_1783,N_335);
nor U3721 (N_3721,N_2345,N_255);
and U3722 (N_3722,N_493,N_1931);
nor U3723 (N_3723,N_813,N_2214);
nand U3724 (N_3724,N_745,N_1638);
and U3725 (N_3725,N_597,N_2069);
or U3726 (N_3726,N_1254,N_314);
xor U3727 (N_3727,N_1741,N_350);
xnor U3728 (N_3728,N_922,N_1966);
nor U3729 (N_3729,N_341,N_1414);
and U3730 (N_3730,N_1014,N_2138);
and U3731 (N_3731,N_2081,N_1416);
xor U3732 (N_3732,N_1534,N_1147);
and U3733 (N_3733,N_1388,N_294);
nor U3734 (N_3734,N_1376,N_894);
or U3735 (N_3735,N_441,N_1330);
xnor U3736 (N_3736,N_547,N_271);
and U3737 (N_3737,N_406,N_1460);
or U3738 (N_3738,N_2354,N_1077);
or U3739 (N_3739,N_1634,N_2409);
or U3740 (N_3740,N_1790,N_2012);
nor U3741 (N_3741,N_2140,N_1705);
nor U3742 (N_3742,N_1709,N_357);
or U3743 (N_3743,N_1051,N_508);
nor U3744 (N_3744,N_2115,N_816);
nor U3745 (N_3745,N_2356,N_1332);
nand U3746 (N_3746,N_1167,N_2048);
or U3747 (N_3747,N_1397,N_2153);
nand U3748 (N_3748,N_2139,N_2053);
or U3749 (N_3749,N_285,N_1005);
nand U3750 (N_3750,N_126,N_384);
xnor U3751 (N_3751,N_2403,N_2490);
xnor U3752 (N_3752,N_1257,N_1945);
and U3753 (N_3753,N_311,N_762);
xor U3754 (N_3754,N_407,N_1552);
xor U3755 (N_3755,N_671,N_542);
xor U3756 (N_3756,N_2094,N_886);
and U3757 (N_3757,N_39,N_2259);
xnor U3758 (N_3758,N_1385,N_545);
xor U3759 (N_3759,N_432,N_481);
or U3760 (N_3760,N_403,N_1191);
nand U3761 (N_3761,N_54,N_515);
nor U3762 (N_3762,N_198,N_2053);
nor U3763 (N_3763,N_2264,N_1610);
or U3764 (N_3764,N_1850,N_588);
xnor U3765 (N_3765,N_2276,N_2348);
xnor U3766 (N_3766,N_2156,N_1108);
or U3767 (N_3767,N_2124,N_1559);
nand U3768 (N_3768,N_2310,N_424);
nor U3769 (N_3769,N_1180,N_155);
and U3770 (N_3770,N_2236,N_961);
or U3771 (N_3771,N_1683,N_2182);
nor U3772 (N_3772,N_348,N_44);
nor U3773 (N_3773,N_794,N_2365);
nand U3774 (N_3774,N_417,N_969);
nand U3775 (N_3775,N_2430,N_1481);
nor U3776 (N_3776,N_736,N_1021);
nand U3777 (N_3777,N_618,N_1174);
nor U3778 (N_3778,N_444,N_1071);
nor U3779 (N_3779,N_1755,N_1063);
and U3780 (N_3780,N_1759,N_1541);
nand U3781 (N_3781,N_542,N_2245);
or U3782 (N_3782,N_1249,N_1149);
or U3783 (N_3783,N_1090,N_997);
xnor U3784 (N_3784,N_861,N_1837);
nor U3785 (N_3785,N_986,N_1807);
xnor U3786 (N_3786,N_565,N_1217);
and U3787 (N_3787,N_1135,N_71);
nand U3788 (N_3788,N_1201,N_13);
nor U3789 (N_3789,N_2095,N_2073);
or U3790 (N_3790,N_889,N_906);
nor U3791 (N_3791,N_1419,N_1397);
nand U3792 (N_3792,N_881,N_1251);
nand U3793 (N_3793,N_867,N_602);
nor U3794 (N_3794,N_296,N_933);
nand U3795 (N_3795,N_1050,N_2096);
nand U3796 (N_3796,N_927,N_2491);
or U3797 (N_3797,N_1463,N_136);
xnor U3798 (N_3798,N_188,N_509);
nand U3799 (N_3799,N_1214,N_319);
nand U3800 (N_3800,N_946,N_1033);
xor U3801 (N_3801,N_1048,N_2435);
xor U3802 (N_3802,N_584,N_43);
nand U3803 (N_3803,N_1887,N_282);
nor U3804 (N_3804,N_2040,N_1915);
and U3805 (N_3805,N_1135,N_3);
and U3806 (N_3806,N_664,N_107);
and U3807 (N_3807,N_59,N_1410);
or U3808 (N_3808,N_810,N_338);
nor U3809 (N_3809,N_953,N_757);
nor U3810 (N_3810,N_1268,N_1605);
nand U3811 (N_3811,N_1401,N_1925);
xnor U3812 (N_3812,N_635,N_1930);
and U3813 (N_3813,N_1640,N_90);
nand U3814 (N_3814,N_875,N_1323);
and U3815 (N_3815,N_2061,N_2283);
and U3816 (N_3816,N_671,N_120);
nand U3817 (N_3817,N_1916,N_1713);
or U3818 (N_3818,N_852,N_765);
and U3819 (N_3819,N_1847,N_1213);
and U3820 (N_3820,N_1403,N_1596);
or U3821 (N_3821,N_1879,N_1081);
or U3822 (N_3822,N_79,N_1239);
and U3823 (N_3823,N_521,N_334);
and U3824 (N_3824,N_1442,N_582);
and U3825 (N_3825,N_2240,N_1693);
nand U3826 (N_3826,N_661,N_1409);
or U3827 (N_3827,N_157,N_2336);
and U3828 (N_3828,N_2082,N_270);
or U3829 (N_3829,N_534,N_115);
or U3830 (N_3830,N_135,N_1084);
nor U3831 (N_3831,N_1998,N_1821);
nor U3832 (N_3832,N_2468,N_2202);
and U3833 (N_3833,N_830,N_483);
and U3834 (N_3834,N_1666,N_1927);
and U3835 (N_3835,N_2327,N_1412);
or U3836 (N_3836,N_624,N_323);
and U3837 (N_3837,N_1003,N_531);
xor U3838 (N_3838,N_1952,N_927);
nand U3839 (N_3839,N_1115,N_997);
or U3840 (N_3840,N_752,N_266);
or U3841 (N_3841,N_220,N_798);
xnor U3842 (N_3842,N_1513,N_2018);
nor U3843 (N_3843,N_400,N_1139);
nand U3844 (N_3844,N_1736,N_1501);
nor U3845 (N_3845,N_914,N_2093);
and U3846 (N_3846,N_2318,N_1014);
nand U3847 (N_3847,N_2274,N_1225);
nor U3848 (N_3848,N_1232,N_1588);
nand U3849 (N_3849,N_2142,N_2257);
or U3850 (N_3850,N_2080,N_2471);
nand U3851 (N_3851,N_905,N_563);
xor U3852 (N_3852,N_932,N_311);
and U3853 (N_3853,N_88,N_39);
nand U3854 (N_3854,N_525,N_1006);
nor U3855 (N_3855,N_1385,N_564);
or U3856 (N_3856,N_2257,N_1570);
and U3857 (N_3857,N_1299,N_207);
or U3858 (N_3858,N_129,N_1887);
nor U3859 (N_3859,N_1398,N_1556);
nor U3860 (N_3860,N_1011,N_2293);
xor U3861 (N_3861,N_2095,N_1543);
nor U3862 (N_3862,N_626,N_2164);
xor U3863 (N_3863,N_1729,N_368);
and U3864 (N_3864,N_62,N_2218);
and U3865 (N_3865,N_224,N_2080);
and U3866 (N_3866,N_1808,N_1641);
or U3867 (N_3867,N_355,N_2452);
nor U3868 (N_3868,N_474,N_497);
and U3869 (N_3869,N_91,N_1720);
and U3870 (N_3870,N_502,N_2435);
and U3871 (N_3871,N_747,N_667);
nand U3872 (N_3872,N_806,N_2442);
nor U3873 (N_3873,N_2457,N_443);
or U3874 (N_3874,N_894,N_898);
nand U3875 (N_3875,N_2209,N_607);
or U3876 (N_3876,N_366,N_634);
xnor U3877 (N_3877,N_1752,N_2230);
xnor U3878 (N_3878,N_5,N_2456);
or U3879 (N_3879,N_1384,N_1042);
and U3880 (N_3880,N_1574,N_171);
or U3881 (N_3881,N_1551,N_1663);
and U3882 (N_3882,N_1528,N_1484);
or U3883 (N_3883,N_1902,N_1836);
nand U3884 (N_3884,N_2452,N_1929);
and U3885 (N_3885,N_2189,N_2353);
nand U3886 (N_3886,N_2022,N_2427);
nand U3887 (N_3887,N_1249,N_2494);
nand U3888 (N_3888,N_369,N_2309);
or U3889 (N_3889,N_1645,N_315);
nand U3890 (N_3890,N_1507,N_1177);
nand U3891 (N_3891,N_1348,N_354);
or U3892 (N_3892,N_1241,N_2030);
nand U3893 (N_3893,N_1892,N_1479);
nor U3894 (N_3894,N_1557,N_1589);
and U3895 (N_3895,N_1511,N_158);
xor U3896 (N_3896,N_452,N_613);
nor U3897 (N_3897,N_1607,N_370);
nand U3898 (N_3898,N_1357,N_1452);
xnor U3899 (N_3899,N_39,N_42);
xnor U3900 (N_3900,N_800,N_259);
or U3901 (N_3901,N_400,N_1985);
nand U3902 (N_3902,N_657,N_1703);
or U3903 (N_3903,N_512,N_2343);
xnor U3904 (N_3904,N_1467,N_2142);
or U3905 (N_3905,N_2494,N_1165);
xnor U3906 (N_3906,N_1239,N_940);
nand U3907 (N_3907,N_1316,N_901);
or U3908 (N_3908,N_2260,N_23);
nor U3909 (N_3909,N_2479,N_2491);
and U3910 (N_3910,N_2178,N_2362);
nand U3911 (N_3911,N_1896,N_1530);
nand U3912 (N_3912,N_1668,N_2122);
or U3913 (N_3913,N_826,N_782);
nand U3914 (N_3914,N_1020,N_302);
or U3915 (N_3915,N_385,N_2462);
nor U3916 (N_3916,N_1754,N_2418);
nor U3917 (N_3917,N_2040,N_210);
or U3918 (N_3918,N_956,N_704);
xor U3919 (N_3919,N_1818,N_1842);
nor U3920 (N_3920,N_1648,N_760);
xnor U3921 (N_3921,N_1856,N_1301);
and U3922 (N_3922,N_1754,N_28);
nor U3923 (N_3923,N_2358,N_2433);
nor U3924 (N_3924,N_1446,N_972);
nor U3925 (N_3925,N_1444,N_1934);
xor U3926 (N_3926,N_1854,N_1464);
nor U3927 (N_3927,N_1763,N_25);
and U3928 (N_3928,N_1299,N_175);
nand U3929 (N_3929,N_196,N_1939);
and U3930 (N_3930,N_2497,N_2044);
or U3931 (N_3931,N_1306,N_195);
nand U3932 (N_3932,N_42,N_1730);
and U3933 (N_3933,N_1494,N_2221);
and U3934 (N_3934,N_2403,N_1487);
or U3935 (N_3935,N_1546,N_2175);
or U3936 (N_3936,N_565,N_1414);
xor U3937 (N_3937,N_459,N_2217);
or U3938 (N_3938,N_2384,N_1745);
nand U3939 (N_3939,N_1627,N_1476);
xnor U3940 (N_3940,N_300,N_1411);
nor U3941 (N_3941,N_1301,N_2240);
and U3942 (N_3942,N_2460,N_1178);
and U3943 (N_3943,N_1822,N_1027);
xnor U3944 (N_3944,N_716,N_304);
xor U3945 (N_3945,N_1183,N_1102);
xnor U3946 (N_3946,N_160,N_721);
xor U3947 (N_3947,N_2327,N_2209);
nor U3948 (N_3948,N_1685,N_2307);
xnor U3949 (N_3949,N_2194,N_2245);
nand U3950 (N_3950,N_2136,N_145);
xnor U3951 (N_3951,N_435,N_1901);
nand U3952 (N_3952,N_1039,N_1422);
xor U3953 (N_3953,N_2467,N_2472);
xnor U3954 (N_3954,N_1809,N_1556);
xor U3955 (N_3955,N_2043,N_2196);
nor U3956 (N_3956,N_2001,N_344);
or U3957 (N_3957,N_2117,N_1319);
nor U3958 (N_3958,N_39,N_674);
or U3959 (N_3959,N_899,N_2089);
nand U3960 (N_3960,N_2111,N_140);
xor U3961 (N_3961,N_954,N_323);
xnor U3962 (N_3962,N_110,N_1798);
xnor U3963 (N_3963,N_2450,N_869);
xor U3964 (N_3964,N_830,N_1589);
nand U3965 (N_3965,N_1284,N_2378);
and U3966 (N_3966,N_1028,N_2425);
xnor U3967 (N_3967,N_1099,N_2428);
and U3968 (N_3968,N_2158,N_406);
and U3969 (N_3969,N_2207,N_1619);
and U3970 (N_3970,N_1861,N_1754);
and U3971 (N_3971,N_469,N_1040);
and U3972 (N_3972,N_1791,N_786);
and U3973 (N_3973,N_2498,N_1608);
nand U3974 (N_3974,N_908,N_2010);
nor U3975 (N_3975,N_1114,N_583);
nand U3976 (N_3976,N_1255,N_1691);
nor U3977 (N_3977,N_1361,N_24);
or U3978 (N_3978,N_459,N_2353);
nand U3979 (N_3979,N_1627,N_495);
and U3980 (N_3980,N_2492,N_1219);
nor U3981 (N_3981,N_2001,N_976);
or U3982 (N_3982,N_157,N_147);
nand U3983 (N_3983,N_1169,N_1187);
xnor U3984 (N_3984,N_327,N_1557);
xnor U3985 (N_3985,N_698,N_340);
nand U3986 (N_3986,N_1502,N_2375);
and U3987 (N_3987,N_528,N_2100);
or U3988 (N_3988,N_1525,N_1772);
nand U3989 (N_3989,N_905,N_566);
and U3990 (N_3990,N_1662,N_1143);
nor U3991 (N_3991,N_1436,N_1334);
xor U3992 (N_3992,N_2497,N_2485);
nand U3993 (N_3993,N_2442,N_897);
or U3994 (N_3994,N_2424,N_32);
nor U3995 (N_3995,N_561,N_2374);
nor U3996 (N_3996,N_1886,N_131);
nand U3997 (N_3997,N_2281,N_1927);
or U3998 (N_3998,N_1376,N_512);
nor U3999 (N_3999,N_57,N_801);
or U4000 (N_4000,N_719,N_2101);
xnor U4001 (N_4001,N_771,N_1429);
nand U4002 (N_4002,N_417,N_1513);
and U4003 (N_4003,N_1969,N_1945);
or U4004 (N_4004,N_88,N_346);
nand U4005 (N_4005,N_1018,N_2219);
nand U4006 (N_4006,N_1662,N_1282);
xnor U4007 (N_4007,N_329,N_2003);
and U4008 (N_4008,N_2046,N_680);
nor U4009 (N_4009,N_839,N_307);
xnor U4010 (N_4010,N_1805,N_2362);
and U4011 (N_4011,N_1826,N_1733);
nand U4012 (N_4012,N_2244,N_1592);
nand U4013 (N_4013,N_1785,N_1662);
nand U4014 (N_4014,N_638,N_2280);
xor U4015 (N_4015,N_1890,N_1224);
and U4016 (N_4016,N_1761,N_1259);
and U4017 (N_4017,N_1351,N_1496);
nor U4018 (N_4018,N_1325,N_1808);
xnor U4019 (N_4019,N_1501,N_1401);
and U4020 (N_4020,N_1461,N_1397);
nand U4021 (N_4021,N_749,N_260);
nor U4022 (N_4022,N_569,N_1929);
nor U4023 (N_4023,N_1730,N_1851);
or U4024 (N_4024,N_580,N_1490);
or U4025 (N_4025,N_1021,N_2373);
or U4026 (N_4026,N_280,N_1914);
or U4027 (N_4027,N_1902,N_2242);
nand U4028 (N_4028,N_2130,N_1498);
nand U4029 (N_4029,N_1442,N_1772);
nand U4030 (N_4030,N_1148,N_1779);
or U4031 (N_4031,N_2249,N_2381);
xor U4032 (N_4032,N_1730,N_1654);
nand U4033 (N_4033,N_593,N_797);
xnor U4034 (N_4034,N_2491,N_123);
nand U4035 (N_4035,N_2281,N_759);
nor U4036 (N_4036,N_2144,N_192);
xnor U4037 (N_4037,N_1935,N_1042);
or U4038 (N_4038,N_1200,N_125);
nor U4039 (N_4039,N_1435,N_1957);
xor U4040 (N_4040,N_2091,N_2345);
and U4041 (N_4041,N_2165,N_1371);
nand U4042 (N_4042,N_2443,N_1875);
nor U4043 (N_4043,N_1658,N_738);
nand U4044 (N_4044,N_196,N_2486);
and U4045 (N_4045,N_2138,N_209);
or U4046 (N_4046,N_177,N_1282);
or U4047 (N_4047,N_1990,N_2397);
nor U4048 (N_4048,N_2328,N_126);
nor U4049 (N_4049,N_1379,N_2096);
nand U4050 (N_4050,N_412,N_818);
nand U4051 (N_4051,N_994,N_448);
xor U4052 (N_4052,N_789,N_1431);
and U4053 (N_4053,N_1940,N_2188);
or U4054 (N_4054,N_1877,N_1520);
nor U4055 (N_4055,N_1197,N_65);
xnor U4056 (N_4056,N_2192,N_2319);
xor U4057 (N_4057,N_426,N_2416);
xor U4058 (N_4058,N_1777,N_870);
nand U4059 (N_4059,N_75,N_2326);
nor U4060 (N_4060,N_654,N_1638);
and U4061 (N_4061,N_204,N_963);
xnor U4062 (N_4062,N_1705,N_38);
and U4063 (N_4063,N_1491,N_975);
and U4064 (N_4064,N_184,N_116);
or U4065 (N_4065,N_1056,N_1651);
nor U4066 (N_4066,N_479,N_1853);
nor U4067 (N_4067,N_125,N_2245);
nor U4068 (N_4068,N_227,N_2415);
nand U4069 (N_4069,N_355,N_86);
and U4070 (N_4070,N_1834,N_594);
xor U4071 (N_4071,N_366,N_1101);
and U4072 (N_4072,N_1740,N_1950);
xnor U4073 (N_4073,N_1849,N_1983);
xor U4074 (N_4074,N_1391,N_288);
nor U4075 (N_4075,N_412,N_2364);
and U4076 (N_4076,N_1403,N_2279);
and U4077 (N_4077,N_103,N_2123);
nand U4078 (N_4078,N_1100,N_516);
nand U4079 (N_4079,N_1373,N_2370);
or U4080 (N_4080,N_921,N_1431);
and U4081 (N_4081,N_788,N_895);
nor U4082 (N_4082,N_2267,N_1086);
nand U4083 (N_4083,N_649,N_1736);
nor U4084 (N_4084,N_595,N_1507);
nand U4085 (N_4085,N_1458,N_465);
or U4086 (N_4086,N_1195,N_642);
nor U4087 (N_4087,N_2219,N_2315);
and U4088 (N_4088,N_1513,N_2280);
and U4089 (N_4089,N_178,N_241);
and U4090 (N_4090,N_2399,N_1746);
nor U4091 (N_4091,N_1993,N_1035);
nor U4092 (N_4092,N_334,N_689);
xnor U4093 (N_4093,N_1736,N_1218);
nand U4094 (N_4094,N_1625,N_1477);
nor U4095 (N_4095,N_417,N_1822);
xor U4096 (N_4096,N_1295,N_1799);
and U4097 (N_4097,N_221,N_2235);
nor U4098 (N_4098,N_1449,N_2281);
or U4099 (N_4099,N_174,N_1320);
or U4100 (N_4100,N_865,N_1041);
and U4101 (N_4101,N_1177,N_1164);
xor U4102 (N_4102,N_128,N_1976);
or U4103 (N_4103,N_2129,N_1536);
xnor U4104 (N_4104,N_984,N_1634);
nand U4105 (N_4105,N_2182,N_1172);
or U4106 (N_4106,N_1028,N_2440);
xor U4107 (N_4107,N_1867,N_1764);
and U4108 (N_4108,N_1952,N_423);
xnor U4109 (N_4109,N_2233,N_1931);
or U4110 (N_4110,N_1111,N_360);
nand U4111 (N_4111,N_1647,N_1087);
nand U4112 (N_4112,N_161,N_2095);
nor U4113 (N_4113,N_2340,N_309);
or U4114 (N_4114,N_1521,N_2439);
xor U4115 (N_4115,N_1513,N_2418);
and U4116 (N_4116,N_955,N_1349);
and U4117 (N_4117,N_41,N_2313);
or U4118 (N_4118,N_2291,N_2145);
nor U4119 (N_4119,N_98,N_1464);
nand U4120 (N_4120,N_1726,N_1024);
or U4121 (N_4121,N_2235,N_422);
nand U4122 (N_4122,N_1017,N_824);
or U4123 (N_4123,N_1842,N_1389);
nand U4124 (N_4124,N_2251,N_1538);
nand U4125 (N_4125,N_807,N_19);
or U4126 (N_4126,N_1380,N_2117);
nand U4127 (N_4127,N_236,N_2075);
xor U4128 (N_4128,N_630,N_1102);
nand U4129 (N_4129,N_952,N_1593);
nor U4130 (N_4130,N_1045,N_2210);
nor U4131 (N_4131,N_30,N_1718);
and U4132 (N_4132,N_1228,N_1738);
nand U4133 (N_4133,N_398,N_324);
xor U4134 (N_4134,N_791,N_243);
nor U4135 (N_4135,N_1407,N_567);
xnor U4136 (N_4136,N_2463,N_762);
and U4137 (N_4137,N_1538,N_1332);
nand U4138 (N_4138,N_2022,N_451);
xor U4139 (N_4139,N_2087,N_859);
xor U4140 (N_4140,N_1840,N_299);
nor U4141 (N_4141,N_1259,N_1195);
or U4142 (N_4142,N_726,N_824);
and U4143 (N_4143,N_1847,N_757);
nand U4144 (N_4144,N_1823,N_1277);
xnor U4145 (N_4145,N_66,N_900);
and U4146 (N_4146,N_251,N_1566);
and U4147 (N_4147,N_1766,N_2286);
or U4148 (N_4148,N_1716,N_2004);
nand U4149 (N_4149,N_616,N_1788);
or U4150 (N_4150,N_2374,N_1195);
nand U4151 (N_4151,N_918,N_1360);
nand U4152 (N_4152,N_334,N_1309);
and U4153 (N_4153,N_1057,N_1512);
nand U4154 (N_4154,N_2148,N_2480);
or U4155 (N_4155,N_1657,N_1041);
nand U4156 (N_4156,N_1610,N_903);
and U4157 (N_4157,N_151,N_783);
xor U4158 (N_4158,N_1022,N_1843);
nor U4159 (N_4159,N_1188,N_2060);
nand U4160 (N_4160,N_503,N_1169);
or U4161 (N_4161,N_2072,N_1050);
xor U4162 (N_4162,N_2014,N_2314);
nand U4163 (N_4163,N_1702,N_1162);
nor U4164 (N_4164,N_960,N_262);
or U4165 (N_4165,N_1799,N_541);
xor U4166 (N_4166,N_1710,N_1750);
and U4167 (N_4167,N_2483,N_1800);
or U4168 (N_4168,N_276,N_98);
and U4169 (N_4169,N_955,N_1257);
nand U4170 (N_4170,N_1102,N_968);
nand U4171 (N_4171,N_604,N_1744);
nor U4172 (N_4172,N_1332,N_1467);
or U4173 (N_4173,N_1566,N_656);
and U4174 (N_4174,N_1713,N_2158);
xnor U4175 (N_4175,N_1898,N_1450);
nor U4176 (N_4176,N_1620,N_522);
nor U4177 (N_4177,N_731,N_2409);
or U4178 (N_4178,N_518,N_2150);
nor U4179 (N_4179,N_562,N_1059);
nor U4180 (N_4180,N_253,N_1668);
nor U4181 (N_4181,N_778,N_1016);
nor U4182 (N_4182,N_1734,N_1621);
and U4183 (N_4183,N_1227,N_579);
or U4184 (N_4184,N_315,N_1092);
and U4185 (N_4185,N_1180,N_923);
nand U4186 (N_4186,N_518,N_886);
or U4187 (N_4187,N_529,N_1637);
or U4188 (N_4188,N_517,N_602);
nor U4189 (N_4189,N_965,N_292);
nand U4190 (N_4190,N_1722,N_1493);
and U4191 (N_4191,N_1789,N_1229);
nand U4192 (N_4192,N_2449,N_2169);
nand U4193 (N_4193,N_56,N_1476);
xnor U4194 (N_4194,N_192,N_1673);
xnor U4195 (N_4195,N_1000,N_1191);
nand U4196 (N_4196,N_1026,N_2481);
and U4197 (N_4197,N_1109,N_1011);
nand U4198 (N_4198,N_1754,N_150);
and U4199 (N_4199,N_2236,N_571);
or U4200 (N_4200,N_1826,N_56);
and U4201 (N_4201,N_2097,N_1231);
nand U4202 (N_4202,N_558,N_1988);
and U4203 (N_4203,N_2247,N_1075);
or U4204 (N_4204,N_1282,N_1416);
or U4205 (N_4205,N_2391,N_39);
xnor U4206 (N_4206,N_2216,N_2173);
or U4207 (N_4207,N_1273,N_1598);
nor U4208 (N_4208,N_1239,N_2410);
xor U4209 (N_4209,N_325,N_2231);
nand U4210 (N_4210,N_1363,N_1731);
nor U4211 (N_4211,N_180,N_814);
or U4212 (N_4212,N_1466,N_1467);
nor U4213 (N_4213,N_2284,N_1796);
and U4214 (N_4214,N_631,N_1339);
and U4215 (N_4215,N_1336,N_96);
or U4216 (N_4216,N_1413,N_2265);
and U4217 (N_4217,N_39,N_1117);
xnor U4218 (N_4218,N_987,N_2284);
and U4219 (N_4219,N_1620,N_2040);
and U4220 (N_4220,N_1585,N_2238);
nand U4221 (N_4221,N_141,N_1125);
xor U4222 (N_4222,N_526,N_174);
or U4223 (N_4223,N_2402,N_630);
xor U4224 (N_4224,N_2490,N_72);
or U4225 (N_4225,N_24,N_635);
nor U4226 (N_4226,N_927,N_32);
or U4227 (N_4227,N_299,N_2063);
nand U4228 (N_4228,N_1473,N_1911);
xnor U4229 (N_4229,N_1101,N_1752);
xnor U4230 (N_4230,N_1577,N_246);
xor U4231 (N_4231,N_606,N_2250);
or U4232 (N_4232,N_1973,N_2019);
xor U4233 (N_4233,N_415,N_626);
or U4234 (N_4234,N_1096,N_41);
nand U4235 (N_4235,N_2041,N_846);
or U4236 (N_4236,N_685,N_761);
nor U4237 (N_4237,N_839,N_1453);
or U4238 (N_4238,N_2030,N_657);
nor U4239 (N_4239,N_990,N_853);
and U4240 (N_4240,N_2179,N_483);
xor U4241 (N_4241,N_308,N_2306);
and U4242 (N_4242,N_1108,N_855);
xor U4243 (N_4243,N_748,N_1314);
or U4244 (N_4244,N_1608,N_699);
xnor U4245 (N_4245,N_611,N_307);
nor U4246 (N_4246,N_2259,N_1234);
nand U4247 (N_4247,N_272,N_1061);
nand U4248 (N_4248,N_360,N_800);
nor U4249 (N_4249,N_678,N_1047);
and U4250 (N_4250,N_748,N_1454);
xnor U4251 (N_4251,N_1775,N_2372);
or U4252 (N_4252,N_273,N_1207);
and U4253 (N_4253,N_99,N_2390);
xor U4254 (N_4254,N_625,N_1192);
and U4255 (N_4255,N_2059,N_2013);
xnor U4256 (N_4256,N_197,N_209);
nand U4257 (N_4257,N_2065,N_214);
or U4258 (N_4258,N_1407,N_527);
nor U4259 (N_4259,N_1262,N_2027);
nor U4260 (N_4260,N_1488,N_2021);
and U4261 (N_4261,N_1842,N_2081);
and U4262 (N_4262,N_1768,N_381);
nor U4263 (N_4263,N_839,N_2493);
and U4264 (N_4264,N_1982,N_633);
nand U4265 (N_4265,N_2346,N_818);
nor U4266 (N_4266,N_433,N_159);
or U4267 (N_4267,N_1132,N_1113);
and U4268 (N_4268,N_1358,N_161);
nor U4269 (N_4269,N_626,N_875);
or U4270 (N_4270,N_357,N_817);
or U4271 (N_4271,N_1334,N_388);
and U4272 (N_4272,N_1796,N_1920);
or U4273 (N_4273,N_909,N_461);
xor U4274 (N_4274,N_1096,N_1141);
nand U4275 (N_4275,N_624,N_797);
and U4276 (N_4276,N_724,N_51);
nand U4277 (N_4277,N_1290,N_1704);
or U4278 (N_4278,N_1272,N_892);
and U4279 (N_4279,N_2397,N_1907);
nand U4280 (N_4280,N_2175,N_1472);
xnor U4281 (N_4281,N_2303,N_1512);
or U4282 (N_4282,N_1439,N_2227);
or U4283 (N_4283,N_1669,N_40);
or U4284 (N_4284,N_2302,N_667);
nand U4285 (N_4285,N_2085,N_2253);
xor U4286 (N_4286,N_230,N_1639);
nand U4287 (N_4287,N_1498,N_171);
xnor U4288 (N_4288,N_860,N_2078);
and U4289 (N_4289,N_1439,N_1882);
or U4290 (N_4290,N_1715,N_79);
nor U4291 (N_4291,N_1508,N_1322);
or U4292 (N_4292,N_2266,N_561);
xnor U4293 (N_4293,N_2120,N_731);
or U4294 (N_4294,N_2226,N_1244);
nand U4295 (N_4295,N_1041,N_2120);
or U4296 (N_4296,N_1717,N_1736);
or U4297 (N_4297,N_2455,N_623);
or U4298 (N_4298,N_616,N_1355);
xor U4299 (N_4299,N_487,N_163);
nor U4300 (N_4300,N_662,N_202);
nand U4301 (N_4301,N_2185,N_1190);
or U4302 (N_4302,N_1512,N_633);
or U4303 (N_4303,N_1075,N_2167);
xnor U4304 (N_4304,N_1598,N_1572);
xor U4305 (N_4305,N_262,N_2121);
and U4306 (N_4306,N_180,N_373);
and U4307 (N_4307,N_844,N_1489);
or U4308 (N_4308,N_1415,N_2455);
and U4309 (N_4309,N_1252,N_882);
or U4310 (N_4310,N_146,N_242);
and U4311 (N_4311,N_361,N_2281);
and U4312 (N_4312,N_340,N_1705);
nand U4313 (N_4313,N_2039,N_2034);
nand U4314 (N_4314,N_1255,N_1268);
and U4315 (N_4315,N_493,N_608);
nor U4316 (N_4316,N_338,N_2457);
xnor U4317 (N_4317,N_2342,N_2036);
and U4318 (N_4318,N_869,N_927);
and U4319 (N_4319,N_2163,N_1394);
nor U4320 (N_4320,N_1053,N_1708);
and U4321 (N_4321,N_1241,N_965);
and U4322 (N_4322,N_727,N_2014);
nand U4323 (N_4323,N_1806,N_1344);
nor U4324 (N_4324,N_1877,N_1643);
xor U4325 (N_4325,N_1711,N_1374);
nor U4326 (N_4326,N_744,N_1206);
or U4327 (N_4327,N_1317,N_2009);
nor U4328 (N_4328,N_2212,N_1667);
and U4329 (N_4329,N_1008,N_251);
or U4330 (N_4330,N_2375,N_1429);
nor U4331 (N_4331,N_1453,N_991);
xor U4332 (N_4332,N_1789,N_1478);
xnor U4333 (N_4333,N_1903,N_793);
or U4334 (N_4334,N_901,N_1094);
xor U4335 (N_4335,N_233,N_811);
and U4336 (N_4336,N_1256,N_2075);
and U4337 (N_4337,N_2033,N_1644);
nand U4338 (N_4338,N_87,N_507);
xnor U4339 (N_4339,N_1326,N_2194);
xnor U4340 (N_4340,N_606,N_306);
or U4341 (N_4341,N_1947,N_2256);
or U4342 (N_4342,N_1635,N_715);
and U4343 (N_4343,N_233,N_345);
nor U4344 (N_4344,N_1831,N_1518);
nor U4345 (N_4345,N_1327,N_509);
nand U4346 (N_4346,N_7,N_1960);
or U4347 (N_4347,N_2268,N_37);
nor U4348 (N_4348,N_1357,N_933);
nor U4349 (N_4349,N_1273,N_1268);
or U4350 (N_4350,N_104,N_633);
nand U4351 (N_4351,N_1777,N_1682);
and U4352 (N_4352,N_546,N_1607);
nand U4353 (N_4353,N_1397,N_2201);
or U4354 (N_4354,N_2386,N_2020);
nor U4355 (N_4355,N_2457,N_1724);
xor U4356 (N_4356,N_365,N_743);
xnor U4357 (N_4357,N_67,N_764);
xnor U4358 (N_4358,N_1946,N_505);
xnor U4359 (N_4359,N_1173,N_2320);
nand U4360 (N_4360,N_714,N_1903);
nand U4361 (N_4361,N_1012,N_1427);
or U4362 (N_4362,N_1635,N_828);
or U4363 (N_4363,N_1824,N_640);
and U4364 (N_4364,N_715,N_605);
and U4365 (N_4365,N_1619,N_1725);
or U4366 (N_4366,N_1733,N_1912);
nand U4367 (N_4367,N_1458,N_1666);
xnor U4368 (N_4368,N_1974,N_1412);
nand U4369 (N_4369,N_2054,N_1108);
or U4370 (N_4370,N_1250,N_1856);
and U4371 (N_4371,N_74,N_354);
xnor U4372 (N_4372,N_63,N_2024);
xor U4373 (N_4373,N_1820,N_949);
and U4374 (N_4374,N_2347,N_917);
or U4375 (N_4375,N_443,N_1580);
and U4376 (N_4376,N_21,N_549);
or U4377 (N_4377,N_806,N_2377);
nor U4378 (N_4378,N_1418,N_1697);
nand U4379 (N_4379,N_2290,N_499);
nor U4380 (N_4380,N_808,N_1378);
or U4381 (N_4381,N_1154,N_1446);
or U4382 (N_4382,N_1856,N_1490);
xor U4383 (N_4383,N_1365,N_2362);
nand U4384 (N_4384,N_390,N_150);
and U4385 (N_4385,N_2139,N_1719);
xor U4386 (N_4386,N_2338,N_1755);
or U4387 (N_4387,N_1466,N_632);
nand U4388 (N_4388,N_1869,N_962);
and U4389 (N_4389,N_496,N_943);
and U4390 (N_4390,N_1852,N_1611);
nand U4391 (N_4391,N_1431,N_1745);
or U4392 (N_4392,N_1942,N_398);
xnor U4393 (N_4393,N_1814,N_795);
nand U4394 (N_4394,N_2284,N_1027);
or U4395 (N_4395,N_752,N_1932);
nand U4396 (N_4396,N_2378,N_1874);
xnor U4397 (N_4397,N_1145,N_2336);
and U4398 (N_4398,N_2016,N_1155);
nand U4399 (N_4399,N_2181,N_2108);
nand U4400 (N_4400,N_5,N_1899);
nor U4401 (N_4401,N_777,N_1137);
or U4402 (N_4402,N_130,N_1587);
nor U4403 (N_4403,N_686,N_194);
xor U4404 (N_4404,N_1377,N_1137);
and U4405 (N_4405,N_1631,N_772);
and U4406 (N_4406,N_1877,N_321);
and U4407 (N_4407,N_378,N_2179);
and U4408 (N_4408,N_2348,N_13);
nand U4409 (N_4409,N_1878,N_2431);
nand U4410 (N_4410,N_1156,N_145);
xnor U4411 (N_4411,N_31,N_558);
xor U4412 (N_4412,N_387,N_938);
and U4413 (N_4413,N_476,N_1149);
xor U4414 (N_4414,N_1485,N_98);
nor U4415 (N_4415,N_559,N_1938);
xnor U4416 (N_4416,N_207,N_1427);
or U4417 (N_4417,N_1899,N_739);
xnor U4418 (N_4418,N_2178,N_606);
xor U4419 (N_4419,N_1562,N_185);
and U4420 (N_4420,N_1903,N_271);
nor U4421 (N_4421,N_2434,N_1040);
or U4422 (N_4422,N_893,N_574);
nand U4423 (N_4423,N_2327,N_2360);
nand U4424 (N_4424,N_1691,N_1097);
nand U4425 (N_4425,N_2124,N_1057);
or U4426 (N_4426,N_327,N_2326);
or U4427 (N_4427,N_401,N_17);
nor U4428 (N_4428,N_1578,N_462);
or U4429 (N_4429,N_1759,N_186);
nand U4430 (N_4430,N_1513,N_495);
nor U4431 (N_4431,N_184,N_2324);
and U4432 (N_4432,N_93,N_383);
or U4433 (N_4433,N_1965,N_639);
xor U4434 (N_4434,N_1413,N_2351);
and U4435 (N_4435,N_625,N_430);
or U4436 (N_4436,N_2059,N_762);
and U4437 (N_4437,N_1271,N_1811);
nor U4438 (N_4438,N_774,N_1514);
xnor U4439 (N_4439,N_1470,N_2297);
and U4440 (N_4440,N_400,N_901);
and U4441 (N_4441,N_171,N_2006);
and U4442 (N_4442,N_1108,N_2006);
or U4443 (N_4443,N_1139,N_652);
nand U4444 (N_4444,N_39,N_1196);
or U4445 (N_4445,N_1721,N_1599);
and U4446 (N_4446,N_639,N_633);
xor U4447 (N_4447,N_1681,N_1558);
or U4448 (N_4448,N_2379,N_754);
and U4449 (N_4449,N_557,N_119);
and U4450 (N_4450,N_1036,N_1815);
nor U4451 (N_4451,N_1702,N_1199);
nor U4452 (N_4452,N_379,N_2010);
nor U4453 (N_4453,N_610,N_897);
nor U4454 (N_4454,N_2050,N_828);
nand U4455 (N_4455,N_1292,N_1722);
xnor U4456 (N_4456,N_1638,N_439);
or U4457 (N_4457,N_1205,N_1538);
and U4458 (N_4458,N_2401,N_2405);
xor U4459 (N_4459,N_2445,N_334);
and U4460 (N_4460,N_1079,N_204);
nand U4461 (N_4461,N_1917,N_2338);
or U4462 (N_4462,N_2063,N_395);
or U4463 (N_4463,N_189,N_2254);
nor U4464 (N_4464,N_1168,N_807);
nand U4465 (N_4465,N_2073,N_2358);
nand U4466 (N_4466,N_574,N_2138);
nand U4467 (N_4467,N_168,N_966);
nor U4468 (N_4468,N_652,N_498);
and U4469 (N_4469,N_857,N_1352);
xnor U4470 (N_4470,N_1634,N_310);
nor U4471 (N_4471,N_682,N_2082);
and U4472 (N_4472,N_734,N_1585);
nor U4473 (N_4473,N_2169,N_469);
nand U4474 (N_4474,N_1593,N_1657);
or U4475 (N_4475,N_330,N_1708);
or U4476 (N_4476,N_1308,N_1386);
or U4477 (N_4477,N_1573,N_2298);
xnor U4478 (N_4478,N_1728,N_883);
nor U4479 (N_4479,N_837,N_809);
nand U4480 (N_4480,N_1131,N_1631);
nand U4481 (N_4481,N_2273,N_335);
nor U4482 (N_4482,N_1336,N_259);
xnor U4483 (N_4483,N_2158,N_935);
and U4484 (N_4484,N_2194,N_1024);
nand U4485 (N_4485,N_1773,N_1064);
xnor U4486 (N_4486,N_2345,N_554);
nor U4487 (N_4487,N_772,N_797);
xor U4488 (N_4488,N_1899,N_1263);
and U4489 (N_4489,N_1144,N_1687);
xor U4490 (N_4490,N_333,N_70);
and U4491 (N_4491,N_1966,N_298);
nand U4492 (N_4492,N_235,N_1556);
xnor U4493 (N_4493,N_1034,N_2194);
and U4494 (N_4494,N_2220,N_868);
and U4495 (N_4495,N_1538,N_1527);
nor U4496 (N_4496,N_1375,N_2133);
nor U4497 (N_4497,N_1424,N_2334);
and U4498 (N_4498,N_561,N_630);
or U4499 (N_4499,N_401,N_67);
xnor U4500 (N_4500,N_689,N_827);
and U4501 (N_4501,N_1612,N_477);
xnor U4502 (N_4502,N_1021,N_2065);
or U4503 (N_4503,N_1094,N_329);
or U4504 (N_4504,N_1125,N_1211);
and U4505 (N_4505,N_407,N_1123);
nand U4506 (N_4506,N_616,N_1499);
and U4507 (N_4507,N_1902,N_938);
or U4508 (N_4508,N_2464,N_300);
nor U4509 (N_4509,N_1790,N_1075);
and U4510 (N_4510,N_315,N_784);
and U4511 (N_4511,N_2133,N_2348);
or U4512 (N_4512,N_87,N_2231);
or U4513 (N_4513,N_502,N_1784);
and U4514 (N_4514,N_143,N_2233);
xor U4515 (N_4515,N_870,N_1011);
or U4516 (N_4516,N_942,N_1427);
xor U4517 (N_4517,N_2056,N_1396);
and U4518 (N_4518,N_239,N_1510);
and U4519 (N_4519,N_454,N_1964);
or U4520 (N_4520,N_1173,N_1703);
nor U4521 (N_4521,N_507,N_469);
nor U4522 (N_4522,N_511,N_2268);
xor U4523 (N_4523,N_1582,N_330);
xor U4524 (N_4524,N_570,N_2096);
and U4525 (N_4525,N_1169,N_1540);
or U4526 (N_4526,N_1642,N_677);
xor U4527 (N_4527,N_2049,N_1138);
nand U4528 (N_4528,N_84,N_1502);
xor U4529 (N_4529,N_1748,N_193);
nand U4530 (N_4530,N_2327,N_996);
or U4531 (N_4531,N_594,N_1925);
nor U4532 (N_4532,N_781,N_1185);
and U4533 (N_4533,N_1490,N_712);
nor U4534 (N_4534,N_1098,N_1425);
xnor U4535 (N_4535,N_2006,N_736);
xor U4536 (N_4536,N_433,N_929);
nand U4537 (N_4537,N_1620,N_104);
xor U4538 (N_4538,N_1368,N_2237);
xor U4539 (N_4539,N_1077,N_759);
nor U4540 (N_4540,N_2070,N_2196);
nor U4541 (N_4541,N_1427,N_120);
nor U4542 (N_4542,N_802,N_1854);
xor U4543 (N_4543,N_1888,N_2377);
nor U4544 (N_4544,N_2497,N_175);
and U4545 (N_4545,N_1654,N_2423);
or U4546 (N_4546,N_808,N_2104);
nand U4547 (N_4547,N_1527,N_1685);
nand U4548 (N_4548,N_46,N_425);
xor U4549 (N_4549,N_833,N_955);
nand U4550 (N_4550,N_85,N_1363);
and U4551 (N_4551,N_2254,N_42);
or U4552 (N_4552,N_1536,N_2115);
or U4553 (N_4553,N_2289,N_157);
or U4554 (N_4554,N_2378,N_16);
xnor U4555 (N_4555,N_966,N_2041);
or U4556 (N_4556,N_779,N_1060);
nand U4557 (N_4557,N_1756,N_2445);
and U4558 (N_4558,N_1507,N_952);
and U4559 (N_4559,N_2210,N_2001);
nor U4560 (N_4560,N_2125,N_1878);
nor U4561 (N_4561,N_2038,N_318);
xor U4562 (N_4562,N_290,N_2264);
nor U4563 (N_4563,N_456,N_542);
nor U4564 (N_4564,N_2171,N_2339);
or U4565 (N_4565,N_1371,N_1945);
nand U4566 (N_4566,N_1811,N_1440);
and U4567 (N_4567,N_868,N_252);
or U4568 (N_4568,N_141,N_1891);
nor U4569 (N_4569,N_1867,N_1930);
and U4570 (N_4570,N_687,N_866);
and U4571 (N_4571,N_1513,N_1836);
nor U4572 (N_4572,N_285,N_653);
nand U4573 (N_4573,N_2099,N_1515);
and U4574 (N_4574,N_899,N_2341);
or U4575 (N_4575,N_417,N_20);
or U4576 (N_4576,N_2466,N_150);
nand U4577 (N_4577,N_1180,N_2265);
nand U4578 (N_4578,N_954,N_1924);
nand U4579 (N_4579,N_1957,N_556);
and U4580 (N_4580,N_432,N_649);
nor U4581 (N_4581,N_1645,N_1411);
xor U4582 (N_4582,N_1604,N_1458);
nor U4583 (N_4583,N_334,N_609);
xor U4584 (N_4584,N_195,N_356);
or U4585 (N_4585,N_678,N_1671);
xnor U4586 (N_4586,N_390,N_1644);
or U4587 (N_4587,N_1306,N_184);
xnor U4588 (N_4588,N_1505,N_1646);
nand U4589 (N_4589,N_2321,N_922);
nand U4590 (N_4590,N_552,N_1853);
or U4591 (N_4591,N_316,N_765);
or U4592 (N_4592,N_1238,N_2108);
and U4593 (N_4593,N_1723,N_131);
nand U4594 (N_4594,N_1455,N_2132);
xor U4595 (N_4595,N_420,N_616);
nand U4596 (N_4596,N_2389,N_699);
and U4597 (N_4597,N_1736,N_437);
xnor U4598 (N_4598,N_1941,N_1148);
nor U4599 (N_4599,N_805,N_1812);
and U4600 (N_4600,N_2306,N_1372);
xor U4601 (N_4601,N_209,N_1782);
nor U4602 (N_4602,N_1283,N_1296);
nor U4603 (N_4603,N_730,N_2495);
xnor U4604 (N_4604,N_1184,N_1631);
xnor U4605 (N_4605,N_1542,N_844);
xnor U4606 (N_4606,N_2446,N_1460);
nor U4607 (N_4607,N_1931,N_1317);
or U4608 (N_4608,N_1883,N_433);
or U4609 (N_4609,N_232,N_1497);
or U4610 (N_4610,N_2402,N_369);
nand U4611 (N_4611,N_1825,N_1266);
nand U4612 (N_4612,N_299,N_1936);
or U4613 (N_4613,N_1320,N_327);
and U4614 (N_4614,N_2435,N_1147);
nand U4615 (N_4615,N_1482,N_1713);
xor U4616 (N_4616,N_1461,N_2244);
or U4617 (N_4617,N_1734,N_1288);
nand U4618 (N_4618,N_402,N_566);
or U4619 (N_4619,N_1395,N_1724);
nor U4620 (N_4620,N_1536,N_1401);
xor U4621 (N_4621,N_1420,N_1190);
or U4622 (N_4622,N_1990,N_253);
and U4623 (N_4623,N_2375,N_1479);
xor U4624 (N_4624,N_1882,N_1487);
xnor U4625 (N_4625,N_67,N_1939);
and U4626 (N_4626,N_2426,N_1614);
nor U4627 (N_4627,N_629,N_1945);
nand U4628 (N_4628,N_1905,N_1204);
xor U4629 (N_4629,N_1994,N_2069);
and U4630 (N_4630,N_1091,N_1690);
or U4631 (N_4631,N_1807,N_1073);
nand U4632 (N_4632,N_1838,N_45);
nand U4633 (N_4633,N_683,N_885);
nand U4634 (N_4634,N_422,N_25);
and U4635 (N_4635,N_389,N_2243);
xor U4636 (N_4636,N_1155,N_2178);
and U4637 (N_4637,N_1074,N_1644);
nor U4638 (N_4638,N_1854,N_422);
and U4639 (N_4639,N_2110,N_1070);
xnor U4640 (N_4640,N_31,N_2169);
nand U4641 (N_4641,N_201,N_485);
xor U4642 (N_4642,N_1332,N_77);
nand U4643 (N_4643,N_1565,N_503);
nand U4644 (N_4644,N_2261,N_714);
nor U4645 (N_4645,N_647,N_1467);
xor U4646 (N_4646,N_1743,N_950);
and U4647 (N_4647,N_784,N_1757);
nand U4648 (N_4648,N_1080,N_51);
xnor U4649 (N_4649,N_1428,N_1915);
nand U4650 (N_4650,N_643,N_1055);
xor U4651 (N_4651,N_23,N_849);
nand U4652 (N_4652,N_2333,N_95);
and U4653 (N_4653,N_1310,N_1391);
xor U4654 (N_4654,N_207,N_99);
or U4655 (N_4655,N_399,N_1914);
nor U4656 (N_4656,N_2378,N_1061);
xnor U4657 (N_4657,N_1384,N_1163);
nor U4658 (N_4658,N_847,N_827);
xnor U4659 (N_4659,N_1190,N_1121);
nand U4660 (N_4660,N_559,N_1720);
and U4661 (N_4661,N_1590,N_1950);
and U4662 (N_4662,N_1487,N_2038);
and U4663 (N_4663,N_72,N_1909);
or U4664 (N_4664,N_1887,N_1260);
and U4665 (N_4665,N_2019,N_1468);
xnor U4666 (N_4666,N_1984,N_2308);
nor U4667 (N_4667,N_1839,N_796);
or U4668 (N_4668,N_675,N_2272);
or U4669 (N_4669,N_2295,N_2073);
nor U4670 (N_4670,N_1957,N_1068);
xnor U4671 (N_4671,N_2073,N_1302);
xor U4672 (N_4672,N_1413,N_1101);
nor U4673 (N_4673,N_1138,N_1652);
nand U4674 (N_4674,N_53,N_1796);
nor U4675 (N_4675,N_1242,N_545);
nor U4676 (N_4676,N_1769,N_521);
or U4677 (N_4677,N_2278,N_1622);
or U4678 (N_4678,N_215,N_334);
or U4679 (N_4679,N_1605,N_2305);
and U4680 (N_4680,N_1757,N_196);
or U4681 (N_4681,N_1568,N_1848);
and U4682 (N_4682,N_2458,N_1910);
xor U4683 (N_4683,N_756,N_548);
nand U4684 (N_4684,N_2101,N_677);
nand U4685 (N_4685,N_892,N_129);
nor U4686 (N_4686,N_716,N_229);
nand U4687 (N_4687,N_1390,N_2058);
or U4688 (N_4688,N_1095,N_887);
xor U4689 (N_4689,N_2108,N_648);
xor U4690 (N_4690,N_2156,N_1379);
and U4691 (N_4691,N_1137,N_239);
and U4692 (N_4692,N_925,N_2159);
or U4693 (N_4693,N_2298,N_2148);
and U4694 (N_4694,N_2062,N_1487);
nand U4695 (N_4695,N_577,N_866);
xor U4696 (N_4696,N_1634,N_975);
nor U4697 (N_4697,N_1903,N_1615);
xnor U4698 (N_4698,N_2001,N_122);
nor U4699 (N_4699,N_376,N_14);
nor U4700 (N_4700,N_1910,N_681);
nand U4701 (N_4701,N_1079,N_2124);
xnor U4702 (N_4702,N_444,N_86);
or U4703 (N_4703,N_433,N_104);
xor U4704 (N_4704,N_4,N_1246);
nand U4705 (N_4705,N_1101,N_2244);
and U4706 (N_4706,N_2344,N_1035);
or U4707 (N_4707,N_1197,N_135);
or U4708 (N_4708,N_350,N_1204);
and U4709 (N_4709,N_2148,N_1785);
or U4710 (N_4710,N_2377,N_2286);
nor U4711 (N_4711,N_2256,N_970);
nor U4712 (N_4712,N_2104,N_1671);
or U4713 (N_4713,N_1950,N_774);
xnor U4714 (N_4714,N_1456,N_994);
nand U4715 (N_4715,N_1776,N_1346);
nand U4716 (N_4716,N_929,N_612);
xor U4717 (N_4717,N_1395,N_1745);
nand U4718 (N_4718,N_1780,N_1916);
or U4719 (N_4719,N_88,N_1338);
or U4720 (N_4720,N_1630,N_281);
nor U4721 (N_4721,N_554,N_2390);
and U4722 (N_4722,N_122,N_844);
xor U4723 (N_4723,N_742,N_445);
nor U4724 (N_4724,N_5,N_1781);
nand U4725 (N_4725,N_1191,N_2166);
or U4726 (N_4726,N_32,N_1856);
xor U4727 (N_4727,N_2428,N_1660);
xor U4728 (N_4728,N_1459,N_1624);
or U4729 (N_4729,N_1908,N_1401);
xnor U4730 (N_4730,N_1450,N_356);
nand U4731 (N_4731,N_1140,N_545);
nor U4732 (N_4732,N_2084,N_2319);
xor U4733 (N_4733,N_1960,N_620);
xnor U4734 (N_4734,N_489,N_385);
or U4735 (N_4735,N_2101,N_1393);
nor U4736 (N_4736,N_747,N_641);
nor U4737 (N_4737,N_2193,N_1505);
nor U4738 (N_4738,N_45,N_1429);
xor U4739 (N_4739,N_1439,N_478);
nor U4740 (N_4740,N_376,N_2006);
xor U4741 (N_4741,N_2224,N_2091);
or U4742 (N_4742,N_81,N_286);
xor U4743 (N_4743,N_1753,N_554);
or U4744 (N_4744,N_1220,N_2402);
nor U4745 (N_4745,N_2244,N_941);
and U4746 (N_4746,N_2300,N_1027);
or U4747 (N_4747,N_370,N_1199);
xnor U4748 (N_4748,N_1477,N_1168);
or U4749 (N_4749,N_1832,N_1998);
xnor U4750 (N_4750,N_2055,N_1378);
nand U4751 (N_4751,N_672,N_1458);
and U4752 (N_4752,N_75,N_2033);
and U4753 (N_4753,N_990,N_1564);
nand U4754 (N_4754,N_70,N_235);
nand U4755 (N_4755,N_1208,N_455);
or U4756 (N_4756,N_939,N_1116);
nand U4757 (N_4757,N_1501,N_1378);
nand U4758 (N_4758,N_956,N_1725);
and U4759 (N_4759,N_432,N_945);
nor U4760 (N_4760,N_1667,N_614);
xnor U4761 (N_4761,N_1100,N_951);
xor U4762 (N_4762,N_284,N_2052);
xor U4763 (N_4763,N_38,N_2426);
or U4764 (N_4764,N_1241,N_1133);
or U4765 (N_4765,N_2363,N_488);
nor U4766 (N_4766,N_1433,N_1558);
nand U4767 (N_4767,N_1302,N_943);
and U4768 (N_4768,N_1351,N_673);
nor U4769 (N_4769,N_1158,N_1548);
xor U4770 (N_4770,N_2161,N_1353);
or U4771 (N_4771,N_1172,N_1346);
and U4772 (N_4772,N_536,N_1396);
nor U4773 (N_4773,N_1060,N_1728);
xnor U4774 (N_4774,N_778,N_1249);
and U4775 (N_4775,N_1063,N_545);
or U4776 (N_4776,N_54,N_1644);
xor U4777 (N_4777,N_310,N_19);
nor U4778 (N_4778,N_1848,N_1551);
nor U4779 (N_4779,N_399,N_1953);
xor U4780 (N_4780,N_1285,N_877);
nand U4781 (N_4781,N_396,N_412);
and U4782 (N_4782,N_1702,N_2356);
nor U4783 (N_4783,N_2253,N_125);
or U4784 (N_4784,N_352,N_1303);
xnor U4785 (N_4785,N_882,N_563);
nand U4786 (N_4786,N_2495,N_1766);
and U4787 (N_4787,N_885,N_2117);
or U4788 (N_4788,N_1235,N_2046);
nand U4789 (N_4789,N_996,N_983);
nor U4790 (N_4790,N_1208,N_587);
nor U4791 (N_4791,N_1485,N_756);
nand U4792 (N_4792,N_627,N_790);
xor U4793 (N_4793,N_90,N_1024);
nor U4794 (N_4794,N_1391,N_915);
or U4795 (N_4795,N_646,N_1862);
xnor U4796 (N_4796,N_690,N_886);
and U4797 (N_4797,N_2425,N_1140);
nor U4798 (N_4798,N_377,N_1030);
or U4799 (N_4799,N_1651,N_398);
or U4800 (N_4800,N_1737,N_1148);
nand U4801 (N_4801,N_2369,N_1139);
and U4802 (N_4802,N_237,N_2201);
nand U4803 (N_4803,N_907,N_1066);
xor U4804 (N_4804,N_481,N_475);
and U4805 (N_4805,N_556,N_461);
xnor U4806 (N_4806,N_1201,N_743);
and U4807 (N_4807,N_183,N_2031);
xnor U4808 (N_4808,N_1990,N_2199);
nand U4809 (N_4809,N_1323,N_350);
nand U4810 (N_4810,N_1073,N_1701);
xnor U4811 (N_4811,N_659,N_1162);
or U4812 (N_4812,N_1454,N_1765);
or U4813 (N_4813,N_449,N_2049);
nand U4814 (N_4814,N_687,N_1812);
nor U4815 (N_4815,N_2037,N_2055);
xor U4816 (N_4816,N_17,N_1706);
nand U4817 (N_4817,N_1658,N_970);
nor U4818 (N_4818,N_1748,N_1507);
nor U4819 (N_4819,N_1224,N_1854);
or U4820 (N_4820,N_2145,N_101);
nor U4821 (N_4821,N_327,N_1178);
nor U4822 (N_4822,N_1436,N_334);
or U4823 (N_4823,N_747,N_1222);
and U4824 (N_4824,N_1646,N_973);
and U4825 (N_4825,N_2364,N_1831);
nor U4826 (N_4826,N_873,N_1459);
nor U4827 (N_4827,N_128,N_522);
and U4828 (N_4828,N_29,N_400);
and U4829 (N_4829,N_1806,N_1357);
nor U4830 (N_4830,N_967,N_1780);
nor U4831 (N_4831,N_1702,N_1456);
and U4832 (N_4832,N_2200,N_1173);
xor U4833 (N_4833,N_2194,N_49);
nand U4834 (N_4834,N_1129,N_348);
xor U4835 (N_4835,N_877,N_728);
nand U4836 (N_4836,N_483,N_559);
nand U4837 (N_4837,N_1426,N_1641);
and U4838 (N_4838,N_651,N_1953);
or U4839 (N_4839,N_1929,N_412);
or U4840 (N_4840,N_2031,N_133);
or U4841 (N_4841,N_499,N_1340);
nand U4842 (N_4842,N_922,N_2192);
nand U4843 (N_4843,N_2246,N_978);
and U4844 (N_4844,N_900,N_1635);
nor U4845 (N_4845,N_1354,N_1614);
or U4846 (N_4846,N_2164,N_16);
and U4847 (N_4847,N_2246,N_287);
xnor U4848 (N_4848,N_1670,N_576);
nor U4849 (N_4849,N_262,N_1319);
nand U4850 (N_4850,N_190,N_382);
and U4851 (N_4851,N_1514,N_803);
and U4852 (N_4852,N_1191,N_2373);
nand U4853 (N_4853,N_1808,N_449);
nand U4854 (N_4854,N_2020,N_564);
or U4855 (N_4855,N_1411,N_1611);
or U4856 (N_4856,N_2133,N_454);
nand U4857 (N_4857,N_1509,N_857);
nand U4858 (N_4858,N_1943,N_1419);
nand U4859 (N_4859,N_204,N_82);
nor U4860 (N_4860,N_322,N_29);
nor U4861 (N_4861,N_321,N_129);
and U4862 (N_4862,N_1126,N_1109);
nor U4863 (N_4863,N_727,N_1827);
and U4864 (N_4864,N_1949,N_48);
nand U4865 (N_4865,N_2338,N_1940);
and U4866 (N_4866,N_1117,N_1532);
and U4867 (N_4867,N_1902,N_1705);
nand U4868 (N_4868,N_1811,N_2274);
and U4869 (N_4869,N_1567,N_45);
and U4870 (N_4870,N_2207,N_1644);
nand U4871 (N_4871,N_444,N_213);
and U4872 (N_4872,N_2061,N_136);
nor U4873 (N_4873,N_1048,N_1860);
or U4874 (N_4874,N_1620,N_1851);
nand U4875 (N_4875,N_2320,N_921);
nor U4876 (N_4876,N_540,N_2114);
and U4877 (N_4877,N_1181,N_2118);
or U4878 (N_4878,N_2391,N_379);
nor U4879 (N_4879,N_305,N_1769);
and U4880 (N_4880,N_2055,N_193);
and U4881 (N_4881,N_24,N_733);
nand U4882 (N_4882,N_977,N_553);
and U4883 (N_4883,N_421,N_1788);
nand U4884 (N_4884,N_1095,N_85);
nand U4885 (N_4885,N_1029,N_2377);
or U4886 (N_4886,N_1236,N_80);
xor U4887 (N_4887,N_993,N_414);
nand U4888 (N_4888,N_1195,N_1562);
or U4889 (N_4889,N_1539,N_262);
or U4890 (N_4890,N_2129,N_1122);
xnor U4891 (N_4891,N_1391,N_339);
and U4892 (N_4892,N_108,N_1180);
nand U4893 (N_4893,N_694,N_665);
and U4894 (N_4894,N_103,N_1606);
nor U4895 (N_4895,N_2015,N_1324);
nor U4896 (N_4896,N_2369,N_9);
and U4897 (N_4897,N_2210,N_1920);
and U4898 (N_4898,N_2366,N_1290);
xnor U4899 (N_4899,N_1235,N_577);
and U4900 (N_4900,N_1301,N_1100);
nand U4901 (N_4901,N_221,N_1177);
or U4902 (N_4902,N_1830,N_481);
nor U4903 (N_4903,N_2029,N_582);
or U4904 (N_4904,N_1335,N_1866);
xnor U4905 (N_4905,N_835,N_1509);
and U4906 (N_4906,N_984,N_813);
xnor U4907 (N_4907,N_1090,N_1332);
xnor U4908 (N_4908,N_2442,N_153);
xor U4909 (N_4909,N_2420,N_2059);
nor U4910 (N_4910,N_2474,N_1243);
and U4911 (N_4911,N_1660,N_338);
nor U4912 (N_4912,N_650,N_2158);
xor U4913 (N_4913,N_603,N_1854);
nor U4914 (N_4914,N_1464,N_1380);
xor U4915 (N_4915,N_694,N_721);
and U4916 (N_4916,N_54,N_414);
or U4917 (N_4917,N_1107,N_330);
or U4918 (N_4918,N_66,N_1754);
and U4919 (N_4919,N_1285,N_2198);
xor U4920 (N_4920,N_1935,N_1749);
or U4921 (N_4921,N_1493,N_339);
or U4922 (N_4922,N_319,N_122);
and U4923 (N_4923,N_445,N_205);
xor U4924 (N_4924,N_2213,N_1962);
nor U4925 (N_4925,N_1207,N_1987);
nor U4926 (N_4926,N_2227,N_922);
or U4927 (N_4927,N_967,N_2419);
or U4928 (N_4928,N_1462,N_510);
nor U4929 (N_4929,N_2182,N_372);
xor U4930 (N_4930,N_1979,N_903);
nor U4931 (N_4931,N_1965,N_793);
xnor U4932 (N_4932,N_1779,N_607);
or U4933 (N_4933,N_584,N_2330);
and U4934 (N_4934,N_179,N_2484);
nor U4935 (N_4935,N_1837,N_651);
nor U4936 (N_4936,N_2346,N_1440);
nand U4937 (N_4937,N_2274,N_293);
xnor U4938 (N_4938,N_663,N_1481);
or U4939 (N_4939,N_1277,N_207);
nand U4940 (N_4940,N_351,N_1359);
xor U4941 (N_4941,N_833,N_662);
and U4942 (N_4942,N_1579,N_432);
and U4943 (N_4943,N_1466,N_1080);
or U4944 (N_4944,N_1343,N_983);
nor U4945 (N_4945,N_853,N_857);
nor U4946 (N_4946,N_566,N_828);
nor U4947 (N_4947,N_596,N_1281);
and U4948 (N_4948,N_393,N_982);
and U4949 (N_4949,N_2124,N_1424);
or U4950 (N_4950,N_1202,N_428);
nor U4951 (N_4951,N_1392,N_487);
nand U4952 (N_4952,N_1776,N_709);
nand U4953 (N_4953,N_2261,N_1008);
and U4954 (N_4954,N_264,N_2480);
and U4955 (N_4955,N_1169,N_1875);
or U4956 (N_4956,N_988,N_2212);
xnor U4957 (N_4957,N_1938,N_1432);
nor U4958 (N_4958,N_1075,N_2015);
xnor U4959 (N_4959,N_490,N_1151);
or U4960 (N_4960,N_65,N_1095);
and U4961 (N_4961,N_2472,N_857);
nand U4962 (N_4962,N_1904,N_573);
nor U4963 (N_4963,N_1381,N_1528);
nor U4964 (N_4964,N_753,N_628);
nor U4965 (N_4965,N_279,N_1510);
nand U4966 (N_4966,N_1558,N_365);
xnor U4967 (N_4967,N_669,N_1451);
nor U4968 (N_4968,N_1875,N_479);
and U4969 (N_4969,N_1188,N_1108);
and U4970 (N_4970,N_609,N_2404);
and U4971 (N_4971,N_146,N_1369);
nand U4972 (N_4972,N_2034,N_1352);
or U4973 (N_4973,N_1787,N_685);
or U4974 (N_4974,N_2156,N_1469);
nand U4975 (N_4975,N_1198,N_2474);
and U4976 (N_4976,N_2303,N_2361);
nand U4977 (N_4977,N_210,N_743);
and U4978 (N_4978,N_2286,N_575);
xor U4979 (N_4979,N_1492,N_1407);
nor U4980 (N_4980,N_920,N_1298);
or U4981 (N_4981,N_1545,N_1032);
and U4982 (N_4982,N_47,N_1867);
xor U4983 (N_4983,N_1394,N_2324);
and U4984 (N_4984,N_876,N_1847);
nand U4985 (N_4985,N_818,N_2209);
and U4986 (N_4986,N_1974,N_1268);
xor U4987 (N_4987,N_342,N_1413);
and U4988 (N_4988,N_1387,N_1285);
nor U4989 (N_4989,N_1793,N_575);
nand U4990 (N_4990,N_666,N_330);
nand U4991 (N_4991,N_2024,N_300);
and U4992 (N_4992,N_792,N_284);
and U4993 (N_4993,N_2410,N_1894);
nand U4994 (N_4994,N_1498,N_1683);
and U4995 (N_4995,N_2296,N_2472);
and U4996 (N_4996,N_1352,N_2439);
nand U4997 (N_4997,N_409,N_1782);
xnor U4998 (N_4998,N_2027,N_432);
xnor U4999 (N_4999,N_664,N_718);
nor UO_0 (O_0,N_3324,N_4636);
xor UO_1 (O_1,N_3680,N_3625);
and UO_2 (O_2,N_2506,N_3382);
or UO_3 (O_3,N_3774,N_3387);
and UO_4 (O_4,N_4397,N_3323);
nor UO_5 (O_5,N_3282,N_3353);
nor UO_6 (O_6,N_2627,N_3326);
nor UO_7 (O_7,N_2696,N_3294);
and UO_8 (O_8,N_3235,N_4980);
xnor UO_9 (O_9,N_3048,N_4800);
nor UO_10 (O_10,N_3844,N_3834);
nand UO_11 (O_11,N_4157,N_4297);
and UO_12 (O_12,N_2568,N_4753);
xor UO_13 (O_13,N_3371,N_3570);
nor UO_14 (O_14,N_4478,N_4952);
nor UO_15 (O_15,N_4039,N_4047);
nand UO_16 (O_16,N_2680,N_3477);
nand UO_17 (O_17,N_3116,N_4685);
and UO_18 (O_18,N_4869,N_3177);
nor UO_19 (O_19,N_3124,N_3937);
and UO_20 (O_20,N_4598,N_2537);
and UO_21 (O_21,N_4369,N_4728);
xnor UO_22 (O_22,N_2517,N_4231);
or UO_23 (O_23,N_3706,N_2853);
nand UO_24 (O_24,N_4664,N_4198);
nand UO_25 (O_25,N_2655,N_4413);
nand UO_26 (O_26,N_4816,N_3370);
and UO_27 (O_27,N_3186,N_4591);
nand UO_28 (O_28,N_2913,N_3645);
nor UO_29 (O_29,N_3474,N_4299);
nand UO_30 (O_30,N_4036,N_3101);
nand UO_31 (O_31,N_4844,N_4782);
xnor UO_32 (O_32,N_4592,N_4220);
xnor UO_33 (O_33,N_4180,N_2702);
nor UO_34 (O_34,N_3169,N_4117);
xor UO_35 (O_35,N_3160,N_3874);
nand UO_36 (O_36,N_2788,N_4549);
nor UO_37 (O_37,N_2812,N_2550);
and UO_38 (O_38,N_4038,N_4358);
xor UO_39 (O_39,N_4799,N_4519);
and UO_40 (O_40,N_3849,N_3777);
and UO_41 (O_41,N_4308,N_4775);
nand UO_42 (O_42,N_2784,N_3531);
and UO_43 (O_43,N_3610,N_3027);
and UO_44 (O_44,N_3084,N_3816);
xnor UO_45 (O_45,N_2722,N_3067);
nand UO_46 (O_46,N_3992,N_4201);
xor UO_47 (O_47,N_3858,N_3879);
nand UO_48 (O_48,N_4814,N_4565);
xor UO_49 (O_49,N_2781,N_3443);
nor UO_50 (O_50,N_3144,N_2755);
and UO_51 (O_51,N_3156,N_3217);
nor UO_52 (O_52,N_4529,N_3333);
and UO_53 (O_53,N_3063,N_3970);
or UO_54 (O_54,N_2964,N_4915);
nor UO_55 (O_55,N_4238,N_2795);
or UO_56 (O_56,N_2530,N_4524);
and UO_57 (O_57,N_3993,N_4264);
or UO_58 (O_58,N_3832,N_2629);
xnor UO_59 (O_59,N_3790,N_4935);
nor UO_60 (O_60,N_4642,N_4373);
or UO_61 (O_61,N_3907,N_3807);
nor UO_62 (O_62,N_4757,N_3032);
xnor UO_63 (O_63,N_4770,N_3737);
or UO_64 (O_64,N_3437,N_2717);
xor UO_65 (O_65,N_3801,N_4964);
and UO_66 (O_66,N_4897,N_3306);
or UO_67 (O_67,N_3327,N_4570);
and UO_68 (O_68,N_2618,N_4443);
nand UO_69 (O_69,N_4416,N_4459);
and UO_70 (O_70,N_2578,N_3936);
xor UO_71 (O_71,N_3661,N_2646);
nor UO_72 (O_72,N_4431,N_4351);
nor UO_73 (O_73,N_3930,N_2986);
and UO_74 (O_74,N_2762,N_4845);
nor UO_75 (O_75,N_2565,N_3276);
nand UO_76 (O_76,N_2871,N_3598);
nor UO_77 (O_77,N_3917,N_4355);
or UO_78 (O_78,N_3595,N_3182);
and UO_79 (O_79,N_4078,N_4994);
nand UO_80 (O_80,N_3329,N_3093);
and UO_81 (O_81,N_3722,N_4452);
xor UO_82 (O_82,N_2922,N_3753);
nand UO_83 (O_83,N_3366,N_3708);
nand UO_84 (O_84,N_3923,N_3533);
or UO_85 (O_85,N_4174,N_4244);
and UO_86 (O_86,N_3127,N_4825);
and UO_87 (O_87,N_3720,N_4925);
nor UO_88 (O_88,N_4631,N_2827);
xor UO_89 (O_89,N_3317,N_3825);
and UO_90 (O_90,N_4891,N_3361);
nand UO_91 (O_91,N_4401,N_2616);
xnor UO_92 (O_92,N_4550,N_4278);
nand UO_93 (O_93,N_4836,N_4058);
xor UO_94 (O_94,N_4634,N_4646);
nand UO_95 (O_95,N_2894,N_3108);
xnor UO_96 (O_96,N_3602,N_4583);
xor UO_97 (O_97,N_2699,N_3897);
xor UO_98 (O_98,N_4284,N_2671);
and UO_99 (O_99,N_2991,N_3931);
or UO_100 (O_100,N_4307,N_3784);
nand UO_101 (O_101,N_3668,N_4933);
xor UO_102 (O_102,N_4268,N_2713);
nor UO_103 (O_103,N_3229,N_3789);
xor UO_104 (O_104,N_2670,N_3339);
xnor UO_105 (O_105,N_4827,N_2924);
nand UO_106 (O_106,N_2636,N_4165);
or UO_107 (O_107,N_2852,N_4257);
nor UO_108 (O_108,N_4917,N_3192);
nand UO_109 (O_109,N_3519,N_4873);
or UO_110 (O_110,N_3428,N_4247);
or UO_111 (O_111,N_2841,N_4745);
nor UO_112 (O_112,N_3195,N_3877);
xor UO_113 (O_113,N_4137,N_4709);
or UO_114 (O_114,N_3113,N_3155);
xor UO_115 (O_115,N_4123,N_4807);
or UO_116 (O_116,N_3647,N_2976);
nand UO_117 (O_117,N_4118,N_3685);
nand UO_118 (O_118,N_4393,N_4637);
or UO_119 (O_119,N_4693,N_2747);
nor UO_120 (O_120,N_3848,N_3054);
nor UO_121 (O_121,N_4419,N_3138);
nor UO_122 (O_122,N_4995,N_3482);
or UO_123 (O_123,N_3337,N_3950);
and UO_124 (O_124,N_3298,N_2911);
and UO_125 (O_125,N_4894,N_4424);
nor UO_126 (O_126,N_2950,N_2849);
and UO_127 (O_127,N_2712,N_3019);
xnor UO_128 (O_128,N_2682,N_3769);
nand UO_129 (O_129,N_3004,N_3297);
or UO_130 (O_130,N_3718,N_4677);
or UO_131 (O_131,N_4436,N_3754);
nand UO_132 (O_132,N_3725,N_4846);
or UO_133 (O_133,N_4639,N_4094);
nand UO_134 (O_134,N_4199,N_4020);
xnor UO_135 (O_135,N_2697,N_3498);
nor UO_136 (O_136,N_2835,N_3886);
xor UO_137 (O_137,N_3111,N_3524);
and UO_138 (O_138,N_3660,N_3075);
and UO_139 (O_139,N_4389,N_3209);
or UO_140 (O_140,N_2608,N_3866);
nand UO_141 (O_141,N_2692,N_3977);
or UO_142 (O_142,N_4507,N_4356);
or UO_143 (O_143,N_4116,N_3176);
nand UO_144 (O_144,N_3049,N_3245);
nand UO_145 (O_145,N_2564,N_3277);
nand UO_146 (O_146,N_3433,N_3266);
nand UO_147 (O_147,N_3827,N_3133);
nand UO_148 (O_148,N_4588,N_3161);
nand UO_149 (O_149,N_2869,N_3320);
xnor UO_150 (O_150,N_2628,N_4889);
nand UO_151 (O_151,N_2933,N_2643);
nor UO_152 (O_152,N_4070,N_4054);
and UO_153 (O_153,N_4906,N_4357);
and UO_154 (O_154,N_2688,N_4148);
or UO_155 (O_155,N_3485,N_4629);
nor UO_156 (O_156,N_4699,N_2899);
nor UO_157 (O_157,N_4811,N_4970);
or UO_158 (O_158,N_4585,N_3582);
nand UO_159 (O_159,N_4331,N_4595);
nand UO_160 (O_160,N_4626,N_2555);
or UO_161 (O_161,N_4830,N_3137);
nand UO_162 (O_162,N_3379,N_4329);
or UO_163 (O_163,N_2554,N_2928);
nor UO_164 (O_164,N_2910,N_2840);
or UO_165 (O_165,N_3744,N_4888);
xor UO_166 (O_166,N_2994,N_4968);
and UO_167 (O_167,N_3928,N_4382);
nand UO_168 (O_168,N_3270,N_4154);
xor UO_169 (O_169,N_3791,N_3034);
or UO_170 (O_170,N_3682,N_3150);
and UO_171 (O_171,N_3171,N_4604);
or UO_172 (O_172,N_4795,N_4217);
or UO_173 (O_173,N_3732,N_4734);
xnor UO_174 (O_174,N_4610,N_3041);
or UO_175 (O_175,N_4105,N_2677);
xnor UO_176 (O_176,N_4212,N_3980);
xnor UO_177 (O_177,N_3525,N_2981);
nand UO_178 (O_178,N_3174,N_4805);
nand UO_179 (O_179,N_3357,N_2553);
xnor UO_180 (O_180,N_4160,N_4142);
and UO_181 (O_181,N_3035,N_2708);
nor UO_182 (O_182,N_4748,N_2740);
nand UO_183 (O_183,N_2657,N_2842);
and UO_184 (O_184,N_2557,N_2562);
nand UO_185 (O_185,N_4421,N_4542);
nand UO_186 (O_186,N_3227,N_2771);
or UO_187 (O_187,N_4143,N_4128);
or UO_188 (O_188,N_4691,N_3461);
or UO_189 (O_189,N_4887,N_2610);
nand UO_190 (O_190,N_2901,N_4527);
xor UO_191 (O_191,N_4193,N_4042);
nor UO_192 (O_192,N_4724,N_3383);
nand UO_193 (O_193,N_2728,N_4912);
xnor UO_194 (O_194,N_3069,N_4226);
xor UO_195 (O_195,N_4023,N_4092);
or UO_196 (O_196,N_4084,N_3629);
and UO_197 (O_197,N_3974,N_2513);
nand UO_198 (O_198,N_4928,N_4121);
nor UO_199 (O_199,N_4780,N_4730);
or UO_200 (O_200,N_4535,N_2949);
or UO_201 (O_201,N_2599,N_4796);
nor UO_202 (O_202,N_3142,N_4975);
nand UO_203 (O_203,N_3822,N_3143);
or UO_204 (O_204,N_3898,N_2700);
and UO_205 (O_205,N_4661,N_3164);
nor UO_206 (O_206,N_3638,N_3080);
or UO_207 (O_207,N_3652,N_3042);
nor UO_208 (O_208,N_2941,N_3766);
nand UO_209 (O_209,N_2996,N_4732);
nor UO_210 (O_210,N_3359,N_4942);
or UO_211 (O_211,N_4697,N_3441);
xor UO_212 (O_212,N_2948,N_3869);
nor UO_213 (O_213,N_4501,N_2515);
or UO_214 (O_214,N_4822,N_2760);
or UO_215 (O_215,N_2822,N_2518);
nor UO_216 (O_216,N_2510,N_2508);
or UO_217 (O_217,N_4909,N_4214);
or UO_218 (O_218,N_4294,N_3508);
xor UO_219 (O_219,N_3698,N_4282);
or UO_220 (O_220,N_4185,N_3495);
nor UO_221 (O_221,N_4867,N_3918);
or UO_222 (O_222,N_2653,N_3283);
or UO_223 (O_223,N_2619,N_2665);
nor UO_224 (O_224,N_3319,N_3120);
nand UO_225 (O_225,N_2567,N_4263);
and UO_226 (O_226,N_3523,N_4705);
or UO_227 (O_227,N_4866,N_3128);
or UO_228 (O_228,N_3062,N_3348);
nor UO_229 (O_229,N_2845,N_3268);
or UO_230 (O_230,N_4031,N_4400);
nand UO_231 (O_231,N_2527,N_4514);
or UO_232 (O_232,N_3559,N_3089);
nor UO_233 (O_233,N_3496,N_4291);
or UO_234 (O_234,N_2779,N_4608);
xnor UO_235 (O_235,N_2973,N_2711);
and UO_236 (O_236,N_4211,N_3749);
xor UO_237 (O_237,N_2525,N_3208);
nand UO_238 (O_238,N_2804,N_4319);
xnor UO_239 (O_239,N_3921,N_3278);
nand UO_240 (O_240,N_2863,N_2701);
xnor UO_241 (O_241,N_3654,N_3236);
or UO_242 (O_242,N_4395,N_4941);
or UO_243 (O_243,N_3967,N_3430);
nor UO_244 (O_244,N_2939,N_3287);
xnor UO_245 (O_245,N_2915,N_4076);
nand UO_246 (O_246,N_4239,N_4960);
nor UO_247 (O_247,N_4609,N_3030);
nand UO_248 (O_248,N_2851,N_2890);
and UO_249 (O_249,N_4051,N_4948);
nand UO_250 (O_250,N_2635,N_2598);
and UO_251 (O_251,N_4531,N_3788);
or UO_252 (O_252,N_4009,N_3521);
nand UO_253 (O_253,N_2566,N_3962);
and UO_254 (O_254,N_2951,N_4376);
xnor UO_255 (O_255,N_3988,N_3863);
xor UO_256 (O_256,N_4835,N_2502);
xor UO_257 (O_257,N_2625,N_3377);
or UO_258 (O_258,N_3580,N_4702);
nor UO_259 (O_259,N_4457,N_3438);
and UO_260 (O_260,N_3157,N_3824);
nor UO_261 (O_261,N_3731,N_2560);
nand UO_262 (O_262,N_4719,N_4593);
nor UO_263 (O_263,N_4806,N_4013);
or UO_264 (O_264,N_4999,N_4033);
xor UO_265 (O_265,N_3767,N_4517);
nand UO_266 (O_266,N_4463,N_4863);
or UO_267 (O_267,N_3597,N_2703);
nand UO_268 (O_268,N_3205,N_4509);
and UO_269 (O_269,N_3085,N_3318);
xor UO_270 (O_270,N_3012,N_2838);
nand UO_271 (O_271,N_4541,N_2685);
and UO_272 (O_272,N_3601,N_2966);
and UO_273 (O_273,N_2607,N_3691);
and UO_274 (O_274,N_3193,N_3210);
or UO_275 (O_275,N_2666,N_4277);
nor UO_276 (O_276,N_4985,N_4015);
and UO_277 (O_277,N_4833,N_4872);
and UO_278 (O_278,N_3587,N_4590);
nor UO_279 (O_279,N_4183,N_3735);
or UO_280 (O_280,N_2729,N_4005);
xor UO_281 (O_281,N_4904,N_4285);
or UO_282 (O_282,N_3552,N_2885);
nand UO_283 (O_283,N_4809,N_2720);
nor UO_284 (O_284,N_3820,N_3105);
and UO_285 (O_285,N_3007,N_4599);
and UO_286 (O_286,N_4972,N_3579);
nand UO_287 (O_287,N_4002,N_2790);
and UO_288 (O_288,N_3417,N_4496);
xor UO_289 (O_289,N_3592,N_4102);
nand UO_290 (O_290,N_3102,N_4254);
or UO_291 (O_291,N_4628,N_3170);
nand UO_292 (O_292,N_4290,N_3369);
xor UO_293 (O_293,N_2673,N_2809);
xor UO_294 (O_294,N_2917,N_4518);
nor UO_295 (O_295,N_3112,N_4756);
or UO_296 (O_296,N_3480,N_3149);
and UO_297 (O_297,N_4113,N_3238);
xor UO_298 (O_298,N_2883,N_4341);
xor UO_299 (O_299,N_4484,N_3983);
or UO_300 (O_300,N_3368,N_3429);
nand UO_301 (O_301,N_4747,N_3960);
or UO_302 (O_302,N_3971,N_3673);
or UO_303 (O_303,N_4893,N_2596);
xor UO_304 (O_304,N_3568,N_2820);
nand UO_305 (O_305,N_2808,N_3384);
xnor UO_306 (O_306,N_3119,N_3079);
and UO_307 (O_307,N_4548,N_3705);
xnor UO_308 (O_308,N_4072,N_4237);
nor UO_309 (O_309,N_2603,N_2766);
nor UO_310 (O_310,N_4515,N_4318);
nand UO_311 (O_311,N_2907,N_4266);
or UO_312 (O_312,N_4119,N_4648);
nand UO_313 (O_313,N_2659,N_2858);
and UO_314 (O_314,N_4536,N_3925);
xnor UO_315 (O_315,N_3234,N_4487);
xor UO_316 (O_316,N_3442,N_3628);
or UO_317 (O_317,N_3742,N_4317);
nor UO_318 (O_318,N_3040,N_4138);
xnor UO_319 (O_319,N_2965,N_4649);
or UO_320 (O_320,N_4630,N_3343);
xor UO_321 (O_321,N_3730,N_4225);
nand UO_322 (O_322,N_2548,N_4956);
and UO_323 (O_323,N_4046,N_4427);
nand UO_324 (O_324,N_2844,N_2668);
xnor UO_325 (O_325,N_4874,N_2806);
xnor UO_326 (O_326,N_4818,N_3426);
nor UO_327 (O_327,N_3322,N_3896);
nand UO_328 (O_328,N_4787,N_4750);
or UO_329 (O_329,N_4108,N_3249);
and UO_330 (O_330,N_3302,N_4717);
and UO_331 (O_331,N_4614,N_3515);
and UO_332 (O_332,N_4572,N_3039);
and UO_333 (O_333,N_3812,N_2985);
and UO_334 (O_334,N_2987,N_3942);
nor UO_335 (O_335,N_4045,N_3292);
or UO_336 (O_336,N_4354,N_3003);
nand UO_337 (O_337,N_3876,N_4169);
nand UO_338 (O_338,N_4486,N_4538);
xor UO_339 (O_339,N_3094,N_2756);
or UO_340 (O_340,N_3542,N_4502);
and UO_341 (O_341,N_4150,N_3483);
xnor UO_342 (O_342,N_4439,N_4003);
nor UO_343 (O_343,N_3091,N_2935);
xor UO_344 (O_344,N_3201,N_4384);
xor UO_345 (O_345,N_2709,N_4301);
nand UO_346 (O_346,N_4575,N_3166);
nor UO_347 (O_347,N_3614,N_3852);
nand UO_348 (O_348,N_4839,N_3232);
xnor UO_349 (O_349,N_3274,N_4205);
and UO_350 (O_350,N_4695,N_4954);
xnor UO_351 (O_351,N_4978,N_3179);
nor UO_352 (O_352,N_4164,N_4241);
nand UO_353 (O_353,N_3364,N_2955);
or UO_354 (O_354,N_2855,N_4044);
or UO_355 (O_355,N_3522,N_2535);
and UO_356 (O_356,N_3553,N_3115);
nor UO_357 (O_357,N_2686,N_4206);
xor UO_358 (O_358,N_4936,N_3255);
nand UO_359 (O_359,N_3271,N_3701);
nor UO_360 (O_360,N_3206,N_2857);
nand UO_361 (O_361,N_4674,N_2676);
nor UO_362 (O_362,N_4428,N_3588);
xnor UO_363 (O_363,N_3664,N_3761);
nor UO_364 (O_364,N_4473,N_4100);
nor UO_365 (O_365,N_2912,N_4735);
nor UO_366 (O_366,N_3460,N_3315);
nand UO_367 (O_367,N_3476,N_2768);
or UO_368 (O_368,N_4445,N_3215);
and UO_369 (O_369,N_2968,N_4763);
nand UO_370 (O_370,N_3471,N_3633);
and UO_371 (O_371,N_3627,N_4191);
nand UO_372 (O_372,N_4601,N_3376);
or UO_373 (O_373,N_3263,N_4703);
nand UO_374 (O_374,N_3478,N_3656);
nor UO_375 (O_375,N_3456,N_4010);
or UO_376 (O_376,N_3358,N_3920);
xnor UO_377 (O_377,N_4817,N_4841);
nand UO_378 (O_378,N_3159,N_3233);
or UO_379 (O_379,N_2946,N_2684);
nand UO_380 (O_380,N_4857,N_2575);
nor UO_381 (O_381,N_4683,N_3847);
and UO_382 (O_382,N_4720,N_3957);
and UO_383 (O_383,N_2810,N_3578);
or UO_384 (O_384,N_3196,N_3662);
xor UO_385 (O_385,N_3821,N_2829);
and UO_386 (O_386,N_3408,N_3823);
xnor UO_387 (O_387,N_4323,N_3565);
xor UO_388 (O_388,N_3051,N_3650);
and UO_389 (O_389,N_3349,N_2814);
and UO_390 (O_390,N_3002,N_2758);
xnor UO_391 (O_391,N_3878,N_3563);
nor UO_392 (O_392,N_2613,N_4151);
nor UO_393 (O_393,N_3615,N_3605);
nor UO_394 (O_394,N_3912,N_3388);
and UO_395 (O_395,N_3810,N_3016);
xnor UO_396 (O_396,N_3231,N_3131);
and UO_397 (O_397,N_2934,N_3681);
nor UO_398 (O_398,N_2916,N_3688);
xor UO_399 (O_399,N_3757,N_2611);
nor UO_400 (O_400,N_3607,N_3979);
nand UO_401 (O_401,N_3487,N_3472);
nand UO_402 (O_402,N_4134,N_2588);
xnor UO_403 (O_403,N_3611,N_4383);
nand UO_404 (O_404,N_3696,N_2538);
nand UO_405 (O_405,N_3505,N_2881);
or UO_406 (O_406,N_4523,N_4188);
and UO_407 (O_407,N_2825,N_3290);
nand UO_408 (O_408,N_4672,N_3172);
xor UO_409 (O_409,N_3489,N_2561);
nor UO_410 (O_410,N_3798,N_4823);
or UO_411 (O_411,N_4934,N_3813);
nor UO_412 (O_412,N_3180,N_2892);
nor UO_413 (O_413,N_3036,N_3053);
xnor UO_414 (O_414,N_3332,N_4603);
xor UO_415 (O_415,N_4361,N_3926);
nand UO_416 (O_416,N_3214,N_4453);
or UO_417 (O_417,N_3944,N_3031);
or UO_418 (O_418,N_3976,N_4513);
and UO_419 (O_419,N_3968,N_3078);
nand UO_420 (O_420,N_3275,N_3316);
nor UO_421 (O_421,N_3871,N_2621);
and UO_422 (O_422,N_4414,N_3644);
nor UO_423 (O_423,N_3783,N_4798);
and UO_424 (O_424,N_3410,N_2642);
nand UO_425 (O_425,N_2736,N_4540);
nor UO_426 (O_426,N_3954,N_4767);
xnor UO_427 (O_427,N_3458,N_4368);
and UO_428 (O_428,N_2925,N_3459);
nor UO_429 (O_429,N_3467,N_3015);
and UO_430 (O_430,N_4371,N_3427);
or UO_431 (O_431,N_3955,N_4792);
or UO_432 (O_432,N_4052,N_3219);
and UO_433 (O_433,N_3103,N_2752);
or UO_434 (O_434,N_2593,N_4265);
or UO_435 (O_435,N_3532,N_3123);
nand UO_436 (O_436,N_2674,N_3399);
or UO_437 (O_437,N_4271,N_3687);
or UO_438 (O_438,N_4402,N_4884);
nor UO_439 (O_439,N_4613,N_2581);
xor UO_440 (O_440,N_4465,N_3518);
nor UO_441 (O_441,N_4000,N_2961);
and UO_442 (O_442,N_3291,N_2944);
or UO_443 (O_443,N_4759,N_4375);
nand UO_444 (O_444,N_2584,N_3941);
xor UO_445 (O_445,N_4563,N_4325);
nand UO_446 (O_446,N_4622,N_2919);
xnor UO_447 (O_447,N_4997,N_4246);
xnor UO_448 (O_448,N_3545,N_4659);
or UO_449 (O_449,N_3488,N_3405);
nand UO_450 (O_450,N_4392,N_2891);
and UO_451 (O_451,N_2866,N_3796);
nor UO_452 (O_452,N_3057,N_3299);
nand UO_453 (O_453,N_2872,N_2932);
or UO_454 (O_454,N_4736,N_4680);
nor UO_455 (O_455,N_3421,N_2706);
nand UO_456 (O_456,N_3295,N_3230);
or UO_457 (O_457,N_4407,N_4049);
xor UO_458 (O_458,N_4449,N_4131);
and UO_459 (O_459,N_3167,N_2799);
or UO_460 (O_460,N_3726,N_4951);
nand UO_461 (O_461,N_3044,N_4377);
nor UO_462 (O_462,N_4666,N_3484);
xnor UO_463 (O_463,N_3000,N_2997);
nor UO_464 (O_464,N_3817,N_4468);
xor UO_465 (O_465,N_3888,N_2647);
xnor UO_466 (O_466,N_4004,N_3136);
nand UO_467 (O_467,N_2571,N_3683);
or UO_468 (O_468,N_3935,N_4528);
and UO_469 (O_469,N_3689,N_3787);
xnor UO_470 (O_470,N_3448,N_4446);
nand UO_471 (O_471,N_4248,N_4554);
nand UO_472 (O_472,N_4670,N_2776);
or UO_473 (O_473,N_4207,N_4923);
xnor UO_474 (O_474,N_4594,N_3905);
nor UO_475 (O_475,N_4611,N_3190);
or UO_476 (O_476,N_3537,N_4236);
and UO_477 (O_477,N_4298,N_4353);
or UO_478 (O_478,N_2573,N_2819);
nand UO_479 (O_479,N_4132,N_2623);
xnor UO_480 (O_480,N_3632,N_3118);
xnor UO_481 (O_481,N_4921,N_2698);
and UO_482 (O_482,N_4851,N_3738);
or UO_483 (O_483,N_3719,N_2854);
and UO_484 (O_484,N_4482,N_4769);
nand UO_485 (O_485,N_2860,N_4162);
nor UO_486 (O_486,N_2743,N_3845);
or UO_487 (O_487,N_4344,N_4438);
and UO_488 (O_488,N_4671,N_3087);
xnor UO_489 (O_489,N_4130,N_3009);
nand UO_490 (O_490,N_2746,N_4098);
nor UO_491 (O_491,N_2521,N_4701);
nor UO_492 (O_492,N_4991,N_3412);
xor UO_493 (O_493,N_2831,N_4927);
and UO_494 (O_494,N_4415,N_4713);
nand UO_495 (O_495,N_4731,N_4442);
nor UO_496 (O_496,N_3207,N_4698);
xnor UO_497 (O_497,N_3856,N_3956);
xnor UO_498 (O_498,N_4017,N_3221);
nor UO_499 (O_499,N_3020,N_2731);
nand UO_500 (O_500,N_3612,N_3591);
or UO_501 (O_501,N_2850,N_2576);
nand UO_502 (O_502,N_3684,N_2690);
and UO_503 (O_503,N_2794,N_4580);
and UO_504 (O_504,N_3864,N_3853);
xnor UO_505 (O_505,N_3741,N_3253);
or UO_506 (O_506,N_2504,N_2615);
and UO_507 (O_507,N_2867,N_3037);
xnor UO_508 (O_508,N_3258,N_2648);
nand UO_509 (O_509,N_4615,N_3280);
nand UO_510 (O_510,N_3224,N_3751);
or UO_511 (O_511,N_3634,N_3286);
or UO_512 (O_512,N_3043,N_4065);
nor UO_513 (O_513,N_2687,N_3997);
or UO_514 (O_514,N_4974,N_2519);
and UO_515 (O_515,N_4469,N_3838);
xnor UO_516 (O_516,N_3703,N_3466);
xnor UO_517 (O_517,N_4152,N_3248);
or UO_518 (O_518,N_4558,N_3511);
xnor UO_519 (O_519,N_4316,N_3314);
xor UO_520 (O_520,N_3659,N_3855);
nor UO_521 (O_521,N_3194,N_3025);
xor UO_522 (O_522,N_3109,N_4172);
xnor UO_523 (O_523,N_4332,N_3400);
or UO_524 (O_524,N_4802,N_4612);
nand UO_525 (O_525,N_3780,N_3422);
nor UO_526 (O_526,N_4914,N_2639);
or UO_527 (O_527,N_4710,N_2846);
and UO_528 (O_528,N_4552,N_3344);
xnor UO_529 (O_529,N_3305,N_3778);
nor UO_530 (O_530,N_4153,N_4129);
xnor UO_531 (O_531,N_4190,N_4255);
or UO_532 (O_532,N_4556,N_3904);
or UO_533 (O_533,N_2859,N_3494);
nor UO_534 (O_534,N_4895,N_4040);
or UO_535 (O_535,N_2732,N_3567);
and UO_536 (O_536,N_4114,N_4202);
nor UO_537 (O_537,N_3547,N_4270);
and UO_538 (O_538,N_2641,N_4423);
nand UO_539 (O_539,N_2787,N_4684);
xnor UO_540 (O_540,N_2914,N_3999);
nor UO_541 (O_541,N_3092,N_2726);
and UO_542 (O_542,N_3924,N_3561);
xnor UO_543 (O_543,N_2602,N_3074);
or UO_544 (O_544,N_3657,N_4454);
nand UO_545 (O_545,N_3076,N_4273);
xnor UO_546 (O_546,N_4352,N_3829);
nand UO_547 (O_547,N_3393,N_3265);
and UO_548 (O_548,N_3055,N_2704);
nand UO_549 (O_549,N_3310,N_3168);
and UO_550 (O_550,N_2876,N_3005);
and UO_551 (O_551,N_3617,N_3504);
and UO_552 (O_552,N_3445,N_4821);
and UO_553 (O_553,N_4641,N_4559);
nand UO_554 (O_554,N_2783,N_3715);
or UO_555 (O_555,N_3342,N_4101);
nor UO_556 (O_556,N_3470,N_4521);
nand UO_557 (O_557,N_2631,N_3946);
and UO_558 (O_558,N_3435,N_4778);
nor UO_559 (O_559,N_3449,N_3585);
nor UO_560 (O_560,N_4115,N_2828);
and UO_561 (O_561,N_3223,N_3158);
and UO_562 (O_562,N_2906,N_4216);
nor UO_563 (O_563,N_2543,N_3911);
nand UO_564 (O_564,N_3146,N_2983);
nor UO_565 (O_565,N_3551,N_3083);
nand UO_566 (O_566,N_2640,N_3973);
or UO_567 (O_567,N_4364,N_4267);
nor UO_568 (O_568,N_3104,N_2563);
xnor UO_569 (O_569,N_3259,N_4426);
and UO_570 (O_570,N_3922,N_4326);
or UO_571 (O_571,N_3746,N_3396);
or UO_572 (O_572,N_3502,N_2927);
nand UO_573 (O_573,N_2970,N_3213);
xnor UO_574 (O_574,N_4173,N_3026);
nor UO_575 (O_575,N_2592,N_3958);
nor UO_576 (O_576,N_2644,N_4362);
nand UO_577 (O_577,N_3404,N_4946);
xor UO_578 (O_578,N_4878,N_4083);
and UO_579 (O_579,N_3296,N_2807);
or UO_580 (O_580,N_3341,N_4466);
or UO_581 (O_581,N_2800,N_4222);
nand UO_582 (O_582,N_3694,N_3616);
and UO_583 (O_583,N_3070,N_3122);
xor UO_584 (O_584,N_2797,N_2847);
xnor UO_585 (O_585,N_4918,N_4633);
nor UO_586 (O_586,N_3700,N_2979);
xor UO_587 (O_587,N_4103,N_2978);
or UO_588 (O_588,N_3184,N_3463);
nand UO_589 (O_589,N_4676,N_4727);
nor UO_590 (O_590,N_2661,N_3831);
and UO_591 (O_591,N_4460,N_4425);
or UO_592 (O_592,N_2716,N_4435);
or UO_593 (O_593,N_3211,N_4675);
or UO_594 (O_594,N_4444,N_2539);
and UO_595 (O_595,N_4722,N_4932);
nor UO_596 (O_596,N_4242,N_3714);
or UO_597 (O_597,N_2759,N_4987);
nor UO_598 (O_598,N_4210,N_2529);
and UO_599 (O_599,N_4215,N_3862);
xnor UO_600 (O_600,N_2909,N_3756);
xnor UO_601 (O_601,N_4314,N_3140);
nand UO_602 (O_602,N_3758,N_4022);
nand UO_603 (O_603,N_2938,N_3875);
or UO_604 (O_604,N_3775,N_2908);
and UO_605 (O_605,N_4322,N_3336);
nand UO_606 (O_606,N_4109,N_2536);
and UO_607 (O_607,N_4447,N_4408);
or UO_608 (O_608,N_4112,N_3902);
nand UO_609 (O_609,N_4067,N_2501);
nand UO_610 (O_610,N_3416,N_4856);
or UO_611 (O_611,N_4882,N_4107);
xor UO_612 (O_612,N_4366,N_4865);
or UO_613 (O_613,N_3892,N_4213);
nand UO_614 (O_614,N_4313,N_4339);
nor UO_615 (O_615,N_3250,N_4880);
xnor UO_616 (O_616,N_4958,N_2826);
and UO_617 (O_617,N_4204,N_2526);
xor UO_618 (O_618,N_4081,N_4082);
or UO_619 (O_619,N_3363,N_2902);
nand UO_620 (O_620,N_3398,N_4913);
or UO_621 (O_621,N_4700,N_3059);
nand UO_622 (O_622,N_3770,N_3338);
nand UO_623 (O_623,N_3527,N_4403);
and UO_624 (O_624,N_3842,N_3927);
xor UO_625 (O_625,N_3165,N_4381);
and UO_626 (O_626,N_4124,N_2937);
nor UO_627 (O_627,N_3468,N_3365);
and UO_628 (O_628,N_3613,N_4854);
and UO_629 (O_629,N_4006,N_3707);
and UO_630 (O_630,N_2764,N_2552);
and UO_631 (O_631,N_2723,N_3064);
nand UO_632 (O_632,N_4197,N_3251);
or UO_633 (O_633,N_3147,N_4690);
and UO_634 (O_634,N_3986,N_4729);
and UO_635 (O_635,N_4643,N_2675);
or UO_636 (O_636,N_4480,N_3649);
and UO_637 (O_637,N_4304,N_3135);
and UO_638 (O_638,N_3362,N_3755);
or UO_639 (O_639,N_4176,N_3436);
nor UO_640 (O_640,N_4462,N_4334);
and UO_641 (O_641,N_3151,N_4347);
and UO_642 (O_642,N_4147,N_4497);
xnor UO_643 (O_643,N_4669,N_3303);
nor UO_644 (O_644,N_4950,N_3695);
nor UO_645 (O_645,N_4892,N_3835);
and UO_646 (O_646,N_3013,N_3929);
or UO_647 (O_647,N_3284,N_4899);
or UO_648 (O_648,N_2980,N_3389);
nor UO_649 (O_649,N_2956,N_4136);
nor UO_650 (O_650,N_4662,N_4283);
and UO_651 (O_651,N_4898,N_4099);
xnor UO_652 (O_652,N_3987,N_4019);
and UO_653 (O_653,N_3709,N_4520);
and UO_654 (O_654,N_2645,N_3352);
or UO_655 (O_655,N_4068,N_4001);
or UO_656 (O_656,N_3289,N_3895);
nand UO_657 (O_657,N_2811,N_4122);
and UO_658 (O_658,N_4522,N_3762);
or UO_659 (O_659,N_2848,N_4440);
nor UO_660 (O_660,N_4587,N_2714);
and UO_661 (O_661,N_4363,N_2638);
and UO_662 (O_662,N_4511,N_4170);
xnor UO_663 (O_663,N_3228,N_3345);
xor UO_664 (O_664,N_3554,N_4908);
and UO_665 (O_665,N_4738,N_4315);
or UO_666 (O_666,N_4064,N_2531);
nand UO_667 (O_667,N_4655,N_2868);
or UO_668 (O_668,N_3622,N_3464);
nor UO_669 (O_669,N_3257,N_4885);
xor UO_670 (O_670,N_2789,N_2780);
nand UO_671 (O_671,N_3916,N_3913);
xor UO_672 (O_672,N_3203,N_3899);
nor UO_673 (O_673,N_2678,N_4739);
and UO_674 (O_674,N_2663,N_4229);
nor UO_675 (O_675,N_3734,N_2751);
nor UO_676 (O_676,N_4765,N_4578);
xnor UO_677 (O_677,N_2614,N_3558);
nor UO_678 (O_678,N_2903,N_4422);
nor UO_679 (O_679,N_3272,N_4619);
and UO_680 (O_680,N_4808,N_4733);
xor UO_681 (O_681,N_4530,N_2900);
nor UO_682 (O_682,N_3843,N_2821);
nand UO_683 (O_683,N_2694,N_3868);
nor UO_684 (O_684,N_3328,N_4012);
nor UO_685 (O_685,N_3608,N_4171);
nor UO_686 (O_686,N_4491,N_3406);
nor UO_687 (O_687,N_2738,N_4557);
and UO_688 (O_688,N_4687,N_3583);
xor UO_689 (O_689,N_2879,N_2511);
or UO_690 (O_690,N_4259,N_3237);
nand UO_691 (O_691,N_3859,N_2651);
nor UO_692 (O_692,N_3555,N_4370);
xnor UO_693 (O_693,N_2654,N_2587);
or UO_694 (O_694,N_4783,N_3978);
nor UO_695 (O_695,N_4577,N_2834);
nand UO_696 (O_696,N_4582,N_3534);
or UO_697 (O_697,N_3453,N_4079);
nand UO_698 (O_698,N_3699,N_4485);
and UO_699 (O_699,N_3402,N_4018);
nand UO_700 (O_700,N_2583,N_3792);
nor UO_701 (O_701,N_4644,N_4493);
or UO_702 (O_702,N_2601,N_3998);
nand UO_703 (O_703,N_3697,N_2739);
and UO_704 (O_704,N_4797,N_2773);
nor UO_705 (O_705,N_3690,N_4617);
or UO_706 (O_706,N_3623,N_4433);
nand UO_707 (O_707,N_2984,N_2597);
or UO_708 (O_708,N_4181,N_4417);
nand UO_709 (O_709,N_3854,N_3618);
and UO_710 (O_710,N_4853,N_3247);
nand UO_711 (O_711,N_3857,N_4223);
xor UO_712 (O_712,N_3097,N_4106);
or UO_713 (O_713,N_3880,N_3273);
nand UO_714 (O_714,N_3743,N_3028);
or UO_715 (O_715,N_4218,N_4476);
or UO_716 (O_716,N_3586,N_2503);
and UO_717 (O_717,N_3033,N_4311);
and UO_718 (O_718,N_4715,N_3304);
xnor UO_719 (O_719,N_3082,N_4831);
nand UO_720 (O_720,N_2801,N_4163);
xnor UO_721 (O_721,N_3850,N_2803);
nor UO_722 (O_722,N_3543,N_3932);
or UO_723 (O_723,N_4043,N_2977);
or UO_724 (O_724,N_4420,N_4744);
nor UO_725 (O_725,N_4820,N_3367);
xnor UO_726 (O_726,N_4320,N_2637);
and UO_727 (O_727,N_4146,N_3071);
or UO_728 (O_728,N_4877,N_3919);
nand UO_729 (O_729,N_4155,N_3096);
nand UO_730 (O_730,N_4688,N_4624);
and UO_731 (O_731,N_2600,N_4472);
xor UO_732 (O_732,N_3038,N_2516);
and UO_733 (O_733,N_3540,N_4929);
nor UO_734 (O_734,N_4961,N_4957);
nor UO_735 (O_735,N_2895,N_3312);
nand UO_736 (O_736,N_2962,N_4272);
xor UO_737 (O_737,N_4803,N_4973);
or UO_738 (O_738,N_4764,N_3704);
or UO_739 (O_739,N_4786,N_2818);
and UO_740 (O_740,N_4864,N_3646);
or UO_741 (O_741,N_2585,N_4875);
and UO_742 (O_742,N_3717,N_4890);
nor UO_743 (O_743,N_3947,N_3199);
xor UO_744 (O_744,N_3117,N_3178);
nor UO_745 (O_745,N_4840,N_2772);
nand UO_746 (O_746,N_2662,N_4938);
or UO_747 (O_747,N_3693,N_3163);
and UO_748 (O_748,N_3395,N_4281);
or UO_749 (O_749,N_3355,N_4088);
xnor UO_750 (O_750,N_2782,N_3011);
and UO_751 (O_751,N_3797,N_3425);
or UO_752 (O_752,N_3951,N_3781);
nand UO_753 (O_753,N_3745,N_4993);
nand UO_754 (O_754,N_3052,N_2887);
and UO_755 (O_755,N_2926,N_4310);
nor UO_756 (O_756,N_3125,N_3492);
or UO_757 (O_757,N_2953,N_3536);
xnor UO_758 (O_758,N_4751,N_4016);
xor UO_759 (O_759,N_2959,N_3462);
or UO_760 (O_760,N_3413,N_3984);
and UO_761 (O_761,N_2707,N_4879);
or UO_762 (O_762,N_4746,N_3447);
nand UO_763 (O_763,N_4406,N_4481);
or UO_764 (O_764,N_4437,N_4860);
nor UO_765 (O_765,N_4777,N_4714);
or UO_766 (O_766,N_3723,N_2920);
nor UO_767 (O_767,N_2577,N_3839);
xnor UO_768 (O_768,N_3148,N_4159);
xnor UO_769 (O_769,N_4396,N_4694);
or UO_770 (O_770,N_4077,N_4156);
xor UO_771 (O_771,N_3637,N_2693);
and UO_772 (O_772,N_2533,N_4754);
nor UO_773 (O_773,N_4668,N_4804);
or UO_774 (O_774,N_3865,N_3804);
nor UO_775 (O_775,N_3331,N_4324);
and UO_776 (O_776,N_2741,N_4842);
or UO_777 (O_777,N_2929,N_2999);
and UO_778 (O_778,N_3513,N_3415);
nor UO_779 (O_779,N_2791,N_2579);
and UO_780 (O_780,N_4926,N_2958);
xor UO_781 (O_781,N_2617,N_2658);
or UO_782 (O_782,N_4771,N_3676);
nor UO_783 (O_783,N_2733,N_4126);
xor UO_784 (O_784,N_3860,N_4387);
or UO_785 (O_785,N_4194,N_4945);
xnor UO_786 (O_786,N_4253,N_2940);
xor UO_787 (O_787,N_4086,N_3154);
or UO_788 (O_788,N_3246,N_4686);
or UO_789 (O_789,N_4258,N_3934);
xnor UO_790 (O_790,N_2864,N_3894);
xor UO_791 (O_791,N_3114,N_3653);
xnor UO_792 (O_792,N_2877,N_3933);
and UO_793 (O_793,N_4508,N_4091);
or UO_794 (O_794,N_2532,N_3571);
and UO_795 (O_795,N_4066,N_4050);
xor UO_796 (O_796,N_2778,N_2520);
and UO_797 (O_797,N_4965,N_4616);
xor UO_798 (O_798,N_4125,N_3254);
xnor UO_799 (O_799,N_4494,N_3562);
and UO_800 (O_800,N_2737,N_3129);
and UO_801 (O_801,N_3346,N_3225);
xor UO_802 (O_802,N_3815,N_4104);
or UO_803 (O_803,N_4766,N_3216);
and UO_804 (O_804,N_4374,N_3240);
nand UO_805 (O_805,N_2522,N_4992);
xor UO_806 (O_806,N_3535,N_3631);
nand UO_807 (O_807,N_4145,N_4014);
or UO_808 (O_808,N_4718,N_3516);
xnor UO_809 (O_809,N_4404,N_4506);
nor UO_810 (O_810,N_2995,N_2649);
and UO_811 (O_811,N_3401,N_4149);
nor UO_812 (O_812,N_3772,N_4429);
nor UO_813 (O_813,N_2960,N_4090);
and UO_814 (O_814,N_4269,N_4221);
nand UO_815 (O_815,N_2505,N_3642);
nor UO_816 (O_816,N_4537,N_4525);
or UO_817 (O_817,N_4063,N_4602);
xor UO_818 (O_818,N_4920,N_3242);
nor UO_819 (O_819,N_3702,N_4790);
nor UO_820 (O_820,N_3473,N_2798);
nand UO_821 (O_821,N_2870,N_4252);
and UO_822 (O_822,N_4567,N_2918);
nand UO_823 (O_823,N_2549,N_3674);
and UO_824 (O_824,N_4041,N_4737);
xnor UO_825 (O_825,N_3455,N_3528);
and UO_826 (O_826,N_4288,N_2769);
or UO_827 (O_827,N_3220,N_4293);
or UO_828 (O_828,N_3187,N_2632);
or UO_829 (O_829,N_4801,N_3782);
or UO_830 (O_830,N_3624,N_4505);
and UO_831 (O_831,N_2969,N_3269);
or UO_832 (O_832,N_3189,N_4489);
nor UO_833 (O_833,N_3218,N_4208);
nor UO_834 (O_834,N_4553,N_2650);
nand UO_835 (O_835,N_2943,N_2993);
nor UO_836 (O_836,N_3499,N_2824);
or UO_837 (O_837,N_3510,N_4458);
xor UO_838 (O_838,N_4276,N_3785);
or UO_839 (O_839,N_3261,N_3351);
and UO_840 (O_840,N_4829,N_4167);
nor UO_841 (O_841,N_3397,N_4367);
nand UO_842 (O_842,N_3557,N_3046);
nor UO_843 (O_843,N_2898,N_4562);
nor UO_844 (O_844,N_3403,N_3759);
and UO_845 (O_845,N_4776,N_2695);
or UO_846 (O_846,N_3548,N_4566);
nor UO_847 (O_847,N_4073,N_3908);
and UO_848 (O_848,N_4944,N_2730);
nor UO_849 (O_849,N_4504,N_2734);
or UO_850 (O_850,N_3018,N_3635);
or UO_851 (O_851,N_4074,N_2582);
nor UO_852 (O_852,N_4461,N_4336);
nor UO_853 (O_853,N_3256,N_3501);
nand UO_854 (O_854,N_4819,N_2609);
nor UO_855 (O_855,N_3134,N_4337);
nand UO_856 (O_856,N_3584,N_4573);
nand UO_857 (O_857,N_3450,N_4903);
nand UO_858 (O_858,N_4346,N_3321);
nand UO_859 (O_859,N_2971,N_2570);
and UO_860 (O_860,N_4605,N_4028);
nor UO_861 (O_861,N_4924,N_4182);
and UO_862 (O_862,N_2652,N_3671);
or UO_863 (O_863,N_4305,N_3301);
xor UO_864 (O_864,N_4779,N_4969);
or UO_865 (O_865,N_4861,N_3981);
nand UO_866 (O_866,N_3001,N_4240);
xor UO_867 (O_867,N_3803,N_3771);
or UO_868 (O_868,N_3811,N_3385);
xor UO_869 (O_869,N_3830,N_4896);
and UO_870 (O_870,N_3915,N_4399);
and UO_871 (O_871,N_4342,N_3963);
xor UO_872 (O_872,N_3764,N_3840);
nand UO_873 (O_873,N_2745,N_3029);
or UO_874 (O_874,N_3975,N_3887);
and UO_875 (O_875,N_4093,N_4579);
nand UO_876 (O_876,N_4195,N_3581);
xor UO_877 (O_877,N_4455,N_2785);
nand UO_878 (O_878,N_3678,N_4192);
and UO_879 (O_879,N_4386,N_3885);
xnor UO_880 (O_880,N_4828,N_4230);
nand UO_881 (O_881,N_3334,N_3900);
or UO_882 (O_882,N_4812,N_3068);
or UO_883 (O_883,N_4510,N_3982);
or UO_884 (O_884,N_3021,N_4474);
or UO_885 (O_885,N_2880,N_4245);
nand UO_886 (O_886,N_4785,N_3910);
nor UO_887 (O_887,N_4791,N_3381);
nand UO_888 (O_888,N_4544,N_4539);
xor UO_889 (O_889,N_3711,N_2594);
nand UO_890 (O_890,N_4350,N_4475);
nor UO_891 (O_891,N_2710,N_4966);
or UO_892 (O_892,N_4916,N_4788);
nor UO_893 (O_893,N_3996,N_4499);
nand UO_894 (O_894,N_2569,N_4256);
xor UO_895 (O_895,N_4186,N_4095);
nand UO_896 (O_896,N_2721,N_2873);
or UO_897 (O_897,N_2604,N_4663);
xor UO_898 (O_898,N_3596,N_3431);
nor UO_899 (O_899,N_4862,N_3058);
and UO_900 (O_900,N_3891,N_3640);
nand UO_901 (O_901,N_4441,N_4900);
nor UO_902 (O_902,N_4772,N_2765);
nand UO_903 (O_903,N_3994,N_2793);
nor UO_904 (O_904,N_4312,N_3424);
and UO_905 (O_905,N_3110,N_3752);
xor UO_906 (O_906,N_2719,N_4607);
nor UO_907 (O_907,N_4287,N_3546);
nor UO_908 (O_908,N_3750,N_3529);
or UO_909 (O_909,N_4062,N_4574);
and UO_910 (O_910,N_3107,N_3795);
nor UO_911 (O_911,N_2830,N_2669);
nand UO_912 (O_912,N_3183,N_3727);
nand UO_913 (O_913,N_3241,N_3390);
or UO_914 (O_914,N_4656,N_3497);
or UO_915 (O_915,N_2630,N_2750);
or UO_916 (O_916,N_3630,N_2839);
nand UO_917 (O_917,N_3658,N_3517);
xnor UO_918 (O_918,N_3881,N_3574);
xor UO_919 (O_919,N_4477,N_3909);
xnor UO_920 (O_920,N_2725,N_4470);
nand UO_921 (O_921,N_3520,N_4127);
nor UO_922 (O_922,N_4651,N_3747);
nor UO_923 (O_923,N_3872,N_4546);
nor UO_924 (O_924,N_2509,N_3686);
or UO_925 (O_925,N_3409,N_3173);
nor UO_926 (O_926,N_4512,N_4080);
and UO_927 (O_927,N_2507,N_3423);
xor UO_928 (O_928,N_3648,N_4623);
xnor UO_929 (O_929,N_3867,N_2817);
and UO_930 (O_930,N_2546,N_4911);
and UO_931 (O_931,N_4303,N_4340);
nand UO_932 (O_932,N_4982,N_3481);
or UO_933 (O_933,N_4233,N_4390);
and UO_934 (O_934,N_3264,N_3636);
nand UO_935 (O_935,N_4029,N_2816);
or UO_936 (O_936,N_4343,N_3375);
or UO_937 (O_937,N_2727,N_4589);
and UO_938 (O_938,N_4711,N_3736);
nand UO_939 (O_939,N_4532,N_4328);
and UO_940 (O_940,N_4168,N_4632);
and UO_941 (O_941,N_2749,N_3469);
and UO_942 (O_942,N_3576,N_4144);
nand UO_943 (O_943,N_4409,N_3826);
and UO_944 (O_944,N_3990,N_4059);
nand UO_945 (O_945,N_4189,N_4859);
or UO_946 (O_946,N_4849,N_4784);
xor UO_947 (O_947,N_3454,N_4834);
nand UO_948 (O_948,N_4922,N_2874);
nor UO_949 (O_949,N_3185,N_3765);
and UO_950 (O_950,N_3940,N_4876);
and UO_951 (O_951,N_4568,N_3643);
nand UO_952 (O_952,N_4551,N_4321);
xor UO_953 (O_953,N_3407,N_4741);
nand UO_954 (O_954,N_2633,N_3162);
and UO_955 (O_955,N_3943,N_4979);
nor UO_956 (O_956,N_4292,N_4576);
or UO_957 (O_957,N_3340,N_2865);
xnor UO_958 (O_958,N_4618,N_3677);
nor UO_959 (O_959,N_3017,N_3260);
nor UO_960 (O_960,N_3870,N_4858);
and UO_961 (O_961,N_3330,N_4762);
xnor UO_962 (O_962,N_3906,N_2786);
xnor UO_963 (O_963,N_3818,N_4280);
and UO_964 (O_964,N_2512,N_4681);
nand UO_965 (O_965,N_4959,N_4372);
and UO_966 (O_966,N_4500,N_4274);
xor UO_967 (O_967,N_3773,N_4410);
or UO_968 (O_968,N_4815,N_2626);
or UO_969 (O_969,N_3573,N_2897);
or UO_970 (O_970,N_2667,N_3202);
nor UO_971 (O_971,N_4749,N_4837);
xor UO_972 (O_972,N_3833,N_2967);
and UO_973 (O_973,N_3077,N_2792);
and UO_974 (O_974,N_3786,N_4638);
and UO_975 (O_975,N_3739,N_3884);
or UO_976 (O_976,N_2748,N_3594);
or UO_977 (O_977,N_4986,N_4855);
nand UO_978 (O_978,N_2875,N_4503);
and UO_979 (O_979,N_2893,N_3419);
nor UO_980 (O_980,N_3465,N_3512);
nand UO_981 (O_981,N_4110,N_4120);
nand UO_982 (O_982,N_2805,N_4309);
xnor UO_983 (O_983,N_2942,N_3800);
nor UO_984 (O_984,N_3619,N_3006);
and UO_985 (O_985,N_4962,N_3903);
and UO_986 (O_986,N_2523,N_4335);
nand UO_987 (O_987,N_4516,N_4665);
xor UO_988 (O_988,N_3808,N_3008);
nand UO_989 (O_989,N_3374,N_3239);
xor UO_990 (O_990,N_3712,N_2921);
nor UO_991 (O_991,N_3444,N_3347);
and UO_992 (O_992,N_4032,N_4349);
and UO_993 (O_993,N_2833,N_4526);
and UO_994 (O_994,N_4471,N_4555);
or UO_995 (O_995,N_4405,N_3564);
and UO_996 (O_996,N_4141,N_3621);
xor UO_997 (O_997,N_4871,N_3953);
nand UO_998 (O_998,N_3836,N_3959);
xor UO_999 (O_999,N_4707,N_3212);
endmodule