module basic_500_3000_500_50_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_100,In_335);
nand U1 (N_1,In_268,In_83);
or U2 (N_2,In_280,In_464);
nand U3 (N_3,In_266,In_6);
nor U4 (N_4,In_462,In_165);
or U5 (N_5,In_105,In_180);
nor U6 (N_6,In_97,In_161);
and U7 (N_7,In_194,In_233);
nand U8 (N_8,In_433,In_444);
and U9 (N_9,In_98,In_236);
nand U10 (N_10,In_206,In_293);
nand U11 (N_11,In_303,In_405);
or U12 (N_12,In_155,In_474);
nor U13 (N_13,In_57,In_213);
and U14 (N_14,In_416,In_488);
nand U15 (N_15,In_21,In_35);
nand U16 (N_16,In_350,In_435);
nand U17 (N_17,In_443,In_459);
or U18 (N_18,In_167,In_11);
and U19 (N_19,In_375,In_204);
or U20 (N_20,In_377,In_480);
nor U21 (N_21,In_492,In_17);
nor U22 (N_22,In_215,In_86);
nor U23 (N_23,In_491,In_470);
and U24 (N_24,In_340,In_185);
and U25 (N_25,In_168,In_113);
and U26 (N_26,In_490,In_445);
or U27 (N_27,In_329,In_338);
and U28 (N_28,In_391,In_395);
nand U29 (N_29,In_239,In_363);
nor U30 (N_30,In_423,In_65);
and U31 (N_31,In_414,In_454);
nand U32 (N_32,In_258,In_412);
nor U33 (N_33,In_326,In_298);
nor U34 (N_34,In_368,In_420);
nand U35 (N_35,In_43,In_149);
nand U36 (N_36,In_288,In_379);
and U37 (N_37,In_138,In_489);
or U38 (N_38,In_425,In_243);
nand U39 (N_39,In_223,In_94);
nor U40 (N_40,In_132,In_409);
xor U41 (N_41,In_345,In_225);
and U42 (N_42,In_121,In_66);
or U43 (N_43,In_34,In_378);
nand U44 (N_44,In_118,In_81);
or U45 (N_45,In_170,In_274);
or U46 (N_46,In_297,In_364);
or U47 (N_47,In_342,In_264);
and U48 (N_48,In_261,In_32);
nand U49 (N_49,In_183,In_212);
nor U50 (N_50,In_332,In_242);
nor U51 (N_51,In_51,In_31);
nor U52 (N_52,In_127,In_201);
or U53 (N_53,In_446,In_278);
or U54 (N_54,In_486,In_166);
and U55 (N_55,In_410,In_199);
nand U56 (N_56,In_214,In_245);
or U57 (N_57,In_90,In_269);
nor U58 (N_58,In_473,In_307);
nor U59 (N_59,In_203,In_354);
nand U60 (N_60,In_358,N_36);
xnor U61 (N_61,In_281,In_262);
and U62 (N_62,N_1,In_485);
and U63 (N_63,In_487,N_53);
nor U64 (N_64,In_41,In_361);
and U65 (N_65,In_402,In_82);
and U66 (N_66,In_343,N_58);
and U67 (N_67,In_426,In_150);
or U68 (N_68,In_62,In_455);
or U69 (N_69,N_6,In_253);
nor U70 (N_70,In_2,In_19);
nor U71 (N_71,In_46,In_394);
nor U72 (N_72,N_39,In_483);
and U73 (N_73,In_219,In_373);
nand U74 (N_74,N_30,In_76);
nand U75 (N_75,In_109,In_408);
nand U76 (N_76,In_353,In_226);
and U77 (N_77,In_388,In_498);
or U78 (N_78,In_305,In_99);
nand U79 (N_79,In_169,In_188);
nor U80 (N_80,In_187,In_23);
nor U81 (N_81,In_115,N_45);
nand U82 (N_82,In_383,In_334);
or U83 (N_83,In_58,In_229);
or U84 (N_84,In_456,In_88);
and U85 (N_85,In_424,In_221);
and U86 (N_86,N_51,In_176);
nor U87 (N_87,N_52,In_207);
and U88 (N_88,In_369,In_385);
nand U89 (N_89,In_277,N_40);
nand U90 (N_90,In_413,In_124);
nand U91 (N_91,In_439,In_60);
nor U92 (N_92,In_69,N_32);
nor U93 (N_93,In_108,In_107);
nand U94 (N_94,In_344,In_119);
nand U95 (N_95,In_427,N_26);
nor U96 (N_96,In_29,In_494);
or U97 (N_97,In_254,In_126);
and U98 (N_98,In_400,In_382);
nand U99 (N_99,In_103,In_4);
or U100 (N_100,In_323,In_370);
or U101 (N_101,In_218,N_33);
nand U102 (N_102,In_217,In_460);
and U103 (N_103,In_355,In_92);
nor U104 (N_104,In_315,N_14);
nand U105 (N_105,N_25,In_144);
and U106 (N_106,In_320,N_22);
nor U107 (N_107,In_74,In_36);
or U108 (N_108,In_45,N_13);
or U109 (N_109,In_135,In_15);
and U110 (N_110,In_417,N_16);
nand U111 (N_111,In_374,In_192);
nor U112 (N_112,In_61,In_68);
and U113 (N_113,In_7,In_175);
or U114 (N_114,In_137,In_227);
or U115 (N_115,In_142,In_208);
or U116 (N_116,In_393,In_428);
nor U117 (N_117,In_259,In_49);
nand U118 (N_118,In_171,In_271);
nor U119 (N_119,N_15,In_285);
and U120 (N_120,In_237,In_292);
nand U121 (N_121,In_461,In_24);
and U122 (N_122,In_406,N_42);
nand U123 (N_123,N_12,In_397);
or U124 (N_124,N_35,In_196);
and U125 (N_125,N_60,N_98);
nor U126 (N_126,In_336,N_105);
nand U127 (N_127,In_389,In_429);
and U128 (N_128,N_59,In_398);
and U129 (N_129,N_96,In_282);
and U130 (N_130,N_69,N_49);
or U131 (N_131,In_22,In_112);
nand U132 (N_132,In_401,In_392);
and U133 (N_133,N_108,N_41);
and U134 (N_134,In_63,N_68);
or U135 (N_135,N_65,N_50);
nand U136 (N_136,In_173,In_312);
nor U137 (N_137,N_63,In_220);
and U138 (N_138,In_321,N_78);
nand U139 (N_139,N_19,In_48);
and U140 (N_140,In_246,In_54);
nand U141 (N_141,In_371,In_482);
nand U142 (N_142,In_447,In_479);
nand U143 (N_143,N_28,In_367);
nor U144 (N_144,In_202,In_133);
nor U145 (N_145,In_154,N_24);
nor U146 (N_146,In_322,N_21);
and U147 (N_147,N_48,N_104);
and U148 (N_148,In_317,In_284);
xnor U149 (N_149,In_195,In_493);
nor U150 (N_150,In_216,N_47);
nor U151 (N_151,In_234,In_174);
and U152 (N_152,N_72,In_430);
nor U153 (N_153,In_440,In_286);
nand U154 (N_154,In_396,In_419);
nor U155 (N_155,N_64,In_466);
nor U156 (N_156,In_178,In_5);
or U157 (N_157,N_97,In_228);
or U158 (N_158,In_316,In_130);
nor U159 (N_159,In_70,N_0);
or U160 (N_160,In_387,In_481);
nor U161 (N_161,In_139,N_110);
nand U162 (N_162,In_28,In_310);
and U163 (N_163,In_177,N_107);
or U164 (N_164,In_327,N_109);
or U165 (N_165,In_380,In_250);
and U166 (N_166,In_294,In_467);
or U167 (N_167,In_131,N_79);
nor U168 (N_168,In_452,In_52);
nor U169 (N_169,In_211,N_44);
nor U170 (N_170,In_341,N_71);
nand U171 (N_171,N_7,In_129);
and U172 (N_172,N_55,In_26);
nor U173 (N_173,N_62,In_104);
nor U174 (N_174,In_265,In_134);
and U175 (N_175,N_119,In_106);
or U176 (N_176,In_13,In_421);
nand U177 (N_177,In_47,In_224);
nand U178 (N_178,In_33,In_325);
nor U179 (N_179,In_230,In_241);
and U180 (N_180,N_91,In_257);
nand U181 (N_181,N_29,In_96);
nand U182 (N_182,N_170,In_181);
or U183 (N_183,In_449,N_88);
or U184 (N_184,In_12,In_93);
nor U185 (N_185,In_164,In_302);
and U186 (N_186,N_133,In_53);
nor U187 (N_187,In_300,N_112);
and U188 (N_188,In_110,In_376);
or U189 (N_189,N_56,In_275);
or U190 (N_190,In_184,N_87);
and U191 (N_191,N_73,N_4);
xnor U192 (N_192,In_95,N_136);
and U193 (N_193,In_497,N_83);
nand U194 (N_194,N_137,In_40);
xnor U195 (N_195,In_55,In_469);
nand U196 (N_196,In_465,In_122);
and U197 (N_197,N_129,In_141);
or U198 (N_198,In_357,N_160);
nand U199 (N_199,In_471,In_306);
and U200 (N_200,In_79,In_102);
nand U201 (N_201,In_289,In_80);
nand U202 (N_202,In_476,N_142);
or U203 (N_203,N_114,N_70);
nand U204 (N_204,In_120,In_160);
nor U205 (N_205,N_126,In_27);
nand U206 (N_206,In_484,In_309);
and U207 (N_207,In_290,In_157);
nand U208 (N_208,In_1,N_154);
or U209 (N_209,In_231,N_143);
or U210 (N_210,In_240,In_200);
nor U211 (N_211,N_149,In_189);
nor U212 (N_212,In_125,N_81);
nand U213 (N_213,N_165,In_372);
nand U214 (N_214,N_115,In_248);
nand U215 (N_215,In_291,In_283);
or U216 (N_216,N_111,In_186);
or U217 (N_217,In_313,In_256);
or U218 (N_218,In_431,N_135);
nand U219 (N_219,In_235,In_356);
or U220 (N_220,N_118,In_251);
and U221 (N_221,N_161,N_138);
or U222 (N_222,N_172,N_124);
nand U223 (N_223,In_287,N_173);
nor U224 (N_224,N_75,In_477);
nand U225 (N_225,N_134,In_50);
nor U226 (N_226,In_123,N_89);
and U227 (N_227,N_166,In_148);
or U228 (N_228,In_232,In_249);
and U229 (N_229,In_89,N_146);
nor U230 (N_230,In_432,In_42);
nor U231 (N_231,In_475,In_56);
nand U232 (N_232,In_111,N_128);
nand U233 (N_233,N_66,N_23);
nor U234 (N_234,N_106,In_9);
nor U235 (N_235,In_386,In_14);
nor U236 (N_236,In_451,In_415);
or U237 (N_237,N_11,N_94);
nand U238 (N_238,N_120,In_450);
nand U239 (N_239,In_468,In_362);
or U240 (N_240,In_72,In_495);
nor U241 (N_241,In_162,In_359);
and U242 (N_242,N_130,N_145);
nor U243 (N_243,N_223,In_67);
or U244 (N_244,N_191,N_167);
or U245 (N_245,N_151,N_3);
or U246 (N_246,N_10,N_122);
nor U247 (N_247,N_155,N_239);
and U248 (N_248,In_348,In_116);
nor U249 (N_249,In_143,In_84);
nand U250 (N_250,In_478,In_318);
or U251 (N_251,In_222,In_472);
or U252 (N_252,In_330,In_349);
and U253 (N_253,In_422,N_90);
and U254 (N_254,In_10,N_37);
or U255 (N_255,In_59,In_337);
or U256 (N_256,In_295,N_188);
nor U257 (N_257,In_30,N_95);
nor U258 (N_258,N_202,In_252);
and U259 (N_259,N_101,In_153);
or U260 (N_260,In_399,N_17);
or U261 (N_261,In_87,In_457);
and U262 (N_262,In_458,In_333);
or U263 (N_263,N_205,In_270);
xnor U264 (N_264,N_211,N_57);
or U265 (N_265,In_365,In_145);
nor U266 (N_266,N_231,N_18);
nor U267 (N_267,N_147,In_441);
and U268 (N_268,N_102,In_38);
and U269 (N_269,In_101,N_20);
or U270 (N_270,In_147,In_390);
and U271 (N_271,N_159,N_117);
xnor U272 (N_272,In_193,In_25);
nor U273 (N_273,In_114,In_411);
xnor U274 (N_274,In_453,In_442);
or U275 (N_275,N_204,In_117);
or U276 (N_276,In_331,N_212);
or U277 (N_277,N_179,N_200);
nand U278 (N_278,N_220,N_150);
nand U279 (N_279,N_5,In_197);
or U280 (N_280,N_80,N_203);
nand U281 (N_281,N_226,N_113);
nand U282 (N_282,N_27,N_183);
nand U283 (N_283,In_366,In_496);
nor U284 (N_284,In_381,In_403);
nand U285 (N_285,N_198,In_152);
and U286 (N_286,In_434,In_247);
nor U287 (N_287,N_208,N_222);
or U288 (N_288,N_169,N_132);
and U289 (N_289,N_34,N_46);
and U290 (N_290,N_92,In_437);
and U291 (N_291,N_121,In_91);
or U292 (N_292,N_235,In_319);
nand U293 (N_293,In_146,N_215);
and U294 (N_294,N_152,N_224);
and U295 (N_295,N_176,N_38);
or U296 (N_296,N_43,N_181);
nor U297 (N_297,N_187,N_67);
nor U298 (N_298,In_0,In_324);
and U299 (N_299,N_230,In_64);
and U300 (N_300,N_175,N_162);
nor U301 (N_301,In_190,N_278);
and U302 (N_302,N_76,N_157);
or U303 (N_303,N_185,N_282);
and U304 (N_304,N_182,N_77);
xnor U305 (N_305,N_156,N_276);
nand U306 (N_306,N_103,In_314);
and U307 (N_307,N_255,In_18);
and U308 (N_308,N_177,N_229);
xor U309 (N_309,N_242,In_75);
nor U310 (N_310,In_198,In_238);
and U311 (N_311,In_37,In_140);
nand U312 (N_312,N_272,In_172);
and U313 (N_313,N_61,N_264);
nand U314 (N_314,N_296,In_418);
nand U315 (N_315,N_74,In_77);
nand U316 (N_316,N_240,In_328);
nor U317 (N_317,N_241,N_299);
nand U318 (N_318,In_276,N_271);
nand U319 (N_319,N_189,N_297);
nand U320 (N_320,N_144,N_195);
nor U321 (N_321,N_284,In_39);
and U322 (N_322,N_256,N_171);
nor U323 (N_323,In_384,N_263);
nand U324 (N_324,N_243,N_273);
and U325 (N_325,N_214,In_296);
or U326 (N_326,N_269,N_116);
or U327 (N_327,N_140,N_199);
nand U328 (N_328,N_186,N_158);
nor U329 (N_329,N_8,N_270);
or U330 (N_330,N_190,In_209);
nor U331 (N_331,N_100,N_31);
nand U332 (N_332,In_71,N_123);
nand U333 (N_333,N_209,N_194);
nor U334 (N_334,N_293,N_236);
or U335 (N_335,In_407,N_86);
or U336 (N_336,N_217,N_287);
nor U337 (N_337,N_210,N_251);
nor U338 (N_338,N_252,N_234);
nor U339 (N_339,N_219,N_193);
and U340 (N_340,N_267,N_253);
or U341 (N_341,N_201,In_463);
and U342 (N_342,In_151,In_311);
and U343 (N_343,N_196,N_285);
nor U344 (N_344,N_125,In_159);
and U345 (N_345,In_73,In_360);
and U346 (N_346,In_78,In_499);
or U347 (N_347,In_263,In_279);
or U348 (N_348,In_44,In_205);
or U349 (N_349,In_156,In_352);
nor U350 (N_350,N_82,N_184);
nand U351 (N_351,In_158,N_54);
nand U352 (N_352,N_294,N_238);
nand U353 (N_353,N_168,N_221);
nand U354 (N_354,In_448,N_274);
nand U355 (N_355,N_85,N_148);
nand U356 (N_356,N_2,N_131);
and U357 (N_357,In_244,In_339);
or U358 (N_358,In_308,N_257);
nor U359 (N_359,N_254,N_197);
xnor U360 (N_360,In_404,N_343);
nor U361 (N_361,N_245,N_232);
and U362 (N_362,N_351,N_266);
or U363 (N_363,N_325,N_93);
nor U364 (N_364,In_438,N_354);
or U365 (N_365,N_340,N_352);
nor U366 (N_366,In_182,N_317);
nand U367 (N_367,N_304,N_213);
or U368 (N_368,N_178,N_356);
nand U369 (N_369,In_273,N_330);
nor U370 (N_370,N_246,N_233);
nand U371 (N_371,N_99,N_225);
nand U372 (N_372,N_348,N_279);
or U373 (N_373,N_289,N_316);
nand U374 (N_374,N_291,In_16);
nor U375 (N_375,In_3,In_163);
nand U376 (N_376,In_255,N_312);
and U377 (N_377,N_308,N_174);
or U378 (N_378,In_260,N_335);
or U379 (N_379,N_206,N_127);
nand U380 (N_380,N_237,N_228);
nor U381 (N_381,N_328,N_265);
or U382 (N_382,N_292,N_290);
nor U383 (N_383,N_345,N_346);
nor U384 (N_384,N_163,N_319);
nand U385 (N_385,N_342,N_277);
nand U386 (N_386,N_153,In_20);
and U387 (N_387,N_216,N_298);
nor U388 (N_388,N_318,In_301);
nor U389 (N_389,In_136,N_281);
nor U390 (N_390,In_85,N_344);
or U391 (N_391,N_337,N_327);
nand U392 (N_392,In_8,N_259);
or U393 (N_393,N_244,N_84);
nor U394 (N_394,N_336,N_306);
and U395 (N_395,N_341,N_313);
nor U396 (N_396,N_314,N_180);
nand U397 (N_397,In_179,In_351);
or U398 (N_398,N_275,In_191);
nor U399 (N_399,N_258,In_346);
and U400 (N_400,In_128,N_283);
and U401 (N_401,N_358,N_350);
and U402 (N_402,N_309,In_347);
nor U403 (N_403,N_192,N_268);
xnor U404 (N_404,N_302,N_326);
nand U405 (N_405,In_436,N_288);
and U406 (N_406,N_300,N_303);
nand U407 (N_407,N_250,In_272);
and U408 (N_408,N_349,N_310);
nand U409 (N_409,N_260,N_249);
nand U410 (N_410,N_332,N_320);
or U411 (N_411,N_359,N_331);
nor U412 (N_412,N_301,N_355);
nand U413 (N_413,N_334,N_322);
nand U414 (N_414,N_295,N_218);
nand U415 (N_415,N_307,N_315);
or U416 (N_416,N_9,N_286);
and U417 (N_417,N_207,N_321);
nor U418 (N_418,N_139,N_333);
and U419 (N_419,N_338,N_261);
and U420 (N_420,N_367,N_397);
nor U421 (N_421,N_372,In_304);
and U422 (N_422,N_227,N_366);
xor U423 (N_423,N_388,N_377);
nor U424 (N_424,N_374,N_311);
xor U425 (N_425,N_419,N_400);
or U426 (N_426,N_373,N_382);
nand U427 (N_427,N_363,N_375);
and U428 (N_428,N_141,N_247);
or U429 (N_429,N_365,N_403);
or U430 (N_430,N_323,N_396);
nor U431 (N_431,N_248,N_324);
nor U432 (N_432,N_395,N_368);
or U433 (N_433,N_418,N_407);
and U434 (N_434,N_364,N_371);
and U435 (N_435,N_357,N_392);
nor U436 (N_436,N_409,N_361);
and U437 (N_437,N_369,N_412);
nor U438 (N_438,N_386,In_267);
or U439 (N_439,N_353,N_390);
or U440 (N_440,N_415,N_347);
nor U441 (N_441,N_381,N_417);
nand U442 (N_442,N_399,N_389);
or U443 (N_443,N_384,N_380);
nor U444 (N_444,In_210,N_404);
nand U445 (N_445,N_280,N_329);
nand U446 (N_446,N_406,N_164);
nand U447 (N_447,N_413,N_416);
or U448 (N_448,N_339,N_410);
nor U449 (N_449,N_383,N_379);
nand U450 (N_450,N_362,N_401);
nor U451 (N_451,N_402,N_262);
and U452 (N_452,N_370,In_299);
nor U453 (N_453,N_393,N_408);
and U454 (N_454,N_305,N_360);
and U455 (N_455,N_378,N_387);
xor U456 (N_456,N_376,N_394);
or U457 (N_457,N_411,N_414);
nor U458 (N_458,N_391,N_398);
nor U459 (N_459,N_405,N_385);
xor U460 (N_460,N_400,N_384);
nand U461 (N_461,N_412,N_404);
and U462 (N_462,N_280,N_305);
nand U463 (N_463,N_262,N_379);
or U464 (N_464,N_366,N_412);
nor U465 (N_465,N_412,N_400);
nand U466 (N_466,N_403,N_386);
or U467 (N_467,N_396,N_390);
nand U468 (N_468,N_374,N_407);
or U469 (N_469,N_375,N_386);
nand U470 (N_470,N_353,N_393);
or U471 (N_471,N_357,N_415);
and U472 (N_472,N_399,N_415);
and U473 (N_473,N_402,N_357);
and U474 (N_474,In_210,N_364);
and U475 (N_475,N_227,N_390);
nand U476 (N_476,In_267,N_405);
or U477 (N_477,N_323,N_390);
and U478 (N_478,N_374,N_413);
and U479 (N_479,N_386,N_376);
xor U480 (N_480,N_446,N_443);
nor U481 (N_481,N_455,N_423);
nand U482 (N_482,N_422,N_465);
or U483 (N_483,N_434,N_438);
and U484 (N_484,N_457,N_475);
and U485 (N_485,N_432,N_468);
xor U486 (N_486,N_431,N_435);
or U487 (N_487,N_449,N_444);
nand U488 (N_488,N_436,N_428);
nand U489 (N_489,N_456,N_441);
nor U490 (N_490,N_472,N_448);
or U491 (N_491,N_460,N_462);
or U492 (N_492,N_447,N_445);
or U493 (N_493,N_450,N_430);
or U494 (N_494,N_461,N_442);
and U495 (N_495,N_473,N_439);
or U496 (N_496,N_459,N_437);
nand U497 (N_497,N_425,N_474);
and U498 (N_498,N_429,N_467);
nand U499 (N_499,N_478,N_471);
nor U500 (N_500,N_433,N_454);
or U501 (N_501,N_420,N_458);
and U502 (N_502,N_477,N_464);
nor U503 (N_503,N_421,N_427);
or U504 (N_504,N_440,N_470);
nor U505 (N_505,N_451,N_476);
nor U506 (N_506,N_466,N_426);
or U507 (N_507,N_469,N_479);
nand U508 (N_508,N_452,N_424);
or U509 (N_509,N_463,N_453);
nand U510 (N_510,N_451,N_420);
nand U511 (N_511,N_420,N_425);
nand U512 (N_512,N_427,N_447);
or U513 (N_513,N_465,N_478);
nand U514 (N_514,N_460,N_423);
nor U515 (N_515,N_447,N_470);
nand U516 (N_516,N_444,N_430);
nor U517 (N_517,N_453,N_477);
nand U518 (N_518,N_472,N_431);
or U519 (N_519,N_470,N_435);
nand U520 (N_520,N_461,N_474);
and U521 (N_521,N_442,N_444);
nor U522 (N_522,N_452,N_473);
nand U523 (N_523,N_465,N_463);
nor U524 (N_524,N_461,N_478);
xor U525 (N_525,N_432,N_471);
nor U526 (N_526,N_433,N_421);
nor U527 (N_527,N_473,N_465);
and U528 (N_528,N_451,N_432);
or U529 (N_529,N_471,N_458);
nor U530 (N_530,N_450,N_474);
nand U531 (N_531,N_435,N_429);
or U532 (N_532,N_435,N_477);
nor U533 (N_533,N_460,N_463);
nor U534 (N_534,N_457,N_435);
nand U535 (N_535,N_474,N_466);
or U536 (N_536,N_473,N_425);
nand U537 (N_537,N_475,N_467);
xnor U538 (N_538,N_429,N_447);
or U539 (N_539,N_431,N_428);
and U540 (N_540,N_496,N_518);
nor U541 (N_541,N_528,N_514);
and U542 (N_542,N_538,N_486);
or U543 (N_543,N_539,N_503);
or U544 (N_544,N_505,N_525);
and U545 (N_545,N_495,N_526);
nand U546 (N_546,N_509,N_488);
xor U547 (N_547,N_516,N_510);
or U548 (N_548,N_533,N_492);
nor U549 (N_549,N_480,N_494);
or U550 (N_550,N_522,N_532);
nor U551 (N_551,N_512,N_497);
or U552 (N_552,N_524,N_519);
nor U553 (N_553,N_530,N_487);
nand U554 (N_554,N_513,N_481);
nor U555 (N_555,N_523,N_537);
nor U556 (N_556,N_527,N_500);
nand U557 (N_557,N_511,N_535);
nand U558 (N_558,N_520,N_485);
nand U559 (N_559,N_506,N_517);
and U560 (N_560,N_529,N_490);
or U561 (N_561,N_502,N_498);
or U562 (N_562,N_531,N_508);
or U563 (N_563,N_507,N_521);
or U564 (N_564,N_501,N_482);
and U565 (N_565,N_499,N_504);
or U566 (N_566,N_491,N_483);
nand U567 (N_567,N_536,N_493);
nand U568 (N_568,N_534,N_489);
or U569 (N_569,N_515,N_484);
and U570 (N_570,N_517,N_511);
nor U571 (N_571,N_522,N_492);
or U572 (N_572,N_535,N_518);
and U573 (N_573,N_494,N_516);
or U574 (N_574,N_486,N_512);
nor U575 (N_575,N_510,N_507);
and U576 (N_576,N_480,N_482);
nand U577 (N_577,N_501,N_494);
nor U578 (N_578,N_530,N_499);
or U579 (N_579,N_486,N_517);
or U580 (N_580,N_511,N_499);
nand U581 (N_581,N_510,N_498);
nand U582 (N_582,N_485,N_493);
or U583 (N_583,N_529,N_524);
xor U584 (N_584,N_512,N_518);
and U585 (N_585,N_526,N_508);
and U586 (N_586,N_485,N_525);
nor U587 (N_587,N_519,N_487);
or U588 (N_588,N_512,N_513);
nor U589 (N_589,N_509,N_482);
or U590 (N_590,N_529,N_538);
nand U591 (N_591,N_511,N_489);
xor U592 (N_592,N_532,N_526);
or U593 (N_593,N_537,N_490);
nor U594 (N_594,N_525,N_534);
and U595 (N_595,N_481,N_521);
nand U596 (N_596,N_483,N_507);
nand U597 (N_597,N_508,N_503);
nand U598 (N_598,N_529,N_497);
nand U599 (N_599,N_520,N_510);
or U600 (N_600,N_588,N_594);
nor U601 (N_601,N_558,N_555);
and U602 (N_602,N_574,N_550);
and U603 (N_603,N_597,N_576);
or U604 (N_604,N_584,N_592);
xor U605 (N_605,N_587,N_554);
nand U606 (N_606,N_563,N_595);
and U607 (N_607,N_582,N_545);
or U608 (N_608,N_571,N_591);
nand U609 (N_609,N_564,N_559);
and U610 (N_610,N_569,N_566);
and U611 (N_611,N_542,N_540);
or U612 (N_612,N_546,N_581);
or U613 (N_613,N_543,N_572);
or U614 (N_614,N_557,N_583);
and U615 (N_615,N_596,N_575);
nor U616 (N_616,N_580,N_549);
nand U617 (N_617,N_552,N_551);
xnor U618 (N_618,N_547,N_599);
nand U619 (N_619,N_560,N_567);
and U620 (N_620,N_541,N_548);
nor U621 (N_621,N_565,N_585);
or U622 (N_622,N_561,N_586);
nand U623 (N_623,N_598,N_562);
nor U624 (N_624,N_570,N_589);
or U625 (N_625,N_568,N_593);
nor U626 (N_626,N_590,N_577);
nor U627 (N_627,N_544,N_553);
or U628 (N_628,N_578,N_579);
or U629 (N_629,N_573,N_556);
or U630 (N_630,N_540,N_599);
nand U631 (N_631,N_545,N_561);
or U632 (N_632,N_578,N_590);
or U633 (N_633,N_567,N_555);
nor U634 (N_634,N_596,N_548);
or U635 (N_635,N_552,N_548);
or U636 (N_636,N_576,N_584);
nor U637 (N_637,N_576,N_545);
nand U638 (N_638,N_549,N_570);
nand U639 (N_639,N_585,N_551);
nor U640 (N_640,N_569,N_583);
nor U641 (N_641,N_553,N_554);
nor U642 (N_642,N_599,N_589);
nor U643 (N_643,N_578,N_572);
nand U644 (N_644,N_579,N_566);
and U645 (N_645,N_569,N_548);
nand U646 (N_646,N_550,N_596);
or U647 (N_647,N_578,N_587);
nor U648 (N_648,N_567,N_586);
nor U649 (N_649,N_570,N_583);
nor U650 (N_650,N_558,N_595);
and U651 (N_651,N_550,N_569);
nand U652 (N_652,N_564,N_578);
nand U653 (N_653,N_549,N_544);
or U654 (N_654,N_563,N_593);
nand U655 (N_655,N_562,N_557);
or U656 (N_656,N_581,N_559);
or U657 (N_657,N_583,N_598);
or U658 (N_658,N_584,N_556);
nand U659 (N_659,N_577,N_569);
nand U660 (N_660,N_643,N_612);
nand U661 (N_661,N_618,N_645);
or U662 (N_662,N_617,N_651);
or U663 (N_663,N_638,N_613);
or U664 (N_664,N_647,N_657);
nand U665 (N_665,N_608,N_626);
or U666 (N_666,N_639,N_640);
and U667 (N_667,N_616,N_635);
and U668 (N_668,N_604,N_607);
or U669 (N_669,N_605,N_601);
nand U670 (N_670,N_614,N_630);
nor U671 (N_671,N_655,N_627);
nand U672 (N_672,N_625,N_624);
xnor U673 (N_673,N_631,N_646);
nand U674 (N_674,N_656,N_603);
or U675 (N_675,N_659,N_644);
nand U676 (N_676,N_648,N_637);
or U677 (N_677,N_632,N_602);
nand U678 (N_678,N_629,N_652);
and U679 (N_679,N_650,N_615);
or U680 (N_680,N_628,N_641);
or U681 (N_681,N_642,N_633);
nor U682 (N_682,N_636,N_654);
xnor U683 (N_683,N_622,N_600);
and U684 (N_684,N_634,N_620);
and U685 (N_685,N_623,N_611);
xnor U686 (N_686,N_610,N_606);
nand U687 (N_687,N_649,N_609);
or U688 (N_688,N_621,N_653);
and U689 (N_689,N_619,N_658);
nor U690 (N_690,N_610,N_628);
nand U691 (N_691,N_622,N_618);
or U692 (N_692,N_604,N_655);
or U693 (N_693,N_634,N_618);
or U694 (N_694,N_616,N_633);
and U695 (N_695,N_616,N_638);
and U696 (N_696,N_648,N_617);
nand U697 (N_697,N_647,N_601);
nand U698 (N_698,N_605,N_607);
and U699 (N_699,N_627,N_612);
and U700 (N_700,N_654,N_614);
or U701 (N_701,N_655,N_644);
and U702 (N_702,N_617,N_619);
and U703 (N_703,N_643,N_659);
and U704 (N_704,N_659,N_654);
and U705 (N_705,N_630,N_652);
nand U706 (N_706,N_614,N_631);
nor U707 (N_707,N_635,N_658);
and U708 (N_708,N_631,N_638);
and U709 (N_709,N_631,N_626);
nand U710 (N_710,N_603,N_614);
xnor U711 (N_711,N_609,N_652);
and U712 (N_712,N_607,N_618);
nor U713 (N_713,N_600,N_650);
nor U714 (N_714,N_644,N_637);
or U715 (N_715,N_650,N_637);
or U716 (N_716,N_639,N_638);
and U717 (N_717,N_647,N_621);
nor U718 (N_718,N_645,N_615);
nand U719 (N_719,N_636,N_602);
or U720 (N_720,N_681,N_684);
xnor U721 (N_721,N_718,N_690);
nor U722 (N_722,N_694,N_688);
and U723 (N_723,N_669,N_708);
nand U724 (N_724,N_719,N_661);
or U725 (N_725,N_695,N_689);
nand U726 (N_726,N_706,N_686);
and U727 (N_727,N_698,N_663);
or U728 (N_728,N_701,N_692);
or U729 (N_729,N_710,N_693);
nor U730 (N_730,N_677,N_680);
nand U731 (N_731,N_716,N_672);
or U732 (N_732,N_682,N_673);
nand U733 (N_733,N_685,N_707);
nand U734 (N_734,N_699,N_667);
nor U735 (N_735,N_691,N_665);
or U736 (N_736,N_664,N_670);
and U737 (N_737,N_711,N_702);
or U738 (N_738,N_666,N_679);
nand U739 (N_739,N_668,N_704);
or U740 (N_740,N_678,N_683);
and U741 (N_741,N_715,N_696);
and U742 (N_742,N_712,N_662);
or U743 (N_743,N_709,N_697);
nand U744 (N_744,N_713,N_687);
nand U745 (N_745,N_703,N_675);
or U746 (N_746,N_674,N_700);
or U747 (N_747,N_660,N_714);
and U748 (N_748,N_717,N_705);
nor U749 (N_749,N_671,N_676);
or U750 (N_750,N_711,N_665);
nand U751 (N_751,N_665,N_705);
and U752 (N_752,N_691,N_694);
nor U753 (N_753,N_687,N_696);
nor U754 (N_754,N_699,N_675);
and U755 (N_755,N_666,N_712);
and U756 (N_756,N_665,N_672);
nor U757 (N_757,N_699,N_664);
or U758 (N_758,N_663,N_671);
nor U759 (N_759,N_705,N_697);
or U760 (N_760,N_697,N_684);
nor U761 (N_761,N_712,N_703);
or U762 (N_762,N_666,N_673);
xnor U763 (N_763,N_708,N_678);
nor U764 (N_764,N_674,N_692);
nor U765 (N_765,N_700,N_667);
nand U766 (N_766,N_708,N_713);
or U767 (N_767,N_681,N_661);
or U768 (N_768,N_664,N_689);
and U769 (N_769,N_697,N_700);
nor U770 (N_770,N_688,N_692);
or U771 (N_771,N_712,N_704);
nor U772 (N_772,N_663,N_711);
nand U773 (N_773,N_712,N_697);
nor U774 (N_774,N_705,N_709);
or U775 (N_775,N_666,N_676);
nand U776 (N_776,N_675,N_714);
nand U777 (N_777,N_662,N_671);
and U778 (N_778,N_660,N_699);
nand U779 (N_779,N_699,N_678);
and U780 (N_780,N_727,N_766);
nor U781 (N_781,N_722,N_721);
nand U782 (N_782,N_767,N_725);
and U783 (N_783,N_732,N_764);
nor U784 (N_784,N_775,N_746);
nor U785 (N_785,N_747,N_759);
and U786 (N_786,N_730,N_763);
or U787 (N_787,N_726,N_737);
or U788 (N_788,N_762,N_768);
or U789 (N_789,N_748,N_745);
nand U790 (N_790,N_761,N_757);
nand U791 (N_791,N_774,N_740);
nor U792 (N_792,N_723,N_738);
nor U793 (N_793,N_734,N_749);
nand U794 (N_794,N_756,N_720);
or U795 (N_795,N_754,N_779);
and U796 (N_796,N_729,N_731);
nor U797 (N_797,N_742,N_728);
and U798 (N_798,N_755,N_772);
nand U799 (N_799,N_751,N_744);
nand U800 (N_800,N_752,N_773);
nor U801 (N_801,N_770,N_760);
nand U802 (N_802,N_724,N_743);
and U803 (N_803,N_753,N_777);
nand U804 (N_804,N_758,N_750);
or U805 (N_805,N_769,N_739);
nor U806 (N_806,N_771,N_741);
nand U807 (N_807,N_733,N_735);
nand U808 (N_808,N_778,N_776);
or U809 (N_809,N_736,N_765);
and U810 (N_810,N_731,N_756);
and U811 (N_811,N_765,N_721);
nand U812 (N_812,N_754,N_767);
nor U813 (N_813,N_730,N_739);
nor U814 (N_814,N_742,N_771);
and U815 (N_815,N_764,N_776);
or U816 (N_816,N_761,N_767);
or U817 (N_817,N_739,N_738);
or U818 (N_818,N_740,N_739);
nor U819 (N_819,N_723,N_753);
and U820 (N_820,N_770,N_779);
or U821 (N_821,N_773,N_777);
and U822 (N_822,N_740,N_742);
and U823 (N_823,N_772,N_722);
nor U824 (N_824,N_726,N_738);
or U825 (N_825,N_734,N_742);
or U826 (N_826,N_729,N_774);
or U827 (N_827,N_738,N_767);
or U828 (N_828,N_760,N_732);
or U829 (N_829,N_740,N_755);
nor U830 (N_830,N_749,N_738);
nor U831 (N_831,N_756,N_730);
or U832 (N_832,N_777,N_774);
nor U833 (N_833,N_762,N_767);
nand U834 (N_834,N_740,N_767);
or U835 (N_835,N_769,N_772);
nor U836 (N_836,N_729,N_773);
nand U837 (N_837,N_746,N_776);
nand U838 (N_838,N_738,N_757);
or U839 (N_839,N_736,N_752);
or U840 (N_840,N_834,N_784);
nor U841 (N_841,N_817,N_786);
nand U842 (N_842,N_780,N_811);
nor U843 (N_843,N_790,N_833);
nor U844 (N_844,N_823,N_813);
nand U845 (N_845,N_793,N_807);
nor U846 (N_846,N_802,N_809);
or U847 (N_847,N_822,N_787);
xor U848 (N_848,N_781,N_791);
and U849 (N_849,N_812,N_800);
and U850 (N_850,N_806,N_820);
nand U851 (N_851,N_827,N_788);
nor U852 (N_852,N_785,N_831);
nor U853 (N_853,N_797,N_815);
or U854 (N_854,N_824,N_792);
xnor U855 (N_855,N_799,N_805);
or U856 (N_856,N_839,N_818);
and U857 (N_857,N_835,N_810);
nand U858 (N_858,N_782,N_816);
nor U859 (N_859,N_796,N_801);
nand U860 (N_860,N_838,N_804);
or U861 (N_861,N_819,N_795);
nor U862 (N_862,N_830,N_837);
nand U863 (N_863,N_836,N_825);
or U864 (N_864,N_829,N_798);
or U865 (N_865,N_828,N_821);
and U866 (N_866,N_803,N_794);
or U867 (N_867,N_808,N_814);
or U868 (N_868,N_783,N_832);
xnor U869 (N_869,N_826,N_789);
nand U870 (N_870,N_799,N_824);
and U871 (N_871,N_790,N_824);
nand U872 (N_872,N_826,N_780);
and U873 (N_873,N_822,N_815);
and U874 (N_874,N_793,N_785);
or U875 (N_875,N_833,N_832);
and U876 (N_876,N_807,N_817);
and U877 (N_877,N_832,N_799);
nor U878 (N_878,N_821,N_798);
xnor U879 (N_879,N_793,N_816);
nand U880 (N_880,N_792,N_804);
and U881 (N_881,N_808,N_792);
and U882 (N_882,N_802,N_793);
nand U883 (N_883,N_821,N_835);
or U884 (N_884,N_830,N_826);
nor U885 (N_885,N_810,N_824);
nand U886 (N_886,N_815,N_798);
and U887 (N_887,N_785,N_821);
nor U888 (N_888,N_783,N_818);
nand U889 (N_889,N_793,N_835);
or U890 (N_890,N_815,N_805);
nor U891 (N_891,N_805,N_838);
nand U892 (N_892,N_810,N_801);
or U893 (N_893,N_783,N_799);
or U894 (N_894,N_827,N_793);
or U895 (N_895,N_839,N_833);
nand U896 (N_896,N_818,N_792);
and U897 (N_897,N_837,N_839);
nand U898 (N_898,N_813,N_825);
nand U899 (N_899,N_828,N_817);
nor U900 (N_900,N_842,N_872);
nand U901 (N_901,N_879,N_878);
nand U902 (N_902,N_846,N_888);
nor U903 (N_903,N_859,N_860);
xnor U904 (N_904,N_857,N_880);
nand U905 (N_905,N_892,N_847);
nand U906 (N_906,N_848,N_877);
or U907 (N_907,N_866,N_887);
nor U908 (N_908,N_840,N_855);
or U909 (N_909,N_881,N_841);
and U910 (N_910,N_899,N_885);
nor U911 (N_911,N_886,N_894);
or U912 (N_912,N_844,N_865);
nand U913 (N_913,N_861,N_871);
and U914 (N_914,N_889,N_875);
and U915 (N_915,N_896,N_870);
nand U916 (N_916,N_884,N_876);
and U917 (N_917,N_849,N_895);
nand U918 (N_918,N_854,N_897);
and U919 (N_919,N_850,N_874);
nand U920 (N_920,N_890,N_863);
and U921 (N_921,N_856,N_868);
or U922 (N_922,N_858,N_891);
or U923 (N_923,N_864,N_893);
nand U924 (N_924,N_867,N_851);
or U925 (N_925,N_845,N_883);
nand U926 (N_926,N_869,N_852);
and U927 (N_927,N_862,N_843);
nand U928 (N_928,N_898,N_873);
and U929 (N_929,N_853,N_882);
nand U930 (N_930,N_845,N_860);
and U931 (N_931,N_878,N_840);
nand U932 (N_932,N_891,N_850);
and U933 (N_933,N_857,N_870);
nand U934 (N_934,N_875,N_886);
xor U935 (N_935,N_850,N_897);
xor U936 (N_936,N_887,N_879);
nor U937 (N_937,N_899,N_867);
or U938 (N_938,N_864,N_895);
nand U939 (N_939,N_873,N_874);
nor U940 (N_940,N_877,N_842);
nand U941 (N_941,N_873,N_879);
and U942 (N_942,N_859,N_885);
or U943 (N_943,N_858,N_882);
nand U944 (N_944,N_861,N_856);
nor U945 (N_945,N_890,N_884);
and U946 (N_946,N_899,N_897);
or U947 (N_947,N_862,N_889);
or U948 (N_948,N_895,N_841);
nand U949 (N_949,N_882,N_844);
and U950 (N_950,N_872,N_895);
and U951 (N_951,N_872,N_892);
nor U952 (N_952,N_892,N_864);
or U953 (N_953,N_892,N_851);
nor U954 (N_954,N_890,N_850);
and U955 (N_955,N_843,N_858);
and U956 (N_956,N_870,N_898);
and U957 (N_957,N_881,N_849);
or U958 (N_958,N_858,N_865);
and U959 (N_959,N_863,N_850);
and U960 (N_960,N_951,N_945);
nand U961 (N_961,N_920,N_940);
or U962 (N_962,N_907,N_928);
and U963 (N_963,N_934,N_926);
nand U964 (N_964,N_950,N_932);
or U965 (N_965,N_931,N_921);
or U966 (N_966,N_922,N_955);
or U967 (N_967,N_930,N_944);
nand U968 (N_968,N_909,N_915);
and U969 (N_969,N_938,N_904);
nand U970 (N_970,N_948,N_943);
and U971 (N_971,N_900,N_957);
nand U972 (N_972,N_947,N_913);
nand U973 (N_973,N_902,N_952);
nand U974 (N_974,N_954,N_942);
nor U975 (N_975,N_901,N_946);
or U976 (N_976,N_935,N_906);
or U977 (N_977,N_916,N_914);
nor U978 (N_978,N_919,N_956);
nand U979 (N_979,N_910,N_903);
or U980 (N_980,N_908,N_927);
and U981 (N_981,N_937,N_911);
and U982 (N_982,N_958,N_959);
nor U983 (N_983,N_905,N_924);
nand U984 (N_984,N_929,N_933);
nand U985 (N_985,N_917,N_918);
nor U986 (N_986,N_949,N_953);
nor U987 (N_987,N_912,N_936);
or U988 (N_988,N_923,N_941);
nand U989 (N_989,N_939,N_925);
or U990 (N_990,N_926,N_905);
or U991 (N_991,N_909,N_955);
or U992 (N_992,N_911,N_932);
or U993 (N_993,N_931,N_930);
or U994 (N_994,N_907,N_952);
xor U995 (N_995,N_939,N_912);
and U996 (N_996,N_905,N_947);
and U997 (N_997,N_927,N_940);
and U998 (N_998,N_954,N_955);
nor U999 (N_999,N_952,N_904);
or U1000 (N_1000,N_952,N_953);
nor U1001 (N_1001,N_926,N_955);
nand U1002 (N_1002,N_941,N_913);
nand U1003 (N_1003,N_957,N_940);
or U1004 (N_1004,N_941,N_905);
nor U1005 (N_1005,N_943,N_956);
nor U1006 (N_1006,N_932,N_904);
and U1007 (N_1007,N_904,N_928);
or U1008 (N_1008,N_934,N_918);
nor U1009 (N_1009,N_929,N_919);
nand U1010 (N_1010,N_943,N_946);
or U1011 (N_1011,N_955,N_908);
or U1012 (N_1012,N_953,N_900);
xnor U1013 (N_1013,N_907,N_954);
and U1014 (N_1014,N_919,N_905);
nand U1015 (N_1015,N_910,N_946);
and U1016 (N_1016,N_927,N_907);
and U1017 (N_1017,N_948,N_932);
nor U1018 (N_1018,N_905,N_913);
and U1019 (N_1019,N_948,N_944);
nor U1020 (N_1020,N_998,N_975);
nand U1021 (N_1021,N_962,N_976);
and U1022 (N_1022,N_1011,N_965);
or U1023 (N_1023,N_971,N_985);
or U1024 (N_1024,N_1013,N_988);
and U1025 (N_1025,N_1018,N_1019);
nor U1026 (N_1026,N_1002,N_997);
nor U1027 (N_1027,N_963,N_992);
nand U1028 (N_1028,N_994,N_993);
nand U1029 (N_1029,N_979,N_986);
nor U1030 (N_1030,N_1012,N_1000);
or U1031 (N_1031,N_1004,N_1014);
nor U1032 (N_1032,N_1015,N_972);
nor U1033 (N_1033,N_967,N_996);
and U1034 (N_1034,N_961,N_1007);
nand U1035 (N_1035,N_970,N_964);
nand U1036 (N_1036,N_987,N_981);
nand U1037 (N_1037,N_978,N_969);
nor U1038 (N_1038,N_989,N_990);
and U1039 (N_1039,N_983,N_973);
or U1040 (N_1040,N_968,N_1001);
and U1041 (N_1041,N_974,N_1005);
nor U1042 (N_1042,N_984,N_1016);
nand U1043 (N_1043,N_960,N_999);
nor U1044 (N_1044,N_980,N_991);
nand U1045 (N_1045,N_1008,N_995);
or U1046 (N_1046,N_1003,N_1006);
and U1047 (N_1047,N_977,N_966);
and U1048 (N_1048,N_1009,N_982);
or U1049 (N_1049,N_1010,N_1017);
and U1050 (N_1050,N_1013,N_971);
or U1051 (N_1051,N_1019,N_972);
nor U1052 (N_1052,N_1011,N_993);
and U1053 (N_1053,N_1000,N_985);
and U1054 (N_1054,N_1016,N_985);
and U1055 (N_1055,N_1007,N_984);
nor U1056 (N_1056,N_965,N_964);
nand U1057 (N_1057,N_1018,N_988);
nand U1058 (N_1058,N_963,N_995);
nand U1059 (N_1059,N_1006,N_1015);
and U1060 (N_1060,N_1012,N_974);
nor U1061 (N_1061,N_999,N_1015);
nor U1062 (N_1062,N_1008,N_1017);
and U1063 (N_1063,N_1005,N_976);
nand U1064 (N_1064,N_1012,N_991);
nor U1065 (N_1065,N_965,N_1014);
nor U1066 (N_1066,N_987,N_1006);
or U1067 (N_1067,N_960,N_985);
and U1068 (N_1068,N_964,N_988);
nor U1069 (N_1069,N_1007,N_970);
or U1070 (N_1070,N_977,N_967);
nand U1071 (N_1071,N_962,N_1006);
and U1072 (N_1072,N_1016,N_966);
nor U1073 (N_1073,N_967,N_1001);
or U1074 (N_1074,N_1000,N_989);
and U1075 (N_1075,N_965,N_984);
and U1076 (N_1076,N_962,N_991);
nand U1077 (N_1077,N_1019,N_986);
and U1078 (N_1078,N_963,N_972);
nand U1079 (N_1079,N_967,N_985);
nor U1080 (N_1080,N_1050,N_1064);
or U1081 (N_1081,N_1046,N_1025);
nor U1082 (N_1082,N_1040,N_1060);
nor U1083 (N_1083,N_1052,N_1070);
and U1084 (N_1084,N_1039,N_1074);
nor U1085 (N_1085,N_1059,N_1068);
or U1086 (N_1086,N_1057,N_1037);
and U1087 (N_1087,N_1026,N_1075);
xor U1088 (N_1088,N_1051,N_1049);
and U1089 (N_1089,N_1078,N_1033);
and U1090 (N_1090,N_1035,N_1027);
nand U1091 (N_1091,N_1042,N_1041);
nand U1092 (N_1092,N_1023,N_1045);
or U1093 (N_1093,N_1038,N_1036);
or U1094 (N_1094,N_1065,N_1072);
and U1095 (N_1095,N_1058,N_1055);
and U1096 (N_1096,N_1047,N_1030);
and U1097 (N_1097,N_1062,N_1066);
nor U1098 (N_1098,N_1043,N_1054);
nor U1099 (N_1099,N_1077,N_1024);
or U1100 (N_1100,N_1028,N_1073);
or U1101 (N_1101,N_1067,N_1076);
or U1102 (N_1102,N_1079,N_1071);
nor U1103 (N_1103,N_1029,N_1022);
and U1104 (N_1104,N_1056,N_1053);
nor U1105 (N_1105,N_1063,N_1020);
or U1106 (N_1106,N_1032,N_1034);
or U1107 (N_1107,N_1069,N_1031);
and U1108 (N_1108,N_1044,N_1021);
or U1109 (N_1109,N_1048,N_1061);
nand U1110 (N_1110,N_1055,N_1068);
and U1111 (N_1111,N_1043,N_1029);
or U1112 (N_1112,N_1045,N_1065);
and U1113 (N_1113,N_1021,N_1049);
and U1114 (N_1114,N_1066,N_1048);
nor U1115 (N_1115,N_1038,N_1078);
nor U1116 (N_1116,N_1071,N_1037);
or U1117 (N_1117,N_1061,N_1052);
nor U1118 (N_1118,N_1044,N_1079);
nor U1119 (N_1119,N_1038,N_1022);
and U1120 (N_1120,N_1041,N_1064);
and U1121 (N_1121,N_1021,N_1059);
and U1122 (N_1122,N_1058,N_1066);
and U1123 (N_1123,N_1023,N_1021);
xor U1124 (N_1124,N_1067,N_1077);
or U1125 (N_1125,N_1044,N_1056);
and U1126 (N_1126,N_1073,N_1040);
or U1127 (N_1127,N_1023,N_1039);
and U1128 (N_1128,N_1021,N_1076);
and U1129 (N_1129,N_1065,N_1036);
nand U1130 (N_1130,N_1070,N_1077);
nor U1131 (N_1131,N_1035,N_1055);
nor U1132 (N_1132,N_1059,N_1071);
nand U1133 (N_1133,N_1074,N_1025);
and U1134 (N_1134,N_1056,N_1077);
nor U1135 (N_1135,N_1074,N_1046);
nand U1136 (N_1136,N_1075,N_1022);
and U1137 (N_1137,N_1042,N_1021);
nand U1138 (N_1138,N_1062,N_1048);
nand U1139 (N_1139,N_1050,N_1076);
nand U1140 (N_1140,N_1084,N_1105);
nor U1141 (N_1141,N_1129,N_1119);
and U1142 (N_1142,N_1083,N_1098);
or U1143 (N_1143,N_1082,N_1101);
and U1144 (N_1144,N_1108,N_1127);
xnor U1145 (N_1145,N_1094,N_1121);
or U1146 (N_1146,N_1136,N_1092);
nor U1147 (N_1147,N_1106,N_1102);
nand U1148 (N_1148,N_1088,N_1131);
and U1149 (N_1149,N_1089,N_1124);
nand U1150 (N_1150,N_1095,N_1103);
or U1151 (N_1151,N_1138,N_1097);
nand U1152 (N_1152,N_1090,N_1117);
nand U1153 (N_1153,N_1116,N_1126);
and U1154 (N_1154,N_1107,N_1133);
and U1155 (N_1155,N_1115,N_1122);
and U1156 (N_1156,N_1111,N_1118);
nor U1157 (N_1157,N_1128,N_1104);
nor U1158 (N_1158,N_1125,N_1114);
and U1159 (N_1159,N_1081,N_1120);
nand U1160 (N_1160,N_1135,N_1113);
and U1161 (N_1161,N_1080,N_1123);
and U1162 (N_1162,N_1110,N_1109);
nor U1163 (N_1163,N_1096,N_1137);
nand U1164 (N_1164,N_1085,N_1130);
or U1165 (N_1165,N_1132,N_1093);
nor U1166 (N_1166,N_1087,N_1086);
and U1167 (N_1167,N_1112,N_1099);
nand U1168 (N_1168,N_1091,N_1139);
and U1169 (N_1169,N_1100,N_1134);
nor U1170 (N_1170,N_1121,N_1135);
or U1171 (N_1171,N_1112,N_1094);
and U1172 (N_1172,N_1134,N_1099);
or U1173 (N_1173,N_1121,N_1098);
or U1174 (N_1174,N_1134,N_1087);
and U1175 (N_1175,N_1125,N_1139);
nor U1176 (N_1176,N_1132,N_1111);
nand U1177 (N_1177,N_1135,N_1088);
and U1178 (N_1178,N_1138,N_1089);
and U1179 (N_1179,N_1139,N_1106);
or U1180 (N_1180,N_1090,N_1137);
nor U1181 (N_1181,N_1112,N_1089);
and U1182 (N_1182,N_1139,N_1082);
nor U1183 (N_1183,N_1121,N_1131);
or U1184 (N_1184,N_1134,N_1131);
or U1185 (N_1185,N_1135,N_1093);
or U1186 (N_1186,N_1117,N_1104);
nor U1187 (N_1187,N_1110,N_1082);
and U1188 (N_1188,N_1109,N_1084);
nand U1189 (N_1189,N_1139,N_1114);
and U1190 (N_1190,N_1118,N_1085);
nor U1191 (N_1191,N_1089,N_1100);
nand U1192 (N_1192,N_1139,N_1108);
and U1193 (N_1193,N_1130,N_1083);
nand U1194 (N_1194,N_1097,N_1121);
nand U1195 (N_1195,N_1107,N_1128);
or U1196 (N_1196,N_1118,N_1112);
and U1197 (N_1197,N_1112,N_1082);
or U1198 (N_1198,N_1131,N_1083);
or U1199 (N_1199,N_1134,N_1107);
and U1200 (N_1200,N_1157,N_1198);
and U1201 (N_1201,N_1145,N_1181);
nor U1202 (N_1202,N_1169,N_1144);
and U1203 (N_1203,N_1195,N_1140);
and U1204 (N_1204,N_1185,N_1192);
nor U1205 (N_1205,N_1196,N_1166);
and U1206 (N_1206,N_1155,N_1175);
nand U1207 (N_1207,N_1183,N_1153);
and U1208 (N_1208,N_1173,N_1199);
nand U1209 (N_1209,N_1171,N_1158);
nor U1210 (N_1210,N_1165,N_1172);
nor U1211 (N_1211,N_1148,N_1186);
nor U1212 (N_1212,N_1193,N_1149);
nor U1213 (N_1213,N_1174,N_1161);
and U1214 (N_1214,N_1177,N_1191);
and U1215 (N_1215,N_1182,N_1159);
nand U1216 (N_1216,N_1146,N_1163);
nor U1217 (N_1217,N_1184,N_1187);
or U1218 (N_1218,N_1190,N_1164);
and U1219 (N_1219,N_1189,N_1150);
or U1220 (N_1220,N_1179,N_1167);
and U1221 (N_1221,N_1154,N_1194);
nand U1222 (N_1222,N_1147,N_1162);
xor U1223 (N_1223,N_1188,N_1156);
and U1224 (N_1224,N_1170,N_1197);
nor U1225 (N_1225,N_1178,N_1160);
and U1226 (N_1226,N_1143,N_1141);
and U1227 (N_1227,N_1176,N_1151);
nor U1228 (N_1228,N_1142,N_1152);
or U1229 (N_1229,N_1180,N_1168);
nor U1230 (N_1230,N_1175,N_1196);
nor U1231 (N_1231,N_1148,N_1155);
xnor U1232 (N_1232,N_1196,N_1149);
nand U1233 (N_1233,N_1170,N_1154);
nand U1234 (N_1234,N_1167,N_1173);
or U1235 (N_1235,N_1187,N_1196);
or U1236 (N_1236,N_1172,N_1149);
nor U1237 (N_1237,N_1183,N_1161);
or U1238 (N_1238,N_1187,N_1172);
nand U1239 (N_1239,N_1174,N_1178);
nor U1240 (N_1240,N_1153,N_1149);
nand U1241 (N_1241,N_1140,N_1177);
nand U1242 (N_1242,N_1179,N_1176);
nand U1243 (N_1243,N_1159,N_1152);
and U1244 (N_1244,N_1146,N_1183);
nand U1245 (N_1245,N_1144,N_1142);
and U1246 (N_1246,N_1178,N_1168);
xnor U1247 (N_1247,N_1182,N_1199);
or U1248 (N_1248,N_1185,N_1169);
nand U1249 (N_1249,N_1186,N_1182);
nor U1250 (N_1250,N_1142,N_1181);
or U1251 (N_1251,N_1186,N_1192);
xnor U1252 (N_1252,N_1168,N_1150);
nor U1253 (N_1253,N_1158,N_1168);
or U1254 (N_1254,N_1183,N_1171);
nand U1255 (N_1255,N_1192,N_1158);
and U1256 (N_1256,N_1163,N_1188);
nor U1257 (N_1257,N_1144,N_1171);
nand U1258 (N_1258,N_1190,N_1199);
nor U1259 (N_1259,N_1147,N_1175);
nand U1260 (N_1260,N_1230,N_1247);
or U1261 (N_1261,N_1212,N_1234);
or U1262 (N_1262,N_1209,N_1224);
nand U1263 (N_1263,N_1238,N_1236);
or U1264 (N_1264,N_1228,N_1258);
or U1265 (N_1265,N_1237,N_1256);
nor U1266 (N_1266,N_1244,N_1242);
or U1267 (N_1267,N_1253,N_1232);
nor U1268 (N_1268,N_1235,N_1208);
or U1269 (N_1269,N_1204,N_1206);
xor U1270 (N_1270,N_1211,N_1240);
nand U1271 (N_1271,N_1223,N_1220);
nand U1272 (N_1272,N_1233,N_1210);
and U1273 (N_1273,N_1255,N_1217);
nand U1274 (N_1274,N_1215,N_1201);
or U1275 (N_1275,N_1246,N_1216);
nand U1276 (N_1276,N_1218,N_1254);
nand U1277 (N_1277,N_1239,N_1243);
or U1278 (N_1278,N_1259,N_1214);
nand U1279 (N_1279,N_1231,N_1221);
or U1280 (N_1280,N_1203,N_1241);
or U1281 (N_1281,N_1245,N_1227);
and U1282 (N_1282,N_1200,N_1251);
nor U1283 (N_1283,N_1226,N_1229);
nand U1284 (N_1284,N_1250,N_1225);
nand U1285 (N_1285,N_1249,N_1213);
and U1286 (N_1286,N_1205,N_1202);
and U1287 (N_1287,N_1222,N_1252);
nand U1288 (N_1288,N_1207,N_1257);
and U1289 (N_1289,N_1219,N_1248);
and U1290 (N_1290,N_1240,N_1216);
nor U1291 (N_1291,N_1212,N_1250);
nor U1292 (N_1292,N_1207,N_1206);
or U1293 (N_1293,N_1232,N_1219);
or U1294 (N_1294,N_1203,N_1251);
or U1295 (N_1295,N_1238,N_1232);
nand U1296 (N_1296,N_1207,N_1231);
or U1297 (N_1297,N_1203,N_1205);
nand U1298 (N_1298,N_1250,N_1259);
and U1299 (N_1299,N_1247,N_1221);
or U1300 (N_1300,N_1230,N_1256);
and U1301 (N_1301,N_1202,N_1233);
nor U1302 (N_1302,N_1244,N_1253);
or U1303 (N_1303,N_1217,N_1223);
nand U1304 (N_1304,N_1221,N_1224);
or U1305 (N_1305,N_1210,N_1238);
and U1306 (N_1306,N_1233,N_1255);
and U1307 (N_1307,N_1254,N_1216);
nor U1308 (N_1308,N_1224,N_1210);
or U1309 (N_1309,N_1246,N_1221);
nand U1310 (N_1310,N_1234,N_1251);
or U1311 (N_1311,N_1259,N_1244);
or U1312 (N_1312,N_1210,N_1254);
or U1313 (N_1313,N_1249,N_1202);
xor U1314 (N_1314,N_1241,N_1244);
nand U1315 (N_1315,N_1259,N_1216);
or U1316 (N_1316,N_1244,N_1226);
or U1317 (N_1317,N_1211,N_1247);
nand U1318 (N_1318,N_1235,N_1257);
nor U1319 (N_1319,N_1224,N_1254);
nor U1320 (N_1320,N_1294,N_1260);
nand U1321 (N_1321,N_1276,N_1283);
or U1322 (N_1322,N_1304,N_1299);
nor U1323 (N_1323,N_1297,N_1293);
or U1324 (N_1324,N_1266,N_1279);
nand U1325 (N_1325,N_1308,N_1309);
nand U1326 (N_1326,N_1314,N_1288);
nor U1327 (N_1327,N_1271,N_1312);
or U1328 (N_1328,N_1267,N_1280);
nand U1329 (N_1329,N_1269,N_1278);
nor U1330 (N_1330,N_1319,N_1291);
nand U1331 (N_1331,N_1302,N_1277);
nand U1332 (N_1332,N_1300,N_1295);
nand U1333 (N_1333,N_1262,N_1261);
nor U1334 (N_1334,N_1284,N_1282);
nor U1335 (N_1335,N_1303,N_1316);
nand U1336 (N_1336,N_1287,N_1305);
and U1337 (N_1337,N_1296,N_1285);
nor U1338 (N_1338,N_1264,N_1290);
or U1339 (N_1339,N_1286,N_1263);
nor U1340 (N_1340,N_1317,N_1268);
or U1341 (N_1341,N_1275,N_1270);
nand U1342 (N_1342,N_1289,N_1281);
nand U1343 (N_1343,N_1306,N_1301);
nor U1344 (N_1344,N_1265,N_1311);
nor U1345 (N_1345,N_1272,N_1298);
nand U1346 (N_1346,N_1273,N_1310);
nand U1347 (N_1347,N_1307,N_1318);
and U1348 (N_1348,N_1315,N_1274);
nor U1349 (N_1349,N_1292,N_1313);
and U1350 (N_1350,N_1263,N_1308);
nand U1351 (N_1351,N_1285,N_1262);
nand U1352 (N_1352,N_1285,N_1313);
and U1353 (N_1353,N_1294,N_1297);
or U1354 (N_1354,N_1260,N_1283);
nor U1355 (N_1355,N_1274,N_1275);
nor U1356 (N_1356,N_1274,N_1271);
and U1357 (N_1357,N_1303,N_1279);
and U1358 (N_1358,N_1281,N_1297);
nand U1359 (N_1359,N_1316,N_1269);
and U1360 (N_1360,N_1315,N_1273);
nand U1361 (N_1361,N_1280,N_1299);
or U1362 (N_1362,N_1273,N_1292);
and U1363 (N_1363,N_1288,N_1290);
nand U1364 (N_1364,N_1319,N_1264);
and U1365 (N_1365,N_1275,N_1280);
nor U1366 (N_1366,N_1300,N_1268);
nand U1367 (N_1367,N_1262,N_1274);
nor U1368 (N_1368,N_1298,N_1310);
nand U1369 (N_1369,N_1314,N_1296);
or U1370 (N_1370,N_1260,N_1267);
or U1371 (N_1371,N_1282,N_1290);
nor U1372 (N_1372,N_1274,N_1284);
or U1373 (N_1373,N_1269,N_1318);
and U1374 (N_1374,N_1264,N_1310);
nor U1375 (N_1375,N_1319,N_1260);
nand U1376 (N_1376,N_1290,N_1301);
and U1377 (N_1377,N_1277,N_1309);
or U1378 (N_1378,N_1266,N_1272);
nor U1379 (N_1379,N_1304,N_1315);
xor U1380 (N_1380,N_1346,N_1364);
and U1381 (N_1381,N_1340,N_1371);
nand U1382 (N_1382,N_1368,N_1344);
nand U1383 (N_1383,N_1320,N_1373);
and U1384 (N_1384,N_1327,N_1338);
or U1385 (N_1385,N_1335,N_1332);
xor U1386 (N_1386,N_1343,N_1326);
nor U1387 (N_1387,N_1339,N_1356);
nor U1388 (N_1388,N_1369,N_1362);
or U1389 (N_1389,N_1352,N_1342);
nor U1390 (N_1390,N_1328,N_1361);
or U1391 (N_1391,N_1370,N_1376);
or U1392 (N_1392,N_1367,N_1354);
or U1393 (N_1393,N_1375,N_1324);
nor U1394 (N_1394,N_1347,N_1360);
nand U1395 (N_1395,N_1329,N_1357);
nand U1396 (N_1396,N_1379,N_1378);
nand U1397 (N_1397,N_1336,N_1374);
nor U1398 (N_1398,N_1333,N_1330);
or U1399 (N_1399,N_1358,N_1323);
nand U1400 (N_1400,N_1355,N_1365);
and U1401 (N_1401,N_1321,N_1363);
nor U1402 (N_1402,N_1322,N_1349);
nor U1403 (N_1403,N_1377,N_1353);
or U1404 (N_1404,N_1359,N_1334);
nand U1405 (N_1405,N_1351,N_1372);
nand U1406 (N_1406,N_1341,N_1366);
and U1407 (N_1407,N_1348,N_1337);
and U1408 (N_1408,N_1345,N_1331);
nand U1409 (N_1409,N_1325,N_1350);
or U1410 (N_1410,N_1367,N_1321);
nor U1411 (N_1411,N_1350,N_1345);
nor U1412 (N_1412,N_1354,N_1360);
or U1413 (N_1413,N_1353,N_1365);
xnor U1414 (N_1414,N_1351,N_1323);
nor U1415 (N_1415,N_1350,N_1354);
and U1416 (N_1416,N_1375,N_1330);
xor U1417 (N_1417,N_1352,N_1324);
xnor U1418 (N_1418,N_1376,N_1330);
nand U1419 (N_1419,N_1365,N_1372);
and U1420 (N_1420,N_1358,N_1326);
or U1421 (N_1421,N_1367,N_1353);
and U1422 (N_1422,N_1368,N_1334);
and U1423 (N_1423,N_1329,N_1335);
nand U1424 (N_1424,N_1364,N_1377);
and U1425 (N_1425,N_1324,N_1363);
or U1426 (N_1426,N_1364,N_1370);
or U1427 (N_1427,N_1336,N_1322);
nor U1428 (N_1428,N_1326,N_1376);
nor U1429 (N_1429,N_1353,N_1338);
nand U1430 (N_1430,N_1340,N_1367);
nor U1431 (N_1431,N_1334,N_1378);
xor U1432 (N_1432,N_1371,N_1331);
nor U1433 (N_1433,N_1365,N_1328);
nor U1434 (N_1434,N_1341,N_1330);
or U1435 (N_1435,N_1359,N_1338);
nor U1436 (N_1436,N_1375,N_1337);
or U1437 (N_1437,N_1338,N_1377);
or U1438 (N_1438,N_1345,N_1357);
nor U1439 (N_1439,N_1362,N_1346);
nand U1440 (N_1440,N_1416,N_1439);
or U1441 (N_1441,N_1406,N_1405);
nor U1442 (N_1442,N_1392,N_1437);
nor U1443 (N_1443,N_1393,N_1384);
nor U1444 (N_1444,N_1429,N_1434);
or U1445 (N_1445,N_1435,N_1421);
nand U1446 (N_1446,N_1423,N_1413);
nand U1447 (N_1447,N_1403,N_1390);
nand U1448 (N_1448,N_1411,N_1382);
or U1449 (N_1449,N_1415,N_1414);
nand U1450 (N_1450,N_1430,N_1419);
nand U1451 (N_1451,N_1387,N_1396);
nand U1452 (N_1452,N_1424,N_1412);
and U1453 (N_1453,N_1425,N_1409);
and U1454 (N_1454,N_1404,N_1431);
nand U1455 (N_1455,N_1398,N_1410);
nand U1456 (N_1456,N_1395,N_1394);
or U1457 (N_1457,N_1389,N_1426);
nand U1458 (N_1458,N_1422,N_1428);
nor U1459 (N_1459,N_1401,N_1432);
and U1460 (N_1460,N_1408,N_1400);
nand U1461 (N_1461,N_1407,N_1399);
nand U1462 (N_1462,N_1433,N_1417);
or U1463 (N_1463,N_1427,N_1388);
and U1464 (N_1464,N_1418,N_1380);
and U1465 (N_1465,N_1381,N_1385);
and U1466 (N_1466,N_1386,N_1383);
nand U1467 (N_1467,N_1391,N_1436);
or U1468 (N_1468,N_1420,N_1397);
and U1469 (N_1469,N_1438,N_1402);
nor U1470 (N_1470,N_1412,N_1384);
or U1471 (N_1471,N_1391,N_1426);
nand U1472 (N_1472,N_1413,N_1405);
and U1473 (N_1473,N_1386,N_1423);
or U1474 (N_1474,N_1419,N_1432);
and U1475 (N_1475,N_1419,N_1406);
nand U1476 (N_1476,N_1386,N_1400);
xor U1477 (N_1477,N_1386,N_1419);
and U1478 (N_1478,N_1423,N_1391);
nor U1479 (N_1479,N_1393,N_1415);
nand U1480 (N_1480,N_1424,N_1427);
and U1481 (N_1481,N_1389,N_1437);
or U1482 (N_1482,N_1393,N_1421);
and U1483 (N_1483,N_1429,N_1408);
nor U1484 (N_1484,N_1404,N_1387);
nor U1485 (N_1485,N_1400,N_1397);
nand U1486 (N_1486,N_1436,N_1413);
or U1487 (N_1487,N_1436,N_1399);
nor U1488 (N_1488,N_1420,N_1414);
and U1489 (N_1489,N_1426,N_1382);
or U1490 (N_1490,N_1394,N_1434);
and U1491 (N_1491,N_1406,N_1417);
nand U1492 (N_1492,N_1414,N_1437);
or U1493 (N_1493,N_1420,N_1381);
and U1494 (N_1494,N_1431,N_1427);
and U1495 (N_1495,N_1381,N_1399);
nor U1496 (N_1496,N_1433,N_1430);
nor U1497 (N_1497,N_1431,N_1430);
and U1498 (N_1498,N_1394,N_1436);
nor U1499 (N_1499,N_1421,N_1404);
nor U1500 (N_1500,N_1440,N_1486);
nor U1501 (N_1501,N_1468,N_1467);
nand U1502 (N_1502,N_1497,N_1474);
and U1503 (N_1503,N_1469,N_1480);
and U1504 (N_1504,N_1496,N_1491);
and U1505 (N_1505,N_1490,N_1457);
and U1506 (N_1506,N_1443,N_1450);
nand U1507 (N_1507,N_1451,N_1482);
or U1508 (N_1508,N_1473,N_1460);
and U1509 (N_1509,N_1495,N_1493);
and U1510 (N_1510,N_1472,N_1456);
nand U1511 (N_1511,N_1477,N_1475);
nand U1512 (N_1512,N_1498,N_1463);
nor U1513 (N_1513,N_1471,N_1481);
or U1514 (N_1514,N_1441,N_1470);
xor U1515 (N_1515,N_1449,N_1494);
and U1516 (N_1516,N_1487,N_1446);
or U1517 (N_1517,N_1478,N_1444);
nor U1518 (N_1518,N_1458,N_1485);
and U1519 (N_1519,N_1461,N_1465);
nor U1520 (N_1520,N_1452,N_1479);
or U1521 (N_1521,N_1492,N_1466);
nor U1522 (N_1522,N_1455,N_1484);
and U1523 (N_1523,N_1454,N_1447);
nand U1524 (N_1524,N_1445,N_1442);
nand U1525 (N_1525,N_1448,N_1453);
and U1526 (N_1526,N_1483,N_1462);
nand U1527 (N_1527,N_1499,N_1459);
or U1528 (N_1528,N_1464,N_1476);
nand U1529 (N_1529,N_1488,N_1489);
nor U1530 (N_1530,N_1456,N_1450);
or U1531 (N_1531,N_1498,N_1499);
or U1532 (N_1532,N_1497,N_1478);
nor U1533 (N_1533,N_1474,N_1460);
and U1534 (N_1534,N_1451,N_1492);
nor U1535 (N_1535,N_1485,N_1467);
xnor U1536 (N_1536,N_1469,N_1466);
nand U1537 (N_1537,N_1484,N_1448);
nand U1538 (N_1538,N_1456,N_1490);
and U1539 (N_1539,N_1499,N_1442);
and U1540 (N_1540,N_1482,N_1465);
and U1541 (N_1541,N_1457,N_1459);
nand U1542 (N_1542,N_1460,N_1499);
or U1543 (N_1543,N_1485,N_1495);
nand U1544 (N_1544,N_1475,N_1490);
or U1545 (N_1545,N_1485,N_1441);
xor U1546 (N_1546,N_1449,N_1443);
and U1547 (N_1547,N_1496,N_1450);
nor U1548 (N_1548,N_1472,N_1483);
nor U1549 (N_1549,N_1454,N_1461);
nor U1550 (N_1550,N_1499,N_1449);
or U1551 (N_1551,N_1485,N_1454);
and U1552 (N_1552,N_1473,N_1459);
nor U1553 (N_1553,N_1462,N_1469);
and U1554 (N_1554,N_1482,N_1469);
nor U1555 (N_1555,N_1483,N_1476);
and U1556 (N_1556,N_1489,N_1462);
or U1557 (N_1557,N_1498,N_1451);
nor U1558 (N_1558,N_1497,N_1487);
nand U1559 (N_1559,N_1491,N_1481);
and U1560 (N_1560,N_1505,N_1534);
or U1561 (N_1561,N_1541,N_1544);
and U1562 (N_1562,N_1506,N_1537);
and U1563 (N_1563,N_1514,N_1557);
or U1564 (N_1564,N_1554,N_1532);
and U1565 (N_1565,N_1529,N_1555);
and U1566 (N_1566,N_1510,N_1533);
and U1567 (N_1567,N_1504,N_1531);
nor U1568 (N_1568,N_1548,N_1549);
or U1569 (N_1569,N_1522,N_1509);
nand U1570 (N_1570,N_1530,N_1519);
and U1571 (N_1571,N_1525,N_1546);
nor U1572 (N_1572,N_1511,N_1520);
nor U1573 (N_1573,N_1551,N_1528);
nand U1574 (N_1574,N_1526,N_1515);
and U1575 (N_1575,N_1527,N_1545);
or U1576 (N_1576,N_1500,N_1535);
nor U1577 (N_1577,N_1513,N_1512);
or U1578 (N_1578,N_1547,N_1518);
nand U1579 (N_1579,N_1543,N_1550);
nor U1580 (N_1580,N_1521,N_1516);
nand U1581 (N_1581,N_1558,N_1507);
and U1582 (N_1582,N_1540,N_1538);
and U1583 (N_1583,N_1501,N_1556);
nor U1584 (N_1584,N_1552,N_1523);
nor U1585 (N_1585,N_1503,N_1553);
nor U1586 (N_1586,N_1542,N_1502);
nor U1587 (N_1587,N_1517,N_1524);
or U1588 (N_1588,N_1536,N_1508);
nor U1589 (N_1589,N_1539,N_1559);
nor U1590 (N_1590,N_1538,N_1530);
and U1591 (N_1591,N_1518,N_1542);
and U1592 (N_1592,N_1546,N_1555);
or U1593 (N_1593,N_1500,N_1510);
nand U1594 (N_1594,N_1546,N_1526);
nor U1595 (N_1595,N_1558,N_1543);
or U1596 (N_1596,N_1540,N_1533);
and U1597 (N_1597,N_1554,N_1505);
and U1598 (N_1598,N_1550,N_1526);
nor U1599 (N_1599,N_1546,N_1500);
nor U1600 (N_1600,N_1542,N_1514);
nor U1601 (N_1601,N_1555,N_1557);
nand U1602 (N_1602,N_1555,N_1523);
and U1603 (N_1603,N_1532,N_1528);
and U1604 (N_1604,N_1542,N_1529);
nor U1605 (N_1605,N_1530,N_1539);
or U1606 (N_1606,N_1508,N_1520);
nand U1607 (N_1607,N_1557,N_1528);
or U1608 (N_1608,N_1521,N_1517);
xor U1609 (N_1609,N_1512,N_1507);
and U1610 (N_1610,N_1524,N_1507);
nand U1611 (N_1611,N_1549,N_1519);
or U1612 (N_1612,N_1544,N_1505);
and U1613 (N_1613,N_1535,N_1518);
nor U1614 (N_1614,N_1515,N_1529);
xnor U1615 (N_1615,N_1539,N_1545);
nor U1616 (N_1616,N_1502,N_1532);
and U1617 (N_1617,N_1534,N_1556);
or U1618 (N_1618,N_1511,N_1519);
or U1619 (N_1619,N_1505,N_1558);
nor U1620 (N_1620,N_1605,N_1611);
or U1621 (N_1621,N_1616,N_1609);
xnor U1622 (N_1622,N_1573,N_1574);
nand U1623 (N_1623,N_1590,N_1572);
and U1624 (N_1624,N_1589,N_1601);
nor U1625 (N_1625,N_1608,N_1586);
nand U1626 (N_1626,N_1618,N_1607);
nor U1627 (N_1627,N_1575,N_1580);
nor U1628 (N_1628,N_1619,N_1612);
and U1629 (N_1629,N_1614,N_1568);
nand U1630 (N_1630,N_1585,N_1561);
nand U1631 (N_1631,N_1613,N_1563);
or U1632 (N_1632,N_1600,N_1591);
nand U1633 (N_1633,N_1604,N_1615);
nand U1634 (N_1634,N_1598,N_1577);
nor U1635 (N_1635,N_1579,N_1584);
or U1636 (N_1636,N_1578,N_1567);
xor U1637 (N_1637,N_1581,N_1571);
and U1638 (N_1638,N_1583,N_1603);
nand U1639 (N_1639,N_1592,N_1565);
or U1640 (N_1640,N_1564,N_1593);
or U1641 (N_1641,N_1599,N_1588);
or U1642 (N_1642,N_1562,N_1569);
and U1643 (N_1643,N_1595,N_1610);
or U1644 (N_1644,N_1566,N_1602);
or U1645 (N_1645,N_1617,N_1596);
and U1646 (N_1646,N_1560,N_1597);
or U1647 (N_1647,N_1582,N_1587);
nand U1648 (N_1648,N_1594,N_1606);
and U1649 (N_1649,N_1570,N_1576);
and U1650 (N_1650,N_1566,N_1617);
and U1651 (N_1651,N_1595,N_1593);
nand U1652 (N_1652,N_1610,N_1580);
nor U1653 (N_1653,N_1569,N_1615);
nand U1654 (N_1654,N_1583,N_1604);
or U1655 (N_1655,N_1615,N_1584);
and U1656 (N_1656,N_1566,N_1613);
and U1657 (N_1657,N_1561,N_1560);
and U1658 (N_1658,N_1592,N_1561);
nand U1659 (N_1659,N_1569,N_1589);
or U1660 (N_1660,N_1579,N_1574);
nand U1661 (N_1661,N_1604,N_1575);
nor U1662 (N_1662,N_1564,N_1599);
nand U1663 (N_1663,N_1616,N_1567);
and U1664 (N_1664,N_1579,N_1560);
and U1665 (N_1665,N_1594,N_1598);
nor U1666 (N_1666,N_1569,N_1598);
xor U1667 (N_1667,N_1583,N_1572);
nor U1668 (N_1668,N_1597,N_1605);
nand U1669 (N_1669,N_1579,N_1615);
nand U1670 (N_1670,N_1613,N_1598);
or U1671 (N_1671,N_1580,N_1607);
or U1672 (N_1672,N_1563,N_1596);
and U1673 (N_1673,N_1592,N_1599);
nand U1674 (N_1674,N_1600,N_1590);
nand U1675 (N_1675,N_1617,N_1609);
xor U1676 (N_1676,N_1587,N_1613);
or U1677 (N_1677,N_1593,N_1606);
nor U1678 (N_1678,N_1608,N_1592);
and U1679 (N_1679,N_1574,N_1591);
nand U1680 (N_1680,N_1626,N_1647);
xnor U1681 (N_1681,N_1622,N_1631);
nor U1682 (N_1682,N_1666,N_1653);
nor U1683 (N_1683,N_1620,N_1674);
nand U1684 (N_1684,N_1663,N_1632);
or U1685 (N_1685,N_1627,N_1667);
xnor U1686 (N_1686,N_1633,N_1655);
nor U1687 (N_1687,N_1669,N_1658);
or U1688 (N_1688,N_1678,N_1664);
nand U1689 (N_1689,N_1679,N_1646);
nand U1690 (N_1690,N_1652,N_1637);
or U1691 (N_1691,N_1665,N_1636);
nor U1692 (N_1692,N_1677,N_1645);
nor U1693 (N_1693,N_1638,N_1648);
nor U1694 (N_1694,N_1650,N_1657);
xor U1695 (N_1695,N_1651,N_1630);
nor U1696 (N_1696,N_1640,N_1670);
nor U1697 (N_1697,N_1641,N_1649);
nand U1698 (N_1698,N_1675,N_1671);
or U1699 (N_1699,N_1642,N_1628);
and U1700 (N_1700,N_1629,N_1621);
nor U1701 (N_1701,N_1676,N_1662);
xor U1702 (N_1702,N_1668,N_1644);
and U1703 (N_1703,N_1659,N_1635);
and U1704 (N_1704,N_1624,N_1625);
and U1705 (N_1705,N_1639,N_1661);
nand U1706 (N_1706,N_1660,N_1623);
nor U1707 (N_1707,N_1656,N_1643);
or U1708 (N_1708,N_1654,N_1634);
or U1709 (N_1709,N_1673,N_1672);
nand U1710 (N_1710,N_1655,N_1649);
nor U1711 (N_1711,N_1670,N_1649);
and U1712 (N_1712,N_1626,N_1648);
nor U1713 (N_1713,N_1627,N_1666);
nand U1714 (N_1714,N_1627,N_1677);
nor U1715 (N_1715,N_1634,N_1679);
nor U1716 (N_1716,N_1670,N_1671);
or U1717 (N_1717,N_1624,N_1627);
and U1718 (N_1718,N_1674,N_1647);
nor U1719 (N_1719,N_1624,N_1677);
nand U1720 (N_1720,N_1639,N_1679);
and U1721 (N_1721,N_1649,N_1678);
nand U1722 (N_1722,N_1637,N_1639);
nand U1723 (N_1723,N_1625,N_1622);
or U1724 (N_1724,N_1635,N_1624);
and U1725 (N_1725,N_1662,N_1644);
or U1726 (N_1726,N_1620,N_1623);
or U1727 (N_1727,N_1650,N_1664);
nor U1728 (N_1728,N_1639,N_1627);
or U1729 (N_1729,N_1629,N_1623);
nor U1730 (N_1730,N_1661,N_1677);
nand U1731 (N_1731,N_1668,N_1651);
nand U1732 (N_1732,N_1675,N_1643);
nand U1733 (N_1733,N_1654,N_1678);
or U1734 (N_1734,N_1657,N_1629);
and U1735 (N_1735,N_1660,N_1627);
and U1736 (N_1736,N_1622,N_1654);
and U1737 (N_1737,N_1646,N_1620);
nand U1738 (N_1738,N_1640,N_1626);
and U1739 (N_1739,N_1638,N_1633);
nand U1740 (N_1740,N_1737,N_1694);
nor U1741 (N_1741,N_1693,N_1689);
nor U1742 (N_1742,N_1736,N_1707);
and U1743 (N_1743,N_1704,N_1721);
and U1744 (N_1744,N_1712,N_1702);
and U1745 (N_1745,N_1723,N_1732);
nand U1746 (N_1746,N_1728,N_1680);
nor U1747 (N_1747,N_1734,N_1700);
or U1748 (N_1748,N_1726,N_1703);
or U1749 (N_1749,N_1738,N_1716);
nand U1750 (N_1750,N_1681,N_1720);
nor U1751 (N_1751,N_1735,N_1698);
xor U1752 (N_1752,N_1691,N_1722);
nor U1753 (N_1753,N_1709,N_1724);
nor U1754 (N_1754,N_1696,N_1690);
or U1755 (N_1755,N_1739,N_1733);
and U1756 (N_1756,N_1687,N_1729);
xnor U1757 (N_1757,N_1711,N_1708);
nor U1758 (N_1758,N_1683,N_1717);
nand U1759 (N_1759,N_1697,N_1706);
nand U1760 (N_1760,N_1695,N_1686);
nor U1761 (N_1761,N_1715,N_1719);
nand U1762 (N_1762,N_1705,N_1727);
or U1763 (N_1763,N_1730,N_1701);
xor U1764 (N_1764,N_1725,N_1684);
nand U1765 (N_1765,N_1682,N_1713);
and U1766 (N_1766,N_1710,N_1699);
and U1767 (N_1767,N_1692,N_1685);
nor U1768 (N_1768,N_1718,N_1688);
or U1769 (N_1769,N_1731,N_1714);
nor U1770 (N_1770,N_1694,N_1723);
nor U1771 (N_1771,N_1684,N_1739);
and U1772 (N_1772,N_1730,N_1738);
and U1773 (N_1773,N_1682,N_1724);
nand U1774 (N_1774,N_1732,N_1718);
nor U1775 (N_1775,N_1721,N_1725);
nand U1776 (N_1776,N_1731,N_1686);
nor U1777 (N_1777,N_1708,N_1690);
and U1778 (N_1778,N_1687,N_1691);
nand U1779 (N_1779,N_1737,N_1717);
or U1780 (N_1780,N_1682,N_1707);
nor U1781 (N_1781,N_1714,N_1736);
or U1782 (N_1782,N_1731,N_1737);
nor U1783 (N_1783,N_1704,N_1685);
nor U1784 (N_1784,N_1691,N_1724);
nand U1785 (N_1785,N_1721,N_1730);
nor U1786 (N_1786,N_1724,N_1730);
and U1787 (N_1787,N_1697,N_1738);
xor U1788 (N_1788,N_1699,N_1723);
nand U1789 (N_1789,N_1739,N_1730);
nor U1790 (N_1790,N_1722,N_1708);
nor U1791 (N_1791,N_1724,N_1703);
or U1792 (N_1792,N_1727,N_1708);
and U1793 (N_1793,N_1727,N_1728);
nor U1794 (N_1794,N_1736,N_1728);
xnor U1795 (N_1795,N_1694,N_1681);
and U1796 (N_1796,N_1723,N_1700);
or U1797 (N_1797,N_1689,N_1702);
or U1798 (N_1798,N_1714,N_1710);
nor U1799 (N_1799,N_1705,N_1711);
or U1800 (N_1800,N_1741,N_1764);
or U1801 (N_1801,N_1773,N_1766);
or U1802 (N_1802,N_1789,N_1750);
nor U1803 (N_1803,N_1794,N_1748);
nor U1804 (N_1804,N_1784,N_1795);
nor U1805 (N_1805,N_1769,N_1746);
nor U1806 (N_1806,N_1787,N_1755);
nand U1807 (N_1807,N_1783,N_1763);
nor U1808 (N_1808,N_1771,N_1786);
and U1809 (N_1809,N_1779,N_1774);
nor U1810 (N_1810,N_1759,N_1745);
or U1811 (N_1811,N_1767,N_1792);
nand U1812 (N_1812,N_1761,N_1747);
and U1813 (N_1813,N_1754,N_1778);
and U1814 (N_1814,N_1799,N_1790);
nand U1815 (N_1815,N_1756,N_1777);
nand U1816 (N_1816,N_1775,N_1791);
or U1817 (N_1817,N_1758,N_1742);
and U1818 (N_1818,N_1753,N_1743);
nor U1819 (N_1819,N_1797,N_1744);
nand U1820 (N_1820,N_1793,N_1760);
and U1821 (N_1821,N_1752,N_1782);
or U1822 (N_1822,N_1788,N_1772);
nor U1823 (N_1823,N_1757,N_1785);
nand U1824 (N_1824,N_1765,N_1751);
nand U1825 (N_1825,N_1768,N_1762);
and U1826 (N_1826,N_1780,N_1796);
or U1827 (N_1827,N_1740,N_1770);
and U1828 (N_1828,N_1798,N_1749);
and U1829 (N_1829,N_1781,N_1776);
nor U1830 (N_1830,N_1747,N_1756);
and U1831 (N_1831,N_1793,N_1744);
nor U1832 (N_1832,N_1799,N_1791);
nor U1833 (N_1833,N_1754,N_1755);
nor U1834 (N_1834,N_1774,N_1790);
and U1835 (N_1835,N_1787,N_1743);
nor U1836 (N_1836,N_1782,N_1762);
and U1837 (N_1837,N_1784,N_1785);
and U1838 (N_1838,N_1791,N_1757);
and U1839 (N_1839,N_1796,N_1792);
nor U1840 (N_1840,N_1766,N_1782);
xor U1841 (N_1841,N_1793,N_1750);
and U1842 (N_1842,N_1747,N_1762);
nand U1843 (N_1843,N_1792,N_1787);
nand U1844 (N_1844,N_1754,N_1749);
and U1845 (N_1845,N_1741,N_1754);
and U1846 (N_1846,N_1783,N_1779);
nor U1847 (N_1847,N_1742,N_1765);
nor U1848 (N_1848,N_1794,N_1786);
or U1849 (N_1849,N_1782,N_1757);
nand U1850 (N_1850,N_1770,N_1767);
nand U1851 (N_1851,N_1768,N_1752);
nand U1852 (N_1852,N_1740,N_1786);
nor U1853 (N_1853,N_1763,N_1742);
nand U1854 (N_1854,N_1746,N_1779);
or U1855 (N_1855,N_1766,N_1799);
or U1856 (N_1856,N_1777,N_1782);
and U1857 (N_1857,N_1771,N_1778);
nor U1858 (N_1858,N_1776,N_1769);
or U1859 (N_1859,N_1797,N_1767);
nand U1860 (N_1860,N_1848,N_1832);
or U1861 (N_1861,N_1858,N_1838);
xor U1862 (N_1862,N_1845,N_1840);
nand U1863 (N_1863,N_1849,N_1821);
nand U1864 (N_1864,N_1830,N_1829);
nand U1865 (N_1865,N_1819,N_1833);
nand U1866 (N_1866,N_1818,N_1844);
nor U1867 (N_1867,N_1811,N_1857);
nor U1868 (N_1868,N_1828,N_1846);
nor U1869 (N_1869,N_1809,N_1808);
or U1870 (N_1870,N_1847,N_1859);
nand U1871 (N_1871,N_1803,N_1851);
and U1872 (N_1872,N_1841,N_1802);
and U1873 (N_1873,N_1805,N_1813);
and U1874 (N_1874,N_1824,N_1827);
nor U1875 (N_1875,N_1816,N_1839);
or U1876 (N_1876,N_1855,N_1825);
or U1877 (N_1877,N_1856,N_1800);
or U1878 (N_1878,N_1814,N_1804);
nand U1879 (N_1879,N_1843,N_1817);
nand U1880 (N_1880,N_1853,N_1852);
and U1881 (N_1881,N_1837,N_1834);
or U1882 (N_1882,N_1823,N_1801);
or U1883 (N_1883,N_1850,N_1854);
nand U1884 (N_1884,N_1810,N_1807);
and U1885 (N_1885,N_1822,N_1826);
nand U1886 (N_1886,N_1815,N_1842);
nor U1887 (N_1887,N_1835,N_1836);
nor U1888 (N_1888,N_1831,N_1812);
nand U1889 (N_1889,N_1820,N_1806);
nor U1890 (N_1890,N_1833,N_1815);
nand U1891 (N_1891,N_1823,N_1856);
nand U1892 (N_1892,N_1848,N_1829);
and U1893 (N_1893,N_1837,N_1803);
or U1894 (N_1894,N_1815,N_1811);
and U1895 (N_1895,N_1838,N_1835);
nand U1896 (N_1896,N_1820,N_1818);
nand U1897 (N_1897,N_1820,N_1836);
and U1898 (N_1898,N_1811,N_1825);
or U1899 (N_1899,N_1833,N_1807);
or U1900 (N_1900,N_1817,N_1812);
or U1901 (N_1901,N_1828,N_1808);
nor U1902 (N_1902,N_1809,N_1801);
nor U1903 (N_1903,N_1852,N_1822);
and U1904 (N_1904,N_1857,N_1808);
and U1905 (N_1905,N_1834,N_1833);
and U1906 (N_1906,N_1826,N_1824);
nand U1907 (N_1907,N_1838,N_1818);
nand U1908 (N_1908,N_1811,N_1851);
nor U1909 (N_1909,N_1838,N_1807);
and U1910 (N_1910,N_1818,N_1854);
or U1911 (N_1911,N_1811,N_1837);
or U1912 (N_1912,N_1836,N_1851);
or U1913 (N_1913,N_1826,N_1857);
or U1914 (N_1914,N_1842,N_1820);
nand U1915 (N_1915,N_1833,N_1806);
nor U1916 (N_1916,N_1844,N_1855);
or U1917 (N_1917,N_1830,N_1835);
and U1918 (N_1918,N_1820,N_1837);
nor U1919 (N_1919,N_1801,N_1837);
or U1920 (N_1920,N_1919,N_1871);
nor U1921 (N_1921,N_1894,N_1907);
nor U1922 (N_1922,N_1903,N_1904);
or U1923 (N_1923,N_1917,N_1918);
nand U1924 (N_1924,N_1909,N_1897);
nor U1925 (N_1925,N_1870,N_1895);
or U1926 (N_1926,N_1901,N_1911);
or U1927 (N_1927,N_1910,N_1892);
nand U1928 (N_1928,N_1868,N_1880);
or U1929 (N_1929,N_1874,N_1872);
nor U1930 (N_1930,N_1912,N_1867);
nand U1931 (N_1931,N_1864,N_1866);
or U1932 (N_1932,N_1915,N_1887);
and U1933 (N_1933,N_1889,N_1908);
nand U1934 (N_1934,N_1876,N_1865);
and U1935 (N_1935,N_1882,N_1869);
nor U1936 (N_1936,N_1888,N_1896);
nand U1937 (N_1937,N_1884,N_1899);
nor U1938 (N_1938,N_1905,N_1890);
nand U1939 (N_1939,N_1862,N_1877);
nor U1940 (N_1940,N_1875,N_1906);
nor U1941 (N_1941,N_1914,N_1873);
and U1942 (N_1942,N_1913,N_1878);
or U1943 (N_1943,N_1861,N_1900);
nor U1944 (N_1944,N_1860,N_1863);
or U1945 (N_1945,N_1885,N_1898);
nor U1946 (N_1946,N_1916,N_1879);
or U1947 (N_1947,N_1893,N_1891);
or U1948 (N_1948,N_1886,N_1883);
and U1949 (N_1949,N_1881,N_1902);
and U1950 (N_1950,N_1863,N_1907);
or U1951 (N_1951,N_1896,N_1905);
and U1952 (N_1952,N_1886,N_1871);
or U1953 (N_1953,N_1873,N_1918);
nand U1954 (N_1954,N_1867,N_1863);
or U1955 (N_1955,N_1870,N_1896);
nand U1956 (N_1956,N_1864,N_1897);
nand U1957 (N_1957,N_1911,N_1887);
or U1958 (N_1958,N_1870,N_1898);
nand U1959 (N_1959,N_1903,N_1916);
nor U1960 (N_1960,N_1891,N_1890);
and U1961 (N_1961,N_1902,N_1867);
and U1962 (N_1962,N_1884,N_1903);
and U1963 (N_1963,N_1876,N_1901);
nor U1964 (N_1964,N_1874,N_1892);
xnor U1965 (N_1965,N_1915,N_1869);
or U1966 (N_1966,N_1915,N_1889);
nand U1967 (N_1967,N_1881,N_1906);
nor U1968 (N_1968,N_1901,N_1879);
nand U1969 (N_1969,N_1878,N_1892);
and U1970 (N_1970,N_1913,N_1914);
nor U1971 (N_1971,N_1871,N_1881);
nor U1972 (N_1972,N_1890,N_1897);
and U1973 (N_1973,N_1903,N_1919);
and U1974 (N_1974,N_1909,N_1877);
nor U1975 (N_1975,N_1880,N_1893);
nor U1976 (N_1976,N_1881,N_1910);
and U1977 (N_1977,N_1900,N_1883);
nand U1978 (N_1978,N_1896,N_1898);
xnor U1979 (N_1979,N_1860,N_1886);
and U1980 (N_1980,N_1942,N_1920);
and U1981 (N_1981,N_1941,N_1958);
nor U1982 (N_1982,N_1949,N_1976);
and U1983 (N_1983,N_1924,N_1964);
and U1984 (N_1984,N_1951,N_1932);
nor U1985 (N_1985,N_1931,N_1947);
nand U1986 (N_1986,N_1938,N_1946);
nand U1987 (N_1987,N_1965,N_1954);
and U1988 (N_1988,N_1975,N_1927);
xnor U1989 (N_1989,N_1933,N_1945);
nand U1990 (N_1990,N_1961,N_1923);
or U1991 (N_1991,N_1926,N_1928);
or U1992 (N_1992,N_1972,N_1930);
and U1993 (N_1993,N_1935,N_1968);
nand U1994 (N_1994,N_1977,N_1921);
or U1995 (N_1995,N_1978,N_1971);
and U1996 (N_1996,N_1953,N_1963);
or U1997 (N_1997,N_1962,N_1929);
and U1998 (N_1998,N_1937,N_1936);
or U1999 (N_1999,N_1967,N_1974);
and U2000 (N_2000,N_1956,N_1957);
nor U2001 (N_2001,N_1960,N_1955);
or U2002 (N_2002,N_1948,N_1943);
nor U2003 (N_2003,N_1922,N_1925);
nand U2004 (N_2004,N_1939,N_1959);
and U2005 (N_2005,N_1950,N_1934);
nor U2006 (N_2006,N_1970,N_1969);
nand U2007 (N_2007,N_1940,N_1979);
nor U2008 (N_2008,N_1973,N_1966);
nand U2009 (N_2009,N_1944,N_1952);
nor U2010 (N_2010,N_1939,N_1941);
nand U2011 (N_2011,N_1942,N_1940);
nand U2012 (N_2012,N_1955,N_1944);
nor U2013 (N_2013,N_1945,N_1932);
or U2014 (N_2014,N_1962,N_1950);
or U2015 (N_2015,N_1940,N_1974);
nand U2016 (N_2016,N_1921,N_1924);
nand U2017 (N_2017,N_1949,N_1938);
and U2018 (N_2018,N_1949,N_1957);
nand U2019 (N_2019,N_1960,N_1965);
and U2020 (N_2020,N_1936,N_1948);
and U2021 (N_2021,N_1934,N_1925);
nand U2022 (N_2022,N_1922,N_1959);
nand U2023 (N_2023,N_1931,N_1943);
nand U2024 (N_2024,N_1955,N_1965);
nand U2025 (N_2025,N_1964,N_1963);
xor U2026 (N_2026,N_1956,N_1967);
nor U2027 (N_2027,N_1957,N_1924);
and U2028 (N_2028,N_1932,N_1971);
nor U2029 (N_2029,N_1975,N_1955);
and U2030 (N_2030,N_1971,N_1938);
and U2031 (N_2031,N_1964,N_1959);
nor U2032 (N_2032,N_1945,N_1928);
nand U2033 (N_2033,N_1922,N_1966);
and U2034 (N_2034,N_1955,N_1959);
nand U2035 (N_2035,N_1960,N_1930);
nand U2036 (N_2036,N_1964,N_1931);
nor U2037 (N_2037,N_1937,N_1928);
nor U2038 (N_2038,N_1970,N_1974);
nor U2039 (N_2039,N_1949,N_1974);
and U2040 (N_2040,N_2007,N_1987);
nand U2041 (N_2041,N_1994,N_1988);
and U2042 (N_2042,N_1999,N_2002);
nor U2043 (N_2043,N_1991,N_1980);
and U2044 (N_2044,N_2017,N_2038);
and U2045 (N_2045,N_2008,N_1986);
nor U2046 (N_2046,N_2022,N_2032);
and U2047 (N_2047,N_1993,N_2036);
or U2048 (N_2048,N_2029,N_2026);
and U2049 (N_2049,N_2000,N_2028);
and U2050 (N_2050,N_1985,N_2003);
or U2051 (N_2051,N_1992,N_2031);
nand U2052 (N_2052,N_2021,N_1998);
or U2053 (N_2053,N_1983,N_2011);
or U2054 (N_2054,N_2010,N_2019);
and U2055 (N_2055,N_2024,N_2037);
or U2056 (N_2056,N_2012,N_2023);
nand U2057 (N_2057,N_1984,N_2001);
nand U2058 (N_2058,N_2009,N_1989);
and U2059 (N_2059,N_2004,N_2027);
and U2060 (N_2060,N_2030,N_1995);
and U2061 (N_2061,N_1997,N_1996);
nor U2062 (N_2062,N_2013,N_2005);
or U2063 (N_2063,N_2020,N_2039);
nand U2064 (N_2064,N_1990,N_2033);
and U2065 (N_2065,N_1982,N_2006);
nand U2066 (N_2066,N_2016,N_2035);
nand U2067 (N_2067,N_2018,N_1981);
nor U2068 (N_2068,N_2034,N_2015);
nor U2069 (N_2069,N_2025,N_2014);
nor U2070 (N_2070,N_2008,N_2025);
and U2071 (N_2071,N_2021,N_2022);
or U2072 (N_2072,N_1986,N_2026);
nand U2073 (N_2073,N_2032,N_1987);
and U2074 (N_2074,N_2001,N_2006);
xor U2075 (N_2075,N_2012,N_2003);
nand U2076 (N_2076,N_2008,N_1991);
or U2077 (N_2077,N_2039,N_2016);
and U2078 (N_2078,N_2008,N_2034);
or U2079 (N_2079,N_2030,N_2001);
nand U2080 (N_2080,N_1999,N_1986);
and U2081 (N_2081,N_1983,N_1998);
nor U2082 (N_2082,N_1989,N_1988);
or U2083 (N_2083,N_2037,N_1996);
and U2084 (N_2084,N_2011,N_2008);
nand U2085 (N_2085,N_1980,N_1998);
and U2086 (N_2086,N_2032,N_2036);
nand U2087 (N_2087,N_2014,N_2028);
nor U2088 (N_2088,N_1997,N_1987);
nor U2089 (N_2089,N_1985,N_2032);
and U2090 (N_2090,N_2029,N_2023);
nor U2091 (N_2091,N_2020,N_2001);
and U2092 (N_2092,N_2002,N_1994);
nor U2093 (N_2093,N_2017,N_1995);
and U2094 (N_2094,N_2007,N_2001);
nand U2095 (N_2095,N_1998,N_2001);
nand U2096 (N_2096,N_1994,N_2001);
nand U2097 (N_2097,N_2030,N_2029);
or U2098 (N_2098,N_2015,N_2030);
and U2099 (N_2099,N_2002,N_2004);
nor U2100 (N_2100,N_2068,N_2073);
or U2101 (N_2101,N_2072,N_2097);
nand U2102 (N_2102,N_2053,N_2076);
nor U2103 (N_2103,N_2044,N_2094);
nor U2104 (N_2104,N_2087,N_2080);
and U2105 (N_2105,N_2054,N_2045);
and U2106 (N_2106,N_2099,N_2066);
nor U2107 (N_2107,N_2091,N_2047);
nand U2108 (N_2108,N_2051,N_2046);
or U2109 (N_2109,N_2075,N_2083);
nor U2110 (N_2110,N_2067,N_2042);
nor U2111 (N_2111,N_2040,N_2086);
and U2112 (N_2112,N_2059,N_2049);
nor U2113 (N_2113,N_2056,N_2043);
nor U2114 (N_2114,N_2078,N_2077);
nand U2115 (N_2115,N_2048,N_2060);
nand U2116 (N_2116,N_2095,N_2071);
nand U2117 (N_2117,N_2070,N_2063);
and U2118 (N_2118,N_2081,N_2085);
or U2119 (N_2119,N_2064,N_2061);
nand U2120 (N_2120,N_2058,N_2065);
nand U2121 (N_2121,N_2057,N_2041);
nand U2122 (N_2122,N_2069,N_2050);
and U2123 (N_2123,N_2092,N_2052);
nand U2124 (N_2124,N_2096,N_2082);
and U2125 (N_2125,N_2098,N_2089);
nand U2126 (N_2126,N_2090,N_2093);
xor U2127 (N_2127,N_2079,N_2084);
nor U2128 (N_2128,N_2088,N_2055);
and U2129 (N_2129,N_2062,N_2074);
nor U2130 (N_2130,N_2084,N_2056);
nor U2131 (N_2131,N_2098,N_2051);
nor U2132 (N_2132,N_2093,N_2053);
or U2133 (N_2133,N_2041,N_2083);
nor U2134 (N_2134,N_2041,N_2096);
or U2135 (N_2135,N_2084,N_2041);
or U2136 (N_2136,N_2094,N_2056);
or U2137 (N_2137,N_2068,N_2099);
and U2138 (N_2138,N_2048,N_2062);
and U2139 (N_2139,N_2049,N_2068);
nor U2140 (N_2140,N_2055,N_2093);
or U2141 (N_2141,N_2074,N_2075);
or U2142 (N_2142,N_2053,N_2073);
and U2143 (N_2143,N_2048,N_2082);
and U2144 (N_2144,N_2060,N_2099);
and U2145 (N_2145,N_2091,N_2064);
nor U2146 (N_2146,N_2052,N_2042);
nor U2147 (N_2147,N_2067,N_2061);
and U2148 (N_2148,N_2046,N_2057);
nor U2149 (N_2149,N_2072,N_2069);
nand U2150 (N_2150,N_2048,N_2099);
nand U2151 (N_2151,N_2055,N_2098);
and U2152 (N_2152,N_2046,N_2070);
xnor U2153 (N_2153,N_2068,N_2094);
nand U2154 (N_2154,N_2076,N_2045);
or U2155 (N_2155,N_2067,N_2085);
and U2156 (N_2156,N_2065,N_2066);
nand U2157 (N_2157,N_2082,N_2091);
or U2158 (N_2158,N_2073,N_2043);
nor U2159 (N_2159,N_2041,N_2042);
or U2160 (N_2160,N_2131,N_2156);
or U2161 (N_2161,N_2108,N_2130);
and U2162 (N_2162,N_2154,N_2122);
or U2163 (N_2163,N_2117,N_2152);
and U2164 (N_2164,N_2157,N_2121);
nor U2165 (N_2165,N_2127,N_2146);
or U2166 (N_2166,N_2119,N_2120);
nor U2167 (N_2167,N_2138,N_2159);
nor U2168 (N_2168,N_2115,N_2113);
nand U2169 (N_2169,N_2141,N_2142);
nor U2170 (N_2170,N_2129,N_2135);
nor U2171 (N_2171,N_2134,N_2144);
and U2172 (N_2172,N_2118,N_2128);
nor U2173 (N_2173,N_2147,N_2103);
nand U2174 (N_2174,N_2143,N_2132);
nor U2175 (N_2175,N_2104,N_2109);
or U2176 (N_2176,N_2139,N_2116);
nor U2177 (N_2177,N_2140,N_2136);
and U2178 (N_2178,N_2100,N_2101);
nand U2179 (N_2179,N_2137,N_2107);
xor U2180 (N_2180,N_2125,N_2105);
or U2181 (N_2181,N_2110,N_2112);
or U2182 (N_2182,N_2150,N_2126);
nor U2183 (N_2183,N_2114,N_2123);
and U2184 (N_2184,N_2153,N_2155);
and U2185 (N_2185,N_2102,N_2145);
nand U2186 (N_2186,N_2149,N_2106);
nand U2187 (N_2187,N_2124,N_2133);
and U2188 (N_2188,N_2151,N_2158);
nand U2189 (N_2189,N_2111,N_2148);
nand U2190 (N_2190,N_2137,N_2109);
nand U2191 (N_2191,N_2149,N_2135);
nand U2192 (N_2192,N_2157,N_2152);
nand U2193 (N_2193,N_2140,N_2104);
and U2194 (N_2194,N_2143,N_2103);
nand U2195 (N_2195,N_2129,N_2152);
nand U2196 (N_2196,N_2106,N_2118);
and U2197 (N_2197,N_2140,N_2130);
and U2198 (N_2198,N_2111,N_2157);
and U2199 (N_2199,N_2120,N_2107);
or U2200 (N_2200,N_2114,N_2106);
and U2201 (N_2201,N_2108,N_2131);
nor U2202 (N_2202,N_2146,N_2159);
or U2203 (N_2203,N_2153,N_2152);
nand U2204 (N_2204,N_2135,N_2132);
and U2205 (N_2205,N_2117,N_2114);
and U2206 (N_2206,N_2142,N_2113);
or U2207 (N_2207,N_2128,N_2136);
or U2208 (N_2208,N_2119,N_2159);
nand U2209 (N_2209,N_2141,N_2106);
and U2210 (N_2210,N_2105,N_2118);
nand U2211 (N_2211,N_2114,N_2122);
and U2212 (N_2212,N_2101,N_2117);
nor U2213 (N_2213,N_2149,N_2110);
and U2214 (N_2214,N_2142,N_2155);
nor U2215 (N_2215,N_2111,N_2156);
or U2216 (N_2216,N_2141,N_2107);
or U2217 (N_2217,N_2104,N_2152);
nor U2218 (N_2218,N_2140,N_2102);
or U2219 (N_2219,N_2108,N_2113);
nor U2220 (N_2220,N_2167,N_2181);
and U2221 (N_2221,N_2165,N_2201);
or U2222 (N_2222,N_2204,N_2196);
or U2223 (N_2223,N_2169,N_2215);
nor U2224 (N_2224,N_2166,N_2192);
or U2225 (N_2225,N_2199,N_2202);
nor U2226 (N_2226,N_2184,N_2174);
nand U2227 (N_2227,N_2172,N_2160);
or U2228 (N_2228,N_2193,N_2179);
or U2229 (N_2229,N_2212,N_2208);
and U2230 (N_2230,N_2188,N_2211);
or U2231 (N_2231,N_2190,N_2171);
nor U2232 (N_2232,N_2207,N_2189);
and U2233 (N_2233,N_2180,N_2163);
nor U2234 (N_2234,N_2219,N_2170);
or U2235 (N_2235,N_2173,N_2176);
nand U2236 (N_2236,N_2217,N_2210);
nand U2237 (N_2237,N_2191,N_2205);
nor U2238 (N_2238,N_2218,N_2203);
and U2239 (N_2239,N_2175,N_2162);
xnor U2240 (N_2240,N_2187,N_2195);
and U2241 (N_2241,N_2200,N_2206);
and U2242 (N_2242,N_2198,N_2164);
or U2243 (N_2243,N_2213,N_2186);
and U2244 (N_2244,N_2168,N_2194);
nand U2245 (N_2245,N_2177,N_2178);
or U2246 (N_2246,N_2197,N_2182);
or U2247 (N_2247,N_2183,N_2214);
or U2248 (N_2248,N_2161,N_2185);
nand U2249 (N_2249,N_2209,N_2216);
and U2250 (N_2250,N_2183,N_2164);
or U2251 (N_2251,N_2197,N_2212);
or U2252 (N_2252,N_2187,N_2216);
and U2253 (N_2253,N_2216,N_2179);
nor U2254 (N_2254,N_2165,N_2176);
or U2255 (N_2255,N_2198,N_2208);
and U2256 (N_2256,N_2192,N_2168);
or U2257 (N_2257,N_2200,N_2179);
nand U2258 (N_2258,N_2182,N_2215);
nor U2259 (N_2259,N_2196,N_2200);
nand U2260 (N_2260,N_2204,N_2160);
nor U2261 (N_2261,N_2219,N_2177);
nor U2262 (N_2262,N_2172,N_2167);
nor U2263 (N_2263,N_2214,N_2165);
nor U2264 (N_2264,N_2170,N_2207);
or U2265 (N_2265,N_2197,N_2185);
or U2266 (N_2266,N_2213,N_2182);
or U2267 (N_2267,N_2181,N_2169);
or U2268 (N_2268,N_2167,N_2186);
or U2269 (N_2269,N_2190,N_2184);
nor U2270 (N_2270,N_2162,N_2173);
or U2271 (N_2271,N_2176,N_2219);
or U2272 (N_2272,N_2187,N_2200);
xnor U2273 (N_2273,N_2193,N_2171);
or U2274 (N_2274,N_2180,N_2201);
nand U2275 (N_2275,N_2173,N_2181);
nand U2276 (N_2276,N_2205,N_2170);
nor U2277 (N_2277,N_2188,N_2197);
nand U2278 (N_2278,N_2166,N_2172);
nor U2279 (N_2279,N_2183,N_2219);
nor U2280 (N_2280,N_2225,N_2257);
or U2281 (N_2281,N_2251,N_2235);
or U2282 (N_2282,N_2278,N_2239);
and U2283 (N_2283,N_2245,N_2271);
nand U2284 (N_2284,N_2227,N_2261);
nand U2285 (N_2285,N_2269,N_2274);
nand U2286 (N_2286,N_2234,N_2268);
nand U2287 (N_2287,N_2242,N_2252);
or U2288 (N_2288,N_2260,N_2279);
and U2289 (N_2289,N_2246,N_2275);
nor U2290 (N_2290,N_2223,N_2256);
and U2291 (N_2291,N_2243,N_2267);
or U2292 (N_2292,N_2277,N_2233);
nor U2293 (N_2293,N_2241,N_2222);
nand U2294 (N_2294,N_2229,N_2236);
or U2295 (N_2295,N_2254,N_2228);
nor U2296 (N_2296,N_2240,N_2250);
and U2297 (N_2297,N_2244,N_2230);
nor U2298 (N_2298,N_2265,N_2237);
nor U2299 (N_2299,N_2263,N_2220);
nor U2300 (N_2300,N_2238,N_2273);
and U2301 (N_2301,N_2249,N_2258);
or U2302 (N_2302,N_2221,N_2226);
nand U2303 (N_2303,N_2270,N_2255);
nand U2304 (N_2304,N_2262,N_2247);
or U2305 (N_2305,N_2248,N_2232);
xor U2306 (N_2306,N_2224,N_2266);
or U2307 (N_2307,N_2264,N_2231);
or U2308 (N_2308,N_2253,N_2276);
and U2309 (N_2309,N_2272,N_2259);
nand U2310 (N_2310,N_2269,N_2237);
and U2311 (N_2311,N_2239,N_2248);
and U2312 (N_2312,N_2251,N_2237);
nor U2313 (N_2313,N_2234,N_2223);
nor U2314 (N_2314,N_2234,N_2240);
and U2315 (N_2315,N_2223,N_2252);
and U2316 (N_2316,N_2275,N_2255);
nand U2317 (N_2317,N_2267,N_2273);
and U2318 (N_2318,N_2231,N_2230);
or U2319 (N_2319,N_2229,N_2275);
xor U2320 (N_2320,N_2244,N_2242);
and U2321 (N_2321,N_2239,N_2222);
or U2322 (N_2322,N_2221,N_2223);
and U2323 (N_2323,N_2256,N_2232);
and U2324 (N_2324,N_2263,N_2271);
or U2325 (N_2325,N_2230,N_2275);
and U2326 (N_2326,N_2234,N_2274);
nor U2327 (N_2327,N_2252,N_2250);
or U2328 (N_2328,N_2260,N_2258);
nor U2329 (N_2329,N_2238,N_2227);
and U2330 (N_2330,N_2261,N_2232);
nand U2331 (N_2331,N_2225,N_2267);
nor U2332 (N_2332,N_2241,N_2258);
nor U2333 (N_2333,N_2234,N_2256);
nor U2334 (N_2334,N_2259,N_2274);
nand U2335 (N_2335,N_2229,N_2269);
or U2336 (N_2336,N_2223,N_2241);
and U2337 (N_2337,N_2258,N_2232);
nand U2338 (N_2338,N_2260,N_2250);
or U2339 (N_2339,N_2279,N_2262);
and U2340 (N_2340,N_2286,N_2322);
nand U2341 (N_2341,N_2293,N_2309);
or U2342 (N_2342,N_2323,N_2280);
nor U2343 (N_2343,N_2318,N_2283);
or U2344 (N_2344,N_2329,N_2303);
nand U2345 (N_2345,N_2319,N_2327);
and U2346 (N_2346,N_2282,N_2288);
or U2347 (N_2347,N_2296,N_2294);
nand U2348 (N_2348,N_2300,N_2307);
nor U2349 (N_2349,N_2339,N_2337);
nand U2350 (N_2350,N_2298,N_2326);
or U2351 (N_2351,N_2281,N_2312);
or U2352 (N_2352,N_2321,N_2302);
and U2353 (N_2353,N_2328,N_2306);
or U2354 (N_2354,N_2297,N_2325);
nand U2355 (N_2355,N_2334,N_2316);
nand U2356 (N_2356,N_2314,N_2305);
nand U2357 (N_2357,N_2295,N_2324);
nand U2358 (N_2358,N_2287,N_2333);
nor U2359 (N_2359,N_2313,N_2301);
or U2360 (N_2360,N_2284,N_2299);
or U2361 (N_2361,N_2317,N_2285);
nand U2362 (N_2362,N_2308,N_2304);
and U2363 (N_2363,N_2315,N_2289);
or U2364 (N_2364,N_2311,N_2332);
or U2365 (N_2365,N_2331,N_2338);
nor U2366 (N_2366,N_2320,N_2292);
or U2367 (N_2367,N_2336,N_2291);
nor U2368 (N_2368,N_2335,N_2290);
and U2369 (N_2369,N_2310,N_2330);
or U2370 (N_2370,N_2333,N_2339);
nand U2371 (N_2371,N_2325,N_2307);
and U2372 (N_2372,N_2317,N_2331);
nor U2373 (N_2373,N_2336,N_2297);
nand U2374 (N_2374,N_2329,N_2299);
nor U2375 (N_2375,N_2297,N_2333);
or U2376 (N_2376,N_2287,N_2296);
nor U2377 (N_2377,N_2294,N_2319);
or U2378 (N_2378,N_2313,N_2282);
nor U2379 (N_2379,N_2299,N_2280);
or U2380 (N_2380,N_2303,N_2326);
and U2381 (N_2381,N_2337,N_2307);
nor U2382 (N_2382,N_2307,N_2288);
or U2383 (N_2383,N_2330,N_2286);
xnor U2384 (N_2384,N_2335,N_2295);
and U2385 (N_2385,N_2327,N_2290);
and U2386 (N_2386,N_2290,N_2316);
nand U2387 (N_2387,N_2281,N_2321);
and U2388 (N_2388,N_2329,N_2338);
nand U2389 (N_2389,N_2307,N_2333);
and U2390 (N_2390,N_2317,N_2316);
nor U2391 (N_2391,N_2339,N_2302);
xnor U2392 (N_2392,N_2334,N_2317);
and U2393 (N_2393,N_2314,N_2321);
and U2394 (N_2394,N_2322,N_2302);
and U2395 (N_2395,N_2328,N_2320);
nand U2396 (N_2396,N_2306,N_2320);
or U2397 (N_2397,N_2293,N_2287);
nor U2398 (N_2398,N_2319,N_2302);
nand U2399 (N_2399,N_2309,N_2299);
or U2400 (N_2400,N_2353,N_2345);
nor U2401 (N_2401,N_2366,N_2399);
or U2402 (N_2402,N_2396,N_2373);
and U2403 (N_2403,N_2344,N_2398);
or U2404 (N_2404,N_2390,N_2350);
xnor U2405 (N_2405,N_2351,N_2383);
nor U2406 (N_2406,N_2343,N_2368);
and U2407 (N_2407,N_2347,N_2369);
nand U2408 (N_2408,N_2382,N_2358);
and U2409 (N_2409,N_2363,N_2374);
xor U2410 (N_2410,N_2365,N_2378);
or U2411 (N_2411,N_2367,N_2379);
nor U2412 (N_2412,N_2340,N_2342);
and U2413 (N_2413,N_2364,N_2357);
or U2414 (N_2414,N_2387,N_2354);
nor U2415 (N_2415,N_2395,N_2375);
nor U2416 (N_2416,N_2392,N_2362);
nand U2417 (N_2417,N_2376,N_2381);
and U2418 (N_2418,N_2397,N_2370);
and U2419 (N_2419,N_2371,N_2360);
xor U2420 (N_2420,N_2361,N_2341);
or U2421 (N_2421,N_2384,N_2348);
nor U2422 (N_2422,N_2346,N_2380);
nand U2423 (N_2423,N_2391,N_2393);
nor U2424 (N_2424,N_2372,N_2389);
and U2425 (N_2425,N_2386,N_2359);
and U2426 (N_2426,N_2394,N_2385);
or U2427 (N_2427,N_2388,N_2352);
or U2428 (N_2428,N_2349,N_2356);
nand U2429 (N_2429,N_2355,N_2377);
and U2430 (N_2430,N_2375,N_2369);
and U2431 (N_2431,N_2342,N_2396);
nand U2432 (N_2432,N_2391,N_2365);
nand U2433 (N_2433,N_2353,N_2348);
nand U2434 (N_2434,N_2374,N_2388);
or U2435 (N_2435,N_2396,N_2390);
nor U2436 (N_2436,N_2383,N_2341);
or U2437 (N_2437,N_2356,N_2383);
nand U2438 (N_2438,N_2372,N_2397);
nor U2439 (N_2439,N_2352,N_2365);
or U2440 (N_2440,N_2359,N_2395);
or U2441 (N_2441,N_2391,N_2379);
and U2442 (N_2442,N_2396,N_2374);
or U2443 (N_2443,N_2394,N_2351);
nand U2444 (N_2444,N_2349,N_2372);
and U2445 (N_2445,N_2388,N_2392);
and U2446 (N_2446,N_2396,N_2372);
or U2447 (N_2447,N_2343,N_2399);
or U2448 (N_2448,N_2386,N_2380);
nand U2449 (N_2449,N_2345,N_2391);
nor U2450 (N_2450,N_2377,N_2375);
and U2451 (N_2451,N_2357,N_2348);
xnor U2452 (N_2452,N_2369,N_2353);
or U2453 (N_2453,N_2394,N_2341);
nor U2454 (N_2454,N_2389,N_2399);
nand U2455 (N_2455,N_2377,N_2346);
nor U2456 (N_2456,N_2382,N_2397);
and U2457 (N_2457,N_2343,N_2355);
nand U2458 (N_2458,N_2345,N_2350);
and U2459 (N_2459,N_2367,N_2396);
or U2460 (N_2460,N_2406,N_2432);
nor U2461 (N_2461,N_2408,N_2459);
nand U2462 (N_2462,N_2430,N_2421);
nand U2463 (N_2463,N_2419,N_2434);
and U2464 (N_2464,N_2410,N_2424);
nand U2465 (N_2465,N_2439,N_2422);
nor U2466 (N_2466,N_2401,N_2423);
or U2467 (N_2467,N_2437,N_2416);
xnor U2468 (N_2468,N_2405,N_2418);
nand U2469 (N_2469,N_2448,N_2457);
and U2470 (N_2470,N_2428,N_2429);
or U2471 (N_2471,N_2454,N_2438);
nand U2472 (N_2472,N_2403,N_2458);
and U2473 (N_2473,N_2414,N_2452);
and U2474 (N_2474,N_2443,N_2451);
nor U2475 (N_2475,N_2425,N_2413);
or U2476 (N_2476,N_2412,N_2435);
and U2477 (N_2477,N_2415,N_2400);
nor U2478 (N_2478,N_2455,N_2450);
nor U2479 (N_2479,N_2447,N_2420);
or U2480 (N_2480,N_2449,N_2441);
nor U2481 (N_2481,N_2417,N_2404);
nand U2482 (N_2482,N_2445,N_2444);
nand U2483 (N_2483,N_2453,N_2442);
or U2484 (N_2484,N_2433,N_2436);
or U2485 (N_2485,N_2426,N_2402);
and U2486 (N_2486,N_2407,N_2431);
or U2487 (N_2487,N_2446,N_2409);
nor U2488 (N_2488,N_2456,N_2440);
nor U2489 (N_2489,N_2427,N_2411);
or U2490 (N_2490,N_2449,N_2415);
and U2491 (N_2491,N_2429,N_2450);
nor U2492 (N_2492,N_2419,N_2459);
nand U2493 (N_2493,N_2404,N_2429);
or U2494 (N_2494,N_2421,N_2425);
and U2495 (N_2495,N_2416,N_2403);
nand U2496 (N_2496,N_2435,N_2414);
and U2497 (N_2497,N_2448,N_2437);
and U2498 (N_2498,N_2426,N_2407);
nand U2499 (N_2499,N_2451,N_2416);
xor U2500 (N_2500,N_2416,N_2450);
and U2501 (N_2501,N_2452,N_2431);
or U2502 (N_2502,N_2448,N_2420);
nand U2503 (N_2503,N_2435,N_2449);
nor U2504 (N_2504,N_2425,N_2416);
nor U2505 (N_2505,N_2404,N_2405);
or U2506 (N_2506,N_2401,N_2441);
nand U2507 (N_2507,N_2449,N_2456);
or U2508 (N_2508,N_2446,N_2420);
nand U2509 (N_2509,N_2421,N_2418);
nand U2510 (N_2510,N_2409,N_2452);
or U2511 (N_2511,N_2401,N_2400);
nor U2512 (N_2512,N_2404,N_2419);
nor U2513 (N_2513,N_2413,N_2402);
and U2514 (N_2514,N_2441,N_2420);
and U2515 (N_2515,N_2434,N_2402);
and U2516 (N_2516,N_2415,N_2456);
and U2517 (N_2517,N_2411,N_2447);
nand U2518 (N_2518,N_2418,N_2453);
nor U2519 (N_2519,N_2453,N_2424);
nor U2520 (N_2520,N_2513,N_2468);
nand U2521 (N_2521,N_2493,N_2463);
or U2522 (N_2522,N_2471,N_2517);
and U2523 (N_2523,N_2462,N_2496);
and U2524 (N_2524,N_2486,N_2469);
nor U2525 (N_2525,N_2488,N_2478);
nand U2526 (N_2526,N_2503,N_2483);
nand U2527 (N_2527,N_2470,N_2489);
xnor U2528 (N_2528,N_2499,N_2514);
or U2529 (N_2529,N_2491,N_2490);
or U2530 (N_2530,N_2508,N_2467);
nand U2531 (N_2531,N_2504,N_2461);
and U2532 (N_2532,N_2485,N_2473);
nand U2533 (N_2533,N_2472,N_2482);
or U2534 (N_2534,N_2495,N_2480);
and U2535 (N_2535,N_2500,N_2518);
or U2536 (N_2536,N_2507,N_2506);
and U2537 (N_2537,N_2501,N_2498);
nand U2538 (N_2538,N_2484,N_2464);
nand U2539 (N_2539,N_2519,N_2502);
and U2540 (N_2540,N_2476,N_2465);
nor U2541 (N_2541,N_2515,N_2512);
and U2542 (N_2542,N_2479,N_2505);
xnor U2543 (N_2543,N_2510,N_2511);
nand U2544 (N_2544,N_2475,N_2497);
and U2545 (N_2545,N_2516,N_2509);
and U2546 (N_2546,N_2494,N_2460);
or U2547 (N_2547,N_2477,N_2474);
nor U2548 (N_2548,N_2481,N_2492);
nor U2549 (N_2549,N_2466,N_2487);
or U2550 (N_2550,N_2515,N_2499);
nand U2551 (N_2551,N_2499,N_2487);
and U2552 (N_2552,N_2479,N_2492);
and U2553 (N_2553,N_2462,N_2481);
or U2554 (N_2554,N_2461,N_2509);
and U2555 (N_2555,N_2485,N_2490);
nand U2556 (N_2556,N_2477,N_2505);
or U2557 (N_2557,N_2497,N_2466);
or U2558 (N_2558,N_2475,N_2518);
nand U2559 (N_2559,N_2480,N_2491);
nand U2560 (N_2560,N_2506,N_2513);
nand U2561 (N_2561,N_2484,N_2479);
nand U2562 (N_2562,N_2516,N_2470);
or U2563 (N_2563,N_2480,N_2469);
nand U2564 (N_2564,N_2462,N_2487);
nor U2565 (N_2565,N_2476,N_2510);
nor U2566 (N_2566,N_2508,N_2476);
and U2567 (N_2567,N_2500,N_2495);
nor U2568 (N_2568,N_2488,N_2461);
and U2569 (N_2569,N_2519,N_2487);
or U2570 (N_2570,N_2470,N_2486);
nand U2571 (N_2571,N_2498,N_2511);
and U2572 (N_2572,N_2485,N_2500);
nand U2573 (N_2573,N_2475,N_2464);
and U2574 (N_2574,N_2472,N_2517);
or U2575 (N_2575,N_2478,N_2503);
or U2576 (N_2576,N_2484,N_2514);
and U2577 (N_2577,N_2509,N_2486);
nor U2578 (N_2578,N_2508,N_2468);
or U2579 (N_2579,N_2509,N_2518);
nand U2580 (N_2580,N_2575,N_2563);
nor U2581 (N_2581,N_2550,N_2553);
and U2582 (N_2582,N_2547,N_2528);
nand U2583 (N_2583,N_2578,N_2574);
nor U2584 (N_2584,N_2546,N_2535);
nor U2585 (N_2585,N_2571,N_2572);
or U2586 (N_2586,N_2576,N_2541);
and U2587 (N_2587,N_2551,N_2562);
nor U2588 (N_2588,N_2554,N_2531);
nand U2589 (N_2589,N_2565,N_2560);
nor U2590 (N_2590,N_2561,N_2543);
or U2591 (N_2591,N_2564,N_2537);
nor U2592 (N_2592,N_2558,N_2567);
and U2593 (N_2593,N_2536,N_2577);
nand U2594 (N_2594,N_2548,N_2570);
nand U2595 (N_2595,N_2542,N_2568);
nand U2596 (N_2596,N_2538,N_2579);
or U2597 (N_2597,N_2534,N_2526);
or U2598 (N_2598,N_2533,N_2525);
and U2599 (N_2599,N_2545,N_2573);
nor U2600 (N_2600,N_2569,N_2530);
nor U2601 (N_2601,N_2520,N_2521);
or U2602 (N_2602,N_2557,N_2555);
nor U2603 (N_2603,N_2539,N_2566);
nand U2604 (N_2604,N_2549,N_2559);
nor U2605 (N_2605,N_2552,N_2540);
or U2606 (N_2606,N_2522,N_2544);
or U2607 (N_2607,N_2524,N_2523);
nand U2608 (N_2608,N_2532,N_2556);
nand U2609 (N_2609,N_2527,N_2529);
nor U2610 (N_2610,N_2563,N_2567);
nand U2611 (N_2611,N_2572,N_2547);
nor U2612 (N_2612,N_2530,N_2549);
nor U2613 (N_2613,N_2529,N_2567);
and U2614 (N_2614,N_2561,N_2525);
and U2615 (N_2615,N_2538,N_2569);
nor U2616 (N_2616,N_2562,N_2576);
and U2617 (N_2617,N_2533,N_2578);
and U2618 (N_2618,N_2565,N_2566);
or U2619 (N_2619,N_2571,N_2575);
and U2620 (N_2620,N_2566,N_2536);
or U2621 (N_2621,N_2559,N_2544);
and U2622 (N_2622,N_2553,N_2560);
and U2623 (N_2623,N_2550,N_2559);
and U2624 (N_2624,N_2567,N_2545);
and U2625 (N_2625,N_2532,N_2524);
and U2626 (N_2626,N_2530,N_2523);
or U2627 (N_2627,N_2565,N_2543);
or U2628 (N_2628,N_2541,N_2536);
nor U2629 (N_2629,N_2554,N_2536);
or U2630 (N_2630,N_2567,N_2556);
nand U2631 (N_2631,N_2568,N_2539);
and U2632 (N_2632,N_2553,N_2574);
nand U2633 (N_2633,N_2547,N_2558);
or U2634 (N_2634,N_2521,N_2546);
or U2635 (N_2635,N_2533,N_2522);
and U2636 (N_2636,N_2566,N_2568);
nand U2637 (N_2637,N_2533,N_2529);
nor U2638 (N_2638,N_2572,N_2567);
and U2639 (N_2639,N_2574,N_2533);
nor U2640 (N_2640,N_2636,N_2611);
and U2641 (N_2641,N_2632,N_2627);
or U2642 (N_2642,N_2607,N_2603);
nor U2643 (N_2643,N_2582,N_2597);
or U2644 (N_2644,N_2629,N_2590);
nor U2645 (N_2645,N_2609,N_2614);
nand U2646 (N_2646,N_2638,N_2588);
nand U2647 (N_2647,N_2591,N_2595);
nor U2648 (N_2648,N_2628,N_2624);
nand U2649 (N_2649,N_2598,N_2620);
xor U2650 (N_2650,N_2608,N_2586);
nor U2651 (N_2651,N_2613,N_2605);
and U2652 (N_2652,N_2615,N_2630);
nand U2653 (N_2653,N_2634,N_2581);
and U2654 (N_2654,N_2610,N_2625);
nand U2655 (N_2655,N_2618,N_2589);
and U2656 (N_2656,N_2593,N_2587);
and U2657 (N_2657,N_2617,N_2639);
and U2658 (N_2658,N_2626,N_2580);
and U2659 (N_2659,N_2622,N_2612);
or U2660 (N_2660,N_2596,N_2599);
or U2661 (N_2661,N_2637,N_2606);
nand U2662 (N_2662,N_2631,N_2623);
or U2663 (N_2663,N_2600,N_2621);
or U2664 (N_2664,N_2619,N_2616);
nor U2665 (N_2665,N_2635,N_2592);
or U2666 (N_2666,N_2584,N_2594);
or U2667 (N_2667,N_2583,N_2602);
or U2668 (N_2668,N_2601,N_2604);
or U2669 (N_2669,N_2585,N_2633);
and U2670 (N_2670,N_2621,N_2629);
and U2671 (N_2671,N_2624,N_2605);
nand U2672 (N_2672,N_2612,N_2611);
nand U2673 (N_2673,N_2588,N_2587);
nand U2674 (N_2674,N_2588,N_2626);
nand U2675 (N_2675,N_2638,N_2585);
nand U2676 (N_2676,N_2612,N_2586);
or U2677 (N_2677,N_2635,N_2630);
nor U2678 (N_2678,N_2606,N_2635);
nand U2679 (N_2679,N_2590,N_2581);
nand U2680 (N_2680,N_2601,N_2607);
nand U2681 (N_2681,N_2583,N_2629);
nand U2682 (N_2682,N_2617,N_2607);
nand U2683 (N_2683,N_2610,N_2635);
and U2684 (N_2684,N_2591,N_2609);
or U2685 (N_2685,N_2591,N_2623);
xor U2686 (N_2686,N_2615,N_2618);
and U2687 (N_2687,N_2625,N_2617);
or U2688 (N_2688,N_2587,N_2634);
nor U2689 (N_2689,N_2603,N_2598);
nand U2690 (N_2690,N_2635,N_2605);
or U2691 (N_2691,N_2619,N_2607);
nand U2692 (N_2692,N_2627,N_2597);
nand U2693 (N_2693,N_2585,N_2590);
nand U2694 (N_2694,N_2626,N_2604);
nand U2695 (N_2695,N_2594,N_2638);
and U2696 (N_2696,N_2580,N_2613);
and U2697 (N_2697,N_2629,N_2610);
or U2698 (N_2698,N_2610,N_2614);
nand U2699 (N_2699,N_2632,N_2639);
nor U2700 (N_2700,N_2645,N_2657);
and U2701 (N_2701,N_2681,N_2690);
nand U2702 (N_2702,N_2641,N_2688);
nor U2703 (N_2703,N_2654,N_2675);
nor U2704 (N_2704,N_2647,N_2656);
and U2705 (N_2705,N_2676,N_2648);
nand U2706 (N_2706,N_2662,N_2670);
and U2707 (N_2707,N_2696,N_2673);
nor U2708 (N_2708,N_2680,N_2698);
and U2709 (N_2709,N_2695,N_2644);
or U2710 (N_2710,N_2682,N_2667);
and U2711 (N_2711,N_2691,N_2699);
or U2712 (N_2712,N_2684,N_2649);
nor U2713 (N_2713,N_2678,N_2646);
and U2714 (N_2714,N_2693,N_2686);
and U2715 (N_2715,N_2689,N_2692);
and U2716 (N_2716,N_2687,N_2672);
nor U2717 (N_2717,N_2642,N_2694);
or U2718 (N_2718,N_2651,N_2664);
and U2719 (N_2719,N_2659,N_2669);
and U2720 (N_2720,N_2677,N_2652);
nand U2721 (N_2721,N_2643,N_2655);
nor U2722 (N_2722,N_2685,N_2661);
nor U2723 (N_2723,N_2665,N_2697);
nor U2724 (N_2724,N_2640,N_2660);
and U2725 (N_2725,N_2671,N_2653);
nor U2726 (N_2726,N_2668,N_2674);
nand U2727 (N_2727,N_2650,N_2658);
and U2728 (N_2728,N_2666,N_2663);
or U2729 (N_2729,N_2683,N_2679);
nor U2730 (N_2730,N_2640,N_2669);
nand U2731 (N_2731,N_2657,N_2641);
xor U2732 (N_2732,N_2687,N_2697);
nand U2733 (N_2733,N_2668,N_2649);
or U2734 (N_2734,N_2670,N_2694);
nand U2735 (N_2735,N_2675,N_2670);
and U2736 (N_2736,N_2647,N_2667);
or U2737 (N_2737,N_2671,N_2646);
nand U2738 (N_2738,N_2690,N_2666);
and U2739 (N_2739,N_2670,N_2681);
or U2740 (N_2740,N_2673,N_2678);
nor U2741 (N_2741,N_2677,N_2646);
nor U2742 (N_2742,N_2667,N_2693);
nand U2743 (N_2743,N_2687,N_2660);
nand U2744 (N_2744,N_2659,N_2661);
and U2745 (N_2745,N_2651,N_2668);
and U2746 (N_2746,N_2667,N_2652);
or U2747 (N_2747,N_2694,N_2648);
nand U2748 (N_2748,N_2698,N_2663);
nand U2749 (N_2749,N_2673,N_2689);
nand U2750 (N_2750,N_2658,N_2655);
and U2751 (N_2751,N_2691,N_2685);
and U2752 (N_2752,N_2690,N_2699);
nor U2753 (N_2753,N_2699,N_2641);
xor U2754 (N_2754,N_2695,N_2663);
or U2755 (N_2755,N_2699,N_2672);
or U2756 (N_2756,N_2672,N_2648);
or U2757 (N_2757,N_2681,N_2654);
and U2758 (N_2758,N_2679,N_2685);
and U2759 (N_2759,N_2664,N_2662);
nor U2760 (N_2760,N_2751,N_2720);
or U2761 (N_2761,N_2735,N_2757);
nand U2762 (N_2762,N_2717,N_2701);
nand U2763 (N_2763,N_2716,N_2700);
nand U2764 (N_2764,N_2750,N_2713);
and U2765 (N_2765,N_2709,N_2712);
nor U2766 (N_2766,N_2744,N_2737);
or U2767 (N_2767,N_2711,N_2724);
nand U2768 (N_2768,N_2726,N_2719);
xnor U2769 (N_2769,N_2759,N_2708);
nor U2770 (N_2770,N_2748,N_2729);
xnor U2771 (N_2771,N_2739,N_2725);
nand U2772 (N_2772,N_2722,N_2758);
nor U2773 (N_2773,N_2738,N_2703);
xor U2774 (N_2774,N_2733,N_2741);
nand U2775 (N_2775,N_2753,N_2728);
nand U2776 (N_2776,N_2756,N_2730);
or U2777 (N_2777,N_2743,N_2704);
nor U2778 (N_2778,N_2715,N_2746);
and U2779 (N_2779,N_2749,N_2734);
or U2780 (N_2780,N_2742,N_2752);
and U2781 (N_2781,N_2706,N_2710);
nand U2782 (N_2782,N_2721,N_2707);
nand U2783 (N_2783,N_2745,N_2714);
xor U2784 (N_2784,N_2740,N_2705);
nand U2785 (N_2785,N_2718,N_2732);
and U2786 (N_2786,N_2723,N_2731);
nand U2787 (N_2787,N_2736,N_2702);
and U2788 (N_2788,N_2727,N_2754);
and U2789 (N_2789,N_2747,N_2755);
nand U2790 (N_2790,N_2711,N_2721);
nand U2791 (N_2791,N_2751,N_2724);
and U2792 (N_2792,N_2711,N_2759);
nor U2793 (N_2793,N_2722,N_2731);
or U2794 (N_2794,N_2746,N_2747);
or U2795 (N_2795,N_2721,N_2705);
and U2796 (N_2796,N_2759,N_2717);
or U2797 (N_2797,N_2748,N_2726);
and U2798 (N_2798,N_2753,N_2756);
and U2799 (N_2799,N_2708,N_2707);
nand U2800 (N_2800,N_2717,N_2729);
nor U2801 (N_2801,N_2711,N_2732);
xor U2802 (N_2802,N_2756,N_2707);
nor U2803 (N_2803,N_2712,N_2756);
or U2804 (N_2804,N_2759,N_2755);
or U2805 (N_2805,N_2750,N_2712);
nor U2806 (N_2806,N_2720,N_2702);
and U2807 (N_2807,N_2752,N_2732);
nand U2808 (N_2808,N_2736,N_2715);
and U2809 (N_2809,N_2748,N_2717);
or U2810 (N_2810,N_2742,N_2733);
and U2811 (N_2811,N_2706,N_2747);
and U2812 (N_2812,N_2712,N_2733);
or U2813 (N_2813,N_2736,N_2725);
and U2814 (N_2814,N_2728,N_2715);
or U2815 (N_2815,N_2702,N_2735);
nand U2816 (N_2816,N_2756,N_2718);
nand U2817 (N_2817,N_2752,N_2736);
nor U2818 (N_2818,N_2743,N_2717);
nor U2819 (N_2819,N_2759,N_2752);
nand U2820 (N_2820,N_2797,N_2817);
or U2821 (N_2821,N_2814,N_2818);
and U2822 (N_2822,N_2777,N_2810);
nor U2823 (N_2823,N_2796,N_2764);
nor U2824 (N_2824,N_2783,N_2779);
or U2825 (N_2825,N_2763,N_2809);
or U2826 (N_2826,N_2771,N_2761);
and U2827 (N_2827,N_2792,N_2781);
and U2828 (N_2828,N_2767,N_2766);
nor U2829 (N_2829,N_2778,N_2782);
nand U2830 (N_2830,N_2785,N_2775);
nand U2831 (N_2831,N_2770,N_2816);
or U2832 (N_2832,N_2798,N_2794);
and U2833 (N_2833,N_2765,N_2784);
nand U2834 (N_2834,N_2800,N_2788);
nor U2835 (N_2835,N_2791,N_2815);
nand U2836 (N_2836,N_2806,N_2802);
or U2837 (N_2837,N_2774,N_2768);
or U2838 (N_2838,N_2786,N_2801);
and U2839 (N_2839,N_2804,N_2762);
nand U2840 (N_2840,N_2803,N_2805);
nor U2841 (N_2841,N_2807,N_2811);
nor U2842 (N_2842,N_2772,N_2813);
nand U2843 (N_2843,N_2808,N_2787);
and U2844 (N_2844,N_2799,N_2760);
nand U2845 (N_2845,N_2780,N_2789);
nor U2846 (N_2846,N_2773,N_2776);
or U2847 (N_2847,N_2795,N_2819);
or U2848 (N_2848,N_2790,N_2769);
or U2849 (N_2849,N_2793,N_2812);
nand U2850 (N_2850,N_2773,N_2804);
nor U2851 (N_2851,N_2798,N_2796);
nand U2852 (N_2852,N_2783,N_2794);
nand U2853 (N_2853,N_2814,N_2775);
nor U2854 (N_2854,N_2810,N_2806);
or U2855 (N_2855,N_2817,N_2814);
and U2856 (N_2856,N_2819,N_2783);
nand U2857 (N_2857,N_2782,N_2780);
and U2858 (N_2858,N_2762,N_2790);
or U2859 (N_2859,N_2802,N_2763);
nor U2860 (N_2860,N_2810,N_2811);
nand U2861 (N_2861,N_2810,N_2779);
or U2862 (N_2862,N_2807,N_2800);
nand U2863 (N_2863,N_2780,N_2794);
nand U2864 (N_2864,N_2784,N_2812);
and U2865 (N_2865,N_2782,N_2767);
nor U2866 (N_2866,N_2761,N_2799);
nand U2867 (N_2867,N_2780,N_2760);
xor U2868 (N_2868,N_2792,N_2805);
nor U2869 (N_2869,N_2815,N_2817);
and U2870 (N_2870,N_2773,N_2817);
or U2871 (N_2871,N_2800,N_2762);
and U2872 (N_2872,N_2800,N_2790);
and U2873 (N_2873,N_2772,N_2768);
nor U2874 (N_2874,N_2811,N_2778);
or U2875 (N_2875,N_2814,N_2799);
nor U2876 (N_2876,N_2815,N_2763);
or U2877 (N_2877,N_2818,N_2791);
xor U2878 (N_2878,N_2767,N_2787);
or U2879 (N_2879,N_2813,N_2805);
nand U2880 (N_2880,N_2858,N_2868);
or U2881 (N_2881,N_2833,N_2844);
or U2882 (N_2882,N_2829,N_2852);
nor U2883 (N_2883,N_2871,N_2873);
nor U2884 (N_2884,N_2848,N_2864);
nand U2885 (N_2885,N_2867,N_2846);
nand U2886 (N_2886,N_2842,N_2824);
nor U2887 (N_2887,N_2835,N_2879);
and U2888 (N_2888,N_2832,N_2838);
nor U2889 (N_2889,N_2825,N_2859);
nor U2890 (N_2890,N_2872,N_2831);
nor U2891 (N_2891,N_2822,N_2821);
or U2892 (N_2892,N_2861,N_2860);
or U2893 (N_2893,N_2830,N_2840);
nor U2894 (N_2894,N_2828,N_2862);
nor U2895 (N_2895,N_2853,N_2869);
nand U2896 (N_2896,N_2854,N_2856);
and U2897 (N_2897,N_2875,N_2865);
nor U2898 (N_2898,N_2836,N_2866);
nor U2899 (N_2899,N_2877,N_2855);
nand U2900 (N_2900,N_2843,N_2837);
and U2901 (N_2901,N_2876,N_2823);
nor U2902 (N_2902,N_2834,N_2874);
nand U2903 (N_2903,N_2851,N_2820);
or U2904 (N_2904,N_2839,N_2870);
or U2905 (N_2905,N_2847,N_2878);
xnor U2906 (N_2906,N_2863,N_2850);
nor U2907 (N_2907,N_2857,N_2845);
and U2908 (N_2908,N_2827,N_2841);
nand U2909 (N_2909,N_2826,N_2849);
nor U2910 (N_2910,N_2820,N_2862);
nor U2911 (N_2911,N_2861,N_2824);
and U2912 (N_2912,N_2873,N_2824);
or U2913 (N_2913,N_2871,N_2834);
or U2914 (N_2914,N_2856,N_2826);
xnor U2915 (N_2915,N_2835,N_2868);
and U2916 (N_2916,N_2868,N_2821);
or U2917 (N_2917,N_2846,N_2851);
nor U2918 (N_2918,N_2855,N_2862);
nor U2919 (N_2919,N_2854,N_2875);
nand U2920 (N_2920,N_2855,N_2852);
nor U2921 (N_2921,N_2852,N_2862);
or U2922 (N_2922,N_2826,N_2850);
nor U2923 (N_2923,N_2874,N_2851);
xnor U2924 (N_2924,N_2872,N_2839);
and U2925 (N_2925,N_2821,N_2862);
nor U2926 (N_2926,N_2854,N_2844);
or U2927 (N_2927,N_2852,N_2860);
xnor U2928 (N_2928,N_2868,N_2879);
nand U2929 (N_2929,N_2839,N_2827);
nand U2930 (N_2930,N_2845,N_2877);
nand U2931 (N_2931,N_2858,N_2852);
and U2932 (N_2932,N_2844,N_2852);
nand U2933 (N_2933,N_2828,N_2843);
nand U2934 (N_2934,N_2853,N_2875);
and U2935 (N_2935,N_2828,N_2848);
nand U2936 (N_2936,N_2845,N_2843);
and U2937 (N_2937,N_2858,N_2872);
or U2938 (N_2938,N_2850,N_2842);
xnor U2939 (N_2939,N_2865,N_2824);
xnor U2940 (N_2940,N_2882,N_2890);
nor U2941 (N_2941,N_2938,N_2933);
and U2942 (N_2942,N_2910,N_2925);
and U2943 (N_2943,N_2916,N_2896);
and U2944 (N_2944,N_2893,N_2892);
xnor U2945 (N_2945,N_2926,N_2904);
nor U2946 (N_2946,N_2935,N_2880);
nor U2947 (N_2947,N_2936,N_2889);
and U2948 (N_2948,N_2923,N_2899);
nor U2949 (N_2949,N_2895,N_2927);
xnor U2950 (N_2950,N_2937,N_2912);
nor U2951 (N_2951,N_2886,N_2883);
xnor U2952 (N_2952,N_2932,N_2888);
nand U2953 (N_2953,N_2934,N_2930);
nor U2954 (N_2954,N_2931,N_2907);
nor U2955 (N_2955,N_2920,N_2928);
nand U2956 (N_2956,N_2902,N_2911);
nor U2957 (N_2957,N_2918,N_2908);
and U2958 (N_2958,N_2913,N_2887);
and U2959 (N_2959,N_2906,N_2897);
nor U2960 (N_2960,N_2898,N_2884);
nor U2961 (N_2961,N_2922,N_2891);
nor U2962 (N_2962,N_2914,N_2900);
and U2963 (N_2963,N_2909,N_2881);
or U2964 (N_2964,N_2885,N_2901);
nand U2965 (N_2965,N_2921,N_2924);
nand U2966 (N_2966,N_2917,N_2915);
and U2967 (N_2967,N_2894,N_2939);
and U2968 (N_2968,N_2905,N_2903);
nor U2969 (N_2969,N_2919,N_2929);
nor U2970 (N_2970,N_2891,N_2892);
xor U2971 (N_2971,N_2939,N_2880);
and U2972 (N_2972,N_2890,N_2918);
xnor U2973 (N_2973,N_2886,N_2890);
nand U2974 (N_2974,N_2901,N_2894);
and U2975 (N_2975,N_2917,N_2916);
and U2976 (N_2976,N_2915,N_2909);
nor U2977 (N_2977,N_2938,N_2884);
nor U2978 (N_2978,N_2900,N_2890);
nand U2979 (N_2979,N_2889,N_2926);
nor U2980 (N_2980,N_2885,N_2937);
nor U2981 (N_2981,N_2910,N_2889);
nor U2982 (N_2982,N_2888,N_2930);
nor U2983 (N_2983,N_2918,N_2920);
nand U2984 (N_2984,N_2889,N_2935);
or U2985 (N_2985,N_2917,N_2919);
and U2986 (N_2986,N_2892,N_2938);
nand U2987 (N_2987,N_2916,N_2918);
and U2988 (N_2988,N_2921,N_2890);
or U2989 (N_2989,N_2893,N_2884);
or U2990 (N_2990,N_2936,N_2930);
or U2991 (N_2991,N_2896,N_2882);
or U2992 (N_2992,N_2880,N_2918);
nor U2993 (N_2993,N_2915,N_2905);
nor U2994 (N_2994,N_2883,N_2896);
nand U2995 (N_2995,N_2923,N_2906);
nor U2996 (N_2996,N_2906,N_2907);
or U2997 (N_2997,N_2901,N_2939);
nor U2998 (N_2998,N_2907,N_2895);
or U2999 (N_2999,N_2917,N_2933);
and UO_0 (O_0,N_2982,N_2950);
nand UO_1 (O_1,N_2979,N_2991);
nor UO_2 (O_2,N_2961,N_2945);
and UO_3 (O_3,N_2942,N_2973);
and UO_4 (O_4,N_2970,N_2993);
nand UO_5 (O_5,N_2952,N_2965);
nor UO_6 (O_6,N_2963,N_2994);
or UO_7 (O_7,N_2940,N_2969);
nor UO_8 (O_8,N_2948,N_2955);
or UO_9 (O_9,N_2987,N_2975);
or UO_10 (O_10,N_2981,N_2960);
nand UO_11 (O_11,N_2944,N_2989);
nand UO_12 (O_12,N_2968,N_2962);
nand UO_13 (O_13,N_2958,N_2990);
and UO_14 (O_14,N_2951,N_2985);
and UO_15 (O_15,N_2947,N_2984);
nor UO_16 (O_16,N_2967,N_2941);
and UO_17 (O_17,N_2980,N_2978);
and UO_18 (O_18,N_2957,N_2949);
or UO_19 (O_19,N_2943,N_2976);
and UO_20 (O_20,N_2966,N_2983);
nand UO_21 (O_21,N_2946,N_2996);
nand UO_22 (O_22,N_2974,N_2964);
nor UO_23 (O_23,N_2986,N_2972);
nor UO_24 (O_24,N_2953,N_2971);
or UO_25 (O_25,N_2988,N_2999);
or UO_26 (O_26,N_2959,N_2954);
nor UO_27 (O_27,N_2956,N_2995);
or UO_28 (O_28,N_2992,N_2998);
and UO_29 (O_29,N_2977,N_2997);
and UO_30 (O_30,N_2985,N_2972);
or UO_31 (O_31,N_2991,N_2996);
and UO_32 (O_32,N_2945,N_2976);
or UO_33 (O_33,N_2965,N_2982);
nor UO_34 (O_34,N_2961,N_2984);
and UO_35 (O_35,N_2942,N_2963);
and UO_36 (O_36,N_2953,N_2981);
or UO_37 (O_37,N_2970,N_2964);
nor UO_38 (O_38,N_2990,N_2999);
and UO_39 (O_39,N_2980,N_2989);
and UO_40 (O_40,N_2986,N_2977);
or UO_41 (O_41,N_2994,N_2987);
nand UO_42 (O_42,N_2999,N_2953);
or UO_43 (O_43,N_2945,N_2949);
and UO_44 (O_44,N_2996,N_2975);
nand UO_45 (O_45,N_2953,N_2988);
nand UO_46 (O_46,N_2946,N_2949);
nand UO_47 (O_47,N_2952,N_2984);
or UO_48 (O_48,N_2944,N_2980);
and UO_49 (O_49,N_2992,N_2949);
and UO_50 (O_50,N_2951,N_2943);
or UO_51 (O_51,N_2994,N_2995);
nand UO_52 (O_52,N_2985,N_2942);
and UO_53 (O_53,N_2999,N_2993);
or UO_54 (O_54,N_2984,N_2959);
or UO_55 (O_55,N_2982,N_2979);
xnor UO_56 (O_56,N_2984,N_2948);
nor UO_57 (O_57,N_2983,N_2950);
nor UO_58 (O_58,N_2946,N_2977);
nand UO_59 (O_59,N_2991,N_2940);
or UO_60 (O_60,N_2974,N_2958);
or UO_61 (O_61,N_2991,N_2971);
and UO_62 (O_62,N_2990,N_2986);
or UO_63 (O_63,N_2994,N_2973);
or UO_64 (O_64,N_2975,N_2974);
and UO_65 (O_65,N_2959,N_2955);
nand UO_66 (O_66,N_2995,N_2971);
and UO_67 (O_67,N_2972,N_2973);
or UO_68 (O_68,N_2947,N_2951);
nand UO_69 (O_69,N_2958,N_2940);
nand UO_70 (O_70,N_2955,N_2970);
and UO_71 (O_71,N_2961,N_2982);
or UO_72 (O_72,N_2975,N_2982);
or UO_73 (O_73,N_2964,N_2994);
and UO_74 (O_74,N_2955,N_2961);
nand UO_75 (O_75,N_2985,N_2987);
nor UO_76 (O_76,N_2948,N_2973);
nand UO_77 (O_77,N_2966,N_2974);
nor UO_78 (O_78,N_2982,N_2963);
or UO_79 (O_79,N_2982,N_2996);
nor UO_80 (O_80,N_2992,N_2981);
nor UO_81 (O_81,N_2978,N_2984);
nand UO_82 (O_82,N_2952,N_2948);
or UO_83 (O_83,N_2940,N_2961);
nand UO_84 (O_84,N_2969,N_2989);
or UO_85 (O_85,N_2952,N_2993);
nand UO_86 (O_86,N_2977,N_2967);
nor UO_87 (O_87,N_2949,N_2996);
nor UO_88 (O_88,N_2991,N_2990);
nand UO_89 (O_89,N_2985,N_2993);
nor UO_90 (O_90,N_2943,N_2945);
nor UO_91 (O_91,N_2987,N_2972);
nor UO_92 (O_92,N_2990,N_2972);
and UO_93 (O_93,N_2970,N_2947);
nand UO_94 (O_94,N_2984,N_2983);
or UO_95 (O_95,N_2958,N_2952);
xnor UO_96 (O_96,N_2980,N_2962);
nor UO_97 (O_97,N_2973,N_2983);
nor UO_98 (O_98,N_2951,N_2984);
nor UO_99 (O_99,N_2987,N_2968);
nand UO_100 (O_100,N_2963,N_2960);
and UO_101 (O_101,N_2984,N_2955);
nand UO_102 (O_102,N_2944,N_2993);
nor UO_103 (O_103,N_2984,N_2954);
or UO_104 (O_104,N_2945,N_2983);
and UO_105 (O_105,N_2968,N_2974);
nor UO_106 (O_106,N_2967,N_2950);
and UO_107 (O_107,N_2980,N_2972);
nor UO_108 (O_108,N_2944,N_2983);
nor UO_109 (O_109,N_2995,N_2997);
nor UO_110 (O_110,N_2987,N_2981);
nor UO_111 (O_111,N_2980,N_2940);
and UO_112 (O_112,N_2994,N_2972);
nor UO_113 (O_113,N_2974,N_2952);
or UO_114 (O_114,N_2981,N_2989);
or UO_115 (O_115,N_2959,N_2957);
nand UO_116 (O_116,N_2951,N_2959);
or UO_117 (O_117,N_2983,N_2963);
and UO_118 (O_118,N_2977,N_2949);
or UO_119 (O_119,N_2953,N_2973);
or UO_120 (O_120,N_2991,N_2975);
nand UO_121 (O_121,N_2941,N_2943);
nand UO_122 (O_122,N_2994,N_2946);
nor UO_123 (O_123,N_2964,N_2998);
nand UO_124 (O_124,N_2973,N_2969);
nor UO_125 (O_125,N_2965,N_2991);
or UO_126 (O_126,N_2981,N_2970);
nor UO_127 (O_127,N_2996,N_2965);
nand UO_128 (O_128,N_2980,N_2977);
nand UO_129 (O_129,N_2973,N_2991);
nor UO_130 (O_130,N_2959,N_2973);
or UO_131 (O_131,N_2992,N_2942);
nor UO_132 (O_132,N_2977,N_2988);
or UO_133 (O_133,N_2989,N_2982);
nand UO_134 (O_134,N_2998,N_2959);
or UO_135 (O_135,N_2940,N_2950);
and UO_136 (O_136,N_2950,N_2999);
and UO_137 (O_137,N_2998,N_2989);
nand UO_138 (O_138,N_2962,N_2958);
or UO_139 (O_139,N_2969,N_2992);
nand UO_140 (O_140,N_2995,N_2970);
and UO_141 (O_141,N_2977,N_2953);
and UO_142 (O_142,N_2954,N_2982);
nand UO_143 (O_143,N_2986,N_2954);
nor UO_144 (O_144,N_2980,N_2982);
and UO_145 (O_145,N_2944,N_2974);
and UO_146 (O_146,N_2950,N_2943);
or UO_147 (O_147,N_2958,N_2968);
nand UO_148 (O_148,N_2958,N_2942);
or UO_149 (O_149,N_2966,N_2964);
or UO_150 (O_150,N_2949,N_2994);
or UO_151 (O_151,N_2961,N_2954);
and UO_152 (O_152,N_2968,N_2953);
nor UO_153 (O_153,N_2967,N_2993);
nor UO_154 (O_154,N_2974,N_2979);
or UO_155 (O_155,N_2986,N_2975);
nand UO_156 (O_156,N_2982,N_2940);
and UO_157 (O_157,N_2943,N_2992);
xor UO_158 (O_158,N_2968,N_2942);
and UO_159 (O_159,N_2966,N_2960);
or UO_160 (O_160,N_2996,N_2992);
nor UO_161 (O_161,N_2986,N_2940);
and UO_162 (O_162,N_2974,N_2990);
and UO_163 (O_163,N_2989,N_2976);
xnor UO_164 (O_164,N_2998,N_2969);
or UO_165 (O_165,N_2959,N_2999);
and UO_166 (O_166,N_2945,N_2962);
and UO_167 (O_167,N_2997,N_2955);
nand UO_168 (O_168,N_2991,N_2944);
or UO_169 (O_169,N_2971,N_2951);
or UO_170 (O_170,N_2964,N_2988);
nor UO_171 (O_171,N_2977,N_2982);
nor UO_172 (O_172,N_2998,N_2943);
nand UO_173 (O_173,N_2970,N_2959);
nor UO_174 (O_174,N_2976,N_2953);
and UO_175 (O_175,N_2955,N_2989);
or UO_176 (O_176,N_2959,N_2978);
and UO_177 (O_177,N_2955,N_2988);
nand UO_178 (O_178,N_2971,N_2945);
or UO_179 (O_179,N_2943,N_2980);
or UO_180 (O_180,N_2977,N_2979);
nand UO_181 (O_181,N_2968,N_2969);
or UO_182 (O_182,N_2948,N_2972);
and UO_183 (O_183,N_2976,N_2997);
or UO_184 (O_184,N_2942,N_2981);
nor UO_185 (O_185,N_2972,N_2950);
and UO_186 (O_186,N_2979,N_2946);
or UO_187 (O_187,N_2982,N_2958);
or UO_188 (O_188,N_2959,N_2974);
nor UO_189 (O_189,N_2965,N_2980);
nand UO_190 (O_190,N_2984,N_2989);
or UO_191 (O_191,N_2956,N_2940);
nand UO_192 (O_192,N_2990,N_2987);
nand UO_193 (O_193,N_2946,N_2990);
nor UO_194 (O_194,N_2944,N_2962);
nor UO_195 (O_195,N_2980,N_2981);
nor UO_196 (O_196,N_2966,N_2973);
and UO_197 (O_197,N_2985,N_2991);
and UO_198 (O_198,N_2978,N_2967);
nand UO_199 (O_199,N_2953,N_2946);
or UO_200 (O_200,N_2989,N_2961);
or UO_201 (O_201,N_2981,N_2943);
nor UO_202 (O_202,N_2963,N_2949);
nand UO_203 (O_203,N_2946,N_2999);
and UO_204 (O_204,N_2963,N_2941);
nor UO_205 (O_205,N_2984,N_2946);
nor UO_206 (O_206,N_2963,N_2965);
and UO_207 (O_207,N_2944,N_2981);
nand UO_208 (O_208,N_2967,N_2962);
nand UO_209 (O_209,N_2958,N_2945);
nor UO_210 (O_210,N_2954,N_2970);
nand UO_211 (O_211,N_2970,N_2967);
or UO_212 (O_212,N_2967,N_2973);
and UO_213 (O_213,N_2948,N_2970);
nand UO_214 (O_214,N_2977,N_2989);
nand UO_215 (O_215,N_2991,N_2954);
nor UO_216 (O_216,N_2967,N_2991);
or UO_217 (O_217,N_2963,N_2956);
and UO_218 (O_218,N_2978,N_2941);
nand UO_219 (O_219,N_2961,N_2943);
nand UO_220 (O_220,N_2992,N_2984);
or UO_221 (O_221,N_2952,N_2979);
nor UO_222 (O_222,N_2970,N_2957);
and UO_223 (O_223,N_2970,N_2988);
and UO_224 (O_224,N_2947,N_2949);
nor UO_225 (O_225,N_2966,N_2977);
nor UO_226 (O_226,N_2964,N_2965);
and UO_227 (O_227,N_2988,N_2975);
nor UO_228 (O_228,N_2967,N_2954);
and UO_229 (O_229,N_2947,N_2995);
or UO_230 (O_230,N_2982,N_2955);
or UO_231 (O_231,N_2940,N_2955);
nor UO_232 (O_232,N_2962,N_2974);
nand UO_233 (O_233,N_2940,N_2964);
nand UO_234 (O_234,N_2975,N_2957);
or UO_235 (O_235,N_2988,N_2976);
and UO_236 (O_236,N_2987,N_2999);
nand UO_237 (O_237,N_2989,N_2956);
or UO_238 (O_238,N_2969,N_2991);
and UO_239 (O_239,N_2989,N_2942);
nand UO_240 (O_240,N_2995,N_2967);
or UO_241 (O_241,N_2989,N_2965);
or UO_242 (O_242,N_2962,N_2989);
nand UO_243 (O_243,N_2952,N_2982);
and UO_244 (O_244,N_2991,N_2961);
or UO_245 (O_245,N_2967,N_2956);
nand UO_246 (O_246,N_2963,N_2975);
and UO_247 (O_247,N_2989,N_2953);
nor UO_248 (O_248,N_2967,N_2994);
and UO_249 (O_249,N_2998,N_2975);
and UO_250 (O_250,N_2957,N_2945);
nand UO_251 (O_251,N_2949,N_2972);
or UO_252 (O_252,N_2952,N_2996);
nor UO_253 (O_253,N_2957,N_2982);
and UO_254 (O_254,N_2993,N_2994);
or UO_255 (O_255,N_2947,N_2979);
nand UO_256 (O_256,N_2999,N_2975);
and UO_257 (O_257,N_2984,N_2945);
or UO_258 (O_258,N_2953,N_2944);
nand UO_259 (O_259,N_2954,N_2950);
xor UO_260 (O_260,N_2944,N_2986);
and UO_261 (O_261,N_2972,N_2958);
nand UO_262 (O_262,N_2970,N_2956);
and UO_263 (O_263,N_2976,N_2948);
and UO_264 (O_264,N_2962,N_2979);
and UO_265 (O_265,N_2970,N_2941);
and UO_266 (O_266,N_2989,N_2960);
or UO_267 (O_267,N_2981,N_2984);
nand UO_268 (O_268,N_2973,N_2961);
and UO_269 (O_269,N_2983,N_2997);
or UO_270 (O_270,N_2943,N_2947);
or UO_271 (O_271,N_2946,N_2970);
nand UO_272 (O_272,N_2989,N_2983);
nand UO_273 (O_273,N_2958,N_2979);
and UO_274 (O_274,N_2958,N_2985);
nor UO_275 (O_275,N_2947,N_2967);
nor UO_276 (O_276,N_2967,N_2969);
nand UO_277 (O_277,N_2993,N_2979);
nand UO_278 (O_278,N_2988,N_2952);
nand UO_279 (O_279,N_2982,N_2944);
or UO_280 (O_280,N_2985,N_2990);
nor UO_281 (O_281,N_2979,N_2971);
or UO_282 (O_282,N_2954,N_2978);
or UO_283 (O_283,N_2973,N_2998);
nand UO_284 (O_284,N_2961,N_2993);
and UO_285 (O_285,N_2976,N_2978);
nor UO_286 (O_286,N_2991,N_2993);
or UO_287 (O_287,N_2958,N_2975);
or UO_288 (O_288,N_2955,N_2954);
nor UO_289 (O_289,N_2971,N_2966);
nor UO_290 (O_290,N_2988,N_2954);
or UO_291 (O_291,N_2992,N_2987);
or UO_292 (O_292,N_2950,N_2951);
nor UO_293 (O_293,N_2988,N_2962);
and UO_294 (O_294,N_2992,N_2966);
nand UO_295 (O_295,N_2972,N_2999);
and UO_296 (O_296,N_2974,N_2946);
nor UO_297 (O_297,N_2969,N_2970);
nor UO_298 (O_298,N_2979,N_2973);
nor UO_299 (O_299,N_2941,N_2979);
and UO_300 (O_300,N_2980,N_2957);
or UO_301 (O_301,N_2973,N_2960);
nand UO_302 (O_302,N_2952,N_2994);
nor UO_303 (O_303,N_2982,N_2967);
or UO_304 (O_304,N_2960,N_2979);
or UO_305 (O_305,N_2999,N_2977);
and UO_306 (O_306,N_2961,N_2972);
and UO_307 (O_307,N_2981,N_2995);
nand UO_308 (O_308,N_2951,N_2998);
and UO_309 (O_309,N_2949,N_2961);
or UO_310 (O_310,N_2962,N_2993);
nor UO_311 (O_311,N_2995,N_2992);
nor UO_312 (O_312,N_2940,N_2973);
nand UO_313 (O_313,N_2980,N_2985);
or UO_314 (O_314,N_2956,N_2994);
nor UO_315 (O_315,N_2969,N_2994);
nand UO_316 (O_316,N_2999,N_2956);
nand UO_317 (O_317,N_2984,N_2974);
or UO_318 (O_318,N_2973,N_2963);
nor UO_319 (O_319,N_2983,N_2987);
and UO_320 (O_320,N_2945,N_2964);
nand UO_321 (O_321,N_2999,N_2966);
nor UO_322 (O_322,N_2977,N_2944);
nand UO_323 (O_323,N_2972,N_2952);
nand UO_324 (O_324,N_2990,N_2993);
nand UO_325 (O_325,N_2993,N_2978);
or UO_326 (O_326,N_2956,N_2984);
nand UO_327 (O_327,N_2980,N_2996);
and UO_328 (O_328,N_2986,N_2980);
nor UO_329 (O_329,N_2961,N_2947);
nor UO_330 (O_330,N_2979,N_2961);
and UO_331 (O_331,N_2991,N_2976);
nor UO_332 (O_332,N_2962,N_2975);
nand UO_333 (O_333,N_2967,N_2966);
xor UO_334 (O_334,N_2980,N_2974);
and UO_335 (O_335,N_2969,N_2954);
nor UO_336 (O_336,N_2967,N_2946);
nand UO_337 (O_337,N_2984,N_2994);
nor UO_338 (O_338,N_2982,N_2962);
nor UO_339 (O_339,N_2950,N_2949);
nand UO_340 (O_340,N_2985,N_2957);
nor UO_341 (O_341,N_2944,N_2952);
or UO_342 (O_342,N_2957,N_2956);
or UO_343 (O_343,N_2967,N_2963);
and UO_344 (O_344,N_2974,N_2977);
and UO_345 (O_345,N_2962,N_2959);
and UO_346 (O_346,N_2969,N_2951);
nor UO_347 (O_347,N_2957,N_2996);
or UO_348 (O_348,N_2954,N_2999);
nand UO_349 (O_349,N_2961,N_2970);
nor UO_350 (O_350,N_2958,N_2999);
nor UO_351 (O_351,N_2941,N_2993);
or UO_352 (O_352,N_2972,N_2956);
and UO_353 (O_353,N_2968,N_2991);
and UO_354 (O_354,N_2957,N_2984);
or UO_355 (O_355,N_2974,N_2949);
nand UO_356 (O_356,N_2989,N_2951);
nand UO_357 (O_357,N_2997,N_2975);
nand UO_358 (O_358,N_2973,N_2975);
xnor UO_359 (O_359,N_2959,N_2975);
and UO_360 (O_360,N_2980,N_2987);
nor UO_361 (O_361,N_2972,N_2954);
nor UO_362 (O_362,N_2990,N_2964);
nor UO_363 (O_363,N_2970,N_2942);
nor UO_364 (O_364,N_2994,N_2945);
nor UO_365 (O_365,N_2964,N_2951);
nor UO_366 (O_366,N_2997,N_2981);
nand UO_367 (O_367,N_2957,N_2942);
nand UO_368 (O_368,N_2991,N_2956);
and UO_369 (O_369,N_2993,N_2954);
nand UO_370 (O_370,N_2997,N_2980);
nand UO_371 (O_371,N_2965,N_2975);
nand UO_372 (O_372,N_2982,N_2974);
nor UO_373 (O_373,N_2950,N_2979);
nand UO_374 (O_374,N_2986,N_2951);
nand UO_375 (O_375,N_2996,N_2942);
nand UO_376 (O_376,N_2957,N_2944);
nor UO_377 (O_377,N_2982,N_2968);
nand UO_378 (O_378,N_2992,N_2953);
or UO_379 (O_379,N_2986,N_2983);
or UO_380 (O_380,N_2963,N_2955);
and UO_381 (O_381,N_2964,N_2979);
and UO_382 (O_382,N_2996,N_2988);
nand UO_383 (O_383,N_2965,N_2946);
nor UO_384 (O_384,N_2943,N_2988);
and UO_385 (O_385,N_2948,N_2997);
nand UO_386 (O_386,N_2946,N_2987);
and UO_387 (O_387,N_2965,N_2969);
nand UO_388 (O_388,N_2998,N_2978);
xnor UO_389 (O_389,N_2987,N_2961);
nand UO_390 (O_390,N_2943,N_2999);
or UO_391 (O_391,N_2957,N_2958);
nor UO_392 (O_392,N_2941,N_2945);
nand UO_393 (O_393,N_2945,N_2973);
or UO_394 (O_394,N_2956,N_2971);
nor UO_395 (O_395,N_2988,N_2947);
nand UO_396 (O_396,N_2993,N_2960);
or UO_397 (O_397,N_2985,N_2956);
or UO_398 (O_398,N_2975,N_2969);
nor UO_399 (O_399,N_2976,N_2944);
and UO_400 (O_400,N_2973,N_2965);
or UO_401 (O_401,N_2975,N_2978);
nand UO_402 (O_402,N_2942,N_2951);
or UO_403 (O_403,N_2992,N_2986);
or UO_404 (O_404,N_2949,N_2962);
nor UO_405 (O_405,N_2976,N_2972);
and UO_406 (O_406,N_2955,N_2983);
nand UO_407 (O_407,N_2992,N_2963);
xor UO_408 (O_408,N_2974,N_2951);
xor UO_409 (O_409,N_2982,N_2948);
and UO_410 (O_410,N_2986,N_2985);
nand UO_411 (O_411,N_2948,N_2945);
and UO_412 (O_412,N_2966,N_2948);
nor UO_413 (O_413,N_2994,N_2978);
nor UO_414 (O_414,N_2967,N_2974);
nor UO_415 (O_415,N_2955,N_2991);
nand UO_416 (O_416,N_2956,N_2950);
or UO_417 (O_417,N_2951,N_2965);
nor UO_418 (O_418,N_2979,N_2953);
or UO_419 (O_419,N_2960,N_2994);
nor UO_420 (O_420,N_2973,N_2951);
or UO_421 (O_421,N_2992,N_2952);
nor UO_422 (O_422,N_2986,N_2995);
nor UO_423 (O_423,N_2951,N_2976);
or UO_424 (O_424,N_2963,N_2978);
nand UO_425 (O_425,N_2974,N_2945);
nand UO_426 (O_426,N_2992,N_2950);
nor UO_427 (O_427,N_2951,N_2941);
or UO_428 (O_428,N_2997,N_2967);
or UO_429 (O_429,N_2976,N_2962);
nor UO_430 (O_430,N_2999,N_2983);
xor UO_431 (O_431,N_2967,N_2952);
or UO_432 (O_432,N_2950,N_2959);
nand UO_433 (O_433,N_2957,N_2960);
or UO_434 (O_434,N_2949,N_2976);
nor UO_435 (O_435,N_2992,N_2956);
nor UO_436 (O_436,N_2995,N_2983);
and UO_437 (O_437,N_2995,N_2940);
and UO_438 (O_438,N_2961,N_2944);
nand UO_439 (O_439,N_2984,N_2990);
nor UO_440 (O_440,N_2999,N_2944);
nand UO_441 (O_441,N_2962,N_2973);
nand UO_442 (O_442,N_2999,N_2995);
nand UO_443 (O_443,N_2977,N_2971);
nand UO_444 (O_444,N_2948,N_2977);
or UO_445 (O_445,N_2993,N_2998);
or UO_446 (O_446,N_2961,N_2980);
nand UO_447 (O_447,N_2962,N_2963);
or UO_448 (O_448,N_2965,N_2972);
nor UO_449 (O_449,N_2978,N_2968);
or UO_450 (O_450,N_2977,N_2984);
nand UO_451 (O_451,N_2963,N_2944);
nor UO_452 (O_452,N_2971,N_2976);
nor UO_453 (O_453,N_2968,N_2997);
xnor UO_454 (O_454,N_2968,N_2998);
nor UO_455 (O_455,N_2985,N_2974);
nor UO_456 (O_456,N_2993,N_2977);
nor UO_457 (O_457,N_2957,N_2998);
nand UO_458 (O_458,N_2943,N_2987);
or UO_459 (O_459,N_2951,N_2949);
nor UO_460 (O_460,N_2950,N_2996);
nor UO_461 (O_461,N_2978,N_2999);
or UO_462 (O_462,N_2996,N_2999);
and UO_463 (O_463,N_2993,N_2973);
and UO_464 (O_464,N_2972,N_2940);
nand UO_465 (O_465,N_2949,N_2955);
or UO_466 (O_466,N_2974,N_2960);
nor UO_467 (O_467,N_2965,N_2976);
or UO_468 (O_468,N_2944,N_2996);
nand UO_469 (O_469,N_2976,N_2980);
and UO_470 (O_470,N_2977,N_2992);
nor UO_471 (O_471,N_2982,N_2992);
or UO_472 (O_472,N_2965,N_2958);
nor UO_473 (O_473,N_2958,N_2967);
or UO_474 (O_474,N_2945,N_2995);
and UO_475 (O_475,N_2979,N_2989);
and UO_476 (O_476,N_2985,N_2994);
xnor UO_477 (O_477,N_2982,N_2966);
and UO_478 (O_478,N_2997,N_2966);
nand UO_479 (O_479,N_2975,N_2956);
and UO_480 (O_480,N_2950,N_2997);
nor UO_481 (O_481,N_2954,N_2974);
nand UO_482 (O_482,N_2977,N_2955);
or UO_483 (O_483,N_2971,N_2988);
and UO_484 (O_484,N_2987,N_2969);
nor UO_485 (O_485,N_2949,N_2956);
nor UO_486 (O_486,N_2978,N_2940);
nor UO_487 (O_487,N_2983,N_2993);
nor UO_488 (O_488,N_2963,N_2943);
or UO_489 (O_489,N_2960,N_2969);
nor UO_490 (O_490,N_2955,N_2962);
and UO_491 (O_491,N_2995,N_2960);
or UO_492 (O_492,N_2996,N_2969);
or UO_493 (O_493,N_2955,N_2999);
nor UO_494 (O_494,N_2970,N_2987);
nand UO_495 (O_495,N_2981,N_2959);
or UO_496 (O_496,N_2949,N_2954);
nand UO_497 (O_497,N_2973,N_2955);
nand UO_498 (O_498,N_2989,N_2952);
nand UO_499 (O_499,N_2960,N_2950);
endmodule