module basic_1500_15000_2000_20_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_731,In_1345);
nor U1 (N_1,In_1411,In_1437);
nor U2 (N_2,In_967,In_692);
and U3 (N_3,In_831,In_348);
or U4 (N_4,In_1043,In_479);
or U5 (N_5,In_243,In_1030);
or U6 (N_6,In_105,In_1099);
and U7 (N_7,In_1493,In_388);
nand U8 (N_8,In_879,In_202);
nand U9 (N_9,In_1313,In_598);
and U10 (N_10,In_309,In_401);
or U11 (N_11,In_296,In_442);
and U12 (N_12,In_686,In_1496);
or U13 (N_13,In_872,In_304);
or U14 (N_14,In_1149,In_757);
nor U15 (N_15,In_594,In_158);
and U16 (N_16,In_678,In_88);
and U17 (N_17,In_1179,In_16);
and U18 (N_18,In_1084,In_793);
xnor U19 (N_19,In_885,In_32);
or U20 (N_20,In_179,In_196);
or U21 (N_21,In_980,In_258);
nand U22 (N_22,In_114,In_293);
and U23 (N_23,In_935,In_228);
or U24 (N_24,In_934,In_742);
nor U25 (N_25,In_1405,In_1262);
or U26 (N_26,In_249,In_252);
nand U27 (N_27,In_1451,In_489);
nor U28 (N_28,In_1176,In_1101);
xnor U29 (N_29,In_968,In_393);
nor U30 (N_30,In_103,In_1060);
and U31 (N_31,In_450,In_1337);
nor U32 (N_32,In_505,In_699);
and U33 (N_33,In_406,In_246);
and U34 (N_34,In_303,In_435);
and U35 (N_35,In_1135,In_1174);
nor U36 (N_36,In_705,In_1432);
or U37 (N_37,In_73,In_527);
and U38 (N_38,In_446,In_382);
or U39 (N_39,In_1377,In_353);
and U40 (N_40,In_1242,In_741);
xnor U41 (N_41,In_1421,In_156);
nor U42 (N_42,In_1086,In_493);
nor U43 (N_43,In_1157,In_1353);
and U44 (N_44,In_449,In_1145);
nand U45 (N_45,In_822,In_0);
nor U46 (N_46,In_1087,In_286);
and U47 (N_47,In_1209,In_932);
and U48 (N_48,In_676,In_1239);
or U49 (N_49,In_1093,In_526);
nor U50 (N_50,In_573,In_805);
and U51 (N_51,In_599,In_1418);
and U52 (N_52,In_1105,In_15);
or U53 (N_53,In_1370,In_274);
xor U54 (N_54,In_83,In_1327);
or U55 (N_55,In_1033,In_94);
and U56 (N_56,In_175,In_1058);
nand U57 (N_57,In_365,In_325);
nor U58 (N_58,In_1357,In_56);
nand U59 (N_59,In_796,In_1203);
nand U60 (N_60,In_936,In_421);
xnor U61 (N_61,In_1119,In_71);
or U62 (N_62,In_1277,In_1061);
nor U63 (N_63,In_1276,In_587);
nor U64 (N_64,In_1160,In_643);
or U65 (N_65,In_910,In_864);
nor U66 (N_66,In_404,In_441);
nand U67 (N_67,In_1106,In_1401);
nand U68 (N_68,In_559,In_132);
and U69 (N_69,In_1029,In_278);
or U70 (N_70,In_545,In_627);
or U71 (N_71,In_1005,In_1409);
xnor U72 (N_72,In_419,In_675);
nand U73 (N_73,In_236,In_862);
or U74 (N_74,In_461,In_738);
nand U75 (N_75,In_1325,In_916);
nor U76 (N_76,In_280,In_646);
or U77 (N_77,In_804,In_564);
nand U78 (N_78,In_1380,In_889);
nand U79 (N_79,In_172,In_499);
nand U80 (N_80,In_955,In_305);
or U81 (N_81,In_597,In_844);
and U82 (N_82,In_591,In_1340);
or U83 (N_83,In_1491,In_1143);
nand U84 (N_84,In_883,In_402);
nor U85 (N_85,In_1214,In_900);
or U86 (N_86,In_496,In_877);
and U87 (N_87,In_336,In_355);
and U88 (N_88,In_1110,In_194);
or U89 (N_89,In_223,In_308);
nor U90 (N_90,In_507,In_562);
or U91 (N_91,In_1481,In_552);
xor U92 (N_92,In_1296,In_170);
nor U93 (N_93,In_550,In_63);
or U94 (N_94,In_111,In_436);
nand U95 (N_95,In_1066,In_1260);
xnor U96 (N_96,In_1386,In_451);
xor U97 (N_97,In_238,In_487);
or U98 (N_98,In_306,In_1495);
nand U99 (N_99,In_574,In_612);
nor U100 (N_100,In_560,In_478);
nor U101 (N_101,In_18,In_1037);
nand U102 (N_102,In_1026,In_174);
nand U103 (N_103,In_65,In_1152);
and U104 (N_104,In_1245,In_19);
or U105 (N_105,In_1236,In_1454);
nor U106 (N_106,In_547,In_1131);
and U107 (N_107,In_328,In_1133);
nor U108 (N_108,In_1216,In_1396);
and U109 (N_109,In_971,In_217);
or U110 (N_110,In_1051,In_1235);
nor U111 (N_111,In_231,In_27);
or U112 (N_112,In_1224,In_1080);
and U113 (N_113,In_80,In_645);
and U114 (N_114,In_1137,In_959);
and U115 (N_115,In_390,In_1427);
and U116 (N_116,In_1439,In_33);
nor U117 (N_117,In_1212,In_1150);
nor U118 (N_118,In_531,In_1420);
nor U119 (N_119,In_892,In_21);
nor U120 (N_120,In_1088,In_984);
nor U121 (N_121,In_273,In_1480);
and U122 (N_122,In_210,In_666);
or U123 (N_123,In_1040,In_1343);
or U124 (N_124,In_1126,In_265);
xnor U125 (N_125,In_1197,In_842);
xor U126 (N_126,In_605,In_1445);
nand U127 (N_127,In_1180,In_47);
xor U128 (N_128,In_437,In_679);
or U129 (N_129,In_656,In_1116);
nand U130 (N_130,In_969,In_1103);
nor U131 (N_131,In_242,In_1098);
or U132 (N_132,In_1447,In_1484);
or U133 (N_133,In_1195,In_122);
nand U134 (N_134,In_448,In_974);
nor U135 (N_135,In_193,In_475);
nor U136 (N_136,In_1402,In_424);
nand U137 (N_137,In_1064,In_1003);
and U138 (N_138,In_595,In_964);
or U139 (N_139,In_1263,In_812);
nand U140 (N_140,In_681,In_50);
nand U141 (N_141,In_606,In_1384);
or U142 (N_142,In_1450,In_11);
nand U143 (N_143,In_908,In_1054);
or U144 (N_144,In_259,In_30);
or U145 (N_145,In_937,In_638);
nand U146 (N_146,In_1290,In_965);
and U147 (N_147,In_44,In_747);
nor U148 (N_148,In_669,In_693);
nand U149 (N_149,In_1142,In_1300);
or U150 (N_150,In_896,In_1258);
and U151 (N_151,In_366,In_878);
nand U152 (N_152,In_513,In_703);
xnor U153 (N_153,In_1122,In_387);
or U154 (N_154,In_1494,In_1354);
nand U155 (N_155,In_765,In_331);
or U156 (N_156,In_98,In_1438);
xor U157 (N_157,In_604,In_57);
and U158 (N_158,In_457,In_84);
xnor U159 (N_159,In_136,In_716);
nor U160 (N_160,In_180,In_60);
and U161 (N_161,In_583,In_1165);
nor U162 (N_162,In_1046,In_986);
nor U163 (N_163,In_1,In_691);
nand U164 (N_164,In_38,In_865);
and U165 (N_165,In_25,In_1229);
or U166 (N_166,In_789,In_557);
xor U167 (N_167,In_727,In_233);
nand U168 (N_168,In_503,In_463);
and U169 (N_169,In_302,In_1207);
nand U170 (N_170,In_921,In_232);
nor U171 (N_171,In_609,In_924);
nand U172 (N_172,In_326,In_465);
and U173 (N_173,In_1077,In_1463);
nor U174 (N_174,In_758,In_1331);
and U175 (N_175,In_1213,In_641);
and U176 (N_176,In_1299,In_241);
nand U177 (N_177,In_400,In_1237);
or U178 (N_178,In_1347,In_754);
xor U179 (N_179,In_225,In_1226);
or U180 (N_180,In_1342,In_584);
or U181 (N_181,In_1014,In_1458);
nor U182 (N_182,In_119,In_1139);
and U183 (N_183,In_1204,In_1415);
nor U184 (N_184,In_1464,In_329);
or U185 (N_185,In_672,In_1023);
nor U186 (N_186,In_288,In_814);
nor U187 (N_187,In_459,In_87);
nor U188 (N_188,In_795,In_702);
and U189 (N_189,In_45,In_632);
or U190 (N_190,In_929,In_130);
nor U191 (N_191,In_1189,In_426);
or U192 (N_192,In_1311,In_820);
or U193 (N_193,In_700,In_1388);
or U194 (N_194,In_784,In_626);
and U195 (N_195,In_311,In_10);
nor U196 (N_196,In_1293,In_1163);
nor U197 (N_197,In_358,In_785);
and U198 (N_198,In_282,In_905);
nor U199 (N_199,In_1444,In_644);
or U200 (N_200,In_1468,In_1292);
and U201 (N_201,In_131,In_96);
nand U202 (N_202,In_1446,In_650);
or U203 (N_203,In_1035,In_420);
or U204 (N_204,In_815,In_659);
nand U205 (N_205,In_698,In_472);
or U206 (N_206,In_100,In_943);
or U207 (N_207,In_704,In_1315);
and U208 (N_208,In_277,In_655);
or U209 (N_209,In_827,In_124);
nor U210 (N_210,In_951,In_1136);
xnor U211 (N_211,In_1452,In_1309);
nor U212 (N_212,In_786,In_1348);
and U213 (N_213,In_657,In_596);
nor U214 (N_214,In_1358,In_1368);
nor U215 (N_215,In_529,In_256);
xnor U216 (N_216,In_77,In_567);
and U217 (N_217,In_760,In_417);
nor U218 (N_218,In_778,In_690);
nor U219 (N_219,In_1413,In_1089);
xnor U220 (N_220,In_1465,In_1238);
nor U221 (N_221,In_1183,In_380);
or U222 (N_222,In_116,In_852);
or U223 (N_223,In_82,In_729);
xor U224 (N_224,In_1498,In_590);
nor U225 (N_225,In_76,In_761);
nor U226 (N_226,In_588,In_1114);
nor U227 (N_227,In_1120,In_226);
or U228 (N_228,In_517,In_37);
nor U229 (N_229,In_722,In_1312);
nor U230 (N_230,In_349,In_1164);
nor U231 (N_231,In_295,In_950);
nor U232 (N_232,In_1367,In_1278);
or U233 (N_233,In_845,In_269);
or U234 (N_234,In_1349,In_482);
and U235 (N_235,In_1021,In_835);
and U236 (N_236,In_664,In_147);
and U237 (N_237,In_49,In_537);
nor U238 (N_238,In_1194,In_1341);
nor U239 (N_239,In_1457,In_1059);
nor U240 (N_240,In_312,In_1400);
nand U241 (N_241,In_931,In_1271);
and U242 (N_242,In_928,In_1250);
and U243 (N_243,In_565,In_887);
or U244 (N_244,In_1109,In_530);
nand U245 (N_245,In_620,In_140);
nor U246 (N_246,In_1156,In_294);
nand U247 (N_247,In_474,In_121);
nand U248 (N_248,In_995,In_771);
and U249 (N_249,In_70,In_40);
nor U250 (N_250,In_1082,In_536);
or U251 (N_251,In_1094,In_405);
nand U252 (N_252,In_1019,In_1339);
xor U253 (N_253,In_637,In_1108);
or U254 (N_254,In_317,In_1208);
nor U255 (N_255,In_99,In_1070);
or U256 (N_256,In_764,In_846);
nor U257 (N_257,In_711,In_1241);
and U258 (N_258,In_185,In_1173);
nor U259 (N_259,In_821,In_586);
nand U260 (N_260,In_720,In_385);
xnor U261 (N_261,In_839,In_989);
or U262 (N_262,In_807,In_790);
nand U263 (N_263,In_1147,In_894);
nand U264 (N_264,In_432,In_724);
nand U265 (N_265,In_263,In_1346);
or U266 (N_266,In_1243,In_79);
or U267 (N_267,In_93,In_123);
and U268 (N_268,In_756,In_851);
xor U269 (N_269,In_797,In_854);
and U270 (N_270,In_991,In_1172);
or U271 (N_271,In_1305,In_1166);
and U272 (N_272,In_628,In_918);
and U273 (N_273,In_445,In_135);
xor U274 (N_274,In_1366,In_1344);
or U275 (N_275,In_1291,In_1187);
or U276 (N_276,In_1304,In_524);
nor U277 (N_277,In_579,In_203);
and U278 (N_278,In_344,In_922);
or U279 (N_279,In_95,In_1141);
nand U280 (N_280,In_701,In_662);
or U281 (N_281,In_652,In_1097);
xor U282 (N_282,In_204,In_268);
nand U283 (N_283,In_625,In_149);
and U284 (N_284,In_395,In_687);
xnor U285 (N_285,In_1459,In_48);
nand U286 (N_286,In_377,In_642);
nand U287 (N_287,In_1298,In_602);
or U288 (N_288,In_391,In_1048);
or U289 (N_289,In_213,In_81);
and U290 (N_290,In_403,In_746);
nor U291 (N_291,In_1443,In_1478);
and U292 (N_292,In_1379,In_696);
and U293 (N_293,In_621,In_818);
nor U294 (N_294,In_281,In_987);
xor U295 (N_295,In_890,In_1310);
and U296 (N_296,In_1319,In_381);
nor U297 (N_297,In_211,In_1230);
or U298 (N_298,In_1350,In_413);
and U299 (N_299,In_585,In_1081);
and U300 (N_300,In_162,In_471);
nand U301 (N_301,In_271,In_600);
nand U302 (N_302,In_1448,In_763);
nor U303 (N_303,In_544,In_773);
or U304 (N_304,In_975,In_1113);
nand U305 (N_305,In_1270,In_1148);
nor U306 (N_306,In_1466,In_873);
xor U307 (N_307,In_1057,In_607);
nand U308 (N_308,In_1028,In_1261);
nand U309 (N_309,In_1361,In_480);
nand U310 (N_310,In_1359,In_428);
or U311 (N_311,In_200,In_398);
and U312 (N_312,In_1118,In_867);
or U313 (N_313,In_292,In_118);
or U314 (N_314,In_164,In_748);
nor U315 (N_315,In_433,In_423);
xnor U316 (N_316,In_26,In_992);
nand U317 (N_317,In_1085,In_399);
nand U318 (N_318,In_553,In_1107);
nor U319 (N_319,In_35,In_775);
or U320 (N_320,In_911,In_1267);
nand U321 (N_321,In_613,In_1419);
or U322 (N_322,In_187,In_825);
nand U323 (N_323,In_234,In_1482);
nand U324 (N_324,In_1025,In_272);
nand U325 (N_325,In_1006,In_1159);
xor U326 (N_326,In_51,In_551);
nor U327 (N_327,In_712,In_580);
or U328 (N_328,In_333,In_221);
xor U329 (N_329,In_1416,In_1100);
nor U330 (N_330,In_376,In_212);
nor U331 (N_331,In_572,In_1111);
and U332 (N_332,In_285,In_1470);
and U333 (N_333,In_569,In_1475);
xnor U334 (N_334,In_346,In_714);
or U335 (N_335,In_1158,In_466);
nand U336 (N_336,In_1042,In_410);
or U337 (N_337,In_1497,In_1000);
or U338 (N_338,In_339,In_514);
nor U339 (N_339,In_337,In_257);
nor U340 (N_340,In_1186,In_332);
nand U341 (N_341,In_1456,In_184);
xor U342 (N_342,In_1335,In_829);
and U343 (N_343,In_1041,In_1168);
nor U344 (N_344,In_321,In_1363);
and U345 (N_345,In_817,In_868);
nand U346 (N_346,In_653,In_237);
or U347 (N_347,In_735,In_1499);
nand U348 (N_348,In_1013,In_427);
nor U349 (N_349,In_725,In_155);
or U350 (N_350,In_338,In_1422);
or U351 (N_351,In_504,In_143);
nand U352 (N_352,In_1223,In_1220);
nand U353 (N_353,In_780,In_484);
and U354 (N_354,In_36,In_1073);
xnor U355 (N_355,In_141,In_276);
nor U356 (N_356,In_31,In_622);
xor U357 (N_357,In_72,In_849);
nand U358 (N_358,In_876,In_1273);
or U359 (N_359,In_619,In_651);
xor U360 (N_360,In_614,In_126);
and U361 (N_361,In_1016,In_859);
and U362 (N_362,In_1193,In_1074);
or U363 (N_363,In_1425,In_709);
nor U364 (N_364,In_299,In_138);
nand U365 (N_365,In_1407,In_481);
xnor U366 (N_366,In_743,In_841);
nand U367 (N_367,In_133,In_161);
nor U368 (N_368,In_654,In_880);
and U369 (N_369,In_1002,In_145);
or U370 (N_370,In_1130,In_561);
and U371 (N_371,In_89,In_1264);
nand U372 (N_372,In_630,In_850);
nor U373 (N_373,In_582,In_1124);
nand U374 (N_374,In_1417,In_1069);
and U375 (N_375,In_518,In_342);
nor U376 (N_376,In_1206,In_1155);
nor U377 (N_377,In_1306,In_830);
nand U378 (N_378,In_1112,In_1217);
nor U379 (N_379,In_159,In_1198);
or U380 (N_380,In_69,In_958);
nand U381 (N_381,In_216,In_1175);
nor U382 (N_382,In_127,In_978);
or U383 (N_383,In_1001,In_335);
and U384 (N_384,In_753,In_781);
or U385 (N_385,In_1225,In_546);
nor U386 (N_386,In_881,In_893);
or U387 (N_387,In_1065,In_1177);
nand U388 (N_388,In_636,In_1265);
or U389 (N_389,In_1392,In_688);
nand U390 (N_390,In_368,In_352);
and U391 (N_391,In_949,In_534);
and U392 (N_392,In_109,In_1397);
and U393 (N_393,In_334,In_1430);
xnor U394 (N_394,In_1259,In_994);
or U395 (N_395,In_1490,In_363);
nor U396 (N_396,In_799,In_521);
nor U397 (N_397,In_22,In_1492);
xor U398 (N_398,In_255,In_146);
nand U399 (N_399,In_491,In_1044);
nand U400 (N_400,In_152,In_188);
nand U401 (N_401,In_362,In_1391);
and U402 (N_402,In_1284,In_575);
xor U403 (N_403,In_168,In_1389);
nor U404 (N_404,In_68,In_832);
or U405 (N_405,In_697,In_895);
or U406 (N_406,In_1153,In_719);
or U407 (N_407,In_52,In_64);
nor U408 (N_408,In_1125,In_813);
and U409 (N_409,In_372,In_708);
nand U410 (N_410,In_74,In_5);
or U411 (N_411,In_307,In_1127);
and U412 (N_412,In_739,In_1485);
and U413 (N_413,In_199,In_1154);
or U414 (N_414,In_1280,In_106);
nand U415 (N_415,In_422,In_195);
and U416 (N_416,In_840,In_904);
nand U417 (N_417,In_374,In_902);
nor U418 (N_418,In_41,In_1072);
nand U419 (N_419,In_1171,In_440);
or U420 (N_420,In_1062,In_235);
nor U421 (N_421,In_1390,In_201);
or U422 (N_422,In_1301,In_150);
nand U423 (N_423,In_919,In_1134);
or U424 (N_424,In_438,In_139);
nand U425 (N_425,In_665,In_1329);
and U426 (N_426,In_717,In_1322);
xnor U427 (N_427,In_1063,In_909);
nor U428 (N_428,In_112,In_251);
and U429 (N_429,In_838,In_540);
and U430 (N_430,In_824,In_1075);
or U431 (N_431,In_137,In_1287);
nor U432 (N_432,In_1162,In_601);
or U433 (N_433,In_668,In_176);
nand U434 (N_434,In_898,In_884);
and U435 (N_435,In_874,In_800);
nand U436 (N_436,In_260,In_189);
or U437 (N_437,In_624,In_454);
xnor U438 (N_438,In_749,In_254);
nand U439 (N_439,In_319,In_1205);
and U440 (N_440,In_367,In_576);
xnor U441 (N_441,In_1055,In_915);
xnor U442 (N_442,In_721,In_882);
and U443 (N_443,In_1442,In_791);
or U444 (N_444,In_954,In_1039);
nand U445 (N_445,In_327,In_283);
and U446 (N_446,In_1371,In_733);
or U447 (N_447,In_85,In_1104);
nor U448 (N_448,In_12,In_97);
nor U449 (N_449,In_740,In_245);
nand U450 (N_450,In_826,In_858);
or U451 (N_451,In_1404,In_855);
nor U452 (N_452,In_1351,In_737);
xnor U453 (N_453,In_819,In_1394);
or U454 (N_454,In_930,In_1102);
and U455 (N_455,In_1308,In_750);
nor U456 (N_456,In_250,In_856);
nand U457 (N_457,In_1281,In_660);
and U458 (N_458,In_1201,In_680);
and U459 (N_459,In_1027,In_983);
or U460 (N_460,In_460,In_1373);
and U461 (N_461,In_439,In_485);
xor U462 (N_462,In_1288,In_1004);
nor U463 (N_463,In_512,In_962);
and U464 (N_464,In_1285,In_1431);
or U465 (N_465,In_171,In_1095);
nand U466 (N_466,In_62,In_3);
and U467 (N_467,In_767,In_1071);
nor U468 (N_468,In_608,In_347);
or U469 (N_469,In_1477,In_616);
nand U470 (N_470,In_1406,In_86);
nor U471 (N_471,In_506,In_107);
nor U472 (N_472,In_418,In_120);
xor U473 (N_473,In_181,In_1476);
nand U474 (N_474,In_431,In_798);
nor U475 (N_475,In_494,In_787);
and U476 (N_476,In_532,In_458);
and U477 (N_477,In_90,In_836);
nor U478 (N_478,In_811,In_270);
and U479 (N_479,In_926,In_356);
or U480 (N_480,In_34,In_316);
xor U481 (N_481,In_988,In_301);
nand U482 (N_482,In_407,In_59);
or U483 (N_483,In_1252,In_945);
or U484 (N_484,In_1453,In_1123);
xnor U485 (N_485,In_520,In_1289);
xor U486 (N_486,In_755,In_808);
or U487 (N_487,In_566,In_554);
or U488 (N_488,In_728,In_351);
xnor U489 (N_489,In_209,In_244);
nor U490 (N_490,In_997,In_154);
and U491 (N_491,In_1188,In_324);
and U492 (N_492,In_519,In_1483);
and U493 (N_493,In_990,In_266);
or U494 (N_494,In_548,In_1018);
nor U495 (N_495,In_134,In_555);
and U496 (N_496,In_870,In_1269);
nand U497 (N_497,In_973,In_415);
or U498 (N_498,In_942,In_917);
nor U499 (N_499,In_1316,In_823);
nand U500 (N_500,In_383,In_1032);
nand U501 (N_501,In_1469,In_730);
nand U502 (N_502,In_713,In_1294);
and U503 (N_503,In_1428,In_13);
or U504 (N_504,In_1362,In_345);
nand U505 (N_505,In_803,In_46);
and U506 (N_506,In_1050,In_695);
and U507 (N_507,In_67,In_1246);
xor U508 (N_508,In_674,In_571);
nor U509 (N_509,In_558,In_1471);
or U510 (N_510,In_470,In_1011);
or U511 (N_511,In_745,In_425);
xnor U512 (N_512,In_538,In_901);
and U513 (N_513,In_501,In_220);
nor U514 (N_514,In_914,In_1372);
nand U515 (N_515,In_92,In_177);
and U516 (N_516,In_952,In_1079);
and U517 (N_517,In_774,In_291);
nand U518 (N_518,In_1192,In_933);
and U519 (N_519,In_768,In_707);
or U520 (N_520,In_783,In_43);
nor U521 (N_521,In_375,In_1283);
and U522 (N_522,In_1017,In_208);
or U523 (N_523,In_469,In_456);
nor U524 (N_524,In_455,In_615);
and U525 (N_525,In_888,In_1196);
nor U526 (N_526,In_24,In_1317);
or U527 (N_527,In_224,In_972);
nand U528 (N_528,In_341,In_411);
nor U529 (N_529,In_611,In_267);
nor U530 (N_530,In_618,In_1360);
nor U531 (N_531,In_563,In_279);
nor U532 (N_532,In_183,In_770);
and U533 (N_533,In_810,In_219);
and U534 (N_534,In_963,In_1254);
nand U535 (N_535,In_631,In_1015);
and U536 (N_536,In_1047,In_766);
or U537 (N_537,In_14,In_1248);
or U538 (N_538,In_364,In_1295);
and U539 (N_539,In_163,In_542);
nand U540 (N_540,In_160,In_1240);
nand U541 (N_541,In_1211,In_290);
or U542 (N_542,In_927,In_734);
nand U543 (N_543,In_359,In_861);
nor U544 (N_544,In_104,In_314);
and U545 (N_545,In_360,In_42);
nand U546 (N_546,In_1474,In_1433);
nor U547 (N_547,In_369,In_169);
nor U548 (N_548,In_1251,In_1024);
nand U549 (N_549,In_677,In_453);
or U550 (N_550,In_744,In_1410);
nor U551 (N_551,In_511,In_833);
xnor U552 (N_552,In_129,In_1191);
and U553 (N_553,In_8,In_502);
xnor U554 (N_554,In_192,In_1436);
nor U555 (N_555,In_1128,In_1320);
nand U556 (N_556,In_912,In_523);
nand U557 (N_557,In_947,In_222);
and U558 (N_558,In_1129,In_323);
and U559 (N_559,In_938,In_1247);
and U560 (N_560,In_685,In_1231);
or U561 (N_561,In_1314,In_1382);
and U562 (N_562,In_802,In_871);
and U563 (N_563,In_452,In_1423);
nor U564 (N_564,In_907,In_186);
nor U565 (N_565,In_467,In_948);
nor U566 (N_566,In_1096,In_1184);
nor U567 (N_567,In_396,In_1479);
nand U568 (N_568,In_148,In_1009);
xor U569 (N_569,In_647,In_1324);
and U570 (N_570,In_2,In_197);
nand U571 (N_571,In_214,In_1441);
nor U572 (N_572,In_957,In_847);
and U573 (N_573,In_1414,In_239);
nor U574 (N_574,In_1334,In_541);
nand U575 (N_575,In_115,In_1227);
nor U576 (N_576,In_476,In_142);
or U577 (N_577,In_1031,In_999);
xor U578 (N_578,In_1092,In_165);
nor U579 (N_579,In_970,In_1266);
nor U580 (N_580,In_492,In_167);
and U581 (N_581,In_777,In_1228);
or U582 (N_582,In_752,In_639);
xnor U583 (N_583,In_287,In_1034);
nand U584 (N_584,In_1012,In_1253);
xor U585 (N_585,In_218,In_1302);
and U586 (N_586,In_1488,In_1369);
and U587 (N_587,In_1144,In_54);
or U588 (N_588,In_429,In_515);
or U589 (N_589,In_102,In_977);
nand U590 (N_590,In_151,In_956);
nor U591 (N_591,In_1233,In_539);
nand U592 (N_592,In_801,In_516);
nor U593 (N_593,In_772,In_1338);
and U594 (N_594,In_198,In_1045);
nor U595 (N_595,In_473,In_117);
or U596 (N_596,In_298,In_284);
nor U597 (N_597,In_1170,In_75);
nand U598 (N_598,In_673,In_173);
nor U599 (N_599,In_718,In_1232);
nor U600 (N_600,In_592,In_1356);
or U601 (N_601,In_939,In_1375);
nor U602 (N_602,In_1091,In_1036);
and U603 (N_603,In_6,In_866);
or U604 (N_604,In_1282,In_617);
nor U605 (N_605,In_649,In_769);
nor U606 (N_606,In_330,In_409);
and U607 (N_607,In_1330,In_350);
nand U608 (N_608,In_414,In_488);
or U609 (N_609,In_663,In_1210);
nor U610 (N_610,In_1374,In_125);
or U611 (N_611,In_510,In_386);
nor U612 (N_612,In_101,In_373);
or U613 (N_613,In_925,In_603);
and U614 (N_614,In_1352,In_1083);
nor U615 (N_615,In_343,In_806);
nor U616 (N_616,In_941,In_1222);
nand U617 (N_617,In_998,In_227);
and U618 (N_618,In_379,In_389);
nor U619 (N_619,In_1395,In_961);
or U620 (N_620,In_78,In_736);
nor U621 (N_621,In_1321,In_464);
xor U622 (N_622,In_178,In_166);
and U623 (N_623,In_495,In_670);
nand U624 (N_624,In_834,In_1383);
or U625 (N_625,In_710,In_853);
xor U626 (N_626,In_683,In_1332);
and U627 (N_627,In_1181,In_1318);
or U628 (N_628,In_1146,In_4);
nor U629 (N_629,In_1182,In_863);
nand U630 (N_630,In_667,In_658);
nand U631 (N_631,In_378,In_1117);
or U632 (N_632,In_1333,In_1167);
nor U633 (N_633,In_1326,In_726);
and U634 (N_634,In_715,In_497);
nand U635 (N_635,In_508,In_897);
and U636 (N_636,In_623,In_1132);
nor U637 (N_637,In_1472,In_1020);
xnor U638 (N_638,In_944,In_58);
xor U639 (N_639,In_1178,In_361);
or U640 (N_640,In_732,In_1249);
or U641 (N_641,In_300,In_1076);
nand U642 (N_642,In_310,In_1440);
nand U643 (N_643,In_477,In_1138);
nand U644 (N_644,In_490,In_1190);
and U645 (N_645,In_253,In_394);
or U646 (N_646,In_1218,In_447);
and U647 (N_647,In_776,In_275);
nor U648 (N_648,In_751,In_430);
and U649 (N_649,In_1008,In_1489);
and U650 (N_650,In_581,In_1403);
or U651 (N_651,In_723,In_468);
xor U652 (N_652,In_1215,In_1387);
and U653 (N_653,In_1473,In_205);
and U654 (N_654,In_1049,In_9);
or U655 (N_655,In_190,In_1408);
nor U656 (N_656,In_1467,In_29);
and U657 (N_657,In_416,In_976);
nor U658 (N_658,In_1393,In_891);
and U659 (N_659,In_1255,In_1381);
nand U660 (N_660,In_313,In_1376);
nor U661 (N_661,In_207,In_1199);
or U662 (N_662,In_543,In_913);
and U663 (N_663,In_91,In_706);
or U664 (N_664,In_1219,In_634);
and U665 (N_665,In_1256,In_108);
or U666 (N_666,In_953,In_20);
xor U667 (N_667,In_661,In_843);
and U668 (N_668,In_7,In_483);
and U669 (N_669,In_689,In_1221);
nor U670 (N_670,In_1275,In_1010);
nand U671 (N_671,In_899,In_857);
nor U672 (N_672,In_788,In_792);
nor U673 (N_673,In_1328,In_1202);
nor U674 (N_674,In_206,In_966);
xor U675 (N_675,In_434,In_1234);
and U676 (N_676,In_875,In_297);
nand U677 (N_677,In_860,In_1455);
nand U678 (N_678,In_610,In_392);
nand U679 (N_679,In_229,In_809);
nor U680 (N_680,In_248,In_869);
nor U681 (N_681,In_1412,In_1434);
nand U682 (N_682,In_577,In_1272);
nor U683 (N_683,In_322,In_1424);
xor U684 (N_684,In_960,In_589);
xor U685 (N_685,In_906,In_837);
nor U686 (N_686,In_1151,In_1185);
nor U687 (N_687,In_264,In_1365);
xnor U688 (N_688,In_1268,In_629);
and U689 (N_689,In_535,In_128);
nor U690 (N_690,In_318,In_215);
nand U691 (N_691,In_1378,In_1462);
xor U692 (N_692,In_39,In_886);
nand U693 (N_693,In_357,In_55);
and U694 (N_694,In_1355,In_549);
and U695 (N_695,In_1121,In_979);
or U696 (N_696,In_1486,In_828);
or U697 (N_697,In_633,In_1398);
or U698 (N_698,In_1429,In_1449);
or U699 (N_699,In_1244,In_635);
nor U700 (N_700,In_1385,In_153);
nor U701 (N_701,In_779,In_578);
nor U702 (N_702,In_500,In_412);
or U703 (N_703,In_443,In_408);
nand U704 (N_704,In_157,In_1364);
and U705 (N_705,In_1169,In_996);
and U706 (N_706,In_247,In_671);
nand U707 (N_707,In_191,In_993);
nor U708 (N_708,In_320,In_384);
nor U709 (N_709,In_354,In_1286);
and U710 (N_710,In_1274,In_230);
nand U711 (N_711,In_759,In_262);
nor U712 (N_712,In_648,In_1460);
or U713 (N_713,In_1307,In_522);
xnor U714 (N_714,In_920,In_240);
nand U715 (N_715,In_1426,In_1068);
and U716 (N_716,In_462,In_509);
nand U717 (N_717,In_1461,In_946);
and U718 (N_718,In_1038,In_182);
nor U719 (N_719,In_486,In_1007);
nor U720 (N_720,In_568,In_1279);
xor U721 (N_721,In_556,In_144);
nand U722 (N_722,In_444,In_1487);
or U723 (N_723,In_1022,In_340);
nand U724 (N_724,In_782,In_370);
or U725 (N_725,In_1140,In_794);
nand U726 (N_726,In_528,In_762);
nand U727 (N_727,In_1303,In_1435);
and U728 (N_728,In_1052,In_498);
xor U729 (N_729,In_940,In_684);
and U730 (N_730,In_682,In_1323);
nor U731 (N_731,In_1297,In_315);
nand U732 (N_732,In_1200,In_110);
nor U733 (N_733,In_1056,In_694);
or U734 (N_734,In_816,In_640);
nand U735 (N_735,In_261,In_113);
or U736 (N_736,In_1257,In_23);
and U737 (N_737,In_1078,In_903);
nor U738 (N_738,In_525,In_17);
nand U739 (N_739,In_1053,In_371);
and U740 (N_740,In_923,In_289);
nand U741 (N_741,In_397,In_53);
and U742 (N_742,In_533,In_981);
nor U743 (N_743,In_1161,In_570);
and U744 (N_744,In_1090,In_1115);
xor U745 (N_745,In_593,In_848);
and U746 (N_746,In_985,In_1399);
or U747 (N_747,In_1336,In_61);
nand U748 (N_748,In_66,In_28);
nor U749 (N_749,In_982,In_1067);
nor U750 (N_750,N_526,N_597);
nand U751 (N_751,N_222,N_480);
or U752 (N_752,N_400,N_633);
xor U753 (N_753,N_225,N_657);
xnor U754 (N_754,N_483,N_94);
nand U755 (N_755,N_116,N_583);
nor U756 (N_756,N_245,N_180);
xnor U757 (N_757,N_614,N_652);
nand U758 (N_758,N_326,N_739);
nand U759 (N_759,N_206,N_64);
or U760 (N_760,N_332,N_691);
nor U761 (N_761,N_638,N_260);
nor U762 (N_762,N_512,N_320);
or U763 (N_763,N_204,N_52);
and U764 (N_764,N_661,N_357);
nor U765 (N_765,N_519,N_188);
and U766 (N_766,N_634,N_108);
and U767 (N_767,N_12,N_574);
nand U768 (N_768,N_655,N_598);
xnor U769 (N_769,N_544,N_256);
or U770 (N_770,N_77,N_61);
xor U771 (N_771,N_187,N_138);
and U772 (N_772,N_417,N_669);
or U773 (N_773,N_28,N_572);
or U774 (N_774,N_586,N_700);
nand U775 (N_775,N_342,N_438);
or U776 (N_776,N_447,N_131);
nand U777 (N_777,N_113,N_535);
nor U778 (N_778,N_653,N_365);
nand U779 (N_779,N_484,N_459);
or U780 (N_780,N_334,N_428);
xor U781 (N_781,N_209,N_271);
nand U782 (N_782,N_153,N_121);
or U783 (N_783,N_193,N_749);
or U784 (N_784,N_608,N_470);
nor U785 (N_785,N_278,N_289);
nand U786 (N_786,N_127,N_549);
nor U787 (N_787,N_377,N_217);
or U788 (N_788,N_62,N_716);
nand U789 (N_789,N_261,N_59);
nor U790 (N_790,N_185,N_351);
nor U791 (N_791,N_635,N_38);
nor U792 (N_792,N_407,N_86);
or U793 (N_793,N_154,N_314);
and U794 (N_794,N_439,N_730);
and U795 (N_795,N_493,N_585);
nor U796 (N_796,N_132,N_75);
nor U797 (N_797,N_522,N_704);
xor U798 (N_798,N_117,N_577);
nor U799 (N_799,N_631,N_401);
nor U800 (N_800,N_403,N_368);
nand U801 (N_801,N_211,N_137);
and U802 (N_802,N_324,N_595);
or U803 (N_803,N_167,N_507);
or U804 (N_804,N_4,N_197);
and U805 (N_805,N_238,N_318);
nor U806 (N_806,N_190,N_729);
or U807 (N_807,N_110,N_710);
and U808 (N_808,N_160,N_444);
or U809 (N_809,N_236,N_562);
nor U810 (N_810,N_199,N_745);
and U811 (N_811,N_63,N_664);
or U812 (N_812,N_252,N_191);
nor U813 (N_813,N_701,N_429);
nor U814 (N_814,N_450,N_508);
or U815 (N_815,N_44,N_24);
nor U816 (N_816,N_492,N_541);
or U817 (N_817,N_99,N_6);
and U818 (N_818,N_605,N_57);
nand U819 (N_819,N_668,N_150);
or U820 (N_820,N_590,N_727);
nand U821 (N_821,N_213,N_416);
and U822 (N_822,N_443,N_556);
nor U823 (N_823,N_321,N_528);
nand U824 (N_824,N_481,N_542);
xnor U825 (N_825,N_354,N_465);
nor U826 (N_826,N_19,N_128);
nor U827 (N_827,N_269,N_221);
or U828 (N_828,N_589,N_37);
nand U829 (N_829,N_249,N_624);
nand U830 (N_830,N_3,N_630);
nand U831 (N_831,N_587,N_262);
or U832 (N_832,N_69,N_546);
and U833 (N_833,N_346,N_699);
and U834 (N_834,N_246,N_208);
or U835 (N_835,N_7,N_425);
or U836 (N_836,N_309,N_731);
or U837 (N_837,N_550,N_472);
or U838 (N_838,N_126,N_297);
or U839 (N_839,N_679,N_579);
or U840 (N_840,N_65,N_384);
or U841 (N_841,N_287,N_461);
nand U842 (N_842,N_97,N_596);
nand U843 (N_843,N_448,N_473);
and U844 (N_844,N_503,N_290);
and U845 (N_845,N_305,N_692);
xnor U846 (N_846,N_125,N_445);
nand U847 (N_847,N_270,N_47);
or U848 (N_848,N_383,N_717);
and U849 (N_849,N_647,N_14);
nor U850 (N_850,N_176,N_42);
and U851 (N_851,N_74,N_198);
or U852 (N_852,N_659,N_494);
or U853 (N_853,N_561,N_628);
nor U854 (N_854,N_708,N_87);
and U855 (N_855,N_665,N_226);
or U856 (N_856,N_747,N_141);
nor U857 (N_857,N_501,N_538);
nand U858 (N_858,N_228,N_607);
xor U859 (N_859,N_98,N_422);
nand U860 (N_860,N_32,N_404);
nor U861 (N_861,N_694,N_636);
and U862 (N_862,N_709,N_353);
nand U863 (N_863,N_142,N_268);
nand U864 (N_864,N_205,N_402);
and U865 (N_865,N_328,N_558);
nor U866 (N_866,N_366,N_722);
nor U867 (N_867,N_105,N_220);
or U868 (N_868,N_548,N_148);
nor U869 (N_869,N_591,N_442);
nor U870 (N_870,N_489,N_70);
and U871 (N_871,N_54,N_158);
nor U872 (N_872,N_742,N_695);
or U873 (N_873,N_467,N_129);
and U874 (N_874,N_606,N_291);
nand U875 (N_875,N_723,N_398);
xor U876 (N_876,N_456,N_705);
or U877 (N_877,N_564,N_499);
nand U878 (N_878,N_39,N_109);
or U879 (N_879,N_323,N_335);
nor U880 (N_880,N_517,N_413);
nand U881 (N_881,N_551,N_49);
nor U882 (N_882,N_660,N_688);
xnor U883 (N_883,N_666,N_455);
nand U884 (N_884,N_474,N_168);
xor U885 (N_885,N_234,N_683);
or U886 (N_886,N_48,N_458);
or U887 (N_887,N_740,N_582);
or U888 (N_888,N_50,N_139);
and U889 (N_889,N_92,N_285);
nand U890 (N_890,N_124,N_725);
and U891 (N_891,N_672,N_183);
nand U892 (N_892,N_331,N_609);
nand U893 (N_893,N_468,N_449);
or U894 (N_894,N_229,N_9);
nor U895 (N_895,N_136,N_737);
or U896 (N_896,N_391,N_495);
nand U897 (N_897,N_122,N_223);
nand U898 (N_898,N_414,N_242);
nand U899 (N_899,N_280,N_68);
and U900 (N_900,N_721,N_560);
nand U901 (N_901,N_84,N_409);
xnor U902 (N_902,N_35,N_741);
nand U903 (N_903,N_179,N_103);
nand U904 (N_904,N_106,N_703);
or U905 (N_905,N_490,N_239);
and U906 (N_906,N_81,N_163);
or U907 (N_907,N_534,N_567);
nor U908 (N_908,N_27,N_311);
and U909 (N_909,N_622,N_184);
nor U910 (N_910,N_568,N_247);
and U911 (N_911,N_543,N_15);
nand U912 (N_912,N_374,N_362);
nor U913 (N_913,N_5,N_319);
nand U914 (N_914,N_540,N_257);
nor U915 (N_915,N_639,N_552);
xnor U916 (N_916,N_157,N_389);
or U917 (N_917,N_482,N_10);
xnor U918 (N_918,N_244,N_649);
or U919 (N_919,N_658,N_79);
or U920 (N_920,N_675,N_82);
nor U921 (N_921,N_378,N_565);
nand U922 (N_922,N_315,N_284);
nand U923 (N_923,N_663,N_258);
and U924 (N_924,N_2,N_527);
xor U925 (N_925,N_189,N_533);
nand U926 (N_926,N_671,N_76);
nand U927 (N_927,N_553,N_619);
nor U928 (N_928,N_302,N_181);
nand U929 (N_929,N_689,N_524);
nand U930 (N_930,N_186,N_557);
nor U931 (N_931,N_580,N_301);
nand U932 (N_932,N_408,N_724);
nand U933 (N_933,N_73,N_118);
and U934 (N_934,N_230,N_300);
nand U935 (N_935,N_219,N_200);
nand U936 (N_936,N_379,N_264);
nand U937 (N_937,N_243,N_599);
nand U938 (N_938,N_485,N_478);
nor U939 (N_939,N_145,N_254);
nor U940 (N_940,N_516,N_90);
and U941 (N_941,N_680,N_216);
and U942 (N_942,N_547,N_146);
or U943 (N_943,N_17,N_194);
or U944 (N_944,N_363,N_93);
or U945 (N_945,N_133,N_78);
or U946 (N_946,N_678,N_58);
nor U947 (N_947,N_397,N_111);
xnor U948 (N_948,N_277,N_738);
or U949 (N_949,N_266,N_496);
xor U950 (N_950,N_693,N_373);
nor U951 (N_951,N_637,N_746);
nand U952 (N_952,N_513,N_613);
and U953 (N_953,N_361,N_441);
or U954 (N_954,N_682,N_308);
xnor U955 (N_955,N_288,N_376);
or U956 (N_956,N_210,N_96);
or U957 (N_957,N_460,N_250);
and U958 (N_958,N_673,N_570);
xor U959 (N_959,N_214,N_276);
nor U960 (N_960,N_684,N_476);
or U961 (N_961,N_263,N_611);
or U962 (N_962,N_317,N_412);
or U963 (N_963,N_676,N_292);
or U964 (N_964,N_156,N_479);
or U965 (N_965,N_107,N_707);
nor U966 (N_966,N_515,N_16);
nand U967 (N_967,N_232,N_571);
nand U968 (N_968,N_151,N_720);
and U969 (N_969,N_498,N_147);
xnor U970 (N_970,N_462,N_510);
nor U971 (N_971,N_382,N_72);
nand U972 (N_972,N_690,N_91);
nor U973 (N_973,N_644,N_601);
nand U974 (N_974,N_347,N_338);
xnor U975 (N_975,N_677,N_715);
nor U976 (N_976,N_140,N_576);
nand U977 (N_977,N_21,N_702);
and U978 (N_978,N_566,N_350);
nand U979 (N_979,N_248,N_454);
and U980 (N_980,N_734,N_646);
or U981 (N_981,N_11,N_618);
xnor U982 (N_982,N_135,N_457);
or U983 (N_983,N_1,N_352);
or U984 (N_984,N_298,N_149);
or U985 (N_985,N_25,N_170);
and U986 (N_986,N_341,N_53);
nand U987 (N_987,N_274,N_420);
or U988 (N_988,N_88,N_192);
nor U989 (N_989,N_275,N_667);
nor U990 (N_990,N_642,N_539);
xnor U991 (N_991,N_279,N_728);
or U992 (N_992,N_640,N_523);
xor U993 (N_993,N_240,N_581);
and U994 (N_994,N_355,N_578);
or U995 (N_995,N_632,N_497);
nor U996 (N_996,N_325,N_51);
or U997 (N_997,N_164,N_603);
and U998 (N_998,N_23,N_477);
and U999 (N_999,N_748,N_253);
nor U1000 (N_1000,N_20,N_686);
nand U1001 (N_1001,N_504,N_303);
nand U1002 (N_1002,N_545,N_344);
or U1003 (N_1003,N_333,N_452);
and U1004 (N_1004,N_395,N_393);
nand U1005 (N_1005,N_343,N_559);
xnor U1006 (N_1006,N_172,N_55);
and U1007 (N_1007,N_101,N_685);
xnor U1008 (N_1008,N_641,N_505);
nor U1009 (N_1009,N_381,N_371);
nand U1010 (N_1010,N_464,N_152);
and U1011 (N_1011,N_85,N_102);
nand U1012 (N_1012,N_427,N_735);
nor U1013 (N_1013,N_712,N_555);
or U1014 (N_1014,N_594,N_744);
nor U1015 (N_1015,N_112,N_313);
nand U1016 (N_1016,N_307,N_612);
nor U1017 (N_1017,N_588,N_327);
nand U1018 (N_1018,N_337,N_475);
nand U1019 (N_1019,N_713,N_215);
or U1020 (N_1020,N_89,N_423);
and U1021 (N_1021,N_178,N_388);
nor U1022 (N_1022,N_625,N_13);
nor U1023 (N_1023,N_60,N_195);
and U1024 (N_1024,N_654,N_251);
and U1025 (N_1025,N_272,N_166);
or U1026 (N_1026,N_584,N_281);
or U1027 (N_1027,N_233,N_529);
nor U1028 (N_1028,N_165,N_592);
and U1029 (N_1029,N_392,N_440);
or U1030 (N_1030,N_536,N_736);
and U1031 (N_1031,N_421,N_95);
or U1032 (N_1032,N_40,N_231);
xor U1033 (N_1033,N_419,N_610);
and U1034 (N_1034,N_143,N_345);
xnor U1035 (N_1035,N_719,N_399);
nor U1036 (N_1036,N_119,N_732);
or U1037 (N_1037,N_506,N_212);
and U1038 (N_1038,N_697,N_711);
or U1039 (N_1039,N_651,N_294);
nor U1040 (N_1040,N_390,N_743);
and U1041 (N_1041,N_364,N_267);
nor U1042 (N_1042,N_573,N_336);
or U1043 (N_1043,N_554,N_159);
and U1044 (N_1044,N_134,N_348);
or U1045 (N_1045,N_626,N_433);
or U1046 (N_1046,N_486,N_563);
nand U1047 (N_1047,N_369,N_726);
and U1048 (N_1048,N_687,N_162);
and U1049 (N_1049,N_123,N_322);
or U1050 (N_1050,N_71,N_33);
or U1051 (N_1051,N_569,N_296);
or U1052 (N_1052,N_537,N_174);
xnor U1053 (N_1053,N_56,N_358);
nor U1054 (N_1054,N_18,N_437);
or U1055 (N_1055,N_80,N_104);
nand U1056 (N_1056,N_161,N_604);
nand U1057 (N_1057,N_340,N_435);
or U1058 (N_1058,N_415,N_463);
nand U1059 (N_1059,N_282,N_130);
and U1060 (N_1060,N_273,N_31);
nor U1061 (N_1061,N_418,N_451);
nand U1062 (N_1062,N_196,N_83);
xor U1063 (N_1063,N_0,N_670);
or U1064 (N_1064,N_629,N_431);
nand U1065 (N_1065,N_367,N_488);
and U1066 (N_1066,N_509,N_171);
and U1067 (N_1067,N_29,N_514);
nor U1068 (N_1068,N_511,N_299);
xnor U1069 (N_1069,N_466,N_175);
nand U1070 (N_1070,N_349,N_255);
and U1071 (N_1071,N_100,N_259);
or U1072 (N_1072,N_66,N_446);
nand U1073 (N_1073,N_356,N_491);
nor U1074 (N_1074,N_426,N_532);
nand U1075 (N_1075,N_406,N_293);
nor U1076 (N_1076,N_681,N_45);
nand U1077 (N_1077,N_283,N_36);
nor U1078 (N_1078,N_432,N_656);
or U1079 (N_1079,N_411,N_410);
nand U1080 (N_1080,N_114,N_593);
nor U1081 (N_1081,N_46,N_617);
xor U1082 (N_1082,N_370,N_372);
nand U1083 (N_1083,N_359,N_203);
nand U1084 (N_1084,N_575,N_202);
nand U1085 (N_1085,N_144,N_43);
xnor U1086 (N_1086,N_602,N_8);
or U1087 (N_1087,N_227,N_306);
nor U1088 (N_1088,N_645,N_265);
or U1089 (N_1089,N_623,N_201);
nor U1090 (N_1090,N_650,N_26);
and U1091 (N_1091,N_696,N_224);
nor U1092 (N_1092,N_304,N_469);
nand U1093 (N_1093,N_430,N_329);
nor U1094 (N_1094,N_471,N_396);
or U1095 (N_1095,N_453,N_487);
xor U1096 (N_1096,N_621,N_173);
and U1097 (N_1097,N_616,N_706);
nand U1098 (N_1098,N_155,N_386);
nand U1099 (N_1099,N_286,N_615);
or U1100 (N_1100,N_237,N_662);
or U1101 (N_1101,N_182,N_22);
nand U1102 (N_1102,N_375,N_235);
nor U1103 (N_1103,N_500,N_310);
nand U1104 (N_1104,N_120,N_674);
nor U1105 (N_1105,N_521,N_525);
nor U1106 (N_1106,N_405,N_502);
and U1107 (N_1107,N_169,N_360);
nor U1108 (N_1108,N_41,N_380);
nand U1109 (N_1109,N_295,N_600);
nor U1110 (N_1110,N_698,N_718);
nand U1111 (N_1111,N_627,N_387);
nand U1112 (N_1112,N_312,N_434);
nand U1113 (N_1113,N_424,N_67);
nor U1114 (N_1114,N_34,N_520);
or U1115 (N_1115,N_385,N_531);
and U1116 (N_1116,N_115,N_394);
and U1117 (N_1117,N_339,N_530);
or U1118 (N_1118,N_30,N_733);
nor U1119 (N_1119,N_620,N_714);
nand U1120 (N_1120,N_218,N_643);
and U1121 (N_1121,N_316,N_648);
and U1122 (N_1122,N_518,N_241);
or U1123 (N_1123,N_207,N_436);
or U1124 (N_1124,N_177,N_330);
nor U1125 (N_1125,N_210,N_421);
nor U1126 (N_1126,N_660,N_709);
nand U1127 (N_1127,N_15,N_49);
nor U1128 (N_1128,N_530,N_355);
nand U1129 (N_1129,N_351,N_451);
and U1130 (N_1130,N_221,N_564);
or U1131 (N_1131,N_306,N_99);
nor U1132 (N_1132,N_428,N_651);
or U1133 (N_1133,N_399,N_553);
nand U1134 (N_1134,N_154,N_518);
or U1135 (N_1135,N_217,N_498);
or U1136 (N_1136,N_251,N_407);
and U1137 (N_1137,N_694,N_422);
nand U1138 (N_1138,N_672,N_79);
nor U1139 (N_1139,N_23,N_439);
xnor U1140 (N_1140,N_534,N_710);
and U1141 (N_1141,N_253,N_78);
and U1142 (N_1142,N_721,N_329);
nor U1143 (N_1143,N_726,N_95);
nor U1144 (N_1144,N_714,N_422);
nand U1145 (N_1145,N_552,N_519);
nand U1146 (N_1146,N_401,N_298);
nand U1147 (N_1147,N_396,N_131);
or U1148 (N_1148,N_430,N_348);
nor U1149 (N_1149,N_690,N_68);
nand U1150 (N_1150,N_79,N_500);
xnor U1151 (N_1151,N_521,N_256);
nand U1152 (N_1152,N_255,N_269);
and U1153 (N_1153,N_700,N_260);
nor U1154 (N_1154,N_316,N_37);
nor U1155 (N_1155,N_583,N_329);
nand U1156 (N_1156,N_199,N_710);
and U1157 (N_1157,N_225,N_666);
or U1158 (N_1158,N_306,N_324);
nand U1159 (N_1159,N_725,N_695);
xor U1160 (N_1160,N_235,N_79);
or U1161 (N_1161,N_537,N_360);
nand U1162 (N_1162,N_214,N_346);
or U1163 (N_1163,N_598,N_226);
nand U1164 (N_1164,N_731,N_238);
nor U1165 (N_1165,N_261,N_375);
or U1166 (N_1166,N_237,N_560);
and U1167 (N_1167,N_188,N_650);
xnor U1168 (N_1168,N_618,N_200);
or U1169 (N_1169,N_640,N_299);
xor U1170 (N_1170,N_472,N_519);
or U1171 (N_1171,N_130,N_375);
nor U1172 (N_1172,N_428,N_641);
or U1173 (N_1173,N_278,N_399);
or U1174 (N_1174,N_115,N_155);
nand U1175 (N_1175,N_199,N_318);
and U1176 (N_1176,N_478,N_405);
nor U1177 (N_1177,N_478,N_527);
or U1178 (N_1178,N_513,N_106);
nand U1179 (N_1179,N_494,N_622);
xnor U1180 (N_1180,N_554,N_664);
nand U1181 (N_1181,N_593,N_718);
and U1182 (N_1182,N_119,N_429);
or U1183 (N_1183,N_558,N_5);
or U1184 (N_1184,N_607,N_728);
xnor U1185 (N_1185,N_259,N_522);
nor U1186 (N_1186,N_684,N_577);
and U1187 (N_1187,N_125,N_509);
or U1188 (N_1188,N_220,N_381);
xor U1189 (N_1189,N_110,N_97);
nand U1190 (N_1190,N_485,N_152);
nor U1191 (N_1191,N_184,N_67);
nor U1192 (N_1192,N_691,N_195);
or U1193 (N_1193,N_565,N_413);
nand U1194 (N_1194,N_6,N_181);
xnor U1195 (N_1195,N_304,N_155);
or U1196 (N_1196,N_157,N_697);
nand U1197 (N_1197,N_619,N_647);
nor U1198 (N_1198,N_129,N_304);
nor U1199 (N_1199,N_55,N_714);
nand U1200 (N_1200,N_380,N_240);
xor U1201 (N_1201,N_18,N_571);
nor U1202 (N_1202,N_45,N_704);
xor U1203 (N_1203,N_708,N_505);
or U1204 (N_1204,N_548,N_325);
nand U1205 (N_1205,N_476,N_397);
or U1206 (N_1206,N_560,N_12);
nand U1207 (N_1207,N_58,N_26);
xor U1208 (N_1208,N_134,N_500);
and U1209 (N_1209,N_491,N_460);
and U1210 (N_1210,N_126,N_533);
nand U1211 (N_1211,N_425,N_420);
nor U1212 (N_1212,N_249,N_440);
nor U1213 (N_1213,N_742,N_126);
nand U1214 (N_1214,N_210,N_333);
nor U1215 (N_1215,N_417,N_604);
xnor U1216 (N_1216,N_190,N_696);
and U1217 (N_1217,N_371,N_257);
or U1218 (N_1218,N_647,N_249);
or U1219 (N_1219,N_111,N_389);
nor U1220 (N_1220,N_591,N_368);
or U1221 (N_1221,N_589,N_12);
and U1222 (N_1222,N_253,N_625);
and U1223 (N_1223,N_325,N_183);
or U1224 (N_1224,N_167,N_634);
nand U1225 (N_1225,N_493,N_714);
or U1226 (N_1226,N_561,N_633);
nor U1227 (N_1227,N_42,N_563);
nor U1228 (N_1228,N_663,N_731);
xor U1229 (N_1229,N_742,N_288);
or U1230 (N_1230,N_212,N_293);
or U1231 (N_1231,N_737,N_198);
or U1232 (N_1232,N_38,N_710);
and U1233 (N_1233,N_440,N_673);
xor U1234 (N_1234,N_223,N_589);
or U1235 (N_1235,N_321,N_621);
nand U1236 (N_1236,N_685,N_512);
and U1237 (N_1237,N_620,N_438);
xor U1238 (N_1238,N_213,N_321);
nand U1239 (N_1239,N_179,N_551);
and U1240 (N_1240,N_186,N_694);
or U1241 (N_1241,N_192,N_512);
or U1242 (N_1242,N_430,N_456);
nor U1243 (N_1243,N_471,N_567);
and U1244 (N_1244,N_364,N_648);
and U1245 (N_1245,N_160,N_107);
nand U1246 (N_1246,N_589,N_91);
nor U1247 (N_1247,N_88,N_49);
nand U1248 (N_1248,N_523,N_615);
xor U1249 (N_1249,N_182,N_525);
and U1250 (N_1250,N_613,N_544);
or U1251 (N_1251,N_554,N_417);
nand U1252 (N_1252,N_656,N_430);
and U1253 (N_1253,N_367,N_596);
and U1254 (N_1254,N_343,N_158);
nand U1255 (N_1255,N_619,N_727);
nor U1256 (N_1256,N_41,N_48);
nand U1257 (N_1257,N_5,N_0);
or U1258 (N_1258,N_78,N_672);
nand U1259 (N_1259,N_31,N_585);
nor U1260 (N_1260,N_318,N_152);
xor U1261 (N_1261,N_657,N_701);
and U1262 (N_1262,N_353,N_646);
or U1263 (N_1263,N_343,N_506);
nand U1264 (N_1264,N_168,N_425);
and U1265 (N_1265,N_39,N_568);
and U1266 (N_1266,N_605,N_713);
nand U1267 (N_1267,N_579,N_132);
nor U1268 (N_1268,N_595,N_142);
or U1269 (N_1269,N_56,N_205);
or U1270 (N_1270,N_457,N_148);
nor U1271 (N_1271,N_677,N_730);
and U1272 (N_1272,N_336,N_714);
xnor U1273 (N_1273,N_109,N_229);
or U1274 (N_1274,N_23,N_307);
and U1275 (N_1275,N_196,N_266);
or U1276 (N_1276,N_635,N_138);
nand U1277 (N_1277,N_4,N_183);
nand U1278 (N_1278,N_455,N_161);
or U1279 (N_1279,N_674,N_522);
nand U1280 (N_1280,N_713,N_177);
xor U1281 (N_1281,N_10,N_360);
xnor U1282 (N_1282,N_635,N_314);
nand U1283 (N_1283,N_656,N_398);
and U1284 (N_1284,N_423,N_690);
or U1285 (N_1285,N_538,N_347);
or U1286 (N_1286,N_3,N_595);
and U1287 (N_1287,N_168,N_288);
nor U1288 (N_1288,N_684,N_76);
and U1289 (N_1289,N_39,N_172);
or U1290 (N_1290,N_730,N_378);
nor U1291 (N_1291,N_85,N_637);
or U1292 (N_1292,N_613,N_247);
nand U1293 (N_1293,N_24,N_670);
nand U1294 (N_1294,N_230,N_521);
and U1295 (N_1295,N_552,N_304);
nand U1296 (N_1296,N_147,N_129);
xor U1297 (N_1297,N_521,N_106);
or U1298 (N_1298,N_380,N_156);
and U1299 (N_1299,N_278,N_622);
nor U1300 (N_1300,N_373,N_274);
xor U1301 (N_1301,N_484,N_203);
or U1302 (N_1302,N_337,N_416);
and U1303 (N_1303,N_74,N_589);
and U1304 (N_1304,N_37,N_59);
or U1305 (N_1305,N_185,N_473);
or U1306 (N_1306,N_562,N_34);
xnor U1307 (N_1307,N_457,N_467);
or U1308 (N_1308,N_352,N_391);
and U1309 (N_1309,N_657,N_594);
and U1310 (N_1310,N_52,N_432);
and U1311 (N_1311,N_168,N_312);
and U1312 (N_1312,N_379,N_16);
or U1313 (N_1313,N_151,N_424);
nor U1314 (N_1314,N_532,N_491);
xor U1315 (N_1315,N_150,N_451);
nand U1316 (N_1316,N_232,N_515);
xor U1317 (N_1317,N_124,N_60);
and U1318 (N_1318,N_527,N_188);
nor U1319 (N_1319,N_160,N_305);
nor U1320 (N_1320,N_545,N_39);
nand U1321 (N_1321,N_111,N_97);
nor U1322 (N_1322,N_26,N_558);
or U1323 (N_1323,N_557,N_441);
xnor U1324 (N_1324,N_157,N_592);
nand U1325 (N_1325,N_325,N_484);
nor U1326 (N_1326,N_640,N_575);
nand U1327 (N_1327,N_143,N_479);
and U1328 (N_1328,N_254,N_679);
or U1329 (N_1329,N_193,N_507);
nor U1330 (N_1330,N_434,N_432);
nor U1331 (N_1331,N_94,N_622);
and U1332 (N_1332,N_626,N_276);
nor U1333 (N_1333,N_8,N_486);
nand U1334 (N_1334,N_649,N_136);
and U1335 (N_1335,N_439,N_674);
xor U1336 (N_1336,N_30,N_464);
and U1337 (N_1337,N_507,N_408);
or U1338 (N_1338,N_383,N_521);
nand U1339 (N_1339,N_331,N_142);
and U1340 (N_1340,N_672,N_516);
nor U1341 (N_1341,N_186,N_126);
and U1342 (N_1342,N_33,N_371);
nor U1343 (N_1343,N_40,N_219);
or U1344 (N_1344,N_248,N_11);
or U1345 (N_1345,N_533,N_672);
nand U1346 (N_1346,N_22,N_712);
nand U1347 (N_1347,N_274,N_648);
and U1348 (N_1348,N_281,N_155);
nand U1349 (N_1349,N_145,N_534);
nor U1350 (N_1350,N_293,N_253);
or U1351 (N_1351,N_377,N_439);
nor U1352 (N_1352,N_554,N_44);
xor U1353 (N_1353,N_114,N_642);
and U1354 (N_1354,N_453,N_707);
nor U1355 (N_1355,N_391,N_291);
and U1356 (N_1356,N_465,N_588);
nand U1357 (N_1357,N_185,N_444);
nand U1358 (N_1358,N_376,N_634);
and U1359 (N_1359,N_384,N_735);
or U1360 (N_1360,N_133,N_648);
nor U1361 (N_1361,N_98,N_574);
or U1362 (N_1362,N_348,N_329);
or U1363 (N_1363,N_94,N_180);
nor U1364 (N_1364,N_644,N_79);
xnor U1365 (N_1365,N_655,N_355);
nor U1366 (N_1366,N_174,N_428);
and U1367 (N_1367,N_314,N_183);
and U1368 (N_1368,N_548,N_66);
xor U1369 (N_1369,N_485,N_536);
nand U1370 (N_1370,N_541,N_572);
or U1371 (N_1371,N_284,N_582);
and U1372 (N_1372,N_211,N_201);
nor U1373 (N_1373,N_648,N_216);
or U1374 (N_1374,N_683,N_358);
nand U1375 (N_1375,N_47,N_363);
nand U1376 (N_1376,N_565,N_682);
nand U1377 (N_1377,N_502,N_746);
and U1378 (N_1378,N_435,N_223);
nand U1379 (N_1379,N_289,N_581);
nand U1380 (N_1380,N_202,N_602);
nand U1381 (N_1381,N_145,N_687);
and U1382 (N_1382,N_0,N_690);
or U1383 (N_1383,N_46,N_439);
or U1384 (N_1384,N_347,N_63);
and U1385 (N_1385,N_506,N_53);
and U1386 (N_1386,N_9,N_546);
nand U1387 (N_1387,N_35,N_377);
and U1388 (N_1388,N_105,N_682);
xor U1389 (N_1389,N_160,N_400);
and U1390 (N_1390,N_472,N_135);
nor U1391 (N_1391,N_449,N_93);
xor U1392 (N_1392,N_497,N_541);
or U1393 (N_1393,N_246,N_406);
and U1394 (N_1394,N_81,N_116);
and U1395 (N_1395,N_448,N_297);
xnor U1396 (N_1396,N_560,N_94);
or U1397 (N_1397,N_125,N_52);
nand U1398 (N_1398,N_655,N_160);
and U1399 (N_1399,N_205,N_142);
and U1400 (N_1400,N_489,N_490);
or U1401 (N_1401,N_304,N_639);
xor U1402 (N_1402,N_700,N_447);
nor U1403 (N_1403,N_529,N_220);
xor U1404 (N_1404,N_598,N_431);
or U1405 (N_1405,N_722,N_206);
xnor U1406 (N_1406,N_158,N_261);
and U1407 (N_1407,N_656,N_508);
nand U1408 (N_1408,N_443,N_276);
nor U1409 (N_1409,N_23,N_435);
and U1410 (N_1410,N_258,N_552);
nor U1411 (N_1411,N_288,N_190);
and U1412 (N_1412,N_392,N_315);
or U1413 (N_1413,N_92,N_334);
nand U1414 (N_1414,N_454,N_440);
nand U1415 (N_1415,N_485,N_637);
and U1416 (N_1416,N_122,N_545);
and U1417 (N_1417,N_273,N_672);
nand U1418 (N_1418,N_583,N_370);
or U1419 (N_1419,N_568,N_689);
nor U1420 (N_1420,N_446,N_407);
nand U1421 (N_1421,N_350,N_502);
or U1422 (N_1422,N_720,N_37);
nand U1423 (N_1423,N_327,N_384);
and U1424 (N_1424,N_128,N_164);
and U1425 (N_1425,N_220,N_330);
nand U1426 (N_1426,N_443,N_246);
nor U1427 (N_1427,N_292,N_460);
and U1428 (N_1428,N_272,N_595);
and U1429 (N_1429,N_424,N_228);
and U1430 (N_1430,N_283,N_295);
nor U1431 (N_1431,N_659,N_255);
nor U1432 (N_1432,N_341,N_483);
and U1433 (N_1433,N_315,N_197);
and U1434 (N_1434,N_635,N_334);
or U1435 (N_1435,N_721,N_214);
nand U1436 (N_1436,N_87,N_309);
nor U1437 (N_1437,N_540,N_599);
nor U1438 (N_1438,N_645,N_706);
nor U1439 (N_1439,N_29,N_7);
nor U1440 (N_1440,N_603,N_349);
or U1441 (N_1441,N_453,N_121);
nor U1442 (N_1442,N_177,N_61);
nand U1443 (N_1443,N_612,N_616);
nand U1444 (N_1444,N_129,N_122);
and U1445 (N_1445,N_679,N_219);
nor U1446 (N_1446,N_579,N_322);
or U1447 (N_1447,N_213,N_729);
or U1448 (N_1448,N_714,N_439);
or U1449 (N_1449,N_2,N_663);
or U1450 (N_1450,N_523,N_87);
xnor U1451 (N_1451,N_460,N_188);
nor U1452 (N_1452,N_111,N_373);
nand U1453 (N_1453,N_222,N_77);
or U1454 (N_1454,N_340,N_251);
or U1455 (N_1455,N_184,N_147);
nor U1456 (N_1456,N_741,N_189);
nor U1457 (N_1457,N_212,N_551);
or U1458 (N_1458,N_376,N_324);
and U1459 (N_1459,N_405,N_509);
or U1460 (N_1460,N_346,N_338);
and U1461 (N_1461,N_197,N_83);
nor U1462 (N_1462,N_189,N_546);
or U1463 (N_1463,N_658,N_45);
nor U1464 (N_1464,N_233,N_707);
nor U1465 (N_1465,N_85,N_629);
nor U1466 (N_1466,N_54,N_6);
or U1467 (N_1467,N_353,N_279);
or U1468 (N_1468,N_9,N_98);
and U1469 (N_1469,N_577,N_535);
nand U1470 (N_1470,N_197,N_627);
or U1471 (N_1471,N_648,N_65);
nor U1472 (N_1472,N_182,N_516);
nand U1473 (N_1473,N_244,N_9);
or U1474 (N_1474,N_16,N_469);
and U1475 (N_1475,N_330,N_747);
nand U1476 (N_1476,N_9,N_67);
or U1477 (N_1477,N_536,N_32);
nand U1478 (N_1478,N_543,N_555);
nand U1479 (N_1479,N_371,N_6);
and U1480 (N_1480,N_722,N_360);
or U1481 (N_1481,N_666,N_81);
and U1482 (N_1482,N_238,N_639);
nand U1483 (N_1483,N_664,N_410);
or U1484 (N_1484,N_387,N_669);
nor U1485 (N_1485,N_241,N_728);
or U1486 (N_1486,N_25,N_229);
nor U1487 (N_1487,N_523,N_726);
xnor U1488 (N_1488,N_459,N_307);
and U1489 (N_1489,N_578,N_645);
nand U1490 (N_1490,N_65,N_52);
and U1491 (N_1491,N_489,N_123);
nor U1492 (N_1492,N_85,N_154);
and U1493 (N_1493,N_713,N_187);
nor U1494 (N_1494,N_633,N_647);
nand U1495 (N_1495,N_547,N_569);
or U1496 (N_1496,N_640,N_109);
and U1497 (N_1497,N_150,N_85);
or U1498 (N_1498,N_478,N_497);
or U1499 (N_1499,N_131,N_46);
or U1500 (N_1500,N_763,N_919);
or U1501 (N_1501,N_1187,N_978);
nand U1502 (N_1502,N_956,N_1400);
or U1503 (N_1503,N_864,N_1072);
or U1504 (N_1504,N_1113,N_1279);
nand U1505 (N_1505,N_1421,N_852);
xor U1506 (N_1506,N_1445,N_1482);
nand U1507 (N_1507,N_800,N_939);
nor U1508 (N_1508,N_1425,N_1273);
nor U1509 (N_1509,N_1050,N_1168);
nor U1510 (N_1510,N_926,N_1357);
and U1511 (N_1511,N_761,N_1474);
nor U1512 (N_1512,N_1239,N_1302);
nand U1513 (N_1513,N_968,N_1033);
nor U1514 (N_1514,N_1061,N_1172);
nor U1515 (N_1515,N_1371,N_1066);
or U1516 (N_1516,N_951,N_798);
nor U1517 (N_1517,N_1136,N_1193);
xnor U1518 (N_1518,N_1032,N_1154);
and U1519 (N_1519,N_1344,N_1151);
nor U1520 (N_1520,N_1486,N_976);
or U1521 (N_1521,N_1060,N_1166);
nor U1522 (N_1522,N_1434,N_899);
xnor U1523 (N_1523,N_981,N_988);
and U1524 (N_1524,N_1000,N_881);
or U1525 (N_1525,N_1386,N_1018);
nand U1526 (N_1526,N_1184,N_883);
and U1527 (N_1527,N_1156,N_1396);
or U1528 (N_1528,N_1441,N_809);
nor U1529 (N_1529,N_778,N_1384);
nand U1530 (N_1530,N_1128,N_994);
nand U1531 (N_1531,N_1017,N_1215);
nand U1532 (N_1532,N_1062,N_921);
xor U1533 (N_1533,N_1360,N_821);
or U1534 (N_1534,N_944,N_1218);
xor U1535 (N_1535,N_1177,N_1256);
and U1536 (N_1536,N_898,N_826);
and U1537 (N_1537,N_1394,N_1467);
and U1538 (N_1538,N_1047,N_1041);
or U1539 (N_1539,N_795,N_1088);
xnor U1540 (N_1540,N_1496,N_1469);
xor U1541 (N_1541,N_992,N_1162);
or U1542 (N_1542,N_758,N_1497);
and U1543 (N_1543,N_995,N_764);
nand U1544 (N_1544,N_1237,N_780);
nand U1545 (N_1545,N_1324,N_1461);
nor U1546 (N_1546,N_891,N_873);
nor U1547 (N_1547,N_1208,N_1373);
xor U1548 (N_1548,N_762,N_816);
nand U1549 (N_1549,N_960,N_886);
nor U1550 (N_1550,N_1163,N_1102);
nor U1551 (N_1551,N_1011,N_1429);
xnor U1552 (N_1552,N_1476,N_1259);
nor U1553 (N_1553,N_1325,N_1406);
or U1554 (N_1554,N_1119,N_1112);
and U1555 (N_1555,N_945,N_950);
nand U1556 (N_1556,N_1268,N_784);
or U1557 (N_1557,N_1439,N_938);
and U1558 (N_1558,N_1432,N_894);
xor U1559 (N_1559,N_1220,N_937);
or U1560 (N_1560,N_833,N_1299);
and U1561 (N_1561,N_1349,N_1448);
and U1562 (N_1562,N_1214,N_837);
nand U1563 (N_1563,N_1035,N_1167);
nand U1564 (N_1564,N_989,N_1457);
nor U1565 (N_1565,N_927,N_811);
or U1566 (N_1566,N_1413,N_1235);
nand U1567 (N_1567,N_815,N_1092);
or U1568 (N_1568,N_1030,N_940);
or U1569 (N_1569,N_757,N_1276);
or U1570 (N_1570,N_949,N_885);
nand U1571 (N_1571,N_1318,N_1219);
nand U1572 (N_1572,N_922,N_839);
or U1573 (N_1573,N_1415,N_1494);
nand U1574 (N_1574,N_842,N_1334);
or U1575 (N_1575,N_1155,N_835);
and U1576 (N_1576,N_1212,N_1340);
or U1577 (N_1577,N_1255,N_1122);
or U1578 (N_1578,N_1328,N_1309);
or U1579 (N_1579,N_916,N_1149);
nand U1580 (N_1580,N_932,N_760);
nand U1581 (N_1581,N_923,N_1191);
and U1582 (N_1582,N_1037,N_1174);
nand U1583 (N_1583,N_772,N_1491);
xnor U1584 (N_1584,N_1206,N_1294);
or U1585 (N_1585,N_1086,N_1307);
and U1586 (N_1586,N_1404,N_1414);
nor U1587 (N_1587,N_998,N_1068);
nor U1588 (N_1588,N_874,N_896);
or U1589 (N_1589,N_828,N_1228);
nor U1590 (N_1590,N_1375,N_1278);
or U1591 (N_1591,N_1372,N_1312);
nand U1592 (N_1592,N_759,N_930);
and U1593 (N_1593,N_860,N_1189);
and U1594 (N_1594,N_977,N_996);
and U1595 (N_1595,N_958,N_790);
or U1596 (N_1596,N_973,N_1153);
nand U1597 (N_1597,N_1192,N_913);
nor U1598 (N_1598,N_1493,N_997);
or U1599 (N_1599,N_1383,N_1269);
and U1600 (N_1600,N_1115,N_1481);
nand U1601 (N_1601,N_831,N_1132);
nand U1602 (N_1602,N_1329,N_1120);
nor U1603 (N_1603,N_1498,N_1169);
nand U1604 (N_1604,N_1225,N_1099);
or U1605 (N_1605,N_1079,N_1171);
and U1606 (N_1606,N_975,N_777);
or U1607 (N_1607,N_955,N_972);
nand U1608 (N_1608,N_1364,N_1101);
or U1609 (N_1609,N_1379,N_1089);
nand U1610 (N_1610,N_1358,N_1277);
xnor U1611 (N_1611,N_857,N_822);
nor U1612 (N_1612,N_1173,N_1094);
and U1613 (N_1613,N_1186,N_1181);
or U1614 (N_1614,N_775,N_1013);
nor U1615 (N_1615,N_771,N_767);
nand U1616 (N_1616,N_752,N_1065);
xnor U1617 (N_1617,N_1117,N_861);
xnor U1618 (N_1618,N_1180,N_1343);
nor U1619 (N_1619,N_1038,N_1222);
nor U1620 (N_1620,N_967,N_903);
or U1621 (N_1621,N_840,N_1296);
nand U1622 (N_1622,N_1209,N_1342);
and U1623 (N_1623,N_877,N_1346);
nand U1624 (N_1624,N_813,N_832);
nor U1625 (N_1625,N_1430,N_1240);
or U1626 (N_1626,N_1361,N_1282);
xnor U1627 (N_1627,N_1407,N_1110);
nand U1628 (N_1628,N_1283,N_1263);
or U1629 (N_1629,N_901,N_925);
nor U1630 (N_1630,N_1285,N_1422);
and U1631 (N_1631,N_1236,N_1080);
and U1632 (N_1632,N_1368,N_1139);
nand U1633 (N_1633,N_855,N_1385);
nand U1634 (N_1634,N_970,N_1367);
xor U1635 (N_1635,N_1217,N_797);
nand U1636 (N_1636,N_1380,N_1232);
and U1637 (N_1637,N_965,N_1316);
nand U1638 (N_1638,N_1025,N_801);
nor U1639 (N_1639,N_1142,N_1241);
nand U1640 (N_1640,N_808,N_1165);
and U1641 (N_1641,N_1160,N_1144);
xnor U1642 (N_1642,N_1459,N_829);
or U1643 (N_1643,N_1103,N_1056);
or U1644 (N_1644,N_1071,N_933);
nand U1645 (N_1645,N_979,N_1034);
nand U1646 (N_1646,N_1007,N_867);
nand U1647 (N_1647,N_1135,N_1393);
and U1648 (N_1648,N_1100,N_1073);
nand U1649 (N_1649,N_1456,N_1387);
xnor U1650 (N_1650,N_1266,N_1444);
xor U1651 (N_1651,N_980,N_1488);
or U1652 (N_1652,N_1322,N_1244);
and U1653 (N_1653,N_1012,N_1319);
nand U1654 (N_1654,N_900,N_850);
nand U1655 (N_1655,N_1303,N_845);
nor U1656 (N_1656,N_1365,N_1287);
nor U1657 (N_1657,N_1004,N_1118);
nor U1658 (N_1658,N_1010,N_1194);
nand U1659 (N_1659,N_1224,N_805);
or U1660 (N_1660,N_1138,N_1433);
and U1661 (N_1661,N_1008,N_966);
or U1662 (N_1662,N_1363,N_1262);
nor U1663 (N_1663,N_1040,N_803);
nand U1664 (N_1664,N_1216,N_1320);
xnor U1665 (N_1665,N_1473,N_1108);
nand U1666 (N_1666,N_1460,N_904);
xnor U1667 (N_1667,N_1016,N_1426);
or U1668 (N_1668,N_1234,N_756);
nor U1669 (N_1669,N_1416,N_1202);
xnor U1670 (N_1670,N_802,N_1024);
xor U1671 (N_1671,N_910,N_1313);
xnor U1672 (N_1672,N_1083,N_889);
nor U1673 (N_1673,N_1021,N_1447);
nor U1674 (N_1674,N_880,N_1435);
nor U1675 (N_1675,N_924,N_1399);
nor U1676 (N_1676,N_1001,N_1029);
nand U1677 (N_1677,N_1350,N_911);
nor U1678 (N_1678,N_1158,N_765);
and U1679 (N_1679,N_1226,N_1391);
or U1680 (N_1680,N_1337,N_1455);
nor U1681 (N_1681,N_1438,N_1348);
and U1682 (N_1682,N_1417,N_1051);
and U1683 (N_1683,N_1145,N_768);
nor U1684 (N_1684,N_1114,N_1454);
and U1685 (N_1685,N_1431,N_1484);
and U1686 (N_1686,N_1339,N_1131);
or U1687 (N_1687,N_953,N_1188);
and U1688 (N_1688,N_830,N_936);
nor U1689 (N_1689,N_1116,N_1419);
xnor U1690 (N_1690,N_1048,N_1200);
and U1691 (N_1691,N_1347,N_893);
nand U1692 (N_1692,N_1267,N_1472);
nor U1693 (N_1693,N_1074,N_1466);
or U1694 (N_1694,N_1070,N_1211);
xor U1695 (N_1695,N_1123,N_1143);
or U1696 (N_1696,N_827,N_865);
and U1697 (N_1697,N_908,N_820);
and U1698 (N_1698,N_1392,N_1341);
and U1699 (N_1699,N_1317,N_844);
nor U1700 (N_1700,N_856,N_1308);
nand U1701 (N_1701,N_1451,N_1264);
xor U1702 (N_1702,N_1362,N_1449);
and U1703 (N_1703,N_750,N_853);
nor U1704 (N_1704,N_1015,N_902);
and U1705 (N_1705,N_1463,N_1111);
nand U1706 (N_1706,N_1293,N_858);
and U1707 (N_1707,N_934,N_1332);
nand U1708 (N_1708,N_818,N_1003);
and U1709 (N_1709,N_1223,N_1125);
nor U1710 (N_1710,N_1067,N_1284);
nor U1711 (N_1711,N_1301,N_1085);
and U1712 (N_1712,N_1398,N_1412);
nor U1713 (N_1713,N_1458,N_1164);
and U1714 (N_1714,N_1077,N_773);
nor U1715 (N_1715,N_793,N_1377);
nor U1716 (N_1716,N_1195,N_1253);
nor U1717 (N_1717,N_1388,N_897);
or U1718 (N_1718,N_1196,N_1082);
nor U1719 (N_1719,N_961,N_917);
xnor U1720 (N_1720,N_1064,N_1331);
and U1721 (N_1721,N_1271,N_1261);
nand U1722 (N_1722,N_1440,N_1275);
nand U1723 (N_1723,N_1055,N_868);
or U1724 (N_1724,N_905,N_1323);
xor U1725 (N_1725,N_1036,N_1159);
nor U1726 (N_1726,N_1280,N_943);
and U1727 (N_1727,N_993,N_1095);
or U1728 (N_1728,N_1436,N_1039);
nor U1729 (N_1729,N_1321,N_1069);
or U1730 (N_1730,N_1298,N_788);
nor U1731 (N_1731,N_1420,N_888);
nand U1732 (N_1732,N_963,N_985);
nand U1733 (N_1733,N_1198,N_1292);
nand U1734 (N_1734,N_952,N_1295);
or U1735 (N_1735,N_942,N_838);
nand U1736 (N_1736,N_1464,N_1479);
xor U1737 (N_1737,N_1306,N_1106);
nor U1738 (N_1738,N_786,N_1242);
nand U1739 (N_1739,N_969,N_1356);
nand U1740 (N_1740,N_834,N_1366);
nand U1741 (N_1741,N_1096,N_876);
xnor U1742 (N_1742,N_1330,N_1270);
and U1743 (N_1743,N_1205,N_1403);
nand U1744 (N_1744,N_1249,N_959);
and U1745 (N_1745,N_841,N_872);
nand U1746 (N_1746,N_1150,N_1028);
nor U1747 (N_1747,N_779,N_1084);
nand U1748 (N_1748,N_1442,N_1097);
nand U1749 (N_1749,N_806,N_812);
or U1750 (N_1750,N_1178,N_1210);
nand U1751 (N_1751,N_1370,N_948);
nor U1752 (N_1752,N_890,N_879);
nand U1753 (N_1753,N_974,N_766);
nor U1754 (N_1754,N_794,N_1471);
and U1755 (N_1755,N_957,N_1045);
nand U1756 (N_1756,N_1126,N_1410);
or U1757 (N_1757,N_1311,N_1201);
or U1758 (N_1758,N_1374,N_1408);
nand U1759 (N_1759,N_920,N_907);
xor U1760 (N_1760,N_1203,N_863);
or U1761 (N_1761,N_1395,N_906);
xnor U1762 (N_1762,N_1063,N_1355);
xnor U1763 (N_1763,N_1245,N_1221);
or U1764 (N_1764,N_1019,N_1152);
and U1765 (N_1765,N_847,N_836);
nor U1766 (N_1766,N_1207,N_1243);
nand U1767 (N_1767,N_1009,N_1170);
and U1768 (N_1768,N_1376,N_1327);
nor U1769 (N_1769,N_1489,N_1495);
or U1770 (N_1770,N_1052,N_755);
or U1771 (N_1771,N_1290,N_791);
and U1772 (N_1772,N_787,N_1251);
nand U1773 (N_1773,N_1310,N_1470);
nor U1774 (N_1774,N_1492,N_1049);
nand U1775 (N_1775,N_1252,N_954);
and U1776 (N_1776,N_1480,N_781);
nor U1777 (N_1777,N_1418,N_971);
nand U1778 (N_1778,N_947,N_986);
or U1779 (N_1779,N_1076,N_875);
or U1780 (N_1780,N_1353,N_892);
and U1781 (N_1781,N_1129,N_1230);
or U1782 (N_1782,N_851,N_1081);
nor U1783 (N_1783,N_1390,N_792);
or U1784 (N_1784,N_895,N_817);
and U1785 (N_1785,N_1258,N_1402);
and U1786 (N_1786,N_1109,N_1104);
nor U1787 (N_1787,N_1254,N_1305);
nor U1788 (N_1788,N_823,N_870);
xnor U1789 (N_1789,N_1176,N_1179);
nor U1790 (N_1790,N_1054,N_1359);
and U1791 (N_1791,N_1190,N_1437);
xor U1792 (N_1792,N_1397,N_1401);
and U1793 (N_1793,N_1314,N_807);
xnor U1794 (N_1794,N_819,N_866);
nor U1795 (N_1795,N_1078,N_1462);
or U1796 (N_1796,N_1427,N_1185);
nand U1797 (N_1797,N_914,N_814);
and U1798 (N_1798,N_1053,N_1022);
or U1799 (N_1799,N_1288,N_1428);
nor U1800 (N_1800,N_871,N_843);
nor U1801 (N_1801,N_846,N_1213);
nor U1802 (N_1802,N_1453,N_1124);
xor U1803 (N_1803,N_1057,N_1199);
nor U1804 (N_1804,N_1197,N_1409);
nor U1805 (N_1805,N_774,N_869);
nand U1806 (N_1806,N_789,N_1059);
or U1807 (N_1807,N_1475,N_982);
or U1808 (N_1808,N_1105,N_824);
xor U1809 (N_1809,N_1443,N_1090);
and U1810 (N_1810,N_1354,N_1140);
or U1811 (N_1811,N_848,N_1075);
and U1812 (N_1812,N_1274,N_1137);
or U1813 (N_1813,N_849,N_946);
nor U1814 (N_1814,N_783,N_1157);
or U1815 (N_1815,N_1248,N_754);
xor U1816 (N_1816,N_782,N_935);
or U1817 (N_1817,N_1093,N_1130);
or U1818 (N_1818,N_1250,N_1351);
or U1819 (N_1819,N_990,N_1183);
or U1820 (N_1820,N_1450,N_1161);
nand U1821 (N_1821,N_1423,N_796);
nor U1822 (N_1822,N_1446,N_1175);
and U1823 (N_1823,N_1091,N_1134);
and U1824 (N_1824,N_770,N_1247);
and U1825 (N_1825,N_1369,N_825);
or U1826 (N_1826,N_1141,N_1023);
or U1827 (N_1827,N_918,N_1424);
nor U1828 (N_1828,N_991,N_1291);
or U1829 (N_1829,N_1336,N_1147);
nand U1830 (N_1830,N_1204,N_1483);
and U1831 (N_1831,N_929,N_1182);
nor U1832 (N_1832,N_1257,N_1382);
nand U1833 (N_1833,N_1002,N_751);
and U1834 (N_1834,N_1272,N_1133);
or U1835 (N_1835,N_1297,N_912);
and U1836 (N_1836,N_1227,N_1026);
nor U1837 (N_1837,N_1014,N_1046);
and U1838 (N_1838,N_1485,N_1148);
nand U1839 (N_1839,N_804,N_1465);
nand U1840 (N_1840,N_1378,N_1478);
xor U1841 (N_1841,N_1005,N_984);
and U1842 (N_1842,N_1487,N_1231);
and U1843 (N_1843,N_1229,N_882);
or U1844 (N_1844,N_964,N_810);
nor U1845 (N_1845,N_962,N_983);
nand U1846 (N_1846,N_854,N_999);
or U1847 (N_1847,N_1326,N_1289);
or U1848 (N_1848,N_1246,N_1300);
xor U1849 (N_1849,N_1338,N_878);
and U1850 (N_1850,N_1304,N_1027);
nand U1851 (N_1851,N_862,N_1031);
nand U1852 (N_1852,N_1490,N_1345);
or U1853 (N_1853,N_987,N_859);
and U1854 (N_1854,N_909,N_1352);
nor U1855 (N_1855,N_1233,N_1043);
and U1856 (N_1856,N_915,N_1468);
and U1857 (N_1857,N_1499,N_1006);
or U1858 (N_1858,N_776,N_1020);
nand U1859 (N_1859,N_769,N_1146);
nand U1860 (N_1860,N_887,N_1107);
nand U1861 (N_1861,N_1405,N_799);
or U1862 (N_1862,N_1315,N_941);
xnor U1863 (N_1863,N_1098,N_1335);
nor U1864 (N_1864,N_1389,N_753);
and U1865 (N_1865,N_1238,N_1452);
nand U1866 (N_1866,N_1127,N_931);
or U1867 (N_1867,N_1087,N_1281);
or U1868 (N_1868,N_884,N_1042);
nand U1869 (N_1869,N_785,N_1381);
nor U1870 (N_1870,N_1411,N_1260);
nor U1871 (N_1871,N_1058,N_1333);
and U1872 (N_1872,N_1044,N_1477);
xor U1873 (N_1873,N_1121,N_928);
xor U1874 (N_1874,N_1286,N_1265);
xnor U1875 (N_1875,N_967,N_1097);
or U1876 (N_1876,N_1120,N_1456);
xor U1877 (N_1877,N_1066,N_1137);
xnor U1878 (N_1878,N_1471,N_862);
and U1879 (N_1879,N_1263,N_1198);
or U1880 (N_1880,N_1495,N_1463);
xor U1881 (N_1881,N_1283,N_1242);
nand U1882 (N_1882,N_1279,N_948);
nor U1883 (N_1883,N_1219,N_1371);
or U1884 (N_1884,N_1474,N_1218);
or U1885 (N_1885,N_1284,N_1349);
nor U1886 (N_1886,N_772,N_886);
xnor U1887 (N_1887,N_981,N_1033);
nor U1888 (N_1888,N_1235,N_1437);
nor U1889 (N_1889,N_1202,N_783);
and U1890 (N_1890,N_1007,N_1241);
or U1891 (N_1891,N_1115,N_1400);
or U1892 (N_1892,N_1254,N_1389);
or U1893 (N_1893,N_1348,N_1120);
xor U1894 (N_1894,N_1079,N_1236);
nor U1895 (N_1895,N_1182,N_1361);
and U1896 (N_1896,N_796,N_1092);
and U1897 (N_1897,N_1254,N_1123);
nand U1898 (N_1898,N_1039,N_1254);
or U1899 (N_1899,N_1088,N_1215);
and U1900 (N_1900,N_1025,N_1375);
or U1901 (N_1901,N_1241,N_790);
or U1902 (N_1902,N_1216,N_1304);
or U1903 (N_1903,N_1464,N_1281);
and U1904 (N_1904,N_1339,N_1399);
xnor U1905 (N_1905,N_817,N_982);
and U1906 (N_1906,N_830,N_962);
or U1907 (N_1907,N_795,N_757);
nand U1908 (N_1908,N_909,N_886);
or U1909 (N_1909,N_1307,N_979);
or U1910 (N_1910,N_983,N_1251);
or U1911 (N_1911,N_1089,N_1037);
and U1912 (N_1912,N_1466,N_795);
or U1913 (N_1913,N_904,N_828);
nand U1914 (N_1914,N_799,N_1493);
or U1915 (N_1915,N_1106,N_1396);
or U1916 (N_1916,N_1442,N_1161);
nand U1917 (N_1917,N_1390,N_1042);
or U1918 (N_1918,N_1418,N_1172);
nor U1919 (N_1919,N_1189,N_1304);
and U1920 (N_1920,N_1075,N_1114);
and U1921 (N_1921,N_1112,N_933);
or U1922 (N_1922,N_890,N_1018);
nand U1923 (N_1923,N_1129,N_1370);
nand U1924 (N_1924,N_768,N_1235);
and U1925 (N_1925,N_1169,N_926);
nor U1926 (N_1926,N_1128,N_785);
and U1927 (N_1927,N_783,N_761);
nor U1928 (N_1928,N_1207,N_1014);
nand U1929 (N_1929,N_1146,N_1170);
nor U1930 (N_1930,N_1356,N_900);
xnor U1931 (N_1931,N_844,N_1024);
nor U1932 (N_1932,N_1418,N_764);
xor U1933 (N_1933,N_959,N_1131);
nand U1934 (N_1934,N_1450,N_1472);
or U1935 (N_1935,N_1061,N_994);
and U1936 (N_1936,N_1449,N_1277);
or U1937 (N_1937,N_968,N_1376);
and U1938 (N_1938,N_1373,N_1247);
xnor U1939 (N_1939,N_835,N_1181);
or U1940 (N_1940,N_1471,N_1457);
nor U1941 (N_1941,N_1037,N_1293);
xnor U1942 (N_1942,N_1306,N_1386);
or U1943 (N_1943,N_1405,N_927);
nor U1944 (N_1944,N_1296,N_984);
nor U1945 (N_1945,N_1262,N_1114);
nor U1946 (N_1946,N_921,N_1380);
nand U1947 (N_1947,N_1146,N_1469);
and U1948 (N_1948,N_1044,N_1269);
and U1949 (N_1949,N_839,N_854);
xor U1950 (N_1950,N_855,N_1089);
or U1951 (N_1951,N_829,N_757);
and U1952 (N_1952,N_844,N_1183);
nand U1953 (N_1953,N_884,N_1496);
and U1954 (N_1954,N_1420,N_1189);
xnor U1955 (N_1955,N_760,N_1124);
nor U1956 (N_1956,N_1151,N_804);
nor U1957 (N_1957,N_1153,N_845);
nor U1958 (N_1958,N_1305,N_1440);
or U1959 (N_1959,N_1206,N_840);
nor U1960 (N_1960,N_977,N_1100);
or U1961 (N_1961,N_944,N_1349);
nand U1962 (N_1962,N_799,N_1409);
nand U1963 (N_1963,N_1372,N_1450);
or U1964 (N_1964,N_1450,N_1337);
or U1965 (N_1965,N_1183,N_1203);
and U1966 (N_1966,N_1304,N_1395);
and U1967 (N_1967,N_1078,N_1465);
nor U1968 (N_1968,N_838,N_1212);
or U1969 (N_1969,N_932,N_1206);
nor U1970 (N_1970,N_1370,N_846);
nor U1971 (N_1971,N_1056,N_1383);
and U1972 (N_1972,N_1494,N_1135);
nor U1973 (N_1973,N_770,N_1027);
nor U1974 (N_1974,N_1076,N_798);
and U1975 (N_1975,N_1340,N_1013);
nand U1976 (N_1976,N_991,N_818);
nor U1977 (N_1977,N_1092,N_1177);
and U1978 (N_1978,N_814,N_958);
or U1979 (N_1979,N_890,N_1050);
nor U1980 (N_1980,N_1397,N_1486);
nor U1981 (N_1981,N_967,N_1394);
or U1982 (N_1982,N_826,N_782);
nor U1983 (N_1983,N_1056,N_1100);
and U1984 (N_1984,N_1033,N_1483);
nor U1985 (N_1985,N_1177,N_1271);
and U1986 (N_1986,N_1022,N_975);
nand U1987 (N_1987,N_838,N_1192);
and U1988 (N_1988,N_1325,N_1298);
nor U1989 (N_1989,N_803,N_1258);
and U1990 (N_1990,N_828,N_1489);
nor U1991 (N_1991,N_1170,N_1338);
or U1992 (N_1992,N_1377,N_1035);
nor U1993 (N_1993,N_845,N_1271);
nand U1994 (N_1994,N_830,N_980);
nand U1995 (N_1995,N_1247,N_1177);
nor U1996 (N_1996,N_1296,N_754);
or U1997 (N_1997,N_1026,N_948);
and U1998 (N_1998,N_1191,N_770);
nor U1999 (N_1999,N_1381,N_980);
and U2000 (N_2000,N_1128,N_808);
or U2001 (N_2001,N_1014,N_1462);
and U2002 (N_2002,N_956,N_1356);
or U2003 (N_2003,N_1116,N_1337);
nor U2004 (N_2004,N_955,N_1422);
or U2005 (N_2005,N_842,N_890);
nor U2006 (N_2006,N_1294,N_1487);
and U2007 (N_2007,N_1284,N_812);
xor U2008 (N_2008,N_1010,N_881);
and U2009 (N_2009,N_823,N_751);
nand U2010 (N_2010,N_1241,N_1032);
and U2011 (N_2011,N_909,N_996);
nor U2012 (N_2012,N_1056,N_1426);
or U2013 (N_2013,N_1076,N_872);
nand U2014 (N_2014,N_1416,N_776);
nor U2015 (N_2015,N_1455,N_933);
or U2016 (N_2016,N_950,N_982);
nand U2017 (N_2017,N_1305,N_1367);
nor U2018 (N_2018,N_873,N_805);
and U2019 (N_2019,N_1239,N_958);
xnor U2020 (N_2020,N_1378,N_1071);
and U2021 (N_2021,N_1459,N_952);
and U2022 (N_2022,N_964,N_1493);
or U2023 (N_2023,N_1157,N_977);
and U2024 (N_2024,N_994,N_1293);
or U2025 (N_2025,N_1163,N_1249);
nand U2026 (N_2026,N_840,N_1114);
nor U2027 (N_2027,N_771,N_914);
or U2028 (N_2028,N_1332,N_1400);
or U2029 (N_2029,N_1411,N_1267);
nand U2030 (N_2030,N_893,N_1159);
or U2031 (N_2031,N_1258,N_1453);
and U2032 (N_2032,N_1425,N_894);
xor U2033 (N_2033,N_1131,N_856);
nand U2034 (N_2034,N_1164,N_1053);
and U2035 (N_2035,N_1221,N_1477);
or U2036 (N_2036,N_911,N_1056);
xnor U2037 (N_2037,N_1328,N_886);
xor U2038 (N_2038,N_1416,N_1338);
or U2039 (N_2039,N_914,N_1153);
nand U2040 (N_2040,N_1434,N_1268);
or U2041 (N_2041,N_1112,N_909);
xnor U2042 (N_2042,N_1465,N_1132);
or U2043 (N_2043,N_1019,N_975);
nor U2044 (N_2044,N_1284,N_839);
nor U2045 (N_2045,N_1263,N_1247);
xor U2046 (N_2046,N_777,N_901);
nand U2047 (N_2047,N_1308,N_1461);
nand U2048 (N_2048,N_775,N_1250);
or U2049 (N_2049,N_1363,N_1107);
and U2050 (N_2050,N_1041,N_847);
xor U2051 (N_2051,N_1089,N_761);
or U2052 (N_2052,N_759,N_1196);
and U2053 (N_2053,N_1496,N_1081);
and U2054 (N_2054,N_906,N_1026);
or U2055 (N_2055,N_1012,N_845);
or U2056 (N_2056,N_1241,N_1456);
or U2057 (N_2057,N_1451,N_1130);
and U2058 (N_2058,N_1497,N_1264);
or U2059 (N_2059,N_782,N_1309);
or U2060 (N_2060,N_1387,N_1020);
nand U2061 (N_2061,N_1319,N_885);
nand U2062 (N_2062,N_895,N_1319);
and U2063 (N_2063,N_769,N_884);
or U2064 (N_2064,N_1382,N_995);
nand U2065 (N_2065,N_895,N_1364);
or U2066 (N_2066,N_884,N_1489);
and U2067 (N_2067,N_1184,N_1198);
nor U2068 (N_2068,N_1477,N_823);
xnor U2069 (N_2069,N_900,N_1019);
or U2070 (N_2070,N_1328,N_1497);
or U2071 (N_2071,N_1273,N_766);
or U2072 (N_2072,N_897,N_1044);
or U2073 (N_2073,N_1387,N_1220);
and U2074 (N_2074,N_793,N_1302);
or U2075 (N_2075,N_1413,N_1172);
and U2076 (N_2076,N_1097,N_1216);
and U2077 (N_2077,N_1337,N_1234);
and U2078 (N_2078,N_1132,N_1226);
nand U2079 (N_2079,N_1493,N_1378);
or U2080 (N_2080,N_1491,N_1008);
or U2081 (N_2081,N_984,N_1290);
nand U2082 (N_2082,N_1270,N_1048);
nor U2083 (N_2083,N_869,N_1137);
nand U2084 (N_2084,N_1361,N_948);
nor U2085 (N_2085,N_873,N_895);
nor U2086 (N_2086,N_1376,N_1077);
nand U2087 (N_2087,N_1220,N_952);
xor U2088 (N_2088,N_1126,N_892);
and U2089 (N_2089,N_805,N_1217);
nand U2090 (N_2090,N_944,N_1009);
and U2091 (N_2091,N_937,N_1025);
nand U2092 (N_2092,N_979,N_1279);
nor U2093 (N_2093,N_1002,N_1155);
nand U2094 (N_2094,N_913,N_1216);
nand U2095 (N_2095,N_1295,N_1422);
nand U2096 (N_2096,N_1064,N_1478);
xor U2097 (N_2097,N_863,N_1171);
nand U2098 (N_2098,N_1004,N_1475);
and U2099 (N_2099,N_1095,N_824);
or U2100 (N_2100,N_964,N_1308);
xor U2101 (N_2101,N_1159,N_1422);
nor U2102 (N_2102,N_1171,N_1035);
or U2103 (N_2103,N_1278,N_1113);
nor U2104 (N_2104,N_831,N_934);
nand U2105 (N_2105,N_1191,N_1234);
nor U2106 (N_2106,N_864,N_1463);
and U2107 (N_2107,N_1067,N_869);
nor U2108 (N_2108,N_1424,N_978);
nor U2109 (N_2109,N_990,N_928);
or U2110 (N_2110,N_1208,N_948);
or U2111 (N_2111,N_986,N_1311);
or U2112 (N_2112,N_1127,N_1265);
xor U2113 (N_2113,N_1117,N_1239);
xor U2114 (N_2114,N_1088,N_1485);
or U2115 (N_2115,N_1266,N_858);
and U2116 (N_2116,N_1031,N_1015);
and U2117 (N_2117,N_754,N_1034);
nand U2118 (N_2118,N_790,N_1066);
xor U2119 (N_2119,N_1004,N_941);
nor U2120 (N_2120,N_980,N_1042);
nor U2121 (N_2121,N_1264,N_1413);
xor U2122 (N_2122,N_1499,N_1092);
nand U2123 (N_2123,N_1181,N_1115);
xor U2124 (N_2124,N_916,N_1340);
xor U2125 (N_2125,N_943,N_1492);
and U2126 (N_2126,N_1359,N_1223);
nor U2127 (N_2127,N_1264,N_1163);
nor U2128 (N_2128,N_850,N_1357);
or U2129 (N_2129,N_1061,N_1283);
and U2130 (N_2130,N_1009,N_887);
nor U2131 (N_2131,N_926,N_951);
or U2132 (N_2132,N_1488,N_1226);
xnor U2133 (N_2133,N_758,N_865);
nor U2134 (N_2134,N_901,N_1436);
nand U2135 (N_2135,N_1166,N_1219);
xor U2136 (N_2136,N_845,N_870);
nand U2137 (N_2137,N_1092,N_956);
nand U2138 (N_2138,N_896,N_1214);
xor U2139 (N_2139,N_1238,N_1161);
nor U2140 (N_2140,N_1142,N_1115);
nand U2141 (N_2141,N_1010,N_1173);
nor U2142 (N_2142,N_1176,N_1013);
and U2143 (N_2143,N_1103,N_1025);
nor U2144 (N_2144,N_1499,N_1145);
and U2145 (N_2145,N_871,N_981);
and U2146 (N_2146,N_1437,N_1341);
and U2147 (N_2147,N_917,N_1086);
or U2148 (N_2148,N_881,N_1282);
nand U2149 (N_2149,N_1166,N_828);
nor U2150 (N_2150,N_1018,N_1405);
xor U2151 (N_2151,N_1010,N_850);
nor U2152 (N_2152,N_916,N_1210);
and U2153 (N_2153,N_774,N_1319);
nor U2154 (N_2154,N_928,N_1129);
nor U2155 (N_2155,N_1306,N_845);
or U2156 (N_2156,N_1387,N_917);
or U2157 (N_2157,N_1471,N_1496);
and U2158 (N_2158,N_1259,N_917);
nand U2159 (N_2159,N_1359,N_1013);
nand U2160 (N_2160,N_1160,N_1229);
nand U2161 (N_2161,N_978,N_1328);
or U2162 (N_2162,N_1148,N_1002);
and U2163 (N_2163,N_1372,N_1202);
or U2164 (N_2164,N_767,N_1049);
nand U2165 (N_2165,N_999,N_1278);
or U2166 (N_2166,N_982,N_1203);
and U2167 (N_2167,N_889,N_947);
nand U2168 (N_2168,N_783,N_856);
nor U2169 (N_2169,N_905,N_1408);
nand U2170 (N_2170,N_1402,N_1014);
nand U2171 (N_2171,N_1475,N_829);
and U2172 (N_2172,N_1224,N_940);
and U2173 (N_2173,N_1218,N_1206);
and U2174 (N_2174,N_785,N_916);
nor U2175 (N_2175,N_1153,N_1480);
and U2176 (N_2176,N_1422,N_1060);
and U2177 (N_2177,N_1211,N_1036);
nor U2178 (N_2178,N_1370,N_980);
or U2179 (N_2179,N_1319,N_1226);
and U2180 (N_2180,N_862,N_1003);
and U2181 (N_2181,N_1391,N_1063);
nor U2182 (N_2182,N_1217,N_1314);
nor U2183 (N_2183,N_772,N_1489);
and U2184 (N_2184,N_1137,N_1049);
or U2185 (N_2185,N_802,N_1074);
and U2186 (N_2186,N_1222,N_1019);
nand U2187 (N_2187,N_1006,N_1166);
nor U2188 (N_2188,N_1121,N_821);
or U2189 (N_2189,N_1380,N_1155);
nor U2190 (N_2190,N_1302,N_1208);
or U2191 (N_2191,N_958,N_918);
nor U2192 (N_2192,N_1108,N_802);
xnor U2193 (N_2193,N_1205,N_1429);
and U2194 (N_2194,N_1027,N_1061);
and U2195 (N_2195,N_1091,N_1322);
or U2196 (N_2196,N_1281,N_1184);
nand U2197 (N_2197,N_1038,N_1302);
xor U2198 (N_2198,N_1246,N_946);
nand U2199 (N_2199,N_1455,N_1434);
nor U2200 (N_2200,N_1165,N_1144);
nor U2201 (N_2201,N_1309,N_815);
and U2202 (N_2202,N_834,N_806);
nand U2203 (N_2203,N_810,N_944);
nand U2204 (N_2204,N_1252,N_1030);
or U2205 (N_2205,N_890,N_1303);
xnor U2206 (N_2206,N_1159,N_1440);
nor U2207 (N_2207,N_827,N_1477);
or U2208 (N_2208,N_793,N_1207);
or U2209 (N_2209,N_812,N_1128);
or U2210 (N_2210,N_1122,N_994);
and U2211 (N_2211,N_1197,N_1397);
and U2212 (N_2212,N_1418,N_1433);
and U2213 (N_2213,N_1076,N_1334);
and U2214 (N_2214,N_1230,N_1397);
or U2215 (N_2215,N_1197,N_811);
nand U2216 (N_2216,N_1348,N_1187);
and U2217 (N_2217,N_1249,N_1157);
nand U2218 (N_2218,N_1061,N_1364);
and U2219 (N_2219,N_1367,N_963);
or U2220 (N_2220,N_1055,N_1288);
nor U2221 (N_2221,N_1275,N_952);
and U2222 (N_2222,N_1058,N_1204);
or U2223 (N_2223,N_825,N_1017);
and U2224 (N_2224,N_928,N_1219);
nor U2225 (N_2225,N_881,N_1018);
or U2226 (N_2226,N_1432,N_1321);
nor U2227 (N_2227,N_921,N_931);
and U2228 (N_2228,N_1095,N_1192);
or U2229 (N_2229,N_899,N_1237);
and U2230 (N_2230,N_1144,N_1075);
nor U2231 (N_2231,N_1139,N_1084);
or U2232 (N_2232,N_1459,N_1008);
nor U2233 (N_2233,N_946,N_1256);
nor U2234 (N_2234,N_791,N_1256);
nor U2235 (N_2235,N_1261,N_1324);
and U2236 (N_2236,N_1158,N_980);
xnor U2237 (N_2237,N_1117,N_943);
and U2238 (N_2238,N_1495,N_1264);
or U2239 (N_2239,N_988,N_1404);
nand U2240 (N_2240,N_1160,N_755);
or U2241 (N_2241,N_1260,N_787);
nand U2242 (N_2242,N_1170,N_833);
or U2243 (N_2243,N_974,N_1485);
xnor U2244 (N_2244,N_836,N_834);
nor U2245 (N_2245,N_1483,N_1266);
nor U2246 (N_2246,N_1005,N_1196);
or U2247 (N_2247,N_850,N_853);
xor U2248 (N_2248,N_1038,N_1342);
or U2249 (N_2249,N_1367,N_1343);
nand U2250 (N_2250,N_1575,N_1984);
xnor U2251 (N_2251,N_2149,N_1811);
nor U2252 (N_2252,N_2203,N_2004);
xnor U2253 (N_2253,N_1578,N_2151);
nor U2254 (N_2254,N_1711,N_2146);
or U2255 (N_2255,N_1620,N_2018);
or U2256 (N_2256,N_1603,N_2034);
nor U2257 (N_2257,N_1874,N_1937);
nand U2258 (N_2258,N_1995,N_1830);
nand U2259 (N_2259,N_2068,N_1738);
nand U2260 (N_2260,N_1566,N_2160);
or U2261 (N_2261,N_1622,N_2135);
xnor U2262 (N_2262,N_1868,N_2168);
xnor U2263 (N_2263,N_2121,N_2162);
xor U2264 (N_2264,N_2042,N_2026);
nor U2265 (N_2265,N_1737,N_1978);
nor U2266 (N_2266,N_2170,N_2182);
nand U2267 (N_2267,N_2049,N_1636);
nor U2268 (N_2268,N_1854,N_2136);
or U2269 (N_2269,N_2092,N_2228);
and U2270 (N_2270,N_1649,N_1843);
and U2271 (N_2271,N_1962,N_2083);
xor U2272 (N_2272,N_1668,N_2081);
or U2273 (N_2273,N_1595,N_2057);
xnor U2274 (N_2274,N_1790,N_1630);
nor U2275 (N_2275,N_2064,N_2046);
or U2276 (N_2276,N_1893,N_1890);
and U2277 (N_2277,N_1697,N_1935);
or U2278 (N_2278,N_2131,N_2184);
nor U2279 (N_2279,N_1562,N_1709);
nor U2280 (N_2280,N_2225,N_1986);
nand U2281 (N_2281,N_1615,N_2015);
and U2282 (N_2282,N_1707,N_2229);
or U2283 (N_2283,N_1550,N_1807);
nand U2284 (N_2284,N_2100,N_1557);
xor U2285 (N_2285,N_2235,N_1524);
nand U2286 (N_2286,N_1989,N_2119);
xnor U2287 (N_2287,N_1678,N_1836);
nand U2288 (N_2288,N_1921,N_2128);
nand U2289 (N_2289,N_1739,N_2012);
nand U2290 (N_2290,N_1777,N_1509);
nor U2291 (N_2291,N_1594,N_1712);
nor U2292 (N_2292,N_1617,N_2189);
nor U2293 (N_2293,N_1934,N_1667);
and U2294 (N_2294,N_1860,N_1585);
nand U2295 (N_2295,N_1663,N_1745);
and U2296 (N_2296,N_1523,N_1928);
and U2297 (N_2297,N_1927,N_2185);
or U2298 (N_2298,N_1968,N_1702);
or U2299 (N_2299,N_2074,N_1520);
nand U2300 (N_2300,N_1583,N_1670);
nor U2301 (N_2301,N_1781,N_2187);
or U2302 (N_2302,N_1983,N_1878);
nand U2303 (N_2303,N_1788,N_2105);
nand U2304 (N_2304,N_1519,N_2080);
nor U2305 (N_2305,N_1784,N_1587);
and U2306 (N_2306,N_1643,N_1846);
xnor U2307 (N_2307,N_2208,N_2242);
nand U2308 (N_2308,N_1882,N_1640);
nor U2309 (N_2309,N_1613,N_2138);
nor U2310 (N_2310,N_1609,N_2056);
and U2311 (N_2311,N_1931,N_1693);
nand U2312 (N_2312,N_1766,N_2161);
and U2313 (N_2313,N_2063,N_1701);
nand U2314 (N_2314,N_1797,N_1941);
and U2315 (N_2315,N_1692,N_2031);
xnor U2316 (N_2316,N_1618,N_1866);
and U2317 (N_2317,N_1817,N_1671);
nor U2318 (N_2318,N_2238,N_2195);
and U2319 (N_2319,N_1875,N_1792);
nand U2320 (N_2320,N_1627,N_1706);
or U2321 (N_2321,N_1515,N_2106);
and U2322 (N_2322,N_1633,N_1803);
and U2323 (N_2323,N_2072,N_1559);
nand U2324 (N_2324,N_2051,N_1919);
nand U2325 (N_2325,N_1824,N_1782);
and U2326 (N_2326,N_1825,N_1828);
and U2327 (N_2327,N_2186,N_1999);
nor U2328 (N_2328,N_1849,N_2102);
nor U2329 (N_2329,N_2115,N_2166);
nor U2330 (N_2330,N_1717,N_1888);
nand U2331 (N_2331,N_1607,N_1954);
nand U2332 (N_2332,N_1602,N_1722);
and U2333 (N_2333,N_1873,N_2023);
or U2334 (N_2334,N_1598,N_2175);
xor U2335 (N_2335,N_1855,N_1565);
or U2336 (N_2336,N_1659,N_1699);
or U2337 (N_2337,N_2163,N_1584);
nor U2338 (N_2338,N_1512,N_2233);
xor U2339 (N_2339,N_1732,N_2231);
nand U2340 (N_2340,N_2103,N_2088);
and U2341 (N_2341,N_2240,N_1577);
nand U2342 (N_2342,N_2156,N_2243);
and U2343 (N_2343,N_1964,N_1965);
nand U2344 (N_2344,N_2247,N_1754);
nand U2345 (N_2345,N_1799,N_2141);
and U2346 (N_2346,N_2027,N_2028);
nor U2347 (N_2347,N_1916,N_2232);
or U2348 (N_2348,N_1818,N_1614);
and U2349 (N_2349,N_1703,N_2043);
nor U2350 (N_2350,N_1780,N_2040);
nor U2351 (N_2351,N_2202,N_1518);
nand U2352 (N_2352,N_1666,N_1642);
or U2353 (N_2353,N_1991,N_1987);
or U2354 (N_2354,N_1650,N_1801);
nor U2355 (N_2355,N_1522,N_1503);
or U2356 (N_2356,N_2221,N_1913);
xnor U2357 (N_2357,N_1975,N_2075);
nor U2358 (N_2358,N_1552,N_2085);
nor U2359 (N_2359,N_2101,N_1911);
nor U2360 (N_2360,N_1880,N_1749);
and U2361 (N_2361,N_1772,N_2142);
xor U2362 (N_2362,N_1853,N_1838);
nand U2363 (N_2363,N_2205,N_2219);
nand U2364 (N_2364,N_1743,N_1548);
or U2365 (N_2365,N_1530,N_1721);
or U2366 (N_2366,N_1705,N_2013);
and U2367 (N_2367,N_1651,N_2155);
nor U2368 (N_2368,N_2108,N_1943);
and U2369 (N_2369,N_2019,N_2198);
nand U2370 (N_2370,N_1885,N_2244);
or U2371 (N_2371,N_1521,N_2126);
and U2372 (N_2372,N_1918,N_2000);
and U2373 (N_2373,N_1776,N_2070);
nand U2374 (N_2374,N_1596,N_1580);
nor U2375 (N_2375,N_2183,N_1540);
or U2376 (N_2376,N_1624,N_2099);
or U2377 (N_2377,N_1778,N_1889);
or U2378 (N_2378,N_1847,N_1944);
nor U2379 (N_2379,N_1741,N_1623);
nor U2380 (N_2380,N_1563,N_1673);
and U2381 (N_2381,N_2022,N_2164);
nand U2382 (N_2382,N_1850,N_2132);
and U2383 (N_2383,N_1635,N_2177);
or U2384 (N_2384,N_1664,N_1684);
and U2385 (N_2385,N_2044,N_1771);
nor U2386 (N_2386,N_1765,N_1735);
and U2387 (N_2387,N_2062,N_1936);
nor U2388 (N_2388,N_2241,N_2098);
nand U2389 (N_2389,N_1974,N_1549);
nor U2390 (N_2390,N_1844,N_1997);
or U2391 (N_2391,N_1794,N_1611);
or U2392 (N_2392,N_1695,N_1959);
or U2393 (N_2393,N_1606,N_1813);
or U2394 (N_2394,N_1894,N_1929);
nor U2395 (N_2395,N_1500,N_2144);
nand U2396 (N_2396,N_1831,N_1629);
nand U2397 (N_2397,N_2196,N_2154);
nor U2398 (N_2398,N_1665,N_1727);
and U2399 (N_2399,N_1861,N_1661);
or U2400 (N_2400,N_2086,N_1698);
nor U2401 (N_2401,N_1800,N_1957);
and U2402 (N_2402,N_2001,N_1837);
or U2403 (N_2403,N_1976,N_1814);
nor U2404 (N_2404,N_1655,N_2130);
or U2405 (N_2405,N_2071,N_1567);
or U2406 (N_2406,N_1730,N_2113);
and U2407 (N_2407,N_1864,N_1718);
xor U2408 (N_2408,N_1648,N_1804);
xnor U2409 (N_2409,N_1715,N_2008);
or U2410 (N_2410,N_2216,N_1605);
and U2411 (N_2411,N_2096,N_2123);
nand U2412 (N_2412,N_2237,N_1869);
nand U2413 (N_2413,N_1536,N_2073);
or U2414 (N_2414,N_1992,N_2214);
nor U2415 (N_2415,N_2143,N_1586);
or U2416 (N_2416,N_1822,N_2201);
or U2417 (N_2417,N_1507,N_1681);
nor U2418 (N_2418,N_2193,N_1988);
or U2419 (N_2419,N_2145,N_2133);
nor U2420 (N_2420,N_1969,N_1841);
nand U2421 (N_2421,N_2147,N_1708);
or U2422 (N_2422,N_1973,N_1763);
nand U2423 (N_2423,N_1758,N_2180);
or U2424 (N_2424,N_1946,N_1502);
and U2425 (N_2425,N_2094,N_1501);
and U2426 (N_2426,N_1856,N_2047);
nor U2427 (N_2427,N_2041,N_1895);
or U2428 (N_2428,N_1544,N_1685);
nor U2429 (N_2429,N_2091,N_2148);
or U2430 (N_2430,N_2035,N_1555);
xor U2431 (N_2431,N_2003,N_1773);
nand U2432 (N_2432,N_2157,N_2179);
nand U2433 (N_2433,N_1917,N_1570);
nor U2434 (N_2434,N_2025,N_1795);
nand U2435 (N_2435,N_2165,N_1915);
xnor U2436 (N_2436,N_1686,N_1631);
nand U2437 (N_2437,N_1553,N_1852);
or U2438 (N_2438,N_1619,N_1528);
xor U2439 (N_2439,N_2117,N_1912);
nor U2440 (N_2440,N_1510,N_1688);
or U2441 (N_2441,N_1653,N_2021);
and U2442 (N_2442,N_1724,N_2090);
nand U2443 (N_2443,N_1508,N_1576);
nand U2444 (N_2444,N_1951,N_1541);
or U2445 (N_2445,N_1808,N_2125);
nand U2446 (N_2446,N_1764,N_1906);
and U2447 (N_2447,N_2212,N_1979);
and U2448 (N_2448,N_1848,N_1641);
nand U2449 (N_2449,N_1647,N_2093);
nor U2450 (N_2450,N_1857,N_1947);
or U2451 (N_2451,N_1687,N_1985);
nand U2452 (N_2452,N_1950,N_1791);
and U2453 (N_2453,N_2110,N_1690);
nor U2454 (N_2454,N_2122,N_1533);
or U2455 (N_2455,N_1700,N_1859);
or U2456 (N_2456,N_1783,N_1592);
or U2457 (N_2457,N_1545,N_2065);
nand U2458 (N_2458,N_1742,N_1821);
and U2459 (N_2459,N_2002,N_2139);
and U2460 (N_2460,N_2078,N_1506);
xnor U2461 (N_2461,N_1940,N_1977);
and U2462 (N_2462,N_1862,N_1704);
nand U2463 (N_2463,N_2152,N_1884);
nand U2464 (N_2464,N_1571,N_1816);
xnor U2465 (N_2465,N_2172,N_2158);
or U2466 (N_2466,N_1908,N_1637);
nand U2467 (N_2467,N_2134,N_1826);
xor U2468 (N_2468,N_1829,N_1560);
or U2469 (N_2469,N_2052,N_1879);
nand U2470 (N_2470,N_1534,N_2084);
nand U2471 (N_2471,N_2217,N_2016);
nand U2472 (N_2472,N_2129,N_1532);
nand U2473 (N_2473,N_1819,N_1672);
nor U2474 (N_2474,N_1774,N_1558);
nand U2475 (N_2475,N_2153,N_1589);
nand U2476 (N_2476,N_1963,N_1714);
nand U2477 (N_2477,N_1827,N_1744);
or U2478 (N_2478,N_1646,N_2178);
nand U2479 (N_2479,N_1677,N_1805);
or U2480 (N_2480,N_1626,N_1531);
or U2481 (N_2481,N_2069,N_1573);
or U2482 (N_2482,N_1812,N_2045);
nor U2483 (N_2483,N_1511,N_1740);
nor U2484 (N_2484,N_1802,N_2248);
or U2485 (N_2485,N_1676,N_1639);
or U2486 (N_2486,N_1632,N_1952);
nor U2487 (N_2487,N_1832,N_2190);
nor U2488 (N_2488,N_2209,N_2124);
and U2489 (N_2489,N_1581,N_1970);
nand U2490 (N_2490,N_2227,N_1517);
xor U2491 (N_2491,N_2181,N_1961);
nor U2492 (N_2492,N_1755,N_1527);
or U2493 (N_2493,N_1863,N_1504);
nor U2494 (N_2494,N_1731,N_1582);
nor U2495 (N_2495,N_2009,N_2245);
or U2496 (N_2496,N_1896,N_2211);
or U2497 (N_2497,N_1657,N_1658);
and U2498 (N_2498,N_2112,N_2006);
and U2499 (N_2499,N_1728,N_2087);
xnor U2500 (N_2500,N_1839,N_2014);
nor U2501 (N_2501,N_1820,N_2082);
and U2502 (N_2502,N_2060,N_1604);
and U2503 (N_2503,N_2118,N_1746);
and U2504 (N_2504,N_1867,N_2039);
or U2505 (N_2505,N_1725,N_1516);
nand U2506 (N_2506,N_1556,N_2033);
nor U2507 (N_2507,N_2206,N_1953);
and U2508 (N_2508,N_1956,N_1948);
and U2509 (N_2509,N_1551,N_1900);
and U2510 (N_2510,N_1770,N_1710);
or U2511 (N_2511,N_2249,N_2222);
nand U2512 (N_2512,N_1910,N_1526);
or U2513 (N_2513,N_2032,N_1591);
or U2514 (N_2514,N_1547,N_2030);
and U2515 (N_2515,N_2053,N_1716);
xnor U2516 (N_2516,N_2192,N_2024);
or U2517 (N_2517,N_2029,N_2114);
xor U2518 (N_2518,N_1726,N_1747);
nor U2519 (N_2519,N_2127,N_2150);
nor U2520 (N_2520,N_1972,N_1621);
and U2521 (N_2521,N_1752,N_1779);
nand U2522 (N_2522,N_1787,N_1966);
and U2523 (N_2523,N_1720,N_1656);
and U2524 (N_2524,N_1967,N_2050);
or U2525 (N_2525,N_1872,N_2174);
nand U2526 (N_2526,N_1662,N_2054);
or U2527 (N_2527,N_1588,N_1568);
xor U2528 (N_2528,N_2224,N_2140);
xnor U2529 (N_2529,N_1719,N_1757);
xnor U2530 (N_2530,N_1924,N_2200);
nand U2531 (N_2531,N_2104,N_1904);
or U2532 (N_2532,N_2223,N_2010);
or U2533 (N_2533,N_1561,N_2020);
xor U2534 (N_2534,N_1903,N_1572);
nand U2535 (N_2535,N_1939,N_1691);
or U2536 (N_2536,N_1682,N_2037);
or U2537 (N_2537,N_1514,N_1922);
or U2538 (N_2538,N_1891,N_2169);
or U2539 (N_2539,N_1981,N_1750);
nor U2540 (N_2540,N_2059,N_1877);
or U2541 (N_2541,N_1579,N_1674);
xor U2542 (N_2542,N_1660,N_2055);
nand U2543 (N_2543,N_2230,N_1926);
nor U2544 (N_2544,N_1842,N_1597);
xnor U2545 (N_2545,N_1753,N_1980);
and U2546 (N_2546,N_2076,N_1881);
nor U2547 (N_2547,N_1851,N_2137);
or U2548 (N_2548,N_1971,N_1767);
nand U2549 (N_2549,N_1535,N_1865);
xnor U2550 (N_2550,N_1652,N_1762);
and U2551 (N_2551,N_1645,N_2239);
xnor U2552 (N_2552,N_1883,N_1513);
nor U2553 (N_2553,N_1525,N_1902);
and U2554 (N_2554,N_1914,N_1871);
or U2555 (N_2555,N_2109,N_1736);
and U2556 (N_2556,N_2079,N_1542);
and U2557 (N_2557,N_2077,N_1590);
and U2558 (N_2558,N_1909,N_2111);
or U2559 (N_2559,N_1612,N_1625);
and U2560 (N_2560,N_1823,N_2191);
or U2561 (N_2561,N_2236,N_2089);
nor U2562 (N_2562,N_1945,N_1608);
xor U2563 (N_2563,N_1769,N_1809);
nand U2564 (N_2564,N_1644,N_1680);
or U2565 (N_2565,N_2171,N_1923);
or U2566 (N_2566,N_1713,N_2116);
and U2567 (N_2567,N_1785,N_1942);
or U2568 (N_2568,N_1564,N_1760);
and U2569 (N_2569,N_1628,N_1796);
and U2570 (N_2570,N_2210,N_1840);
xor U2571 (N_2571,N_2188,N_1675);
nor U2572 (N_2572,N_2061,N_1759);
or U2573 (N_2573,N_1810,N_2173);
xor U2574 (N_2574,N_1798,N_2011);
or U2575 (N_2575,N_1599,N_1616);
xnor U2576 (N_2576,N_2246,N_2207);
xor U2577 (N_2577,N_2017,N_1505);
xnor U2578 (N_2578,N_1733,N_1990);
nand U2579 (N_2579,N_1543,N_1634);
or U2580 (N_2580,N_2007,N_1876);
or U2581 (N_2581,N_1815,N_2176);
nand U2582 (N_2582,N_1960,N_2215);
nand U2583 (N_2583,N_1887,N_2213);
nand U2584 (N_2584,N_2048,N_1696);
xnor U2585 (N_2585,N_1932,N_2220);
nand U2586 (N_2586,N_1793,N_1925);
nor U2587 (N_2587,N_1892,N_1654);
nor U2588 (N_2588,N_2038,N_1554);
nand U2589 (N_2589,N_1679,N_2226);
nor U2590 (N_2590,N_1574,N_2058);
xnor U2591 (N_2591,N_1833,N_1569);
nor U2592 (N_2592,N_1529,N_1899);
nand U2593 (N_2593,N_1694,N_2159);
nor U2594 (N_2594,N_1898,N_1761);
nand U2595 (N_2595,N_2036,N_1897);
xnor U2596 (N_2596,N_2120,N_2194);
or U2597 (N_2597,N_1870,N_1958);
or U2598 (N_2598,N_1901,N_1930);
or U2599 (N_2599,N_1689,N_1748);
nor U2600 (N_2600,N_1593,N_1982);
nand U2601 (N_2601,N_1734,N_1601);
or U2602 (N_2602,N_1539,N_1537);
or U2603 (N_2603,N_1610,N_1786);
or U2604 (N_2604,N_1886,N_1905);
or U2605 (N_2605,N_1669,N_1858);
nand U2606 (N_2606,N_1806,N_2095);
nor U2607 (N_2607,N_2167,N_2218);
and U2608 (N_2608,N_2005,N_2066);
nor U2609 (N_2609,N_2067,N_1907);
nor U2610 (N_2610,N_2197,N_1920);
xor U2611 (N_2611,N_1546,N_2234);
and U2612 (N_2612,N_1683,N_1768);
nor U2613 (N_2613,N_1775,N_1538);
nand U2614 (N_2614,N_1751,N_1993);
or U2615 (N_2615,N_1949,N_1933);
nand U2616 (N_2616,N_1835,N_1756);
or U2617 (N_2617,N_2097,N_2107);
xnor U2618 (N_2618,N_2199,N_1834);
or U2619 (N_2619,N_1994,N_1729);
nor U2620 (N_2620,N_1996,N_1789);
nand U2621 (N_2621,N_2204,N_1938);
and U2622 (N_2622,N_1600,N_1638);
or U2623 (N_2623,N_1845,N_1955);
nand U2624 (N_2624,N_1998,N_1723);
or U2625 (N_2625,N_2174,N_1725);
or U2626 (N_2626,N_1628,N_1642);
nor U2627 (N_2627,N_1790,N_1674);
or U2628 (N_2628,N_1699,N_1902);
or U2629 (N_2629,N_1820,N_1601);
nand U2630 (N_2630,N_2154,N_1956);
and U2631 (N_2631,N_1789,N_1982);
or U2632 (N_2632,N_1742,N_1557);
and U2633 (N_2633,N_2241,N_1995);
or U2634 (N_2634,N_1966,N_1672);
nand U2635 (N_2635,N_2147,N_1825);
nor U2636 (N_2636,N_2145,N_2161);
and U2637 (N_2637,N_2151,N_2155);
or U2638 (N_2638,N_2186,N_2182);
or U2639 (N_2639,N_2037,N_1623);
or U2640 (N_2640,N_1873,N_2150);
xnor U2641 (N_2641,N_2141,N_1926);
nor U2642 (N_2642,N_2020,N_2119);
and U2643 (N_2643,N_1845,N_2218);
or U2644 (N_2644,N_1506,N_2212);
or U2645 (N_2645,N_1555,N_1808);
xor U2646 (N_2646,N_1980,N_2129);
and U2647 (N_2647,N_1751,N_1931);
nand U2648 (N_2648,N_1666,N_1554);
nor U2649 (N_2649,N_1943,N_1541);
or U2650 (N_2650,N_1631,N_1882);
nand U2651 (N_2651,N_1756,N_2112);
or U2652 (N_2652,N_1710,N_2108);
nand U2653 (N_2653,N_1713,N_1751);
and U2654 (N_2654,N_1609,N_1838);
xnor U2655 (N_2655,N_1575,N_2027);
nor U2656 (N_2656,N_1621,N_1603);
or U2657 (N_2657,N_1581,N_1796);
or U2658 (N_2658,N_2052,N_1608);
nand U2659 (N_2659,N_1529,N_2052);
or U2660 (N_2660,N_1901,N_2171);
and U2661 (N_2661,N_1973,N_1863);
and U2662 (N_2662,N_1852,N_2037);
nor U2663 (N_2663,N_1521,N_1761);
and U2664 (N_2664,N_2169,N_1989);
nor U2665 (N_2665,N_2005,N_1651);
or U2666 (N_2666,N_2137,N_2068);
nor U2667 (N_2667,N_2132,N_1929);
nand U2668 (N_2668,N_1728,N_1533);
or U2669 (N_2669,N_1844,N_1984);
and U2670 (N_2670,N_1671,N_1833);
nand U2671 (N_2671,N_1857,N_1586);
nor U2672 (N_2672,N_2183,N_1720);
or U2673 (N_2673,N_2131,N_2123);
and U2674 (N_2674,N_2132,N_2111);
xor U2675 (N_2675,N_1826,N_1891);
or U2676 (N_2676,N_1750,N_1819);
or U2677 (N_2677,N_1578,N_1762);
nand U2678 (N_2678,N_1996,N_2051);
nor U2679 (N_2679,N_1803,N_2075);
nor U2680 (N_2680,N_1627,N_1711);
xnor U2681 (N_2681,N_1819,N_2046);
nor U2682 (N_2682,N_2194,N_1840);
or U2683 (N_2683,N_2165,N_1628);
and U2684 (N_2684,N_1881,N_1911);
or U2685 (N_2685,N_2037,N_2043);
or U2686 (N_2686,N_2091,N_1648);
and U2687 (N_2687,N_2040,N_1815);
nand U2688 (N_2688,N_1769,N_2172);
nor U2689 (N_2689,N_2176,N_2141);
or U2690 (N_2690,N_1775,N_1658);
xnor U2691 (N_2691,N_1763,N_1976);
nand U2692 (N_2692,N_1540,N_2152);
nand U2693 (N_2693,N_1908,N_2209);
and U2694 (N_2694,N_2084,N_2229);
nand U2695 (N_2695,N_1528,N_1689);
nand U2696 (N_2696,N_1958,N_2167);
and U2697 (N_2697,N_1601,N_2032);
xor U2698 (N_2698,N_1990,N_1920);
nand U2699 (N_2699,N_1631,N_1924);
or U2700 (N_2700,N_1699,N_1874);
and U2701 (N_2701,N_2154,N_2198);
or U2702 (N_2702,N_1719,N_2086);
nor U2703 (N_2703,N_1719,N_2010);
nor U2704 (N_2704,N_1801,N_2072);
nand U2705 (N_2705,N_1777,N_1913);
or U2706 (N_2706,N_2065,N_1797);
and U2707 (N_2707,N_1901,N_1744);
nand U2708 (N_2708,N_1561,N_2123);
or U2709 (N_2709,N_1868,N_1920);
or U2710 (N_2710,N_1858,N_2152);
nand U2711 (N_2711,N_1813,N_1610);
nor U2712 (N_2712,N_1871,N_1793);
and U2713 (N_2713,N_1514,N_1715);
nor U2714 (N_2714,N_1746,N_1638);
nand U2715 (N_2715,N_1680,N_1924);
or U2716 (N_2716,N_1776,N_1821);
nand U2717 (N_2717,N_1587,N_2165);
or U2718 (N_2718,N_2142,N_2060);
nand U2719 (N_2719,N_1798,N_1868);
or U2720 (N_2720,N_1802,N_1825);
nand U2721 (N_2721,N_1527,N_2110);
xnor U2722 (N_2722,N_1911,N_2152);
nor U2723 (N_2723,N_2071,N_1979);
or U2724 (N_2724,N_2205,N_1503);
or U2725 (N_2725,N_1820,N_2214);
or U2726 (N_2726,N_1893,N_2212);
nor U2727 (N_2727,N_1867,N_1693);
and U2728 (N_2728,N_1632,N_2200);
xnor U2729 (N_2729,N_2247,N_1614);
or U2730 (N_2730,N_1584,N_1597);
xor U2731 (N_2731,N_1779,N_2019);
nor U2732 (N_2732,N_1578,N_1990);
or U2733 (N_2733,N_2223,N_1985);
or U2734 (N_2734,N_1591,N_1667);
nand U2735 (N_2735,N_2150,N_1649);
nand U2736 (N_2736,N_2115,N_1511);
xor U2737 (N_2737,N_1780,N_1795);
xnor U2738 (N_2738,N_1562,N_1843);
or U2739 (N_2739,N_1654,N_1567);
or U2740 (N_2740,N_1923,N_1710);
nand U2741 (N_2741,N_1612,N_1836);
or U2742 (N_2742,N_2199,N_1844);
nand U2743 (N_2743,N_1553,N_2244);
xor U2744 (N_2744,N_2174,N_1786);
or U2745 (N_2745,N_1916,N_1723);
and U2746 (N_2746,N_1922,N_1808);
nand U2747 (N_2747,N_1559,N_1570);
or U2748 (N_2748,N_1623,N_1622);
nor U2749 (N_2749,N_1875,N_2118);
nand U2750 (N_2750,N_2058,N_1956);
or U2751 (N_2751,N_2199,N_1634);
nand U2752 (N_2752,N_2055,N_1700);
xnor U2753 (N_2753,N_1646,N_1938);
nand U2754 (N_2754,N_1819,N_1804);
nand U2755 (N_2755,N_1576,N_1641);
nor U2756 (N_2756,N_1815,N_1543);
or U2757 (N_2757,N_1949,N_2134);
or U2758 (N_2758,N_1868,N_2209);
nor U2759 (N_2759,N_1817,N_1988);
nand U2760 (N_2760,N_2090,N_2024);
nor U2761 (N_2761,N_1695,N_1510);
nor U2762 (N_2762,N_1765,N_1543);
or U2763 (N_2763,N_1510,N_1849);
nor U2764 (N_2764,N_2126,N_1960);
and U2765 (N_2765,N_2141,N_1763);
nand U2766 (N_2766,N_1815,N_1732);
nand U2767 (N_2767,N_2032,N_1862);
or U2768 (N_2768,N_1916,N_1614);
and U2769 (N_2769,N_2117,N_2242);
nor U2770 (N_2770,N_2247,N_1957);
nand U2771 (N_2771,N_1887,N_2203);
nand U2772 (N_2772,N_1549,N_1740);
and U2773 (N_2773,N_2070,N_2120);
or U2774 (N_2774,N_1563,N_2050);
nand U2775 (N_2775,N_1717,N_1905);
nor U2776 (N_2776,N_1745,N_1962);
xor U2777 (N_2777,N_1747,N_2145);
nor U2778 (N_2778,N_1766,N_1958);
xor U2779 (N_2779,N_2001,N_2172);
xor U2780 (N_2780,N_1890,N_1589);
nand U2781 (N_2781,N_2117,N_1637);
nand U2782 (N_2782,N_1696,N_1890);
and U2783 (N_2783,N_1696,N_1711);
xnor U2784 (N_2784,N_1724,N_1953);
nand U2785 (N_2785,N_1668,N_1521);
nand U2786 (N_2786,N_1878,N_1658);
or U2787 (N_2787,N_1907,N_2158);
or U2788 (N_2788,N_2241,N_1526);
nor U2789 (N_2789,N_1686,N_1916);
and U2790 (N_2790,N_2001,N_1808);
and U2791 (N_2791,N_2175,N_1743);
nor U2792 (N_2792,N_2011,N_2062);
and U2793 (N_2793,N_1521,N_1800);
and U2794 (N_2794,N_2056,N_2060);
nand U2795 (N_2795,N_2137,N_1721);
nand U2796 (N_2796,N_2195,N_1636);
nor U2797 (N_2797,N_2158,N_2222);
nor U2798 (N_2798,N_1568,N_2046);
and U2799 (N_2799,N_1652,N_1505);
nor U2800 (N_2800,N_1604,N_1990);
or U2801 (N_2801,N_1975,N_1524);
and U2802 (N_2802,N_1554,N_1851);
and U2803 (N_2803,N_1859,N_2031);
nand U2804 (N_2804,N_1820,N_1851);
nand U2805 (N_2805,N_2013,N_2184);
nand U2806 (N_2806,N_1801,N_1677);
xor U2807 (N_2807,N_1688,N_1641);
or U2808 (N_2808,N_1890,N_1699);
xnor U2809 (N_2809,N_1588,N_2029);
nand U2810 (N_2810,N_1952,N_1860);
nand U2811 (N_2811,N_1600,N_2013);
and U2812 (N_2812,N_1918,N_2245);
or U2813 (N_2813,N_1580,N_1860);
nand U2814 (N_2814,N_1560,N_1716);
nand U2815 (N_2815,N_1801,N_2146);
nand U2816 (N_2816,N_2006,N_1923);
nor U2817 (N_2817,N_1794,N_1530);
or U2818 (N_2818,N_1620,N_1783);
or U2819 (N_2819,N_2204,N_1961);
xnor U2820 (N_2820,N_1806,N_2236);
nand U2821 (N_2821,N_1861,N_1537);
or U2822 (N_2822,N_1751,N_1655);
or U2823 (N_2823,N_2243,N_1721);
nand U2824 (N_2824,N_2157,N_2114);
nand U2825 (N_2825,N_1699,N_1504);
and U2826 (N_2826,N_2061,N_1845);
and U2827 (N_2827,N_1789,N_2068);
or U2828 (N_2828,N_1743,N_2236);
and U2829 (N_2829,N_1735,N_2187);
or U2830 (N_2830,N_2224,N_2190);
and U2831 (N_2831,N_2027,N_1814);
xnor U2832 (N_2832,N_1849,N_1848);
and U2833 (N_2833,N_1683,N_2188);
or U2834 (N_2834,N_1949,N_1979);
xor U2835 (N_2835,N_1991,N_1939);
nor U2836 (N_2836,N_2147,N_1951);
nor U2837 (N_2837,N_1587,N_1925);
nand U2838 (N_2838,N_2114,N_1756);
nand U2839 (N_2839,N_1693,N_2162);
or U2840 (N_2840,N_1723,N_2235);
nor U2841 (N_2841,N_1665,N_1600);
or U2842 (N_2842,N_2188,N_2148);
xnor U2843 (N_2843,N_2227,N_1815);
or U2844 (N_2844,N_2185,N_2114);
nand U2845 (N_2845,N_1679,N_2231);
and U2846 (N_2846,N_1878,N_1831);
nand U2847 (N_2847,N_1625,N_1684);
nand U2848 (N_2848,N_1688,N_1716);
xnor U2849 (N_2849,N_2006,N_2035);
xor U2850 (N_2850,N_2181,N_2120);
nor U2851 (N_2851,N_1976,N_1881);
nand U2852 (N_2852,N_2061,N_2184);
or U2853 (N_2853,N_2047,N_1765);
nand U2854 (N_2854,N_2032,N_1724);
nor U2855 (N_2855,N_1535,N_2216);
and U2856 (N_2856,N_2008,N_1514);
or U2857 (N_2857,N_1721,N_1897);
nor U2858 (N_2858,N_2173,N_2116);
or U2859 (N_2859,N_1857,N_2221);
nor U2860 (N_2860,N_2162,N_1655);
and U2861 (N_2861,N_1551,N_1923);
and U2862 (N_2862,N_1678,N_2054);
nor U2863 (N_2863,N_1766,N_1554);
nor U2864 (N_2864,N_2018,N_2044);
nand U2865 (N_2865,N_2214,N_1598);
and U2866 (N_2866,N_1943,N_2156);
nand U2867 (N_2867,N_1701,N_2027);
nor U2868 (N_2868,N_1594,N_2231);
and U2869 (N_2869,N_1500,N_2019);
nand U2870 (N_2870,N_1580,N_2181);
or U2871 (N_2871,N_2090,N_1576);
nand U2872 (N_2872,N_1876,N_1722);
and U2873 (N_2873,N_1741,N_1537);
and U2874 (N_2874,N_1561,N_1935);
and U2875 (N_2875,N_1689,N_1721);
nor U2876 (N_2876,N_1537,N_2136);
nor U2877 (N_2877,N_1880,N_2227);
and U2878 (N_2878,N_1862,N_1576);
xnor U2879 (N_2879,N_1681,N_1858);
nand U2880 (N_2880,N_1806,N_2132);
nand U2881 (N_2881,N_2031,N_1567);
and U2882 (N_2882,N_1878,N_2192);
or U2883 (N_2883,N_1997,N_1730);
nand U2884 (N_2884,N_2206,N_2012);
xnor U2885 (N_2885,N_2054,N_2147);
or U2886 (N_2886,N_1530,N_1781);
and U2887 (N_2887,N_1645,N_2099);
and U2888 (N_2888,N_1949,N_2015);
nor U2889 (N_2889,N_2164,N_1607);
or U2890 (N_2890,N_1515,N_1537);
nor U2891 (N_2891,N_1689,N_1895);
and U2892 (N_2892,N_1921,N_1764);
xor U2893 (N_2893,N_1984,N_1602);
nor U2894 (N_2894,N_1894,N_1775);
and U2895 (N_2895,N_1856,N_2014);
or U2896 (N_2896,N_2238,N_2163);
or U2897 (N_2897,N_1977,N_1764);
or U2898 (N_2898,N_2039,N_1769);
and U2899 (N_2899,N_1542,N_2183);
or U2900 (N_2900,N_1886,N_1517);
xor U2901 (N_2901,N_1517,N_2181);
and U2902 (N_2902,N_1528,N_1524);
or U2903 (N_2903,N_1828,N_1776);
xnor U2904 (N_2904,N_2156,N_2085);
and U2905 (N_2905,N_1525,N_2236);
nand U2906 (N_2906,N_1533,N_1612);
or U2907 (N_2907,N_1820,N_1714);
nor U2908 (N_2908,N_1553,N_1876);
nor U2909 (N_2909,N_2190,N_1501);
and U2910 (N_2910,N_1932,N_2073);
and U2911 (N_2911,N_1634,N_2170);
nor U2912 (N_2912,N_2181,N_1769);
or U2913 (N_2913,N_2223,N_1757);
and U2914 (N_2914,N_1579,N_1545);
nand U2915 (N_2915,N_1577,N_2081);
and U2916 (N_2916,N_1660,N_2102);
and U2917 (N_2917,N_2111,N_1575);
and U2918 (N_2918,N_2218,N_1515);
or U2919 (N_2919,N_1526,N_1681);
nor U2920 (N_2920,N_2068,N_2193);
xnor U2921 (N_2921,N_1706,N_1622);
and U2922 (N_2922,N_2134,N_2141);
nor U2923 (N_2923,N_2216,N_1716);
and U2924 (N_2924,N_1978,N_1860);
xor U2925 (N_2925,N_1525,N_1757);
nor U2926 (N_2926,N_1626,N_1848);
and U2927 (N_2927,N_2243,N_1910);
or U2928 (N_2928,N_2179,N_1774);
nand U2929 (N_2929,N_1853,N_2202);
and U2930 (N_2930,N_1807,N_1885);
nand U2931 (N_2931,N_2045,N_1515);
nor U2932 (N_2932,N_2129,N_1839);
or U2933 (N_2933,N_1845,N_1930);
xor U2934 (N_2934,N_2041,N_1599);
xnor U2935 (N_2935,N_1601,N_1808);
nor U2936 (N_2936,N_1675,N_1591);
nor U2937 (N_2937,N_1545,N_2004);
nor U2938 (N_2938,N_1726,N_1824);
nand U2939 (N_2939,N_1692,N_1524);
xor U2940 (N_2940,N_1992,N_1795);
and U2941 (N_2941,N_1869,N_1588);
nor U2942 (N_2942,N_1505,N_2169);
nand U2943 (N_2943,N_1555,N_2142);
nand U2944 (N_2944,N_1981,N_1581);
or U2945 (N_2945,N_2186,N_1938);
nand U2946 (N_2946,N_1777,N_1654);
nand U2947 (N_2947,N_1582,N_1789);
and U2948 (N_2948,N_2170,N_1565);
nor U2949 (N_2949,N_2104,N_2032);
nand U2950 (N_2950,N_1555,N_1531);
nand U2951 (N_2951,N_2043,N_1831);
nand U2952 (N_2952,N_2017,N_1887);
or U2953 (N_2953,N_2219,N_2232);
or U2954 (N_2954,N_2103,N_1692);
or U2955 (N_2955,N_1798,N_2172);
nor U2956 (N_2956,N_1589,N_2179);
and U2957 (N_2957,N_1789,N_1934);
nand U2958 (N_2958,N_1782,N_1958);
xor U2959 (N_2959,N_1647,N_1940);
nand U2960 (N_2960,N_2043,N_1779);
and U2961 (N_2961,N_1791,N_2249);
xnor U2962 (N_2962,N_2017,N_2232);
nand U2963 (N_2963,N_2159,N_2070);
nor U2964 (N_2964,N_1542,N_1666);
and U2965 (N_2965,N_1514,N_1535);
nor U2966 (N_2966,N_1696,N_1947);
or U2967 (N_2967,N_1815,N_1590);
and U2968 (N_2968,N_1790,N_2170);
or U2969 (N_2969,N_1970,N_2247);
and U2970 (N_2970,N_2033,N_1655);
nor U2971 (N_2971,N_1719,N_1762);
or U2972 (N_2972,N_1658,N_1571);
nand U2973 (N_2973,N_2236,N_1998);
nand U2974 (N_2974,N_1931,N_1563);
nor U2975 (N_2975,N_2132,N_1747);
nand U2976 (N_2976,N_1557,N_2085);
or U2977 (N_2977,N_1561,N_1889);
and U2978 (N_2978,N_1686,N_1832);
and U2979 (N_2979,N_1793,N_1557);
nand U2980 (N_2980,N_2044,N_1695);
or U2981 (N_2981,N_2071,N_2173);
xor U2982 (N_2982,N_1531,N_1928);
xor U2983 (N_2983,N_1690,N_1902);
xor U2984 (N_2984,N_1938,N_1589);
or U2985 (N_2985,N_1940,N_2157);
and U2986 (N_2986,N_1884,N_1622);
nand U2987 (N_2987,N_1602,N_1760);
nor U2988 (N_2988,N_1860,N_2124);
nor U2989 (N_2989,N_1552,N_2161);
or U2990 (N_2990,N_1688,N_1827);
nor U2991 (N_2991,N_1846,N_2231);
nand U2992 (N_2992,N_2108,N_2208);
and U2993 (N_2993,N_2063,N_1530);
and U2994 (N_2994,N_1788,N_2247);
or U2995 (N_2995,N_1899,N_1800);
and U2996 (N_2996,N_1680,N_1928);
and U2997 (N_2997,N_1592,N_1612);
and U2998 (N_2998,N_1946,N_2046);
xnor U2999 (N_2999,N_1745,N_1560);
nor U3000 (N_3000,N_2506,N_2325);
nor U3001 (N_3001,N_2756,N_2768);
xnor U3002 (N_3002,N_2332,N_2329);
and U3003 (N_3003,N_2645,N_2790);
nor U3004 (N_3004,N_2922,N_2838);
nand U3005 (N_3005,N_2599,N_2615);
or U3006 (N_3006,N_2289,N_2327);
nand U3007 (N_3007,N_2356,N_2488);
or U3008 (N_3008,N_2914,N_2284);
and U3009 (N_3009,N_2633,N_2830);
or U3010 (N_3010,N_2871,N_2405);
and U3011 (N_3011,N_2279,N_2341);
nor U3012 (N_3012,N_2354,N_2555);
and U3013 (N_3013,N_2557,N_2545);
nor U3014 (N_3014,N_2779,N_2292);
and U3015 (N_3015,N_2607,N_2932);
and U3016 (N_3016,N_2981,N_2268);
nor U3017 (N_3017,N_2259,N_2643);
nor U3018 (N_3018,N_2467,N_2847);
nor U3019 (N_3019,N_2589,N_2305);
and U3020 (N_3020,N_2269,N_2721);
nor U3021 (N_3021,N_2996,N_2631);
and U3022 (N_3022,N_2666,N_2478);
and U3023 (N_3023,N_2926,N_2740);
nand U3024 (N_3024,N_2373,N_2472);
nand U3025 (N_3025,N_2972,N_2919);
and U3026 (N_3026,N_2445,N_2497);
nand U3027 (N_3027,N_2888,N_2784);
or U3028 (N_3028,N_2890,N_2808);
or U3029 (N_3029,N_2852,N_2858);
nand U3030 (N_3030,N_2788,N_2308);
nor U3031 (N_3031,N_2767,N_2271);
or U3032 (N_3032,N_2664,N_2530);
or U3033 (N_3033,N_2343,N_2860);
nand U3034 (N_3034,N_2939,N_2892);
or U3035 (N_3035,N_2413,N_2464);
or U3036 (N_3036,N_2693,N_2263);
nor U3037 (N_3037,N_2920,N_2391);
nand U3038 (N_3038,N_2969,N_2657);
nor U3039 (N_3039,N_2782,N_2274);
or U3040 (N_3040,N_2569,N_2570);
or U3041 (N_3041,N_2702,N_2764);
or U3042 (N_3042,N_2436,N_2821);
nor U3043 (N_3043,N_2708,N_2621);
nor U3044 (N_3044,N_2603,N_2825);
nand U3045 (N_3045,N_2287,N_2965);
nand U3046 (N_3046,N_2612,N_2850);
and U3047 (N_3047,N_2966,N_2805);
nor U3048 (N_3048,N_2519,N_2826);
and U3049 (N_3049,N_2902,N_2425);
nor U3050 (N_3050,N_2995,N_2711);
nor U3051 (N_3051,N_2617,N_2558);
or U3052 (N_3052,N_2339,N_2994);
nor U3053 (N_3053,N_2820,N_2430);
nor U3054 (N_3054,N_2353,N_2251);
and U3055 (N_3055,N_2574,N_2345);
or U3056 (N_3056,N_2604,N_2900);
xnor U3057 (N_3057,N_2931,N_2309);
nor U3058 (N_3058,N_2508,N_2526);
nand U3059 (N_3059,N_2416,N_2677);
and U3060 (N_3060,N_2917,N_2550);
nand U3061 (N_3061,N_2444,N_2845);
nand U3062 (N_3062,N_2906,N_2322);
nand U3063 (N_3063,N_2691,N_2781);
nand U3064 (N_3064,N_2567,N_2727);
and U3065 (N_3065,N_2722,N_2682);
nor U3066 (N_3066,N_2465,N_2371);
or U3067 (N_3067,N_2815,N_2359);
or U3068 (N_3068,N_2831,N_2446);
xnor U3069 (N_3069,N_2809,N_2449);
or U3070 (N_3070,N_2773,N_2774);
nor U3071 (N_3071,N_2819,N_2522);
nor U3072 (N_3072,N_2877,N_2726);
and U3073 (N_3073,N_2568,N_2429);
nand U3074 (N_3074,N_2584,N_2523);
and U3075 (N_3075,N_2964,N_2793);
and U3076 (N_3076,N_2894,N_2942);
nand U3077 (N_3077,N_2739,N_2576);
or U3078 (N_3078,N_2806,N_2870);
or U3079 (N_3079,N_2447,N_2915);
and U3080 (N_3080,N_2907,N_2281);
or U3081 (N_3081,N_2559,N_2629);
nor U3082 (N_3082,N_2531,N_2843);
or U3083 (N_3083,N_2623,N_2672);
nor U3084 (N_3084,N_2921,N_2959);
nand U3085 (N_3085,N_2505,N_2383);
xor U3086 (N_3086,N_2823,N_2544);
nor U3087 (N_3087,N_2392,N_2620);
or U3088 (N_3088,N_2312,N_2285);
xnor U3089 (N_3089,N_2338,N_2386);
nand U3090 (N_3090,N_2792,N_2524);
and U3091 (N_3091,N_2419,N_2798);
xnor U3092 (N_3092,N_2466,N_2833);
nor U3093 (N_3093,N_2968,N_2539);
nor U3094 (N_3094,N_2647,N_2262);
nand U3095 (N_3095,N_2634,N_2290);
or U3096 (N_3096,N_2818,N_2750);
and U3097 (N_3097,N_2801,N_2554);
and U3098 (N_3098,N_2415,N_2389);
and U3099 (N_3099,N_2717,N_2882);
nand U3100 (N_3100,N_2546,N_2492);
nand U3101 (N_3101,N_2883,N_2283);
or U3102 (N_3102,N_2837,N_2667);
or U3103 (N_3103,N_2998,N_2605);
or U3104 (N_3104,N_2802,N_2443);
and U3105 (N_3105,N_2491,N_2674);
nand U3106 (N_3106,N_2680,N_2730);
nand U3107 (N_3107,N_2957,N_2493);
nor U3108 (N_3108,N_2639,N_2381);
nand U3109 (N_3109,N_2849,N_2579);
and U3110 (N_3110,N_2736,N_2291);
nand U3111 (N_3111,N_2282,N_2923);
nor U3112 (N_3112,N_2362,N_2898);
or U3113 (N_3113,N_2899,N_2310);
or U3114 (N_3114,N_2328,N_2538);
nand U3115 (N_3115,N_2804,N_2824);
nand U3116 (N_3116,N_2699,N_2908);
or U3117 (N_3117,N_2575,N_2811);
nor U3118 (N_3118,N_2650,N_2712);
xnor U3119 (N_3119,N_2771,N_2697);
nor U3120 (N_3120,N_2953,N_2384);
nand U3121 (N_3121,N_2766,N_2857);
nor U3122 (N_3122,N_2377,N_2580);
nor U3123 (N_3123,N_2844,N_2810);
nand U3124 (N_3124,N_2380,N_2961);
nand U3125 (N_3125,N_2897,N_2397);
or U3126 (N_3126,N_2746,N_2765);
nand U3127 (N_3127,N_2601,N_2885);
nand U3128 (N_3128,N_2927,N_2758);
nor U3129 (N_3129,N_2757,N_2695);
nor U3130 (N_3130,N_2912,N_2970);
xnor U3131 (N_3131,N_2542,N_2496);
or U3132 (N_3132,N_2935,N_2709);
or U3133 (N_3133,N_2433,N_2437);
xnor U3134 (N_3134,N_2363,N_2839);
xor U3135 (N_3135,N_2280,N_2533);
or U3136 (N_3136,N_2264,N_2979);
and U3137 (N_3137,N_2404,N_2668);
or U3138 (N_3138,N_2596,N_2720);
or U3139 (N_3139,N_2461,N_2817);
xnor U3140 (N_3140,N_2333,N_2591);
nor U3141 (N_3141,N_2340,N_2909);
and U3142 (N_3142,N_2762,N_2528);
nor U3143 (N_3143,N_2592,N_2307);
xnor U3144 (N_3144,N_2412,N_2684);
nand U3145 (N_3145,N_2370,N_2347);
and U3146 (N_3146,N_2342,N_2257);
nand U3147 (N_3147,N_2618,N_2454);
and U3148 (N_3148,N_2301,N_2753);
nand U3149 (N_3149,N_2813,N_2626);
nor U3150 (N_3150,N_2770,N_2648);
or U3151 (N_3151,N_2611,N_2663);
or U3152 (N_3152,N_2613,N_2848);
and U3153 (N_3153,N_2669,N_2432);
nand U3154 (N_3154,N_2532,N_2982);
and U3155 (N_3155,N_2375,N_2480);
and U3156 (N_3156,N_2933,N_2946);
or U3157 (N_3157,N_2686,N_2481);
and U3158 (N_3158,N_2518,N_2660);
xor U3159 (N_3159,N_2457,N_2929);
and U3160 (N_3160,N_2703,N_2266);
or U3161 (N_3161,N_2253,N_2427);
nand U3162 (N_3162,N_2265,N_2759);
nor U3163 (N_3163,N_2398,N_2423);
xnor U3164 (N_3164,N_2500,N_2675);
nor U3165 (N_3165,N_2529,N_2896);
and U3166 (N_3166,N_2962,N_2256);
nor U3167 (N_3167,N_2955,N_2318);
nand U3168 (N_3168,N_2350,N_2975);
or U3169 (N_3169,N_2477,N_2878);
and U3170 (N_3170,N_2807,N_2780);
or U3171 (N_3171,N_2600,N_2346);
or U3172 (N_3172,N_2864,N_2330);
or U3173 (N_3173,N_2978,N_2842);
nor U3174 (N_3174,N_2796,N_2448);
or U3175 (N_3175,N_2938,N_2832);
nor U3176 (N_3176,N_2960,N_2549);
and U3177 (N_3177,N_2479,N_2989);
nand U3178 (N_3178,N_2595,N_2597);
nor U3179 (N_3179,N_2988,N_2869);
or U3180 (N_3180,N_2853,N_2999);
xnor U3181 (N_3181,N_2361,N_2936);
nor U3182 (N_3182,N_2434,N_2930);
or U3183 (N_3183,N_2344,N_2872);
nor U3184 (N_3184,N_2315,N_2886);
xnor U3185 (N_3185,N_2879,N_2521);
nor U3186 (N_3186,N_2747,N_2656);
and U3187 (N_3187,N_2904,N_2484);
or U3188 (N_3188,N_2928,N_2856);
and U3189 (N_3189,N_2321,N_2945);
nor U3190 (N_3190,N_2816,N_2822);
nor U3191 (N_3191,N_2512,N_2352);
nor U3192 (N_3192,N_2777,N_2934);
xor U3193 (N_3193,N_2385,N_2619);
xnor U3194 (N_3194,N_2867,N_2608);
nor U3195 (N_3195,N_2622,N_2561);
and U3196 (N_3196,N_2442,N_2649);
nand U3197 (N_3197,N_2803,N_2566);
or U3198 (N_3198,N_2763,N_2258);
nand U3199 (N_3199,N_2772,N_2379);
nand U3200 (N_3200,N_2889,N_2866);
nand U3201 (N_3201,N_2951,N_2735);
xnor U3202 (N_3202,N_2458,N_2646);
nand U3203 (N_3203,N_2299,N_2737);
nand U3204 (N_3204,N_2723,N_2644);
nand U3205 (N_3205,N_2336,N_2452);
nand U3206 (N_3206,N_2653,N_2725);
nor U3207 (N_3207,N_2714,N_2536);
or U3208 (N_3208,N_2367,N_2502);
or U3209 (N_3209,N_2630,N_2468);
or U3210 (N_3210,N_2873,N_2827);
xor U3211 (N_3211,N_2859,N_2992);
or U3212 (N_3212,N_2625,N_2628);
and U3213 (N_3213,N_2571,N_2698);
nand U3214 (N_3214,N_2455,N_2688);
and U3215 (N_3215,N_2991,N_2689);
and U3216 (N_3216,N_2378,N_2734);
and U3217 (N_3217,N_2537,N_2658);
and U3218 (N_3218,N_2351,N_2731);
or U3219 (N_3219,N_2394,N_2577);
nand U3220 (N_3220,N_2627,N_2700);
or U3221 (N_3221,N_2562,N_2276);
or U3222 (N_3222,N_2706,N_2286);
nor U3223 (N_3223,N_2509,N_2901);
nand U3224 (N_3224,N_2854,N_2453);
or U3225 (N_3225,N_2498,N_2511);
or U3226 (N_3226,N_2947,N_2704);
or U3227 (N_3227,N_2475,N_2918);
nor U3228 (N_3228,N_2593,N_2884);
nand U3229 (N_3229,N_2635,N_2729);
or U3230 (N_3230,N_2260,N_2364);
nand U3231 (N_3231,N_2895,N_2642);
and U3232 (N_3232,N_2761,N_2516);
nor U3233 (N_3233,N_2977,N_2993);
and U3234 (N_3234,N_2690,N_2463);
or U3235 (N_3235,N_2952,N_2297);
and U3236 (N_3236,N_2738,N_2705);
and U3237 (N_3237,N_2659,N_2598);
nand U3238 (N_3238,N_2451,N_2250);
xor U3239 (N_3239,N_2937,N_2293);
nor U3240 (N_3240,N_2482,N_2624);
xor U3241 (N_3241,N_2476,N_2535);
nor U3242 (N_3242,N_2581,N_2679);
xor U3243 (N_3243,N_2718,N_2426);
and U3244 (N_3244,N_2973,N_2469);
and U3245 (N_3245,N_2984,N_2582);
and U3246 (N_3246,N_2948,N_2585);
and U3247 (N_3247,N_2829,N_2944);
or U3248 (N_3248,N_2489,N_2670);
xor U3249 (N_3249,N_2317,N_2462);
and U3250 (N_3250,N_2606,N_2846);
or U3251 (N_3251,N_2754,N_2812);
xnor U3252 (N_3252,N_2349,N_2610);
xor U3253 (N_3253,N_2671,N_2525);
and U3254 (N_3254,N_2678,N_2278);
or U3255 (N_3255,N_2683,N_2594);
nand U3256 (N_3256,N_2514,N_2971);
nand U3257 (N_3257,N_2685,N_2785);
or U3258 (N_3258,N_2835,N_2696);
and U3259 (N_3259,N_2775,N_2715);
and U3260 (N_3260,N_2387,N_2910);
nor U3261 (N_3261,N_2424,N_2641);
and U3262 (N_3262,N_2547,N_2428);
or U3263 (N_3263,N_2980,N_2368);
or U3264 (N_3264,N_2862,N_2323);
and U3265 (N_3265,N_2787,N_2602);
or U3266 (N_3266,N_2751,N_2943);
and U3267 (N_3267,N_2662,N_2441);
nor U3268 (N_3268,N_2490,N_2913);
nand U3269 (N_3269,N_2795,N_2541);
nor U3270 (N_3270,N_2778,N_2540);
nand U3271 (N_3271,N_2302,N_2732);
nand U3272 (N_3272,N_2789,N_2572);
or U3273 (N_3273,N_2654,N_2288);
nand U3274 (N_3274,N_2507,N_2431);
or U3275 (N_3275,N_2252,N_2314);
nor U3276 (N_3276,N_2728,N_2861);
nand U3277 (N_3277,N_2422,N_2485);
nor U3278 (N_3278,N_2661,N_2316);
and U3279 (N_3279,N_2483,N_2390);
or U3280 (N_3280,N_2504,N_2865);
nand U3281 (N_3281,N_2421,N_2553);
and U3282 (N_3282,N_2355,N_2471);
and U3283 (N_3283,N_2438,N_2296);
or U3284 (N_3284,N_2494,N_2456);
nand U3285 (N_3285,N_2655,N_2609);
and U3286 (N_3286,N_2941,N_2949);
nand U3287 (N_3287,N_2408,N_2313);
or U3288 (N_3288,N_2275,N_2640);
nor U3289 (N_3289,N_2828,N_2724);
nand U3290 (N_3290,N_2956,N_2543);
and U3291 (N_3291,N_2573,N_2836);
and U3292 (N_3292,N_2255,N_2578);
xnor U3293 (N_3293,N_2414,N_2636);
nor U3294 (N_3294,N_2474,N_2783);
and U3295 (N_3295,N_2513,N_2755);
or U3296 (N_3296,N_2517,N_2406);
and U3297 (N_3297,N_2834,N_2303);
or U3298 (N_3298,N_2967,N_2748);
or U3299 (N_3299,N_2319,N_2687);
nor U3300 (N_3300,N_2743,N_2916);
nor U3301 (N_3301,N_2337,N_2254);
and U3302 (N_3302,N_2924,N_2560);
or U3303 (N_3303,N_2940,N_2749);
or U3304 (N_3304,N_2963,N_2791);
and U3305 (N_3305,N_2331,N_2794);
and U3306 (N_3306,N_2410,N_2388);
and U3307 (N_3307,N_2357,N_2903);
nor U3308 (N_3308,N_2893,N_2399);
nor U3309 (N_3309,N_2395,N_2365);
xnor U3310 (N_3310,N_2692,N_2614);
or U3311 (N_3311,N_2974,N_2334);
and U3312 (N_3312,N_2745,N_2769);
or U3313 (N_3313,N_2501,N_2814);
xor U3314 (N_3314,N_2588,N_2719);
and U3315 (N_3315,N_2707,N_2986);
xor U3316 (N_3316,N_2417,N_2887);
or U3317 (N_3317,N_2744,N_2273);
or U3318 (N_3318,N_2440,N_2710);
or U3319 (N_3319,N_2905,N_2551);
or U3320 (N_3320,N_2372,N_2470);
and U3321 (N_3321,N_2997,N_2976);
and U3322 (N_3322,N_2407,N_2374);
or U3323 (N_3323,N_2376,N_2632);
nor U3324 (N_3324,N_2358,N_2401);
nor U3325 (N_3325,N_2676,N_2786);
or U3326 (N_3326,N_2925,N_2486);
and U3327 (N_3327,N_2270,N_2515);
nand U3328 (N_3328,N_2335,N_2295);
or U3329 (N_3329,N_2741,N_2420);
nor U3330 (N_3330,N_2300,N_2400);
nor U3331 (N_3331,N_2393,N_2495);
or U3332 (N_3332,N_2418,N_2348);
or U3333 (N_3333,N_2510,N_2760);
nand U3334 (N_3334,N_2713,N_2681);
nor U3335 (N_3335,N_2587,N_2435);
nand U3336 (N_3336,N_2651,N_2366);
nor U3337 (N_3337,N_2797,N_2586);
and U3338 (N_3338,N_2564,N_2563);
nand U3339 (N_3339,N_2637,N_2851);
or U3340 (N_3340,N_2460,N_2742);
and U3341 (N_3341,N_2985,N_2396);
and U3342 (N_3342,N_2776,N_2868);
or U3343 (N_3343,N_2459,N_2439);
nand U3344 (N_3344,N_2527,N_2382);
nor U3345 (N_3345,N_2548,N_2841);
or U3346 (N_3346,N_2911,N_2590);
nor U3347 (N_3347,N_2320,N_2616);
or U3348 (N_3348,N_2298,N_2450);
and U3349 (N_3349,N_2473,N_2369);
xor U3350 (N_3350,N_2499,N_2294);
or U3351 (N_3351,N_2881,N_2673);
or U3352 (N_3352,N_2277,N_2503);
nor U3353 (N_3353,N_2520,N_2487);
and U3354 (N_3354,N_2272,N_2950);
nor U3355 (N_3355,N_2733,N_2752);
nand U3356 (N_3356,N_2261,N_2652);
nand U3357 (N_3357,N_2326,N_2583);
or U3358 (N_3358,N_2306,N_2311);
nand U3359 (N_3359,N_2409,N_2987);
nand U3360 (N_3360,N_2876,N_2875);
or U3361 (N_3361,N_2701,N_2565);
nor U3362 (N_3362,N_2799,N_2411);
nor U3363 (N_3363,N_2360,N_2855);
nor U3364 (N_3364,N_2638,N_2304);
nand U3365 (N_3365,N_2874,N_2403);
or U3366 (N_3366,N_2556,N_2800);
nand U3367 (N_3367,N_2534,N_2267);
nand U3368 (N_3368,N_2840,N_2716);
xor U3369 (N_3369,N_2402,N_2891);
or U3370 (N_3370,N_2552,N_2665);
xnor U3371 (N_3371,N_2863,N_2983);
nor U3372 (N_3372,N_2880,N_2954);
nand U3373 (N_3373,N_2694,N_2990);
or U3374 (N_3374,N_2324,N_2958);
xor U3375 (N_3375,N_2660,N_2705);
nand U3376 (N_3376,N_2710,N_2362);
nand U3377 (N_3377,N_2725,N_2920);
xnor U3378 (N_3378,N_2934,N_2699);
nor U3379 (N_3379,N_2717,N_2366);
or U3380 (N_3380,N_2829,N_2374);
nor U3381 (N_3381,N_2273,N_2518);
and U3382 (N_3382,N_2357,N_2800);
nor U3383 (N_3383,N_2880,N_2743);
or U3384 (N_3384,N_2546,N_2253);
and U3385 (N_3385,N_2694,N_2812);
xor U3386 (N_3386,N_2643,N_2874);
or U3387 (N_3387,N_2668,N_2706);
or U3388 (N_3388,N_2350,N_2751);
nand U3389 (N_3389,N_2656,N_2978);
nand U3390 (N_3390,N_2833,N_2288);
nand U3391 (N_3391,N_2608,N_2421);
or U3392 (N_3392,N_2465,N_2756);
nand U3393 (N_3393,N_2797,N_2884);
nand U3394 (N_3394,N_2800,N_2891);
nor U3395 (N_3395,N_2725,N_2926);
and U3396 (N_3396,N_2999,N_2504);
nor U3397 (N_3397,N_2299,N_2496);
nor U3398 (N_3398,N_2736,N_2250);
nand U3399 (N_3399,N_2731,N_2455);
and U3400 (N_3400,N_2952,N_2352);
nor U3401 (N_3401,N_2326,N_2794);
nor U3402 (N_3402,N_2276,N_2659);
or U3403 (N_3403,N_2258,N_2287);
or U3404 (N_3404,N_2733,N_2580);
nor U3405 (N_3405,N_2421,N_2517);
and U3406 (N_3406,N_2783,N_2718);
and U3407 (N_3407,N_2507,N_2797);
nor U3408 (N_3408,N_2826,N_2313);
and U3409 (N_3409,N_2842,N_2781);
nor U3410 (N_3410,N_2775,N_2627);
and U3411 (N_3411,N_2470,N_2534);
nor U3412 (N_3412,N_2339,N_2900);
and U3413 (N_3413,N_2723,N_2633);
and U3414 (N_3414,N_2262,N_2871);
nor U3415 (N_3415,N_2661,N_2967);
or U3416 (N_3416,N_2888,N_2487);
nor U3417 (N_3417,N_2730,N_2455);
xor U3418 (N_3418,N_2284,N_2884);
nor U3419 (N_3419,N_2608,N_2488);
nor U3420 (N_3420,N_2838,N_2523);
nand U3421 (N_3421,N_2809,N_2839);
nor U3422 (N_3422,N_2917,N_2924);
nor U3423 (N_3423,N_2482,N_2502);
nand U3424 (N_3424,N_2836,N_2739);
nand U3425 (N_3425,N_2522,N_2583);
nand U3426 (N_3426,N_2694,N_2497);
nor U3427 (N_3427,N_2790,N_2782);
nor U3428 (N_3428,N_2521,N_2618);
nor U3429 (N_3429,N_2676,N_2312);
or U3430 (N_3430,N_2948,N_2265);
and U3431 (N_3431,N_2752,N_2795);
xor U3432 (N_3432,N_2805,N_2419);
nor U3433 (N_3433,N_2587,N_2304);
nor U3434 (N_3434,N_2460,N_2411);
nand U3435 (N_3435,N_2854,N_2702);
and U3436 (N_3436,N_2753,N_2276);
nor U3437 (N_3437,N_2469,N_2390);
and U3438 (N_3438,N_2786,N_2749);
nand U3439 (N_3439,N_2725,N_2959);
xor U3440 (N_3440,N_2779,N_2879);
or U3441 (N_3441,N_2729,N_2341);
or U3442 (N_3442,N_2382,N_2908);
or U3443 (N_3443,N_2705,N_2786);
and U3444 (N_3444,N_2336,N_2836);
nor U3445 (N_3445,N_2690,N_2448);
nor U3446 (N_3446,N_2613,N_2997);
and U3447 (N_3447,N_2875,N_2641);
xnor U3448 (N_3448,N_2438,N_2385);
xor U3449 (N_3449,N_2922,N_2846);
or U3450 (N_3450,N_2851,N_2610);
and U3451 (N_3451,N_2632,N_2477);
or U3452 (N_3452,N_2726,N_2973);
or U3453 (N_3453,N_2384,N_2562);
nand U3454 (N_3454,N_2375,N_2670);
nand U3455 (N_3455,N_2777,N_2282);
nor U3456 (N_3456,N_2439,N_2569);
or U3457 (N_3457,N_2821,N_2850);
nand U3458 (N_3458,N_2966,N_2799);
or U3459 (N_3459,N_2438,N_2810);
xnor U3460 (N_3460,N_2348,N_2747);
and U3461 (N_3461,N_2763,N_2467);
nand U3462 (N_3462,N_2559,N_2688);
nor U3463 (N_3463,N_2695,N_2787);
or U3464 (N_3464,N_2788,N_2589);
and U3465 (N_3465,N_2746,N_2953);
or U3466 (N_3466,N_2369,N_2443);
and U3467 (N_3467,N_2775,N_2582);
or U3468 (N_3468,N_2449,N_2726);
nor U3469 (N_3469,N_2840,N_2906);
nor U3470 (N_3470,N_2287,N_2492);
nor U3471 (N_3471,N_2416,N_2714);
nor U3472 (N_3472,N_2983,N_2847);
or U3473 (N_3473,N_2550,N_2379);
or U3474 (N_3474,N_2266,N_2647);
xnor U3475 (N_3475,N_2586,N_2732);
or U3476 (N_3476,N_2926,N_2692);
or U3477 (N_3477,N_2947,N_2528);
and U3478 (N_3478,N_2895,N_2347);
or U3479 (N_3479,N_2491,N_2935);
nand U3480 (N_3480,N_2612,N_2536);
nand U3481 (N_3481,N_2619,N_2861);
nor U3482 (N_3482,N_2912,N_2752);
or U3483 (N_3483,N_2456,N_2997);
nand U3484 (N_3484,N_2635,N_2961);
nor U3485 (N_3485,N_2350,N_2908);
and U3486 (N_3486,N_2591,N_2969);
or U3487 (N_3487,N_2381,N_2445);
or U3488 (N_3488,N_2477,N_2381);
or U3489 (N_3489,N_2276,N_2501);
nor U3490 (N_3490,N_2518,N_2910);
or U3491 (N_3491,N_2441,N_2348);
or U3492 (N_3492,N_2347,N_2628);
xnor U3493 (N_3493,N_2780,N_2281);
nor U3494 (N_3494,N_2746,N_2847);
nand U3495 (N_3495,N_2496,N_2607);
nor U3496 (N_3496,N_2872,N_2361);
and U3497 (N_3497,N_2354,N_2320);
nand U3498 (N_3498,N_2449,N_2306);
and U3499 (N_3499,N_2774,N_2500);
and U3500 (N_3500,N_2908,N_2493);
or U3501 (N_3501,N_2609,N_2941);
or U3502 (N_3502,N_2719,N_2850);
and U3503 (N_3503,N_2655,N_2639);
nand U3504 (N_3504,N_2706,N_2648);
nor U3505 (N_3505,N_2655,N_2632);
or U3506 (N_3506,N_2892,N_2544);
nand U3507 (N_3507,N_2470,N_2556);
and U3508 (N_3508,N_2475,N_2660);
nor U3509 (N_3509,N_2255,N_2884);
nand U3510 (N_3510,N_2495,N_2713);
and U3511 (N_3511,N_2514,N_2917);
or U3512 (N_3512,N_2454,N_2748);
and U3513 (N_3513,N_2271,N_2666);
nand U3514 (N_3514,N_2279,N_2614);
nor U3515 (N_3515,N_2609,N_2560);
nand U3516 (N_3516,N_2984,N_2725);
and U3517 (N_3517,N_2474,N_2308);
nor U3518 (N_3518,N_2482,N_2619);
nor U3519 (N_3519,N_2814,N_2987);
or U3520 (N_3520,N_2261,N_2998);
nor U3521 (N_3521,N_2656,N_2378);
and U3522 (N_3522,N_2772,N_2745);
or U3523 (N_3523,N_2613,N_2638);
nor U3524 (N_3524,N_2643,N_2377);
xor U3525 (N_3525,N_2365,N_2350);
nor U3526 (N_3526,N_2310,N_2439);
and U3527 (N_3527,N_2980,N_2785);
or U3528 (N_3528,N_2678,N_2549);
or U3529 (N_3529,N_2512,N_2918);
nor U3530 (N_3530,N_2632,N_2796);
nor U3531 (N_3531,N_2671,N_2418);
and U3532 (N_3532,N_2730,N_2665);
nand U3533 (N_3533,N_2307,N_2396);
nand U3534 (N_3534,N_2295,N_2488);
nand U3535 (N_3535,N_2309,N_2886);
nand U3536 (N_3536,N_2874,N_2671);
nand U3537 (N_3537,N_2358,N_2490);
nand U3538 (N_3538,N_2642,N_2464);
nor U3539 (N_3539,N_2543,N_2334);
or U3540 (N_3540,N_2843,N_2372);
nor U3541 (N_3541,N_2495,N_2636);
nand U3542 (N_3542,N_2499,N_2937);
nand U3543 (N_3543,N_2495,N_2453);
nor U3544 (N_3544,N_2542,N_2663);
and U3545 (N_3545,N_2789,N_2911);
nor U3546 (N_3546,N_2528,N_2491);
xor U3547 (N_3547,N_2880,N_2998);
nor U3548 (N_3548,N_2620,N_2708);
nor U3549 (N_3549,N_2785,N_2891);
or U3550 (N_3550,N_2747,N_2571);
or U3551 (N_3551,N_2349,N_2884);
or U3552 (N_3552,N_2579,N_2279);
and U3553 (N_3553,N_2444,N_2269);
nand U3554 (N_3554,N_2899,N_2957);
nand U3555 (N_3555,N_2473,N_2440);
or U3556 (N_3556,N_2990,N_2759);
and U3557 (N_3557,N_2946,N_2581);
xor U3558 (N_3558,N_2411,N_2478);
nand U3559 (N_3559,N_2462,N_2269);
and U3560 (N_3560,N_2726,N_2909);
xnor U3561 (N_3561,N_2698,N_2254);
and U3562 (N_3562,N_2884,N_2616);
nor U3563 (N_3563,N_2289,N_2593);
and U3564 (N_3564,N_2281,N_2459);
xor U3565 (N_3565,N_2958,N_2458);
or U3566 (N_3566,N_2457,N_2711);
and U3567 (N_3567,N_2888,N_2643);
xnor U3568 (N_3568,N_2948,N_2567);
nor U3569 (N_3569,N_2349,N_2649);
or U3570 (N_3570,N_2787,N_2593);
or U3571 (N_3571,N_2757,N_2498);
nand U3572 (N_3572,N_2710,N_2707);
nand U3573 (N_3573,N_2884,N_2997);
xor U3574 (N_3574,N_2915,N_2739);
or U3575 (N_3575,N_2986,N_2854);
nand U3576 (N_3576,N_2967,N_2801);
nand U3577 (N_3577,N_2474,N_2399);
or U3578 (N_3578,N_2899,N_2756);
nor U3579 (N_3579,N_2281,N_2798);
nand U3580 (N_3580,N_2534,N_2951);
nor U3581 (N_3581,N_2592,N_2545);
and U3582 (N_3582,N_2424,N_2616);
or U3583 (N_3583,N_2762,N_2469);
nor U3584 (N_3584,N_2280,N_2570);
or U3585 (N_3585,N_2520,N_2684);
and U3586 (N_3586,N_2460,N_2763);
or U3587 (N_3587,N_2393,N_2437);
or U3588 (N_3588,N_2274,N_2770);
nand U3589 (N_3589,N_2397,N_2686);
or U3590 (N_3590,N_2325,N_2487);
and U3591 (N_3591,N_2732,N_2690);
and U3592 (N_3592,N_2713,N_2557);
nand U3593 (N_3593,N_2734,N_2774);
or U3594 (N_3594,N_2455,N_2412);
or U3595 (N_3595,N_2940,N_2862);
or U3596 (N_3596,N_2367,N_2604);
xor U3597 (N_3597,N_2789,N_2757);
or U3598 (N_3598,N_2469,N_2801);
or U3599 (N_3599,N_2333,N_2661);
nand U3600 (N_3600,N_2304,N_2922);
nor U3601 (N_3601,N_2259,N_2790);
and U3602 (N_3602,N_2779,N_2593);
or U3603 (N_3603,N_2356,N_2361);
or U3604 (N_3604,N_2372,N_2518);
nor U3605 (N_3605,N_2899,N_2557);
nor U3606 (N_3606,N_2521,N_2773);
and U3607 (N_3607,N_2670,N_2291);
nand U3608 (N_3608,N_2471,N_2912);
and U3609 (N_3609,N_2303,N_2947);
nand U3610 (N_3610,N_2899,N_2338);
nor U3611 (N_3611,N_2986,N_2965);
and U3612 (N_3612,N_2782,N_2381);
or U3613 (N_3613,N_2663,N_2881);
or U3614 (N_3614,N_2954,N_2569);
xnor U3615 (N_3615,N_2295,N_2597);
xnor U3616 (N_3616,N_2842,N_2302);
or U3617 (N_3617,N_2696,N_2276);
nand U3618 (N_3618,N_2557,N_2418);
xor U3619 (N_3619,N_2618,N_2574);
nand U3620 (N_3620,N_2928,N_2971);
or U3621 (N_3621,N_2979,N_2511);
or U3622 (N_3622,N_2948,N_2584);
nand U3623 (N_3623,N_2396,N_2490);
and U3624 (N_3624,N_2878,N_2455);
nand U3625 (N_3625,N_2378,N_2488);
nor U3626 (N_3626,N_2549,N_2551);
or U3627 (N_3627,N_2720,N_2714);
nor U3628 (N_3628,N_2586,N_2523);
or U3629 (N_3629,N_2260,N_2375);
nor U3630 (N_3630,N_2631,N_2929);
or U3631 (N_3631,N_2707,N_2932);
nor U3632 (N_3632,N_2432,N_2461);
xnor U3633 (N_3633,N_2409,N_2831);
or U3634 (N_3634,N_2872,N_2528);
and U3635 (N_3635,N_2846,N_2636);
or U3636 (N_3636,N_2706,N_2804);
nor U3637 (N_3637,N_2598,N_2669);
nor U3638 (N_3638,N_2969,N_2492);
nand U3639 (N_3639,N_2359,N_2706);
nand U3640 (N_3640,N_2280,N_2489);
nor U3641 (N_3641,N_2781,N_2628);
or U3642 (N_3642,N_2814,N_2848);
or U3643 (N_3643,N_2743,N_2660);
or U3644 (N_3644,N_2983,N_2522);
nor U3645 (N_3645,N_2501,N_2726);
and U3646 (N_3646,N_2476,N_2905);
nor U3647 (N_3647,N_2338,N_2907);
and U3648 (N_3648,N_2286,N_2841);
or U3649 (N_3649,N_2918,N_2977);
nand U3650 (N_3650,N_2501,N_2974);
and U3651 (N_3651,N_2575,N_2995);
nor U3652 (N_3652,N_2810,N_2857);
nand U3653 (N_3653,N_2619,N_2998);
xnor U3654 (N_3654,N_2709,N_2963);
nor U3655 (N_3655,N_2724,N_2719);
nand U3656 (N_3656,N_2479,N_2642);
xor U3657 (N_3657,N_2384,N_2709);
nand U3658 (N_3658,N_2490,N_2738);
and U3659 (N_3659,N_2886,N_2399);
and U3660 (N_3660,N_2583,N_2493);
or U3661 (N_3661,N_2379,N_2623);
nand U3662 (N_3662,N_2806,N_2250);
or U3663 (N_3663,N_2744,N_2830);
nand U3664 (N_3664,N_2608,N_2545);
nor U3665 (N_3665,N_2998,N_2629);
or U3666 (N_3666,N_2694,N_2618);
and U3667 (N_3667,N_2653,N_2307);
or U3668 (N_3668,N_2709,N_2260);
nand U3669 (N_3669,N_2818,N_2361);
nor U3670 (N_3670,N_2481,N_2609);
or U3671 (N_3671,N_2358,N_2785);
and U3672 (N_3672,N_2598,N_2648);
or U3673 (N_3673,N_2888,N_2363);
nor U3674 (N_3674,N_2708,N_2700);
nor U3675 (N_3675,N_2663,N_2650);
or U3676 (N_3676,N_2641,N_2307);
and U3677 (N_3677,N_2257,N_2820);
or U3678 (N_3678,N_2809,N_2524);
nor U3679 (N_3679,N_2952,N_2418);
or U3680 (N_3680,N_2398,N_2791);
or U3681 (N_3681,N_2593,N_2772);
or U3682 (N_3682,N_2357,N_2517);
nand U3683 (N_3683,N_2859,N_2429);
nor U3684 (N_3684,N_2585,N_2817);
xor U3685 (N_3685,N_2970,N_2884);
and U3686 (N_3686,N_2426,N_2474);
and U3687 (N_3687,N_2751,N_2274);
or U3688 (N_3688,N_2654,N_2851);
nand U3689 (N_3689,N_2549,N_2636);
nand U3690 (N_3690,N_2616,N_2430);
xor U3691 (N_3691,N_2353,N_2536);
or U3692 (N_3692,N_2571,N_2822);
nor U3693 (N_3693,N_2706,N_2609);
nand U3694 (N_3694,N_2783,N_2494);
and U3695 (N_3695,N_2516,N_2765);
xnor U3696 (N_3696,N_2947,N_2662);
or U3697 (N_3697,N_2579,N_2415);
nor U3698 (N_3698,N_2303,N_2483);
nand U3699 (N_3699,N_2535,N_2264);
and U3700 (N_3700,N_2326,N_2435);
nand U3701 (N_3701,N_2740,N_2626);
and U3702 (N_3702,N_2591,N_2808);
nor U3703 (N_3703,N_2917,N_2599);
nand U3704 (N_3704,N_2700,N_2925);
or U3705 (N_3705,N_2328,N_2304);
or U3706 (N_3706,N_2752,N_2498);
nor U3707 (N_3707,N_2918,N_2683);
nor U3708 (N_3708,N_2528,N_2619);
or U3709 (N_3709,N_2774,N_2485);
nand U3710 (N_3710,N_2332,N_2997);
nor U3711 (N_3711,N_2797,N_2635);
xnor U3712 (N_3712,N_2861,N_2781);
xor U3713 (N_3713,N_2431,N_2272);
nor U3714 (N_3714,N_2728,N_2919);
nor U3715 (N_3715,N_2727,N_2849);
or U3716 (N_3716,N_2878,N_2726);
xnor U3717 (N_3717,N_2319,N_2587);
or U3718 (N_3718,N_2605,N_2531);
nor U3719 (N_3719,N_2468,N_2890);
nor U3720 (N_3720,N_2446,N_2503);
nor U3721 (N_3721,N_2690,N_2705);
nor U3722 (N_3722,N_2426,N_2616);
or U3723 (N_3723,N_2863,N_2643);
and U3724 (N_3724,N_2299,N_2487);
nand U3725 (N_3725,N_2291,N_2920);
or U3726 (N_3726,N_2471,N_2653);
or U3727 (N_3727,N_2984,N_2676);
xor U3728 (N_3728,N_2528,N_2843);
or U3729 (N_3729,N_2763,N_2757);
or U3730 (N_3730,N_2509,N_2583);
and U3731 (N_3731,N_2560,N_2739);
nand U3732 (N_3732,N_2686,N_2668);
nor U3733 (N_3733,N_2597,N_2928);
nor U3734 (N_3734,N_2899,N_2453);
nand U3735 (N_3735,N_2978,N_2958);
nand U3736 (N_3736,N_2781,N_2347);
and U3737 (N_3737,N_2734,N_2648);
and U3738 (N_3738,N_2255,N_2875);
xor U3739 (N_3739,N_2373,N_2669);
nand U3740 (N_3740,N_2621,N_2475);
nor U3741 (N_3741,N_2983,N_2674);
or U3742 (N_3742,N_2575,N_2643);
nand U3743 (N_3743,N_2999,N_2363);
nand U3744 (N_3744,N_2899,N_2824);
nand U3745 (N_3745,N_2469,N_2811);
nor U3746 (N_3746,N_2854,N_2308);
nor U3747 (N_3747,N_2991,N_2318);
nor U3748 (N_3748,N_2796,N_2310);
nand U3749 (N_3749,N_2349,N_2551);
xor U3750 (N_3750,N_3376,N_3747);
or U3751 (N_3751,N_3555,N_3606);
or U3752 (N_3752,N_3120,N_3419);
nor U3753 (N_3753,N_3647,N_3038);
and U3754 (N_3754,N_3674,N_3610);
xor U3755 (N_3755,N_3371,N_3638);
or U3756 (N_3756,N_3730,N_3514);
nor U3757 (N_3757,N_3204,N_3065);
xnor U3758 (N_3758,N_3517,N_3289);
nor U3759 (N_3759,N_3279,N_3278);
nand U3760 (N_3760,N_3636,N_3567);
or U3761 (N_3761,N_3700,N_3098);
nor U3762 (N_3762,N_3563,N_3598);
and U3763 (N_3763,N_3218,N_3242);
nor U3764 (N_3764,N_3551,N_3334);
nor U3765 (N_3765,N_3400,N_3125);
and U3766 (N_3766,N_3281,N_3126);
or U3767 (N_3767,N_3169,N_3485);
and U3768 (N_3768,N_3620,N_3663);
or U3769 (N_3769,N_3630,N_3446);
and U3770 (N_3770,N_3471,N_3192);
xor U3771 (N_3771,N_3560,N_3541);
xnor U3772 (N_3772,N_3359,N_3687);
xor U3773 (N_3773,N_3602,N_3091);
nand U3774 (N_3774,N_3263,N_3338);
and U3775 (N_3775,N_3679,N_3503);
and U3776 (N_3776,N_3507,N_3618);
nor U3777 (N_3777,N_3059,N_3423);
nand U3778 (N_3778,N_3484,N_3629);
and U3779 (N_3779,N_3321,N_3354);
or U3780 (N_3780,N_3073,N_3720);
nor U3781 (N_3781,N_3414,N_3088);
nand U3782 (N_3782,N_3383,N_3302);
nand U3783 (N_3783,N_3511,N_3239);
xnor U3784 (N_3784,N_3078,N_3593);
nand U3785 (N_3785,N_3264,N_3481);
nor U3786 (N_3786,N_3592,N_3559);
nand U3787 (N_3787,N_3340,N_3019);
and U3788 (N_3788,N_3693,N_3637);
nor U3789 (N_3789,N_3584,N_3083);
or U3790 (N_3790,N_3196,N_3733);
nand U3791 (N_3791,N_3314,N_3228);
or U3792 (N_3792,N_3544,N_3549);
and U3793 (N_3793,N_3272,N_3205);
or U3794 (N_3794,N_3474,N_3617);
nand U3795 (N_3795,N_3112,N_3713);
nor U3796 (N_3796,N_3303,N_3722);
nand U3797 (N_3797,N_3554,N_3472);
or U3798 (N_3798,N_3666,N_3685);
nand U3799 (N_3799,N_3327,N_3389);
nor U3800 (N_3800,N_3487,N_3600);
nand U3801 (N_3801,N_3171,N_3684);
and U3802 (N_3802,N_3235,N_3313);
or U3803 (N_3803,N_3717,N_3105);
and U3804 (N_3804,N_3022,N_3273);
and U3805 (N_3805,N_3699,N_3057);
nand U3806 (N_3806,N_3249,N_3193);
and U3807 (N_3807,N_3129,N_3548);
and U3808 (N_3808,N_3203,N_3615);
nand U3809 (N_3809,N_3569,N_3649);
and U3810 (N_3810,N_3587,N_3737);
nand U3811 (N_3811,N_3144,N_3360);
nor U3812 (N_3812,N_3374,N_3741);
nor U3813 (N_3813,N_3124,N_3486);
or U3814 (N_3814,N_3337,N_3308);
nor U3815 (N_3815,N_3363,N_3052);
nand U3816 (N_3816,N_3451,N_3246);
or U3817 (N_3817,N_3325,N_3734);
xnor U3818 (N_3818,N_3590,N_3678);
nor U3819 (N_3819,N_3634,N_3266);
and U3820 (N_3820,N_3149,N_3189);
or U3821 (N_3821,N_3257,N_3058);
or U3822 (N_3822,N_3574,N_3633);
and U3823 (N_3823,N_3342,N_3448);
nor U3824 (N_3824,N_3632,N_3403);
nand U3825 (N_3825,N_3388,N_3292);
or U3826 (N_3826,N_3682,N_3491);
or U3827 (N_3827,N_3015,N_3147);
nand U3828 (N_3828,N_3355,N_3441);
xnor U3829 (N_3829,N_3702,N_3568);
or U3830 (N_3830,N_3522,N_3081);
nor U3831 (N_3831,N_3168,N_3456);
nor U3832 (N_3832,N_3709,N_3255);
nor U3833 (N_3833,N_3130,N_3050);
and U3834 (N_3834,N_3454,N_3447);
or U3835 (N_3835,N_3061,N_3316);
xnor U3836 (N_3836,N_3046,N_3558);
and U3837 (N_3837,N_3082,N_3163);
or U3838 (N_3838,N_3552,N_3557);
xor U3839 (N_3839,N_3449,N_3418);
nand U3840 (N_3840,N_3406,N_3179);
nand U3841 (N_3841,N_3166,N_3183);
and U3842 (N_3842,N_3056,N_3036);
nor U3843 (N_3843,N_3000,N_3089);
nand U3844 (N_3844,N_3521,N_3213);
or U3845 (N_3845,N_3294,N_3387);
nor U3846 (N_3846,N_3542,N_3227);
nor U3847 (N_3847,N_3018,N_3562);
xnor U3848 (N_3848,N_3433,N_3500);
nand U3849 (N_3849,N_3366,N_3087);
and U3850 (N_3850,N_3373,N_3062);
or U3851 (N_3851,N_3698,N_3466);
nand U3852 (N_3852,N_3137,N_3245);
nor U3853 (N_3853,N_3177,N_3288);
and U3854 (N_3854,N_3651,N_3247);
xnor U3855 (N_3855,N_3121,N_3128);
and U3856 (N_3856,N_3119,N_3431);
xnor U3857 (N_3857,N_3681,N_3346);
and U3858 (N_3858,N_3706,N_3315);
xor U3859 (N_3859,N_3131,N_3026);
or U3860 (N_3860,N_3650,N_3599);
or U3861 (N_3861,N_3002,N_3368);
and U3862 (N_3862,N_3386,N_3348);
nand U3863 (N_3863,N_3318,N_3404);
or U3864 (N_3864,N_3677,N_3014);
or U3865 (N_3865,N_3537,N_3113);
or U3866 (N_3866,N_3580,N_3181);
nor U3867 (N_3867,N_3626,N_3017);
nand U3868 (N_3868,N_3208,N_3728);
xnor U3869 (N_3869,N_3006,N_3194);
or U3870 (N_3870,N_3233,N_3207);
nand U3871 (N_3871,N_3270,N_3241);
nor U3872 (N_3872,N_3035,N_3442);
and U3873 (N_3873,N_3528,N_3547);
and U3874 (N_3874,N_3106,N_3165);
and U3875 (N_3875,N_3583,N_3076);
nor U3876 (N_3876,N_3627,N_3379);
nand U3877 (N_3877,N_3727,N_3077);
and U3878 (N_3878,N_3069,N_3164);
nor U3879 (N_3879,N_3284,N_3275);
nor U3880 (N_3880,N_3529,N_3200);
or U3881 (N_3881,N_3322,N_3480);
nand U3882 (N_3882,N_3276,N_3084);
nand U3883 (N_3883,N_3524,N_3619);
or U3884 (N_3884,N_3539,N_3495);
nor U3885 (N_3885,N_3254,N_3465);
or U3886 (N_3886,N_3170,N_3156);
nor U3887 (N_3887,N_3132,N_3066);
or U3888 (N_3888,N_3140,N_3101);
or U3889 (N_3889,N_3286,N_3417);
nor U3890 (N_3890,N_3477,N_3624);
or U3891 (N_3891,N_3402,N_3519);
and U3892 (N_3892,N_3182,N_3075);
or U3893 (N_3893,N_3304,N_3439);
or U3894 (N_3894,N_3043,N_3185);
and U3895 (N_3895,N_3657,N_3351);
nor U3896 (N_3896,N_3582,N_3155);
nor U3897 (N_3897,N_3108,N_3097);
and U3898 (N_3898,N_3297,N_3306);
nor U3899 (N_3899,N_3209,N_3642);
nand U3900 (N_3900,N_3060,N_3455);
or U3901 (N_3901,N_3492,N_3463);
and U3902 (N_3902,N_3109,N_3040);
nand U3903 (N_3903,N_3478,N_3708);
xnor U3904 (N_3904,N_3296,N_3738);
or U3905 (N_3905,N_3329,N_3178);
nor U3906 (N_3906,N_3437,N_3186);
and U3907 (N_3907,N_3392,N_3691);
or U3908 (N_3908,N_3021,N_3326);
and U3909 (N_3909,N_3613,N_3482);
xor U3910 (N_3910,N_3070,N_3152);
nand U3911 (N_3911,N_3307,N_3319);
or U3912 (N_3912,N_3746,N_3664);
or U3913 (N_3913,N_3413,N_3496);
nor U3914 (N_3914,N_3210,N_3725);
and U3915 (N_3915,N_3148,N_3694);
xnor U3916 (N_3916,N_3680,N_3071);
or U3917 (N_3917,N_3042,N_3635);
nand U3918 (N_3918,N_3659,N_3285);
nor U3919 (N_3919,N_3133,N_3470);
and U3920 (N_3920,N_3440,N_3425);
and U3921 (N_3921,N_3714,N_3538);
nand U3922 (N_3922,N_3715,N_3742);
nand U3923 (N_3923,N_3039,N_3645);
and U3924 (N_3924,N_3102,N_3009);
nand U3925 (N_3925,N_3622,N_3339);
and U3926 (N_3926,N_3578,N_3690);
and U3927 (N_3927,N_3460,N_3029);
or U3928 (N_3928,N_3639,N_3653);
nand U3929 (N_3929,N_3187,N_3377);
nor U3930 (N_3930,N_3670,N_3258);
or U3931 (N_3931,N_3175,N_3094);
nor U3932 (N_3932,N_3628,N_3526);
nor U3933 (N_3933,N_3453,N_3291);
nor U3934 (N_3934,N_3719,N_3689);
and U3935 (N_3935,N_3525,N_3216);
nand U3936 (N_3936,N_3369,N_3411);
or U3937 (N_3937,N_3350,N_3357);
nor U3938 (N_3938,N_3141,N_3260);
or U3939 (N_3939,N_3609,N_3004);
and U3940 (N_3940,N_3310,N_3001);
and U3941 (N_3941,N_3723,N_3508);
and U3942 (N_3942,N_3498,N_3430);
and U3943 (N_3943,N_3668,N_3143);
nor U3944 (N_3944,N_3608,N_3745);
and U3945 (N_3945,N_3122,N_3489);
nand U3946 (N_3946,N_3041,N_3420);
nor U3947 (N_3947,N_3652,N_3435);
nor U3948 (N_3948,N_3362,N_3324);
nor U3949 (N_3949,N_3581,N_3409);
xnor U3950 (N_3950,N_3244,N_3748);
nor U3951 (N_3951,N_3660,N_3665);
or U3952 (N_3952,N_3044,N_3654);
or U3953 (N_3953,N_3261,N_3585);
and U3954 (N_3954,N_3153,N_3396);
and U3955 (N_3955,N_3243,N_3100);
or U3956 (N_3956,N_3221,N_3023);
nor U3957 (N_3957,N_3703,N_3516);
and U3958 (N_3958,N_3546,N_3607);
and U3959 (N_3959,N_3184,N_3412);
or U3960 (N_3960,N_3215,N_3399);
or U3961 (N_3961,N_3127,N_3398);
xor U3962 (N_3962,N_3556,N_3509);
nand U3963 (N_3963,N_3696,N_3384);
or U3964 (N_3964,N_3422,N_3658);
nor U3965 (N_3965,N_3385,N_3621);
and U3966 (N_3966,N_3110,N_3683);
nor U3967 (N_3967,N_3375,N_3565);
or U3968 (N_3968,N_3332,N_3145);
nand U3969 (N_3969,N_3601,N_3028);
nor U3970 (N_3970,N_3219,N_3483);
and U3971 (N_3971,N_3237,N_3214);
and U3972 (N_3972,N_3176,N_3111);
nor U3973 (N_3973,N_3103,N_3151);
and U3974 (N_3974,N_3661,N_3701);
nor U3975 (N_3975,N_3107,N_3012);
nand U3976 (N_3976,N_3229,N_3739);
nor U3977 (N_3977,N_3005,N_3048);
or U3978 (N_3978,N_3157,N_3232);
nor U3979 (N_3979,N_3162,N_3595);
nand U3980 (N_3980,N_3697,N_3224);
or U3981 (N_3981,N_3139,N_3320);
nand U3982 (N_3982,N_3330,N_3055);
nor U3983 (N_3983,N_3072,N_3518);
nor U3984 (N_3984,N_3729,N_3504);
or U3985 (N_3985,N_3053,N_3494);
nand U3986 (N_3986,N_3008,N_3735);
xnor U3987 (N_3987,N_3298,N_3416);
and U3988 (N_3988,N_3054,N_3301);
nand U3989 (N_3989,N_3150,N_3501);
nor U3990 (N_3990,N_3190,N_3450);
nor U3991 (N_3991,N_3438,N_3669);
nand U3992 (N_3992,N_3506,N_3676);
xnor U3993 (N_3993,N_3591,N_3049);
and U3994 (N_3994,N_3003,N_3217);
and U3995 (N_3995,N_3570,N_3499);
xor U3996 (N_3996,N_3372,N_3114);
or U3997 (N_3997,N_3238,N_3705);
xor U3998 (N_3998,N_3533,N_3535);
nor U3999 (N_3999,N_3475,N_3010);
or U4000 (N_4000,N_3045,N_3047);
or U4001 (N_4001,N_3530,N_3154);
xor U4002 (N_4002,N_3561,N_3586);
xnor U4003 (N_4003,N_3458,N_3199);
nand U4004 (N_4004,N_3295,N_3180);
or U4005 (N_4005,N_3007,N_3274);
nand U4006 (N_4006,N_3349,N_3724);
nand U4007 (N_4007,N_3085,N_3718);
nor U4008 (N_4008,N_3434,N_3031);
nand U4009 (N_4009,N_3024,N_3749);
xor U4010 (N_4010,N_3536,N_3074);
xor U4011 (N_4011,N_3367,N_3160);
xor U4012 (N_4012,N_3250,N_3716);
or U4013 (N_4013,N_3589,N_3299);
nand U4014 (N_4014,N_3352,N_3051);
and U4015 (N_4015,N_3142,N_3079);
nor U4016 (N_4016,N_3365,N_3201);
or U4017 (N_4017,N_3280,N_3033);
nor U4018 (N_4018,N_3515,N_3265);
nand U4019 (N_4019,N_3159,N_3577);
or U4020 (N_4020,N_3711,N_3493);
nand U4021 (N_4021,N_3356,N_3603);
nand U4022 (N_4022,N_3063,N_3612);
or U4023 (N_4023,N_3573,N_3656);
nor U4024 (N_4024,N_3335,N_3673);
nand U4025 (N_4025,N_3464,N_3197);
nand U4026 (N_4026,N_3672,N_3667);
nor U4027 (N_4027,N_3259,N_3364);
nor U4028 (N_4028,N_3345,N_3220);
xnor U4029 (N_4029,N_3283,N_3428);
and U4030 (N_4030,N_3631,N_3116);
and U4031 (N_4031,N_3712,N_3740);
and U4032 (N_4032,N_3347,N_3476);
xor U4033 (N_4033,N_3462,N_3025);
and U4034 (N_4034,N_3370,N_3115);
xor U4035 (N_4035,N_3744,N_3277);
nand U4036 (N_4036,N_3134,N_3623);
xnor U4037 (N_4037,N_3067,N_3421);
nor U4038 (N_4038,N_3344,N_3675);
and U4039 (N_4039,N_3614,N_3096);
nand U4040 (N_4040,N_3037,N_3692);
nor U4041 (N_4041,N_3721,N_3671);
nor U4042 (N_4042,N_3564,N_3034);
or U4043 (N_4043,N_3251,N_3161);
and U4044 (N_4044,N_3020,N_3625);
nor U4045 (N_4045,N_3211,N_3510);
xnor U4046 (N_4046,N_3271,N_3011);
xnor U4047 (N_4047,N_3473,N_3118);
nand U4048 (N_4048,N_3688,N_3443);
nand U4049 (N_4049,N_3234,N_3467);
and U4050 (N_4050,N_3575,N_3424);
nor U4051 (N_4051,N_3571,N_3490);
nor U4052 (N_4052,N_3191,N_3445);
nor U4053 (N_4053,N_3545,N_3604);
xnor U4054 (N_4054,N_3093,N_3566);
and U4055 (N_4055,N_3240,N_3256);
and U4056 (N_4056,N_3269,N_3452);
xnor U4057 (N_4057,N_3479,N_3174);
nand U4058 (N_4058,N_3328,N_3410);
or U4059 (N_4059,N_3236,N_3596);
and U4060 (N_4060,N_3016,N_3092);
or U4061 (N_4061,N_3534,N_3226);
and U4062 (N_4062,N_3262,N_3086);
and U4063 (N_4063,N_3282,N_3378);
xor U4064 (N_4064,N_3188,N_3731);
nor U4065 (N_4065,N_3695,N_3172);
nand U4066 (N_4066,N_3550,N_3146);
nand U4067 (N_4067,N_3401,N_3576);
nor U4068 (N_4068,N_3605,N_3527);
or U4069 (N_4069,N_3531,N_3341);
nor U4070 (N_4070,N_3646,N_3643);
nand U4071 (N_4071,N_3225,N_3312);
nor U4072 (N_4072,N_3206,N_3644);
nand U4073 (N_4073,N_3095,N_3427);
and U4074 (N_4074,N_3597,N_3594);
nand U4075 (N_4075,N_3173,N_3394);
xnor U4076 (N_4076,N_3253,N_3391);
or U4077 (N_4077,N_3686,N_3502);
and U4078 (N_4078,N_3468,N_3198);
nand U4079 (N_4079,N_3287,N_3030);
nor U4080 (N_4080,N_3268,N_3353);
or U4081 (N_4081,N_3395,N_3138);
nand U4082 (N_4082,N_3432,N_3202);
and U4083 (N_4083,N_3361,N_3611);
and U4084 (N_4084,N_3343,N_3382);
nand U4085 (N_4085,N_3223,N_3013);
nor U4086 (N_4086,N_3123,N_3640);
xor U4087 (N_4087,N_3405,N_3252);
nor U4088 (N_4088,N_3704,N_3540);
xnor U4089 (N_4089,N_3064,N_3743);
or U4090 (N_4090,N_3497,N_3381);
and U4091 (N_4091,N_3358,N_3553);
or U4092 (N_4092,N_3212,N_3532);
xor U4093 (N_4093,N_3457,N_3512);
or U4094 (N_4094,N_3662,N_3641);
xor U4095 (N_4095,N_3393,N_3230);
nor U4096 (N_4096,N_3415,N_3158);
or U4097 (N_4097,N_3380,N_3736);
and U4098 (N_4098,N_3397,N_3309);
and U4099 (N_4099,N_3616,N_3135);
nor U4100 (N_4100,N_3588,N_3104);
nand U4101 (N_4101,N_3331,N_3436);
or U4102 (N_4102,N_3513,N_3267);
nand U4103 (N_4103,N_3222,N_3080);
or U4104 (N_4104,N_3290,N_3543);
or U4105 (N_4105,N_3461,N_3136);
and U4106 (N_4106,N_3710,N_3293);
nand U4107 (N_4107,N_3333,N_3469);
xnor U4108 (N_4108,N_3648,N_3429);
and U4109 (N_4109,N_3707,N_3090);
or U4110 (N_4110,N_3336,N_3407);
nor U4111 (N_4111,N_3579,N_3231);
or U4112 (N_4112,N_3572,N_3655);
nand U4113 (N_4113,N_3311,N_3426);
nand U4114 (N_4114,N_3117,N_3167);
nand U4115 (N_4115,N_3408,N_3726);
nor U4116 (N_4116,N_3099,N_3520);
and U4117 (N_4117,N_3505,N_3317);
and U4118 (N_4118,N_3248,N_3032);
nor U4119 (N_4119,N_3732,N_3068);
nor U4120 (N_4120,N_3300,N_3523);
nand U4121 (N_4121,N_3195,N_3390);
nand U4122 (N_4122,N_3027,N_3305);
xnor U4123 (N_4123,N_3323,N_3444);
nand U4124 (N_4124,N_3459,N_3488);
and U4125 (N_4125,N_3733,N_3614);
or U4126 (N_4126,N_3379,N_3116);
and U4127 (N_4127,N_3308,N_3165);
nand U4128 (N_4128,N_3259,N_3012);
and U4129 (N_4129,N_3062,N_3430);
nor U4130 (N_4130,N_3576,N_3357);
nand U4131 (N_4131,N_3701,N_3180);
nor U4132 (N_4132,N_3364,N_3727);
and U4133 (N_4133,N_3493,N_3452);
nand U4134 (N_4134,N_3180,N_3606);
nand U4135 (N_4135,N_3296,N_3111);
or U4136 (N_4136,N_3024,N_3655);
nand U4137 (N_4137,N_3150,N_3042);
nand U4138 (N_4138,N_3166,N_3632);
and U4139 (N_4139,N_3670,N_3740);
nand U4140 (N_4140,N_3045,N_3357);
nand U4141 (N_4141,N_3308,N_3526);
nand U4142 (N_4142,N_3736,N_3451);
nand U4143 (N_4143,N_3661,N_3186);
nand U4144 (N_4144,N_3642,N_3262);
nor U4145 (N_4145,N_3338,N_3530);
nand U4146 (N_4146,N_3191,N_3511);
nor U4147 (N_4147,N_3704,N_3198);
and U4148 (N_4148,N_3147,N_3182);
and U4149 (N_4149,N_3509,N_3266);
or U4150 (N_4150,N_3376,N_3192);
and U4151 (N_4151,N_3385,N_3348);
nor U4152 (N_4152,N_3234,N_3715);
nor U4153 (N_4153,N_3568,N_3225);
and U4154 (N_4154,N_3281,N_3604);
nand U4155 (N_4155,N_3625,N_3029);
and U4156 (N_4156,N_3651,N_3337);
nand U4157 (N_4157,N_3677,N_3659);
nor U4158 (N_4158,N_3521,N_3304);
and U4159 (N_4159,N_3245,N_3028);
nor U4160 (N_4160,N_3562,N_3052);
nor U4161 (N_4161,N_3584,N_3590);
and U4162 (N_4162,N_3522,N_3520);
or U4163 (N_4163,N_3417,N_3249);
nor U4164 (N_4164,N_3278,N_3488);
nor U4165 (N_4165,N_3186,N_3110);
nand U4166 (N_4166,N_3054,N_3036);
and U4167 (N_4167,N_3296,N_3645);
or U4168 (N_4168,N_3011,N_3553);
or U4169 (N_4169,N_3655,N_3436);
or U4170 (N_4170,N_3073,N_3341);
xor U4171 (N_4171,N_3096,N_3652);
or U4172 (N_4172,N_3066,N_3503);
and U4173 (N_4173,N_3013,N_3039);
nand U4174 (N_4174,N_3415,N_3632);
nand U4175 (N_4175,N_3594,N_3526);
nor U4176 (N_4176,N_3479,N_3716);
and U4177 (N_4177,N_3102,N_3050);
nor U4178 (N_4178,N_3436,N_3606);
or U4179 (N_4179,N_3718,N_3560);
and U4180 (N_4180,N_3264,N_3451);
nand U4181 (N_4181,N_3371,N_3461);
nand U4182 (N_4182,N_3078,N_3175);
nor U4183 (N_4183,N_3250,N_3592);
or U4184 (N_4184,N_3448,N_3220);
and U4185 (N_4185,N_3056,N_3412);
nand U4186 (N_4186,N_3191,N_3680);
nor U4187 (N_4187,N_3307,N_3383);
nor U4188 (N_4188,N_3027,N_3673);
or U4189 (N_4189,N_3083,N_3131);
or U4190 (N_4190,N_3577,N_3300);
or U4191 (N_4191,N_3585,N_3560);
nand U4192 (N_4192,N_3322,N_3506);
nand U4193 (N_4193,N_3358,N_3149);
or U4194 (N_4194,N_3089,N_3691);
nand U4195 (N_4195,N_3001,N_3386);
nand U4196 (N_4196,N_3275,N_3094);
nor U4197 (N_4197,N_3698,N_3057);
nand U4198 (N_4198,N_3543,N_3195);
or U4199 (N_4199,N_3270,N_3394);
and U4200 (N_4200,N_3597,N_3286);
nand U4201 (N_4201,N_3103,N_3313);
xor U4202 (N_4202,N_3363,N_3024);
and U4203 (N_4203,N_3002,N_3478);
or U4204 (N_4204,N_3022,N_3114);
or U4205 (N_4205,N_3377,N_3531);
or U4206 (N_4206,N_3416,N_3639);
or U4207 (N_4207,N_3570,N_3089);
and U4208 (N_4208,N_3670,N_3519);
or U4209 (N_4209,N_3252,N_3342);
nor U4210 (N_4210,N_3045,N_3009);
nand U4211 (N_4211,N_3213,N_3060);
nand U4212 (N_4212,N_3510,N_3707);
or U4213 (N_4213,N_3560,N_3378);
nand U4214 (N_4214,N_3349,N_3269);
or U4215 (N_4215,N_3731,N_3613);
and U4216 (N_4216,N_3430,N_3033);
nand U4217 (N_4217,N_3302,N_3640);
and U4218 (N_4218,N_3142,N_3566);
or U4219 (N_4219,N_3736,N_3252);
nor U4220 (N_4220,N_3595,N_3108);
nor U4221 (N_4221,N_3080,N_3522);
nand U4222 (N_4222,N_3559,N_3297);
nand U4223 (N_4223,N_3561,N_3713);
and U4224 (N_4224,N_3175,N_3532);
nor U4225 (N_4225,N_3703,N_3314);
nor U4226 (N_4226,N_3039,N_3087);
nand U4227 (N_4227,N_3112,N_3014);
and U4228 (N_4228,N_3423,N_3712);
nand U4229 (N_4229,N_3007,N_3397);
and U4230 (N_4230,N_3056,N_3335);
xor U4231 (N_4231,N_3431,N_3273);
nor U4232 (N_4232,N_3445,N_3435);
or U4233 (N_4233,N_3734,N_3327);
xnor U4234 (N_4234,N_3191,N_3371);
and U4235 (N_4235,N_3356,N_3435);
nand U4236 (N_4236,N_3116,N_3716);
nor U4237 (N_4237,N_3615,N_3074);
nand U4238 (N_4238,N_3150,N_3428);
nor U4239 (N_4239,N_3124,N_3319);
and U4240 (N_4240,N_3366,N_3290);
or U4241 (N_4241,N_3344,N_3671);
xnor U4242 (N_4242,N_3377,N_3668);
or U4243 (N_4243,N_3632,N_3158);
nor U4244 (N_4244,N_3515,N_3735);
or U4245 (N_4245,N_3419,N_3458);
and U4246 (N_4246,N_3026,N_3619);
nand U4247 (N_4247,N_3088,N_3412);
nand U4248 (N_4248,N_3489,N_3676);
nand U4249 (N_4249,N_3030,N_3600);
nor U4250 (N_4250,N_3230,N_3187);
nand U4251 (N_4251,N_3516,N_3397);
nor U4252 (N_4252,N_3566,N_3451);
and U4253 (N_4253,N_3186,N_3630);
nand U4254 (N_4254,N_3577,N_3314);
and U4255 (N_4255,N_3422,N_3586);
nand U4256 (N_4256,N_3491,N_3618);
and U4257 (N_4257,N_3634,N_3087);
nor U4258 (N_4258,N_3612,N_3628);
nand U4259 (N_4259,N_3298,N_3711);
and U4260 (N_4260,N_3237,N_3568);
nand U4261 (N_4261,N_3545,N_3264);
nor U4262 (N_4262,N_3311,N_3304);
and U4263 (N_4263,N_3693,N_3579);
and U4264 (N_4264,N_3037,N_3181);
and U4265 (N_4265,N_3025,N_3004);
nor U4266 (N_4266,N_3076,N_3313);
nor U4267 (N_4267,N_3715,N_3388);
and U4268 (N_4268,N_3551,N_3584);
nand U4269 (N_4269,N_3579,N_3478);
or U4270 (N_4270,N_3342,N_3676);
and U4271 (N_4271,N_3329,N_3306);
or U4272 (N_4272,N_3021,N_3647);
or U4273 (N_4273,N_3171,N_3231);
nand U4274 (N_4274,N_3012,N_3330);
or U4275 (N_4275,N_3391,N_3180);
xnor U4276 (N_4276,N_3655,N_3418);
nand U4277 (N_4277,N_3151,N_3048);
and U4278 (N_4278,N_3416,N_3557);
nor U4279 (N_4279,N_3132,N_3458);
nand U4280 (N_4280,N_3506,N_3136);
or U4281 (N_4281,N_3392,N_3522);
xnor U4282 (N_4282,N_3281,N_3004);
nor U4283 (N_4283,N_3058,N_3054);
or U4284 (N_4284,N_3683,N_3737);
nor U4285 (N_4285,N_3602,N_3727);
and U4286 (N_4286,N_3525,N_3061);
and U4287 (N_4287,N_3328,N_3491);
nand U4288 (N_4288,N_3026,N_3418);
nor U4289 (N_4289,N_3225,N_3021);
and U4290 (N_4290,N_3683,N_3147);
and U4291 (N_4291,N_3643,N_3011);
or U4292 (N_4292,N_3416,N_3088);
or U4293 (N_4293,N_3702,N_3349);
nor U4294 (N_4294,N_3597,N_3262);
nor U4295 (N_4295,N_3084,N_3472);
nand U4296 (N_4296,N_3438,N_3017);
nand U4297 (N_4297,N_3427,N_3521);
or U4298 (N_4298,N_3249,N_3086);
nor U4299 (N_4299,N_3496,N_3134);
nand U4300 (N_4300,N_3102,N_3294);
nand U4301 (N_4301,N_3449,N_3196);
nor U4302 (N_4302,N_3482,N_3235);
nor U4303 (N_4303,N_3593,N_3556);
nand U4304 (N_4304,N_3135,N_3019);
or U4305 (N_4305,N_3010,N_3095);
xnor U4306 (N_4306,N_3351,N_3399);
nand U4307 (N_4307,N_3368,N_3620);
and U4308 (N_4308,N_3414,N_3260);
nor U4309 (N_4309,N_3208,N_3370);
nor U4310 (N_4310,N_3495,N_3636);
or U4311 (N_4311,N_3383,N_3252);
nor U4312 (N_4312,N_3695,N_3302);
and U4313 (N_4313,N_3620,N_3483);
or U4314 (N_4314,N_3670,N_3226);
nor U4315 (N_4315,N_3094,N_3242);
nor U4316 (N_4316,N_3424,N_3456);
and U4317 (N_4317,N_3155,N_3585);
nor U4318 (N_4318,N_3227,N_3041);
and U4319 (N_4319,N_3734,N_3699);
and U4320 (N_4320,N_3452,N_3293);
nor U4321 (N_4321,N_3180,N_3140);
and U4322 (N_4322,N_3053,N_3388);
nand U4323 (N_4323,N_3472,N_3066);
xnor U4324 (N_4324,N_3553,N_3500);
or U4325 (N_4325,N_3603,N_3396);
nor U4326 (N_4326,N_3507,N_3125);
or U4327 (N_4327,N_3311,N_3292);
or U4328 (N_4328,N_3206,N_3009);
and U4329 (N_4329,N_3601,N_3715);
nand U4330 (N_4330,N_3615,N_3712);
and U4331 (N_4331,N_3177,N_3437);
nand U4332 (N_4332,N_3191,N_3347);
or U4333 (N_4333,N_3244,N_3259);
and U4334 (N_4334,N_3364,N_3439);
and U4335 (N_4335,N_3073,N_3177);
nor U4336 (N_4336,N_3537,N_3590);
or U4337 (N_4337,N_3399,N_3490);
nor U4338 (N_4338,N_3337,N_3619);
nand U4339 (N_4339,N_3646,N_3214);
nand U4340 (N_4340,N_3564,N_3582);
xnor U4341 (N_4341,N_3494,N_3219);
nand U4342 (N_4342,N_3702,N_3274);
nand U4343 (N_4343,N_3097,N_3459);
or U4344 (N_4344,N_3682,N_3305);
nand U4345 (N_4345,N_3413,N_3125);
nor U4346 (N_4346,N_3227,N_3140);
nor U4347 (N_4347,N_3474,N_3506);
nand U4348 (N_4348,N_3361,N_3358);
and U4349 (N_4349,N_3285,N_3587);
nand U4350 (N_4350,N_3604,N_3728);
and U4351 (N_4351,N_3167,N_3544);
and U4352 (N_4352,N_3014,N_3336);
or U4353 (N_4353,N_3719,N_3328);
and U4354 (N_4354,N_3026,N_3552);
nand U4355 (N_4355,N_3009,N_3469);
nand U4356 (N_4356,N_3266,N_3619);
nor U4357 (N_4357,N_3726,N_3069);
and U4358 (N_4358,N_3400,N_3165);
nand U4359 (N_4359,N_3622,N_3102);
xor U4360 (N_4360,N_3637,N_3418);
and U4361 (N_4361,N_3310,N_3690);
nor U4362 (N_4362,N_3315,N_3346);
or U4363 (N_4363,N_3435,N_3116);
nor U4364 (N_4364,N_3235,N_3376);
or U4365 (N_4365,N_3691,N_3261);
nor U4366 (N_4366,N_3423,N_3199);
nand U4367 (N_4367,N_3071,N_3026);
nor U4368 (N_4368,N_3363,N_3155);
or U4369 (N_4369,N_3382,N_3312);
and U4370 (N_4370,N_3191,N_3094);
nand U4371 (N_4371,N_3146,N_3511);
nand U4372 (N_4372,N_3437,N_3735);
and U4373 (N_4373,N_3656,N_3690);
nand U4374 (N_4374,N_3575,N_3595);
or U4375 (N_4375,N_3065,N_3280);
and U4376 (N_4376,N_3739,N_3663);
and U4377 (N_4377,N_3723,N_3711);
nand U4378 (N_4378,N_3090,N_3744);
or U4379 (N_4379,N_3630,N_3377);
xor U4380 (N_4380,N_3700,N_3653);
and U4381 (N_4381,N_3487,N_3147);
nor U4382 (N_4382,N_3547,N_3129);
nor U4383 (N_4383,N_3427,N_3514);
or U4384 (N_4384,N_3046,N_3255);
or U4385 (N_4385,N_3657,N_3608);
or U4386 (N_4386,N_3515,N_3457);
nand U4387 (N_4387,N_3623,N_3189);
or U4388 (N_4388,N_3085,N_3736);
nor U4389 (N_4389,N_3629,N_3641);
and U4390 (N_4390,N_3604,N_3434);
xor U4391 (N_4391,N_3330,N_3089);
nand U4392 (N_4392,N_3071,N_3087);
and U4393 (N_4393,N_3043,N_3188);
or U4394 (N_4394,N_3128,N_3584);
nand U4395 (N_4395,N_3744,N_3627);
xor U4396 (N_4396,N_3571,N_3097);
or U4397 (N_4397,N_3601,N_3348);
and U4398 (N_4398,N_3100,N_3439);
and U4399 (N_4399,N_3047,N_3646);
xnor U4400 (N_4400,N_3197,N_3647);
or U4401 (N_4401,N_3171,N_3468);
and U4402 (N_4402,N_3678,N_3354);
nor U4403 (N_4403,N_3624,N_3199);
nand U4404 (N_4404,N_3162,N_3190);
or U4405 (N_4405,N_3547,N_3214);
nor U4406 (N_4406,N_3073,N_3336);
or U4407 (N_4407,N_3543,N_3384);
nor U4408 (N_4408,N_3123,N_3418);
xor U4409 (N_4409,N_3415,N_3613);
or U4410 (N_4410,N_3384,N_3203);
nand U4411 (N_4411,N_3718,N_3225);
or U4412 (N_4412,N_3238,N_3723);
nor U4413 (N_4413,N_3732,N_3148);
xnor U4414 (N_4414,N_3448,N_3381);
nor U4415 (N_4415,N_3206,N_3064);
nand U4416 (N_4416,N_3036,N_3062);
nor U4417 (N_4417,N_3237,N_3147);
and U4418 (N_4418,N_3199,N_3173);
xor U4419 (N_4419,N_3294,N_3502);
nand U4420 (N_4420,N_3736,N_3526);
nor U4421 (N_4421,N_3171,N_3211);
nor U4422 (N_4422,N_3540,N_3299);
and U4423 (N_4423,N_3375,N_3506);
nor U4424 (N_4424,N_3308,N_3410);
nor U4425 (N_4425,N_3079,N_3261);
nand U4426 (N_4426,N_3455,N_3697);
xnor U4427 (N_4427,N_3305,N_3623);
nor U4428 (N_4428,N_3731,N_3643);
and U4429 (N_4429,N_3140,N_3345);
nand U4430 (N_4430,N_3706,N_3724);
xor U4431 (N_4431,N_3533,N_3057);
and U4432 (N_4432,N_3082,N_3216);
or U4433 (N_4433,N_3417,N_3358);
xor U4434 (N_4434,N_3021,N_3380);
nand U4435 (N_4435,N_3369,N_3310);
xor U4436 (N_4436,N_3351,N_3500);
or U4437 (N_4437,N_3361,N_3460);
or U4438 (N_4438,N_3059,N_3714);
and U4439 (N_4439,N_3403,N_3029);
nand U4440 (N_4440,N_3622,N_3692);
and U4441 (N_4441,N_3301,N_3465);
nand U4442 (N_4442,N_3655,N_3317);
nor U4443 (N_4443,N_3227,N_3603);
or U4444 (N_4444,N_3054,N_3135);
or U4445 (N_4445,N_3598,N_3463);
nor U4446 (N_4446,N_3311,N_3186);
and U4447 (N_4447,N_3543,N_3222);
and U4448 (N_4448,N_3712,N_3095);
nor U4449 (N_4449,N_3044,N_3548);
or U4450 (N_4450,N_3713,N_3159);
nand U4451 (N_4451,N_3588,N_3742);
nor U4452 (N_4452,N_3556,N_3225);
nand U4453 (N_4453,N_3505,N_3417);
nor U4454 (N_4454,N_3251,N_3257);
nor U4455 (N_4455,N_3702,N_3286);
or U4456 (N_4456,N_3039,N_3660);
xor U4457 (N_4457,N_3485,N_3130);
nor U4458 (N_4458,N_3643,N_3337);
nor U4459 (N_4459,N_3638,N_3174);
or U4460 (N_4460,N_3095,N_3250);
or U4461 (N_4461,N_3657,N_3510);
nand U4462 (N_4462,N_3377,N_3473);
nand U4463 (N_4463,N_3469,N_3308);
or U4464 (N_4464,N_3051,N_3692);
nand U4465 (N_4465,N_3628,N_3384);
nor U4466 (N_4466,N_3206,N_3655);
or U4467 (N_4467,N_3034,N_3553);
nor U4468 (N_4468,N_3575,N_3413);
nor U4469 (N_4469,N_3641,N_3256);
xor U4470 (N_4470,N_3131,N_3296);
or U4471 (N_4471,N_3327,N_3516);
nor U4472 (N_4472,N_3005,N_3462);
nand U4473 (N_4473,N_3565,N_3190);
and U4474 (N_4474,N_3233,N_3397);
nor U4475 (N_4475,N_3729,N_3470);
nand U4476 (N_4476,N_3356,N_3068);
nor U4477 (N_4477,N_3061,N_3154);
nand U4478 (N_4478,N_3277,N_3407);
or U4479 (N_4479,N_3421,N_3623);
nand U4480 (N_4480,N_3539,N_3510);
and U4481 (N_4481,N_3548,N_3699);
nor U4482 (N_4482,N_3250,N_3683);
nor U4483 (N_4483,N_3471,N_3256);
nand U4484 (N_4484,N_3165,N_3275);
nor U4485 (N_4485,N_3555,N_3737);
or U4486 (N_4486,N_3615,N_3348);
and U4487 (N_4487,N_3679,N_3417);
nand U4488 (N_4488,N_3490,N_3226);
nor U4489 (N_4489,N_3459,N_3349);
nand U4490 (N_4490,N_3715,N_3286);
nor U4491 (N_4491,N_3466,N_3177);
or U4492 (N_4492,N_3184,N_3312);
and U4493 (N_4493,N_3670,N_3333);
nor U4494 (N_4494,N_3749,N_3419);
nor U4495 (N_4495,N_3557,N_3244);
and U4496 (N_4496,N_3244,N_3403);
nor U4497 (N_4497,N_3054,N_3172);
nand U4498 (N_4498,N_3695,N_3350);
xor U4499 (N_4499,N_3427,N_3718);
or U4500 (N_4500,N_3843,N_4360);
nand U4501 (N_4501,N_3924,N_3757);
nor U4502 (N_4502,N_4419,N_4468);
or U4503 (N_4503,N_4424,N_3912);
or U4504 (N_4504,N_4238,N_3778);
nand U4505 (N_4505,N_4160,N_4322);
and U4506 (N_4506,N_3902,N_3806);
nand U4507 (N_4507,N_4261,N_4191);
nor U4508 (N_4508,N_3878,N_4306);
or U4509 (N_4509,N_4162,N_3911);
nor U4510 (N_4510,N_4056,N_3852);
or U4511 (N_4511,N_3764,N_4005);
nor U4512 (N_4512,N_4091,N_4019);
xnor U4513 (N_4513,N_3846,N_4287);
nor U4514 (N_4514,N_3922,N_4230);
nor U4515 (N_4515,N_4179,N_3782);
and U4516 (N_4516,N_3957,N_4198);
nand U4517 (N_4517,N_3802,N_3947);
and U4518 (N_4518,N_4095,N_3800);
nand U4519 (N_4519,N_4460,N_4368);
or U4520 (N_4520,N_4436,N_3986);
xor U4521 (N_4521,N_3917,N_4265);
nand U4522 (N_4522,N_4213,N_4301);
xnor U4523 (N_4523,N_4262,N_4202);
nor U4524 (N_4524,N_4080,N_4188);
and U4525 (N_4525,N_4439,N_3941);
and U4526 (N_4526,N_4237,N_3990);
nand U4527 (N_4527,N_3876,N_4099);
and U4528 (N_4528,N_3855,N_3956);
and U4529 (N_4529,N_4048,N_4105);
or U4530 (N_4530,N_4331,N_4383);
nor U4531 (N_4531,N_4067,N_4232);
nor U4532 (N_4532,N_3873,N_3938);
nand U4533 (N_4533,N_4467,N_3798);
nor U4534 (N_4534,N_4189,N_4248);
nor U4535 (N_4535,N_4352,N_3927);
nor U4536 (N_4536,N_4243,N_3996);
and U4537 (N_4537,N_4380,N_4081);
and U4538 (N_4538,N_4258,N_3942);
nand U4539 (N_4539,N_3867,N_4327);
nor U4540 (N_4540,N_4039,N_4022);
and U4541 (N_4541,N_4055,N_4144);
and U4542 (N_4542,N_4425,N_3831);
nor U4543 (N_4543,N_4354,N_4351);
or U4544 (N_4544,N_4061,N_3905);
nor U4545 (N_4545,N_3835,N_3788);
nor U4546 (N_4546,N_4033,N_4498);
or U4547 (N_4547,N_4486,N_4494);
nor U4548 (N_4548,N_3756,N_4480);
nand U4549 (N_4549,N_3860,N_4373);
nand U4550 (N_4550,N_4381,N_4429);
nand U4551 (N_4551,N_4324,N_4187);
and U4552 (N_4552,N_4129,N_3827);
and U4553 (N_4553,N_4259,N_4200);
nand U4554 (N_4554,N_3889,N_3842);
nand U4555 (N_4555,N_4348,N_4307);
xor U4556 (N_4556,N_4323,N_4483);
nand U4557 (N_4557,N_3752,N_4330);
and U4558 (N_4558,N_4207,N_3926);
nand U4559 (N_4559,N_3780,N_3854);
nand U4560 (N_4560,N_4314,N_3863);
nand U4561 (N_4561,N_3892,N_4141);
nand U4562 (N_4562,N_4403,N_4406);
nor U4563 (N_4563,N_3933,N_4010);
nand U4564 (N_4564,N_4362,N_4251);
nand U4565 (N_4565,N_4343,N_4288);
or U4566 (N_4566,N_4041,N_4418);
nor U4567 (N_4567,N_4122,N_4153);
or U4568 (N_4568,N_4441,N_4195);
nor U4569 (N_4569,N_4266,N_4297);
xnor U4570 (N_4570,N_3883,N_4020);
or U4571 (N_4571,N_4002,N_3960);
nor U4572 (N_4572,N_3971,N_4245);
nor U4573 (N_4573,N_4206,N_4004);
nand U4574 (N_4574,N_4316,N_4131);
and U4575 (N_4575,N_3944,N_4071);
or U4576 (N_4576,N_4282,N_4278);
nand U4577 (N_4577,N_4180,N_3750);
and U4578 (N_4578,N_3862,N_3916);
or U4579 (N_4579,N_4374,N_4044);
and U4580 (N_4580,N_3840,N_4392);
nor U4581 (N_4581,N_3858,N_4239);
or U4582 (N_4582,N_3871,N_4130);
nor U4583 (N_4583,N_4084,N_4047);
or U4584 (N_4584,N_3880,N_4367);
nor U4585 (N_4585,N_3921,N_4092);
nor U4586 (N_4586,N_4066,N_4231);
nand U4587 (N_4587,N_4384,N_4434);
nor U4588 (N_4588,N_4397,N_4300);
and U4589 (N_4589,N_3787,N_4499);
xor U4590 (N_4590,N_3950,N_3784);
nor U4591 (N_4591,N_4390,N_4456);
nor U4592 (N_4592,N_4219,N_4274);
and U4593 (N_4593,N_4021,N_4221);
nand U4594 (N_4594,N_3887,N_4457);
or U4595 (N_4595,N_4059,N_4063);
nand U4596 (N_4596,N_4125,N_4378);
nor U4597 (N_4597,N_4442,N_4489);
or U4598 (N_4598,N_3789,N_4358);
nor U4599 (N_4599,N_3805,N_4340);
nor U4600 (N_4600,N_4190,N_4495);
nand U4601 (N_4601,N_4437,N_4224);
nor U4602 (N_4602,N_4026,N_4275);
or U4603 (N_4603,N_3810,N_3949);
or U4604 (N_4604,N_4032,N_4208);
nand U4605 (N_4605,N_4347,N_4484);
and U4606 (N_4606,N_3998,N_4050);
nor U4607 (N_4607,N_3868,N_4292);
nand U4608 (N_4608,N_4427,N_4074);
nor U4609 (N_4609,N_4433,N_3803);
and U4610 (N_4610,N_4075,N_3962);
or U4611 (N_4611,N_4396,N_4319);
and U4612 (N_4612,N_4291,N_3919);
xor U4613 (N_4613,N_3847,N_4242);
nor U4614 (N_4614,N_4375,N_3943);
and U4615 (N_4615,N_4379,N_4276);
xor U4616 (N_4616,N_4305,N_4270);
nand U4617 (N_4617,N_4445,N_4488);
xnor U4618 (N_4618,N_4103,N_3859);
nor U4619 (N_4619,N_4106,N_4393);
or U4620 (N_4620,N_4088,N_3899);
or U4621 (N_4621,N_4249,N_3755);
nor U4622 (N_4622,N_4009,N_4165);
or U4623 (N_4623,N_3797,N_3965);
nor U4624 (N_4624,N_4235,N_4446);
nor U4625 (N_4625,N_4459,N_4264);
nor U4626 (N_4626,N_4108,N_4449);
and U4627 (N_4627,N_4387,N_3837);
or U4628 (N_4628,N_4082,N_3995);
nand U4629 (N_4629,N_3754,N_3759);
nor U4630 (N_4630,N_4415,N_4176);
or U4631 (N_4631,N_4426,N_4487);
xnor U4632 (N_4632,N_3761,N_3991);
nor U4633 (N_4633,N_3848,N_4127);
or U4634 (N_4634,N_4205,N_4199);
or U4635 (N_4635,N_4365,N_3825);
nor U4636 (N_4636,N_3839,N_3885);
and U4637 (N_4637,N_4097,N_4283);
or U4638 (N_4638,N_4151,N_3801);
xnor U4639 (N_4639,N_4051,N_3774);
or U4640 (N_4640,N_4169,N_3970);
nand U4641 (N_4641,N_4057,N_4400);
and U4642 (N_4642,N_3771,N_4220);
and U4643 (N_4643,N_4196,N_4104);
nor U4644 (N_4644,N_4184,N_3935);
and U4645 (N_4645,N_4172,N_3909);
nand U4646 (N_4646,N_4110,N_4045);
and U4647 (N_4647,N_4014,N_4293);
and U4648 (N_4648,N_4211,N_4173);
and U4649 (N_4649,N_4234,N_4253);
nor U4650 (N_4650,N_4015,N_4453);
or U4651 (N_4651,N_4277,N_4431);
and U4652 (N_4652,N_3973,N_4000);
or U4653 (N_4653,N_4223,N_4273);
nor U4654 (N_4654,N_3898,N_4147);
or U4655 (N_4655,N_3896,N_4133);
and U4656 (N_4656,N_4268,N_3785);
nor U4657 (N_4657,N_4395,N_4318);
nand U4658 (N_4658,N_3779,N_3999);
and U4659 (N_4659,N_4236,N_4333);
or U4660 (N_4660,N_3851,N_3882);
nor U4661 (N_4661,N_4413,N_3984);
nor U4662 (N_4662,N_4119,N_4254);
or U4663 (N_4663,N_4115,N_4335);
nand U4664 (N_4664,N_4185,N_3866);
and U4665 (N_4665,N_4073,N_3946);
nor U4666 (N_4666,N_3870,N_4289);
nand U4667 (N_4667,N_3961,N_4012);
and U4668 (N_4668,N_4201,N_3963);
nor U4669 (N_4669,N_3823,N_3983);
nand U4670 (N_4670,N_3793,N_3813);
nor U4671 (N_4671,N_4295,N_4194);
and U4672 (N_4672,N_3817,N_4077);
nor U4673 (N_4673,N_3792,N_4309);
and U4674 (N_4674,N_3895,N_4336);
nor U4675 (N_4675,N_4177,N_4136);
or U4676 (N_4676,N_4040,N_4369);
nand U4677 (N_4677,N_4222,N_4053);
xor U4678 (N_4678,N_4438,N_3969);
nand U4679 (N_4679,N_4093,N_4370);
and U4680 (N_4680,N_3891,N_4428);
nor U4681 (N_4681,N_3822,N_4152);
nand U4682 (N_4682,N_4281,N_3972);
nor U4683 (N_4683,N_4170,N_4027);
nor U4684 (N_4684,N_4017,N_4443);
or U4685 (N_4685,N_3979,N_3799);
nand U4686 (N_4686,N_4256,N_3888);
and U4687 (N_4687,N_4113,N_4462);
xor U4688 (N_4688,N_4416,N_4361);
nor U4689 (N_4689,N_4430,N_4070);
nand U4690 (N_4690,N_3952,N_4475);
nand U4691 (N_4691,N_3934,N_4338);
and U4692 (N_4692,N_4035,N_4356);
nand U4693 (N_4693,N_3811,N_3829);
and U4694 (N_4694,N_3791,N_4156);
and U4695 (N_4695,N_4308,N_4226);
nand U4696 (N_4696,N_3903,N_3923);
xor U4697 (N_4697,N_4043,N_4124);
and U4698 (N_4698,N_4046,N_3959);
nor U4699 (N_4699,N_4025,N_4466);
and U4700 (N_4700,N_3932,N_3978);
or U4701 (N_4701,N_3980,N_3836);
and U4702 (N_4702,N_4294,N_3818);
nor U4703 (N_4703,N_4143,N_3948);
nand U4704 (N_4704,N_3890,N_4357);
or U4705 (N_4705,N_4377,N_3987);
nor U4706 (N_4706,N_4037,N_4345);
or U4707 (N_4707,N_3906,N_3872);
nor U4708 (N_4708,N_3945,N_3790);
nand U4709 (N_4709,N_4272,N_4317);
nand U4710 (N_4710,N_4279,N_4038);
xnor U4711 (N_4711,N_4072,N_3874);
nand U4712 (N_4712,N_3992,N_3920);
nand U4713 (N_4713,N_4315,N_4328);
nor U4714 (N_4714,N_4497,N_3830);
nand U4715 (N_4715,N_4491,N_4036);
and U4716 (N_4716,N_4342,N_4089);
xnor U4717 (N_4717,N_4477,N_3897);
nor U4718 (N_4718,N_4132,N_4376);
nand U4719 (N_4719,N_4386,N_4158);
nand U4720 (N_4720,N_4079,N_4042);
nor U4721 (N_4721,N_4112,N_4126);
or U4722 (N_4722,N_4204,N_4420);
and U4723 (N_4723,N_4006,N_4432);
nor U4724 (N_4724,N_4086,N_4321);
nor U4725 (N_4725,N_4087,N_4109);
nor U4726 (N_4726,N_4182,N_4410);
or U4727 (N_4727,N_3781,N_4094);
nor U4728 (N_4728,N_3849,N_4366);
and U4729 (N_4729,N_4472,N_4461);
nor U4730 (N_4730,N_4470,N_4178);
nand U4731 (N_4731,N_3856,N_4490);
nor U4732 (N_4732,N_4128,N_4161);
nand U4733 (N_4733,N_4142,N_4139);
nand U4734 (N_4734,N_4018,N_3915);
or U4735 (N_4735,N_3940,N_4382);
xor U4736 (N_4736,N_4155,N_4450);
nor U4737 (N_4737,N_3853,N_4479);
nor U4738 (N_4738,N_3988,N_3770);
nor U4739 (N_4739,N_4463,N_4263);
nor U4740 (N_4740,N_4031,N_4447);
and U4741 (N_4741,N_4471,N_4102);
xnor U4742 (N_4742,N_4257,N_4454);
xnor U4743 (N_4743,N_4422,N_4062);
nor U4744 (N_4744,N_4313,N_4229);
or U4745 (N_4745,N_4280,N_3964);
or U4746 (N_4746,N_4003,N_4101);
nor U4747 (N_4747,N_3884,N_3834);
nand U4748 (N_4748,N_4421,N_4118);
nor U4749 (N_4749,N_4083,N_3864);
and U4750 (N_4750,N_4150,N_3953);
and U4751 (N_4751,N_4203,N_4225);
nor U4752 (N_4752,N_4214,N_3767);
and U4753 (N_4753,N_4469,N_4341);
nor U4754 (N_4754,N_4455,N_4210);
and U4755 (N_4755,N_3861,N_4355);
and U4756 (N_4756,N_4135,N_4304);
and U4757 (N_4757,N_4078,N_4052);
nor U4758 (N_4758,N_4496,N_3908);
and U4759 (N_4759,N_4121,N_4148);
and U4760 (N_4760,N_4337,N_4209);
nand U4761 (N_4761,N_4116,N_4228);
nand U4762 (N_4762,N_4216,N_4164);
nand U4763 (N_4763,N_3763,N_3869);
and U4764 (N_4764,N_3777,N_3966);
or U4765 (N_4765,N_4286,N_4407);
nor U4766 (N_4766,N_3804,N_4123);
nand U4767 (N_4767,N_4054,N_3775);
or U4768 (N_4768,N_3844,N_4371);
nand U4769 (N_4769,N_4154,N_4117);
nand U4770 (N_4770,N_4267,N_4412);
nand U4771 (N_4771,N_4476,N_3808);
nand U4772 (N_4772,N_3751,N_4485);
nor U4773 (N_4773,N_4269,N_4167);
and U4774 (N_4774,N_4311,N_3931);
or U4775 (N_4775,N_4284,N_3958);
nand U4776 (N_4776,N_3981,N_4398);
and U4777 (N_4777,N_3955,N_4320);
nor U4778 (N_4778,N_4016,N_4492);
or U4779 (N_4779,N_4007,N_4334);
nand U4780 (N_4780,N_3914,N_4440);
or U4781 (N_4781,N_4183,N_4023);
and U4782 (N_4782,N_3796,N_4458);
or U4783 (N_4783,N_4448,N_4409);
or U4784 (N_4784,N_3881,N_4252);
or U4785 (N_4785,N_3765,N_4329);
and U4786 (N_4786,N_4138,N_4149);
and U4787 (N_4787,N_3795,N_3809);
nand U4788 (N_4788,N_3993,N_4385);
nor U4789 (N_4789,N_4478,N_4029);
nor U4790 (N_4790,N_4192,N_4008);
or U4791 (N_4791,N_4417,N_4064);
or U4792 (N_4792,N_4404,N_4058);
nand U4793 (N_4793,N_4303,N_4250);
and U4794 (N_4794,N_4473,N_4111);
or U4795 (N_4795,N_3967,N_4186);
or U4796 (N_4796,N_3812,N_3814);
xor U4797 (N_4797,N_4060,N_4326);
or U4798 (N_4798,N_4452,N_3982);
nand U4799 (N_4799,N_3893,N_3994);
xor U4800 (N_4800,N_3894,N_4096);
nor U4801 (N_4801,N_3828,N_3794);
nor U4802 (N_4802,N_4298,N_3877);
nor U4803 (N_4803,N_4451,N_4193);
or U4804 (N_4804,N_3753,N_3786);
nor U4805 (N_4805,N_4372,N_4114);
and U4806 (N_4806,N_3819,N_3939);
or U4807 (N_4807,N_4049,N_4171);
nand U4808 (N_4808,N_3768,N_4140);
or U4809 (N_4809,N_3821,N_4069);
or U4810 (N_4810,N_3766,N_4076);
xor U4811 (N_4811,N_4065,N_4068);
and U4812 (N_4812,N_4464,N_4181);
or U4813 (N_4813,N_4405,N_4359);
nor U4814 (N_4814,N_4174,N_3776);
xnor U4815 (N_4815,N_4241,N_3833);
or U4816 (N_4816,N_4145,N_3815);
or U4817 (N_4817,N_4163,N_4402);
and U4818 (N_4818,N_3783,N_4481);
nand U4819 (N_4819,N_4325,N_4271);
nor U4820 (N_4820,N_3904,N_4030);
nand U4821 (N_4821,N_4474,N_4098);
and U4822 (N_4822,N_3968,N_4246);
nor U4823 (N_4823,N_4260,N_3930);
and U4824 (N_4824,N_3773,N_3769);
nand U4825 (N_4825,N_4100,N_4310);
and U4826 (N_4826,N_4332,N_3886);
nand U4827 (N_4827,N_4107,N_4296);
nor U4828 (N_4828,N_4394,N_4364);
nand U4829 (N_4829,N_4290,N_3936);
and U4830 (N_4830,N_4389,N_4227);
nand U4831 (N_4831,N_4085,N_3850);
or U4832 (N_4832,N_3824,N_4166);
nor U4833 (N_4833,N_4244,N_3901);
xor U4834 (N_4834,N_4011,N_3976);
and U4835 (N_4835,N_4482,N_4255);
and U4836 (N_4836,N_4465,N_3875);
nand U4837 (N_4837,N_3985,N_3918);
nor U4838 (N_4838,N_3954,N_4408);
nor U4839 (N_4839,N_3845,N_3977);
nor U4840 (N_4840,N_4299,N_4120);
nor U4841 (N_4841,N_3826,N_4175);
nor U4842 (N_4842,N_3832,N_4401);
and U4843 (N_4843,N_4399,N_3838);
nand U4844 (N_4844,N_4411,N_4024);
or U4845 (N_4845,N_3762,N_4353);
or U4846 (N_4846,N_4344,N_4414);
or U4847 (N_4847,N_3816,N_4493);
and U4848 (N_4848,N_4212,N_4197);
and U4849 (N_4849,N_4339,N_3910);
or U4850 (N_4850,N_3928,N_3900);
or U4851 (N_4851,N_3951,N_3907);
and U4852 (N_4852,N_4423,N_3997);
or U4853 (N_4853,N_3879,N_4312);
nand U4854 (N_4854,N_4217,N_4350);
and U4855 (N_4855,N_3857,N_4233);
nor U4856 (N_4856,N_4346,N_3772);
and U4857 (N_4857,N_4001,N_3974);
xor U4858 (N_4858,N_4146,N_3975);
or U4859 (N_4859,N_4349,N_3989);
or U4860 (N_4860,N_4247,N_3807);
or U4861 (N_4861,N_4090,N_4240);
or U4862 (N_4862,N_4134,N_4168);
nor U4863 (N_4863,N_4157,N_3925);
or U4864 (N_4864,N_3760,N_4013);
or U4865 (N_4865,N_4444,N_4218);
xnor U4866 (N_4866,N_4285,N_3929);
nand U4867 (N_4867,N_4435,N_3820);
xnor U4868 (N_4868,N_3937,N_3913);
nor U4869 (N_4869,N_4028,N_4034);
nor U4870 (N_4870,N_4391,N_4137);
or U4871 (N_4871,N_4302,N_4215);
or U4872 (N_4872,N_4159,N_3865);
or U4873 (N_4873,N_3758,N_3841);
nand U4874 (N_4874,N_4363,N_4388);
xnor U4875 (N_4875,N_4130,N_4350);
or U4876 (N_4876,N_4345,N_4286);
and U4877 (N_4877,N_4081,N_4424);
nor U4878 (N_4878,N_4166,N_3916);
nand U4879 (N_4879,N_3938,N_4417);
and U4880 (N_4880,N_4391,N_4069);
and U4881 (N_4881,N_3963,N_4313);
nand U4882 (N_4882,N_4168,N_4051);
nor U4883 (N_4883,N_3950,N_3929);
and U4884 (N_4884,N_4079,N_3867);
xor U4885 (N_4885,N_4329,N_4056);
and U4886 (N_4886,N_3986,N_4071);
nand U4887 (N_4887,N_3787,N_4163);
and U4888 (N_4888,N_4146,N_4266);
nand U4889 (N_4889,N_3980,N_4069);
nor U4890 (N_4890,N_3850,N_4276);
nor U4891 (N_4891,N_3892,N_4054);
or U4892 (N_4892,N_4287,N_4129);
nand U4893 (N_4893,N_4296,N_3856);
nand U4894 (N_4894,N_3927,N_4409);
or U4895 (N_4895,N_4058,N_4340);
or U4896 (N_4896,N_3925,N_4434);
nor U4897 (N_4897,N_4016,N_4382);
and U4898 (N_4898,N_4184,N_3776);
nand U4899 (N_4899,N_4002,N_4197);
xnor U4900 (N_4900,N_3891,N_3886);
nand U4901 (N_4901,N_4199,N_4348);
and U4902 (N_4902,N_4064,N_4308);
nand U4903 (N_4903,N_4200,N_3755);
nor U4904 (N_4904,N_4039,N_4030);
nor U4905 (N_4905,N_4057,N_4492);
or U4906 (N_4906,N_3789,N_3795);
xnor U4907 (N_4907,N_3918,N_4123);
nor U4908 (N_4908,N_3830,N_4367);
nor U4909 (N_4909,N_3796,N_4492);
and U4910 (N_4910,N_4042,N_4240);
xor U4911 (N_4911,N_3956,N_4041);
nor U4912 (N_4912,N_3893,N_4346);
and U4913 (N_4913,N_3881,N_4139);
nor U4914 (N_4914,N_4403,N_4424);
nor U4915 (N_4915,N_3877,N_4233);
xor U4916 (N_4916,N_4127,N_4271);
nand U4917 (N_4917,N_4450,N_4018);
nor U4918 (N_4918,N_3826,N_3927);
or U4919 (N_4919,N_4047,N_4423);
and U4920 (N_4920,N_4215,N_4014);
nand U4921 (N_4921,N_4266,N_4007);
or U4922 (N_4922,N_3927,N_4125);
nand U4923 (N_4923,N_4110,N_4458);
nor U4924 (N_4924,N_3776,N_4038);
nand U4925 (N_4925,N_4481,N_4427);
and U4926 (N_4926,N_4281,N_4077);
nor U4927 (N_4927,N_3781,N_3779);
nor U4928 (N_4928,N_4463,N_4311);
and U4929 (N_4929,N_3852,N_4277);
nor U4930 (N_4930,N_4245,N_4263);
and U4931 (N_4931,N_4385,N_4003);
or U4932 (N_4932,N_4052,N_3839);
nor U4933 (N_4933,N_4244,N_3914);
and U4934 (N_4934,N_3805,N_3817);
and U4935 (N_4935,N_4094,N_3890);
nand U4936 (N_4936,N_3773,N_4196);
and U4937 (N_4937,N_4044,N_3981);
nand U4938 (N_4938,N_4406,N_4303);
or U4939 (N_4939,N_3944,N_3973);
or U4940 (N_4940,N_4486,N_3956);
and U4941 (N_4941,N_4194,N_4154);
nor U4942 (N_4942,N_3936,N_4031);
or U4943 (N_4943,N_4269,N_4014);
and U4944 (N_4944,N_3882,N_3787);
nand U4945 (N_4945,N_3968,N_4295);
xor U4946 (N_4946,N_4477,N_4093);
and U4947 (N_4947,N_4112,N_3927);
nor U4948 (N_4948,N_4187,N_4332);
nand U4949 (N_4949,N_3773,N_3786);
and U4950 (N_4950,N_4099,N_3905);
nor U4951 (N_4951,N_4454,N_4061);
nand U4952 (N_4952,N_3774,N_4180);
nor U4953 (N_4953,N_4366,N_4469);
nor U4954 (N_4954,N_4014,N_3851);
xnor U4955 (N_4955,N_3917,N_4030);
nand U4956 (N_4956,N_3831,N_4215);
nor U4957 (N_4957,N_4311,N_4428);
and U4958 (N_4958,N_4089,N_3863);
and U4959 (N_4959,N_4477,N_3814);
nor U4960 (N_4960,N_3963,N_4216);
nor U4961 (N_4961,N_3783,N_3982);
nor U4962 (N_4962,N_4385,N_4139);
nor U4963 (N_4963,N_4095,N_3813);
nand U4964 (N_4964,N_4143,N_3791);
xnor U4965 (N_4965,N_4044,N_3873);
nor U4966 (N_4966,N_3936,N_3775);
nor U4967 (N_4967,N_4012,N_3885);
or U4968 (N_4968,N_4247,N_4498);
and U4969 (N_4969,N_3756,N_4225);
or U4970 (N_4970,N_3822,N_4228);
nand U4971 (N_4971,N_3938,N_4441);
nor U4972 (N_4972,N_3850,N_4243);
nor U4973 (N_4973,N_4096,N_4037);
and U4974 (N_4974,N_4173,N_3885);
or U4975 (N_4975,N_4076,N_4072);
nor U4976 (N_4976,N_4371,N_3767);
and U4977 (N_4977,N_4327,N_4046);
or U4978 (N_4978,N_4468,N_4244);
xnor U4979 (N_4979,N_4083,N_4169);
xnor U4980 (N_4980,N_4168,N_4063);
and U4981 (N_4981,N_4108,N_3808);
nor U4982 (N_4982,N_4304,N_4166);
or U4983 (N_4983,N_4315,N_3852);
or U4984 (N_4984,N_4141,N_3925);
or U4985 (N_4985,N_4260,N_4248);
and U4986 (N_4986,N_3864,N_3809);
or U4987 (N_4987,N_4231,N_4202);
or U4988 (N_4988,N_4034,N_3959);
nand U4989 (N_4989,N_3983,N_4162);
nand U4990 (N_4990,N_4157,N_4105);
nor U4991 (N_4991,N_4265,N_3826);
nand U4992 (N_4992,N_4347,N_4317);
nand U4993 (N_4993,N_4208,N_3931);
and U4994 (N_4994,N_4094,N_4301);
xnor U4995 (N_4995,N_4120,N_4460);
or U4996 (N_4996,N_4082,N_4163);
or U4997 (N_4997,N_3809,N_3926);
xnor U4998 (N_4998,N_3752,N_3845);
nand U4999 (N_4999,N_3996,N_4078);
and U5000 (N_5000,N_3755,N_4134);
or U5001 (N_5001,N_4145,N_3765);
and U5002 (N_5002,N_3783,N_4476);
or U5003 (N_5003,N_4474,N_4209);
xor U5004 (N_5004,N_3776,N_4140);
and U5005 (N_5005,N_4453,N_4357);
and U5006 (N_5006,N_4285,N_4361);
nor U5007 (N_5007,N_4262,N_3935);
nand U5008 (N_5008,N_4102,N_3893);
or U5009 (N_5009,N_4099,N_4201);
and U5010 (N_5010,N_4039,N_3875);
and U5011 (N_5011,N_3772,N_4004);
or U5012 (N_5012,N_4427,N_4328);
or U5013 (N_5013,N_3856,N_3886);
nand U5014 (N_5014,N_4368,N_4173);
nand U5015 (N_5015,N_4457,N_4185);
xnor U5016 (N_5016,N_4157,N_4054);
nor U5017 (N_5017,N_4438,N_3820);
and U5018 (N_5018,N_4288,N_3966);
xor U5019 (N_5019,N_4013,N_4077);
nor U5020 (N_5020,N_3888,N_4305);
and U5021 (N_5021,N_4271,N_3769);
nand U5022 (N_5022,N_4136,N_3808);
or U5023 (N_5023,N_3974,N_4481);
or U5024 (N_5024,N_4024,N_4396);
xor U5025 (N_5025,N_4497,N_4280);
nand U5026 (N_5026,N_4149,N_4270);
and U5027 (N_5027,N_3952,N_4314);
and U5028 (N_5028,N_4117,N_4422);
nor U5029 (N_5029,N_4483,N_4309);
or U5030 (N_5030,N_3795,N_4185);
and U5031 (N_5031,N_4223,N_4476);
nand U5032 (N_5032,N_4336,N_4289);
or U5033 (N_5033,N_4098,N_3827);
nor U5034 (N_5034,N_4017,N_4406);
and U5035 (N_5035,N_4244,N_4405);
and U5036 (N_5036,N_4274,N_4179);
and U5037 (N_5037,N_3871,N_3969);
nand U5038 (N_5038,N_4048,N_4085);
xnor U5039 (N_5039,N_4160,N_3912);
and U5040 (N_5040,N_4054,N_3945);
nor U5041 (N_5041,N_4123,N_3856);
nand U5042 (N_5042,N_4249,N_3982);
nor U5043 (N_5043,N_3970,N_4468);
nand U5044 (N_5044,N_3976,N_4345);
or U5045 (N_5045,N_4367,N_3926);
or U5046 (N_5046,N_4175,N_4282);
and U5047 (N_5047,N_4094,N_4186);
or U5048 (N_5048,N_3810,N_3801);
nand U5049 (N_5049,N_4313,N_3838);
or U5050 (N_5050,N_4383,N_3769);
or U5051 (N_5051,N_4170,N_4262);
xnor U5052 (N_5052,N_3777,N_4255);
nand U5053 (N_5053,N_4104,N_4200);
nand U5054 (N_5054,N_3879,N_4014);
nor U5055 (N_5055,N_3750,N_4438);
or U5056 (N_5056,N_4050,N_4153);
nor U5057 (N_5057,N_4162,N_3984);
nand U5058 (N_5058,N_3861,N_4353);
or U5059 (N_5059,N_4434,N_4402);
or U5060 (N_5060,N_3994,N_4387);
nor U5061 (N_5061,N_3825,N_4225);
nor U5062 (N_5062,N_4036,N_4046);
nand U5063 (N_5063,N_3806,N_4345);
nor U5064 (N_5064,N_4431,N_3896);
or U5065 (N_5065,N_3837,N_4378);
or U5066 (N_5066,N_4290,N_4055);
or U5067 (N_5067,N_4422,N_4320);
nor U5068 (N_5068,N_3932,N_3956);
nor U5069 (N_5069,N_3999,N_3771);
nand U5070 (N_5070,N_4249,N_4167);
nand U5071 (N_5071,N_4389,N_4133);
or U5072 (N_5072,N_4374,N_4295);
or U5073 (N_5073,N_3783,N_4104);
nor U5074 (N_5074,N_3802,N_3941);
and U5075 (N_5075,N_4221,N_3840);
nor U5076 (N_5076,N_4336,N_4349);
or U5077 (N_5077,N_4238,N_3798);
and U5078 (N_5078,N_4494,N_4290);
nor U5079 (N_5079,N_3863,N_4178);
xor U5080 (N_5080,N_3949,N_4361);
or U5081 (N_5081,N_4481,N_4468);
and U5082 (N_5082,N_4224,N_3982);
and U5083 (N_5083,N_3881,N_3820);
or U5084 (N_5084,N_4085,N_3773);
and U5085 (N_5085,N_3849,N_4327);
and U5086 (N_5086,N_4419,N_3771);
or U5087 (N_5087,N_4184,N_4279);
or U5088 (N_5088,N_3850,N_3775);
and U5089 (N_5089,N_4291,N_3830);
and U5090 (N_5090,N_4092,N_4033);
or U5091 (N_5091,N_4283,N_3932);
or U5092 (N_5092,N_3817,N_3766);
and U5093 (N_5093,N_3809,N_4052);
xnor U5094 (N_5094,N_4279,N_3752);
and U5095 (N_5095,N_4214,N_4489);
nand U5096 (N_5096,N_3915,N_3886);
or U5097 (N_5097,N_3974,N_4380);
or U5098 (N_5098,N_4033,N_3862);
and U5099 (N_5099,N_4282,N_4411);
nand U5100 (N_5100,N_4282,N_3909);
and U5101 (N_5101,N_4056,N_4362);
nand U5102 (N_5102,N_3866,N_3787);
xor U5103 (N_5103,N_3953,N_3863);
nand U5104 (N_5104,N_3999,N_4427);
nor U5105 (N_5105,N_3994,N_3835);
nand U5106 (N_5106,N_4349,N_4480);
nor U5107 (N_5107,N_4387,N_4204);
nand U5108 (N_5108,N_3859,N_4040);
and U5109 (N_5109,N_4497,N_4154);
and U5110 (N_5110,N_4070,N_4322);
or U5111 (N_5111,N_4425,N_3791);
nor U5112 (N_5112,N_4498,N_4293);
nand U5113 (N_5113,N_4389,N_4328);
nand U5114 (N_5114,N_3875,N_3854);
and U5115 (N_5115,N_4155,N_4302);
or U5116 (N_5116,N_4334,N_3985);
and U5117 (N_5117,N_4251,N_4384);
or U5118 (N_5118,N_4040,N_4190);
xor U5119 (N_5119,N_4143,N_3780);
or U5120 (N_5120,N_3949,N_3750);
nor U5121 (N_5121,N_4080,N_3841);
nand U5122 (N_5122,N_3799,N_3887);
or U5123 (N_5123,N_3871,N_3930);
or U5124 (N_5124,N_3950,N_4215);
nor U5125 (N_5125,N_4004,N_4164);
or U5126 (N_5126,N_3953,N_4428);
nand U5127 (N_5127,N_3912,N_4434);
or U5128 (N_5128,N_4046,N_4208);
nand U5129 (N_5129,N_4491,N_4322);
nor U5130 (N_5130,N_4214,N_4497);
nand U5131 (N_5131,N_4125,N_4444);
xnor U5132 (N_5132,N_4473,N_4132);
or U5133 (N_5133,N_4424,N_3792);
or U5134 (N_5134,N_4149,N_3886);
nand U5135 (N_5135,N_3867,N_3919);
nand U5136 (N_5136,N_3920,N_3944);
nor U5137 (N_5137,N_4163,N_4120);
or U5138 (N_5138,N_4320,N_3961);
or U5139 (N_5139,N_4168,N_4431);
nor U5140 (N_5140,N_4064,N_3836);
and U5141 (N_5141,N_4225,N_3918);
or U5142 (N_5142,N_4277,N_4157);
nand U5143 (N_5143,N_4391,N_4239);
and U5144 (N_5144,N_4107,N_3818);
or U5145 (N_5145,N_4371,N_4103);
or U5146 (N_5146,N_4232,N_4025);
and U5147 (N_5147,N_4093,N_4017);
or U5148 (N_5148,N_3932,N_4051);
nor U5149 (N_5149,N_3988,N_4439);
nand U5150 (N_5150,N_4054,N_4425);
or U5151 (N_5151,N_4154,N_4147);
and U5152 (N_5152,N_4262,N_3881);
xor U5153 (N_5153,N_4356,N_4061);
nor U5154 (N_5154,N_3900,N_4438);
nor U5155 (N_5155,N_4338,N_3912);
nand U5156 (N_5156,N_4460,N_3801);
xor U5157 (N_5157,N_3761,N_4163);
or U5158 (N_5158,N_4204,N_4233);
or U5159 (N_5159,N_4229,N_4298);
or U5160 (N_5160,N_3879,N_4319);
nand U5161 (N_5161,N_4283,N_4116);
nor U5162 (N_5162,N_4394,N_4452);
and U5163 (N_5163,N_4494,N_3928);
xor U5164 (N_5164,N_4081,N_4401);
nor U5165 (N_5165,N_4252,N_3765);
xor U5166 (N_5166,N_4452,N_4141);
and U5167 (N_5167,N_3922,N_4485);
nand U5168 (N_5168,N_4391,N_4274);
nor U5169 (N_5169,N_3872,N_3959);
and U5170 (N_5170,N_3852,N_4117);
and U5171 (N_5171,N_3779,N_4093);
xor U5172 (N_5172,N_4426,N_4258);
or U5173 (N_5173,N_4445,N_4031);
or U5174 (N_5174,N_4071,N_3808);
nand U5175 (N_5175,N_3771,N_3927);
and U5176 (N_5176,N_3975,N_3964);
and U5177 (N_5177,N_3942,N_4081);
nand U5178 (N_5178,N_3958,N_3900);
nor U5179 (N_5179,N_4121,N_4297);
xnor U5180 (N_5180,N_3989,N_4188);
or U5181 (N_5181,N_4225,N_4420);
nand U5182 (N_5182,N_4288,N_4316);
and U5183 (N_5183,N_3961,N_3979);
and U5184 (N_5184,N_4139,N_4410);
nor U5185 (N_5185,N_4197,N_3978);
nand U5186 (N_5186,N_4075,N_4290);
and U5187 (N_5187,N_4209,N_3831);
nand U5188 (N_5188,N_4385,N_4163);
nand U5189 (N_5189,N_3878,N_3920);
nand U5190 (N_5190,N_4454,N_3993);
nand U5191 (N_5191,N_3846,N_4290);
and U5192 (N_5192,N_3886,N_3944);
and U5193 (N_5193,N_4285,N_3791);
nand U5194 (N_5194,N_4042,N_4212);
and U5195 (N_5195,N_4111,N_3836);
and U5196 (N_5196,N_4275,N_4367);
or U5197 (N_5197,N_4108,N_4071);
xnor U5198 (N_5198,N_4427,N_3825);
and U5199 (N_5199,N_4261,N_4241);
nand U5200 (N_5200,N_4050,N_4431);
nand U5201 (N_5201,N_3833,N_4088);
nor U5202 (N_5202,N_4045,N_4013);
nand U5203 (N_5203,N_4086,N_4243);
and U5204 (N_5204,N_4413,N_3859);
and U5205 (N_5205,N_4167,N_4325);
or U5206 (N_5206,N_4057,N_4103);
nor U5207 (N_5207,N_4417,N_4243);
nor U5208 (N_5208,N_4215,N_4225);
nand U5209 (N_5209,N_3862,N_3972);
nand U5210 (N_5210,N_3754,N_3763);
or U5211 (N_5211,N_3833,N_4355);
nand U5212 (N_5212,N_4345,N_3996);
or U5213 (N_5213,N_4044,N_4085);
xor U5214 (N_5214,N_4123,N_4439);
nor U5215 (N_5215,N_4220,N_4271);
xor U5216 (N_5216,N_4236,N_4270);
nand U5217 (N_5217,N_4466,N_3889);
or U5218 (N_5218,N_3895,N_4263);
xnor U5219 (N_5219,N_4476,N_4291);
or U5220 (N_5220,N_4110,N_4168);
and U5221 (N_5221,N_4054,N_3754);
and U5222 (N_5222,N_3940,N_3998);
and U5223 (N_5223,N_3774,N_4320);
nor U5224 (N_5224,N_4383,N_3857);
or U5225 (N_5225,N_4047,N_4281);
or U5226 (N_5226,N_4138,N_4178);
nor U5227 (N_5227,N_4466,N_4272);
and U5228 (N_5228,N_4068,N_4252);
and U5229 (N_5229,N_3964,N_4225);
nand U5230 (N_5230,N_3798,N_3797);
or U5231 (N_5231,N_4114,N_4001);
or U5232 (N_5232,N_4234,N_3830);
nand U5233 (N_5233,N_3790,N_3763);
nor U5234 (N_5234,N_3969,N_4233);
nor U5235 (N_5235,N_3914,N_4086);
nand U5236 (N_5236,N_4027,N_4002);
or U5237 (N_5237,N_4425,N_3757);
or U5238 (N_5238,N_4137,N_4436);
xnor U5239 (N_5239,N_4053,N_4308);
nor U5240 (N_5240,N_4107,N_4178);
and U5241 (N_5241,N_4081,N_3906);
and U5242 (N_5242,N_3904,N_4218);
xnor U5243 (N_5243,N_3926,N_4035);
or U5244 (N_5244,N_4128,N_3939);
nand U5245 (N_5245,N_4416,N_3911);
nand U5246 (N_5246,N_4404,N_4123);
and U5247 (N_5247,N_3997,N_4115);
or U5248 (N_5248,N_4198,N_3914);
and U5249 (N_5249,N_4301,N_4317);
nor U5250 (N_5250,N_5199,N_4983);
or U5251 (N_5251,N_5150,N_4782);
nand U5252 (N_5252,N_5098,N_5170);
nor U5253 (N_5253,N_4834,N_4584);
and U5254 (N_5254,N_4916,N_4747);
nand U5255 (N_5255,N_5180,N_4577);
xnor U5256 (N_5256,N_5100,N_5084);
and U5257 (N_5257,N_4849,N_5018);
nand U5258 (N_5258,N_4912,N_4836);
nor U5259 (N_5259,N_5169,N_4940);
and U5260 (N_5260,N_5207,N_5174);
nand U5261 (N_5261,N_4814,N_4588);
nand U5262 (N_5262,N_4926,N_5079);
nor U5263 (N_5263,N_5037,N_4874);
nor U5264 (N_5264,N_5177,N_4969);
or U5265 (N_5265,N_5022,N_4633);
or U5266 (N_5266,N_4761,N_4949);
xnor U5267 (N_5267,N_4530,N_5017);
xnor U5268 (N_5268,N_4925,N_4629);
xor U5269 (N_5269,N_4739,N_4723);
or U5270 (N_5270,N_5095,N_4552);
or U5271 (N_5271,N_4928,N_4649);
nor U5272 (N_5272,N_4707,N_5025);
or U5273 (N_5273,N_4920,N_5183);
nand U5274 (N_5274,N_4578,N_4771);
xnor U5275 (N_5275,N_4958,N_4915);
nand U5276 (N_5276,N_5141,N_4770);
and U5277 (N_5277,N_4561,N_5146);
or U5278 (N_5278,N_4564,N_4944);
nor U5279 (N_5279,N_5126,N_4837);
nor U5280 (N_5280,N_4955,N_4568);
and U5281 (N_5281,N_5237,N_4807);
and U5282 (N_5282,N_4891,N_5056);
nor U5283 (N_5283,N_4674,N_4914);
or U5284 (N_5284,N_4556,N_4678);
xor U5285 (N_5285,N_4877,N_5078);
xnor U5286 (N_5286,N_4878,N_5165);
and U5287 (N_5287,N_4541,N_4742);
or U5288 (N_5288,N_5092,N_4614);
xor U5289 (N_5289,N_4850,N_4979);
nand U5290 (N_5290,N_4795,N_4858);
or U5291 (N_5291,N_4731,N_5233);
nor U5292 (N_5292,N_4722,N_4519);
nor U5293 (N_5293,N_4845,N_5039);
or U5294 (N_5294,N_4816,N_5023);
and U5295 (N_5295,N_4655,N_4562);
nor U5296 (N_5296,N_5052,N_5154);
or U5297 (N_5297,N_4996,N_4968);
and U5298 (N_5298,N_4610,N_4734);
nand U5299 (N_5299,N_4937,N_5038);
and U5300 (N_5300,N_5239,N_4957);
nand U5301 (N_5301,N_4804,N_4802);
and U5302 (N_5302,N_4607,N_4744);
and U5303 (N_5303,N_5124,N_5107);
nor U5304 (N_5304,N_4531,N_4886);
and U5305 (N_5305,N_4605,N_5195);
nor U5306 (N_5306,N_4775,N_5031);
or U5307 (N_5307,N_5216,N_4870);
and U5308 (N_5308,N_4794,N_4786);
and U5309 (N_5309,N_5064,N_4772);
nor U5310 (N_5310,N_4812,N_5134);
nor U5311 (N_5311,N_4576,N_4583);
nand U5312 (N_5312,N_4835,N_4557);
and U5313 (N_5313,N_4932,N_4948);
xor U5314 (N_5314,N_4791,N_5116);
nand U5315 (N_5315,N_4999,N_4977);
or U5316 (N_5316,N_4729,N_4660);
or U5317 (N_5317,N_4543,N_4662);
or U5318 (N_5318,N_4820,N_4934);
and U5319 (N_5319,N_4799,N_5155);
and U5320 (N_5320,N_5227,N_5244);
nand U5321 (N_5321,N_5228,N_5118);
xnor U5322 (N_5322,N_4535,N_4567);
and U5323 (N_5323,N_5226,N_4696);
nor U5324 (N_5324,N_4666,N_4512);
and U5325 (N_5325,N_5058,N_5119);
or U5326 (N_5326,N_4751,N_4560);
xnor U5327 (N_5327,N_4887,N_5127);
or U5328 (N_5328,N_4581,N_5247);
and U5329 (N_5329,N_5062,N_5162);
and U5330 (N_5330,N_5070,N_4652);
nor U5331 (N_5331,N_4600,N_4943);
or U5332 (N_5332,N_4901,N_5212);
and U5333 (N_5333,N_5220,N_5171);
or U5334 (N_5334,N_5158,N_5222);
xor U5335 (N_5335,N_4956,N_4621);
or U5336 (N_5336,N_4762,N_4670);
xnor U5337 (N_5337,N_4749,N_4873);
or U5338 (N_5338,N_4532,N_4505);
xnor U5339 (N_5339,N_4963,N_4709);
nand U5340 (N_5340,N_4683,N_5179);
and U5341 (N_5341,N_5219,N_4755);
or U5342 (N_5342,N_4947,N_4563);
nor U5343 (N_5343,N_4654,N_5202);
nand U5344 (N_5344,N_4668,N_4767);
and U5345 (N_5345,N_5043,N_4718);
nand U5346 (N_5346,N_4672,N_4608);
or U5347 (N_5347,N_4743,N_4766);
or U5348 (N_5348,N_4951,N_4641);
and U5349 (N_5349,N_4950,N_4647);
or U5350 (N_5350,N_4974,N_4753);
nand U5351 (N_5351,N_4504,N_5235);
nand U5352 (N_5352,N_4981,N_4656);
nor U5353 (N_5353,N_5218,N_5131);
nand U5354 (N_5354,N_5080,N_5196);
or U5355 (N_5355,N_4871,N_4622);
or U5356 (N_5356,N_4876,N_5099);
nand U5357 (N_5357,N_4645,N_4521);
and U5358 (N_5358,N_4857,N_4788);
or U5359 (N_5359,N_4803,N_4975);
and U5360 (N_5360,N_4680,N_4516);
and U5361 (N_5361,N_5164,N_4922);
nand U5362 (N_5362,N_5013,N_4919);
and U5363 (N_5363,N_5113,N_4756);
nor U5364 (N_5364,N_4569,N_5000);
and U5365 (N_5365,N_4571,N_5125);
and U5366 (N_5366,N_5168,N_4590);
or U5367 (N_5367,N_4900,N_5190);
nor U5368 (N_5368,N_4980,N_5024);
or U5369 (N_5369,N_4965,N_5230);
or U5370 (N_5370,N_4995,N_4677);
and U5371 (N_5371,N_5248,N_4663);
or U5372 (N_5372,N_4710,N_5152);
and U5373 (N_5373,N_4936,N_4801);
xnor U5374 (N_5374,N_5065,N_4898);
or U5375 (N_5375,N_4962,N_4537);
nor U5376 (N_5376,N_4574,N_4748);
xnor U5377 (N_5377,N_4808,N_4973);
and U5378 (N_5378,N_4502,N_4661);
nor U5379 (N_5379,N_5192,N_4851);
nor U5380 (N_5380,N_5012,N_4904);
nand U5381 (N_5381,N_4597,N_5057);
xor U5382 (N_5382,N_4931,N_4517);
nor U5383 (N_5383,N_4524,N_4905);
nor U5384 (N_5384,N_4635,N_4752);
and U5385 (N_5385,N_4800,N_5225);
and U5386 (N_5386,N_4902,N_4736);
or U5387 (N_5387,N_5175,N_4503);
nand U5388 (N_5388,N_4550,N_4889);
xnor U5389 (N_5389,N_5145,N_5121);
or U5390 (N_5390,N_4509,N_5209);
nand U5391 (N_5391,N_4759,N_4695);
or U5392 (N_5392,N_4903,N_5087);
nor U5393 (N_5393,N_4927,N_4826);
and U5394 (N_5394,N_4859,N_5123);
or U5395 (N_5395,N_5231,N_4658);
and U5396 (N_5396,N_4872,N_4664);
nor U5397 (N_5397,N_4544,N_5198);
and U5398 (N_5398,N_5243,N_5019);
nor U5399 (N_5399,N_5001,N_4684);
nor U5400 (N_5400,N_4997,N_4785);
nor U5401 (N_5401,N_4982,N_4539);
or U5402 (N_5402,N_4885,N_5120);
nor U5403 (N_5403,N_4637,N_4908);
nand U5404 (N_5404,N_4650,N_4976);
or U5405 (N_5405,N_4860,N_4685);
and U5406 (N_5406,N_5197,N_4619);
and U5407 (N_5407,N_5185,N_4783);
nand U5408 (N_5408,N_5232,N_4513);
and U5409 (N_5409,N_4838,N_4642);
or U5410 (N_5410,N_4768,N_4899);
and U5411 (N_5411,N_4548,N_4894);
and U5412 (N_5412,N_4793,N_5030);
nor U5413 (N_5413,N_5090,N_4805);
and U5414 (N_5414,N_4594,N_5004);
or U5415 (N_5415,N_5149,N_4700);
and U5416 (N_5416,N_5096,N_5033);
and U5417 (N_5417,N_4776,N_5073);
nand U5418 (N_5418,N_5105,N_4865);
nor U5419 (N_5419,N_5094,N_4853);
nand U5420 (N_5420,N_4843,N_4972);
or U5421 (N_5421,N_5035,N_4525);
nor U5422 (N_5422,N_4618,N_4985);
or U5423 (N_5423,N_4689,N_4945);
and U5424 (N_5424,N_4881,N_5083);
nand U5425 (N_5425,N_4699,N_5009);
nand U5426 (N_5426,N_4713,N_4546);
and U5427 (N_5427,N_4551,N_4702);
xor U5428 (N_5428,N_5234,N_4798);
nand U5429 (N_5429,N_4971,N_4646);
nand U5430 (N_5430,N_4632,N_4690);
nor U5431 (N_5431,N_4825,N_5224);
or U5432 (N_5432,N_4848,N_4716);
nand U5433 (N_5433,N_4828,N_5172);
and U5434 (N_5434,N_4986,N_4549);
nand U5435 (N_5435,N_5173,N_4724);
nand U5436 (N_5436,N_4827,N_4855);
xnor U5437 (N_5437,N_5122,N_4818);
nor U5438 (N_5438,N_4523,N_4946);
or U5439 (N_5439,N_5028,N_4765);
or U5440 (N_5440,N_5114,N_5130);
or U5441 (N_5441,N_4964,N_4844);
nor U5442 (N_5442,N_4676,N_4579);
and U5443 (N_5443,N_5238,N_4994);
and U5444 (N_5444,N_4725,N_5111);
and U5445 (N_5445,N_4693,N_5045);
and U5446 (N_5446,N_4792,N_4721);
nand U5447 (N_5447,N_4712,N_5157);
and U5448 (N_5448,N_4869,N_4789);
nor U5449 (N_5449,N_5159,N_4659);
or U5450 (N_5450,N_4510,N_5178);
or U5451 (N_5451,N_4806,N_4960);
xor U5452 (N_5452,N_4784,N_4728);
xnor U5453 (N_5453,N_4854,N_4592);
and U5454 (N_5454,N_4617,N_5129);
and U5455 (N_5455,N_4778,N_4813);
nand U5456 (N_5456,N_5211,N_5215);
nor U5457 (N_5457,N_4604,N_5191);
and U5458 (N_5458,N_4711,N_4763);
nand U5459 (N_5459,N_4547,N_4634);
nand U5460 (N_5460,N_4984,N_4821);
or U5461 (N_5461,N_4954,N_4745);
and U5462 (N_5462,N_4679,N_5132);
and U5463 (N_5463,N_4918,N_4738);
xnor U5464 (N_5464,N_4686,N_5074);
or U5465 (N_5465,N_5151,N_5068);
or U5466 (N_5466,N_5214,N_4787);
nor U5467 (N_5467,N_4575,N_4720);
nand U5468 (N_5468,N_4780,N_4582);
or U5469 (N_5469,N_5048,N_4671);
xor U5470 (N_5470,N_4609,N_4832);
nand U5471 (N_5471,N_5104,N_4913);
or U5472 (N_5472,N_4796,N_4625);
nand U5473 (N_5473,N_4890,N_5036);
nand U5474 (N_5474,N_4687,N_4697);
nand U5475 (N_5475,N_5072,N_5088);
or U5476 (N_5476,N_4536,N_5042);
or U5477 (N_5477,N_4911,N_4884);
or U5478 (N_5478,N_4847,N_4760);
nand U5479 (N_5479,N_5176,N_4846);
nand U5480 (N_5480,N_4545,N_4566);
nor U5481 (N_5481,N_4856,N_4506);
nor U5482 (N_5482,N_5201,N_5147);
and U5483 (N_5483,N_5143,N_4555);
nand U5484 (N_5484,N_4777,N_4852);
or U5485 (N_5485,N_5186,N_4917);
nand U5486 (N_5486,N_4735,N_4893);
nor U5487 (N_5487,N_4511,N_5040);
xor U5488 (N_5488,N_4602,N_4737);
nor U5489 (N_5489,N_4809,N_4669);
nor U5490 (N_5490,N_4892,N_5246);
nor U5491 (N_5491,N_4630,N_4703);
xnor U5492 (N_5492,N_5139,N_4998);
nor U5493 (N_5493,N_5229,N_4640);
nand U5494 (N_5494,N_4682,N_4623);
and U5495 (N_5495,N_4790,N_4624);
xor U5496 (N_5496,N_5067,N_4559);
and U5497 (N_5497,N_4528,N_4830);
xor U5498 (N_5498,N_5140,N_4741);
nor U5499 (N_5499,N_4714,N_4500);
and U5500 (N_5500,N_5051,N_5245);
xor U5501 (N_5501,N_4921,N_5187);
and U5502 (N_5502,N_4888,N_4585);
nand U5503 (N_5503,N_5066,N_4797);
nor U5504 (N_5504,N_4540,N_4839);
nand U5505 (N_5505,N_4615,N_4616);
nor U5506 (N_5506,N_4701,N_4518);
nand U5507 (N_5507,N_5213,N_4638);
nand U5508 (N_5508,N_5054,N_5206);
nor U5509 (N_5509,N_4819,N_5110);
nand U5510 (N_5510,N_5049,N_4875);
nor U5511 (N_5511,N_4817,N_4740);
xor U5512 (N_5512,N_5076,N_4961);
or U5513 (N_5513,N_5027,N_5005);
and U5514 (N_5514,N_5046,N_4620);
and U5515 (N_5515,N_4598,N_4757);
nor U5516 (N_5516,N_4715,N_4599);
nor U5517 (N_5517,N_4823,N_4591);
nand U5518 (N_5518,N_4930,N_5204);
nor U5519 (N_5519,N_5117,N_4681);
and U5520 (N_5520,N_4935,N_5137);
xor U5521 (N_5521,N_4589,N_5029);
or U5522 (N_5522,N_4522,N_4596);
xnor U5523 (N_5523,N_5091,N_5106);
and U5524 (N_5524,N_4508,N_4730);
xor U5525 (N_5525,N_4942,N_4811);
nand U5526 (N_5526,N_4673,N_4570);
and U5527 (N_5527,N_4626,N_5184);
or U5528 (N_5528,N_5205,N_5240);
or U5529 (N_5529,N_4520,N_5026);
nor U5530 (N_5530,N_5142,N_5167);
nor U5531 (N_5531,N_5016,N_4527);
and U5532 (N_5532,N_5020,N_5182);
nand U5533 (N_5533,N_4978,N_4572);
nor U5534 (N_5534,N_4657,N_4705);
or U5535 (N_5535,N_4933,N_4636);
nand U5536 (N_5536,N_5181,N_5103);
nor U5537 (N_5537,N_5002,N_4769);
and U5538 (N_5538,N_4580,N_5010);
and U5539 (N_5539,N_4907,N_5102);
nand U5540 (N_5540,N_4959,N_5200);
and U5541 (N_5541,N_5093,N_4515);
nor U5542 (N_5542,N_4953,N_5208);
and U5543 (N_5543,N_4829,N_4929);
xor U5544 (N_5544,N_4606,N_4704);
nand U5545 (N_5545,N_5148,N_4558);
and U5546 (N_5546,N_4727,N_4708);
or U5547 (N_5547,N_4732,N_5041);
nor U5548 (N_5548,N_4627,N_5210);
nor U5549 (N_5549,N_5249,N_4868);
and U5550 (N_5550,N_4896,N_5101);
nand U5551 (N_5551,N_4653,N_5161);
or U5552 (N_5552,N_4565,N_5108);
nor U5553 (N_5553,N_5060,N_4861);
or U5554 (N_5554,N_5189,N_5144);
xor U5555 (N_5555,N_4613,N_5003);
and U5556 (N_5556,N_4692,N_4746);
xnor U5557 (N_5557,N_4906,N_4651);
or U5558 (N_5558,N_4992,N_4758);
nand U5559 (N_5559,N_4824,N_5241);
nor U5560 (N_5560,N_5085,N_4750);
nand U5561 (N_5561,N_5236,N_4601);
nor U5562 (N_5562,N_4967,N_5194);
or U5563 (N_5563,N_5086,N_4773);
nor U5564 (N_5564,N_5008,N_4810);
nand U5565 (N_5565,N_4612,N_4923);
nand U5566 (N_5566,N_4815,N_4573);
nand U5567 (N_5567,N_5021,N_4688);
nor U5568 (N_5568,N_4822,N_4970);
and U5569 (N_5569,N_5193,N_5109);
xor U5570 (N_5570,N_4533,N_4754);
xnor U5571 (N_5571,N_5156,N_4526);
nand U5572 (N_5572,N_4507,N_4726);
and U5573 (N_5573,N_4833,N_5007);
nor U5574 (N_5574,N_4866,N_5135);
nand U5575 (N_5575,N_5014,N_4764);
nand U5576 (N_5576,N_4542,N_4840);
nand U5577 (N_5577,N_4534,N_4648);
nand U5578 (N_5578,N_4966,N_4991);
nand U5579 (N_5579,N_4595,N_4939);
nand U5580 (N_5580,N_5059,N_4779);
nand U5581 (N_5581,N_5011,N_5055);
nor U5582 (N_5582,N_5050,N_5032);
nor U5583 (N_5583,N_4593,N_4628);
nand U5584 (N_5584,N_4987,N_5112);
xor U5585 (N_5585,N_5188,N_4694);
nor U5586 (N_5586,N_4538,N_4611);
and U5587 (N_5587,N_4842,N_5077);
or U5588 (N_5588,N_4988,N_4501);
or U5589 (N_5589,N_4895,N_4880);
nand U5590 (N_5590,N_5138,N_4924);
xnor U5591 (N_5591,N_4774,N_4675);
and U5592 (N_5592,N_4879,N_4719);
or U5593 (N_5593,N_4990,N_5242);
nand U5594 (N_5594,N_5015,N_4883);
nand U5595 (N_5595,N_4553,N_4665);
or U5596 (N_5596,N_5047,N_5115);
or U5597 (N_5597,N_5153,N_4882);
and U5598 (N_5598,N_5097,N_4781);
nand U5599 (N_5599,N_4952,N_5163);
nor U5600 (N_5600,N_4603,N_5006);
or U5601 (N_5601,N_5217,N_4909);
nor U5602 (N_5602,N_5075,N_5203);
or U5603 (N_5603,N_4831,N_4639);
and U5604 (N_5604,N_4554,N_4529);
nor U5605 (N_5605,N_5166,N_5128);
nand U5606 (N_5606,N_5089,N_4989);
nand U5607 (N_5607,N_4863,N_5061);
nor U5608 (N_5608,N_4514,N_4587);
xor U5609 (N_5609,N_5221,N_5136);
or U5610 (N_5610,N_4586,N_4667);
or U5611 (N_5611,N_4698,N_4644);
and U5612 (N_5612,N_5063,N_4733);
or U5613 (N_5613,N_4643,N_5160);
nor U5614 (N_5614,N_4631,N_4938);
nor U5615 (N_5615,N_4867,N_4897);
and U5616 (N_5616,N_5081,N_5133);
nand U5617 (N_5617,N_5223,N_4993);
and U5618 (N_5618,N_4864,N_4910);
and U5619 (N_5619,N_4717,N_4841);
and U5620 (N_5620,N_5034,N_5082);
and U5621 (N_5621,N_5069,N_5053);
and U5622 (N_5622,N_5044,N_4862);
or U5623 (N_5623,N_4941,N_4691);
or U5624 (N_5624,N_5071,N_4706);
or U5625 (N_5625,N_4662,N_4876);
or U5626 (N_5626,N_4621,N_5096);
or U5627 (N_5627,N_4607,N_4907);
nor U5628 (N_5628,N_4511,N_5211);
and U5629 (N_5629,N_4663,N_5202);
nor U5630 (N_5630,N_5095,N_4638);
nor U5631 (N_5631,N_4734,N_5238);
or U5632 (N_5632,N_4761,N_4619);
and U5633 (N_5633,N_4950,N_4710);
nand U5634 (N_5634,N_5234,N_5170);
or U5635 (N_5635,N_5072,N_5242);
xor U5636 (N_5636,N_4606,N_4819);
nor U5637 (N_5637,N_4788,N_5110);
xor U5638 (N_5638,N_5142,N_5148);
and U5639 (N_5639,N_4604,N_4535);
nand U5640 (N_5640,N_4768,N_4616);
or U5641 (N_5641,N_4851,N_4877);
nor U5642 (N_5642,N_4576,N_4784);
nand U5643 (N_5643,N_4504,N_5039);
nor U5644 (N_5644,N_4538,N_5216);
and U5645 (N_5645,N_5011,N_4993);
nand U5646 (N_5646,N_4652,N_4976);
or U5647 (N_5647,N_4698,N_4583);
or U5648 (N_5648,N_4767,N_4823);
nor U5649 (N_5649,N_4757,N_4707);
nand U5650 (N_5650,N_4619,N_4671);
nand U5651 (N_5651,N_4924,N_4846);
or U5652 (N_5652,N_4954,N_5046);
nand U5653 (N_5653,N_4845,N_4972);
and U5654 (N_5654,N_5016,N_5067);
nand U5655 (N_5655,N_4819,N_4539);
and U5656 (N_5656,N_5248,N_4766);
xor U5657 (N_5657,N_4977,N_4515);
nor U5658 (N_5658,N_4881,N_4539);
nand U5659 (N_5659,N_4636,N_5089);
and U5660 (N_5660,N_4539,N_5104);
or U5661 (N_5661,N_5164,N_4542);
nand U5662 (N_5662,N_4675,N_5031);
and U5663 (N_5663,N_4946,N_5009);
or U5664 (N_5664,N_4807,N_4884);
nor U5665 (N_5665,N_5136,N_4608);
nand U5666 (N_5666,N_4570,N_4606);
and U5667 (N_5667,N_4758,N_4771);
xor U5668 (N_5668,N_5055,N_4557);
and U5669 (N_5669,N_4739,N_4710);
and U5670 (N_5670,N_5178,N_4809);
xor U5671 (N_5671,N_5062,N_5040);
and U5672 (N_5672,N_4839,N_4860);
and U5673 (N_5673,N_5117,N_4939);
nand U5674 (N_5674,N_4581,N_5141);
nand U5675 (N_5675,N_4744,N_4678);
and U5676 (N_5676,N_5126,N_4848);
nor U5677 (N_5677,N_4988,N_4788);
or U5678 (N_5678,N_4537,N_5056);
and U5679 (N_5679,N_4881,N_4569);
nor U5680 (N_5680,N_4599,N_5040);
and U5681 (N_5681,N_4927,N_5030);
xor U5682 (N_5682,N_4721,N_4584);
nand U5683 (N_5683,N_5049,N_4659);
nand U5684 (N_5684,N_4718,N_4511);
xor U5685 (N_5685,N_4562,N_4540);
xor U5686 (N_5686,N_5074,N_5217);
nand U5687 (N_5687,N_4672,N_5176);
or U5688 (N_5688,N_5066,N_4610);
or U5689 (N_5689,N_5125,N_5024);
nand U5690 (N_5690,N_5042,N_5033);
xor U5691 (N_5691,N_4683,N_4511);
xor U5692 (N_5692,N_5085,N_4644);
nor U5693 (N_5693,N_5011,N_5086);
and U5694 (N_5694,N_5133,N_4787);
or U5695 (N_5695,N_4753,N_5242);
nand U5696 (N_5696,N_5183,N_4824);
nand U5697 (N_5697,N_5118,N_4888);
nand U5698 (N_5698,N_4984,N_4521);
nor U5699 (N_5699,N_5112,N_4595);
and U5700 (N_5700,N_4583,N_5142);
nor U5701 (N_5701,N_5154,N_4970);
and U5702 (N_5702,N_4532,N_4858);
and U5703 (N_5703,N_4817,N_4528);
nor U5704 (N_5704,N_4627,N_5051);
or U5705 (N_5705,N_4864,N_4697);
xnor U5706 (N_5706,N_5030,N_5211);
and U5707 (N_5707,N_4533,N_4661);
or U5708 (N_5708,N_5099,N_4595);
nand U5709 (N_5709,N_5028,N_4684);
xnor U5710 (N_5710,N_5024,N_4855);
nand U5711 (N_5711,N_4898,N_4713);
and U5712 (N_5712,N_5213,N_4628);
nand U5713 (N_5713,N_4512,N_5113);
or U5714 (N_5714,N_4821,N_4657);
nor U5715 (N_5715,N_4642,N_5243);
nand U5716 (N_5716,N_4647,N_5212);
nor U5717 (N_5717,N_4526,N_5155);
nand U5718 (N_5718,N_5104,N_4976);
or U5719 (N_5719,N_5213,N_5170);
or U5720 (N_5720,N_4926,N_5244);
nand U5721 (N_5721,N_4625,N_5137);
nor U5722 (N_5722,N_4933,N_5001);
and U5723 (N_5723,N_4671,N_4614);
or U5724 (N_5724,N_4540,N_5023);
nand U5725 (N_5725,N_4747,N_5082);
and U5726 (N_5726,N_5002,N_4753);
or U5727 (N_5727,N_4856,N_4766);
nand U5728 (N_5728,N_5163,N_4956);
or U5729 (N_5729,N_5188,N_4598);
nand U5730 (N_5730,N_4679,N_4776);
nand U5731 (N_5731,N_5239,N_4623);
nand U5732 (N_5732,N_5188,N_4672);
and U5733 (N_5733,N_4856,N_4787);
nor U5734 (N_5734,N_5050,N_4886);
and U5735 (N_5735,N_5149,N_5051);
or U5736 (N_5736,N_4899,N_4733);
or U5737 (N_5737,N_5103,N_4922);
nand U5738 (N_5738,N_4908,N_5235);
and U5739 (N_5739,N_5125,N_5190);
nor U5740 (N_5740,N_5187,N_4580);
or U5741 (N_5741,N_4724,N_4816);
nor U5742 (N_5742,N_4822,N_5082);
nor U5743 (N_5743,N_4601,N_4974);
and U5744 (N_5744,N_4990,N_5043);
xnor U5745 (N_5745,N_5007,N_5197);
and U5746 (N_5746,N_4567,N_5130);
or U5747 (N_5747,N_4997,N_4616);
nand U5748 (N_5748,N_5020,N_5032);
nand U5749 (N_5749,N_4786,N_4820);
and U5750 (N_5750,N_5023,N_5082);
nor U5751 (N_5751,N_4531,N_4938);
nand U5752 (N_5752,N_5240,N_5226);
nand U5753 (N_5753,N_4626,N_4905);
or U5754 (N_5754,N_4811,N_5032);
and U5755 (N_5755,N_5140,N_4881);
or U5756 (N_5756,N_4852,N_4986);
or U5757 (N_5757,N_4805,N_5232);
xnor U5758 (N_5758,N_4845,N_5148);
and U5759 (N_5759,N_5221,N_4721);
and U5760 (N_5760,N_4559,N_4779);
nor U5761 (N_5761,N_5170,N_4964);
nor U5762 (N_5762,N_4574,N_5153);
or U5763 (N_5763,N_4669,N_5081);
nand U5764 (N_5764,N_4531,N_4629);
nand U5765 (N_5765,N_4612,N_4653);
nand U5766 (N_5766,N_5111,N_5220);
nor U5767 (N_5767,N_5044,N_5091);
or U5768 (N_5768,N_4557,N_4763);
xnor U5769 (N_5769,N_4793,N_4826);
nor U5770 (N_5770,N_4878,N_4595);
or U5771 (N_5771,N_4578,N_5101);
nand U5772 (N_5772,N_4677,N_4768);
nor U5773 (N_5773,N_5102,N_5061);
xnor U5774 (N_5774,N_4660,N_4917);
nand U5775 (N_5775,N_4515,N_4804);
nor U5776 (N_5776,N_4981,N_5209);
and U5777 (N_5777,N_4968,N_4505);
nand U5778 (N_5778,N_4704,N_4503);
and U5779 (N_5779,N_4502,N_4703);
nand U5780 (N_5780,N_4824,N_4589);
nor U5781 (N_5781,N_5008,N_4947);
nor U5782 (N_5782,N_4983,N_4779);
or U5783 (N_5783,N_5174,N_4914);
or U5784 (N_5784,N_4556,N_4955);
nand U5785 (N_5785,N_5217,N_4667);
nor U5786 (N_5786,N_5202,N_4782);
and U5787 (N_5787,N_4618,N_4950);
nand U5788 (N_5788,N_5235,N_4596);
nor U5789 (N_5789,N_4538,N_5084);
and U5790 (N_5790,N_5150,N_4513);
or U5791 (N_5791,N_4691,N_4722);
nor U5792 (N_5792,N_4813,N_4788);
nand U5793 (N_5793,N_4910,N_5078);
nor U5794 (N_5794,N_4670,N_5082);
nand U5795 (N_5795,N_4531,N_4971);
nand U5796 (N_5796,N_4632,N_4521);
nor U5797 (N_5797,N_5153,N_4559);
and U5798 (N_5798,N_4830,N_4509);
nand U5799 (N_5799,N_4804,N_4645);
nor U5800 (N_5800,N_4800,N_5021);
or U5801 (N_5801,N_4829,N_4928);
xor U5802 (N_5802,N_4679,N_5224);
and U5803 (N_5803,N_5047,N_5160);
and U5804 (N_5804,N_4655,N_4874);
xor U5805 (N_5805,N_5128,N_5218);
or U5806 (N_5806,N_5137,N_4724);
nand U5807 (N_5807,N_4727,N_4996);
nor U5808 (N_5808,N_4797,N_5232);
xnor U5809 (N_5809,N_4858,N_4974);
nand U5810 (N_5810,N_4772,N_4963);
nor U5811 (N_5811,N_5194,N_4910);
nor U5812 (N_5812,N_5244,N_4618);
and U5813 (N_5813,N_4824,N_5126);
nor U5814 (N_5814,N_5244,N_4886);
nor U5815 (N_5815,N_5110,N_5103);
or U5816 (N_5816,N_5236,N_4960);
and U5817 (N_5817,N_5121,N_4585);
nand U5818 (N_5818,N_5050,N_4851);
nand U5819 (N_5819,N_4902,N_5054);
or U5820 (N_5820,N_4502,N_4769);
xnor U5821 (N_5821,N_4900,N_4799);
nand U5822 (N_5822,N_4642,N_5175);
nand U5823 (N_5823,N_4811,N_4567);
and U5824 (N_5824,N_4608,N_5085);
and U5825 (N_5825,N_5077,N_4975);
nor U5826 (N_5826,N_4730,N_5003);
or U5827 (N_5827,N_4682,N_4997);
nand U5828 (N_5828,N_4764,N_4832);
xor U5829 (N_5829,N_4949,N_5108);
xor U5830 (N_5830,N_5131,N_5165);
and U5831 (N_5831,N_4558,N_4675);
nor U5832 (N_5832,N_4789,N_5038);
xor U5833 (N_5833,N_5193,N_5234);
or U5834 (N_5834,N_4760,N_5179);
xnor U5835 (N_5835,N_4675,N_5224);
nor U5836 (N_5836,N_4730,N_4697);
or U5837 (N_5837,N_5221,N_5053);
or U5838 (N_5838,N_5101,N_4691);
nand U5839 (N_5839,N_5144,N_5098);
nand U5840 (N_5840,N_4741,N_5008);
and U5841 (N_5841,N_4786,N_4787);
nor U5842 (N_5842,N_4988,N_4866);
and U5843 (N_5843,N_4653,N_4522);
nand U5844 (N_5844,N_5139,N_5004);
or U5845 (N_5845,N_4848,N_4950);
nand U5846 (N_5846,N_5230,N_5155);
and U5847 (N_5847,N_4870,N_4892);
nand U5848 (N_5848,N_4975,N_4921);
or U5849 (N_5849,N_4571,N_4970);
xor U5850 (N_5850,N_5015,N_5001);
nand U5851 (N_5851,N_4703,N_5022);
or U5852 (N_5852,N_4987,N_4948);
or U5853 (N_5853,N_4566,N_4575);
or U5854 (N_5854,N_5035,N_4843);
nand U5855 (N_5855,N_5009,N_4804);
nand U5856 (N_5856,N_4668,N_4792);
or U5857 (N_5857,N_4913,N_5044);
nand U5858 (N_5858,N_4567,N_4880);
xor U5859 (N_5859,N_5234,N_4858);
nor U5860 (N_5860,N_5051,N_5017);
or U5861 (N_5861,N_4707,N_5071);
or U5862 (N_5862,N_4838,N_5226);
xnor U5863 (N_5863,N_5003,N_4694);
nand U5864 (N_5864,N_4894,N_4628);
or U5865 (N_5865,N_4513,N_4877);
and U5866 (N_5866,N_4565,N_4505);
nor U5867 (N_5867,N_4686,N_5188);
or U5868 (N_5868,N_4539,N_4589);
or U5869 (N_5869,N_4882,N_4928);
nand U5870 (N_5870,N_4558,N_4831);
nor U5871 (N_5871,N_5074,N_4972);
nand U5872 (N_5872,N_5012,N_4799);
and U5873 (N_5873,N_5154,N_4699);
and U5874 (N_5874,N_5063,N_4653);
or U5875 (N_5875,N_4511,N_4876);
xnor U5876 (N_5876,N_5108,N_4893);
and U5877 (N_5877,N_4513,N_4885);
and U5878 (N_5878,N_5163,N_5147);
nor U5879 (N_5879,N_4916,N_4822);
nor U5880 (N_5880,N_4972,N_4848);
and U5881 (N_5881,N_5043,N_4588);
xor U5882 (N_5882,N_4762,N_5136);
and U5883 (N_5883,N_4862,N_5169);
and U5884 (N_5884,N_4652,N_4847);
and U5885 (N_5885,N_4832,N_4701);
xor U5886 (N_5886,N_4886,N_5033);
nand U5887 (N_5887,N_4637,N_4785);
nand U5888 (N_5888,N_4644,N_5174);
nor U5889 (N_5889,N_5228,N_4948);
or U5890 (N_5890,N_4695,N_5091);
xor U5891 (N_5891,N_4541,N_4838);
nor U5892 (N_5892,N_5134,N_4810);
nor U5893 (N_5893,N_4994,N_4867);
or U5894 (N_5894,N_4514,N_5096);
nor U5895 (N_5895,N_5063,N_4800);
and U5896 (N_5896,N_4719,N_4968);
and U5897 (N_5897,N_4791,N_4977);
nor U5898 (N_5898,N_4893,N_4857);
nand U5899 (N_5899,N_5007,N_4592);
nor U5900 (N_5900,N_4915,N_5066);
nor U5901 (N_5901,N_5234,N_4543);
nor U5902 (N_5902,N_4695,N_4791);
or U5903 (N_5903,N_5062,N_4717);
and U5904 (N_5904,N_4976,N_5198);
or U5905 (N_5905,N_5058,N_4630);
or U5906 (N_5906,N_5186,N_5162);
or U5907 (N_5907,N_4620,N_4935);
nand U5908 (N_5908,N_4873,N_4988);
xnor U5909 (N_5909,N_4577,N_4696);
and U5910 (N_5910,N_5107,N_5114);
and U5911 (N_5911,N_5054,N_4821);
xor U5912 (N_5912,N_4542,N_5122);
nand U5913 (N_5913,N_5142,N_4683);
xnor U5914 (N_5914,N_4637,N_4880);
or U5915 (N_5915,N_4929,N_4559);
nor U5916 (N_5916,N_4597,N_4882);
nand U5917 (N_5917,N_5006,N_5051);
xor U5918 (N_5918,N_4935,N_4704);
xnor U5919 (N_5919,N_4849,N_5202);
and U5920 (N_5920,N_4644,N_4508);
xor U5921 (N_5921,N_5108,N_4513);
or U5922 (N_5922,N_4510,N_5049);
nand U5923 (N_5923,N_4555,N_4856);
or U5924 (N_5924,N_4569,N_4973);
nor U5925 (N_5925,N_4789,N_4800);
and U5926 (N_5926,N_4598,N_4630);
or U5927 (N_5927,N_5045,N_4607);
nand U5928 (N_5928,N_4939,N_4752);
and U5929 (N_5929,N_5183,N_5224);
and U5930 (N_5930,N_5045,N_4546);
nand U5931 (N_5931,N_4788,N_4901);
or U5932 (N_5932,N_5236,N_4817);
nor U5933 (N_5933,N_4888,N_5120);
nand U5934 (N_5934,N_4746,N_4502);
or U5935 (N_5935,N_4577,N_5121);
nand U5936 (N_5936,N_4693,N_4618);
nand U5937 (N_5937,N_4596,N_4563);
nor U5938 (N_5938,N_5019,N_4961);
nand U5939 (N_5939,N_5177,N_4932);
nor U5940 (N_5940,N_4792,N_4628);
nand U5941 (N_5941,N_4568,N_4907);
nand U5942 (N_5942,N_5127,N_4503);
nand U5943 (N_5943,N_5238,N_4764);
or U5944 (N_5944,N_5000,N_5174);
and U5945 (N_5945,N_4788,N_4892);
and U5946 (N_5946,N_4987,N_4674);
nor U5947 (N_5947,N_5241,N_4589);
nor U5948 (N_5948,N_4651,N_4588);
nand U5949 (N_5949,N_4838,N_5002);
nor U5950 (N_5950,N_5030,N_5128);
xnor U5951 (N_5951,N_4834,N_4759);
or U5952 (N_5952,N_5112,N_5211);
nand U5953 (N_5953,N_5045,N_4737);
nor U5954 (N_5954,N_4756,N_5120);
and U5955 (N_5955,N_5037,N_5195);
and U5956 (N_5956,N_4687,N_5161);
nor U5957 (N_5957,N_4656,N_4839);
nor U5958 (N_5958,N_5080,N_5090);
and U5959 (N_5959,N_4529,N_4703);
and U5960 (N_5960,N_5117,N_5170);
nor U5961 (N_5961,N_4682,N_5006);
nand U5962 (N_5962,N_4696,N_5231);
and U5963 (N_5963,N_5006,N_4714);
and U5964 (N_5964,N_5050,N_4892);
and U5965 (N_5965,N_4872,N_4836);
and U5966 (N_5966,N_4755,N_4893);
nor U5967 (N_5967,N_4625,N_4915);
and U5968 (N_5968,N_5202,N_5196);
and U5969 (N_5969,N_5148,N_5207);
or U5970 (N_5970,N_4898,N_4837);
nand U5971 (N_5971,N_5094,N_5085);
nor U5972 (N_5972,N_4744,N_4988);
nor U5973 (N_5973,N_5211,N_4885);
or U5974 (N_5974,N_4608,N_5239);
nor U5975 (N_5975,N_4738,N_5175);
or U5976 (N_5976,N_5242,N_5158);
and U5977 (N_5977,N_5163,N_4665);
nand U5978 (N_5978,N_4737,N_4967);
or U5979 (N_5979,N_5036,N_4682);
xor U5980 (N_5980,N_5205,N_4898);
xor U5981 (N_5981,N_5045,N_4651);
nand U5982 (N_5982,N_4747,N_4884);
xor U5983 (N_5983,N_4522,N_4657);
nand U5984 (N_5984,N_5031,N_5234);
and U5985 (N_5985,N_4854,N_5173);
nor U5986 (N_5986,N_5035,N_4882);
nand U5987 (N_5987,N_4770,N_4545);
and U5988 (N_5988,N_4819,N_5055);
xor U5989 (N_5989,N_4515,N_4917);
xor U5990 (N_5990,N_5194,N_4791);
or U5991 (N_5991,N_4532,N_4773);
or U5992 (N_5992,N_4659,N_4620);
xor U5993 (N_5993,N_4913,N_4788);
xor U5994 (N_5994,N_4762,N_4695);
or U5995 (N_5995,N_4969,N_4515);
xor U5996 (N_5996,N_5064,N_4992);
and U5997 (N_5997,N_4997,N_4791);
or U5998 (N_5998,N_4929,N_4505);
and U5999 (N_5999,N_4502,N_5083);
nand U6000 (N_6000,N_5789,N_5965);
and U6001 (N_6001,N_5498,N_5794);
and U6002 (N_6002,N_5730,N_5329);
nand U6003 (N_6003,N_5637,N_5301);
or U6004 (N_6004,N_5929,N_5455);
and U6005 (N_6005,N_5825,N_5355);
nor U6006 (N_6006,N_5641,N_5812);
or U6007 (N_6007,N_5733,N_5697);
nor U6008 (N_6008,N_5341,N_5468);
nand U6009 (N_6009,N_5738,N_5454);
and U6010 (N_6010,N_5257,N_5363);
nor U6011 (N_6011,N_5264,N_5484);
and U6012 (N_6012,N_5673,N_5419);
and U6013 (N_6013,N_5792,N_5376);
nor U6014 (N_6014,N_5763,N_5610);
or U6015 (N_6015,N_5816,N_5334);
or U6016 (N_6016,N_5584,N_5880);
nand U6017 (N_6017,N_5384,N_5606);
and U6018 (N_6018,N_5426,N_5749);
xor U6019 (N_6019,N_5715,N_5586);
nand U6020 (N_6020,N_5488,N_5342);
or U6021 (N_6021,N_5845,N_5971);
and U6022 (N_6022,N_5872,N_5949);
nand U6023 (N_6023,N_5897,N_5937);
nand U6024 (N_6024,N_5955,N_5809);
and U6025 (N_6025,N_5959,N_5609);
and U6026 (N_6026,N_5473,N_5755);
nand U6027 (N_6027,N_5983,N_5420);
nor U6028 (N_6028,N_5439,N_5267);
xnor U6029 (N_6029,N_5948,N_5817);
and U6030 (N_6030,N_5311,N_5492);
nand U6031 (N_6031,N_5408,N_5481);
and U6032 (N_6032,N_5616,N_5296);
or U6033 (N_6033,N_5379,N_5521);
nand U6034 (N_6034,N_5486,N_5266);
and U6035 (N_6035,N_5654,N_5427);
and U6036 (N_6036,N_5386,N_5768);
nor U6037 (N_6037,N_5953,N_5469);
nand U6038 (N_6038,N_5644,N_5935);
xor U6039 (N_6039,N_5819,N_5698);
nor U6040 (N_6040,N_5428,N_5784);
nand U6041 (N_6041,N_5592,N_5387);
nor U6042 (N_6042,N_5875,N_5448);
nor U6043 (N_6043,N_5307,N_5546);
nor U6044 (N_6044,N_5599,N_5289);
nor U6045 (N_6045,N_5677,N_5414);
or U6046 (N_6046,N_5745,N_5326);
or U6047 (N_6047,N_5262,N_5905);
nor U6048 (N_6048,N_5568,N_5801);
and U6049 (N_6049,N_5828,N_5936);
xor U6050 (N_6050,N_5751,N_5635);
nand U6051 (N_6051,N_5932,N_5783);
nand U6052 (N_6052,N_5518,N_5740);
xnor U6053 (N_6053,N_5761,N_5399);
or U6054 (N_6054,N_5696,N_5890);
and U6055 (N_6055,N_5645,N_5798);
nand U6056 (N_6056,N_5862,N_5618);
or U6057 (N_6057,N_5848,N_5833);
and U6058 (N_6058,N_5594,N_5602);
nand U6059 (N_6059,N_5779,N_5631);
nor U6060 (N_6060,N_5831,N_5829);
xnor U6061 (N_6061,N_5914,N_5791);
or U6062 (N_6062,N_5559,N_5578);
and U6063 (N_6063,N_5441,N_5500);
and U6064 (N_6064,N_5847,N_5709);
nor U6065 (N_6065,N_5368,N_5560);
nand U6066 (N_6066,N_5892,N_5389);
or U6067 (N_6067,N_5354,N_5417);
nor U6068 (N_6068,N_5748,N_5575);
nor U6069 (N_6069,N_5974,N_5646);
xor U6070 (N_6070,N_5997,N_5858);
nor U6071 (N_6071,N_5418,N_5256);
or U6072 (N_6072,N_5806,N_5515);
xnor U6073 (N_6073,N_5873,N_5667);
xor U6074 (N_6074,N_5450,N_5879);
and U6075 (N_6075,N_5917,N_5512);
nand U6076 (N_6076,N_5786,N_5352);
and U6077 (N_6077,N_5619,N_5920);
or U6078 (N_6078,N_5605,N_5639);
nor U6079 (N_6079,N_5429,N_5760);
or U6080 (N_6080,N_5550,N_5841);
and U6081 (N_6081,N_5561,N_5462);
xor U6082 (N_6082,N_5315,N_5885);
nand U6083 (N_6083,N_5291,N_5972);
or U6084 (N_6084,N_5889,N_5634);
xor U6085 (N_6085,N_5297,N_5514);
or U6086 (N_6086,N_5854,N_5620);
or U6087 (N_6087,N_5482,N_5451);
or U6088 (N_6088,N_5331,N_5799);
xnor U6089 (N_6089,N_5336,N_5440);
nor U6090 (N_6090,N_5981,N_5343);
and U6091 (N_6091,N_5520,N_5375);
and U6092 (N_6092,N_5501,N_5703);
nand U6093 (N_6093,N_5623,N_5907);
or U6094 (N_6094,N_5773,N_5431);
nand U6095 (N_6095,N_5765,N_5995);
or U6096 (N_6096,N_5716,N_5479);
and U6097 (N_6097,N_5403,N_5700);
and U6098 (N_6098,N_5571,N_5871);
or U6099 (N_6099,N_5360,N_5523);
xor U6100 (N_6100,N_5344,N_5538);
and U6101 (N_6101,N_5886,N_5485);
nand U6102 (N_6102,N_5593,N_5516);
and U6103 (N_6103,N_5710,N_5701);
nand U6104 (N_6104,N_5320,N_5377);
nand U6105 (N_6105,N_5392,N_5367);
xnor U6106 (N_6106,N_5306,N_5757);
or U6107 (N_6107,N_5969,N_5916);
or U6108 (N_6108,N_5928,N_5585);
nor U6109 (N_6109,N_5347,N_5261);
or U6110 (N_6110,N_5911,N_5985);
or U6111 (N_6111,N_5390,N_5883);
and U6112 (N_6112,N_5393,N_5857);
or U6113 (N_6113,N_5321,N_5443);
nor U6114 (N_6114,N_5310,N_5690);
nand U6115 (N_6115,N_5975,N_5723);
nand U6116 (N_6116,N_5470,N_5933);
or U6117 (N_6117,N_5976,N_5737);
xor U6118 (N_6118,N_5708,N_5365);
nand U6119 (N_6119,N_5569,N_5445);
nand U6120 (N_6120,N_5899,N_5581);
nand U6121 (N_6121,N_5351,N_5931);
nand U6122 (N_6122,N_5864,N_5596);
xnor U6123 (N_6123,N_5699,N_5284);
xnor U6124 (N_6124,N_5502,N_5555);
xnor U6125 (N_6125,N_5430,N_5295);
xnor U6126 (N_6126,N_5836,N_5589);
or U6127 (N_6127,N_5902,N_5391);
nand U6128 (N_6128,N_5668,N_5632);
xor U6129 (N_6129,N_5630,N_5565);
nor U6130 (N_6130,N_5826,N_5533);
or U6131 (N_6131,N_5660,N_5588);
nand U6132 (N_6132,N_5478,N_5908);
or U6133 (N_6133,N_5532,N_5280);
xnor U6134 (N_6134,N_5572,N_5778);
nand U6135 (N_6135,N_5407,N_5741);
and U6136 (N_6136,N_5640,N_5952);
nor U6137 (N_6137,N_5622,N_5950);
xnor U6138 (N_6138,N_5545,N_5265);
nor U6139 (N_6139,N_5290,N_5642);
and U6140 (N_6140,N_5688,N_5834);
nor U6141 (N_6141,N_5747,N_5540);
xor U6142 (N_6142,N_5601,N_5651);
and U6143 (N_6143,N_5867,N_5713);
and U6144 (N_6144,N_5672,N_5624);
nand U6145 (N_6145,N_5877,N_5480);
or U6146 (N_6146,N_5827,N_5662);
nor U6147 (N_6147,N_5780,N_5424);
xnor U6148 (N_6148,N_5554,N_5612);
nor U6149 (N_6149,N_5666,N_5796);
and U6150 (N_6150,N_5706,N_5777);
or U6151 (N_6151,N_5904,N_5977);
nand U6152 (N_6152,N_5814,N_5562);
nor U6153 (N_6153,N_5869,N_5608);
nand U6154 (N_6154,N_5566,N_5465);
and U6155 (N_6155,N_5332,N_5647);
and U6156 (N_6156,N_5874,N_5918);
and U6157 (N_6157,N_5434,N_5319);
or U6158 (N_6158,N_5402,N_5775);
and U6159 (N_6159,N_5542,N_5675);
and U6160 (N_6160,N_5963,N_5832);
nand U6161 (N_6161,N_5444,N_5525);
and U6162 (N_6162,N_5659,N_5882);
nand U6163 (N_6163,N_5382,N_5461);
or U6164 (N_6164,N_5494,N_5915);
xor U6165 (N_6165,N_5281,N_5556);
and U6166 (N_6166,N_5309,N_5781);
nand U6167 (N_6167,N_5553,N_5397);
xor U6168 (N_6168,N_5271,N_5693);
and U6169 (N_6169,N_5923,N_5275);
or U6170 (N_6170,N_5856,N_5544);
or U6171 (N_6171,N_5711,N_5998);
or U6172 (N_6172,N_5425,N_5984);
or U6173 (N_6173,N_5754,N_5452);
and U6174 (N_6174,N_5563,N_5721);
nor U6175 (N_6175,N_5852,N_5496);
and U6176 (N_6176,N_5279,N_5270);
and U6177 (N_6177,N_5650,N_5591);
and U6178 (N_6178,N_5686,N_5878);
nor U6179 (N_6179,N_5943,N_5548);
and U6180 (N_6180,N_5850,N_5416);
nor U6181 (N_6181,N_5868,N_5800);
nand U6182 (N_6182,N_5898,N_5476);
nand U6183 (N_6183,N_5724,N_5614);
or U6184 (N_6184,N_5349,N_5986);
and U6185 (N_6185,N_5681,N_5962);
nor U6186 (N_6186,N_5576,N_5661);
xor U6187 (N_6187,N_5727,N_5442);
or U6188 (N_6188,N_5671,N_5348);
xor U6189 (N_6189,N_5638,N_5860);
nand U6190 (N_6190,N_5394,N_5835);
or U6191 (N_6191,N_5837,N_5992);
and U6192 (N_6192,N_5299,N_5327);
or U6193 (N_6193,N_5453,N_5517);
nor U6194 (N_6194,N_5795,N_5855);
and U6195 (N_6195,N_5894,N_5466);
nand U6196 (N_6196,N_5305,N_5689);
nor U6197 (N_6197,N_5964,N_5859);
nor U6198 (N_6198,N_5939,N_5930);
and U6199 (N_6199,N_5657,N_5655);
or U6200 (N_6200,N_5771,N_5467);
nor U6201 (N_6201,N_5557,N_5954);
and U6202 (N_6202,N_5278,N_5579);
nand U6203 (N_6203,N_5406,N_5958);
and U6204 (N_6204,N_5273,N_5372);
or U6205 (N_6205,N_5263,N_5495);
or U6206 (N_6206,N_5643,N_5752);
nand U6207 (N_6207,N_5312,N_5742);
nand U6208 (N_6208,N_5398,N_5802);
nand U6209 (N_6209,N_5472,N_5600);
or U6210 (N_6210,N_5282,N_5790);
xor U6211 (N_6211,N_5269,N_5491);
and U6212 (N_6212,N_5314,N_5471);
and U6213 (N_6213,N_5753,N_5356);
nor U6214 (N_6214,N_5410,N_5663);
nand U6215 (N_6215,N_5611,N_5919);
nor U6216 (N_6216,N_5447,N_5395);
or U6217 (N_6217,N_5358,N_5813);
and U6218 (N_6218,N_5731,N_5401);
or U6219 (N_6219,N_5830,N_5449);
or U6220 (N_6220,N_5861,N_5695);
or U6221 (N_6221,N_5989,N_5712);
xor U6222 (N_6222,N_5357,N_5505);
and U6223 (N_6223,N_5912,N_5843);
and U6224 (N_6224,N_5423,N_5400);
or U6225 (N_6225,N_5457,N_5346);
or U6226 (N_6226,N_5255,N_5824);
or U6227 (N_6227,N_5866,N_5519);
xnor U6228 (N_6228,N_5938,N_5328);
or U6229 (N_6229,N_5947,N_5539);
and U6230 (N_6230,N_5820,N_5330);
xor U6231 (N_6231,N_5968,N_5300);
or U6232 (N_6232,N_5421,N_5887);
nand U6233 (N_6233,N_5613,N_5322);
and U6234 (N_6234,N_5973,N_5957);
nor U6235 (N_6235,N_5552,N_5736);
and U6236 (N_6236,N_5364,N_5718);
nand U6237 (N_6237,N_5260,N_5702);
xnor U6238 (N_6238,N_5808,N_5547);
or U6239 (N_6239,N_5353,N_5531);
xnor U6240 (N_6240,N_5477,N_5527);
xor U6241 (N_6241,N_5359,N_5822);
xor U6242 (N_6242,N_5411,N_5361);
nor U6243 (N_6243,N_5744,N_5374);
nor U6244 (N_6244,N_5369,N_5463);
or U6245 (N_6245,N_5339,N_5549);
nor U6246 (N_6246,N_5762,N_5770);
nor U6247 (N_6247,N_5253,N_5621);
and U6248 (N_6248,N_5735,N_5422);
nand U6249 (N_6249,N_5254,N_5536);
and U6250 (N_6250,N_5595,N_5884);
and U6251 (N_6251,N_5870,N_5685);
xnor U6252 (N_6252,N_5910,N_5750);
nand U6253 (N_6253,N_5979,N_5926);
and U6254 (N_6254,N_5629,N_5893);
nand U6255 (N_6255,N_5793,N_5259);
xnor U6256 (N_6256,N_5653,N_5670);
nor U6257 (N_6257,N_5682,N_5728);
nor U6258 (N_6258,N_5530,N_5287);
nor U6259 (N_6259,N_5844,N_5627);
and U6260 (N_6260,N_5991,N_5464);
and U6261 (N_6261,N_5507,N_5967);
xnor U6262 (N_6262,N_5316,N_5446);
or U6263 (N_6263,N_5318,N_5625);
or U6264 (N_6264,N_5804,N_5604);
xnor U6265 (N_6265,N_5865,N_5674);
and U6266 (N_6266,N_5815,N_5522);
or U6267 (N_6267,N_5597,N_5842);
or U6268 (N_6268,N_5966,N_5526);
nand U6269 (N_6269,N_5694,N_5978);
nand U6270 (N_6270,N_5782,N_5982);
nor U6271 (N_6271,N_5683,N_5787);
nor U6272 (N_6272,N_5338,N_5934);
nor U6273 (N_6273,N_5388,N_5940);
and U6274 (N_6274,N_5286,N_5283);
nor U6275 (N_6275,N_5927,N_5506);
nor U6276 (N_6276,N_5853,N_5456);
xor U6277 (N_6277,N_5308,N_5720);
and U6278 (N_6278,N_5996,N_5810);
nand U6279 (N_6279,N_5385,N_5340);
or U6280 (N_6280,N_5764,N_5906);
nand U6281 (N_6281,N_5324,N_5922);
and U6282 (N_6282,N_5304,N_5537);
and U6283 (N_6283,N_5941,N_5493);
or U6284 (N_6284,N_5725,N_5881);
xor U6285 (N_6285,N_5846,N_5717);
and U6286 (N_6286,N_5726,N_5524);
nor U6287 (N_6287,N_5704,N_5292);
nor U6288 (N_6288,N_5590,N_5475);
or U6289 (N_6289,N_5756,N_5438);
xor U6290 (N_6290,N_5876,N_5692);
nand U6291 (N_6291,N_5656,N_5691);
nor U6292 (N_6292,N_5381,N_5851);
nand U6293 (N_6293,N_5636,N_5714);
or U6294 (N_6294,N_5302,N_5337);
or U6295 (N_6295,N_5960,N_5511);
nand U6296 (N_6296,N_5776,N_5652);
and U6297 (N_6297,N_5293,N_5900);
or U6298 (N_6298,N_5432,N_5288);
and U6299 (N_6299,N_5946,N_5513);
xor U6300 (N_6300,N_5251,N_5433);
xnor U6301 (N_6301,N_5528,N_5298);
or U6302 (N_6302,N_5628,N_5838);
nor U6303 (N_6303,N_5676,N_5658);
or U6304 (N_6304,N_5785,N_5503);
nand U6305 (N_6305,N_5490,N_5366);
and U6306 (N_6306,N_5404,N_5437);
or U6307 (N_6307,N_5317,N_5633);
nor U6308 (N_6308,N_5679,N_5603);
xnor U6309 (N_6309,N_5722,N_5333);
nand U6310 (N_6310,N_5598,N_5350);
xnor U6311 (N_6311,N_5891,N_5474);
nor U6312 (N_6312,N_5587,N_5945);
or U6313 (N_6313,N_5797,N_5925);
or U6314 (N_6314,N_5313,N_5807);
or U6315 (N_6315,N_5805,N_5617);
or U6316 (N_6316,N_5276,N_5504);
or U6317 (N_6317,N_5459,N_5896);
nor U6318 (N_6318,N_5483,N_5951);
nand U6319 (N_6319,N_5436,N_5743);
and U6320 (N_6320,N_5258,N_5487);
nor U6321 (N_6321,N_5788,N_5956);
and U6322 (N_6322,N_5766,N_5615);
and U6323 (N_6323,N_5913,N_5409);
nor U6324 (N_6324,N_5510,N_5396);
or U6325 (N_6325,N_5460,N_5987);
or U6326 (N_6326,N_5811,N_5497);
nor U6327 (N_6327,N_5567,N_5551);
nand U6328 (N_6328,N_5648,N_5415);
and U6329 (N_6329,N_5574,N_5458);
and U6330 (N_6330,N_5285,N_5580);
and U6331 (N_6331,N_5509,N_5325);
and U6332 (N_6332,N_5803,N_5849);
and U6333 (N_6333,N_5734,N_5863);
and U6334 (N_6334,N_5895,N_5303);
and U6335 (N_6335,N_5564,N_5970);
and U6336 (N_6336,N_5818,N_5570);
and U6337 (N_6337,N_5921,N_5274);
xor U6338 (N_6338,N_5924,N_5335);
or U6339 (N_6339,N_5294,N_5999);
nor U6340 (N_6340,N_5888,N_5345);
nand U6341 (N_6341,N_5371,N_5994);
nor U6342 (N_6342,N_5732,N_5373);
or U6343 (N_6343,N_5383,N_5665);
nand U6344 (N_6344,N_5669,N_5903);
xor U6345 (N_6345,N_5739,N_5573);
nand U6346 (N_6346,N_5435,N_5362);
nand U6347 (N_6347,N_5678,N_5534);
and U6348 (N_6348,N_5543,N_5909);
and U6349 (N_6349,N_5839,N_5268);
and U6350 (N_6350,N_5489,N_5582);
nand U6351 (N_6351,N_5942,N_5769);
nand U6352 (N_6352,N_5626,N_5664);
xnor U6353 (N_6353,N_5840,N_5250);
nand U6354 (N_6354,N_5541,N_5583);
or U6355 (N_6355,N_5961,N_5323);
or U6356 (N_6356,N_5508,N_5774);
nor U6357 (N_6357,N_5993,N_5980);
xor U6358 (N_6358,N_5607,N_5988);
nor U6359 (N_6359,N_5705,N_5746);
nand U6360 (N_6360,N_5767,N_5729);
nand U6361 (N_6361,N_5277,N_5823);
and U6362 (N_6362,N_5707,N_5558);
nor U6363 (N_6363,N_5772,N_5687);
or U6364 (N_6364,N_5412,N_5413);
nor U6365 (N_6365,N_5759,N_5529);
nand U6366 (N_6366,N_5821,N_5405);
nand U6367 (N_6367,N_5577,N_5901);
nor U6368 (N_6368,N_5719,N_5499);
or U6369 (N_6369,N_5380,N_5990);
nand U6370 (N_6370,N_5378,N_5680);
or U6371 (N_6371,N_5758,N_5944);
and U6372 (N_6372,N_5649,N_5535);
or U6373 (N_6373,N_5684,N_5272);
nor U6374 (N_6374,N_5370,N_5252);
or U6375 (N_6375,N_5838,N_5692);
or U6376 (N_6376,N_5465,N_5865);
nand U6377 (N_6377,N_5641,N_5713);
or U6378 (N_6378,N_5763,N_5567);
nor U6379 (N_6379,N_5617,N_5887);
nor U6380 (N_6380,N_5730,N_5889);
nand U6381 (N_6381,N_5274,N_5740);
xnor U6382 (N_6382,N_5432,N_5795);
xor U6383 (N_6383,N_5794,N_5508);
nand U6384 (N_6384,N_5497,N_5458);
or U6385 (N_6385,N_5954,N_5744);
and U6386 (N_6386,N_5932,N_5969);
nor U6387 (N_6387,N_5787,N_5539);
xor U6388 (N_6388,N_5749,N_5302);
and U6389 (N_6389,N_5488,N_5780);
nor U6390 (N_6390,N_5707,N_5460);
and U6391 (N_6391,N_5456,N_5691);
or U6392 (N_6392,N_5964,N_5868);
and U6393 (N_6393,N_5452,N_5753);
or U6394 (N_6394,N_5900,N_5756);
and U6395 (N_6395,N_5421,N_5904);
nand U6396 (N_6396,N_5946,N_5972);
or U6397 (N_6397,N_5972,N_5979);
or U6398 (N_6398,N_5621,N_5269);
or U6399 (N_6399,N_5916,N_5458);
and U6400 (N_6400,N_5743,N_5663);
nor U6401 (N_6401,N_5286,N_5496);
xnor U6402 (N_6402,N_5622,N_5270);
nand U6403 (N_6403,N_5483,N_5360);
nor U6404 (N_6404,N_5257,N_5269);
and U6405 (N_6405,N_5311,N_5270);
nand U6406 (N_6406,N_5948,N_5968);
and U6407 (N_6407,N_5826,N_5456);
nand U6408 (N_6408,N_5820,N_5988);
xor U6409 (N_6409,N_5621,N_5915);
nand U6410 (N_6410,N_5889,N_5990);
nand U6411 (N_6411,N_5404,N_5624);
or U6412 (N_6412,N_5780,N_5458);
nor U6413 (N_6413,N_5880,N_5778);
nor U6414 (N_6414,N_5266,N_5255);
nor U6415 (N_6415,N_5873,N_5500);
and U6416 (N_6416,N_5798,N_5554);
nor U6417 (N_6417,N_5294,N_5319);
and U6418 (N_6418,N_5937,N_5454);
xor U6419 (N_6419,N_5796,N_5380);
xor U6420 (N_6420,N_5345,N_5904);
nand U6421 (N_6421,N_5973,N_5738);
or U6422 (N_6422,N_5771,N_5557);
or U6423 (N_6423,N_5254,N_5912);
nor U6424 (N_6424,N_5444,N_5710);
nor U6425 (N_6425,N_5627,N_5952);
nor U6426 (N_6426,N_5263,N_5578);
nor U6427 (N_6427,N_5782,N_5446);
nand U6428 (N_6428,N_5288,N_5905);
and U6429 (N_6429,N_5389,N_5269);
nor U6430 (N_6430,N_5383,N_5644);
nor U6431 (N_6431,N_5377,N_5267);
nor U6432 (N_6432,N_5530,N_5388);
xnor U6433 (N_6433,N_5795,N_5564);
nor U6434 (N_6434,N_5382,N_5433);
nand U6435 (N_6435,N_5909,N_5755);
and U6436 (N_6436,N_5741,N_5892);
and U6437 (N_6437,N_5315,N_5549);
or U6438 (N_6438,N_5446,N_5920);
xor U6439 (N_6439,N_5933,N_5408);
nand U6440 (N_6440,N_5788,N_5388);
or U6441 (N_6441,N_5426,N_5953);
nand U6442 (N_6442,N_5970,N_5252);
nor U6443 (N_6443,N_5592,N_5500);
and U6444 (N_6444,N_5970,N_5438);
nand U6445 (N_6445,N_5965,N_5743);
or U6446 (N_6446,N_5830,N_5321);
nor U6447 (N_6447,N_5942,N_5777);
or U6448 (N_6448,N_5373,N_5698);
nand U6449 (N_6449,N_5468,N_5403);
or U6450 (N_6450,N_5659,N_5349);
nand U6451 (N_6451,N_5784,N_5296);
nor U6452 (N_6452,N_5730,N_5332);
and U6453 (N_6453,N_5476,N_5866);
nor U6454 (N_6454,N_5928,N_5582);
nor U6455 (N_6455,N_5483,N_5603);
or U6456 (N_6456,N_5255,N_5443);
and U6457 (N_6457,N_5308,N_5566);
nor U6458 (N_6458,N_5636,N_5902);
xor U6459 (N_6459,N_5416,N_5350);
nand U6460 (N_6460,N_5454,N_5346);
or U6461 (N_6461,N_5511,N_5576);
or U6462 (N_6462,N_5931,N_5715);
nor U6463 (N_6463,N_5949,N_5603);
nor U6464 (N_6464,N_5635,N_5601);
nor U6465 (N_6465,N_5462,N_5628);
or U6466 (N_6466,N_5733,N_5707);
nand U6467 (N_6467,N_5989,N_5835);
nand U6468 (N_6468,N_5529,N_5802);
nor U6469 (N_6469,N_5678,N_5469);
nand U6470 (N_6470,N_5303,N_5798);
and U6471 (N_6471,N_5495,N_5698);
nor U6472 (N_6472,N_5556,N_5967);
and U6473 (N_6473,N_5361,N_5712);
nor U6474 (N_6474,N_5941,N_5968);
nand U6475 (N_6475,N_5834,N_5331);
nand U6476 (N_6476,N_5673,N_5541);
xor U6477 (N_6477,N_5774,N_5985);
nor U6478 (N_6478,N_5912,N_5520);
and U6479 (N_6479,N_5557,N_5742);
nor U6480 (N_6480,N_5383,N_5351);
or U6481 (N_6481,N_5467,N_5623);
or U6482 (N_6482,N_5904,N_5535);
nand U6483 (N_6483,N_5910,N_5287);
nor U6484 (N_6484,N_5622,N_5684);
or U6485 (N_6485,N_5911,N_5260);
or U6486 (N_6486,N_5513,N_5250);
nand U6487 (N_6487,N_5885,N_5464);
nand U6488 (N_6488,N_5477,N_5492);
nand U6489 (N_6489,N_5836,N_5609);
and U6490 (N_6490,N_5553,N_5369);
or U6491 (N_6491,N_5361,N_5757);
nand U6492 (N_6492,N_5873,N_5994);
and U6493 (N_6493,N_5894,N_5457);
nand U6494 (N_6494,N_5837,N_5500);
nor U6495 (N_6495,N_5603,N_5473);
nand U6496 (N_6496,N_5741,N_5624);
xor U6497 (N_6497,N_5490,N_5781);
nand U6498 (N_6498,N_5964,N_5735);
nor U6499 (N_6499,N_5587,N_5492);
and U6500 (N_6500,N_5862,N_5551);
and U6501 (N_6501,N_5840,N_5841);
nor U6502 (N_6502,N_5963,N_5321);
and U6503 (N_6503,N_5950,N_5660);
nand U6504 (N_6504,N_5824,N_5906);
nand U6505 (N_6505,N_5626,N_5547);
and U6506 (N_6506,N_5460,N_5979);
or U6507 (N_6507,N_5941,N_5272);
nor U6508 (N_6508,N_5532,N_5984);
or U6509 (N_6509,N_5595,N_5755);
and U6510 (N_6510,N_5398,N_5783);
nand U6511 (N_6511,N_5799,N_5497);
nand U6512 (N_6512,N_5302,N_5297);
and U6513 (N_6513,N_5924,N_5568);
nand U6514 (N_6514,N_5811,N_5726);
nor U6515 (N_6515,N_5277,N_5397);
nor U6516 (N_6516,N_5865,N_5580);
or U6517 (N_6517,N_5900,N_5263);
and U6518 (N_6518,N_5390,N_5725);
or U6519 (N_6519,N_5622,N_5590);
nand U6520 (N_6520,N_5435,N_5853);
nor U6521 (N_6521,N_5827,N_5493);
nor U6522 (N_6522,N_5783,N_5770);
or U6523 (N_6523,N_5625,N_5513);
or U6524 (N_6524,N_5440,N_5723);
and U6525 (N_6525,N_5881,N_5877);
xnor U6526 (N_6526,N_5818,N_5654);
nand U6527 (N_6527,N_5910,N_5605);
xnor U6528 (N_6528,N_5359,N_5946);
or U6529 (N_6529,N_5564,N_5635);
nor U6530 (N_6530,N_5506,N_5352);
and U6531 (N_6531,N_5446,N_5674);
nor U6532 (N_6532,N_5819,N_5545);
nand U6533 (N_6533,N_5370,N_5539);
nor U6534 (N_6534,N_5386,N_5484);
xnor U6535 (N_6535,N_5340,N_5618);
nand U6536 (N_6536,N_5579,N_5858);
or U6537 (N_6537,N_5797,N_5837);
nand U6538 (N_6538,N_5274,N_5850);
or U6539 (N_6539,N_5965,N_5528);
nand U6540 (N_6540,N_5545,N_5397);
nand U6541 (N_6541,N_5377,N_5358);
or U6542 (N_6542,N_5260,N_5721);
and U6543 (N_6543,N_5840,N_5275);
or U6544 (N_6544,N_5960,N_5497);
or U6545 (N_6545,N_5979,N_5302);
xor U6546 (N_6546,N_5380,N_5964);
nand U6547 (N_6547,N_5682,N_5911);
nand U6548 (N_6548,N_5851,N_5790);
and U6549 (N_6549,N_5444,N_5978);
nor U6550 (N_6550,N_5480,N_5471);
xor U6551 (N_6551,N_5541,N_5646);
nand U6552 (N_6552,N_5799,N_5547);
or U6553 (N_6553,N_5463,N_5922);
and U6554 (N_6554,N_5668,N_5895);
nand U6555 (N_6555,N_5729,N_5608);
and U6556 (N_6556,N_5530,N_5948);
nor U6557 (N_6557,N_5755,N_5571);
nand U6558 (N_6558,N_5398,N_5934);
and U6559 (N_6559,N_5901,N_5415);
nor U6560 (N_6560,N_5813,N_5885);
or U6561 (N_6561,N_5421,N_5579);
and U6562 (N_6562,N_5934,N_5769);
nor U6563 (N_6563,N_5271,N_5817);
xor U6564 (N_6564,N_5291,N_5763);
nor U6565 (N_6565,N_5394,N_5302);
nor U6566 (N_6566,N_5640,N_5975);
nor U6567 (N_6567,N_5938,N_5340);
and U6568 (N_6568,N_5945,N_5667);
or U6569 (N_6569,N_5743,N_5929);
or U6570 (N_6570,N_5421,N_5271);
or U6571 (N_6571,N_5411,N_5286);
nor U6572 (N_6572,N_5514,N_5870);
and U6573 (N_6573,N_5703,N_5474);
xnor U6574 (N_6574,N_5765,N_5646);
and U6575 (N_6575,N_5660,N_5646);
nand U6576 (N_6576,N_5590,N_5383);
or U6577 (N_6577,N_5624,N_5516);
nor U6578 (N_6578,N_5449,N_5868);
nor U6579 (N_6579,N_5698,N_5294);
nand U6580 (N_6580,N_5837,N_5627);
nor U6581 (N_6581,N_5566,N_5632);
and U6582 (N_6582,N_5860,N_5777);
nand U6583 (N_6583,N_5814,N_5308);
nand U6584 (N_6584,N_5554,N_5889);
or U6585 (N_6585,N_5702,N_5745);
nand U6586 (N_6586,N_5476,N_5985);
nand U6587 (N_6587,N_5581,N_5758);
and U6588 (N_6588,N_5411,N_5846);
and U6589 (N_6589,N_5452,N_5695);
and U6590 (N_6590,N_5745,N_5936);
and U6591 (N_6591,N_5785,N_5574);
or U6592 (N_6592,N_5635,N_5922);
nor U6593 (N_6593,N_5934,N_5929);
and U6594 (N_6594,N_5586,N_5327);
and U6595 (N_6595,N_5724,N_5627);
or U6596 (N_6596,N_5837,N_5319);
nor U6597 (N_6597,N_5940,N_5697);
nand U6598 (N_6598,N_5838,N_5820);
nor U6599 (N_6599,N_5398,N_5699);
xnor U6600 (N_6600,N_5952,N_5810);
and U6601 (N_6601,N_5308,N_5586);
or U6602 (N_6602,N_5872,N_5268);
nand U6603 (N_6603,N_5496,N_5719);
and U6604 (N_6604,N_5863,N_5569);
nor U6605 (N_6605,N_5259,N_5335);
nor U6606 (N_6606,N_5431,N_5912);
or U6607 (N_6607,N_5524,N_5353);
and U6608 (N_6608,N_5925,N_5736);
and U6609 (N_6609,N_5473,N_5605);
nor U6610 (N_6610,N_5445,N_5652);
and U6611 (N_6611,N_5605,N_5443);
xor U6612 (N_6612,N_5887,N_5290);
nor U6613 (N_6613,N_5324,N_5857);
or U6614 (N_6614,N_5375,N_5589);
or U6615 (N_6615,N_5269,N_5321);
nor U6616 (N_6616,N_5746,N_5480);
nor U6617 (N_6617,N_5724,N_5929);
nand U6618 (N_6618,N_5307,N_5464);
or U6619 (N_6619,N_5302,N_5456);
or U6620 (N_6620,N_5720,N_5852);
or U6621 (N_6621,N_5977,N_5941);
nor U6622 (N_6622,N_5818,N_5431);
nand U6623 (N_6623,N_5401,N_5504);
nor U6624 (N_6624,N_5989,N_5713);
nand U6625 (N_6625,N_5658,N_5813);
and U6626 (N_6626,N_5637,N_5867);
nand U6627 (N_6627,N_5267,N_5622);
nand U6628 (N_6628,N_5284,N_5499);
nand U6629 (N_6629,N_5780,N_5502);
nand U6630 (N_6630,N_5531,N_5869);
or U6631 (N_6631,N_5990,N_5693);
or U6632 (N_6632,N_5839,N_5983);
nand U6633 (N_6633,N_5997,N_5998);
or U6634 (N_6634,N_5728,N_5408);
nor U6635 (N_6635,N_5850,N_5308);
and U6636 (N_6636,N_5781,N_5704);
and U6637 (N_6637,N_5999,N_5742);
and U6638 (N_6638,N_5964,N_5582);
nand U6639 (N_6639,N_5569,N_5698);
nand U6640 (N_6640,N_5976,N_5517);
nor U6641 (N_6641,N_5779,N_5837);
or U6642 (N_6642,N_5688,N_5721);
or U6643 (N_6643,N_5838,N_5695);
nand U6644 (N_6644,N_5420,N_5352);
and U6645 (N_6645,N_5450,N_5974);
or U6646 (N_6646,N_5713,N_5547);
nor U6647 (N_6647,N_5761,N_5751);
nor U6648 (N_6648,N_5427,N_5870);
or U6649 (N_6649,N_5298,N_5836);
or U6650 (N_6650,N_5440,N_5919);
and U6651 (N_6651,N_5757,N_5843);
nand U6652 (N_6652,N_5894,N_5677);
and U6653 (N_6653,N_5680,N_5892);
nand U6654 (N_6654,N_5683,N_5437);
xor U6655 (N_6655,N_5807,N_5909);
nor U6656 (N_6656,N_5914,N_5745);
or U6657 (N_6657,N_5266,N_5555);
nor U6658 (N_6658,N_5531,N_5737);
nand U6659 (N_6659,N_5638,N_5331);
and U6660 (N_6660,N_5279,N_5331);
nor U6661 (N_6661,N_5537,N_5262);
and U6662 (N_6662,N_5660,N_5527);
nor U6663 (N_6663,N_5769,N_5576);
xnor U6664 (N_6664,N_5619,N_5862);
or U6665 (N_6665,N_5999,N_5289);
nor U6666 (N_6666,N_5341,N_5257);
and U6667 (N_6667,N_5657,N_5379);
nand U6668 (N_6668,N_5369,N_5921);
nand U6669 (N_6669,N_5502,N_5611);
nor U6670 (N_6670,N_5429,N_5412);
or U6671 (N_6671,N_5937,N_5887);
xnor U6672 (N_6672,N_5704,N_5919);
and U6673 (N_6673,N_5429,N_5669);
nand U6674 (N_6674,N_5283,N_5884);
and U6675 (N_6675,N_5369,N_5441);
and U6676 (N_6676,N_5776,N_5475);
nand U6677 (N_6677,N_5419,N_5862);
and U6678 (N_6678,N_5483,N_5547);
nor U6679 (N_6679,N_5822,N_5801);
and U6680 (N_6680,N_5644,N_5697);
nor U6681 (N_6681,N_5541,N_5692);
or U6682 (N_6682,N_5435,N_5789);
nand U6683 (N_6683,N_5784,N_5678);
and U6684 (N_6684,N_5386,N_5876);
xnor U6685 (N_6685,N_5920,N_5583);
nor U6686 (N_6686,N_5441,N_5931);
nor U6687 (N_6687,N_5629,N_5977);
or U6688 (N_6688,N_5910,N_5930);
xor U6689 (N_6689,N_5945,N_5349);
nand U6690 (N_6690,N_5501,N_5287);
and U6691 (N_6691,N_5515,N_5428);
and U6692 (N_6692,N_5294,N_5290);
or U6693 (N_6693,N_5267,N_5844);
and U6694 (N_6694,N_5676,N_5388);
and U6695 (N_6695,N_5853,N_5632);
or U6696 (N_6696,N_5280,N_5679);
nand U6697 (N_6697,N_5376,N_5624);
or U6698 (N_6698,N_5587,N_5453);
or U6699 (N_6699,N_5824,N_5340);
and U6700 (N_6700,N_5853,N_5617);
nand U6701 (N_6701,N_5958,N_5630);
nor U6702 (N_6702,N_5388,N_5760);
and U6703 (N_6703,N_5439,N_5351);
xor U6704 (N_6704,N_5952,N_5730);
and U6705 (N_6705,N_5746,N_5355);
or U6706 (N_6706,N_5948,N_5442);
xnor U6707 (N_6707,N_5392,N_5751);
nor U6708 (N_6708,N_5517,N_5731);
nand U6709 (N_6709,N_5789,N_5921);
or U6710 (N_6710,N_5917,N_5589);
or U6711 (N_6711,N_5922,N_5548);
or U6712 (N_6712,N_5511,N_5983);
or U6713 (N_6713,N_5735,N_5763);
or U6714 (N_6714,N_5785,N_5611);
nor U6715 (N_6715,N_5577,N_5338);
xor U6716 (N_6716,N_5821,N_5937);
nor U6717 (N_6717,N_5839,N_5321);
and U6718 (N_6718,N_5536,N_5545);
nand U6719 (N_6719,N_5727,N_5257);
nand U6720 (N_6720,N_5637,N_5821);
or U6721 (N_6721,N_5974,N_5401);
xor U6722 (N_6722,N_5466,N_5993);
nand U6723 (N_6723,N_5775,N_5561);
xnor U6724 (N_6724,N_5774,N_5341);
nor U6725 (N_6725,N_5403,N_5593);
and U6726 (N_6726,N_5455,N_5592);
nor U6727 (N_6727,N_5607,N_5606);
nor U6728 (N_6728,N_5561,N_5487);
or U6729 (N_6729,N_5694,N_5426);
and U6730 (N_6730,N_5887,N_5363);
xnor U6731 (N_6731,N_5916,N_5390);
and U6732 (N_6732,N_5612,N_5800);
xor U6733 (N_6733,N_5260,N_5510);
xor U6734 (N_6734,N_5644,N_5787);
nor U6735 (N_6735,N_5941,N_5794);
nand U6736 (N_6736,N_5458,N_5599);
and U6737 (N_6737,N_5474,N_5873);
xnor U6738 (N_6738,N_5726,N_5934);
nor U6739 (N_6739,N_5877,N_5535);
or U6740 (N_6740,N_5323,N_5336);
nor U6741 (N_6741,N_5410,N_5801);
nand U6742 (N_6742,N_5983,N_5798);
or U6743 (N_6743,N_5759,N_5293);
and U6744 (N_6744,N_5307,N_5347);
nand U6745 (N_6745,N_5510,N_5990);
and U6746 (N_6746,N_5466,N_5311);
and U6747 (N_6747,N_5870,N_5948);
nand U6748 (N_6748,N_5280,N_5987);
and U6749 (N_6749,N_5284,N_5604);
nor U6750 (N_6750,N_6071,N_6533);
nor U6751 (N_6751,N_6381,N_6484);
nor U6752 (N_6752,N_6293,N_6523);
and U6753 (N_6753,N_6371,N_6699);
nor U6754 (N_6754,N_6445,N_6069);
nor U6755 (N_6755,N_6472,N_6491);
and U6756 (N_6756,N_6573,N_6019);
nand U6757 (N_6757,N_6142,N_6626);
nand U6758 (N_6758,N_6229,N_6539);
nor U6759 (N_6759,N_6544,N_6553);
nor U6760 (N_6760,N_6543,N_6407);
or U6761 (N_6761,N_6174,N_6106);
nand U6762 (N_6762,N_6119,N_6058);
nor U6763 (N_6763,N_6661,N_6046);
and U6764 (N_6764,N_6546,N_6648);
nand U6765 (N_6765,N_6285,N_6576);
nor U6766 (N_6766,N_6329,N_6040);
and U6767 (N_6767,N_6207,N_6726);
xnor U6768 (N_6768,N_6324,N_6365);
nor U6769 (N_6769,N_6487,N_6683);
and U6770 (N_6770,N_6203,N_6141);
nand U6771 (N_6771,N_6720,N_6340);
and U6772 (N_6772,N_6298,N_6688);
nand U6773 (N_6773,N_6509,N_6149);
or U6774 (N_6774,N_6101,N_6458);
or U6775 (N_6775,N_6137,N_6330);
nor U6776 (N_6776,N_6043,N_6538);
xor U6777 (N_6777,N_6386,N_6346);
nand U6778 (N_6778,N_6166,N_6712);
or U6779 (N_6779,N_6332,N_6112);
xnor U6780 (N_6780,N_6701,N_6182);
nand U6781 (N_6781,N_6746,N_6524);
nor U6782 (N_6782,N_6702,N_6376);
nand U6783 (N_6783,N_6256,N_6646);
or U6784 (N_6784,N_6429,N_6385);
and U6785 (N_6785,N_6505,N_6372);
or U6786 (N_6786,N_6603,N_6246);
or U6787 (N_6787,N_6640,N_6263);
and U6788 (N_6788,N_6569,N_6557);
and U6789 (N_6789,N_6123,N_6579);
and U6790 (N_6790,N_6219,N_6074);
xor U6791 (N_6791,N_6225,N_6389);
nor U6792 (N_6792,N_6098,N_6453);
nor U6793 (N_6793,N_6247,N_6086);
xnor U6794 (N_6794,N_6451,N_6190);
or U6795 (N_6795,N_6259,N_6710);
nand U6796 (N_6796,N_6162,N_6618);
nand U6797 (N_6797,N_6047,N_6695);
and U6798 (N_6798,N_6282,N_6159);
xor U6799 (N_6799,N_6657,N_6287);
xnor U6800 (N_6800,N_6614,N_6067);
xor U6801 (N_6801,N_6335,N_6305);
and U6802 (N_6802,N_6144,N_6191);
nor U6803 (N_6803,N_6439,N_6474);
and U6804 (N_6804,N_6696,N_6420);
xor U6805 (N_6805,N_6239,N_6303);
and U6806 (N_6806,N_6029,N_6313);
and U6807 (N_6807,N_6664,N_6322);
xnor U6808 (N_6808,N_6627,N_6541);
or U6809 (N_6809,N_6093,N_6555);
nor U6810 (N_6810,N_6638,N_6438);
or U6811 (N_6811,N_6440,N_6268);
nor U6812 (N_6812,N_6321,N_6405);
and U6813 (N_6813,N_6584,N_6483);
or U6814 (N_6814,N_6673,N_6168);
and U6815 (N_6815,N_6201,N_6022);
nor U6816 (N_6816,N_6070,N_6411);
xor U6817 (N_6817,N_6030,N_6350);
nand U6818 (N_6818,N_6110,N_6104);
and U6819 (N_6819,N_6631,N_6749);
and U6820 (N_6820,N_6449,N_6547);
nand U6821 (N_6821,N_6124,N_6412);
or U6822 (N_6822,N_6488,N_6248);
and U6823 (N_6823,N_6577,N_6408);
or U6824 (N_6824,N_6575,N_6489);
nand U6825 (N_6825,N_6624,N_6619);
nor U6826 (N_6826,N_6645,N_6473);
and U6827 (N_6827,N_6187,N_6223);
or U6828 (N_6828,N_6361,N_6276);
and U6829 (N_6829,N_6588,N_6196);
xor U6830 (N_6830,N_6060,N_6525);
nor U6831 (N_6831,N_6306,N_6002);
and U6832 (N_6832,N_6426,N_6333);
and U6833 (N_6833,N_6369,N_6520);
or U6834 (N_6834,N_6529,N_6602);
or U6835 (N_6835,N_6561,N_6336);
and U6836 (N_6836,N_6609,N_6629);
and U6837 (N_6837,N_6200,N_6568);
nor U6838 (N_6838,N_6367,N_6265);
nor U6839 (N_6839,N_6507,N_6585);
and U6840 (N_6840,N_6097,N_6692);
nand U6841 (N_6841,N_6658,N_6084);
and U6842 (N_6842,N_6033,N_6051);
nor U6843 (N_6843,N_6202,N_6642);
nand U6844 (N_6844,N_6279,N_6226);
xor U6845 (N_6845,N_6528,N_6500);
nor U6846 (N_6846,N_6522,N_6028);
nor U6847 (N_6847,N_6551,N_6402);
xor U6848 (N_6848,N_6393,N_6460);
nor U6849 (N_6849,N_6558,N_6072);
nand U6850 (N_6850,N_6077,N_6493);
or U6851 (N_6851,N_6610,N_6406);
and U6852 (N_6852,N_6003,N_6537);
xnor U6853 (N_6853,N_6267,N_6742);
nor U6854 (N_6854,N_6671,N_6020);
nor U6855 (N_6855,N_6281,N_6660);
nor U6856 (N_6856,N_6452,N_6274);
xnor U6857 (N_6857,N_6620,N_6700);
nor U6858 (N_6858,N_6179,N_6722);
nor U6859 (N_6859,N_6125,N_6231);
xnor U6860 (N_6860,N_6652,N_6153);
nor U6861 (N_6861,N_6514,N_6630);
and U6862 (N_6862,N_6266,N_6542);
or U6863 (N_6863,N_6680,N_6616);
and U6864 (N_6864,N_6192,N_6503);
nor U6865 (N_6865,N_6235,N_6118);
nor U6866 (N_6866,N_6230,N_6552);
nand U6867 (N_6867,N_6001,N_6146);
nand U6868 (N_6868,N_6475,N_6283);
nand U6869 (N_6869,N_6165,N_6158);
nand U6870 (N_6870,N_6581,N_6601);
or U6871 (N_6871,N_6253,N_6087);
nand U6872 (N_6872,N_6075,N_6327);
or U6873 (N_6873,N_6092,N_6476);
nand U6874 (N_6874,N_6669,N_6150);
and U6875 (N_6875,N_6733,N_6422);
and U6876 (N_6876,N_6743,N_6740);
nand U6877 (N_6877,N_6210,N_6467);
or U6878 (N_6878,N_6387,N_6309);
and U6879 (N_6879,N_6338,N_6513);
or U6880 (N_6880,N_6024,N_6341);
nand U6881 (N_6881,N_6056,N_6025);
or U6882 (N_6882,N_6587,N_6310);
or U6883 (N_6883,N_6594,N_6213);
nand U6884 (N_6884,N_6470,N_6674);
nand U6885 (N_6885,N_6425,N_6010);
nand U6886 (N_6886,N_6015,N_6085);
or U6887 (N_6887,N_6462,N_6723);
xnor U6888 (N_6888,N_6506,N_6578);
nand U6889 (N_6889,N_6744,N_6731);
and U6890 (N_6890,N_6271,N_6250);
or U6891 (N_6891,N_6478,N_6184);
nor U6892 (N_6892,N_6531,N_6394);
xnor U6893 (N_6893,N_6611,N_6741);
nor U6894 (N_6894,N_6049,N_6454);
nand U6895 (N_6895,N_6607,N_6252);
and U6896 (N_6896,N_6353,N_6319);
and U6897 (N_6897,N_6549,N_6679);
nor U6898 (N_6898,N_6510,N_6604);
nand U6899 (N_6899,N_6628,N_6502);
nor U6900 (N_6900,N_6380,N_6666);
nand U6901 (N_6901,N_6277,N_6126);
xor U6902 (N_6902,N_6388,N_6048);
or U6903 (N_6903,N_6042,N_6721);
nor U6904 (N_6904,N_6649,N_6532);
and U6905 (N_6905,N_6308,N_6677);
and U6906 (N_6906,N_6099,N_6635);
nor U6907 (N_6907,N_6090,N_6466);
and U6908 (N_6908,N_6227,N_6291);
nor U6909 (N_6909,N_6436,N_6176);
xnor U6910 (N_6910,N_6006,N_6540);
or U6911 (N_6911,N_6157,N_6495);
nor U6912 (N_6912,N_6115,N_6299);
or U6913 (N_6913,N_6288,N_6297);
nand U6914 (N_6914,N_6732,N_6665);
xnor U6915 (N_6915,N_6189,N_6073);
xnor U6916 (N_6916,N_6181,N_6081);
and U6917 (N_6917,N_6136,N_6691);
nand U6918 (N_6918,N_6398,N_6325);
or U6919 (N_6919,N_6185,N_6005);
nand U6920 (N_6920,N_6416,N_6356);
nand U6921 (N_6921,N_6378,N_6254);
nand U6922 (N_6922,N_6143,N_6521);
or U6923 (N_6923,N_6217,N_6622);
nor U6924 (N_6924,N_6140,N_6441);
xor U6925 (N_6925,N_6014,N_6486);
nor U6926 (N_6926,N_6280,N_6261);
and U6927 (N_6927,N_6262,N_6345);
and U6928 (N_6928,N_6401,N_6197);
and U6929 (N_6929,N_6206,N_6608);
xnor U6930 (N_6930,N_6471,N_6709);
and U6931 (N_6931,N_6214,N_6082);
and U6932 (N_6932,N_6396,N_6275);
nor U6933 (N_6933,N_6103,N_6148);
or U6934 (N_6934,N_6719,N_6032);
or U6935 (N_6935,N_6698,N_6636);
or U6936 (N_6936,N_6632,N_6655);
nand U6937 (N_6937,N_6164,N_6316);
nand U6938 (N_6938,N_6560,N_6373);
or U6939 (N_6939,N_6013,N_6504);
and U6940 (N_6940,N_6132,N_6572);
and U6941 (N_6941,N_6102,N_6328);
or U6942 (N_6942,N_6044,N_6461);
nor U6943 (N_6943,N_6704,N_6116);
or U6944 (N_6944,N_6562,N_6747);
or U6945 (N_6945,N_6120,N_6053);
and U6946 (N_6946,N_6595,N_6108);
or U6947 (N_6947,N_6526,N_6034);
nor U6948 (N_6948,N_6129,N_6432);
nand U6949 (N_6949,N_6039,N_6130);
nand U6950 (N_6950,N_6375,N_6138);
nor U6951 (N_6951,N_6667,N_6270);
and U6952 (N_6952,N_6447,N_6516);
and U6953 (N_6953,N_6748,N_6415);
nand U6954 (N_6954,N_6403,N_6334);
nand U6955 (N_6955,N_6662,N_6243);
nor U6956 (N_6956,N_6545,N_6041);
nand U6957 (N_6957,N_6357,N_6427);
nor U6958 (N_6958,N_6131,N_6519);
nand U6959 (N_6959,N_6613,N_6697);
nor U6960 (N_6960,N_6715,N_6347);
and U6961 (N_6961,N_6559,N_6301);
and U6962 (N_6962,N_6094,N_6713);
nand U6963 (N_6963,N_6343,N_6314);
nand U6964 (N_6964,N_6482,N_6417);
and U6965 (N_6965,N_6269,N_6349);
and U6966 (N_6966,N_6065,N_6292);
and U6967 (N_6967,N_6566,N_6121);
xnor U6968 (N_6968,N_6433,N_6724);
nand U6969 (N_6969,N_6175,N_6255);
or U6970 (N_6970,N_6621,N_6320);
and U6971 (N_6971,N_6021,N_6377);
and U6972 (N_6972,N_6161,N_6366);
or U6973 (N_6973,N_6606,N_6016);
and U6974 (N_6974,N_6193,N_6567);
or U6975 (N_6975,N_6479,N_6413);
nor U6976 (N_6976,N_6171,N_6705);
nor U6977 (N_6977,N_6435,N_6331);
or U6978 (N_6978,N_6038,N_6342);
nand U6979 (N_6979,N_6586,N_6233);
nor U6980 (N_6980,N_6362,N_6195);
and U6981 (N_6981,N_6012,N_6681);
or U6982 (N_6982,N_6026,N_6729);
and U6983 (N_6983,N_6515,N_6163);
nor U6984 (N_6984,N_6391,N_6249);
or U6985 (N_6985,N_6736,N_6107);
nand U6986 (N_6986,N_6392,N_6465);
and U6987 (N_6987,N_6668,N_6000);
xnor U6988 (N_6988,N_6169,N_6672);
xor U6989 (N_6989,N_6273,N_6083);
nand U6990 (N_6990,N_6605,N_6374);
nor U6991 (N_6991,N_6221,N_6311);
nand U6992 (N_6992,N_6512,N_6199);
and U6993 (N_6993,N_6463,N_6264);
and U6994 (N_6994,N_6404,N_6198);
or U6995 (N_6995,N_6068,N_6091);
nand U6996 (N_6996,N_6527,N_6469);
and U6997 (N_6997,N_6205,N_6570);
and U6998 (N_6998,N_6556,N_6257);
or U6999 (N_6999,N_6428,N_6080);
and U7000 (N_7000,N_6355,N_6204);
nor U7001 (N_7001,N_6592,N_6004);
and U7002 (N_7002,N_6591,N_6617);
xor U7003 (N_7003,N_6061,N_6653);
or U7004 (N_7004,N_6589,N_6490);
or U7005 (N_7005,N_6368,N_6414);
nand U7006 (N_7006,N_6656,N_6088);
and U7007 (N_7007,N_6258,N_6236);
or U7008 (N_7008,N_6064,N_6364);
nand U7009 (N_7009,N_6127,N_6634);
nand U7010 (N_7010,N_6154,N_6639);
nand U7011 (N_7011,N_6468,N_6155);
nand U7012 (N_7012,N_6718,N_6734);
or U7013 (N_7013,N_6456,N_6326);
nor U7014 (N_7014,N_6352,N_6260);
nand U7015 (N_7015,N_6497,N_6222);
nand U7016 (N_7016,N_6009,N_6745);
and U7017 (N_7017,N_6173,N_6105);
and U7018 (N_7018,N_6582,N_6739);
or U7019 (N_7019,N_6641,N_6430);
nor U7020 (N_7020,N_6443,N_6054);
xor U7021 (N_7021,N_6272,N_6459);
nor U7022 (N_7022,N_6384,N_6714);
and U7023 (N_7023,N_6237,N_6152);
nor U7024 (N_7024,N_6348,N_6464);
and U7025 (N_7025,N_6687,N_6289);
nand U7026 (N_7026,N_6117,N_6096);
xor U7027 (N_7027,N_6597,N_6596);
or U7028 (N_7028,N_6593,N_6290);
xnor U7029 (N_7029,N_6481,N_6686);
nor U7030 (N_7030,N_6062,N_6725);
nor U7031 (N_7031,N_6409,N_6703);
nand U7032 (N_7032,N_6172,N_6300);
and U7033 (N_7033,N_6114,N_6534);
nand U7034 (N_7034,N_6654,N_6218);
nand U7035 (N_7035,N_6706,N_6499);
nand U7036 (N_7036,N_6302,N_6111);
xor U7037 (N_7037,N_6563,N_6359);
and U7038 (N_7038,N_6045,N_6612);
nand U7039 (N_7039,N_6344,N_6518);
and U7040 (N_7040,N_6007,N_6650);
or U7041 (N_7041,N_6211,N_6216);
or U7042 (N_7042,N_6018,N_6063);
or U7043 (N_7043,N_6598,N_6390);
nand U7044 (N_7044,N_6496,N_6244);
or U7045 (N_7045,N_6676,N_6424);
or U7046 (N_7046,N_6057,N_6337);
or U7047 (N_7047,N_6682,N_6180);
or U7048 (N_7048,N_6564,N_6550);
xor U7049 (N_7049,N_6444,N_6078);
and U7050 (N_7050,N_6437,N_6183);
and U7051 (N_7051,N_6050,N_6615);
or U7052 (N_7052,N_6383,N_6304);
and U7053 (N_7053,N_6147,N_6188);
or U7054 (N_7054,N_6177,N_6419);
nand U7055 (N_7055,N_6625,N_6633);
xnor U7056 (N_7056,N_6663,N_6224);
nand U7057 (N_7057,N_6446,N_6295);
nor U7058 (N_7058,N_6738,N_6241);
nor U7059 (N_7059,N_6590,N_6643);
and U7060 (N_7060,N_6678,N_6315);
nand U7061 (N_7061,N_6448,N_6035);
and U7062 (N_7062,N_6599,N_6511);
nor U7063 (N_7063,N_6023,N_6535);
or U7064 (N_7064,N_6240,N_6194);
or U7065 (N_7065,N_6135,N_6251);
and U7066 (N_7066,N_6220,N_6059);
nand U7067 (N_7067,N_6457,N_6717);
xnor U7068 (N_7068,N_6637,N_6727);
and U7069 (N_7069,N_6017,N_6477);
xor U7070 (N_7070,N_6670,N_6156);
or U7071 (N_7071,N_6530,N_6685);
and U7072 (N_7072,N_6455,N_6730);
nand U7073 (N_7073,N_6410,N_6134);
or U7074 (N_7074,N_6339,N_6675);
nor U7075 (N_7075,N_6128,N_6382);
or U7076 (N_7076,N_6351,N_6238);
nand U7077 (N_7077,N_6690,N_6354);
and U7078 (N_7078,N_6418,N_6312);
or U7079 (N_7079,N_6360,N_6508);
xnor U7080 (N_7080,N_6728,N_6571);
and U7081 (N_7081,N_6066,N_6716);
nand U7082 (N_7082,N_6395,N_6370);
nor U7083 (N_7083,N_6517,N_6212);
and U7084 (N_7084,N_6399,N_6139);
or U7085 (N_7085,N_6036,N_6109);
nand U7086 (N_7086,N_6076,N_6442);
and U7087 (N_7087,N_6284,N_6079);
nor U7088 (N_7088,N_6423,N_6554);
and U7089 (N_7089,N_6548,N_6167);
nor U7090 (N_7090,N_6494,N_6689);
or U7091 (N_7091,N_6160,N_6095);
nor U7092 (N_7092,N_6294,N_6400);
nand U7093 (N_7093,N_6100,N_6318);
or U7094 (N_7094,N_6580,N_6286);
nand U7095 (N_7095,N_6278,N_6737);
nor U7096 (N_7096,N_6089,N_6651);
nand U7097 (N_7097,N_6208,N_6151);
or U7098 (N_7098,N_6379,N_6170);
and U7099 (N_7099,N_6234,N_6565);
nand U7100 (N_7100,N_6178,N_6145);
nor U7101 (N_7101,N_6323,N_6501);
and U7102 (N_7102,N_6485,N_6659);
or U7103 (N_7103,N_6431,N_6694);
or U7104 (N_7104,N_6421,N_6209);
nand U7105 (N_7105,N_6583,N_6052);
nand U7106 (N_7106,N_6623,N_6480);
nand U7107 (N_7107,N_6574,N_6113);
or U7108 (N_7108,N_6644,N_6307);
nor U7109 (N_7109,N_6397,N_6358);
or U7110 (N_7110,N_6647,N_6711);
nor U7111 (N_7111,N_6031,N_6498);
and U7112 (N_7112,N_6215,N_6363);
nand U7113 (N_7113,N_6133,N_6600);
nor U7114 (N_7114,N_6707,N_6055);
nor U7115 (N_7115,N_6011,N_6186);
and U7116 (N_7116,N_6536,N_6684);
nand U7117 (N_7117,N_6242,N_6708);
and U7118 (N_7118,N_6228,N_6245);
nor U7119 (N_7119,N_6735,N_6450);
xor U7120 (N_7120,N_6027,N_6296);
nand U7121 (N_7121,N_6492,N_6232);
and U7122 (N_7122,N_6693,N_6037);
or U7123 (N_7123,N_6317,N_6122);
nor U7124 (N_7124,N_6434,N_6008);
and U7125 (N_7125,N_6554,N_6073);
or U7126 (N_7126,N_6052,N_6387);
nand U7127 (N_7127,N_6502,N_6467);
and U7128 (N_7128,N_6144,N_6418);
or U7129 (N_7129,N_6138,N_6562);
or U7130 (N_7130,N_6619,N_6217);
nand U7131 (N_7131,N_6057,N_6371);
nand U7132 (N_7132,N_6256,N_6219);
nand U7133 (N_7133,N_6657,N_6229);
nand U7134 (N_7134,N_6482,N_6220);
or U7135 (N_7135,N_6147,N_6312);
nand U7136 (N_7136,N_6360,N_6591);
nand U7137 (N_7137,N_6324,N_6450);
and U7138 (N_7138,N_6707,N_6175);
and U7139 (N_7139,N_6017,N_6386);
nand U7140 (N_7140,N_6626,N_6499);
xnor U7141 (N_7141,N_6509,N_6014);
or U7142 (N_7142,N_6523,N_6231);
nand U7143 (N_7143,N_6252,N_6468);
or U7144 (N_7144,N_6414,N_6083);
and U7145 (N_7145,N_6664,N_6011);
and U7146 (N_7146,N_6446,N_6688);
or U7147 (N_7147,N_6086,N_6221);
nand U7148 (N_7148,N_6226,N_6313);
nor U7149 (N_7149,N_6019,N_6516);
nor U7150 (N_7150,N_6558,N_6239);
nor U7151 (N_7151,N_6221,N_6156);
nand U7152 (N_7152,N_6646,N_6458);
or U7153 (N_7153,N_6526,N_6686);
and U7154 (N_7154,N_6747,N_6624);
and U7155 (N_7155,N_6676,N_6369);
nor U7156 (N_7156,N_6228,N_6625);
nor U7157 (N_7157,N_6673,N_6440);
nor U7158 (N_7158,N_6332,N_6667);
nor U7159 (N_7159,N_6198,N_6212);
or U7160 (N_7160,N_6503,N_6396);
nor U7161 (N_7161,N_6516,N_6087);
xor U7162 (N_7162,N_6064,N_6236);
or U7163 (N_7163,N_6721,N_6358);
and U7164 (N_7164,N_6404,N_6096);
or U7165 (N_7165,N_6131,N_6476);
nor U7166 (N_7166,N_6539,N_6329);
or U7167 (N_7167,N_6361,N_6059);
nor U7168 (N_7168,N_6571,N_6471);
and U7169 (N_7169,N_6351,N_6317);
xnor U7170 (N_7170,N_6027,N_6293);
or U7171 (N_7171,N_6255,N_6500);
nand U7172 (N_7172,N_6204,N_6542);
xnor U7173 (N_7173,N_6457,N_6582);
and U7174 (N_7174,N_6076,N_6623);
nor U7175 (N_7175,N_6508,N_6052);
or U7176 (N_7176,N_6151,N_6055);
and U7177 (N_7177,N_6297,N_6512);
or U7178 (N_7178,N_6439,N_6736);
nor U7179 (N_7179,N_6662,N_6346);
nor U7180 (N_7180,N_6061,N_6294);
and U7181 (N_7181,N_6298,N_6675);
nand U7182 (N_7182,N_6084,N_6556);
nor U7183 (N_7183,N_6371,N_6091);
and U7184 (N_7184,N_6230,N_6529);
nor U7185 (N_7185,N_6014,N_6452);
and U7186 (N_7186,N_6192,N_6253);
nor U7187 (N_7187,N_6456,N_6229);
xnor U7188 (N_7188,N_6677,N_6614);
nand U7189 (N_7189,N_6475,N_6204);
nor U7190 (N_7190,N_6068,N_6633);
or U7191 (N_7191,N_6221,N_6333);
nor U7192 (N_7192,N_6537,N_6438);
nor U7193 (N_7193,N_6087,N_6351);
nand U7194 (N_7194,N_6183,N_6079);
nor U7195 (N_7195,N_6742,N_6326);
or U7196 (N_7196,N_6337,N_6250);
nor U7197 (N_7197,N_6015,N_6313);
xor U7198 (N_7198,N_6244,N_6233);
or U7199 (N_7199,N_6053,N_6388);
nand U7200 (N_7200,N_6362,N_6431);
nand U7201 (N_7201,N_6465,N_6331);
xor U7202 (N_7202,N_6285,N_6687);
and U7203 (N_7203,N_6252,N_6683);
or U7204 (N_7204,N_6251,N_6550);
nor U7205 (N_7205,N_6500,N_6318);
and U7206 (N_7206,N_6297,N_6345);
or U7207 (N_7207,N_6244,N_6075);
nor U7208 (N_7208,N_6288,N_6044);
nand U7209 (N_7209,N_6171,N_6432);
or U7210 (N_7210,N_6153,N_6612);
nor U7211 (N_7211,N_6496,N_6259);
nor U7212 (N_7212,N_6065,N_6642);
or U7213 (N_7213,N_6057,N_6024);
and U7214 (N_7214,N_6470,N_6299);
and U7215 (N_7215,N_6228,N_6210);
xor U7216 (N_7216,N_6112,N_6037);
nand U7217 (N_7217,N_6463,N_6357);
and U7218 (N_7218,N_6467,N_6597);
and U7219 (N_7219,N_6304,N_6361);
and U7220 (N_7220,N_6223,N_6282);
nor U7221 (N_7221,N_6119,N_6725);
nor U7222 (N_7222,N_6635,N_6286);
and U7223 (N_7223,N_6004,N_6489);
or U7224 (N_7224,N_6314,N_6674);
xnor U7225 (N_7225,N_6121,N_6387);
nand U7226 (N_7226,N_6318,N_6182);
nand U7227 (N_7227,N_6046,N_6464);
nor U7228 (N_7228,N_6520,N_6182);
and U7229 (N_7229,N_6644,N_6161);
nand U7230 (N_7230,N_6698,N_6246);
nor U7231 (N_7231,N_6344,N_6293);
or U7232 (N_7232,N_6227,N_6643);
xnor U7233 (N_7233,N_6231,N_6399);
nor U7234 (N_7234,N_6322,N_6545);
xnor U7235 (N_7235,N_6017,N_6272);
nor U7236 (N_7236,N_6051,N_6362);
and U7237 (N_7237,N_6329,N_6012);
xnor U7238 (N_7238,N_6744,N_6365);
and U7239 (N_7239,N_6113,N_6037);
nor U7240 (N_7240,N_6440,N_6595);
xor U7241 (N_7241,N_6347,N_6460);
nor U7242 (N_7242,N_6399,N_6150);
nand U7243 (N_7243,N_6634,N_6619);
nand U7244 (N_7244,N_6651,N_6601);
nand U7245 (N_7245,N_6570,N_6152);
xor U7246 (N_7246,N_6135,N_6229);
and U7247 (N_7247,N_6409,N_6181);
or U7248 (N_7248,N_6517,N_6131);
nand U7249 (N_7249,N_6592,N_6669);
or U7250 (N_7250,N_6423,N_6139);
or U7251 (N_7251,N_6525,N_6418);
or U7252 (N_7252,N_6228,N_6481);
and U7253 (N_7253,N_6465,N_6460);
nor U7254 (N_7254,N_6074,N_6594);
or U7255 (N_7255,N_6230,N_6607);
nor U7256 (N_7256,N_6295,N_6091);
nor U7257 (N_7257,N_6449,N_6269);
nor U7258 (N_7258,N_6480,N_6241);
or U7259 (N_7259,N_6552,N_6691);
nand U7260 (N_7260,N_6732,N_6441);
and U7261 (N_7261,N_6449,N_6073);
nor U7262 (N_7262,N_6075,N_6040);
and U7263 (N_7263,N_6462,N_6564);
or U7264 (N_7264,N_6026,N_6327);
nor U7265 (N_7265,N_6086,N_6452);
nand U7266 (N_7266,N_6371,N_6578);
xor U7267 (N_7267,N_6390,N_6071);
nor U7268 (N_7268,N_6653,N_6304);
nor U7269 (N_7269,N_6073,N_6539);
nor U7270 (N_7270,N_6509,N_6353);
or U7271 (N_7271,N_6206,N_6272);
nand U7272 (N_7272,N_6510,N_6285);
xnor U7273 (N_7273,N_6593,N_6381);
nand U7274 (N_7274,N_6671,N_6260);
nor U7275 (N_7275,N_6474,N_6504);
or U7276 (N_7276,N_6173,N_6638);
or U7277 (N_7277,N_6175,N_6162);
xor U7278 (N_7278,N_6181,N_6404);
or U7279 (N_7279,N_6556,N_6660);
or U7280 (N_7280,N_6069,N_6596);
nor U7281 (N_7281,N_6693,N_6573);
xnor U7282 (N_7282,N_6341,N_6502);
xnor U7283 (N_7283,N_6112,N_6262);
and U7284 (N_7284,N_6521,N_6429);
or U7285 (N_7285,N_6614,N_6173);
nand U7286 (N_7286,N_6290,N_6049);
and U7287 (N_7287,N_6169,N_6741);
nor U7288 (N_7288,N_6330,N_6126);
xor U7289 (N_7289,N_6223,N_6197);
nand U7290 (N_7290,N_6737,N_6105);
or U7291 (N_7291,N_6109,N_6485);
and U7292 (N_7292,N_6681,N_6337);
or U7293 (N_7293,N_6113,N_6190);
xnor U7294 (N_7294,N_6108,N_6544);
nand U7295 (N_7295,N_6252,N_6731);
nor U7296 (N_7296,N_6722,N_6646);
and U7297 (N_7297,N_6416,N_6035);
and U7298 (N_7298,N_6208,N_6432);
xor U7299 (N_7299,N_6061,N_6001);
or U7300 (N_7300,N_6073,N_6735);
xnor U7301 (N_7301,N_6121,N_6500);
nor U7302 (N_7302,N_6368,N_6481);
and U7303 (N_7303,N_6026,N_6328);
nand U7304 (N_7304,N_6297,N_6133);
nor U7305 (N_7305,N_6732,N_6128);
or U7306 (N_7306,N_6532,N_6478);
nor U7307 (N_7307,N_6202,N_6350);
and U7308 (N_7308,N_6573,N_6341);
and U7309 (N_7309,N_6597,N_6425);
nor U7310 (N_7310,N_6276,N_6539);
nor U7311 (N_7311,N_6398,N_6435);
nand U7312 (N_7312,N_6119,N_6377);
nor U7313 (N_7313,N_6278,N_6082);
xor U7314 (N_7314,N_6188,N_6098);
or U7315 (N_7315,N_6672,N_6490);
or U7316 (N_7316,N_6445,N_6448);
or U7317 (N_7317,N_6439,N_6397);
nand U7318 (N_7318,N_6014,N_6243);
nor U7319 (N_7319,N_6414,N_6124);
and U7320 (N_7320,N_6062,N_6046);
nand U7321 (N_7321,N_6278,N_6492);
nand U7322 (N_7322,N_6587,N_6253);
nand U7323 (N_7323,N_6029,N_6439);
or U7324 (N_7324,N_6125,N_6510);
nor U7325 (N_7325,N_6068,N_6204);
nor U7326 (N_7326,N_6459,N_6038);
nand U7327 (N_7327,N_6035,N_6712);
nand U7328 (N_7328,N_6556,N_6696);
nor U7329 (N_7329,N_6272,N_6673);
and U7330 (N_7330,N_6299,N_6220);
nand U7331 (N_7331,N_6229,N_6687);
and U7332 (N_7332,N_6310,N_6291);
or U7333 (N_7333,N_6443,N_6517);
nand U7334 (N_7334,N_6104,N_6684);
and U7335 (N_7335,N_6516,N_6298);
xnor U7336 (N_7336,N_6056,N_6464);
xor U7337 (N_7337,N_6214,N_6154);
or U7338 (N_7338,N_6594,N_6349);
xnor U7339 (N_7339,N_6392,N_6115);
or U7340 (N_7340,N_6686,N_6509);
and U7341 (N_7341,N_6260,N_6490);
xor U7342 (N_7342,N_6497,N_6096);
or U7343 (N_7343,N_6361,N_6273);
or U7344 (N_7344,N_6438,N_6236);
xnor U7345 (N_7345,N_6383,N_6537);
nor U7346 (N_7346,N_6422,N_6624);
or U7347 (N_7347,N_6722,N_6064);
and U7348 (N_7348,N_6649,N_6307);
nor U7349 (N_7349,N_6329,N_6692);
or U7350 (N_7350,N_6116,N_6670);
xnor U7351 (N_7351,N_6652,N_6018);
nand U7352 (N_7352,N_6723,N_6130);
or U7353 (N_7353,N_6587,N_6058);
nand U7354 (N_7354,N_6502,N_6407);
xnor U7355 (N_7355,N_6249,N_6472);
nor U7356 (N_7356,N_6455,N_6558);
nand U7357 (N_7357,N_6706,N_6391);
nor U7358 (N_7358,N_6035,N_6257);
or U7359 (N_7359,N_6407,N_6308);
nand U7360 (N_7360,N_6414,N_6278);
or U7361 (N_7361,N_6379,N_6110);
and U7362 (N_7362,N_6586,N_6093);
nor U7363 (N_7363,N_6661,N_6264);
and U7364 (N_7364,N_6282,N_6729);
and U7365 (N_7365,N_6476,N_6032);
nor U7366 (N_7366,N_6428,N_6271);
nor U7367 (N_7367,N_6254,N_6075);
nand U7368 (N_7368,N_6684,N_6230);
nand U7369 (N_7369,N_6404,N_6467);
and U7370 (N_7370,N_6454,N_6108);
and U7371 (N_7371,N_6356,N_6183);
nand U7372 (N_7372,N_6438,N_6163);
and U7373 (N_7373,N_6647,N_6091);
xor U7374 (N_7374,N_6444,N_6509);
nand U7375 (N_7375,N_6259,N_6370);
nand U7376 (N_7376,N_6712,N_6681);
nor U7377 (N_7377,N_6244,N_6418);
or U7378 (N_7378,N_6581,N_6441);
nand U7379 (N_7379,N_6013,N_6723);
nand U7380 (N_7380,N_6429,N_6443);
or U7381 (N_7381,N_6166,N_6061);
nand U7382 (N_7382,N_6000,N_6732);
nand U7383 (N_7383,N_6628,N_6479);
and U7384 (N_7384,N_6070,N_6162);
and U7385 (N_7385,N_6560,N_6265);
or U7386 (N_7386,N_6354,N_6666);
nand U7387 (N_7387,N_6510,N_6184);
nand U7388 (N_7388,N_6476,N_6575);
and U7389 (N_7389,N_6164,N_6078);
or U7390 (N_7390,N_6255,N_6482);
nor U7391 (N_7391,N_6554,N_6348);
nand U7392 (N_7392,N_6544,N_6305);
xnor U7393 (N_7393,N_6446,N_6651);
xnor U7394 (N_7394,N_6725,N_6419);
nor U7395 (N_7395,N_6555,N_6196);
xnor U7396 (N_7396,N_6070,N_6196);
and U7397 (N_7397,N_6399,N_6609);
and U7398 (N_7398,N_6283,N_6137);
nor U7399 (N_7399,N_6680,N_6568);
nand U7400 (N_7400,N_6748,N_6107);
nor U7401 (N_7401,N_6366,N_6615);
and U7402 (N_7402,N_6339,N_6046);
xnor U7403 (N_7403,N_6289,N_6100);
nand U7404 (N_7404,N_6368,N_6460);
nand U7405 (N_7405,N_6510,N_6119);
and U7406 (N_7406,N_6217,N_6603);
nand U7407 (N_7407,N_6297,N_6714);
xnor U7408 (N_7408,N_6387,N_6679);
or U7409 (N_7409,N_6468,N_6078);
and U7410 (N_7410,N_6312,N_6212);
nor U7411 (N_7411,N_6349,N_6083);
nor U7412 (N_7412,N_6586,N_6259);
or U7413 (N_7413,N_6668,N_6580);
or U7414 (N_7414,N_6347,N_6171);
or U7415 (N_7415,N_6536,N_6637);
or U7416 (N_7416,N_6551,N_6429);
nor U7417 (N_7417,N_6610,N_6314);
nand U7418 (N_7418,N_6109,N_6650);
nor U7419 (N_7419,N_6390,N_6072);
or U7420 (N_7420,N_6505,N_6554);
and U7421 (N_7421,N_6527,N_6258);
and U7422 (N_7422,N_6424,N_6074);
xor U7423 (N_7423,N_6420,N_6216);
and U7424 (N_7424,N_6005,N_6722);
or U7425 (N_7425,N_6469,N_6104);
and U7426 (N_7426,N_6699,N_6301);
nor U7427 (N_7427,N_6661,N_6248);
nor U7428 (N_7428,N_6663,N_6237);
nand U7429 (N_7429,N_6039,N_6330);
nand U7430 (N_7430,N_6593,N_6086);
nor U7431 (N_7431,N_6732,N_6568);
nor U7432 (N_7432,N_6142,N_6729);
nand U7433 (N_7433,N_6200,N_6384);
nand U7434 (N_7434,N_6046,N_6393);
xnor U7435 (N_7435,N_6172,N_6201);
or U7436 (N_7436,N_6259,N_6393);
nand U7437 (N_7437,N_6564,N_6477);
xnor U7438 (N_7438,N_6128,N_6594);
or U7439 (N_7439,N_6509,N_6320);
and U7440 (N_7440,N_6197,N_6678);
nand U7441 (N_7441,N_6539,N_6030);
nand U7442 (N_7442,N_6674,N_6572);
and U7443 (N_7443,N_6733,N_6584);
nand U7444 (N_7444,N_6659,N_6427);
nand U7445 (N_7445,N_6180,N_6197);
nor U7446 (N_7446,N_6235,N_6019);
and U7447 (N_7447,N_6007,N_6670);
and U7448 (N_7448,N_6630,N_6620);
nand U7449 (N_7449,N_6723,N_6566);
nor U7450 (N_7450,N_6544,N_6238);
or U7451 (N_7451,N_6191,N_6277);
and U7452 (N_7452,N_6744,N_6112);
and U7453 (N_7453,N_6375,N_6037);
nand U7454 (N_7454,N_6444,N_6492);
nor U7455 (N_7455,N_6397,N_6498);
or U7456 (N_7456,N_6136,N_6339);
or U7457 (N_7457,N_6598,N_6094);
or U7458 (N_7458,N_6035,N_6558);
or U7459 (N_7459,N_6155,N_6156);
and U7460 (N_7460,N_6394,N_6636);
nor U7461 (N_7461,N_6211,N_6717);
nor U7462 (N_7462,N_6037,N_6440);
nand U7463 (N_7463,N_6544,N_6600);
or U7464 (N_7464,N_6731,N_6066);
nand U7465 (N_7465,N_6722,N_6426);
nand U7466 (N_7466,N_6490,N_6319);
nor U7467 (N_7467,N_6466,N_6642);
and U7468 (N_7468,N_6178,N_6736);
nor U7469 (N_7469,N_6312,N_6556);
nor U7470 (N_7470,N_6166,N_6319);
and U7471 (N_7471,N_6145,N_6646);
nand U7472 (N_7472,N_6651,N_6697);
or U7473 (N_7473,N_6723,N_6335);
nor U7474 (N_7474,N_6129,N_6277);
or U7475 (N_7475,N_6419,N_6108);
nor U7476 (N_7476,N_6049,N_6481);
xor U7477 (N_7477,N_6528,N_6359);
xnor U7478 (N_7478,N_6390,N_6420);
and U7479 (N_7479,N_6502,N_6151);
or U7480 (N_7480,N_6623,N_6270);
or U7481 (N_7481,N_6655,N_6480);
nand U7482 (N_7482,N_6274,N_6326);
nand U7483 (N_7483,N_6172,N_6464);
and U7484 (N_7484,N_6617,N_6058);
nand U7485 (N_7485,N_6734,N_6048);
nand U7486 (N_7486,N_6450,N_6188);
and U7487 (N_7487,N_6615,N_6469);
nand U7488 (N_7488,N_6507,N_6365);
nor U7489 (N_7489,N_6029,N_6168);
nor U7490 (N_7490,N_6713,N_6628);
or U7491 (N_7491,N_6537,N_6215);
or U7492 (N_7492,N_6093,N_6163);
or U7493 (N_7493,N_6347,N_6107);
xor U7494 (N_7494,N_6158,N_6367);
or U7495 (N_7495,N_6379,N_6302);
nand U7496 (N_7496,N_6505,N_6722);
and U7497 (N_7497,N_6664,N_6274);
nor U7498 (N_7498,N_6537,N_6516);
nand U7499 (N_7499,N_6711,N_6085);
and U7500 (N_7500,N_7252,N_7448);
xnor U7501 (N_7501,N_7301,N_6756);
nor U7502 (N_7502,N_7186,N_7456);
or U7503 (N_7503,N_7450,N_7294);
or U7504 (N_7504,N_7395,N_6846);
or U7505 (N_7505,N_7173,N_7002);
nand U7506 (N_7506,N_6886,N_7164);
or U7507 (N_7507,N_6927,N_7220);
and U7508 (N_7508,N_7290,N_7113);
nor U7509 (N_7509,N_7352,N_7457);
and U7510 (N_7510,N_7063,N_7052);
nand U7511 (N_7511,N_7179,N_6992);
nand U7512 (N_7512,N_7099,N_6961);
xor U7513 (N_7513,N_7488,N_7243);
nor U7514 (N_7514,N_7137,N_7271);
nor U7515 (N_7515,N_6754,N_7462);
nor U7516 (N_7516,N_6903,N_6928);
xnor U7517 (N_7517,N_7427,N_6883);
and U7518 (N_7518,N_7327,N_7171);
nand U7519 (N_7519,N_7483,N_7471);
and U7520 (N_7520,N_7323,N_7348);
and U7521 (N_7521,N_7480,N_6847);
or U7522 (N_7522,N_7041,N_7221);
nand U7523 (N_7523,N_6974,N_7151);
nand U7524 (N_7524,N_7429,N_6769);
nand U7525 (N_7525,N_7245,N_7250);
xor U7526 (N_7526,N_7496,N_6983);
and U7527 (N_7527,N_6854,N_7085);
nand U7528 (N_7528,N_7307,N_7414);
xnor U7529 (N_7529,N_6750,N_7108);
nor U7530 (N_7530,N_7451,N_7343);
nor U7531 (N_7531,N_6791,N_6773);
nor U7532 (N_7532,N_6996,N_6822);
and U7533 (N_7533,N_7117,N_7268);
nand U7534 (N_7534,N_7042,N_7053);
nor U7535 (N_7535,N_6863,N_6957);
or U7536 (N_7536,N_6884,N_7235);
nor U7537 (N_7537,N_6840,N_7421);
nand U7538 (N_7538,N_7124,N_6971);
and U7539 (N_7539,N_6829,N_7435);
nor U7540 (N_7540,N_6765,N_6782);
xor U7541 (N_7541,N_6856,N_7350);
nor U7542 (N_7542,N_6826,N_7198);
nand U7543 (N_7543,N_7407,N_7094);
xnor U7544 (N_7544,N_6965,N_7300);
nor U7545 (N_7545,N_7400,N_7434);
nand U7546 (N_7546,N_7358,N_7060);
nand U7547 (N_7547,N_6838,N_6799);
or U7548 (N_7548,N_7375,N_7230);
nand U7549 (N_7549,N_7396,N_6953);
nor U7550 (N_7550,N_6873,N_7177);
and U7551 (N_7551,N_6875,N_6979);
or U7552 (N_7552,N_6841,N_6923);
nand U7553 (N_7553,N_7494,N_7283);
or U7554 (N_7554,N_6760,N_7383);
xnor U7555 (N_7555,N_7026,N_6810);
or U7556 (N_7556,N_6850,N_7285);
and U7557 (N_7557,N_7364,N_6817);
and U7558 (N_7558,N_6946,N_7382);
nor U7559 (N_7559,N_7191,N_6805);
nand U7560 (N_7560,N_7184,N_6955);
nor U7561 (N_7561,N_7325,N_7266);
nand U7562 (N_7562,N_7253,N_6786);
and U7563 (N_7563,N_6945,N_6894);
nand U7564 (N_7564,N_7188,N_7234);
and U7565 (N_7565,N_6929,N_6792);
xor U7566 (N_7566,N_7430,N_7167);
nand U7567 (N_7567,N_6998,N_7201);
or U7568 (N_7568,N_7411,N_6950);
and U7569 (N_7569,N_7306,N_7463);
xnor U7570 (N_7570,N_7373,N_7147);
nor U7571 (N_7571,N_7438,N_7021);
xor U7572 (N_7572,N_7247,N_7155);
nand U7573 (N_7573,N_7013,N_6866);
and U7574 (N_7574,N_7485,N_7455);
or U7575 (N_7575,N_6888,N_7029);
and U7576 (N_7576,N_7061,N_7114);
nor U7577 (N_7577,N_6755,N_7009);
nand U7578 (N_7578,N_7410,N_6823);
and U7579 (N_7579,N_7461,N_7134);
and U7580 (N_7580,N_7102,N_7474);
nor U7581 (N_7581,N_7418,N_7272);
and U7582 (N_7582,N_7062,N_6959);
and U7583 (N_7583,N_6778,N_6892);
nand U7584 (N_7584,N_7016,N_7491);
nand U7585 (N_7585,N_7412,N_7340);
or U7586 (N_7586,N_7424,N_7088);
xor U7587 (N_7587,N_7187,N_6993);
nor U7588 (N_7588,N_7467,N_7401);
or U7589 (N_7589,N_7490,N_6942);
nor U7590 (N_7590,N_7317,N_7073);
or U7591 (N_7591,N_7329,N_7154);
or U7592 (N_7592,N_7444,N_7215);
nand U7593 (N_7593,N_7354,N_7443);
nor U7594 (N_7594,N_7050,N_7034);
nand U7595 (N_7595,N_7032,N_7116);
or U7596 (N_7596,N_7022,N_7043);
xnor U7597 (N_7597,N_7078,N_7111);
nor U7598 (N_7598,N_6815,N_6989);
xnor U7599 (N_7599,N_7189,N_6776);
nor U7600 (N_7600,N_7428,N_7075);
or U7601 (N_7601,N_6868,N_6816);
or U7602 (N_7602,N_7148,N_7242);
nand U7603 (N_7603,N_7241,N_7058);
nand U7604 (N_7604,N_7292,N_6939);
or U7605 (N_7605,N_6807,N_7399);
and U7606 (N_7606,N_7464,N_6811);
nand U7607 (N_7607,N_7475,N_7105);
nor U7608 (N_7608,N_7251,N_6970);
or U7609 (N_7609,N_7479,N_6862);
or U7610 (N_7610,N_7129,N_7036);
nor U7611 (N_7611,N_6844,N_7087);
or U7612 (N_7612,N_7093,N_7020);
or U7613 (N_7613,N_6848,N_6907);
or U7614 (N_7614,N_7135,N_7387);
xnor U7615 (N_7615,N_6858,N_6855);
xnor U7616 (N_7616,N_7007,N_7370);
or U7617 (N_7617,N_6980,N_6766);
nor U7618 (N_7618,N_7205,N_7442);
and U7619 (N_7619,N_6908,N_6825);
nor U7620 (N_7620,N_6801,N_7472);
and U7621 (N_7621,N_6882,N_7083);
nor U7622 (N_7622,N_7279,N_6896);
xnor U7623 (N_7623,N_7153,N_7328);
nand U7624 (N_7624,N_6885,N_7112);
nor U7625 (N_7625,N_6762,N_7469);
nand U7626 (N_7626,N_7057,N_7367);
or U7627 (N_7627,N_7195,N_7107);
and U7628 (N_7628,N_6917,N_7006);
and U7629 (N_7629,N_7059,N_6870);
or U7630 (N_7630,N_7000,N_7084);
nand U7631 (N_7631,N_7017,N_7183);
nor U7632 (N_7632,N_6851,N_6981);
nand U7633 (N_7633,N_6877,N_6872);
nor U7634 (N_7634,N_7366,N_6947);
xor U7635 (N_7635,N_7030,N_7152);
and U7636 (N_7636,N_7180,N_7371);
or U7637 (N_7637,N_6865,N_7048);
or U7638 (N_7638,N_7118,N_7489);
or U7639 (N_7639,N_7357,N_6861);
and U7640 (N_7640,N_7031,N_7257);
xnor U7641 (N_7641,N_7047,N_7012);
or U7642 (N_7642,N_7406,N_7288);
and U7643 (N_7643,N_6804,N_7092);
nor U7644 (N_7644,N_6770,N_7132);
xor U7645 (N_7645,N_6753,N_6914);
or U7646 (N_7646,N_7403,N_7123);
or U7647 (N_7647,N_7299,N_7273);
or U7648 (N_7648,N_7284,N_6781);
or U7649 (N_7649,N_6975,N_7206);
nor U7650 (N_7650,N_7281,N_7368);
and U7651 (N_7651,N_7238,N_7003);
nand U7652 (N_7652,N_7244,N_7498);
or U7653 (N_7653,N_7199,N_7100);
or U7654 (N_7654,N_6797,N_7361);
and U7655 (N_7655,N_7072,N_7374);
and U7656 (N_7656,N_6982,N_7004);
nor U7657 (N_7657,N_7404,N_7274);
xor U7658 (N_7658,N_7381,N_7495);
nor U7659 (N_7659,N_6839,N_7385);
or U7660 (N_7660,N_7265,N_6969);
or U7661 (N_7661,N_7440,N_7321);
nand U7662 (N_7662,N_7351,N_7138);
xnor U7663 (N_7663,N_7228,N_7332);
or U7664 (N_7664,N_6964,N_7202);
nor U7665 (N_7665,N_7207,N_7419);
and U7666 (N_7666,N_7293,N_6808);
nor U7667 (N_7667,N_6911,N_6915);
nor U7668 (N_7668,N_7033,N_6900);
nand U7669 (N_7669,N_7477,N_6785);
xnor U7670 (N_7670,N_6788,N_7260);
or U7671 (N_7671,N_6830,N_7453);
nand U7672 (N_7672,N_7181,N_7203);
nand U7673 (N_7673,N_7222,N_6941);
xor U7674 (N_7674,N_7096,N_7185);
or U7675 (N_7675,N_6832,N_7001);
or U7676 (N_7676,N_6890,N_7255);
or U7677 (N_7677,N_7277,N_7125);
or U7678 (N_7678,N_6889,N_7344);
or U7679 (N_7679,N_7077,N_7433);
xor U7680 (N_7680,N_7143,N_7018);
nand U7681 (N_7681,N_7178,N_6921);
nor U7682 (N_7682,N_7101,N_6887);
or U7683 (N_7683,N_7109,N_7169);
and U7684 (N_7684,N_6906,N_7054);
or U7685 (N_7685,N_7158,N_6940);
nand U7686 (N_7686,N_6800,N_7011);
or U7687 (N_7687,N_7263,N_7345);
or U7688 (N_7688,N_6876,N_7342);
nor U7689 (N_7689,N_6835,N_6904);
or U7690 (N_7690,N_6794,N_7445);
xnor U7691 (N_7691,N_7226,N_6834);
nor U7692 (N_7692,N_7303,N_7156);
nand U7693 (N_7693,N_7209,N_6930);
and U7694 (N_7694,N_6818,N_6952);
and U7695 (N_7695,N_7286,N_6925);
and U7696 (N_7696,N_7338,N_7076);
and U7697 (N_7697,N_7311,N_6775);
or U7698 (N_7698,N_7454,N_6968);
or U7699 (N_7699,N_7055,N_7090);
and U7700 (N_7700,N_6936,N_7175);
xor U7701 (N_7701,N_7259,N_7081);
nand U7702 (N_7702,N_6779,N_6771);
nor U7703 (N_7703,N_6912,N_6764);
and U7704 (N_7704,N_7258,N_6819);
or U7705 (N_7705,N_6789,N_7333);
nand U7706 (N_7706,N_7024,N_7097);
xor U7707 (N_7707,N_7027,N_7256);
and U7708 (N_7708,N_7380,N_6757);
and U7709 (N_7709,N_6871,N_6898);
and U7710 (N_7710,N_6780,N_7231);
nor U7711 (N_7711,N_7409,N_7334);
and U7712 (N_7712,N_7145,N_7349);
or U7713 (N_7713,N_7104,N_7240);
xor U7714 (N_7714,N_6878,N_6767);
nor U7715 (N_7715,N_6933,N_7216);
xor U7716 (N_7716,N_6820,N_7172);
and U7717 (N_7717,N_6976,N_7160);
nor U7718 (N_7718,N_7356,N_6763);
nor U7719 (N_7719,N_7074,N_7170);
and U7720 (N_7720,N_7282,N_7405);
xor U7721 (N_7721,N_7459,N_7008);
nand U7722 (N_7722,N_7478,N_7149);
nor U7723 (N_7723,N_7131,N_6798);
nor U7724 (N_7724,N_7389,N_7355);
or U7725 (N_7725,N_7128,N_6951);
and U7726 (N_7726,N_7261,N_7233);
or U7727 (N_7727,N_6956,N_6902);
nand U7728 (N_7728,N_6948,N_6836);
and U7729 (N_7729,N_7388,N_7064);
and U7730 (N_7730,N_7377,N_6938);
nor U7731 (N_7731,N_7197,N_6853);
and U7732 (N_7732,N_6893,N_7497);
or U7733 (N_7733,N_7136,N_7103);
and U7734 (N_7734,N_7331,N_6920);
or U7735 (N_7735,N_6901,N_6772);
or U7736 (N_7736,N_7067,N_7079);
nand U7737 (N_7737,N_7229,N_7082);
or U7738 (N_7738,N_7378,N_7213);
nand U7739 (N_7739,N_6897,N_7210);
or U7740 (N_7740,N_7436,N_6913);
or U7741 (N_7741,N_7095,N_7441);
xnor U7742 (N_7742,N_7417,N_7130);
nor U7743 (N_7743,N_6919,N_7318);
and U7744 (N_7744,N_7248,N_7165);
nor U7745 (N_7745,N_7425,N_6999);
nand U7746 (N_7746,N_7360,N_7308);
and U7747 (N_7747,N_7174,N_7468);
or U7748 (N_7748,N_6963,N_7280);
nand U7749 (N_7749,N_6995,N_7142);
or U7750 (N_7750,N_6899,N_7275);
nand U7751 (N_7751,N_7014,N_7264);
or U7752 (N_7752,N_7304,N_7010);
and U7753 (N_7753,N_7359,N_7365);
xor U7754 (N_7754,N_6879,N_7267);
xor U7755 (N_7755,N_7449,N_7319);
and U7756 (N_7756,N_6960,N_6849);
and U7757 (N_7757,N_6935,N_7019);
or U7758 (N_7758,N_6958,N_6944);
and U7759 (N_7759,N_6937,N_7347);
nor U7760 (N_7760,N_6783,N_7484);
or U7761 (N_7761,N_7316,N_7499);
or U7762 (N_7762,N_7163,N_7068);
nor U7763 (N_7763,N_7040,N_7056);
nand U7764 (N_7764,N_7394,N_6802);
xor U7765 (N_7765,N_6795,N_6926);
and U7766 (N_7766,N_7091,N_7106);
and U7767 (N_7767,N_6833,N_7446);
nor U7768 (N_7768,N_7420,N_7150);
nand U7769 (N_7769,N_6905,N_7326);
nand U7770 (N_7770,N_7372,N_6949);
xnor U7771 (N_7771,N_6852,N_7098);
nand U7772 (N_7772,N_6977,N_7402);
or U7773 (N_7773,N_7276,N_7289);
nand U7774 (N_7774,N_7071,N_7127);
nand U7775 (N_7775,N_7126,N_7162);
nand U7776 (N_7776,N_7080,N_7139);
or U7777 (N_7777,N_7437,N_7422);
nand U7778 (N_7778,N_7346,N_7362);
nor U7779 (N_7779,N_7470,N_6891);
or U7780 (N_7780,N_6978,N_7341);
nand U7781 (N_7781,N_7298,N_7159);
and U7782 (N_7782,N_6813,N_6984);
and U7783 (N_7783,N_7270,N_7232);
nor U7784 (N_7784,N_7295,N_6831);
nor U7785 (N_7785,N_7335,N_7214);
nand U7786 (N_7786,N_7320,N_7376);
nand U7787 (N_7787,N_6828,N_7391);
nor U7788 (N_7788,N_7465,N_7168);
and U7789 (N_7789,N_7431,N_7296);
nor U7790 (N_7790,N_7119,N_6759);
nand U7791 (N_7791,N_7144,N_6931);
nor U7792 (N_7792,N_7493,N_7458);
nand U7793 (N_7793,N_7069,N_7302);
and U7794 (N_7794,N_7416,N_7190);
or U7795 (N_7795,N_7432,N_7035);
nor U7796 (N_7796,N_7146,N_6934);
nand U7797 (N_7797,N_7314,N_7278);
nor U7798 (N_7798,N_6790,N_7262);
nor U7799 (N_7799,N_6784,N_7310);
or U7800 (N_7800,N_6967,N_7120);
or U7801 (N_7801,N_6752,N_6843);
xor U7802 (N_7802,N_7313,N_6809);
nand U7803 (N_7803,N_6972,N_7386);
nand U7804 (N_7804,N_6814,N_6758);
xor U7805 (N_7805,N_7208,N_7487);
or U7806 (N_7806,N_6803,N_7397);
nand U7807 (N_7807,N_7415,N_7045);
and U7808 (N_7808,N_7161,N_7223);
nor U7809 (N_7809,N_7196,N_7037);
nor U7810 (N_7810,N_7312,N_7028);
nor U7811 (N_7811,N_7212,N_7269);
nand U7812 (N_7812,N_6932,N_6774);
or U7813 (N_7813,N_7051,N_7413);
and U7814 (N_7814,N_6954,N_6880);
nand U7815 (N_7815,N_7460,N_7339);
nor U7816 (N_7816,N_7481,N_7423);
and U7817 (N_7817,N_7254,N_7140);
or U7818 (N_7818,N_7249,N_7287);
and U7819 (N_7819,N_7086,N_7291);
nand U7820 (N_7820,N_7211,N_7049);
and U7821 (N_7821,N_7336,N_6864);
nand U7822 (N_7822,N_6869,N_7426);
nand U7823 (N_7823,N_7353,N_6962);
and U7824 (N_7824,N_7392,N_6997);
nor U7825 (N_7825,N_6988,N_6918);
nor U7826 (N_7826,N_6909,N_6859);
and U7827 (N_7827,N_7070,N_7157);
nor U7828 (N_7828,N_7141,N_7297);
or U7829 (N_7829,N_7217,N_7039);
nand U7830 (N_7830,N_6777,N_7066);
or U7831 (N_7831,N_7315,N_7218);
or U7832 (N_7832,N_7393,N_6860);
or U7833 (N_7833,N_7398,N_7015);
nor U7834 (N_7834,N_7246,N_6986);
and U7835 (N_7835,N_7492,N_6806);
or U7836 (N_7836,N_6837,N_7239);
or U7837 (N_7837,N_7193,N_6827);
nand U7838 (N_7838,N_7005,N_6973);
or U7839 (N_7839,N_7182,N_6994);
xor U7840 (N_7840,N_7447,N_6924);
and U7841 (N_7841,N_7473,N_7482);
or U7842 (N_7842,N_7237,N_6990);
nand U7843 (N_7843,N_6812,N_6987);
nand U7844 (N_7844,N_6751,N_6916);
and U7845 (N_7845,N_6985,N_7322);
nand U7846 (N_7846,N_7452,N_7408);
xor U7847 (N_7847,N_7236,N_6796);
or U7848 (N_7848,N_7133,N_7204);
and U7849 (N_7849,N_7390,N_7224);
nor U7850 (N_7850,N_6966,N_7227);
nand U7851 (N_7851,N_7379,N_7486);
nor U7852 (N_7852,N_7384,N_7121);
or U7853 (N_7853,N_7466,N_7065);
or U7854 (N_7854,N_6857,N_6793);
or U7855 (N_7855,N_7089,N_7025);
and U7856 (N_7856,N_7439,N_6881);
nand U7857 (N_7857,N_6821,N_6910);
nor U7858 (N_7858,N_6845,N_7192);
and U7859 (N_7859,N_7200,N_7176);
nor U7860 (N_7860,N_6824,N_7023);
and U7861 (N_7861,N_7194,N_6842);
and U7862 (N_7862,N_6768,N_7225);
nand U7863 (N_7863,N_7110,N_7330);
nor U7864 (N_7864,N_7038,N_7122);
xnor U7865 (N_7865,N_6787,N_7369);
or U7866 (N_7866,N_7337,N_7363);
or U7867 (N_7867,N_6943,N_7166);
nor U7868 (N_7868,N_7309,N_7046);
or U7869 (N_7869,N_7305,N_6761);
and U7870 (N_7870,N_7044,N_6922);
nor U7871 (N_7871,N_6895,N_7324);
nor U7872 (N_7872,N_7476,N_6991);
nor U7873 (N_7873,N_6867,N_7219);
nor U7874 (N_7874,N_7115,N_6874);
and U7875 (N_7875,N_7147,N_6998);
nand U7876 (N_7876,N_7009,N_6921);
nor U7877 (N_7877,N_7017,N_7254);
or U7878 (N_7878,N_6841,N_6889);
or U7879 (N_7879,N_7206,N_7147);
nand U7880 (N_7880,N_7367,N_6900);
or U7881 (N_7881,N_7069,N_6773);
and U7882 (N_7882,N_7314,N_6755);
xnor U7883 (N_7883,N_6917,N_6879);
nor U7884 (N_7884,N_7456,N_7224);
or U7885 (N_7885,N_6978,N_7086);
or U7886 (N_7886,N_7486,N_7437);
or U7887 (N_7887,N_6808,N_7467);
nand U7888 (N_7888,N_7093,N_7065);
and U7889 (N_7889,N_7445,N_7101);
nand U7890 (N_7890,N_7065,N_7186);
nand U7891 (N_7891,N_6910,N_6848);
and U7892 (N_7892,N_7397,N_6795);
or U7893 (N_7893,N_7195,N_7488);
and U7894 (N_7894,N_7244,N_6780);
and U7895 (N_7895,N_6880,N_7495);
nand U7896 (N_7896,N_7178,N_7208);
and U7897 (N_7897,N_7046,N_7364);
or U7898 (N_7898,N_7332,N_7313);
nor U7899 (N_7899,N_7018,N_6949);
nor U7900 (N_7900,N_6779,N_7302);
xor U7901 (N_7901,N_6762,N_6920);
nand U7902 (N_7902,N_7260,N_6765);
nor U7903 (N_7903,N_7134,N_7283);
xor U7904 (N_7904,N_6771,N_7258);
or U7905 (N_7905,N_7285,N_7381);
nor U7906 (N_7906,N_7131,N_7084);
nor U7907 (N_7907,N_7152,N_7226);
nor U7908 (N_7908,N_6950,N_7341);
and U7909 (N_7909,N_7471,N_7200);
nor U7910 (N_7910,N_7374,N_7177);
nor U7911 (N_7911,N_6845,N_7219);
nand U7912 (N_7912,N_7074,N_7312);
nor U7913 (N_7913,N_6887,N_7166);
xor U7914 (N_7914,N_6925,N_6787);
nand U7915 (N_7915,N_7112,N_7437);
nor U7916 (N_7916,N_7408,N_6994);
and U7917 (N_7917,N_7107,N_6953);
nand U7918 (N_7918,N_7112,N_6887);
nor U7919 (N_7919,N_7101,N_7209);
or U7920 (N_7920,N_6871,N_6869);
nor U7921 (N_7921,N_7318,N_6942);
nor U7922 (N_7922,N_7389,N_7086);
nand U7923 (N_7923,N_7200,N_6900);
nor U7924 (N_7924,N_7208,N_6905);
xnor U7925 (N_7925,N_6750,N_7443);
or U7926 (N_7926,N_7275,N_7362);
nand U7927 (N_7927,N_7217,N_7400);
nand U7928 (N_7928,N_7423,N_7107);
and U7929 (N_7929,N_7237,N_6969);
xnor U7930 (N_7930,N_7043,N_7028);
nor U7931 (N_7931,N_7451,N_7492);
or U7932 (N_7932,N_7002,N_6948);
nor U7933 (N_7933,N_7497,N_7180);
and U7934 (N_7934,N_7438,N_7214);
nor U7935 (N_7935,N_7494,N_7413);
nor U7936 (N_7936,N_7001,N_7431);
xnor U7937 (N_7937,N_6925,N_7082);
nand U7938 (N_7938,N_6777,N_7201);
and U7939 (N_7939,N_7409,N_7374);
nor U7940 (N_7940,N_7492,N_7207);
nor U7941 (N_7941,N_7059,N_7226);
nor U7942 (N_7942,N_6780,N_6896);
or U7943 (N_7943,N_7491,N_7326);
and U7944 (N_7944,N_7054,N_7494);
nand U7945 (N_7945,N_7087,N_7492);
or U7946 (N_7946,N_7267,N_7291);
and U7947 (N_7947,N_6939,N_7347);
nand U7948 (N_7948,N_6950,N_7125);
and U7949 (N_7949,N_7138,N_7153);
or U7950 (N_7950,N_6957,N_6788);
or U7951 (N_7951,N_6866,N_6965);
nor U7952 (N_7952,N_7377,N_7292);
and U7953 (N_7953,N_6792,N_7078);
xor U7954 (N_7954,N_7280,N_6830);
and U7955 (N_7955,N_6899,N_7040);
or U7956 (N_7956,N_7295,N_7192);
nor U7957 (N_7957,N_7131,N_7259);
nand U7958 (N_7958,N_6876,N_6778);
nor U7959 (N_7959,N_7145,N_7081);
xnor U7960 (N_7960,N_7406,N_7165);
and U7961 (N_7961,N_7484,N_6828);
nor U7962 (N_7962,N_7214,N_6858);
or U7963 (N_7963,N_7204,N_6869);
xnor U7964 (N_7964,N_7481,N_7378);
nand U7965 (N_7965,N_6999,N_7452);
or U7966 (N_7966,N_7079,N_7288);
nor U7967 (N_7967,N_7090,N_7185);
nand U7968 (N_7968,N_7411,N_7331);
or U7969 (N_7969,N_7321,N_7268);
or U7970 (N_7970,N_6948,N_6894);
or U7971 (N_7971,N_7142,N_6959);
or U7972 (N_7972,N_7434,N_7181);
and U7973 (N_7973,N_6796,N_7159);
and U7974 (N_7974,N_6783,N_6894);
nand U7975 (N_7975,N_7488,N_7016);
nor U7976 (N_7976,N_7300,N_7434);
nor U7977 (N_7977,N_6964,N_7132);
and U7978 (N_7978,N_7260,N_7420);
xor U7979 (N_7979,N_7315,N_7131);
nor U7980 (N_7980,N_6814,N_7361);
and U7981 (N_7981,N_7158,N_7287);
nor U7982 (N_7982,N_7030,N_6757);
xor U7983 (N_7983,N_7125,N_7224);
and U7984 (N_7984,N_7461,N_7157);
nand U7985 (N_7985,N_6850,N_6917);
nand U7986 (N_7986,N_7352,N_7059);
nor U7987 (N_7987,N_7021,N_6878);
nand U7988 (N_7988,N_7273,N_6872);
nor U7989 (N_7989,N_7226,N_7189);
xor U7990 (N_7990,N_6900,N_7419);
nor U7991 (N_7991,N_7279,N_7329);
nor U7992 (N_7992,N_7485,N_6866);
and U7993 (N_7993,N_7365,N_7306);
or U7994 (N_7994,N_6776,N_7304);
or U7995 (N_7995,N_7138,N_6994);
and U7996 (N_7996,N_7037,N_6881);
nor U7997 (N_7997,N_6984,N_6793);
xnor U7998 (N_7998,N_6861,N_6827);
xnor U7999 (N_7999,N_6952,N_7320);
or U8000 (N_8000,N_6843,N_7401);
or U8001 (N_8001,N_7088,N_7235);
nor U8002 (N_8002,N_7459,N_7227);
and U8003 (N_8003,N_7332,N_7464);
and U8004 (N_8004,N_6990,N_7354);
nand U8005 (N_8005,N_6929,N_6974);
and U8006 (N_8006,N_7202,N_6773);
or U8007 (N_8007,N_7073,N_7374);
nand U8008 (N_8008,N_7134,N_7246);
and U8009 (N_8009,N_7177,N_6834);
and U8010 (N_8010,N_7499,N_7191);
or U8011 (N_8011,N_7001,N_7472);
nor U8012 (N_8012,N_6856,N_6795);
nand U8013 (N_8013,N_7135,N_7072);
xnor U8014 (N_8014,N_6846,N_6968);
nand U8015 (N_8015,N_7148,N_6836);
or U8016 (N_8016,N_7450,N_6957);
or U8017 (N_8017,N_6810,N_7053);
nand U8018 (N_8018,N_7381,N_6974);
nand U8019 (N_8019,N_7125,N_7330);
nand U8020 (N_8020,N_7298,N_7268);
and U8021 (N_8021,N_7326,N_6989);
or U8022 (N_8022,N_7120,N_6768);
and U8023 (N_8023,N_7347,N_6930);
and U8024 (N_8024,N_7069,N_7402);
or U8025 (N_8025,N_7093,N_6914);
xor U8026 (N_8026,N_6944,N_7398);
or U8027 (N_8027,N_7338,N_7221);
nand U8028 (N_8028,N_6981,N_7336);
and U8029 (N_8029,N_6764,N_7256);
or U8030 (N_8030,N_7175,N_7024);
nand U8031 (N_8031,N_7218,N_7460);
nand U8032 (N_8032,N_6868,N_6777);
or U8033 (N_8033,N_6877,N_7334);
xor U8034 (N_8034,N_7473,N_7052);
or U8035 (N_8035,N_7120,N_7277);
and U8036 (N_8036,N_7323,N_7242);
or U8037 (N_8037,N_6833,N_7286);
or U8038 (N_8038,N_7356,N_6769);
nand U8039 (N_8039,N_7089,N_6784);
or U8040 (N_8040,N_7351,N_6853);
nor U8041 (N_8041,N_6961,N_7120);
or U8042 (N_8042,N_7442,N_7414);
nor U8043 (N_8043,N_7472,N_7168);
nor U8044 (N_8044,N_7483,N_6827);
nand U8045 (N_8045,N_7326,N_6981);
nand U8046 (N_8046,N_7364,N_7117);
and U8047 (N_8047,N_7446,N_7396);
nor U8048 (N_8048,N_7374,N_6960);
nand U8049 (N_8049,N_7051,N_7270);
xor U8050 (N_8050,N_7287,N_6977);
and U8051 (N_8051,N_7295,N_7254);
xor U8052 (N_8052,N_7268,N_6849);
and U8053 (N_8053,N_6764,N_6826);
or U8054 (N_8054,N_7341,N_7486);
or U8055 (N_8055,N_6989,N_7479);
nor U8056 (N_8056,N_6809,N_6894);
and U8057 (N_8057,N_7242,N_7341);
and U8058 (N_8058,N_7061,N_7146);
nor U8059 (N_8059,N_7303,N_7232);
nor U8060 (N_8060,N_7438,N_6875);
nor U8061 (N_8061,N_7086,N_6968);
nand U8062 (N_8062,N_7320,N_6818);
or U8063 (N_8063,N_6790,N_7258);
and U8064 (N_8064,N_7046,N_7378);
or U8065 (N_8065,N_7438,N_7039);
or U8066 (N_8066,N_7252,N_7449);
or U8067 (N_8067,N_7037,N_6924);
and U8068 (N_8068,N_7450,N_7279);
nand U8069 (N_8069,N_7160,N_7336);
or U8070 (N_8070,N_6979,N_6797);
nand U8071 (N_8071,N_6847,N_7408);
or U8072 (N_8072,N_7430,N_7481);
nor U8073 (N_8073,N_6887,N_6975);
or U8074 (N_8074,N_7188,N_6941);
xnor U8075 (N_8075,N_6823,N_6766);
and U8076 (N_8076,N_6971,N_7492);
nor U8077 (N_8077,N_7454,N_6762);
nor U8078 (N_8078,N_7338,N_7038);
nand U8079 (N_8079,N_7463,N_6972);
nand U8080 (N_8080,N_7326,N_6973);
or U8081 (N_8081,N_7423,N_6977);
and U8082 (N_8082,N_6809,N_6838);
nor U8083 (N_8083,N_7056,N_6813);
or U8084 (N_8084,N_7254,N_7123);
nand U8085 (N_8085,N_7437,N_7070);
or U8086 (N_8086,N_6887,N_6982);
nor U8087 (N_8087,N_6781,N_7070);
or U8088 (N_8088,N_7481,N_7450);
nand U8089 (N_8089,N_6965,N_7289);
or U8090 (N_8090,N_7309,N_7431);
nand U8091 (N_8091,N_7487,N_6798);
or U8092 (N_8092,N_7280,N_6844);
xnor U8093 (N_8093,N_7117,N_7059);
and U8094 (N_8094,N_6818,N_7222);
nand U8095 (N_8095,N_7118,N_7284);
nor U8096 (N_8096,N_7327,N_6855);
nor U8097 (N_8097,N_6959,N_6867);
xor U8098 (N_8098,N_7310,N_7152);
and U8099 (N_8099,N_7066,N_7256);
nand U8100 (N_8100,N_6976,N_6815);
or U8101 (N_8101,N_7218,N_7354);
and U8102 (N_8102,N_7166,N_7087);
and U8103 (N_8103,N_7084,N_6961);
nand U8104 (N_8104,N_7145,N_6938);
or U8105 (N_8105,N_7467,N_6946);
nor U8106 (N_8106,N_7068,N_6828);
nand U8107 (N_8107,N_6799,N_6975);
or U8108 (N_8108,N_6963,N_7010);
and U8109 (N_8109,N_7420,N_7451);
or U8110 (N_8110,N_6800,N_7128);
and U8111 (N_8111,N_6883,N_7089);
nor U8112 (N_8112,N_7362,N_6972);
xnor U8113 (N_8113,N_7226,N_7384);
nor U8114 (N_8114,N_7212,N_7308);
or U8115 (N_8115,N_6963,N_6780);
or U8116 (N_8116,N_6775,N_7421);
and U8117 (N_8117,N_7464,N_7457);
or U8118 (N_8118,N_7262,N_7313);
nor U8119 (N_8119,N_6812,N_7376);
nand U8120 (N_8120,N_7497,N_7340);
or U8121 (N_8121,N_7396,N_6808);
or U8122 (N_8122,N_7011,N_7487);
nor U8123 (N_8123,N_7033,N_7211);
and U8124 (N_8124,N_6940,N_6759);
or U8125 (N_8125,N_7457,N_6811);
nand U8126 (N_8126,N_7114,N_6763);
nand U8127 (N_8127,N_7178,N_7498);
and U8128 (N_8128,N_6906,N_7270);
nand U8129 (N_8129,N_6797,N_6938);
or U8130 (N_8130,N_7058,N_7334);
nand U8131 (N_8131,N_7194,N_7120);
xnor U8132 (N_8132,N_6991,N_7355);
xnor U8133 (N_8133,N_6855,N_7378);
or U8134 (N_8134,N_6941,N_7121);
and U8135 (N_8135,N_6792,N_7390);
or U8136 (N_8136,N_7137,N_7314);
and U8137 (N_8137,N_7293,N_7330);
or U8138 (N_8138,N_6791,N_6857);
xor U8139 (N_8139,N_7459,N_7312);
or U8140 (N_8140,N_6936,N_6975);
or U8141 (N_8141,N_7311,N_6904);
and U8142 (N_8142,N_7427,N_7245);
xor U8143 (N_8143,N_7317,N_7074);
nor U8144 (N_8144,N_7034,N_6760);
nor U8145 (N_8145,N_6808,N_7020);
nand U8146 (N_8146,N_7277,N_7011);
nor U8147 (N_8147,N_6963,N_6967);
nand U8148 (N_8148,N_7289,N_7084);
xor U8149 (N_8149,N_6976,N_7044);
xnor U8150 (N_8150,N_7398,N_7140);
nor U8151 (N_8151,N_7213,N_7217);
nor U8152 (N_8152,N_6949,N_6940);
nand U8153 (N_8153,N_6950,N_6804);
nor U8154 (N_8154,N_7347,N_6836);
or U8155 (N_8155,N_6761,N_6817);
or U8156 (N_8156,N_6848,N_7186);
nor U8157 (N_8157,N_7479,N_7372);
xnor U8158 (N_8158,N_7341,N_7179);
nor U8159 (N_8159,N_6822,N_6932);
and U8160 (N_8160,N_6778,N_7053);
xor U8161 (N_8161,N_7331,N_6941);
and U8162 (N_8162,N_7019,N_7014);
nor U8163 (N_8163,N_7266,N_7241);
nand U8164 (N_8164,N_7413,N_6923);
and U8165 (N_8165,N_6787,N_7196);
nand U8166 (N_8166,N_7245,N_7485);
nand U8167 (N_8167,N_7203,N_7146);
and U8168 (N_8168,N_6886,N_7030);
nor U8169 (N_8169,N_6815,N_7131);
and U8170 (N_8170,N_7301,N_7200);
and U8171 (N_8171,N_6751,N_7328);
or U8172 (N_8172,N_7310,N_6965);
and U8173 (N_8173,N_6774,N_7231);
nand U8174 (N_8174,N_7138,N_6851);
and U8175 (N_8175,N_7122,N_6944);
and U8176 (N_8176,N_7391,N_7193);
or U8177 (N_8177,N_7367,N_7060);
or U8178 (N_8178,N_7365,N_7130);
and U8179 (N_8179,N_6931,N_6965);
and U8180 (N_8180,N_7486,N_7403);
or U8181 (N_8181,N_7402,N_6902);
and U8182 (N_8182,N_6914,N_7425);
nor U8183 (N_8183,N_6778,N_7279);
and U8184 (N_8184,N_7314,N_7007);
and U8185 (N_8185,N_7038,N_7283);
nand U8186 (N_8186,N_7262,N_7026);
xnor U8187 (N_8187,N_7254,N_6928);
and U8188 (N_8188,N_7273,N_6818);
nand U8189 (N_8189,N_7378,N_7035);
xnor U8190 (N_8190,N_7025,N_6913);
nor U8191 (N_8191,N_7247,N_7086);
or U8192 (N_8192,N_7067,N_6986);
nand U8193 (N_8193,N_7039,N_6969);
nand U8194 (N_8194,N_6758,N_6938);
and U8195 (N_8195,N_7472,N_7287);
and U8196 (N_8196,N_7038,N_7468);
and U8197 (N_8197,N_7359,N_7328);
and U8198 (N_8198,N_7071,N_6816);
nand U8199 (N_8199,N_7451,N_6826);
and U8200 (N_8200,N_6988,N_7254);
nand U8201 (N_8201,N_7114,N_7147);
and U8202 (N_8202,N_7353,N_7262);
nand U8203 (N_8203,N_7467,N_7470);
nand U8204 (N_8204,N_6988,N_7318);
or U8205 (N_8205,N_7351,N_7296);
or U8206 (N_8206,N_7401,N_6760);
nor U8207 (N_8207,N_6763,N_7395);
nand U8208 (N_8208,N_6861,N_6894);
nor U8209 (N_8209,N_6979,N_7308);
xor U8210 (N_8210,N_6885,N_6859);
nor U8211 (N_8211,N_7156,N_7379);
or U8212 (N_8212,N_6883,N_6866);
and U8213 (N_8213,N_7388,N_6901);
or U8214 (N_8214,N_6769,N_7498);
nand U8215 (N_8215,N_7495,N_6968);
or U8216 (N_8216,N_7133,N_7169);
nand U8217 (N_8217,N_7361,N_7077);
or U8218 (N_8218,N_7180,N_6839);
nor U8219 (N_8219,N_7286,N_6966);
or U8220 (N_8220,N_7248,N_7072);
and U8221 (N_8221,N_6971,N_7353);
nand U8222 (N_8222,N_6755,N_7160);
and U8223 (N_8223,N_6912,N_7082);
nor U8224 (N_8224,N_7210,N_6823);
or U8225 (N_8225,N_7469,N_7242);
and U8226 (N_8226,N_6753,N_7449);
nand U8227 (N_8227,N_6809,N_6815);
nand U8228 (N_8228,N_6904,N_7349);
xnor U8229 (N_8229,N_6980,N_6829);
and U8230 (N_8230,N_6874,N_7398);
nor U8231 (N_8231,N_7347,N_7301);
nor U8232 (N_8232,N_7178,N_7407);
nor U8233 (N_8233,N_6760,N_7063);
nand U8234 (N_8234,N_7387,N_7302);
nor U8235 (N_8235,N_7241,N_7098);
xor U8236 (N_8236,N_6891,N_7234);
nor U8237 (N_8237,N_7062,N_6769);
xnor U8238 (N_8238,N_6793,N_7391);
or U8239 (N_8239,N_7145,N_6939);
or U8240 (N_8240,N_6937,N_7089);
or U8241 (N_8241,N_6986,N_7046);
and U8242 (N_8242,N_6944,N_6786);
and U8243 (N_8243,N_7139,N_7408);
or U8244 (N_8244,N_7390,N_7421);
nor U8245 (N_8245,N_7475,N_6846);
nor U8246 (N_8246,N_7259,N_7120);
nand U8247 (N_8247,N_7237,N_7395);
nand U8248 (N_8248,N_7236,N_7047);
and U8249 (N_8249,N_7145,N_6838);
and U8250 (N_8250,N_8046,N_8058);
xor U8251 (N_8251,N_8123,N_7881);
nor U8252 (N_8252,N_7557,N_7984);
or U8253 (N_8253,N_7636,N_8141);
and U8254 (N_8254,N_7656,N_8009);
or U8255 (N_8255,N_8179,N_7589);
or U8256 (N_8256,N_8202,N_8011);
or U8257 (N_8257,N_7781,N_7552);
and U8258 (N_8258,N_7555,N_7757);
nand U8259 (N_8259,N_7564,N_7987);
xor U8260 (N_8260,N_7538,N_8002);
and U8261 (N_8261,N_7504,N_7872);
nor U8262 (N_8262,N_7730,N_7674);
and U8263 (N_8263,N_8027,N_7959);
and U8264 (N_8264,N_7698,N_7767);
or U8265 (N_8265,N_8135,N_7820);
or U8266 (N_8266,N_7610,N_7775);
or U8267 (N_8267,N_7944,N_8216);
and U8268 (N_8268,N_8186,N_7653);
xnor U8269 (N_8269,N_7854,N_8088);
xnor U8270 (N_8270,N_7714,N_7624);
nor U8271 (N_8271,N_7956,N_7704);
or U8272 (N_8272,N_7793,N_7533);
nor U8273 (N_8273,N_7584,N_7873);
nor U8274 (N_8274,N_7623,N_7889);
nor U8275 (N_8275,N_7751,N_7599);
and U8276 (N_8276,N_8114,N_7553);
or U8277 (N_8277,N_7921,N_7967);
and U8278 (N_8278,N_7927,N_7539);
or U8279 (N_8279,N_8144,N_7885);
and U8280 (N_8280,N_7541,N_8020);
nor U8281 (N_8281,N_7819,N_8134);
and U8282 (N_8282,N_7996,N_8077);
and U8283 (N_8283,N_8013,N_7681);
and U8284 (N_8284,N_7783,N_7619);
nor U8285 (N_8285,N_7855,N_8143);
xnor U8286 (N_8286,N_7894,N_7990);
nand U8287 (N_8287,N_7567,N_7663);
nor U8288 (N_8288,N_7722,N_8070);
nand U8289 (N_8289,N_7680,N_7766);
nand U8290 (N_8290,N_8197,N_7771);
and U8291 (N_8291,N_7926,N_7932);
and U8292 (N_8292,N_8040,N_7897);
and U8293 (N_8293,N_7871,N_7705);
xnor U8294 (N_8294,N_7596,N_8075);
nor U8295 (N_8295,N_7514,N_7842);
nand U8296 (N_8296,N_7887,N_7969);
nor U8297 (N_8297,N_7856,N_7699);
xor U8298 (N_8298,N_7831,N_7510);
nor U8299 (N_8299,N_7579,N_7594);
or U8300 (N_8300,N_7601,N_7840);
or U8301 (N_8301,N_8231,N_7817);
nand U8302 (N_8302,N_8066,N_8158);
and U8303 (N_8303,N_8124,N_7867);
and U8304 (N_8304,N_7938,N_8110);
or U8305 (N_8305,N_8049,N_7665);
nand U8306 (N_8306,N_7878,N_8122);
or U8307 (N_8307,N_7675,N_7554);
or U8308 (N_8308,N_7968,N_8223);
nand U8309 (N_8309,N_8029,N_8157);
nor U8310 (N_8310,N_7837,N_7958);
and U8311 (N_8311,N_7648,N_8015);
xor U8312 (N_8312,N_7587,N_8248);
and U8313 (N_8313,N_7655,N_7522);
nand U8314 (N_8314,N_7506,N_7687);
nor U8315 (N_8315,N_8221,N_7558);
and U8316 (N_8316,N_7691,N_7773);
nor U8317 (N_8317,N_7768,N_7518);
nand U8318 (N_8318,N_8208,N_7795);
nor U8319 (N_8319,N_7641,N_7616);
and U8320 (N_8320,N_7975,N_8206);
nor U8321 (N_8321,N_7772,N_7642);
and U8322 (N_8322,N_7713,N_7947);
or U8323 (N_8323,N_7633,N_8025);
and U8324 (N_8324,N_7791,N_7798);
nand U8325 (N_8325,N_8104,N_8005);
xor U8326 (N_8326,N_8083,N_7801);
and U8327 (N_8327,N_7891,N_8230);
nor U8328 (N_8328,N_8021,N_8160);
xor U8329 (N_8329,N_7779,N_7563);
and U8330 (N_8330,N_7852,N_7622);
nand U8331 (N_8331,N_8125,N_8050);
nand U8332 (N_8332,N_8218,N_8003);
nand U8333 (N_8333,N_8149,N_8076);
nor U8334 (N_8334,N_8051,N_8116);
nand U8335 (N_8335,N_8026,N_7754);
or U8336 (N_8336,N_8128,N_8138);
and U8337 (N_8337,N_7529,N_7832);
and U8338 (N_8338,N_8156,N_7924);
and U8339 (N_8339,N_7738,N_8227);
and U8340 (N_8340,N_7809,N_8220);
nor U8341 (N_8341,N_8081,N_7915);
or U8342 (N_8342,N_8080,N_7708);
and U8343 (N_8343,N_7937,N_8209);
nand U8344 (N_8344,N_7950,N_8101);
nand U8345 (N_8345,N_8213,N_7526);
xor U8346 (N_8346,N_7803,N_7581);
or U8347 (N_8347,N_8071,N_7933);
or U8348 (N_8348,N_8243,N_7695);
xnor U8349 (N_8349,N_8217,N_7918);
xor U8350 (N_8350,N_7976,N_7569);
xnor U8351 (N_8351,N_8033,N_7711);
or U8352 (N_8352,N_7764,N_7718);
and U8353 (N_8353,N_7753,N_8224);
and U8354 (N_8354,N_7978,N_7945);
nor U8355 (N_8355,N_8096,N_7732);
or U8356 (N_8356,N_7672,N_7605);
nand U8357 (N_8357,N_7707,N_7870);
nor U8358 (N_8358,N_7902,N_8182);
xor U8359 (N_8359,N_7841,N_7979);
xor U8360 (N_8360,N_7865,N_8048);
or U8361 (N_8361,N_7570,N_8131);
or U8362 (N_8362,N_7759,N_7621);
and U8363 (N_8363,N_8043,N_8226);
nor U8364 (N_8364,N_8140,N_7515);
and U8365 (N_8365,N_7828,N_8107);
or U8366 (N_8366,N_8247,N_7527);
xnor U8367 (N_8367,N_8152,N_7556);
xnor U8368 (N_8368,N_7661,N_8205);
and U8369 (N_8369,N_7747,N_7729);
and U8370 (N_8370,N_8103,N_7728);
and U8371 (N_8371,N_7760,N_7613);
or U8372 (N_8372,N_7940,N_7580);
xnor U8373 (N_8373,N_8161,N_8063);
xnor U8374 (N_8374,N_8094,N_7907);
nor U8375 (N_8375,N_7964,N_8053);
or U8376 (N_8376,N_7849,N_7574);
nor U8377 (N_8377,N_8000,N_8185);
or U8378 (N_8378,N_8065,N_7544);
nor U8379 (N_8379,N_7784,N_7762);
or U8380 (N_8380,N_7995,N_7628);
nor U8381 (N_8381,N_7774,N_7758);
nor U8382 (N_8382,N_7678,N_7890);
nor U8383 (N_8383,N_7998,N_7943);
nand U8384 (N_8384,N_7649,N_7516);
and U8385 (N_8385,N_8069,N_7595);
nor U8386 (N_8386,N_7548,N_7612);
nand U8387 (N_8387,N_8201,N_7863);
nand U8388 (N_8388,N_7954,N_8031);
or U8389 (N_8389,N_7712,N_8064);
xor U8390 (N_8390,N_7919,N_7805);
or U8391 (N_8391,N_8042,N_8052);
xnor U8392 (N_8392,N_7833,N_7733);
and U8393 (N_8393,N_7765,N_7573);
or U8394 (N_8394,N_8191,N_7512);
and U8395 (N_8395,N_8057,N_7866);
and U8396 (N_8396,N_7814,N_8242);
and U8397 (N_8397,N_7788,N_7972);
nor U8398 (N_8398,N_7593,N_7912);
and U8399 (N_8399,N_7720,N_7668);
and U8400 (N_8400,N_7647,N_7503);
or U8401 (N_8401,N_7960,N_8097);
and U8402 (N_8402,N_7607,N_7934);
nand U8403 (N_8403,N_8087,N_7966);
nand U8404 (N_8404,N_7716,N_8199);
nor U8405 (N_8405,N_8060,N_8079);
or U8406 (N_8406,N_7789,N_8045);
nand U8407 (N_8407,N_7845,N_7688);
nand U8408 (N_8408,N_7869,N_8006);
xor U8409 (N_8409,N_7682,N_8238);
and U8410 (N_8410,N_7710,N_8115);
and U8411 (N_8411,N_7726,N_8095);
nand U8412 (N_8412,N_7614,N_7925);
and U8413 (N_8413,N_7685,N_7637);
or U8414 (N_8414,N_7723,N_7739);
nor U8415 (N_8415,N_8105,N_7715);
nor U8416 (N_8416,N_8241,N_7536);
nand U8417 (N_8417,N_7755,N_7994);
nand U8418 (N_8418,N_7741,N_7606);
nor U8419 (N_8419,N_8092,N_7982);
and U8420 (N_8420,N_7868,N_7531);
nand U8421 (N_8421,N_7756,N_7684);
nand U8422 (N_8422,N_7821,N_7929);
nand U8423 (N_8423,N_7946,N_7598);
nand U8424 (N_8424,N_7922,N_7517);
nor U8425 (N_8425,N_7550,N_8085);
and U8426 (N_8426,N_8237,N_8176);
nand U8427 (N_8427,N_7876,N_8139);
or U8428 (N_8428,N_7701,N_8084);
xor U8429 (N_8429,N_7737,N_7794);
or U8430 (N_8430,N_7540,N_7836);
nand U8431 (N_8431,N_7640,N_8038);
nor U8432 (N_8432,N_7689,N_7903);
nor U8433 (N_8433,N_8056,N_7963);
nand U8434 (N_8434,N_7901,N_7886);
xor U8435 (N_8435,N_7991,N_7585);
nor U8436 (N_8436,N_7635,N_7879);
and U8437 (N_8437,N_7900,N_7931);
nand U8438 (N_8438,N_7740,N_8165);
nand U8439 (N_8439,N_7534,N_8137);
or U8440 (N_8440,N_7654,N_7939);
nor U8441 (N_8441,N_7874,N_8155);
or U8442 (N_8442,N_7559,N_7860);
nand U8443 (N_8443,N_8181,N_8246);
nand U8444 (N_8444,N_8148,N_7692);
nor U8445 (N_8445,N_8166,N_7898);
or U8446 (N_8446,N_8136,N_7683);
nor U8447 (N_8447,N_8187,N_8012);
nand U8448 (N_8448,N_7858,N_7965);
nor U8449 (N_8449,N_8229,N_8178);
and U8450 (N_8450,N_7914,N_8037);
and U8451 (N_8451,N_7864,N_8034);
and U8452 (N_8452,N_7706,N_7571);
xor U8453 (N_8453,N_7752,N_7829);
and U8454 (N_8454,N_7697,N_8121);
or U8455 (N_8455,N_7952,N_7962);
nand U8456 (N_8456,N_8210,N_8059);
xnor U8457 (N_8457,N_8118,N_8112);
or U8458 (N_8458,N_8062,N_7839);
xor U8459 (N_8459,N_7799,N_8130);
or U8460 (N_8460,N_7844,N_7620);
or U8461 (N_8461,N_8102,N_7508);
nor U8462 (N_8462,N_7575,N_8041);
and U8463 (N_8463,N_7500,N_7909);
or U8464 (N_8464,N_7896,N_7851);
nand U8465 (N_8465,N_7877,N_8047);
nand U8466 (N_8466,N_7631,N_7935);
and U8467 (N_8467,N_8035,N_7778);
nor U8468 (N_8468,N_8174,N_7749);
nand U8469 (N_8469,N_7677,N_8100);
nand U8470 (N_8470,N_7744,N_8126);
nor U8471 (N_8471,N_8219,N_7746);
or U8472 (N_8472,N_8239,N_7634);
nand U8473 (N_8473,N_8108,N_7560);
nor U8474 (N_8474,N_7770,N_8163);
nand U8475 (N_8475,N_7735,N_8117);
and U8476 (N_8476,N_7660,N_8171);
or U8477 (N_8477,N_8129,N_7702);
or U8478 (N_8478,N_8189,N_7911);
and U8479 (N_8479,N_8010,N_7651);
and U8480 (N_8480,N_7818,N_7857);
nand U8481 (N_8481,N_7630,N_8222);
nand U8482 (N_8482,N_7812,N_7602);
nand U8483 (N_8483,N_8167,N_8198);
nor U8484 (N_8484,N_7615,N_7742);
nand U8485 (N_8485,N_7676,N_7736);
and U8486 (N_8486,N_7629,N_8151);
or U8487 (N_8487,N_7645,N_7673);
or U8488 (N_8488,N_7727,N_7523);
nand U8489 (N_8489,N_7505,N_7908);
and U8490 (N_8490,N_8172,N_8039);
nor U8491 (N_8491,N_8232,N_7520);
or U8492 (N_8492,N_7892,N_7731);
and U8493 (N_8493,N_7600,N_7928);
or U8494 (N_8494,N_7884,N_8196);
or U8495 (N_8495,N_7662,N_7528);
and U8496 (N_8496,N_7917,N_7748);
and U8497 (N_8497,N_7893,N_8061);
or U8498 (N_8498,N_7999,N_7882);
and U8499 (N_8499,N_8180,N_7511);
or U8500 (N_8500,N_7834,N_7690);
and U8501 (N_8501,N_7895,N_8240);
and U8502 (N_8502,N_7547,N_7566);
and U8503 (N_8503,N_7721,N_7618);
nor U8504 (N_8504,N_8036,N_8169);
nor U8505 (N_8505,N_7980,N_8098);
nor U8506 (N_8506,N_8091,N_7530);
and U8507 (N_8507,N_8120,N_7862);
nand U8508 (N_8508,N_8211,N_8200);
xnor U8509 (N_8509,N_7543,N_8132);
nand U8510 (N_8510,N_7734,N_8111);
or U8511 (N_8511,N_8195,N_7743);
nand U8512 (N_8512,N_7955,N_8228);
nor U8513 (N_8513,N_7827,N_7646);
or U8514 (N_8514,N_8067,N_8023);
nor U8515 (N_8515,N_7906,N_7804);
nor U8516 (N_8516,N_8030,N_8004);
xnor U8517 (N_8517,N_7509,N_8072);
or U8518 (N_8518,N_7830,N_8127);
and U8519 (N_8519,N_7627,N_7745);
or U8520 (N_8520,N_7502,N_7992);
and U8521 (N_8521,N_7666,N_8207);
nor U8522 (N_8522,N_8147,N_7597);
and U8523 (N_8523,N_8109,N_7923);
xnor U8524 (N_8524,N_7883,N_8212);
or U8525 (N_8525,N_7659,N_7703);
nand U8526 (N_8526,N_7810,N_7973);
nand U8527 (N_8527,N_7686,N_8204);
xnor U8528 (N_8528,N_8162,N_8008);
and U8529 (N_8529,N_7591,N_8073);
nand U8530 (N_8530,N_8089,N_7905);
or U8531 (N_8531,N_8173,N_8074);
nand U8532 (N_8532,N_7671,N_7546);
nand U8533 (N_8533,N_8183,N_7643);
or U8534 (N_8534,N_7951,N_7551);
nand U8535 (N_8535,N_7565,N_7985);
nand U8536 (N_8536,N_7658,N_7549);
nand U8537 (N_8537,N_7904,N_7709);
or U8538 (N_8538,N_8018,N_7875);
nor U8539 (N_8539,N_7850,N_8014);
and U8540 (N_8540,N_7519,N_7724);
nand U8541 (N_8541,N_7626,N_8168);
nor U8542 (N_8542,N_7604,N_8054);
or U8543 (N_8543,N_7993,N_7521);
nand U8544 (N_8544,N_7590,N_7582);
and U8545 (N_8545,N_7910,N_8153);
nor U8546 (N_8546,N_7941,N_7562);
and U8547 (N_8547,N_7761,N_8017);
and U8548 (N_8548,N_7838,N_7763);
xnor U8549 (N_8549,N_7786,N_7792);
nor U8550 (N_8550,N_8099,N_7880);
nor U8551 (N_8551,N_7670,N_7608);
nor U8552 (N_8552,N_7657,N_7561);
nor U8553 (N_8553,N_7532,N_7750);
nor U8554 (N_8554,N_7787,N_7777);
nor U8555 (N_8555,N_7669,N_7576);
or U8556 (N_8556,N_7835,N_7989);
or U8557 (N_8557,N_7785,N_7823);
or U8558 (N_8558,N_7667,N_8225);
or U8559 (N_8559,N_7578,N_7815);
and U8560 (N_8560,N_7638,N_7806);
or U8561 (N_8561,N_7816,N_8170);
and U8562 (N_8562,N_7961,N_7942);
or U8563 (N_8563,N_7679,N_7916);
nor U8564 (N_8564,N_8214,N_7513);
nand U8565 (N_8565,N_8078,N_8175);
nor U8566 (N_8566,N_7652,N_7825);
nand U8567 (N_8567,N_7577,N_7853);
nand U8568 (N_8568,N_7811,N_7800);
or U8569 (N_8569,N_7780,N_8001);
and U8570 (N_8570,N_7650,N_7501);
xor U8571 (N_8571,N_7700,N_7986);
xor U8572 (N_8572,N_7848,N_8028);
nand U8573 (N_8573,N_7797,N_8235);
nor U8574 (N_8574,N_8236,N_7936);
and U8575 (N_8575,N_8154,N_7537);
xnor U8576 (N_8576,N_7535,N_7769);
and U8577 (N_8577,N_8159,N_7953);
xor U8578 (N_8578,N_7639,N_8164);
nand U8579 (N_8579,N_7611,N_7782);
and U8580 (N_8580,N_7725,N_7644);
nand U8581 (N_8581,N_8133,N_8024);
xnor U8582 (N_8582,N_8106,N_7572);
and U8583 (N_8583,N_7957,N_8192);
nor U8584 (N_8584,N_8086,N_7822);
nand U8585 (N_8585,N_8234,N_7588);
or U8586 (N_8586,N_7861,N_7586);
nand U8587 (N_8587,N_8193,N_7949);
or U8588 (N_8588,N_7592,N_7808);
or U8589 (N_8589,N_8044,N_7997);
nor U8590 (N_8590,N_7847,N_7846);
and U8591 (N_8591,N_8068,N_8188);
nand U8592 (N_8592,N_8142,N_8119);
nand U8593 (N_8593,N_7583,N_7790);
or U8594 (N_8594,N_8249,N_8177);
or U8595 (N_8595,N_7983,N_8032);
or U8596 (N_8596,N_7948,N_7988);
or U8597 (N_8597,N_8113,N_8146);
nand U8598 (N_8598,N_8190,N_7826);
nor U8599 (N_8599,N_7920,N_8194);
nand U8600 (N_8600,N_7609,N_7507);
nand U8601 (N_8601,N_7977,N_7568);
nor U8602 (N_8602,N_7796,N_8203);
and U8603 (N_8603,N_7776,N_7632);
and U8604 (N_8604,N_7813,N_7899);
or U8605 (N_8605,N_7981,N_7524);
nand U8606 (N_8606,N_8055,N_8019);
nand U8607 (N_8607,N_7824,N_8150);
xnor U8608 (N_8608,N_7802,N_7971);
nand U8609 (N_8609,N_7603,N_8016);
nor U8610 (N_8610,N_8007,N_7694);
xnor U8611 (N_8611,N_7717,N_7859);
nor U8612 (N_8612,N_7664,N_7807);
or U8613 (N_8613,N_7696,N_7974);
nand U8614 (N_8614,N_7545,N_8145);
or U8615 (N_8615,N_7617,N_7693);
and U8616 (N_8616,N_7930,N_8082);
and U8617 (N_8617,N_7625,N_7525);
or U8618 (N_8618,N_8245,N_8093);
or U8619 (N_8619,N_7913,N_8215);
or U8620 (N_8620,N_8184,N_8090);
or U8621 (N_8621,N_7843,N_7719);
nand U8622 (N_8622,N_8233,N_7542);
nor U8623 (N_8623,N_7970,N_8244);
nor U8624 (N_8624,N_8022,N_7888);
xnor U8625 (N_8625,N_8226,N_7642);
nor U8626 (N_8626,N_7689,N_7758);
nor U8627 (N_8627,N_7624,N_7740);
nor U8628 (N_8628,N_7759,N_8213);
and U8629 (N_8629,N_8046,N_7952);
or U8630 (N_8630,N_7502,N_8193);
and U8631 (N_8631,N_8125,N_7772);
xnor U8632 (N_8632,N_7833,N_8180);
nor U8633 (N_8633,N_7692,N_7602);
and U8634 (N_8634,N_7704,N_8056);
nand U8635 (N_8635,N_7991,N_8207);
and U8636 (N_8636,N_7567,N_8165);
and U8637 (N_8637,N_8025,N_7650);
nand U8638 (N_8638,N_7906,N_7589);
or U8639 (N_8639,N_7908,N_7625);
nand U8640 (N_8640,N_7550,N_8057);
nand U8641 (N_8641,N_8222,N_7647);
nor U8642 (N_8642,N_7939,N_7761);
or U8643 (N_8643,N_7572,N_7804);
or U8644 (N_8644,N_7599,N_7715);
nand U8645 (N_8645,N_7820,N_7888);
or U8646 (N_8646,N_7537,N_8032);
and U8647 (N_8647,N_7845,N_8214);
or U8648 (N_8648,N_7761,N_7728);
nand U8649 (N_8649,N_8089,N_7568);
and U8650 (N_8650,N_7843,N_7562);
or U8651 (N_8651,N_8174,N_7788);
nand U8652 (N_8652,N_7854,N_7926);
and U8653 (N_8653,N_7829,N_7507);
or U8654 (N_8654,N_7716,N_7688);
or U8655 (N_8655,N_7720,N_7671);
nand U8656 (N_8656,N_7773,N_7959);
and U8657 (N_8657,N_8042,N_7747);
and U8658 (N_8658,N_7897,N_7601);
nor U8659 (N_8659,N_8209,N_7830);
xnor U8660 (N_8660,N_7969,N_7760);
xnor U8661 (N_8661,N_7509,N_7588);
and U8662 (N_8662,N_8166,N_7677);
nor U8663 (N_8663,N_8133,N_7521);
nand U8664 (N_8664,N_8161,N_8125);
nand U8665 (N_8665,N_8092,N_8149);
xor U8666 (N_8666,N_7876,N_7755);
and U8667 (N_8667,N_7788,N_8122);
and U8668 (N_8668,N_7595,N_7877);
nor U8669 (N_8669,N_7828,N_7954);
nand U8670 (N_8670,N_8007,N_8237);
and U8671 (N_8671,N_7513,N_7833);
or U8672 (N_8672,N_7509,N_7861);
and U8673 (N_8673,N_7936,N_7938);
nand U8674 (N_8674,N_7864,N_7699);
nor U8675 (N_8675,N_7795,N_7536);
or U8676 (N_8676,N_7869,N_7703);
nor U8677 (N_8677,N_7783,N_8237);
and U8678 (N_8678,N_8179,N_7842);
or U8679 (N_8679,N_7739,N_7710);
or U8680 (N_8680,N_7649,N_7668);
or U8681 (N_8681,N_7587,N_8028);
nand U8682 (N_8682,N_8133,N_7814);
and U8683 (N_8683,N_8109,N_7859);
xnor U8684 (N_8684,N_7623,N_8160);
nor U8685 (N_8685,N_8045,N_7930);
or U8686 (N_8686,N_7859,N_7890);
or U8687 (N_8687,N_7994,N_7613);
or U8688 (N_8688,N_8248,N_7602);
nand U8689 (N_8689,N_8210,N_7581);
nor U8690 (N_8690,N_7979,N_7708);
or U8691 (N_8691,N_7911,N_8227);
and U8692 (N_8692,N_8108,N_8179);
or U8693 (N_8693,N_7500,N_7994);
and U8694 (N_8694,N_8225,N_8061);
nor U8695 (N_8695,N_8160,N_7915);
and U8696 (N_8696,N_7591,N_7781);
or U8697 (N_8697,N_8188,N_7705);
nor U8698 (N_8698,N_7694,N_7741);
nand U8699 (N_8699,N_7901,N_7582);
and U8700 (N_8700,N_8069,N_7818);
nand U8701 (N_8701,N_8192,N_7570);
and U8702 (N_8702,N_7844,N_8009);
nor U8703 (N_8703,N_7878,N_7710);
or U8704 (N_8704,N_8078,N_8217);
and U8705 (N_8705,N_7528,N_8014);
or U8706 (N_8706,N_8006,N_7570);
nor U8707 (N_8707,N_7797,N_8166);
and U8708 (N_8708,N_8123,N_7667);
and U8709 (N_8709,N_7612,N_7752);
nor U8710 (N_8710,N_8074,N_7695);
or U8711 (N_8711,N_7719,N_7579);
xor U8712 (N_8712,N_8013,N_7725);
xnor U8713 (N_8713,N_7974,N_7724);
nand U8714 (N_8714,N_7862,N_7768);
or U8715 (N_8715,N_8147,N_7627);
nand U8716 (N_8716,N_7552,N_7656);
or U8717 (N_8717,N_7696,N_7581);
nand U8718 (N_8718,N_8228,N_8025);
nor U8719 (N_8719,N_7776,N_8199);
and U8720 (N_8720,N_8108,N_8127);
nand U8721 (N_8721,N_7595,N_7984);
xnor U8722 (N_8722,N_7909,N_8078);
and U8723 (N_8723,N_7899,N_8225);
and U8724 (N_8724,N_7793,N_8082);
nand U8725 (N_8725,N_7866,N_8179);
and U8726 (N_8726,N_7755,N_7955);
nand U8727 (N_8727,N_7554,N_8228);
nor U8728 (N_8728,N_8064,N_7512);
or U8729 (N_8729,N_8087,N_8139);
nor U8730 (N_8730,N_7897,N_7840);
nand U8731 (N_8731,N_8040,N_7700);
nor U8732 (N_8732,N_7857,N_7866);
and U8733 (N_8733,N_7719,N_8210);
nor U8734 (N_8734,N_7833,N_8086);
xnor U8735 (N_8735,N_8187,N_7724);
nand U8736 (N_8736,N_7502,N_7622);
xnor U8737 (N_8737,N_7920,N_7537);
nand U8738 (N_8738,N_7882,N_7576);
nor U8739 (N_8739,N_7881,N_7571);
and U8740 (N_8740,N_7790,N_7564);
or U8741 (N_8741,N_8174,N_8245);
or U8742 (N_8742,N_7641,N_8029);
and U8743 (N_8743,N_7841,N_8175);
xnor U8744 (N_8744,N_8037,N_7633);
nor U8745 (N_8745,N_7896,N_7945);
nand U8746 (N_8746,N_7841,N_7844);
or U8747 (N_8747,N_8093,N_7666);
or U8748 (N_8748,N_7976,N_7522);
nor U8749 (N_8749,N_7805,N_8172);
nand U8750 (N_8750,N_7954,N_7690);
nor U8751 (N_8751,N_7541,N_8230);
nand U8752 (N_8752,N_7739,N_7745);
and U8753 (N_8753,N_8175,N_7785);
or U8754 (N_8754,N_7510,N_7721);
nor U8755 (N_8755,N_8042,N_8166);
xnor U8756 (N_8756,N_7966,N_7869);
nor U8757 (N_8757,N_8054,N_7837);
nand U8758 (N_8758,N_8153,N_8145);
or U8759 (N_8759,N_7956,N_8145);
nand U8760 (N_8760,N_7736,N_8068);
or U8761 (N_8761,N_8212,N_7981);
and U8762 (N_8762,N_7957,N_7828);
nand U8763 (N_8763,N_7940,N_7826);
nor U8764 (N_8764,N_7685,N_7690);
nor U8765 (N_8765,N_8129,N_7565);
or U8766 (N_8766,N_7844,N_8171);
and U8767 (N_8767,N_7779,N_7614);
nand U8768 (N_8768,N_7929,N_8202);
or U8769 (N_8769,N_7627,N_8073);
nand U8770 (N_8770,N_7852,N_7748);
nor U8771 (N_8771,N_7835,N_7732);
nand U8772 (N_8772,N_8095,N_7562);
and U8773 (N_8773,N_7517,N_7511);
or U8774 (N_8774,N_7763,N_7774);
nand U8775 (N_8775,N_8008,N_7560);
and U8776 (N_8776,N_7558,N_7791);
or U8777 (N_8777,N_7533,N_7707);
nand U8778 (N_8778,N_8096,N_7733);
or U8779 (N_8779,N_7807,N_8245);
nand U8780 (N_8780,N_7589,N_8115);
nor U8781 (N_8781,N_8225,N_7756);
or U8782 (N_8782,N_7996,N_7516);
and U8783 (N_8783,N_7903,N_7692);
and U8784 (N_8784,N_8128,N_8223);
and U8785 (N_8785,N_7634,N_7738);
nor U8786 (N_8786,N_7632,N_8140);
or U8787 (N_8787,N_7791,N_7831);
nand U8788 (N_8788,N_8234,N_8197);
or U8789 (N_8789,N_7670,N_7535);
and U8790 (N_8790,N_8013,N_7836);
or U8791 (N_8791,N_8181,N_7569);
nand U8792 (N_8792,N_7857,N_8026);
nor U8793 (N_8793,N_7980,N_7760);
or U8794 (N_8794,N_7877,N_7947);
or U8795 (N_8795,N_7848,N_8139);
xnor U8796 (N_8796,N_7715,N_8100);
nor U8797 (N_8797,N_8035,N_7962);
and U8798 (N_8798,N_7851,N_8143);
or U8799 (N_8799,N_7982,N_7601);
nand U8800 (N_8800,N_8034,N_7704);
nor U8801 (N_8801,N_7722,N_7638);
nand U8802 (N_8802,N_7835,N_8090);
and U8803 (N_8803,N_7600,N_7733);
nand U8804 (N_8804,N_7654,N_7778);
nor U8805 (N_8805,N_8124,N_7639);
nand U8806 (N_8806,N_7898,N_7594);
xnor U8807 (N_8807,N_7555,N_8240);
and U8808 (N_8808,N_8117,N_8185);
or U8809 (N_8809,N_8002,N_7718);
nor U8810 (N_8810,N_7974,N_8048);
or U8811 (N_8811,N_8213,N_8048);
or U8812 (N_8812,N_8238,N_7987);
and U8813 (N_8813,N_7923,N_8188);
xor U8814 (N_8814,N_7902,N_7518);
or U8815 (N_8815,N_7954,N_8246);
or U8816 (N_8816,N_7510,N_7839);
nand U8817 (N_8817,N_7560,N_7924);
or U8818 (N_8818,N_8136,N_8226);
nand U8819 (N_8819,N_7954,N_7927);
and U8820 (N_8820,N_7679,N_8026);
and U8821 (N_8821,N_7672,N_8026);
or U8822 (N_8822,N_7536,N_8008);
nor U8823 (N_8823,N_7620,N_7611);
and U8824 (N_8824,N_7658,N_7714);
and U8825 (N_8825,N_8139,N_7505);
xnor U8826 (N_8826,N_7508,N_8059);
nand U8827 (N_8827,N_7749,N_8075);
xor U8828 (N_8828,N_8010,N_8075);
and U8829 (N_8829,N_7879,N_7705);
or U8830 (N_8830,N_8061,N_7614);
and U8831 (N_8831,N_7517,N_7803);
nor U8832 (N_8832,N_8189,N_8097);
nor U8833 (N_8833,N_8099,N_7698);
nor U8834 (N_8834,N_8018,N_7865);
nand U8835 (N_8835,N_7594,N_7557);
nor U8836 (N_8836,N_7671,N_7579);
nor U8837 (N_8837,N_8138,N_7745);
nor U8838 (N_8838,N_7961,N_8095);
xor U8839 (N_8839,N_7747,N_7979);
xnor U8840 (N_8840,N_8180,N_7676);
nor U8841 (N_8841,N_7768,N_7840);
and U8842 (N_8842,N_7641,N_7592);
or U8843 (N_8843,N_7525,N_7560);
nand U8844 (N_8844,N_8077,N_7937);
and U8845 (N_8845,N_7856,N_7598);
and U8846 (N_8846,N_7835,N_7570);
nor U8847 (N_8847,N_7605,N_8233);
nand U8848 (N_8848,N_7625,N_8045);
and U8849 (N_8849,N_8232,N_7672);
or U8850 (N_8850,N_7677,N_7832);
nor U8851 (N_8851,N_8239,N_7869);
nand U8852 (N_8852,N_7605,N_7970);
nand U8853 (N_8853,N_8184,N_7854);
nor U8854 (N_8854,N_7916,N_8212);
and U8855 (N_8855,N_7638,N_7974);
nor U8856 (N_8856,N_7730,N_8071);
nand U8857 (N_8857,N_8122,N_7703);
nor U8858 (N_8858,N_7956,N_8196);
and U8859 (N_8859,N_7502,N_8238);
nor U8860 (N_8860,N_7534,N_7958);
nor U8861 (N_8861,N_7555,N_8100);
and U8862 (N_8862,N_8149,N_8204);
and U8863 (N_8863,N_8229,N_7835);
nand U8864 (N_8864,N_7943,N_7994);
or U8865 (N_8865,N_7503,N_7666);
nand U8866 (N_8866,N_7658,N_7593);
nand U8867 (N_8867,N_7674,N_7890);
xor U8868 (N_8868,N_7506,N_7621);
xor U8869 (N_8869,N_7909,N_8080);
or U8870 (N_8870,N_8238,N_8210);
nor U8871 (N_8871,N_8141,N_7964);
nand U8872 (N_8872,N_7817,N_7680);
nor U8873 (N_8873,N_7600,N_8028);
and U8874 (N_8874,N_8231,N_8024);
nor U8875 (N_8875,N_7627,N_8059);
nand U8876 (N_8876,N_7888,N_7690);
and U8877 (N_8877,N_7508,N_7672);
nor U8878 (N_8878,N_7710,N_7866);
xnor U8879 (N_8879,N_7908,N_8139);
and U8880 (N_8880,N_7500,N_8073);
xor U8881 (N_8881,N_7956,N_8048);
nor U8882 (N_8882,N_8013,N_7559);
nand U8883 (N_8883,N_7678,N_7788);
nor U8884 (N_8884,N_7740,N_8042);
or U8885 (N_8885,N_8009,N_7653);
xor U8886 (N_8886,N_8177,N_7566);
xnor U8887 (N_8887,N_7641,N_7502);
nand U8888 (N_8888,N_7767,N_8236);
xor U8889 (N_8889,N_8049,N_8218);
and U8890 (N_8890,N_8193,N_8111);
nor U8891 (N_8891,N_7894,N_8221);
nand U8892 (N_8892,N_7826,N_7891);
or U8893 (N_8893,N_7865,N_7713);
nand U8894 (N_8894,N_7655,N_7567);
xnor U8895 (N_8895,N_7559,N_8115);
and U8896 (N_8896,N_8052,N_7986);
nor U8897 (N_8897,N_7853,N_7894);
or U8898 (N_8898,N_7812,N_8055);
nand U8899 (N_8899,N_7918,N_7993);
nor U8900 (N_8900,N_7991,N_7709);
and U8901 (N_8901,N_7772,N_7911);
xnor U8902 (N_8902,N_7650,N_7981);
nor U8903 (N_8903,N_7536,N_8100);
xor U8904 (N_8904,N_8220,N_7603);
nor U8905 (N_8905,N_7970,N_7869);
and U8906 (N_8906,N_7510,N_7737);
xnor U8907 (N_8907,N_7643,N_7564);
and U8908 (N_8908,N_8011,N_7917);
or U8909 (N_8909,N_7680,N_8034);
or U8910 (N_8910,N_7506,N_8071);
nand U8911 (N_8911,N_7855,N_7510);
xor U8912 (N_8912,N_8186,N_7506);
nor U8913 (N_8913,N_7669,N_7793);
and U8914 (N_8914,N_7559,N_8110);
nor U8915 (N_8915,N_7790,N_8166);
or U8916 (N_8916,N_7714,N_8053);
and U8917 (N_8917,N_7517,N_7617);
nor U8918 (N_8918,N_8051,N_8125);
xnor U8919 (N_8919,N_7707,N_7605);
and U8920 (N_8920,N_7551,N_7895);
nor U8921 (N_8921,N_7995,N_7632);
or U8922 (N_8922,N_8154,N_7586);
nand U8923 (N_8923,N_7870,N_7860);
and U8924 (N_8924,N_7860,N_7744);
nor U8925 (N_8925,N_8052,N_7714);
and U8926 (N_8926,N_8133,N_7864);
xor U8927 (N_8927,N_7850,N_7882);
xnor U8928 (N_8928,N_7880,N_7864);
or U8929 (N_8929,N_7589,N_8038);
nor U8930 (N_8930,N_7694,N_7589);
or U8931 (N_8931,N_8195,N_7979);
nor U8932 (N_8932,N_7781,N_7978);
and U8933 (N_8933,N_7882,N_7650);
nand U8934 (N_8934,N_7818,N_7996);
nor U8935 (N_8935,N_7751,N_7965);
or U8936 (N_8936,N_7889,N_8213);
xor U8937 (N_8937,N_8206,N_8004);
nor U8938 (N_8938,N_7815,N_7884);
nand U8939 (N_8939,N_8072,N_8104);
nand U8940 (N_8940,N_8226,N_7675);
or U8941 (N_8941,N_7789,N_7697);
nand U8942 (N_8942,N_7880,N_7577);
nor U8943 (N_8943,N_7829,N_8083);
and U8944 (N_8944,N_7549,N_7604);
nand U8945 (N_8945,N_7697,N_7995);
nand U8946 (N_8946,N_7543,N_8181);
xnor U8947 (N_8947,N_8011,N_7791);
or U8948 (N_8948,N_7608,N_8226);
xor U8949 (N_8949,N_7967,N_7767);
nor U8950 (N_8950,N_7991,N_8179);
xnor U8951 (N_8951,N_7952,N_7678);
xor U8952 (N_8952,N_7628,N_7740);
nor U8953 (N_8953,N_8083,N_8098);
or U8954 (N_8954,N_8037,N_7568);
and U8955 (N_8955,N_7863,N_7665);
nand U8956 (N_8956,N_7953,N_8078);
xor U8957 (N_8957,N_7787,N_7584);
and U8958 (N_8958,N_7508,N_8174);
and U8959 (N_8959,N_7647,N_7579);
and U8960 (N_8960,N_7938,N_7849);
and U8961 (N_8961,N_7582,N_7633);
or U8962 (N_8962,N_8021,N_8228);
nand U8963 (N_8963,N_7758,N_8061);
and U8964 (N_8964,N_8200,N_7619);
nor U8965 (N_8965,N_8223,N_8059);
and U8966 (N_8966,N_8217,N_7670);
or U8967 (N_8967,N_7871,N_8056);
and U8968 (N_8968,N_7557,N_7680);
nand U8969 (N_8969,N_7605,N_8228);
and U8970 (N_8970,N_7696,N_7539);
nor U8971 (N_8971,N_8067,N_8140);
xor U8972 (N_8972,N_7816,N_7872);
or U8973 (N_8973,N_7809,N_7985);
nor U8974 (N_8974,N_8183,N_7547);
and U8975 (N_8975,N_7835,N_7983);
nand U8976 (N_8976,N_8159,N_7535);
nand U8977 (N_8977,N_7521,N_8081);
and U8978 (N_8978,N_8164,N_7869);
or U8979 (N_8979,N_7677,N_7686);
or U8980 (N_8980,N_7741,N_7549);
nor U8981 (N_8981,N_7530,N_7556);
nand U8982 (N_8982,N_7669,N_7594);
nand U8983 (N_8983,N_7802,N_7926);
xnor U8984 (N_8984,N_8121,N_7625);
nand U8985 (N_8985,N_7945,N_7926);
or U8986 (N_8986,N_7527,N_7610);
and U8987 (N_8987,N_7860,N_8155);
xnor U8988 (N_8988,N_7693,N_7507);
nand U8989 (N_8989,N_8034,N_7560);
or U8990 (N_8990,N_7806,N_8206);
nand U8991 (N_8991,N_7523,N_7677);
or U8992 (N_8992,N_7797,N_7789);
nand U8993 (N_8993,N_7568,N_8233);
and U8994 (N_8994,N_7950,N_8246);
and U8995 (N_8995,N_7791,N_7954);
nand U8996 (N_8996,N_8215,N_7737);
nand U8997 (N_8997,N_7873,N_7988);
and U8998 (N_8998,N_7561,N_7880);
nor U8999 (N_8999,N_7791,N_7879);
nand U9000 (N_9000,N_8904,N_8760);
or U9001 (N_9001,N_8511,N_8629);
xnor U9002 (N_9002,N_8764,N_8360);
nand U9003 (N_9003,N_8982,N_8630);
nor U9004 (N_9004,N_8504,N_8663);
and U9005 (N_9005,N_8279,N_8495);
and U9006 (N_9006,N_8297,N_8706);
nand U9007 (N_9007,N_8774,N_8509);
nand U9008 (N_9008,N_8618,N_8428);
and U9009 (N_9009,N_8666,N_8540);
nor U9010 (N_9010,N_8841,N_8470);
nor U9011 (N_9011,N_8315,N_8259);
nor U9012 (N_9012,N_8843,N_8411);
xnor U9013 (N_9013,N_8580,N_8874);
nor U9014 (N_9014,N_8709,N_8754);
xor U9015 (N_9015,N_8672,N_8961);
nor U9016 (N_9016,N_8445,N_8976);
nor U9017 (N_9017,N_8688,N_8349);
and U9018 (N_9018,N_8742,N_8409);
nand U9019 (N_9019,N_8311,N_8788);
nand U9020 (N_9020,N_8912,N_8382);
or U9021 (N_9021,N_8680,N_8738);
xor U9022 (N_9022,N_8467,N_8925);
nand U9023 (N_9023,N_8942,N_8549);
nand U9024 (N_9024,N_8930,N_8386);
or U9025 (N_9025,N_8779,N_8269);
nand U9026 (N_9026,N_8389,N_8363);
nor U9027 (N_9027,N_8842,N_8955);
and U9028 (N_9028,N_8408,N_8547);
and U9029 (N_9029,N_8512,N_8447);
nand U9030 (N_9030,N_8572,N_8330);
nor U9031 (N_9031,N_8763,N_8271);
and U9032 (N_9032,N_8426,N_8857);
or U9033 (N_9033,N_8864,N_8953);
nor U9034 (N_9034,N_8808,N_8868);
nor U9035 (N_9035,N_8286,N_8775);
or U9036 (N_9036,N_8260,N_8883);
or U9037 (N_9037,N_8784,N_8937);
and U9038 (N_9038,N_8909,N_8451);
and U9039 (N_9039,N_8280,N_8728);
nand U9040 (N_9040,N_8635,N_8308);
nor U9041 (N_9041,N_8477,N_8807);
and U9042 (N_9042,N_8254,N_8829);
xnor U9043 (N_9043,N_8612,N_8785);
or U9044 (N_9044,N_8866,N_8673);
or U9045 (N_9045,N_8422,N_8703);
nor U9046 (N_9046,N_8812,N_8573);
nand U9047 (N_9047,N_8380,N_8402);
nor U9048 (N_9048,N_8491,N_8570);
and U9049 (N_9049,N_8561,N_8616);
or U9050 (N_9050,N_8412,N_8318);
nor U9051 (N_9051,N_8989,N_8362);
and U9052 (N_9052,N_8959,N_8285);
nand U9053 (N_9053,N_8834,N_8933);
xor U9054 (N_9054,N_8737,N_8908);
nand U9055 (N_9055,N_8610,N_8876);
nor U9056 (N_9056,N_8480,N_8585);
and U9057 (N_9057,N_8820,N_8598);
nor U9058 (N_9058,N_8861,N_8458);
and U9059 (N_9059,N_8740,N_8708);
and U9060 (N_9060,N_8916,N_8801);
or U9061 (N_9061,N_8979,N_8985);
nor U9062 (N_9062,N_8892,N_8523);
nand U9063 (N_9063,N_8867,N_8948);
nand U9064 (N_9064,N_8498,N_8981);
nand U9065 (N_9065,N_8697,N_8606);
and U9066 (N_9066,N_8965,N_8716);
nor U9067 (N_9067,N_8499,N_8323);
nor U9068 (N_9068,N_8278,N_8614);
and U9069 (N_9069,N_8443,N_8604);
nand U9070 (N_9070,N_8622,N_8678);
nand U9071 (N_9071,N_8939,N_8533);
nand U9072 (N_9072,N_8729,N_8685);
nor U9073 (N_9073,N_8488,N_8272);
or U9074 (N_9074,N_8655,N_8320);
nor U9075 (N_9075,N_8634,N_8994);
nand U9076 (N_9076,N_8682,N_8593);
nand U9077 (N_9077,N_8450,N_8823);
nor U9078 (N_9078,N_8291,N_8448);
nand U9079 (N_9079,N_8287,N_8446);
nand U9080 (N_9080,N_8795,N_8670);
nand U9081 (N_9081,N_8911,N_8759);
xor U9082 (N_9082,N_8336,N_8956);
nor U9083 (N_9083,N_8435,N_8407);
or U9084 (N_9084,N_8677,N_8684);
nor U9085 (N_9085,N_8569,N_8814);
nand U9086 (N_9086,N_8466,N_8691);
nand U9087 (N_9087,N_8800,N_8802);
and U9088 (N_9088,N_8700,N_8873);
nand U9089 (N_9089,N_8919,N_8356);
nand U9090 (N_9090,N_8437,N_8973);
nand U9091 (N_9091,N_8563,N_8299);
nor U9092 (N_9092,N_8421,N_8815);
nor U9093 (N_9093,N_8387,N_8313);
and U9094 (N_9094,N_8510,N_8300);
nor U9095 (N_9095,N_8681,N_8657);
and U9096 (N_9096,N_8350,N_8932);
nor U9097 (N_9097,N_8776,N_8649);
or U9098 (N_9098,N_8772,N_8967);
nand U9099 (N_9099,N_8340,N_8722);
nor U9100 (N_9100,N_8496,N_8791);
nor U9101 (N_9101,N_8913,N_8543);
or U9102 (N_9102,N_8717,N_8895);
or U9103 (N_9103,N_8662,N_8381);
and U9104 (N_9104,N_8970,N_8995);
and U9105 (N_9105,N_8720,N_8958);
nor U9106 (N_9106,N_8719,N_8416);
and U9107 (N_9107,N_8534,N_8661);
and U9108 (N_9108,N_8319,N_8838);
nor U9109 (N_9109,N_8565,N_8951);
nand U9110 (N_9110,N_8645,N_8264);
xor U9111 (N_9111,N_8632,N_8597);
nor U9112 (N_9112,N_8877,N_8928);
nor U9113 (N_9113,N_8332,N_8420);
or U9114 (N_9114,N_8902,N_8718);
and U9115 (N_9115,N_8705,N_8879);
xor U9116 (N_9116,N_8805,N_8993);
nand U9117 (N_9117,N_8980,N_8393);
xnor U9118 (N_9118,N_8513,N_8749);
nor U9119 (N_9119,N_8465,N_8871);
and U9120 (N_9120,N_8659,N_8701);
and U9121 (N_9121,N_8745,N_8949);
xor U9122 (N_9122,N_8463,N_8265);
nor U9123 (N_9123,N_8810,N_8564);
or U9124 (N_9124,N_8735,N_8261);
or U9125 (N_9125,N_8853,N_8743);
nand U9126 (N_9126,N_8787,N_8762);
nor U9127 (N_9127,N_8266,N_8793);
nor U9128 (N_9128,N_8858,N_8583);
nor U9129 (N_9129,N_8508,N_8650);
nand U9130 (N_9130,N_8859,N_8686);
or U9131 (N_9131,N_8438,N_8997);
or U9132 (N_9132,N_8875,N_8889);
nand U9133 (N_9133,N_8669,N_8314);
xor U9134 (N_9134,N_8817,N_8986);
nand U9135 (N_9135,N_8526,N_8256);
nor U9136 (N_9136,N_8768,N_8660);
or U9137 (N_9137,N_8777,N_8984);
xor U9138 (N_9138,N_8358,N_8436);
and U9139 (N_9139,N_8419,N_8460);
nor U9140 (N_9140,N_8490,N_8884);
and U9141 (N_9141,N_8628,N_8761);
nand U9142 (N_9142,N_8675,N_8922);
or U9143 (N_9143,N_8579,N_8766);
nor U9144 (N_9144,N_8794,N_8452);
and U9145 (N_9145,N_8298,N_8651);
or U9146 (N_9146,N_8289,N_8890);
or U9147 (N_9147,N_8501,N_8502);
xor U9148 (N_9148,N_8668,N_8975);
nand U9149 (N_9149,N_8366,N_8963);
or U9150 (N_9150,N_8770,N_8331);
xnor U9151 (N_9151,N_8600,N_8590);
nor U9152 (N_9152,N_8905,N_8252);
nor U9153 (N_9153,N_8926,N_8878);
and U9154 (N_9154,N_8489,N_8397);
or U9155 (N_9155,N_8893,N_8778);
xnor U9156 (N_9156,N_8557,N_8410);
nor U9157 (N_9157,N_8920,N_8530);
nand U9158 (N_9158,N_8957,N_8934);
nor U9159 (N_9159,N_8746,N_8797);
and U9160 (N_9160,N_8813,N_8591);
or U9161 (N_9161,N_8667,N_8636);
nand U9162 (N_9162,N_8845,N_8427);
xor U9163 (N_9163,N_8275,N_8560);
or U9164 (N_9164,N_8907,N_8918);
nor U9165 (N_9165,N_8442,N_8457);
or U9166 (N_9166,N_8255,N_8839);
xnor U9167 (N_9167,N_8505,N_8282);
nor U9168 (N_9168,N_8620,N_8702);
or U9169 (N_9169,N_8648,N_8929);
nor U9170 (N_9170,N_8977,N_8303);
and U9171 (N_9171,N_8506,N_8277);
and U9172 (N_9172,N_8587,N_8545);
nand U9173 (N_9173,N_8947,N_8444);
nor U9174 (N_9174,N_8676,N_8528);
nor U9175 (N_9175,N_8273,N_8485);
nand U9176 (N_9176,N_8824,N_8307);
nand U9177 (N_9177,N_8752,N_8609);
nand U9178 (N_9178,N_8840,N_8556);
nand U9179 (N_9179,N_8696,N_8695);
nor U9180 (N_9180,N_8576,N_8462);
and U9181 (N_9181,N_8617,N_8832);
nor U9182 (N_9182,N_8596,N_8964);
nor U9183 (N_9183,N_8941,N_8476);
xor U9184 (N_9184,N_8699,N_8479);
and U9185 (N_9185,N_8693,N_8322);
nand U9186 (N_9186,N_8773,N_8855);
or U9187 (N_9187,N_8687,N_8836);
nor U9188 (N_9188,N_8990,N_8383);
nand U9189 (N_9189,N_8268,N_8730);
nand U9190 (N_9190,N_8586,N_8992);
nor U9191 (N_9191,N_8847,N_8454);
nand U9192 (N_9192,N_8921,N_8558);
nand U9193 (N_9193,N_8423,N_8969);
nand U9194 (N_9194,N_8983,N_8581);
or U9195 (N_9195,N_8413,N_8346);
nor U9196 (N_9196,N_8370,N_8653);
and U9197 (N_9197,N_8430,N_8769);
nand U9198 (N_9198,N_8385,N_8809);
nor U9199 (N_9199,N_8333,N_8846);
nor U9200 (N_9200,N_8559,N_8848);
and U9201 (N_9201,N_8398,N_8384);
xor U9202 (N_9202,N_8747,N_8935);
nor U9203 (N_9203,N_8721,N_8999);
xnor U9204 (N_9204,N_8619,N_8455);
or U9205 (N_9205,N_8379,N_8471);
or U9206 (N_9206,N_8945,N_8732);
xor U9207 (N_9207,N_8830,N_8588);
nor U9208 (N_9208,N_8664,N_8539);
or U9209 (N_9209,N_8344,N_8689);
nand U9210 (N_9210,N_8850,N_8825);
and U9211 (N_9211,N_8414,N_8494);
and U9212 (N_9212,N_8262,N_8552);
and U9213 (N_9213,N_8365,N_8631);
and U9214 (N_9214,N_8584,N_8345);
and U9215 (N_9215,N_8492,N_8882);
xnor U9216 (N_9216,N_8253,N_8301);
or U9217 (N_9217,N_8923,N_8852);
and U9218 (N_9218,N_8734,N_8514);
xnor U9219 (N_9219,N_8633,N_8736);
xnor U9220 (N_9220,N_8903,N_8270);
nand U9221 (N_9221,N_8475,N_8373);
or U9222 (N_9222,N_8683,N_8578);
xor U9223 (N_9223,N_8627,N_8487);
nand U9224 (N_9224,N_8711,N_8723);
nor U9225 (N_9225,N_8962,N_8783);
or U9226 (N_9226,N_8364,N_8715);
and U9227 (N_9227,N_8405,N_8537);
nand U9228 (N_9228,N_8944,N_8637);
nor U9229 (N_9229,N_8910,N_8425);
xor U9230 (N_9230,N_8671,N_8731);
nor U9231 (N_9231,N_8267,N_8603);
or U9232 (N_9232,N_8522,N_8639);
or U9233 (N_9233,N_8390,N_8434);
and U9234 (N_9234,N_8404,N_8396);
and U9235 (N_9235,N_8625,N_8304);
nor U9236 (N_9236,N_8656,N_8707);
and U9237 (N_9237,N_8520,N_8283);
nand U9238 (N_9238,N_8251,N_8726);
or U9239 (N_9239,N_8592,N_8357);
nor U9240 (N_9240,N_8595,N_8615);
and U9241 (N_9241,N_8865,N_8546);
and U9242 (N_9242,N_8521,N_8541);
or U9243 (N_9243,N_8833,N_8429);
or U9244 (N_9244,N_8374,N_8439);
xnor U9245 (N_9245,N_8854,N_8258);
and U9246 (N_9246,N_8361,N_8453);
nand U9247 (N_9247,N_8863,N_8325);
or U9248 (N_9248,N_8647,N_8324);
nand U9249 (N_9249,N_8359,N_8611);
or U9250 (N_9250,N_8607,N_8601);
nor U9251 (N_9251,N_8338,N_8638);
xnor U9252 (N_9252,N_8862,N_8869);
nand U9253 (N_9253,N_8594,N_8341);
nor U9254 (N_9254,N_8765,N_8792);
nand U9255 (N_9255,N_8885,N_8403);
nand U9256 (N_9256,N_8621,N_8901);
and U9257 (N_9257,N_8417,N_8551);
or U9258 (N_9258,N_8725,N_8469);
and U9259 (N_9259,N_8544,N_8449);
nand U9260 (N_9260,N_8288,N_8328);
xnor U9261 (N_9261,N_8555,N_8658);
nor U9262 (N_9262,N_8987,N_8767);
xnor U9263 (N_9263,N_8294,N_8566);
or U9264 (N_9264,N_8516,N_8899);
nor U9265 (N_9265,N_8310,N_8727);
and U9266 (N_9266,N_8713,N_8828);
nor U9267 (N_9267,N_8468,N_8352);
nand U9268 (N_9268,N_8507,N_8654);
nand U9269 (N_9269,N_8527,N_8623);
nor U9270 (N_9270,N_8844,N_8679);
nand U9271 (N_9271,N_8582,N_8938);
nand U9272 (N_9272,N_8827,N_8860);
xor U9273 (N_9273,N_8991,N_8394);
nand U9274 (N_9274,N_8900,N_8851);
and U9275 (N_9275,N_8602,N_8296);
or U9276 (N_9276,N_8305,N_8837);
xor U9277 (N_9277,N_8295,N_8940);
and U9278 (N_9278,N_8531,N_8281);
nor U9279 (N_9279,N_8898,N_8372);
xnor U9280 (N_9280,N_8757,N_8665);
nor U9281 (N_9281,N_8309,N_8816);
or U9282 (N_9282,N_8724,N_8326);
or U9283 (N_9283,N_8881,N_8532);
or U9284 (N_9284,N_8971,N_8302);
xor U9285 (N_9285,N_8355,N_8486);
and U9286 (N_9286,N_8811,N_8339);
or U9287 (N_9287,N_8642,N_8712);
nand U9288 (N_9288,N_8433,N_8401);
or U9289 (N_9289,N_8376,N_8478);
nand U9290 (N_9290,N_8400,N_8978);
nor U9291 (N_9291,N_8798,N_8589);
or U9292 (N_9292,N_8367,N_8274);
nor U9293 (N_9293,N_8914,N_8782);
nor U9294 (N_9294,N_8368,N_8574);
or U9295 (N_9295,N_8786,N_8529);
and U9296 (N_9296,N_8316,N_8554);
xnor U9297 (N_9297,N_8756,N_8431);
or U9298 (N_9298,N_8826,N_8497);
and U9299 (N_9299,N_8406,N_8950);
nand U9300 (N_9300,N_8896,N_8870);
nand U9301 (N_9301,N_8790,N_8263);
nand U9302 (N_9302,N_8996,N_8392);
or U9303 (N_9303,N_8250,N_8484);
nand U9304 (N_9304,N_8388,N_8348);
xor U9305 (N_9305,N_8542,N_8714);
and U9306 (N_9306,N_8375,N_8988);
or U9307 (N_9307,N_8456,N_8292);
nand U9308 (N_9308,N_8652,N_8399);
nor U9309 (N_9309,N_8440,N_8891);
nor U9310 (N_9310,N_8329,N_8536);
and U9311 (N_9311,N_8796,N_8966);
nor U9312 (N_9312,N_8519,N_8644);
nand U9313 (N_9313,N_8518,N_8674);
nor U9314 (N_9314,N_8755,N_8822);
nand U9315 (N_9315,N_8441,N_8924);
or U9316 (N_9316,N_8831,N_8998);
nand U9317 (N_9317,N_8474,N_8733);
or U9318 (N_9318,N_8771,N_8354);
nor U9319 (N_9319,N_8472,N_8351);
nand U9320 (N_9320,N_8550,N_8290);
xnor U9321 (N_9321,N_8974,N_8568);
nor U9322 (N_9322,N_8897,N_8646);
and U9323 (N_9323,N_8887,N_8337);
or U9324 (N_9324,N_8626,N_8293);
nor U9325 (N_9325,N_8915,N_8517);
or U9326 (N_9326,N_8327,N_8880);
or U9327 (N_9327,N_8821,N_8758);
or U9328 (N_9328,N_8424,N_8943);
or U9329 (N_9329,N_8751,N_8312);
nand U9330 (N_9330,N_8548,N_8567);
and U9331 (N_9331,N_8524,N_8321);
nor U9332 (N_9332,N_8799,N_8806);
nor U9333 (N_9333,N_8334,N_8538);
nand U9334 (N_9334,N_8481,N_8936);
and U9335 (N_9335,N_8804,N_8780);
or U9336 (N_9336,N_8483,N_8335);
nor U9337 (N_9337,N_8503,N_8599);
or U9338 (N_9338,N_8690,N_8927);
nand U9339 (N_9339,N_8753,N_8692);
nand U9340 (N_9340,N_8571,N_8317);
or U9341 (N_9341,N_8605,N_8835);
nand U9342 (N_9342,N_8972,N_8432);
or U9343 (N_9343,N_8704,N_8415);
nand U9344 (N_9344,N_8640,N_8347);
nand U9345 (N_9345,N_8553,N_8562);
xor U9346 (N_9346,N_8894,N_8371);
or U9347 (N_9347,N_8946,N_8461);
and U9348 (N_9348,N_8624,N_8306);
and U9349 (N_9349,N_8750,N_8391);
xor U9350 (N_9350,N_8952,N_8525);
nand U9351 (N_9351,N_8856,N_8643);
and U9352 (N_9352,N_8710,N_8917);
nand U9353 (N_9353,N_8613,N_8608);
nor U9354 (N_9354,N_8739,N_8748);
or U9355 (N_9355,N_8284,N_8369);
xor U9356 (N_9356,N_8698,N_8342);
nor U9357 (N_9357,N_8577,N_8931);
and U9358 (N_9358,N_8493,N_8849);
nor U9359 (N_9359,N_8641,N_8515);
or U9360 (N_9360,N_8818,N_8343);
or U9361 (N_9361,N_8694,N_8353);
and U9362 (N_9362,N_8803,N_8781);
and U9363 (N_9363,N_8500,N_8535);
xor U9364 (N_9364,N_8744,N_8276);
xor U9365 (N_9365,N_8872,N_8819);
xor U9366 (N_9366,N_8418,N_8464);
nand U9367 (N_9367,N_8395,N_8575);
nand U9368 (N_9368,N_8459,N_8482);
and U9369 (N_9369,N_8741,N_8473);
nor U9370 (N_9370,N_8257,N_8954);
and U9371 (N_9371,N_8888,N_8789);
and U9372 (N_9372,N_8378,N_8906);
and U9373 (N_9373,N_8886,N_8968);
nor U9374 (N_9374,N_8960,N_8377);
nor U9375 (N_9375,N_8755,N_8693);
and U9376 (N_9376,N_8944,N_8646);
or U9377 (N_9377,N_8966,N_8597);
xor U9378 (N_9378,N_8893,N_8317);
nor U9379 (N_9379,N_8469,N_8410);
and U9380 (N_9380,N_8850,N_8465);
nand U9381 (N_9381,N_8522,N_8606);
or U9382 (N_9382,N_8988,N_8504);
or U9383 (N_9383,N_8715,N_8974);
nand U9384 (N_9384,N_8685,N_8482);
nor U9385 (N_9385,N_8391,N_8399);
or U9386 (N_9386,N_8351,N_8969);
or U9387 (N_9387,N_8291,N_8363);
and U9388 (N_9388,N_8567,N_8713);
nand U9389 (N_9389,N_8796,N_8269);
nand U9390 (N_9390,N_8945,N_8809);
nand U9391 (N_9391,N_8279,N_8763);
xor U9392 (N_9392,N_8536,N_8639);
nor U9393 (N_9393,N_8539,N_8898);
or U9394 (N_9394,N_8531,N_8418);
nor U9395 (N_9395,N_8500,N_8567);
or U9396 (N_9396,N_8835,N_8335);
or U9397 (N_9397,N_8471,N_8307);
xnor U9398 (N_9398,N_8425,N_8601);
xor U9399 (N_9399,N_8389,N_8780);
nand U9400 (N_9400,N_8823,N_8342);
xnor U9401 (N_9401,N_8409,N_8820);
nor U9402 (N_9402,N_8633,N_8395);
xor U9403 (N_9403,N_8789,N_8972);
and U9404 (N_9404,N_8301,N_8779);
or U9405 (N_9405,N_8482,N_8714);
or U9406 (N_9406,N_8328,N_8338);
nor U9407 (N_9407,N_8708,N_8341);
and U9408 (N_9408,N_8781,N_8306);
or U9409 (N_9409,N_8653,N_8512);
and U9410 (N_9410,N_8896,N_8297);
and U9411 (N_9411,N_8456,N_8293);
or U9412 (N_9412,N_8821,N_8844);
or U9413 (N_9413,N_8847,N_8489);
nand U9414 (N_9414,N_8438,N_8298);
nor U9415 (N_9415,N_8366,N_8567);
nand U9416 (N_9416,N_8915,N_8281);
or U9417 (N_9417,N_8803,N_8448);
and U9418 (N_9418,N_8972,N_8728);
and U9419 (N_9419,N_8260,N_8588);
nor U9420 (N_9420,N_8913,N_8449);
and U9421 (N_9421,N_8342,N_8849);
nor U9422 (N_9422,N_8873,N_8319);
or U9423 (N_9423,N_8783,N_8261);
xnor U9424 (N_9424,N_8571,N_8285);
or U9425 (N_9425,N_8585,N_8563);
or U9426 (N_9426,N_8264,N_8458);
or U9427 (N_9427,N_8385,N_8912);
and U9428 (N_9428,N_8597,N_8944);
or U9429 (N_9429,N_8693,N_8307);
nand U9430 (N_9430,N_8695,N_8309);
and U9431 (N_9431,N_8480,N_8760);
nor U9432 (N_9432,N_8600,N_8825);
nand U9433 (N_9433,N_8786,N_8293);
or U9434 (N_9434,N_8416,N_8654);
nor U9435 (N_9435,N_8904,N_8402);
and U9436 (N_9436,N_8345,N_8624);
and U9437 (N_9437,N_8766,N_8344);
and U9438 (N_9438,N_8735,N_8611);
and U9439 (N_9439,N_8980,N_8795);
or U9440 (N_9440,N_8482,N_8259);
nand U9441 (N_9441,N_8326,N_8726);
nor U9442 (N_9442,N_8979,N_8375);
xor U9443 (N_9443,N_8736,N_8286);
nand U9444 (N_9444,N_8713,N_8554);
or U9445 (N_9445,N_8628,N_8810);
or U9446 (N_9446,N_8957,N_8558);
nor U9447 (N_9447,N_8735,N_8581);
or U9448 (N_9448,N_8960,N_8990);
nand U9449 (N_9449,N_8841,N_8463);
or U9450 (N_9450,N_8509,N_8301);
and U9451 (N_9451,N_8612,N_8564);
nor U9452 (N_9452,N_8348,N_8482);
nor U9453 (N_9453,N_8650,N_8334);
nand U9454 (N_9454,N_8537,N_8539);
or U9455 (N_9455,N_8684,N_8532);
nand U9456 (N_9456,N_8589,N_8445);
nor U9457 (N_9457,N_8457,N_8489);
or U9458 (N_9458,N_8806,N_8777);
or U9459 (N_9459,N_8686,N_8595);
nor U9460 (N_9460,N_8446,N_8509);
nand U9461 (N_9461,N_8355,N_8416);
nor U9462 (N_9462,N_8512,N_8601);
or U9463 (N_9463,N_8704,N_8420);
and U9464 (N_9464,N_8267,N_8436);
nor U9465 (N_9465,N_8548,N_8996);
nand U9466 (N_9466,N_8608,N_8698);
xnor U9467 (N_9467,N_8446,N_8457);
nand U9468 (N_9468,N_8698,N_8668);
nand U9469 (N_9469,N_8321,N_8527);
nor U9470 (N_9470,N_8513,N_8594);
xor U9471 (N_9471,N_8659,N_8974);
and U9472 (N_9472,N_8338,N_8504);
or U9473 (N_9473,N_8603,N_8799);
or U9474 (N_9474,N_8568,N_8438);
nor U9475 (N_9475,N_8310,N_8909);
nor U9476 (N_9476,N_8776,N_8595);
nand U9477 (N_9477,N_8554,N_8932);
nand U9478 (N_9478,N_8619,N_8944);
nor U9479 (N_9479,N_8661,N_8781);
nand U9480 (N_9480,N_8972,N_8583);
or U9481 (N_9481,N_8310,N_8751);
and U9482 (N_9482,N_8802,N_8647);
nand U9483 (N_9483,N_8519,N_8661);
xor U9484 (N_9484,N_8466,N_8774);
nand U9485 (N_9485,N_8529,N_8411);
nor U9486 (N_9486,N_8495,N_8526);
and U9487 (N_9487,N_8735,N_8805);
xnor U9488 (N_9488,N_8970,N_8781);
xor U9489 (N_9489,N_8525,N_8479);
and U9490 (N_9490,N_8378,N_8807);
nand U9491 (N_9491,N_8495,N_8290);
or U9492 (N_9492,N_8955,N_8992);
xor U9493 (N_9493,N_8471,N_8458);
nor U9494 (N_9494,N_8398,N_8535);
nor U9495 (N_9495,N_8835,N_8411);
and U9496 (N_9496,N_8506,N_8830);
nand U9497 (N_9497,N_8986,N_8798);
nand U9498 (N_9498,N_8336,N_8547);
nor U9499 (N_9499,N_8820,N_8500);
nand U9500 (N_9500,N_8554,N_8587);
nor U9501 (N_9501,N_8880,N_8341);
and U9502 (N_9502,N_8637,N_8576);
nor U9503 (N_9503,N_8717,N_8309);
or U9504 (N_9504,N_8663,N_8931);
or U9505 (N_9505,N_8991,N_8884);
nand U9506 (N_9506,N_8875,N_8747);
nand U9507 (N_9507,N_8332,N_8525);
or U9508 (N_9508,N_8266,N_8510);
nor U9509 (N_9509,N_8711,N_8516);
nand U9510 (N_9510,N_8972,N_8543);
or U9511 (N_9511,N_8524,N_8251);
nor U9512 (N_9512,N_8378,N_8574);
nor U9513 (N_9513,N_8280,N_8708);
or U9514 (N_9514,N_8972,N_8848);
and U9515 (N_9515,N_8432,N_8693);
nand U9516 (N_9516,N_8416,N_8849);
or U9517 (N_9517,N_8778,N_8395);
or U9518 (N_9518,N_8502,N_8559);
nor U9519 (N_9519,N_8961,N_8728);
and U9520 (N_9520,N_8630,N_8269);
nor U9521 (N_9521,N_8718,N_8832);
xor U9522 (N_9522,N_8377,N_8502);
xnor U9523 (N_9523,N_8774,N_8558);
and U9524 (N_9524,N_8464,N_8498);
nor U9525 (N_9525,N_8777,N_8431);
or U9526 (N_9526,N_8785,N_8892);
and U9527 (N_9527,N_8834,N_8258);
nor U9528 (N_9528,N_8268,N_8917);
nand U9529 (N_9529,N_8497,N_8541);
nand U9530 (N_9530,N_8884,N_8685);
xor U9531 (N_9531,N_8575,N_8397);
nand U9532 (N_9532,N_8912,N_8575);
nor U9533 (N_9533,N_8253,N_8281);
nand U9534 (N_9534,N_8329,N_8935);
and U9535 (N_9535,N_8685,N_8598);
nand U9536 (N_9536,N_8274,N_8368);
nor U9537 (N_9537,N_8494,N_8385);
nor U9538 (N_9538,N_8590,N_8540);
or U9539 (N_9539,N_8526,N_8368);
nor U9540 (N_9540,N_8365,N_8711);
nor U9541 (N_9541,N_8593,N_8815);
nor U9542 (N_9542,N_8973,N_8444);
xnor U9543 (N_9543,N_8710,N_8444);
nand U9544 (N_9544,N_8546,N_8729);
nor U9545 (N_9545,N_8636,N_8862);
nand U9546 (N_9546,N_8379,N_8908);
xnor U9547 (N_9547,N_8807,N_8289);
nor U9548 (N_9548,N_8269,N_8290);
and U9549 (N_9549,N_8649,N_8252);
nand U9550 (N_9550,N_8981,N_8379);
nor U9551 (N_9551,N_8883,N_8879);
and U9552 (N_9552,N_8856,N_8272);
nor U9553 (N_9553,N_8621,N_8679);
nor U9554 (N_9554,N_8472,N_8269);
or U9555 (N_9555,N_8622,N_8601);
xnor U9556 (N_9556,N_8515,N_8696);
or U9557 (N_9557,N_8749,N_8700);
nor U9558 (N_9558,N_8545,N_8670);
nor U9559 (N_9559,N_8536,N_8927);
and U9560 (N_9560,N_8327,N_8899);
nor U9561 (N_9561,N_8301,N_8643);
and U9562 (N_9562,N_8957,N_8300);
nor U9563 (N_9563,N_8624,N_8878);
nor U9564 (N_9564,N_8766,N_8445);
or U9565 (N_9565,N_8837,N_8631);
and U9566 (N_9566,N_8620,N_8707);
nand U9567 (N_9567,N_8678,N_8564);
xnor U9568 (N_9568,N_8333,N_8616);
nor U9569 (N_9569,N_8375,N_8617);
or U9570 (N_9570,N_8584,N_8706);
nand U9571 (N_9571,N_8487,N_8643);
and U9572 (N_9572,N_8318,N_8977);
nand U9573 (N_9573,N_8625,N_8438);
nand U9574 (N_9574,N_8770,N_8387);
nor U9575 (N_9575,N_8341,N_8895);
xor U9576 (N_9576,N_8943,N_8652);
nor U9577 (N_9577,N_8778,N_8646);
and U9578 (N_9578,N_8873,N_8258);
or U9579 (N_9579,N_8299,N_8686);
nand U9580 (N_9580,N_8800,N_8484);
and U9581 (N_9581,N_8763,N_8485);
nor U9582 (N_9582,N_8964,N_8874);
or U9583 (N_9583,N_8980,N_8452);
nor U9584 (N_9584,N_8626,N_8437);
or U9585 (N_9585,N_8747,N_8545);
nor U9586 (N_9586,N_8476,N_8620);
and U9587 (N_9587,N_8767,N_8837);
nand U9588 (N_9588,N_8453,N_8489);
nor U9589 (N_9589,N_8349,N_8398);
nand U9590 (N_9590,N_8303,N_8268);
nand U9591 (N_9591,N_8358,N_8333);
and U9592 (N_9592,N_8929,N_8669);
nand U9593 (N_9593,N_8899,N_8549);
nor U9594 (N_9594,N_8370,N_8615);
xor U9595 (N_9595,N_8994,N_8829);
nand U9596 (N_9596,N_8353,N_8359);
nand U9597 (N_9597,N_8348,N_8557);
xor U9598 (N_9598,N_8787,N_8259);
nor U9599 (N_9599,N_8912,N_8447);
nand U9600 (N_9600,N_8929,N_8616);
nor U9601 (N_9601,N_8548,N_8867);
xor U9602 (N_9602,N_8975,N_8844);
nor U9603 (N_9603,N_8946,N_8827);
nand U9604 (N_9604,N_8285,N_8801);
xnor U9605 (N_9605,N_8620,N_8988);
nor U9606 (N_9606,N_8492,N_8746);
nor U9607 (N_9607,N_8782,N_8624);
nand U9608 (N_9608,N_8655,N_8889);
or U9609 (N_9609,N_8975,N_8661);
xnor U9610 (N_9610,N_8519,N_8470);
and U9611 (N_9611,N_8944,N_8602);
and U9612 (N_9612,N_8977,N_8702);
and U9613 (N_9613,N_8811,N_8597);
or U9614 (N_9614,N_8729,N_8778);
nand U9615 (N_9615,N_8791,N_8696);
nand U9616 (N_9616,N_8493,N_8625);
and U9617 (N_9617,N_8499,N_8570);
and U9618 (N_9618,N_8639,N_8730);
and U9619 (N_9619,N_8736,N_8516);
nor U9620 (N_9620,N_8343,N_8288);
xor U9621 (N_9621,N_8905,N_8528);
xnor U9622 (N_9622,N_8662,N_8279);
nand U9623 (N_9623,N_8674,N_8263);
or U9624 (N_9624,N_8326,N_8757);
and U9625 (N_9625,N_8998,N_8969);
or U9626 (N_9626,N_8736,N_8612);
nand U9627 (N_9627,N_8951,N_8719);
or U9628 (N_9628,N_8403,N_8979);
nor U9629 (N_9629,N_8579,N_8624);
nor U9630 (N_9630,N_8657,N_8891);
xor U9631 (N_9631,N_8735,N_8292);
and U9632 (N_9632,N_8476,N_8856);
nand U9633 (N_9633,N_8496,N_8535);
or U9634 (N_9634,N_8674,N_8323);
nor U9635 (N_9635,N_8960,N_8261);
or U9636 (N_9636,N_8826,N_8431);
or U9637 (N_9637,N_8323,N_8313);
and U9638 (N_9638,N_8560,N_8564);
nand U9639 (N_9639,N_8696,N_8808);
and U9640 (N_9640,N_8421,N_8449);
xnor U9641 (N_9641,N_8777,N_8637);
nor U9642 (N_9642,N_8403,N_8761);
or U9643 (N_9643,N_8698,N_8817);
nor U9644 (N_9644,N_8480,N_8723);
xnor U9645 (N_9645,N_8271,N_8516);
or U9646 (N_9646,N_8869,N_8265);
nor U9647 (N_9647,N_8534,N_8797);
nor U9648 (N_9648,N_8404,N_8622);
or U9649 (N_9649,N_8395,N_8598);
or U9650 (N_9650,N_8459,N_8456);
and U9651 (N_9651,N_8404,N_8800);
nand U9652 (N_9652,N_8706,N_8448);
nand U9653 (N_9653,N_8905,N_8367);
or U9654 (N_9654,N_8419,N_8326);
or U9655 (N_9655,N_8798,N_8612);
and U9656 (N_9656,N_8966,N_8891);
and U9657 (N_9657,N_8721,N_8585);
or U9658 (N_9658,N_8701,N_8263);
nand U9659 (N_9659,N_8699,N_8642);
and U9660 (N_9660,N_8333,N_8332);
or U9661 (N_9661,N_8566,N_8731);
nand U9662 (N_9662,N_8271,N_8742);
xnor U9663 (N_9663,N_8281,N_8560);
and U9664 (N_9664,N_8654,N_8492);
xor U9665 (N_9665,N_8873,N_8327);
xnor U9666 (N_9666,N_8264,N_8615);
nand U9667 (N_9667,N_8396,N_8272);
and U9668 (N_9668,N_8859,N_8702);
and U9669 (N_9669,N_8267,N_8420);
or U9670 (N_9670,N_8312,N_8428);
and U9671 (N_9671,N_8529,N_8590);
nor U9672 (N_9672,N_8343,N_8540);
nand U9673 (N_9673,N_8940,N_8988);
and U9674 (N_9674,N_8845,N_8887);
nand U9675 (N_9675,N_8430,N_8968);
and U9676 (N_9676,N_8805,N_8657);
or U9677 (N_9677,N_8516,N_8662);
or U9678 (N_9678,N_8939,N_8321);
or U9679 (N_9679,N_8940,N_8756);
and U9680 (N_9680,N_8524,N_8408);
or U9681 (N_9681,N_8371,N_8560);
and U9682 (N_9682,N_8615,N_8696);
nor U9683 (N_9683,N_8585,N_8614);
nand U9684 (N_9684,N_8627,N_8458);
nand U9685 (N_9685,N_8649,N_8424);
nand U9686 (N_9686,N_8476,N_8387);
and U9687 (N_9687,N_8741,N_8508);
or U9688 (N_9688,N_8911,N_8836);
and U9689 (N_9689,N_8924,N_8935);
nand U9690 (N_9690,N_8928,N_8746);
nand U9691 (N_9691,N_8409,N_8965);
nand U9692 (N_9692,N_8873,N_8474);
nor U9693 (N_9693,N_8396,N_8427);
nand U9694 (N_9694,N_8410,N_8521);
xor U9695 (N_9695,N_8912,N_8675);
and U9696 (N_9696,N_8808,N_8537);
nor U9697 (N_9697,N_8441,N_8778);
xor U9698 (N_9698,N_8682,N_8479);
nand U9699 (N_9699,N_8509,N_8773);
nor U9700 (N_9700,N_8937,N_8678);
or U9701 (N_9701,N_8941,N_8544);
and U9702 (N_9702,N_8266,N_8468);
and U9703 (N_9703,N_8990,N_8339);
nor U9704 (N_9704,N_8570,N_8321);
xnor U9705 (N_9705,N_8505,N_8922);
xor U9706 (N_9706,N_8610,N_8355);
nor U9707 (N_9707,N_8793,N_8856);
or U9708 (N_9708,N_8535,N_8866);
and U9709 (N_9709,N_8410,N_8562);
and U9710 (N_9710,N_8375,N_8587);
nand U9711 (N_9711,N_8831,N_8600);
nand U9712 (N_9712,N_8400,N_8563);
nand U9713 (N_9713,N_8463,N_8890);
and U9714 (N_9714,N_8603,N_8567);
or U9715 (N_9715,N_8589,N_8296);
and U9716 (N_9716,N_8844,N_8294);
nand U9717 (N_9717,N_8315,N_8634);
nand U9718 (N_9718,N_8899,N_8449);
and U9719 (N_9719,N_8810,N_8835);
nand U9720 (N_9720,N_8372,N_8520);
nand U9721 (N_9721,N_8618,N_8927);
or U9722 (N_9722,N_8647,N_8469);
or U9723 (N_9723,N_8315,N_8499);
and U9724 (N_9724,N_8454,N_8558);
nand U9725 (N_9725,N_8464,N_8991);
and U9726 (N_9726,N_8649,N_8346);
nor U9727 (N_9727,N_8484,N_8503);
or U9728 (N_9728,N_8345,N_8366);
and U9729 (N_9729,N_8777,N_8843);
or U9730 (N_9730,N_8340,N_8981);
nand U9731 (N_9731,N_8489,N_8772);
nor U9732 (N_9732,N_8760,N_8616);
and U9733 (N_9733,N_8675,N_8291);
and U9734 (N_9734,N_8640,N_8901);
or U9735 (N_9735,N_8801,N_8666);
nand U9736 (N_9736,N_8508,N_8873);
nor U9737 (N_9737,N_8457,N_8424);
nand U9738 (N_9738,N_8427,N_8822);
nor U9739 (N_9739,N_8986,N_8536);
xor U9740 (N_9740,N_8941,N_8928);
nor U9741 (N_9741,N_8663,N_8581);
nor U9742 (N_9742,N_8621,N_8309);
nand U9743 (N_9743,N_8367,N_8420);
and U9744 (N_9744,N_8497,N_8619);
nand U9745 (N_9745,N_8571,N_8682);
or U9746 (N_9746,N_8658,N_8454);
or U9747 (N_9747,N_8523,N_8497);
xnor U9748 (N_9748,N_8980,N_8266);
nor U9749 (N_9749,N_8746,N_8573);
or U9750 (N_9750,N_9236,N_9147);
nand U9751 (N_9751,N_9096,N_9567);
nor U9752 (N_9752,N_9102,N_9228);
and U9753 (N_9753,N_9749,N_9615);
and U9754 (N_9754,N_9085,N_9705);
nor U9755 (N_9755,N_9437,N_9552);
and U9756 (N_9756,N_9033,N_9470);
and U9757 (N_9757,N_9691,N_9222);
or U9758 (N_9758,N_9141,N_9081);
nand U9759 (N_9759,N_9010,N_9646);
nand U9760 (N_9760,N_9494,N_9038);
nor U9761 (N_9761,N_9082,N_9016);
nand U9762 (N_9762,N_9233,N_9592);
or U9763 (N_9763,N_9678,N_9075);
nor U9764 (N_9764,N_9602,N_9162);
nor U9765 (N_9765,N_9306,N_9544);
and U9766 (N_9766,N_9279,N_9617);
or U9767 (N_9767,N_9373,N_9040);
and U9768 (N_9768,N_9153,N_9628);
nand U9769 (N_9769,N_9686,N_9748);
and U9770 (N_9770,N_9507,N_9625);
nand U9771 (N_9771,N_9323,N_9583);
nor U9772 (N_9772,N_9298,N_9369);
nand U9773 (N_9773,N_9384,N_9716);
or U9774 (N_9774,N_9501,N_9274);
xnor U9775 (N_9775,N_9217,N_9256);
or U9776 (N_9776,N_9019,N_9513);
and U9777 (N_9777,N_9317,N_9376);
and U9778 (N_9778,N_9562,N_9670);
or U9779 (N_9779,N_9297,N_9121);
nor U9780 (N_9780,N_9607,N_9395);
nand U9781 (N_9781,N_9512,N_9639);
nand U9782 (N_9782,N_9215,N_9407);
xnor U9783 (N_9783,N_9740,N_9537);
nand U9784 (N_9784,N_9619,N_9028);
and U9785 (N_9785,N_9420,N_9166);
or U9786 (N_9786,N_9148,N_9101);
nor U9787 (N_9787,N_9597,N_9269);
nor U9788 (N_9788,N_9098,N_9047);
nor U9789 (N_9789,N_9084,N_9363);
nand U9790 (N_9790,N_9076,N_9720);
nor U9791 (N_9791,N_9108,N_9527);
or U9792 (N_9792,N_9574,N_9163);
or U9793 (N_9793,N_9219,N_9123);
xor U9794 (N_9794,N_9444,N_9186);
and U9795 (N_9795,N_9079,N_9568);
or U9796 (N_9796,N_9471,N_9286);
nand U9797 (N_9797,N_9432,N_9064);
nor U9798 (N_9798,N_9232,N_9000);
or U9799 (N_9799,N_9611,N_9252);
nor U9800 (N_9800,N_9709,N_9667);
and U9801 (N_9801,N_9368,N_9331);
nor U9802 (N_9802,N_9711,N_9227);
or U9803 (N_9803,N_9177,N_9090);
nor U9804 (N_9804,N_9195,N_9546);
or U9805 (N_9805,N_9659,N_9253);
or U9806 (N_9806,N_9169,N_9724);
and U9807 (N_9807,N_9721,N_9396);
or U9808 (N_9808,N_9041,N_9579);
or U9809 (N_9809,N_9487,N_9402);
and U9810 (N_9810,N_9151,N_9594);
nor U9811 (N_9811,N_9220,N_9208);
and U9812 (N_9812,N_9155,N_9235);
and U9813 (N_9813,N_9080,N_9638);
xor U9814 (N_9814,N_9509,N_9747);
nor U9815 (N_9815,N_9685,N_9367);
and U9816 (N_9816,N_9677,N_9290);
nor U9817 (N_9817,N_9077,N_9735);
or U9818 (N_9818,N_9534,N_9493);
and U9819 (N_9819,N_9743,N_9436);
or U9820 (N_9820,N_9308,N_9003);
nor U9821 (N_9821,N_9392,N_9673);
nor U9822 (N_9822,N_9372,N_9431);
xnor U9823 (N_9823,N_9245,N_9401);
or U9824 (N_9824,N_9438,N_9456);
nor U9825 (N_9825,N_9429,N_9281);
or U9826 (N_9826,N_9706,N_9058);
xor U9827 (N_9827,N_9347,N_9107);
xor U9828 (N_9828,N_9135,N_9455);
nor U9829 (N_9829,N_9015,N_9504);
nand U9830 (N_9830,N_9741,N_9205);
and U9831 (N_9831,N_9035,N_9626);
nand U9832 (N_9832,N_9114,N_9127);
nor U9833 (N_9833,N_9422,N_9557);
nand U9834 (N_9834,N_9325,N_9543);
nand U9835 (N_9835,N_9655,N_9074);
xor U9836 (N_9836,N_9426,N_9138);
nor U9837 (N_9837,N_9196,N_9553);
or U9838 (N_9838,N_9318,N_9599);
or U9839 (N_9839,N_9020,N_9311);
and U9840 (N_9840,N_9669,N_9320);
and U9841 (N_9841,N_9604,N_9581);
and U9842 (N_9842,N_9353,N_9578);
nand U9843 (N_9843,N_9689,N_9476);
nor U9844 (N_9844,N_9259,N_9199);
nor U9845 (N_9845,N_9443,N_9405);
and U9846 (N_9846,N_9343,N_9337);
xor U9847 (N_9847,N_9315,N_9616);
and U9848 (N_9848,N_9404,N_9414);
nor U9849 (N_9849,N_9461,N_9103);
nand U9850 (N_9850,N_9702,N_9417);
or U9851 (N_9851,N_9278,N_9660);
and U9852 (N_9852,N_9575,N_9067);
nand U9853 (N_9853,N_9653,N_9486);
and U9854 (N_9854,N_9137,N_9412);
nand U9855 (N_9855,N_9459,N_9267);
xnor U9856 (N_9856,N_9351,N_9563);
or U9857 (N_9857,N_9004,N_9388);
nand U9858 (N_9858,N_9571,N_9072);
or U9859 (N_9859,N_9460,N_9582);
xor U9860 (N_9860,N_9230,N_9591);
or U9861 (N_9861,N_9484,N_9265);
or U9862 (N_9862,N_9654,N_9111);
nor U9863 (N_9863,N_9416,N_9188);
or U9864 (N_9864,N_9039,N_9737);
nor U9865 (N_9865,N_9387,N_9334);
or U9866 (N_9866,N_9301,N_9545);
nand U9867 (N_9867,N_9231,N_9349);
and U9868 (N_9868,N_9167,N_9425);
nand U9869 (N_9869,N_9419,N_9503);
or U9870 (N_9870,N_9475,N_9719);
nor U9871 (N_9871,N_9451,N_9131);
and U9872 (N_9872,N_9239,N_9187);
or U9873 (N_9873,N_9309,N_9251);
nor U9874 (N_9874,N_9009,N_9088);
xor U9875 (N_9875,N_9261,N_9056);
nor U9876 (N_9876,N_9356,N_9549);
or U9877 (N_9877,N_9738,N_9474);
nor U9878 (N_9878,N_9435,N_9360);
nand U9879 (N_9879,N_9596,N_9365);
xnor U9880 (N_9880,N_9694,N_9590);
and U9881 (N_9881,N_9700,N_9531);
nand U9882 (N_9882,N_9120,N_9464);
nand U9883 (N_9883,N_9620,N_9270);
nor U9884 (N_9884,N_9099,N_9658);
nor U9885 (N_9885,N_9168,N_9674);
and U9886 (N_9886,N_9313,N_9011);
or U9887 (N_9887,N_9031,N_9715);
and U9888 (N_9888,N_9661,N_9069);
or U9889 (N_9889,N_9371,N_9164);
nor U9890 (N_9890,N_9515,N_9091);
nand U9891 (N_9891,N_9022,N_9324);
nor U9892 (N_9892,N_9725,N_9050);
nor U9893 (N_9893,N_9296,N_9642);
nor U9894 (N_9894,N_9283,N_9176);
xnor U9895 (N_9895,N_9466,N_9282);
nand U9896 (N_9896,N_9478,N_9303);
xor U9897 (N_9897,N_9714,N_9154);
nor U9898 (N_9898,N_9021,N_9518);
and U9899 (N_9899,N_9338,N_9586);
xnor U9900 (N_9900,N_9379,N_9183);
nand U9901 (N_9901,N_9200,N_9248);
nand U9902 (N_9902,N_9555,N_9644);
nand U9903 (N_9903,N_9558,N_9535);
or U9904 (N_9904,N_9139,N_9389);
or U9905 (N_9905,N_9406,N_9564);
nor U9906 (N_9906,N_9733,N_9649);
nor U9907 (N_9907,N_9304,N_9526);
and U9908 (N_9908,N_9173,N_9449);
nand U9909 (N_9909,N_9226,N_9539);
nand U9910 (N_9910,N_9624,N_9608);
and U9911 (N_9911,N_9410,N_9601);
and U9912 (N_9912,N_9722,N_9284);
or U9913 (N_9913,N_9745,N_9631);
nor U9914 (N_9914,N_9580,N_9223);
and U9915 (N_9915,N_9089,N_9002);
nor U9916 (N_9916,N_9275,N_9394);
xor U9917 (N_9917,N_9397,N_9502);
nor U9918 (N_9918,N_9012,N_9057);
nand U9919 (N_9919,N_9124,N_9676);
and U9920 (N_9920,N_9051,N_9152);
nor U9921 (N_9921,N_9292,N_9472);
nand U9922 (N_9922,N_9603,N_9190);
xor U9923 (N_9923,N_9354,N_9744);
nor U9924 (N_9924,N_9062,N_9598);
nand U9925 (N_9925,N_9656,N_9143);
or U9926 (N_9926,N_9211,N_9481);
nor U9927 (N_9927,N_9746,N_9541);
nand U9928 (N_9928,N_9201,N_9565);
or U9929 (N_9929,N_9034,N_9496);
nor U9930 (N_9930,N_9189,N_9480);
xnor U9931 (N_9931,N_9636,N_9713);
nor U9932 (N_9932,N_9448,N_9358);
and U9933 (N_9933,N_9178,N_9623);
and U9934 (N_9934,N_9375,N_9008);
xor U9935 (N_9935,N_9287,N_9238);
or U9936 (N_9936,N_9520,N_9447);
nor U9937 (N_9937,N_9209,N_9731);
nand U9938 (N_9938,N_9648,N_9693);
and U9939 (N_9939,N_9122,N_9453);
and U9940 (N_9940,N_9119,N_9680);
xor U9941 (N_9941,N_9637,N_9584);
nand U9942 (N_9942,N_9357,N_9548);
xnor U9943 (N_9943,N_9030,N_9145);
nand U9944 (N_9944,N_9622,N_9027);
nor U9945 (N_9945,N_9174,N_9202);
nor U9946 (N_9946,N_9576,N_9696);
nand U9947 (N_9947,N_9385,N_9156);
nand U9948 (N_9948,N_9634,N_9730);
nor U9949 (N_9949,N_9718,N_9662);
nand U9950 (N_9950,N_9382,N_9577);
and U9951 (N_9951,N_9643,N_9117);
or U9952 (N_9952,N_9723,N_9078);
or U9953 (N_9953,N_9408,N_9411);
or U9954 (N_9954,N_9398,N_9441);
nor U9955 (N_9955,N_9013,N_9687);
nor U9956 (N_9956,N_9043,N_9630);
or U9957 (N_9957,N_9467,N_9364);
nor U9958 (N_9958,N_9497,N_9052);
nand U9959 (N_9959,N_9247,N_9682);
or U9960 (N_9960,N_9328,N_9633);
nor U9961 (N_9961,N_9066,N_9529);
or U9962 (N_9962,N_9029,N_9116);
nor U9963 (N_9963,N_9403,N_9295);
xnor U9964 (N_9964,N_9488,N_9427);
nand U9965 (N_9965,N_9508,N_9194);
and U9966 (N_9966,N_9490,N_9130);
nor U9967 (N_9967,N_9479,N_9516);
nand U9968 (N_9968,N_9260,N_9126);
nand U9969 (N_9969,N_9609,N_9136);
nand U9970 (N_9970,N_9024,N_9149);
and U9971 (N_9971,N_9469,N_9439);
or U9972 (N_9972,N_9005,N_9273);
xor U9973 (N_9973,N_9629,N_9344);
xor U9974 (N_9974,N_9665,N_9255);
and U9975 (N_9975,N_9172,N_9310);
nor U9976 (N_9976,N_9105,N_9129);
nand U9977 (N_9977,N_9510,N_9418);
nand U9978 (N_9978,N_9302,N_9218);
xnor U9979 (N_9979,N_9386,N_9554);
or U9980 (N_9980,N_9442,N_9048);
or U9981 (N_9981,N_9044,N_9359);
and U9982 (N_9982,N_9133,N_9161);
or U9983 (N_9983,N_9647,N_9006);
xnor U9984 (N_9984,N_9225,N_9146);
and U9985 (N_9985,N_9180,N_9125);
nor U9986 (N_9986,N_9593,N_9113);
nor U9987 (N_9987,N_9538,N_9316);
and U9988 (N_9988,N_9198,N_9073);
nor U9989 (N_9989,N_9229,N_9366);
nand U9990 (N_9990,N_9551,N_9452);
nand U9991 (N_9991,N_9258,N_9063);
nand U9992 (N_9992,N_9703,N_9109);
xor U9993 (N_9993,N_9684,N_9632);
nor U9994 (N_9994,N_9519,N_9652);
xnor U9995 (N_9995,N_9547,N_9068);
or U9996 (N_9996,N_9413,N_9645);
and U9997 (N_9997,N_9492,N_9224);
nor U9998 (N_9998,N_9300,N_9672);
nor U9999 (N_9999,N_9112,N_9536);
or U10000 (N_10000,N_9335,N_9289);
and U10001 (N_10001,N_9561,N_9339);
and U10002 (N_10002,N_9485,N_9635);
nor U10003 (N_10003,N_9206,N_9556);
and U10004 (N_10004,N_9179,N_9540);
nand U10005 (N_10005,N_9134,N_9707);
nor U10006 (N_10006,N_9327,N_9499);
or U10007 (N_10007,N_9621,N_9681);
nor U10008 (N_10008,N_9679,N_9506);
or U10009 (N_10009,N_9065,N_9175);
or U10010 (N_10010,N_9588,N_9511);
nor U10011 (N_10011,N_9465,N_9184);
nor U10012 (N_10012,N_9695,N_9093);
and U10013 (N_10013,N_9237,N_9061);
nor U10014 (N_10014,N_9450,N_9675);
and U10015 (N_10015,N_9560,N_9651);
nand U10016 (N_10016,N_9342,N_9244);
nor U10017 (N_10017,N_9482,N_9573);
nand U10018 (N_10018,N_9525,N_9158);
nor U10019 (N_10019,N_9350,N_9514);
and U10020 (N_10020,N_9160,N_9104);
nand U10021 (N_10021,N_9585,N_9517);
and U10022 (N_10022,N_9042,N_9374);
or U10023 (N_10023,N_9037,N_9701);
nand U10024 (N_10024,N_9213,N_9370);
or U10025 (N_10025,N_9348,N_9291);
nand U10026 (N_10026,N_9277,N_9729);
nor U10027 (N_10027,N_9212,N_9393);
nand U10028 (N_10028,N_9717,N_9106);
nand U10029 (N_10029,N_9060,N_9692);
nand U10030 (N_10030,N_9268,N_9234);
nand U10031 (N_10031,N_9293,N_9566);
or U10032 (N_10032,N_9587,N_9032);
and U10033 (N_10033,N_9118,N_9262);
and U10034 (N_10034,N_9036,N_9346);
and U10035 (N_10035,N_9266,N_9380);
nand U10036 (N_10036,N_9528,N_9390);
nand U10037 (N_10037,N_9627,N_9263);
and U10038 (N_10038,N_9522,N_9288);
nor U10039 (N_10039,N_9663,N_9440);
and U10040 (N_10040,N_9362,N_9391);
nand U10041 (N_10041,N_9142,N_9115);
nand U10042 (N_10042,N_9250,N_9664);
or U10043 (N_10043,N_9181,N_9415);
and U10044 (N_10044,N_9710,N_9462);
xnor U10045 (N_10045,N_9312,N_9683);
and U10046 (N_10046,N_9421,N_9704);
nand U10047 (N_10047,N_9100,N_9246);
or U10048 (N_10048,N_9688,N_9092);
nand U10049 (N_10049,N_9197,N_9613);
nand U10050 (N_10050,N_9221,N_9171);
nand U10051 (N_10051,N_9477,N_9589);
nor U10052 (N_10052,N_9192,N_9017);
or U10053 (N_10053,N_9473,N_9666);
xor U10054 (N_10054,N_9204,N_9428);
nand U10055 (N_10055,N_9150,N_9378);
nand U10056 (N_10056,N_9018,N_9249);
nand U10057 (N_10057,N_9600,N_9739);
nand U10058 (N_10058,N_9144,N_9657);
nor U10059 (N_10059,N_9214,N_9569);
nor U10060 (N_10060,N_9305,N_9157);
nand U10061 (N_10061,N_9400,N_9500);
nand U10062 (N_10062,N_9742,N_9322);
nand U10063 (N_10063,N_9326,N_9614);
nor U10064 (N_10064,N_9521,N_9505);
nor U10065 (N_10065,N_9053,N_9399);
or U10066 (N_10066,N_9650,N_9285);
or U10067 (N_10067,N_9110,N_9430);
nand U10068 (N_10068,N_9671,N_9299);
or U10069 (N_10069,N_9340,N_9336);
and U10070 (N_10070,N_9445,N_9468);
xor U10071 (N_10071,N_9314,N_9023);
nand U10072 (N_10072,N_9446,N_9610);
or U10073 (N_10073,N_9330,N_9612);
nand U10074 (N_10074,N_9532,N_9046);
or U10075 (N_10075,N_9345,N_9458);
nand U10076 (N_10076,N_9054,N_9457);
nor U10077 (N_10077,N_9708,N_9203);
or U10078 (N_10078,N_9207,N_9128);
or U10079 (N_10079,N_9071,N_9045);
nor U10080 (N_10080,N_9240,N_9025);
or U10081 (N_10081,N_9559,N_9498);
nand U10082 (N_10082,N_9690,N_9381);
or U10083 (N_10083,N_9726,N_9618);
or U10084 (N_10084,N_9550,N_9533);
nand U10085 (N_10085,N_9524,N_9332);
nand U10086 (N_10086,N_9094,N_9132);
nand U10087 (N_10087,N_9007,N_9495);
nand U10088 (N_10088,N_9086,N_9170);
or U10089 (N_10089,N_9606,N_9595);
nand U10090 (N_10090,N_9319,N_9185);
nand U10091 (N_10091,N_9454,N_9434);
nand U10092 (N_10092,N_9605,N_9329);
and U10093 (N_10093,N_9083,N_9254);
or U10094 (N_10094,N_9276,N_9732);
or U10095 (N_10095,N_9165,N_9483);
or U10096 (N_10096,N_9489,N_9423);
nor U10097 (N_10097,N_9523,N_9242);
and U10098 (N_10098,N_9241,N_9272);
nand U10099 (N_10099,N_9307,N_9049);
nand U10100 (N_10100,N_9210,N_9697);
nor U10101 (N_10101,N_9191,N_9699);
nand U10102 (N_10102,N_9321,N_9409);
and U10103 (N_10103,N_9698,N_9333);
or U10104 (N_10104,N_9001,N_9216);
nor U10105 (N_10105,N_9140,N_9355);
and U10106 (N_10106,N_9352,N_9361);
and U10107 (N_10107,N_9728,N_9736);
nand U10108 (N_10108,N_9182,N_9640);
and U10109 (N_10109,N_9280,N_9070);
and U10110 (N_10110,N_9377,N_9087);
and U10111 (N_10111,N_9159,N_9055);
nor U10112 (N_10112,N_9341,N_9095);
nand U10113 (N_10113,N_9294,N_9463);
and U10114 (N_10114,N_9572,N_9668);
xnor U10115 (N_10115,N_9097,N_9257);
and U10116 (N_10116,N_9014,N_9530);
nor U10117 (N_10117,N_9271,N_9712);
nor U10118 (N_10118,N_9491,N_9734);
or U10119 (N_10119,N_9727,N_9542);
nor U10120 (N_10120,N_9424,N_9570);
and U10121 (N_10121,N_9264,N_9059);
and U10122 (N_10122,N_9193,N_9641);
nor U10123 (N_10123,N_9026,N_9433);
nor U10124 (N_10124,N_9243,N_9383);
nand U10125 (N_10125,N_9318,N_9703);
nand U10126 (N_10126,N_9581,N_9638);
xor U10127 (N_10127,N_9275,N_9350);
nor U10128 (N_10128,N_9288,N_9589);
nand U10129 (N_10129,N_9282,N_9700);
and U10130 (N_10130,N_9497,N_9630);
and U10131 (N_10131,N_9121,N_9663);
and U10132 (N_10132,N_9735,N_9721);
or U10133 (N_10133,N_9234,N_9359);
xor U10134 (N_10134,N_9713,N_9741);
nand U10135 (N_10135,N_9131,N_9588);
nor U10136 (N_10136,N_9739,N_9025);
and U10137 (N_10137,N_9217,N_9341);
or U10138 (N_10138,N_9725,N_9588);
and U10139 (N_10139,N_9152,N_9158);
nand U10140 (N_10140,N_9020,N_9169);
nor U10141 (N_10141,N_9234,N_9142);
or U10142 (N_10142,N_9570,N_9258);
and U10143 (N_10143,N_9340,N_9421);
nand U10144 (N_10144,N_9670,N_9358);
nor U10145 (N_10145,N_9368,N_9653);
nor U10146 (N_10146,N_9043,N_9580);
or U10147 (N_10147,N_9239,N_9489);
nand U10148 (N_10148,N_9247,N_9488);
nand U10149 (N_10149,N_9037,N_9578);
and U10150 (N_10150,N_9140,N_9493);
nor U10151 (N_10151,N_9701,N_9145);
or U10152 (N_10152,N_9424,N_9162);
or U10153 (N_10153,N_9077,N_9700);
nand U10154 (N_10154,N_9184,N_9523);
or U10155 (N_10155,N_9255,N_9144);
nand U10156 (N_10156,N_9611,N_9144);
nor U10157 (N_10157,N_9688,N_9061);
and U10158 (N_10158,N_9382,N_9257);
xor U10159 (N_10159,N_9547,N_9275);
nor U10160 (N_10160,N_9331,N_9096);
nand U10161 (N_10161,N_9702,N_9030);
and U10162 (N_10162,N_9332,N_9370);
or U10163 (N_10163,N_9467,N_9558);
xnor U10164 (N_10164,N_9480,N_9112);
and U10165 (N_10165,N_9237,N_9012);
nor U10166 (N_10166,N_9198,N_9012);
or U10167 (N_10167,N_9562,N_9358);
or U10168 (N_10168,N_9087,N_9158);
xor U10169 (N_10169,N_9453,N_9342);
nor U10170 (N_10170,N_9511,N_9357);
nor U10171 (N_10171,N_9734,N_9685);
nand U10172 (N_10172,N_9088,N_9136);
nor U10173 (N_10173,N_9719,N_9028);
or U10174 (N_10174,N_9177,N_9355);
nand U10175 (N_10175,N_9675,N_9152);
or U10176 (N_10176,N_9679,N_9688);
or U10177 (N_10177,N_9363,N_9584);
and U10178 (N_10178,N_9105,N_9155);
nand U10179 (N_10179,N_9641,N_9061);
or U10180 (N_10180,N_9081,N_9118);
xor U10181 (N_10181,N_9452,N_9407);
nor U10182 (N_10182,N_9282,N_9212);
or U10183 (N_10183,N_9650,N_9078);
nand U10184 (N_10184,N_9286,N_9351);
or U10185 (N_10185,N_9083,N_9641);
nand U10186 (N_10186,N_9342,N_9438);
xnor U10187 (N_10187,N_9178,N_9604);
xnor U10188 (N_10188,N_9191,N_9514);
and U10189 (N_10189,N_9032,N_9208);
nor U10190 (N_10190,N_9235,N_9194);
xor U10191 (N_10191,N_9097,N_9547);
nand U10192 (N_10192,N_9426,N_9713);
and U10193 (N_10193,N_9615,N_9338);
nand U10194 (N_10194,N_9367,N_9284);
nand U10195 (N_10195,N_9053,N_9004);
and U10196 (N_10196,N_9436,N_9741);
nor U10197 (N_10197,N_9698,N_9108);
and U10198 (N_10198,N_9504,N_9237);
or U10199 (N_10199,N_9358,N_9090);
xnor U10200 (N_10200,N_9120,N_9598);
xor U10201 (N_10201,N_9604,N_9171);
or U10202 (N_10202,N_9139,N_9253);
and U10203 (N_10203,N_9280,N_9281);
and U10204 (N_10204,N_9105,N_9279);
or U10205 (N_10205,N_9630,N_9645);
or U10206 (N_10206,N_9403,N_9215);
and U10207 (N_10207,N_9204,N_9525);
and U10208 (N_10208,N_9152,N_9383);
and U10209 (N_10209,N_9327,N_9107);
xor U10210 (N_10210,N_9281,N_9268);
and U10211 (N_10211,N_9062,N_9240);
xor U10212 (N_10212,N_9307,N_9413);
nand U10213 (N_10213,N_9140,N_9356);
and U10214 (N_10214,N_9389,N_9395);
or U10215 (N_10215,N_9352,N_9290);
nand U10216 (N_10216,N_9585,N_9334);
or U10217 (N_10217,N_9463,N_9508);
or U10218 (N_10218,N_9160,N_9192);
and U10219 (N_10219,N_9007,N_9449);
and U10220 (N_10220,N_9529,N_9622);
or U10221 (N_10221,N_9454,N_9707);
xor U10222 (N_10222,N_9049,N_9239);
nor U10223 (N_10223,N_9110,N_9314);
or U10224 (N_10224,N_9678,N_9442);
nor U10225 (N_10225,N_9608,N_9240);
nand U10226 (N_10226,N_9180,N_9671);
nand U10227 (N_10227,N_9658,N_9260);
and U10228 (N_10228,N_9116,N_9390);
nand U10229 (N_10229,N_9739,N_9369);
nand U10230 (N_10230,N_9035,N_9705);
nor U10231 (N_10231,N_9427,N_9334);
nand U10232 (N_10232,N_9696,N_9090);
and U10233 (N_10233,N_9598,N_9140);
or U10234 (N_10234,N_9367,N_9668);
or U10235 (N_10235,N_9362,N_9160);
or U10236 (N_10236,N_9666,N_9684);
or U10237 (N_10237,N_9511,N_9318);
nand U10238 (N_10238,N_9218,N_9047);
or U10239 (N_10239,N_9068,N_9010);
nand U10240 (N_10240,N_9642,N_9036);
nor U10241 (N_10241,N_9145,N_9500);
nor U10242 (N_10242,N_9434,N_9301);
xnor U10243 (N_10243,N_9577,N_9638);
xnor U10244 (N_10244,N_9649,N_9016);
nor U10245 (N_10245,N_9086,N_9101);
nand U10246 (N_10246,N_9513,N_9437);
and U10247 (N_10247,N_9722,N_9221);
xnor U10248 (N_10248,N_9591,N_9427);
xnor U10249 (N_10249,N_9663,N_9145);
nand U10250 (N_10250,N_9732,N_9047);
xor U10251 (N_10251,N_9438,N_9739);
nand U10252 (N_10252,N_9181,N_9229);
nor U10253 (N_10253,N_9053,N_9202);
or U10254 (N_10254,N_9406,N_9637);
nor U10255 (N_10255,N_9695,N_9730);
and U10256 (N_10256,N_9465,N_9373);
xor U10257 (N_10257,N_9484,N_9718);
and U10258 (N_10258,N_9261,N_9199);
or U10259 (N_10259,N_9134,N_9524);
or U10260 (N_10260,N_9160,N_9690);
and U10261 (N_10261,N_9548,N_9104);
and U10262 (N_10262,N_9445,N_9529);
and U10263 (N_10263,N_9625,N_9551);
and U10264 (N_10264,N_9403,N_9016);
or U10265 (N_10265,N_9730,N_9132);
and U10266 (N_10266,N_9036,N_9543);
and U10267 (N_10267,N_9412,N_9441);
nor U10268 (N_10268,N_9385,N_9096);
nor U10269 (N_10269,N_9001,N_9282);
nand U10270 (N_10270,N_9018,N_9208);
and U10271 (N_10271,N_9584,N_9674);
nor U10272 (N_10272,N_9515,N_9511);
nand U10273 (N_10273,N_9597,N_9025);
or U10274 (N_10274,N_9540,N_9665);
and U10275 (N_10275,N_9706,N_9619);
and U10276 (N_10276,N_9220,N_9490);
xor U10277 (N_10277,N_9041,N_9039);
xnor U10278 (N_10278,N_9469,N_9079);
and U10279 (N_10279,N_9683,N_9729);
nor U10280 (N_10280,N_9620,N_9106);
and U10281 (N_10281,N_9197,N_9423);
nand U10282 (N_10282,N_9104,N_9709);
and U10283 (N_10283,N_9571,N_9101);
xor U10284 (N_10284,N_9199,N_9248);
and U10285 (N_10285,N_9402,N_9505);
and U10286 (N_10286,N_9278,N_9163);
nor U10287 (N_10287,N_9016,N_9488);
nand U10288 (N_10288,N_9486,N_9548);
nor U10289 (N_10289,N_9173,N_9277);
or U10290 (N_10290,N_9560,N_9548);
nor U10291 (N_10291,N_9349,N_9540);
nor U10292 (N_10292,N_9000,N_9049);
xor U10293 (N_10293,N_9607,N_9035);
or U10294 (N_10294,N_9120,N_9075);
nand U10295 (N_10295,N_9557,N_9731);
nor U10296 (N_10296,N_9525,N_9199);
nand U10297 (N_10297,N_9245,N_9511);
nand U10298 (N_10298,N_9051,N_9094);
nand U10299 (N_10299,N_9245,N_9278);
nand U10300 (N_10300,N_9637,N_9287);
and U10301 (N_10301,N_9648,N_9287);
or U10302 (N_10302,N_9485,N_9064);
nand U10303 (N_10303,N_9298,N_9101);
and U10304 (N_10304,N_9450,N_9152);
xnor U10305 (N_10305,N_9027,N_9645);
xnor U10306 (N_10306,N_9399,N_9604);
or U10307 (N_10307,N_9261,N_9444);
nor U10308 (N_10308,N_9119,N_9081);
and U10309 (N_10309,N_9656,N_9452);
xnor U10310 (N_10310,N_9170,N_9240);
nand U10311 (N_10311,N_9690,N_9261);
nand U10312 (N_10312,N_9566,N_9716);
xnor U10313 (N_10313,N_9319,N_9162);
or U10314 (N_10314,N_9673,N_9642);
nand U10315 (N_10315,N_9532,N_9531);
and U10316 (N_10316,N_9661,N_9660);
and U10317 (N_10317,N_9350,N_9215);
nand U10318 (N_10318,N_9197,N_9595);
nand U10319 (N_10319,N_9539,N_9734);
nor U10320 (N_10320,N_9710,N_9233);
nor U10321 (N_10321,N_9000,N_9203);
nand U10322 (N_10322,N_9315,N_9144);
nand U10323 (N_10323,N_9574,N_9707);
nor U10324 (N_10324,N_9243,N_9101);
nand U10325 (N_10325,N_9060,N_9368);
and U10326 (N_10326,N_9119,N_9661);
nand U10327 (N_10327,N_9164,N_9557);
nand U10328 (N_10328,N_9678,N_9454);
and U10329 (N_10329,N_9747,N_9353);
or U10330 (N_10330,N_9052,N_9420);
or U10331 (N_10331,N_9435,N_9387);
and U10332 (N_10332,N_9717,N_9023);
nor U10333 (N_10333,N_9590,N_9441);
nand U10334 (N_10334,N_9103,N_9109);
nand U10335 (N_10335,N_9748,N_9167);
nand U10336 (N_10336,N_9542,N_9657);
nor U10337 (N_10337,N_9039,N_9008);
xor U10338 (N_10338,N_9659,N_9578);
nand U10339 (N_10339,N_9322,N_9634);
or U10340 (N_10340,N_9127,N_9399);
or U10341 (N_10341,N_9578,N_9542);
and U10342 (N_10342,N_9652,N_9087);
nor U10343 (N_10343,N_9016,N_9056);
nand U10344 (N_10344,N_9138,N_9471);
and U10345 (N_10345,N_9295,N_9616);
or U10346 (N_10346,N_9341,N_9009);
nand U10347 (N_10347,N_9375,N_9683);
nand U10348 (N_10348,N_9308,N_9661);
and U10349 (N_10349,N_9251,N_9204);
nor U10350 (N_10350,N_9741,N_9158);
or U10351 (N_10351,N_9498,N_9602);
or U10352 (N_10352,N_9370,N_9404);
or U10353 (N_10353,N_9423,N_9478);
nor U10354 (N_10354,N_9421,N_9320);
or U10355 (N_10355,N_9133,N_9167);
xnor U10356 (N_10356,N_9411,N_9564);
nand U10357 (N_10357,N_9456,N_9419);
and U10358 (N_10358,N_9387,N_9218);
or U10359 (N_10359,N_9074,N_9542);
and U10360 (N_10360,N_9610,N_9663);
xnor U10361 (N_10361,N_9219,N_9409);
nand U10362 (N_10362,N_9109,N_9570);
nor U10363 (N_10363,N_9300,N_9095);
or U10364 (N_10364,N_9575,N_9476);
or U10365 (N_10365,N_9117,N_9329);
and U10366 (N_10366,N_9427,N_9671);
nand U10367 (N_10367,N_9694,N_9335);
and U10368 (N_10368,N_9012,N_9691);
and U10369 (N_10369,N_9214,N_9561);
or U10370 (N_10370,N_9581,N_9045);
nor U10371 (N_10371,N_9519,N_9024);
nor U10372 (N_10372,N_9389,N_9446);
nor U10373 (N_10373,N_9209,N_9076);
nor U10374 (N_10374,N_9071,N_9022);
nand U10375 (N_10375,N_9338,N_9359);
nor U10376 (N_10376,N_9505,N_9142);
nor U10377 (N_10377,N_9075,N_9497);
or U10378 (N_10378,N_9601,N_9002);
nand U10379 (N_10379,N_9628,N_9156);
and U10380 (N_10380,N_9297,N_9686);
and U10381 (N_10381,N_9598,N_9720);
or U10382 (N_10382,N_9720,N_9481);
nand U10383 (N_10383,N_9398,N_9594);
xor U10384 (N_10384,N_9739,N_9145);
and U10385 (N_10385,N_9740,N_9610);
nand U10386 (N_10386,N_9080,N_9315);
or U10387 (N_10387,N_9264,N_9194);
or U10388 (N_10388,N_9702,N_9103);
or U10389 (N_10389,N_9281,N_9079);
and U10390 (N_10390,N_9338,N_9315);
or U10391 (N_10391,N_9048,N_9324);
nor U10392 (N_10392,N_9177,N_9356);
and U10393 (N_10393,N_9643,N_9305);
xor U10394 (N_10394,N_9616,N_9204);
and U10395 (N_10395,N_9561,N_9648);
nor U10396 (N_10396,N_9405,N_9409);
and U10397 (N_10397,N_9448,N_9665);
and U10398 (N_10398,N_9428,N_9172);
and U10399 (N_10399,N_9009,N_9498);
and U10400 (N_10400,N_9305,N_9160);
xnor U10401 (N_10401,N_9356,N_9322);
and U10402 (N_10402,N_9590,N_9450);
or U10403 (N_10403,N_9694,N_9043);
nor U10404 (N_10404,N_9272,N_9445);
nand U10405 (N_10405,N_9361,N_9007);
or U10406 (N_10406,N_9485,N_9670);
nor U10407 (N_10407,N_9553,N_9244);
and U10408 (N_10408,N_9534,N_9653);
or U10409 (N_10409,N_9392,N_9277);
or U10410 (N_10410,N_9204,N_9141);
nor U10411 (N_10411,N_9492,N_9577);
nand U10412 (N_10412,N_9405,N_9506);
or U10413 (N_10413,N_9201,N_9486);
xor U10414 (N_10414,N_9533,N_9579);
or U10415 (N_10415,N_9250,N_9246);
nand U10416 (N_10416,N_9426,N_9571);
or U10417 (N_10417,N_9509,N_9522);
or U10418 (N_10418,N_9584,N_9687);
or U10419 (N_10419,N_9487,N_9721);
nand U10420 (N_10420,N_9476,N_9182);
nor U10421 (N_10421,N_9023,N_9471);
nor U10422 (N_10422,N_9638,N_9140);
and U10423 (N_10423,N_9530,N_9702);
nor U10424 (N_10424,N_9706,N_9488);
or U10425 (N_10425,N_9460,N_9032);
nand U10426 (N_10426,N_9535,N_9577);
or U10427 (N_10427,N_9497,N_9018);
nor U10428 (N_10428,N_9279,N_9515);
nor U10429 (N_10429,N_9034,N_9529);
xor U10430 (N_10430,N_9330,N_9396);
nand U10431 (N_10431,N_9340,N_9105);
and U10432 (N_10432,N_9161,N_9251);
nor U10433 (N_10433,N_9218,N_9300);
and U10434 (N_10434,N_9632,N_9425);
nand U10435 (N_10435,N_9702,N_9001);
nand U10436 (N_10436,N_9336,N_9028);
nand U10437 (N_10437,N_9334,N_9027);
and U10438 (N_10438,N_9582,N_9614);
nand U10439 (N_10439,N_9542,N_9064);
and U10440 (N_10440,N_9134,N_9502);
nand U10441 (N_10441,N_9066,N_9587);
nand U10442 (N_10442,N_9281,N_9608);
and U10443 (N_10443,N_9426,N_9067);
or U10444 (N_10444,N_9494,N_9060);
nor U10445 (N_10445,N_9221,N_9691);
nand U10446 (N_10446,N_9383,N_9272);
and U10447 (N_10447,N_9565,N_9389);
nor U10448 (N_10448,N_9307,N_9064);
nor U10449 (N_10449,N_9598,N_9445);
and U10450 (N_10450,N_9690,N_9510);
xnor U10451 (N_10451,N_9254,N_9068);
or U10452 (N_10452,N_9120,N_9257);
and U10453 (N_10453,N_9532,N_9521);
or U10454 (N_10454,N_9285,N_9699);
and U10455 (N_10455,N_9560,N_9397);
or U10456 (N_10456,N_9743,N_9252);
nand U10457 (N_10457,N_9227,N_9234);
and U10458 (N_10458,N_9407,N_9648);
or U10459 (N_10459,N_9268,N_9511);
and U10460 (N_10460,N_9568,N_9646);
or U10461 (N_10461,N_9173,N_9342);
nand U10462 (N_10462,N_9189,N_9370);
and U10463 (N_10463,N_9584,N_9486);
nor U10464 (N_10464,N_9060,N_9446);
nor U10465 (N_10465,N_9440,N_9400);
or U10466 (N_10466,N_9188,N_9478);
and U10467 (N_10467,N_9555,N_9106);
or U10468 (N_10468,N_9538,N_9700);
nand U10469 (N_10469,N_9054,N_9253);
xnor U10470 (N_10470,N_9127,N_9077);
nor U10471 (N_10471,N_9081,N_9300);
nor U10472 (N_10472,N_9748,N_9742);
nor U10473 (N_10473,N_9559,N_9667);
nand U10474 (N_10474,N_9345,N_9506);
nand U10475 (N_10475,N_9051,N_9098);
and U10476 (N_10476,N_9300,N_9674);
or U10477 (N_10477,N_9642,N_9132);
nand U10478 (N_10478,N_9545,N_9513);
nor U10479 (N_10479,N_9023,N_9443);
xnor U10480 (N_10480,N_9455,N_9388);
nand U10481 (N_10481,N_9316,N_9614);
nand U10482 (N_10482,N_9082,N_9350);
nor U10483 (N_10483,N_9538,N_9455);
and U10484 (N_10484,N_9136,N_9227);
nor U10485 (N_10485,N_9407,N_9118);
xor U10486 (N_10486,N_9436,N_9019);
and U10487 (N_10487,N_9350,N_9588);
nand U10488 (N_10488,N_9645,N_9066);
and U10489 (N_10489,N_9147,N_9534);
nand U10490 (N_10490,N_9408,N_9156);
or U10491 (N_10491,N_9049,N_9416);
xnor U10492 (N_10492,N_9194,N_9564);
xor U10493 (N_10493,N_9394,N_9031);
nand U10494 (N_10494,N_9528,N_9688);
or U10495 (N_10495,N_9137,N_9048);
nand U10496 (N_10496,N_9738,N_9054);
nand U10497 (N_10497,N_9331,N_9065);
nand U10498 (N_10498,N_9260,N_9414);
nand U10499 (N_10499,N_9521,N_9382);
xnor U10500 (N_10500,N_9823,N_10415);
or U10501 (N_10501,N_10290,N_10391);
and U10502 (N_10502,N_9907,N_10017);
nand U10503 (N_10503,N_10354,N_10154);
nor U10504 (N_10504,N_9860,N_10029);
and U10505 (N_10505,N_9792,N_10034);
nor U10506 (N_10506,N_9958,N_9906);
or U10507 (N_10507,N_10148,N_9764);
nand U10508 (N_10508,N_10123,N_10045);
xor U10509 (N_10509,N_10485,N_10367);
nor U10510 (N_10510,N_10112,N_9867);
and U10511 (N_10511,N_10206,N_10442);
xor U10512 (N_10512,N_10271,N_10159);
or U10513 (N_10513,N_9911,N_10357);
nand U10514 (N_10514,N_10014,N_10342);
and U10515 (N_10515,N_10224,N_10220);
xor U10516 (N_10516,N_10050,N_9847);
nor U10517 (N_10517,N_10347,N_10333);
nor U10518 (N_10518,N_10022,N_9924);
or U10519 (N_10519,N_10261,N_10423);
or U10520 (N_10520,N_10132,N_10096);
and U10521 (N_10521,N_10279,N_10173);
or U10522 (N_10522,N_10008,N_9772);
nor U10523 (N_10523,N_10340,N_9771);
nor U10524 (N_10524,N_10293,N_10169);
and U10525 (N_10525,N_9954,N_10153);
nor U10526 (N_10526,N_10401,N_9796);
xor U10527 (N_10527,N_9755,N_10002);
nor U10528 (N_10528,N_10098,N_9839);
and U10529 (N_10529,N_10052,N_9935);
xnor U10530 (N_10530,N_9899,N_9926);
nor U10531 (N_10531,N_10370,N_10270);
nor U10532 (N_10532,N_10300,N_10193);
nand U10533 (N_10533,N_10111,N_9840);
nand U10534 (N_10534,N_9876,N_10468);
nand U10535 (N_10535,N_9993,N_10072);
xnor U10536 (N_10536,N_10127,N_10387);
and U10537 (N_10537,N_10479,N_10419);
nand U10538 (N_10538,N_10021,N_9846);
and U10539 (N_10539,N_9952,N_10144);
nand U10540 (N_10540,N_9870,N_10283);
nor U10541 (N_10541,N_9830,N_10495);
xnor U10542 (N_10542,N_10336,N_10307);
or U10543 (N_10543,N_10023,N_10103);
xor U10544 (N_10544,N_10164,N_10094);
xor U10545 (N_10545,N_10025,N_10348);
and U10546 (N_10546,N_10202,N_10126);
and U10547 (N_10547,N_9941,N_10332);
or U10548 (N_10548,N_10092,N_10260);
nor U10549 (N_10549,N_10185,N_9841);
nor U10550 (N_10550,N_10305,N_9939);
or U10551 (N_10551,N_10309,N_10124);
or U10552 (N_10552,N_10175,N_10047);
and U10553 (N_10553,N_10128,N_10301);
nand U10554 (N_10554,N_10219,N_9797);
nor U10555 (N_10555,N_9916,N_10470);
nand U10556 (N_10556,N_9799,N_10440);
nor U10557 (N_10557,N_10484,N_9866);
nor U10558 (N_10558,N_9963,N_10026);
nor U10559 (N_10559,N_10188,N_10337);
nor U10560 (N_10560,N_10353,N_10061);
nor U10561 (N_10561,N_10156,N_9855);
and U10562 (N_10562,N_10000,N_9931);
nand U10563 (N_10563,N_10344,N_9971);
and U10564 (N_10564,N_10257,N_10091);
nand U10565 (N_10565,N_10474,N_10068);
or U10566 (N_10566,N_10100,N_10447);
or U10567 (N_10567,N_9765,N_9854);
nand U10568 (N_10568,N_9877,N_10041);
or U10569 (N_10569,N_9978,N_10011);
and U10570 (N_10570,N_9972,N_9888);
and U10571 (N_10571,N_10432,N_9836);
xor U10572 (N_10572,N_10198,N_9992);
nand U10573 (N_10573,N_9933,N_10411);
nand U10574 (N_10574,N_10480,N_10295);
nand U10575 (N_10575,N_10358,N_10325);
nand U10576 (N_10576,N_10276,N_10245);
nand U10577 (N_10577,N_10491,N_10174);
or U10578 (N_10578,N_10109,N_9957);
nor U10579 (N_10579,N_10006,N_10472);
or U10580 (N_10580,N_10161,N_10125);
and U10581 (N_10581,N_10272,N_10339);
nor U10582 (N_10582,N_9842,N_10262);
and U10583 (N_10583,N_10248,N_9912);
nand U10584 (N_10584,N_9998,N_10298);
nand U10585 (N_10585,N_9778,N_10375);
and U10586 (N_10586,N_9761,N_9875);
or U10587 (N_10587,N_10143,N_10464);
or U10588 (N_10588,N_9955,N_10314);
xnor U10589 (N_10589,N_9790,N_10388);
and U10590 (N_10590,N_10190,N_10294);
and U10591 (N_10591,N_10253,N_9983);
or U10592 (N_10592,N_10494,N_9930);
or U10593 (N_10593,N_10089,N_10121);
or U10594 (N_10594,N_10256,N_10117);
and U10595 (N_10595,N_10114,N_10330);
or U10596 (N_10596,N_10238,N_10379);
nor U10597 (N_10597,N_10386,N_10216);
nor U10598 (N_10598,N_10497,N_10405);
nor U10599 (N_10599,N_10394,N_10268);
nor U10600 (N_10600,N_10247,N_10212);
or U10601 (N_10601,N_9902,N_9780);
nor U10602 (N_10602,N_10054,N_10278);
nand U10603 (N_10603,N_10095,N_10493);
or U10604 (N_10604,N_9945,N_9980);
nor U10605 (N_10605,N_10383,N_10194);
and U10606 (N_10606,N_10304,N_9757);
and U10607 (N_10607,N_10178,N_9759);
nand U10608 (N_10608,N_10044,N_9834);
nor U10609 (N_10609,N_9921,N_9874);
nor U10610 (N_10610,N_10399,N_10449);
or U10611 (N_10611,N_9868,N_10032);
nor U10612 (N_10612,N_9758,N_10016);
xor U10613 (N_10613,N_9903,N_10018);
and U10614 (N_10614,N_9787,N_9970);
nor U10615 (N_10615,N_9934,N_10077);
nand U10616 (N_10616,N_10404,N_9756);
xnor U10617 (N_10617,N_10088,N_10019);
and U10618 (N_10618,N_10452,N_9813);
nor U10619 (N_10619,N_10020,N_10312);
nand U10620 (N_10620,N_9820,N_10446);
or U10621 (N_10621,N_9807,N_10122);
and U10622 (N_10622,N_9962,N_10141);
and U10623 (N_10623,N_10181,N_10180);
nand U10624 (N_10624,N_10350,N_9959);
or U10625 (N_10625,N_10250,N_10208);
nor U10626 (N_10626,N_10297,N_10177);
nor U10627 (N_10627,N_9995,N_10302);
or U10628 (N_10628,N_9750,N_9785);
and U10629 (N_10629,N_10074,N_10051);
xnor U10630 (N_10630,N_10010,N_9946);
nor U10631 (N_10631,N_10036,N_10139);
nand U10632 (N_10632,N_10361,N_10073);
xor U10633 (N_10633,N_10443,N_10269);
or U10634 (N_10634,N_9852,N_9897);
and U10635 (N_10635,N_10385,N_10459);
xor U10636 (N_10636,N_10013,N_9811);
nand U10637 (N_10637,N_9783,N_10078);
or U10638 (N_10638,N_9966,N_10274);
xnor U10639 (N_10639,N_10456,N_9975);
or U10640 (N_10640,N_9753,N_10263);
nor U10641 (N_10641,N_10498,N_10430);
nor U10642 (N_10642,N_10346,N_10137);
and U10643 (N_10643,N_10113,N_10012);
nand U10644 (N_10644,N_10209,N_10280);
and U10645 (N_10645,N_10064,N_10338);
xnor U10646 (N_10646,N_10203,N_10267);
xnor U10647 (N_10647,N_10049,N_10395);
and U10648 (N_10648,N_10106,N_9828);
xor U10649 (N_10649,N_9843,N_9893);
nor U10650 (N_10650,N_10053,N_10058);
and U10651 (N_10651,N_9894,N_9887);
nor U10652 (N_10652,N_9968,N_10412);
nand U10653 (N_10653,N_10378,N_9806);
or U10654 (N_10654,N_10351,N_10421);
and U10655 (N_10655,N_9999,N_9858);
nand U10656 (N_10656,N_9965,N_10093);
xor U10657 (N_10657,N_10402,N_9918);
or U10658 (N_10658,N_10184,N_10217);
or U10659 (N_10659,N_10223,N_9956);
nand U10660 (N_10660,N_10226,N_10075);
or U10661 (N_10661,N_10368,N_9949);
and U10662 (N_10662,N_10063,N_9851);
nand U10663 (N_10663,N_10135,N_10056);
or U10664 (N_10664,N_10225,N_9832);
nor U10665 (N_10665,N_10249,N_9985);
nor U10666 (N_10666,N_10234,N_10084);
or U10667 (N_10667,N_9882,N_10176);
or U10668 (N_10668,N_9929,N_10145);
nor U10669 (N_10669,N_9950,N_10197);
and U10670 (N_10670,N_10436,N_10062);
and U10671 (N_10671,N_10237,N_10398);
and U10672 (N_10672,N_10211,N_10060);
and U10673 (N_10673,N_10318,N_10487);
nor U10674 (N_10674,N_10321,N_9768);
xnor U10675 (N_10675,N_9879,N_10201);
nor U10676 (N_10676,N_9896,N_9873);
nor U10677 (N_10677,N_10119,N_9831);
and U10678 (N_10678,N_10129,N_9908);
nand U10679 (N_10679,N_9937,N_10258);
nor U10680 (N_10680,N_10373,N_10408);
xor U10681 (N_10681,N_10489,N_9816);
and U10682 (N_10682,N_10067,N_10458);
or U10683 (N_10683,N_9845,N_10384);
nor U10684 (N_10684,N_10429,N_9850);
nor U10685 (N_10685,N_9793,N_9782);
and U10686 (N_10686,N_9981,N_10273);
nor U10687 (N_10687,N_10200,N_10087);
nor U10688 (N_10688,N_10229,N_10133);
or U10689 (N_10689,N_10120,N_9789);
nand U10690 (N_10690,N_10031,N_10365);
nor U10691 (N_10691,N_9984,N_10228);
and U10692 (N_10692,N_10242,N_10310);
and U10693 (N_10693,N_9862,N_10439);
and U10694 (N_10694,N_10005,N_10140);
nor U10695 (N_10695,N_9751,N_9794);
and U10696 (N_10696,N_10231,N_10170);
and U10697 (N_10697,N_9996,N_9821);
nand U10698 (N_10698,N_9986,N_10469);
xnor U10699 (N_10699,N_10186,N_10210);
and U10700 (N_10700,N_10167,N_10035);
or U10701 (N_10701,N_10326,N_10065);
nor U10702 (N_10702,N_10289,N_10466);
nand U10703 (N_10703,N_10311,N_9943);
and U10704 (N_10704,N_10213,N_10414);
or U10705 (N_10705,N_9967,N_9809);
and U10706 (N_10706,N_10406,N_9767);
nor U10707 (N_10707,N_9754,N_9878);
nor U10708 (N_10708,N_9788,N_9923);
nor U10709 (N_10709,N_10028,N_9914);
and U10710 (N_10710,N_10199,N_9863);
nand U10711 (N_10711,N_10003,N_10254);
nand U10712 (N_10712,N_9779,N_10196);
nor U10713 (N_10713,N_9776,N_9936);
nor U10714 (N_10714,N_9786,N_10130);
and U10715 (N_10715,N_9824,N_10157);
nand U10716 (N_10716,N_9803,N_9762);
and U10717 (N_10717,N_10434,N_9990);
and U10718 (N_10718,N_9770,N_10343);
or U10719 (N_10719,N_10291,N_10460);
nand U10720 (N_10720,N_10481,N_10080);
nand U10721 (N_10721,N_10259,N_10235);
nand U10722 (N_10722,N_10475,N_10163);
xnor U10723 (N_10723,N_10150,N_10371);
nand U10724 (N_10724,N_9915,N_10187);
and U10725 (N_10725,N_10451,N_10090);
or U10726 (N_10726,N_10376,N_10482);
and U10727 (N_10727,N_10478,N_10264);
or U10728 (N_10728,N_10457,N_10461);
or U10729 (N_10729,N_9976,N_10407);
nand U10730 (N_10730,N_9883,N_9837);
nand U10731 (N_10731,N_9818,N_10319);
and U10732 (N_10732,N_10382,N_10366);
and U10733 (N_10733,N_10349,N_9919);
or U10734 (N_10734,N_9977,N_9808);
xor U10735 (N_10735,N_10277,N_10400);
xor U10736 (N_10736,N_10374,N_10313);
nor U10737 (N_10737,N_10476,N_10204);
nor U10738 (N_10738,N_9922,N_9861);
and U10739 (N_10739,N_10168,N_9829);
nand U10740 (N_10740,N_10038,N_10115);
or U10741 (N_10741,N_10102,N_10138);
or U10742 (N_10742,N_10059,N_10046);
and U10743 (N_10743,N_10299,N_9835);
nor U10744 (N_10744,N_10246,N_10403);
nand U10745 (N_10745,N_10205,N_10207);
xor U10746 (N_10746,N_10425,N_9784);
and U10747 (N_10747,N_10191,N_10147);
nor U10748 (N_10748,N_10473,N_10316);
and U10749 (N_10749,N_10490,N_10004);
nor U10750 (N_10750,N_9880,N_10409);
nand U10751 (N_10751,N_9856,N_10435);
nor U10752 (N_10752,N_9760,N_10037);
or U10753 (N_10753,N_10364,N_10255);
nand U10754 (N_10754,N_9920,N_10463);
nand U10755 (N_10755,N_10438,N_9942);
nor U10756 (N_10756,N_10030,N_10331);
nor U10757 (N_10757,N_9815,N_10431);
nand U10758 (N_10758,N_10007,N_10303);
or U10759 (N_10759,N_9827,N_10134);
or U10760 (N_10760,N_10467,N_9951);
or U10761 (N_10761,N_10081,N_10445);
nand U10762 (N_10762,N_10043,N_9795);
and U10763 (N_10763,N_10486,N_9865);
nand U10764 (N_10764,N_9889,N_10107);
or U10765 (N_10765,N_10101,N_9801);
nor U10766 (N_10766,N_10162,N_9844);
nand U10767 (N_10767,N_10413,N_9775);
nor U10768 (N_10768,N_10306,N_9773);
nor U10769 (N_10769,N_9777,N_10397);
nor U10770 (N_10770,N_10057,N_9913);
xnor U10771 (N_10771,N_9871,N_10070);
or U10772 (N_10772,N_10099,N_10104);
and U10773 (N_10773,N_10221,N_9890);
nand U10774 (N_10774,N_10182,N_9961);
nand U10775 (N_10775,N_9812,N_9940);
and U10776 (N_10776,N_9987,N_9769);
or U10777 (N_10777,N_10142,N_9800);
xor U10778 (N_10778,N_10239,N_10243);
nor U10779 (N_10779,N_9960,N_10069);
nor U10780 (N_10780,N_9798,N_9989);
or U10781 (N_10781,N_10322,N_10222);
and U10782 (N_10782,N_10418,N_10389);
or U10783 (N_10783,N_10040,N_9932);
nand U10784 (N_10784,N_9825,N_10252);
nor U10785 (N_10785,N_9763,N_10377);
nand U10786 (N_10786,N_10359,N_10328);
or U10787 (N_10787,N_10426,N_10172);
nand U10788 (N_10788,N_10288,N_10158);
and U10789 (N_10789,N_9822,N_10136);
xor U10790 (N_10790,N_10323,N_10183);
nand U10791 (N_10791,N_9859,N_10317);
nand U10792 (N_10792,N_10227,N_10083);
nand U10793 (N_10793,N_10362,N_10232);
or U10794 (N_10794,N_10393,N_10450);
or U10795 (N_10795,N_10082,N_9791);
nand U10796 (N_10796,N_10085,N_9857);
nor U10797 (N_10797,N_9781,N_10455);
xnor U10798 (N_10798,N_10009,N_9994);
and U10799 (N_10799,N_10496,N_10492);
nor U10800 (N_10800,N_9814,N_9938);
and U10801 (N_10801,N_10427,N_10390);
nor U10802 (N_10802,N_10499,N_9927);
nor U10803 (N_10803,N_10422,N_10275);
nand U10804 (N_10804,N_10477,N_10024);
and U10805 (N_10805,N_10355,N_10352);
nor U10806 (N_10806,N_10441,N_10166);
nor U10807 (N_10807,N_10152,N_10381);
nor U10808 (N_10808,N_9853,N_10327);
nand U10809 (N_10809,N_10287,N_10066);
xnor U10810 (N_10810,N_9953,N_10392);
and U10811 (N_10811,N_10146,N_9869);
nand U10812 (N_10812,N_9805,N_9925);
nor U10813 (N_10813,N_9895,N_10097);
and U10814 (N_10814,N_10039,N_10195);
and U10815 (N_10815,N_9838,N_10448);
nand U10816 (N_10816,N_10233,N_10462);
nor U10817 (N_10817,N_9982,N_10110);
nand U10818 (N_10818,N_9804,N_10433);
or U10819 (N_10819,N_9802,N_9944);
nand U10820 (N_10820,N_10165,N_10428);
xor U10821 (N_10821,N_9752,N_10179);
or U10822 (N_10822,N_10315,N_10324);
or U10823 (N_10823,N_9886,N_10214);
and U10824 (N_10824,N_10192,N_10266);
nand U10825 (N_10825,N_10241,N_10380);
nor U10826 (N_10826,N_10437,N_10453);
or U10827 (N_10827,N_10396,N_10282);
or U10828 (N_10828,N_10076,N_9892);
nand U10829 (N_10829,N_9928,N_9898);
nand U10830 (N_10830,N_10015,N_10244);
nor U10831 (N_10831,N_9904,N_10345);
xor U10832 (N_10832,N_9833,N_10483);
and U10833 (N_10833,N_9881,N_9891);
and U10834 (N_10834,N_9900,N_9969);
nor U10835 (N_10835,N_10329,N_9948);
and U10836 (N_10836,N_10218,N_9901);
nand U10837 (N_10837,N_9974,N_10420);
or U10838 (N_10838,N_10471,N_10251);
nand U10839 (N_10839,N_10369,N_10160);
and U10840 (N_10840,N_10334,N_10055);
nor U10841 (N_10841,N_10001,N_10488);
nand U10842 (N_10842,N_10189,N_10308);
xnor U10843 (N_10843,N_9997,N_10410);
and U10844 (N_10844,N_10285,N_10292);
nor U10845 (N_10845,N_10149,N_10424);
and U10846 (N_10846,N_10240,N_10363);
nand U10847 (N_10847,N_10108,N_10116);
nor U10848 (N_10848,N_9917,N_9817);
nor U10849 (N_10849,N_10230,N_10118);
and U10850 (N_10850,N_9973,N_9864);
or U10851 (N_10851,N_10042,N_10444);
nand U10852 (N_10852,N_10027,N_10171);
nor U10853 (N_10853,N_10465,N_10417);
nand U10854 (N_10854,N_10360,N_9884);
or U10855 (N_10855,N_9947,N_9848);
or U10856 (N_10856,N_10372,N_10071);
nand U10857 (N_10857,N_10215,N_9885);
nor U10858 (N_10858,N_10335,N_10236);
and U10859 (N_10859,N_9910,N_10033);
nor U10860 (N_10860,N_10086,N_9979);
and U10861 (N_10861,N_10105,N_9810);
nand U10862 (N_10862,N_9819,N_9909);
and U10863 (N_10863,N_9991,N_10284);
and U10864 (N_10864,N_9872,N_10286);
or U10865 (N_10865,N_10151,N_10265);
or U10866 (N_10866,N_10296,N_10454);
or U10867 (N_10867,N_10356,N_10079);
nor U10868 (N_10868,N_9988,N_9826);
nand U10869 (N_10869,N_10341,N_10048);
or U10870 (N_10870,N_9905,N_10281);
nand U10871 (N_10871,N_10155,N_9964);
nand U10872 (N_10872,N_9849,N_9774);
xnor U10873 (N_10873,N_10131,N_9766);
nand U10874 (N_10874,N_10416,N_10320);
or U10875 (N_10875,N_9979,N_10016);
and U10876 (N_10876,N_10218,N_10392);
or U10877 (N_10877,N_9954,N_10097);
and U10878 (N_10878,N_9954,N_10326);
and U10879 (N_10879,N_10072,N_9750);
and U10880 (N_10880,N_10231,N_10328);
or U10881 (N_10881,N_9869,N_9887);
and U10882 (N_10882,N_10089,N_10027);
nand U10883 (N_10883,N_9827,N_10245);
xnor U10884 (N_10884,N_10178,N_9783);
xnor U10885 (N_10885,N_10220,N_9981);
or U10886 (N_10886,N_10355,N_10046);
nor U10887 (N_10887,N_10161,N_10406);
nor U10888 (N_10888,N_10087,N_10049);
or U10889 (N_10889,N_10473,N_10281);
and U10890 (N_10890,N_10458,N_9934);
and U10891 (N_10891,N_9999,N_10018);
or U10892 (N_10892,N_10022,N_10410);
or U10893 (N_10893,N_10103,N_10212);
nand U10894 (N_10894,N_9767,N_9878);
nand U10895 (N_10895,N_9783,N_10256);
nand U10896 (N_10896,N_9869,N_10347);
or U10897 (N_10897,N_9863,N_9751);
or U10898 (N_10898,N_10018,N_10056);
nor U10899 (N_10899,N_10132,N_9865);
nor U10900 (N_10900,N_10425,N_9973);
nor U10901 (N_10901,N_10305,N_10147);
or U10902 (N_10902,N_10229,N_9946);
nand U10903 (N_10903,N_10393,N_10279);
nand U10904 (N_10904,N_10471,N_10479);
and U10905 (N_10905,N_9851,N_10058);
nand U10906 (N_10906,N_9885,N_9869);
nand U10907 (N_10907,N_9982,N_10286);
or U10908 (N_10908,N_10219,N_9850);
nor U10909 (N_10909,N_9912,N_9762);
or U10910 (N_10910,N_9905,N_9833);
nor U10911 (N_10911,N_9915,N_10180);
nand U10912 (N_10912,N_10271,N_10304);
and U10913 (N_10913,N_9750,N_10418);
nand U10914 (N_10914,N_9805,N_10194);
nor U10915 (N_10915,N_9769,N_9960);
nand U10916 (N_10916,N_10007,N_9868);
nor U10917 (N_10917,N_10441,N_10075);
nor U10918 (N_10918,N_10342,N_10179);
nor U10919 (N_10919,N_9946,N_10422);
xnor U10920 (N_10920,N_9900,N_9820);
or U10921 (N_10921,N_10265,N_10005);
and U10922 (N_10922,N_9757,N_9812);
nor U10923 (N_10923,N_9764,N_10437);
nor U10924 (N_10924,N_9841,N_10174);
xor U10925 (N_10925,N_10071,N_10438);
or U10926 (N_10926,N_10135,N_10371);
or U10927 (N_10927,N_9789,N_10369);
xnor U10928 (N_10928,N_10110,N_9797);
or U10929 (N_10929,N_10443,N_10455);
and U10930 (N_10930,N_9994,N_9932);
nand U10931 (N_10931,N_10258,N_9994);
or U10932 (N_10932,N_10143,N_10026);
xor U10933 (N_10933,N_10114,N_10245);
nand U10934 (N_10934,N_10286,N_9842);
and U10935 (N_10935,N_9840,N_9862);
nand U10936 (N_10936,N_10235,N_10163);
or U10937 (N_10937,N_10420,N_9802);
nor U10938 (N_10938,N_10364,N_9814);
or U10939 (N_10939,N_10180,N_9893);
nor U10940 (N_10940,N_9970,N_9756);
nor U10941 (N_10941,N_10309,N_10111);
and U10942 (N_10942,N_9870,N_9885);
and U10943 (N_10943,N_10107,N_10460);
nand U10944 (N_10944,N_10071,N_9789);
xnor U10945 (N_10945,N_10224,N_10035);
nand U10946 (N_10946,N_10177,N_10068);
xnor U10947 (N_10947,N_9873,N_9979);
nand U10948 (N_10948,N_10082,N_9981);
nand U10949 (N_10949,N_10440,N_10392);
nand U10950 (N_10950,N_10193,N_10444);
or U10951 (N_10951,N_10237,N_10102);
nor U10952 (N_10952,N_10002,N_10398);
nor U10953 (N_10953,N_10456,N_9946);
nor U10954 (N_10954,N_9906,N_10283);
or U10955 (N_10955,N_10334,N_9770);
nor U10956 (N_10956,N_10346,N_10264);
xnor U10957 (N_10957,N_10371,N_10341);
xor U10958 (N_10958,N_10454,N_9803);
nand U10959 (N_10959,N_10242,N_10312);
nor U10960 (N_10960,N_10432,N_9810);
or U10961 (N_10961,N_10235,N_10455);
nand U10962 (N_10962,N_10307,N_9941);
nand U10963 (N_10963,N_9803,N_10212);
or U10964 (N_10964,N_10437,N_10083);
nand U10965 (N_10965,N_9807,N_10392);
nand U10966 (N_10966,N_10283,N_9806);
nor U10967 (N_10967,N_10186,N_10396);
nand U10968 (N_10968,N_10071,N_10444);
nor U10969 (N_10969,N_10360,N_10395);
or U10970 (N_10970,N_10282,N_9939);
nor U10971 (N_10971,N_9930,N_10397);
nor U10972 (N_10972,N_10068,N_10479);
nor U10973 (N_10973,N_10129,N_10080);
nor U10974 (N_10974,N_9925,N_9797);
or U10975 (N_10975,N_10104,N_10033);
and U10976 (N_10976,N_9802,N_10279);
nor U10977 (N_10977,N_10381,N_9918);
or U10978 (N_10978,N_9838,N_10450);
or U10979 (N_10979,N_9755,N_10203);
nor U10980 (N_10980,N_10432,N_10227);
nor U10981 (N_10981,N_10187,N_10337);
and U10982 (N_10982,N_9872,N_9789);
or U10983 (N_10983,N_10105,N_10216);
nand U10984 (N_10984,N_10092,N_10310);
xnor U10985 (N_10985,N_10098,N_10209);
nor U10986 (N_10986,N_9916,N_10198);
and U10987 (N_10987,N_9962,N_9773);
or U10988 (N_10988,N_9961,N_10118);
or U10989 (N_10989,N_10437,N_9759);
and U10990 (N_10990,N_10255,N_10272);
and U10991 (N_10991,N_10367,N_9922);
xnor U10992 (N_10992,N_9986,N_10420);
nand U10993 (N_10993,N_9921,N_10324);
nand U10994 (N_10994,N_10397,N_9945);
nand U10995 (N_10995,N_10215,N_10403);
and U10996 (N_10996,N_10309,N_9765);
nor U10997 (N_10997,N_9875,N_10436);
nand U10998 (N_10998,N_9759,N_10046);
xnor U10999 (N_10999,N_10168,N_10475);
nor U11000 (N_11000,N_10245,N_10468);
xor U11001 (N_11001,N_10370,N_9908);
or U11002 (N_11002,N_10249,N_10264);
or U11003 (N_11003,N_10335,N_9932);
and U11004 (N_11004,N_10225,N_10373);
or U11005 (N_11005,N_10162,N_9799);
nor U11006 (N_11006,N_10008,N_10253);
xnor U11007 (N_11007,N_10474,N_9843);
or U11008 (N_11008,N_9784,N_9835);
or U11009 (N_11009,N_9993,N_10355);
nor U11010 (N_11010,N_9930,N_9914);
and U11011 (N_11011,N_9926,N_10304);
and U11012 (N_11012,N_9971,N_10153);
nor U11013 (N_11013,N_9950,N_10437);
nor U11014 (N_11014,N_9767,N_10123);
or U11015 (N_11015,N_9989,N_9774);
or U11016 (N_11016,N_10097,N_10375);
or U11017 (N_11017,N_10251,N_10463);
or U11018 (N_11018,N_9874,N_9753);
nand U11019 (N_11019,N_10408,N_9798);
nor U11020 (N_11020,N_10244,N_10462);
nor U11021 (N_11021,N_9985,N_9760);
nand U11022 (N_11022,N_10349,N_10035);
nand U11023 (N_11023,N_9889,N_9752);
nor U11024 (N_11024,N_10276,N_10387);
nor U11025 (N_11025,N_10108,N_10068);
nand U11026 (N_11026,N_10193,N_10131);
or U11027 (N_11027,N_9957,N_10408);
or U11028 (N_11028,N_10168,N_9880);
nor U11029 (N_11029,N_10168,N_9968);
or U11030 (N_11030,N_10071,N_10315);
nand U11031 (N_11031,N_10493,N_10460);
xor U11032 (N_11032,N_10428,N_10150);
and U11033 (N_11033,N_9848,N_9786);
nor U11034 (N_11034,N_9889,N_9899);
or U11035 (N_11035,N_9997,N_10158);
and U11036 (N_11036,N_10473,N_10191);
nor U11037 (N_11037,N_10317,N_9810);
xnor U11038 (N_11038,N_10106,N_9970);
and U11039 (N_11039,N_10377,N_10062);
and U11040 (N_11040,N_9927,N_10079);
nor U11041 (N_11041,N_9771,N_10116);
nand U11042 (N_11042,N_10242,N_10015);
nor U11043 (N_11043,N_10288,N_9822);
and U11044 (N_11044,N_9857,N_9935);
and U11045 (N_11045,N_10349,N_9835);
and U11046 (N_11046,N_10005,N_9931);
nor U11047 (N_11047,N_10445,N_10016);
nand U11048 (N_11048,N_10219,N_10213);
and U11049 (N_11049,N_10348,N_10399);
or U11050 (N_11050,N_10439,N_10278);
nand U11051 (N_11051,N_10328,N_10324);
or U11052 (N_11052,N_9907,N_10074);
and U11053 (N_11053,N_10248,N_10052);
or U11054 (N_11054,N_10335,N_10268);
xor U11055 (N_11055,N_10212,N_10399);
and U11056 (N_11056,N_10210,N_9992);
or U11057 (N_11057,N_9910,N_10232);
and U11058 (N_11058,N_10188,N_9887);
nand U11059 (N_11059,N_10475,N_10060);
nand U11060 (N_11060,N_9857,N_10488);
or U11061 (N_11061,N_10441,N_9780);
or U11062 (N_11062,N_10255,N_10163);
or U11063 (N_11063,N_10056,N_10377);
nand U11064 (N_11064,N_9895,N_10277);
and U11065 (N_11065,N_10098,N_10096);
nand U11066 (N_11066,N_9919,N_10435);
nand U11067 (N_11067,N_10077,N_10125);
and U11068 (N_11068,N_9870,N_10134);
nand U11069 (N_11069,N_10176,N_10384);
nand U11070 (N_11070,N_10141,N_10423);
and U11071 (N_11071,N_9800,N_9795);
nor U11072 (N_11072,N_10020,N_9862);
nor U11073 (N_11073,N_10315,N_10186);
nor U11074 (N_11074,N_10125,N_9775);
nand U11075 (N_11075,N_9798,N_10075);
or U11076 (N_11076,N_10289,N_9897);
nor U11077 (N_11077,N_9780,N_10179);
or U11078 (N_11078,N_10294,N_10027);
nor U11079 (N_11079,N_9830,N_10408);
nand U11080 (N_11080,N_10446,N_10370);
nand U11081 (N_11081,N_10284,N_9907);
nor U11082 (N_11082,N_9757,N_10128);
nor U11083 (N_11083,N_10216,N_10424);
nor U11084 (N_11084,N_10052,N_10258);
nor U11085 (N_11085,N_10289,N_10003);
nor U11086 (N_11086,N_9926,N_10084);
and U11087 (N_11087,N_10189,N_9870);
and U11088 (N_11088,N_10001,N_9927);
xnor U11089 (N_11089,N_10395,N_9825);
or U11090 (N_11090,N_10399,N_10339);
or U11091 (N_11091,N_10376,N_10430);
and U11092 (N_11092,N_10468,N_9792);
or U11093 (N_11093,N_10036,N_9807);
and U11094 (N_11094,N_9892,N_9766);
and U11095 (N_11095,N_10306,N_10222);
nand U11096 (N_11096,N_10177,N_10390);
or U11097 (N_11097,N_10389,N_10303);
or U11098 (N_11098,N_10184,N_10404);
or U11099 (N_11099,N_10188,N_10079);
or U11100 (N_11100,N_10481,N_9971);
and U11101 (N_11101,N_10398,N_9873);
and U11102 (N_11102,N_10370,N_10241);
nand U11103 (N_11103,N_10045,N_9954);
nor U11104 (N_11104,N_10000,N_10298);
nand U11105 (N_11105,N_9808,N_9972);
and U11106 (N_11106,N_10344,N_9961);
xor U11107 (N_11107,N_9806,N_9777);
nand U11108 (N_11108,N_10384,N_9980);
or U11109 (N_11109,N_10077,N_9882);
nor U11110 (N_11110,N_10139,N_10328);
and U11111 (N_11111,N_9988,N_10362);
nor U11112 (N_11112,N_10034,N_9841);
and U11113 (N_11113,N_9994,N_9867);
nand U11114 (N_11114,N_9982,N_9764);
or U11115 (N_11115,N_10169,N_9921);
or U11116 (N_11116,N_10076,N_9945);
xnor U11117 (N_11117,N_10281,N_10000);
nor U11118 (N_11118,N_10049,N_9893);
nand U11119 (N_11119,N_9920,N_10120);
xor U11120 (N_11120,N_10167,N_10176);
and U11121 (N_11121,N_9957,N_10223);
and U11122 (N_11122,N_10437,N_9816);
and U11123 (N_11123,N_9836,N_10174);
or U11124 (N_11124,N_10128,N_10351);
or U11125 (N_11125,N_9983,N_9845);
nor U11126 (N_11126,N_9974,N_10481);
nor U11127 (N_11127,N_10476,N_9852);
or U11128 (N_11128,N_10432,N_9825);
or U11129 (N_11129,N_10350,N_10147);
nor U11130 (N_11130,N_10031,N_9901);
nand U11131 (N_11131,N_10247,N_10366);
and U11132 (N_11132,N_10118,N_9814);
nor U11133 (N_11133,N_10216,N_10393);
nor U11134 (N_11134,N_10072,N_10092);
and U11135 (N_11135,N_9820,N_9972);
or U11136 (N_11136,N_9879,N_9925);
and U11137 (N_11137,N_10421,N_10355);
nor U11138 (N_11138,N_9976,N_9822);
nand U11139 (N_11139,N_9982,N_9875);
nor U11140 (N_11140,N_10497,N_9939);
and U11141 (N_11141,N_10113,N_10222);
nand U11142 (N_11142,N_9827,N_10182);
nand U11143 (N_11143,N_10012,N_10134);
nor U11144 (N_11144,N_10072,N_10356);
nor U11145 (N_11145,N_10400,N_10348);
nor U11146 (N_11146,N_9984,N_9919);
nand U11147 (N_11147,N_10475,N_9888);
nor U11148 (N_11148,N_9859,N_10223);
nor U11149 (N_11149,N_10455,N_10005);
nand U11150 (N_11150,N_9900,N_9989);
or U11151 (N_11151,N_10011,N_9802);
or U11152 (N_11152,N_10429,N_9827);
nor U11153 (N_11153,N_9889,N_10153);
or U11154 (N_11154,N_10414,N_10218);
and U11155 (N_11155,N_10301,N_9906);
xor U11156 (N_11156,N_9895,N_10067);
or U11157 (N_11157,N_10392,N_10204);
nand U11158 (N_11158,N_10425,N_10175);
nor U11159 (N_11159,N_9979,N_10480);
nor U11160 (N_11160,N_10486,N_10019);
nand U11161 (N_11161,N_10382,N_10163);
nor U11162 (N_11162,N_10418,N_10357);
xnor U11163 (N_11163,N_10006,N_9853);
nor U11164 (N_11164,N_10446,N_10401);
xnor U11165 (N_11165,N_10429,N_10148);
nor U11166 (N_11166,N_10396,N_10409);
and U11167 (N_11167,N_10087,N_9867);
nand U11168 (N_11168,N_10365,N_9866);
nor U11169 (N_11169,N_10123,N_10281);
xnor U11170 (N_11170,N_9833,N_10484);
nand U11171 (N_11171,N_9861,N_10107);
nand U11172 (N_11172,N_10254,N_9926);
and U11173 (N_11173,N_10459,N_9778);
and U11174 (N_11174,N_10090,N_10198);
or U11175 (N_11175,N_10080,N_10333);
nor U11176 (N_11176,N_10042,N_10345);
nor U11177 (N_11177,N_9837,N_10482);
nor U11178 (N_11178,N_9767,N_10301);
and U11179 (N_11179,N_10282,N_10349);
xor U11180 (N_11180,N_10238,N_10066);
nor U11181 (N_11181,N_10272,N_10142);
and U11182 (N_11182,N_10457,N_10459);
or U11183 (N_11183,N_9803,N_10338);
and U11184 (N_11184,N_10488,N_10486);
xor U11185 (N_11185,N_9767,N_9954);
and U11186 (N_11186,N_9824,N_9902);
and U11187 (N_11187,N_10337,N_10101);
nand U11188 (N_11188,N_10320,N_10253);
and U11189 (N_11189,N_10481,N_10031);
xor U11190 (N_11190,N_10344,N_10148);
nor U11191 (N_11191,N_9874,N_9867);
or U11192 (N_11192,N_10363,N_9936);
or U11193 (N_11193,N_10115,N_9880);
nand U11194 (N_11194,N_10321,N_10447);
and U11195 (N_11195,N_10328,N_10295);
nand U11196 (N_11196,N_10088,N_10412);
or U11197 (N_11197,N_10418,N_9945);
nand U11198 (N_11198,N_10057,N_10446);
and U11199 (N_11199,N_10317,N_10200);
nor U11200 (N_11200,N_9853,N_10020);
nand U11201 (N_11201,N_10304,N_10061);
nand U11202 (N_11202,N_9828,N_9867);
and U11203 (N_11203,N_9764,N_10129);
nor U11204 (N_11204,N_10257,N_10329);
nor U11205 (N_11205,N_10445,N_10350);
or U11206 (N_11206,N_10241,N_10352);
and U11207 (N_11207,N_10161,N_10042);
nand U11208 (N_11208,N_9830,N_10031);
nand U11209 (N_11209,N_9924,N_9774);
or U11210 (N_11210,N_10076,N_10005);
nor U11211 (N_11211,N_9938,N_10475);
or U11212 (N_11212,N_9839,N_10095);
nand U11213 (N_11213,N_10297,N_10279);
and U11214 (N_11214,N_10082,N_10261);
nand U11215 (N_11215,N_10063,N_9850);
nand U11216 (N_11216,N_10422,N_9849);
or U11217 (N_11217,N_9811,N_10062);
and U11218 (N_11218,N_10027,N_10367);
or U11219 (N_11219,N_10499,N_10072);
or U11220 (N_11220,N_9990,N_9819);
nor U11221 (N_11221,N_9866,N_10036);
nor U11222 (N_11222,N_10446,N_9928);
or U11223 (N_11223,N_10464,N_10495);
or U11224 (N_11224,N_10165,N_10392);
nor U11225 (N_11225,N_9809,N_10371);
nor U11226 (N_11226,N_10043,N_10384);
and U11227 (N_11227,N_10337,N_10312);
or U11228 (N_11228,N_9865,N_10029);
nor U11229 (N_11229,N_10346,N_10147);
nand U11230 (N_11230,N_10177,N_9777);
and U11231 (N_11231,N_10294,N_10280);
and U11232 (N_11232,N_10267,N_9970);
and U11233 (N_11233,N_10214,N_9771);
nand U11234 (N_11234,N_9911,N_10385);
or U11235 (N_11235,N_10207,N_10386);
nor U11236 (N_11236,N_9772,N_10231);
nand U11237 (N_11237,N_9836,N_10231);
xnor U11238 (N_11238,N_9895,N_10392);
or U11239 (N_11239,N_10227,N_9778);
nand U11240 (N_11240,N_10361,N_10368);
or U11241 (N_11241,N_9852,N_10490);
or U11242 (N_11242,N_9808,N_10318);
and U11243 (N_11243,N_10422,N_10244);
nand U11244 (N_11244,N_10297,N_10243);
or U11245 (N_11245,N_10394,N_10374);
xor U11246 (N_11246,N_10399,N_10362);
and U11247 (N_11247,N_9903,N_9910);
and U11248 (N_11248,N_10251,N_10324);
and U11249 (N_11249,N_9763,N_9880);
and U11250 (N_11250,N_10643,N_10532);
and U11251 (N_11251,N_10540,N_10870);
or U11252 (N_11252,N_11089,N_11099);
nor U11253 (N_11253,N_11234,N_10700);
nand U11254 (N_11254,N_11070,N_10738);
or U11255 (N_11255,N_10929,N_11035);
nor U11256 (N_11256,N_10732,N_10910);
nor U11257 (N_11257,N_11025,N_11131);
nor U11258 (N_11258,N_11181,N_10786);
nand U11259 (N_11259,N_11076,N_10845);
nor U11260 (N_11260,N_10855,N_10974);
nand U11261 (N_11261,N_10940,N_10504);
nand U11262 (N_11262,N_10515,N_11156);
or U11263 (N_11263,N_11227,N_11188);
nor U11264 (N_11264,N_11196,N_11249);
and U11265 (N_11265,N_10511,N_10521);
nand U11266 (N_11266,N_10911,N_10885);
and U11267 (N_11267,N_11244,N_10905);
xnor U11268 (N_11268,N_11215,N_10780);
nand U11269 (N_11269,N_11246,N_10634);
nor U11270 (N_11270,N_10606,N_10967);
nor U11271 (N_11271,N_10691,N_11218);
nand U11272 (N_11272,N_11153,N_11157);
and U11273 (N_11273,N_10567,N_11186);
or U11274 (N_11274,N_10985,N_10657);
nand U11275 (N_11275,N_10604,N_10919);
xor U11276 (N_11276,N_11136,N_10562);
nand U11277 (N_11277,N_10564,N_10512);
or U11278 (N_11278,N_10640,N_11170);
and U11279 (N_11279,N_11116,N_11229);
nand U11280 (N_11280,N_11243,N_11010);
or U11281 (N_11281,N_10728,N_11117);
nor U11282 (N_11282,N_10825,N_10617);
nand U11283 (N_11283,N_10956,N_11111);
nand U11284 (N_11284,N_10693,N_10707);
or U11285 (N_11285,N_10698,N_11128);
or U11286 (N_11286,N_10601,N_10734);
or U11287 (N_11287,N_10976,N_10687);
nor U11288 (N_11288,N_11033,N_11164);
or U11289 (N_11289,N_11032,N_11064);
or U11290 (N_11290,N_10986,N_11062);
and U11291 (N_11291,N_10755,N_10810);
and U11292 (N_11292,N_10864,N_10569);
nand U11293 (N_11293,N_10716,N_10970);
nor U11294 (N_11294,N_10850,N_11160);
nor U11295 (N_11295,N_10580,N_11014);
nor U11296 (N_11296,N_10658,N_11109);
nand U11297 (N_11297,N_10662,N_10995);
and U11298 (N_11298,N_10774,N_10748);
and U11299 (N_11299,N_11187,N_10607);
nor U11300 (N_11300,N_10610,N_10706);
or U11301 (N_11301,N_10808,N_10575);
or U11302 (N_11302,N_11171,N_10740);
xor U11303 (N_11303,N_10804,N_10922);
or U11304 (N_11304,N_10868,N_10697);
nor U11305 (N_11305,N_10730,N_10923);
and U11306 (N_11306,N_10649,N_10867);
nor U11307 (N_11307,N_10705,N_10824);
and U11308 (N_11308,N_10600,N_10928);
nand U11309 (N_11309,N_10899,N_11114);
and U11310 (N_11310,N_10623,N_10949);
nor U11311 (N_11311,N_10816,N_10796);
nor U11312 (N_11312,N_10684,N_10865);
or U11313 (N_11313,N_11067,N_10669);
nand U11314 (N_11314,N_10921,N_11237);
nor U11315 (N_11315,N_10914,N_11007);
nand U11316 (N_11316,N_11021,N_11066);
nor U11317 (N_11317,N_10689,N_10988);
nand U11318 (N_11318,N_10819,N_10888);
xnor U11319 (N_11319,N_11130,N_10987);
nand U11320 (N_11320,N_11209,N_10508);
or U11321 (N_11321,N_10813,N_10803);
nand U11322 (N_11322,N_11073,N_10686);
nor U11323 (N_11323,N_10663,N_10869);
and U11324 (N_11324,N_10677,N_11219);
nand U11325 (N_11325,N_10841,N_11204);
nor U11326 (N_11326,N_10572,N_11221);
nand U11327 (N_11327,N_11036,N_11100);
xor U11328 (N_11328,N_11094,N_10602);
xor U11329 (N_11329,N_10638,N_10652);
xnor U11330 (N_11330,N_11077,N_11048);
or U11331 (N_11331,N_10696,N_10584);
nand U11332 (N_11332,N_11024,N_10828);
or U11333 (N_11333,N_10635,N_11200);
or U11334 (N_11334,N_11096,N_10761);
and U11335 (N_11335,N_10509,N_11151);
or U11336 (N_11336,N_10616,N_11217);
or U11337 (N_11337,N_10563,N_10539);
nor U11338 (N_11338,N_10901,N_11009);
and U11339 (N_11339,N_11084,N_10797);
xnor U11340 (N_11340,N_10897,N_11046);
nor U11341 (N_11341,N_10546,N_10861);
nand U11342 (N_11342,N_11242,N_10637);
and U11343 (N_11343,N_11051,N_10958);
nor U11344 (N_11344,N_10534,N_11052);
nand U11345 (N_11345,N_11197,N_10903);
nor U11346 (N_11346,N_10993,N_10944);
xor U11347 (N_11347,N_11163,N_10720);
and U11348 (N_11348,N_11239,N_10785);
nand U11349 (N_11349,N_11068,N_11125);
nand U11350 (N_11350,N_10592,N_10822);
nor U11351 (N_11351,N_10846,N_11095);
nor U11352 (N_11352,N_10514,N_10975);
nand U11353 (N_11353,N_11055,N_10847);
nor U11354 (N_11354,N_10613,N_10984);
and U11355 (N_11355,N_11030,N_10737);
or U11356 (N_11356,N_10891,N_11090);
or U11357 (N_11357,N_10962,N_11016);
nor U11358 (N_11358,N_10630,N_11003);
or U11359 (N_11359,N_11149,N_11248);
and U11360 (N_11360,N_10555,N_11056);
nor U11361 (N_11361,N_10605,N_10904);
or U11362 (N_11362,N_10530,N_10680);
nor U11363 (N_11363,N_10772,N_10595);
or U11364 (N_11364,N_10969,N_10844);
xor U11365 (N_11365,N_10908,N_10971);
nand U11366 (N_11366,N_10588,N_10980);
nand U11367 (N_11367,N_10682,N_10832);
xnor U11368 (N_11368,N_10551,N_11231);
and U11369 (N_11369,N_10858,N_10729);
nor U11370 (N_11370,N_10754,N_11023);
or U11371 (N_11371,N_10934,N_10943);
nand U11372 (N_11372,N_10760,N_10671);
and U11373 (N_11373,N_10945,N_10957);
nand U11374 (N_11374,N_10895,N_10890);
xnor U11375 (N_11375,N_10789,N_10766);
and U11376 (N_11376,N_10577,N_10982);
nand U11377 (N_11377,N_11106,N_11103);
nand U11378 (N_11378,N_11223,N_10947);
nor U11379 (N_11379,N_10880,N_11150);
nor U11380 (N_11380,N_10665,N_10821);
xor U11381 (N_11381,N_10747,N_10547);
nand U11382 (N_11382,N_10714,N_11207);
nor U11383 (N_11383,N_10673,N_11083);
nand U11384 (N_11384,N_10552,N_10852);
or U11385 (N_11385,N_10875,N_10827);
nor U11386 (N_11386,N_10717,N_11137);
and U11387 (N_11387,N_10763,N_10834);
nand U11388 (N_11388,N_10953,N_10955);
xor U11389 (N_11389,N_10675,N_11148);
nor U11390 (N_11390,N_11178,N_10571);
or U11391 (N_11391,N_10526,N_10653);
or U11392 (N_11392,N_10543,N_10719);
nor U11393 (N_11393,N_10873,N_10725);
or U11394 (N_11394,N_10833,N_10863);
nand U11395 (N_11395,N_10773,N_10710);
and U11396 (N_11396,N_11122,N_11166);
nor U11397 (N_11397,N_10859,N_10536);
nand U11398 (N_11398,N_11082,N_10907);
nor U11399 (N_11399,N_10690,N_11026);
or U11400 (N_11400,N_10744,N_10603);
nor U11401 (N_11401,N_11069,N_10860);
and U11402 (N_11402,N_11185,N_10633);
xnor U11403 (N_11403,N_11044,N_11102);
or U11404 (N_11404,N_10527,N_11133);
or U11405 (N_11405,N_10933,N_10624);
and U11406 (N_11406,N_11074,N_10507);
or U11407 (N_11407,N_10681,N_10502);
xor U11408 (N_11408,N_11142,N_11140);
or U11409 (N_11409,N_11230,N_10735);
or U11410 (N_11410,N_10593,N_11220);
and U11411 (N_11411,N_11013,N_10642);
and U11412 (N_11412,N_10742,N_10902);
nand U11413 (N_11413,N_10784,N_11245);
and U11414 (N_11414,N_10884,N_11011);
nor U11415 (N_11415,N_10722,N_10599);
and U11416 (N_11416,N_10764,N_10959);
nor U11417 (N_11417,N_10900,N_10983);
or U11418 (N_11418,N_11205,N_10779);
nor U11419 (N_11419,N_10924,N_11034);
nand U11420 (N_11420,N_11183,N_11155);
xnor U11421 (N_11421,N_10886,N_11132);
and U11422 (N_11422,N_10629,N_11097);
xor U11423 (N_11423,N_11216,N_10777);
or U11424 (N_11424,N_10752,N_10583);
xnor U11425 (N_11425,N_10879,N_11028);
xnor U11426 (N_11426,N_10505,N_10589);
nand U11427 (N_11427,N_10582,N_10915);
and U11428 (N_11428,N_10538,N_10506);
or U11429 (N_11429,N_11079,N_11123);
xor U11430 (N_11430,N_10767,N_10800);
nor U11431 (N_11431,N_10759,N_10793);
nand U11432 (N_11432,N_10501,N_10932);
or U11433 (N_11433,N_10654,N_10553);
and U11434 (N_11434,N_10749,N_11158);
xor U11435 (N_11435,N_10938,N_10570);
or U11436 (N_11436,N_11210,N_11192);
and U11437 (N_11437,N_10802,N_10645);
nand U11438 (N_11438,N_11127,N_10598);
nand U11439 (N_11439,N_11061,N_10826);
or U11440 (N_11440,N_10990,N_10812);
nand U11441 (N_11441,N_10718,N_10936);
xor U11442 (N_11442,N_11000,N_11112);
or U11443 (N_11443,N_10715,N_11017);
nand U11444 (N_11444,N_10762,N_10733);
nand U11445 (N_11445,N_11161,N_10997);
and U11446 (N_11446,N_10618,N_10529);
and U11447 (N_11447,N_10712,N_10776);
nand U11448 (N_11448,N_10765,N_10631);
or U11449 (N_11449,N_10731,N_11105);
and U11450 (N_11450,N_10787,N_11180);
nand U11451 (N_11451,N_10843,N_10920);
and U11452 (N_11452,N_10661,N_10842);
nor U11453 (N_11453,N_11147,N_10650);
and U11454 (N_11454,N_10952,N_10704);
and U11455 (N_11455,N_11047,N_10794);
and U11456 (N_11456,N_10926,N_10678);
nand U11457 (N_11457,N_11247,N_11004);
nand U11458 (N_11458,N_11154,N_10753);
xor U11459 (N_11459,N_10966,N_10882);
or U11460 (N_11460,N_10524,N_10801);
nor U11461 (N_11461,N_11169,N_11029);
nand U11462 (N_11462,N_11177,N_10622);
or U11463 (N_11463,N_10636,N_10670);
or U11464 (N_11464,N_10612,N_10964);
nand U11465 (N_11465,N_10892,N_10913);
or U11466 (N_11466,N_10877,N_10961);
or U11467 (N_11467,N_10711,N_10778);
and U11468 (N_11468,N_10835,N_10586);
xnor U11469 (N_11469,N_10830,N_10836);
nor U11470 (N_11470,N_10646,N_10587);
or U11471 (N_11471,N_10792,N_10896);
or U11472 (N_11472,N_10806,N_10666);
or U11473 (N_11473,N_10664,N_10609);
or U11474 (N_11474,N_10676,N_11015);
nor U11475 (N_11475,N_10790,N_10639);
nor U11476 (N_11476,N_10541,N_10769);
nand U11477 (N_11477,N_11087,N_10566);
nand U11478 (N_11478,N_11198,N_10724);
nand U11479 (N_11479,N_10655,N_10608);
nand U11480 (N_11480,N_10965,N_10770);
or U11481 (N_11481,N_11050,N_10831);
nor U11482 (N_11482,N_11054,N_10840);
nor U11483 (N_11483,N_10672,N_10517);
xnor U11484 (N_11484,N_10817,N_10513);
nand U11485 (N_11485,N_10556,N_10708);
nand U11486 (N_11486,N_11081,N_10935);
nand U11487 (N_11487,N_10849,N_10626);
nand U11488 (N_11488,N_10627,N_10739);
nor U11489 (N_11489,N_10620,N_11093);
and U11490 (N_11490,N_10736,N_11174);
and U11491 (N_11491,N_10992,N_11080);
nor U11492 (N_11492,N_11020,N_11037);
nor U11493 (N_11493,N_10838,N_10781);
and U11494 (N_11494,N_10948,N_10519);
nand U11495 (N_11495,N_11228,N_11049);
or U11496 (N_11496,N_10917,N_10573);
nand U11497 (N_11497,N_11232,N_11195);
or U11498 (N_11498,N_10916,N_10893);
and U11499 (N_11499,N_11031,N_11129);
or U11500 (N_11500,N_10931,N_11213);
or U11501 (N_11501,N_11175,N_10795);
or U11502 (N_11502,N_10815,N_11135);
and U11503 (N_11503,N_10918,N_10578);
or U11504 (N_11504,N_10741,N_10644);
xnor U11505 (N_11505,N_10548,N_11152);
nand U11506 (N_11506,N_10510,N_11235);
or U11507 (N_11507,N_10520,N_10667);
nor U11508 (N_11508,N_10743,N_11065);
nor U11509 (N_11509,N_10909,N_10701);
nor U11510 (N_11510,N_10783,N_10963);
nor U11511 (N_11511,N_10937,N_10648);
or U11512 (N_11512,N_10898,N_10619);
and U11513 (N_11513,N_10788,N_11222);
nor U11514 (N_11514,N_11072,N_10590);
and U11515 (N_11515,N_10925,N_10615);
or U11516 (N_11516,N_10503,N_10876);
or U11517 (N_11517,N_11118,N_10565);
nor U11518 (N_11518,N_11040,N_10839);
and U11519 (N_11519,N_10621,N_10574);
and U11520 (N_11520,N_11039,N_10894);
or U11521 (N_11521,N_11233,N_11058);
nand U11522 (N_11522,N_11238,N_10721);
and U11523 (N_11523,N_11193,N_10713);
and U11524 (N_11524,N_11168,N_10791);
and U11525 (N_11525,N_11063,N_10668);
xnor U11526 (N_11526,N_10625,N_10887);
and U11527 (N_11527,N_10756,N_10641);
and U11528 (N_11528,N_10853,N_11098);
or U11529 (N_11529,N_11086,N_10856);
xor U11530 (N_11530,N_10878,N_10751);
and U11531 (N_11531,N_10874,N_11194);
or U11532 (N_11532,N_11124,N_11173);
and U11533 (N_11533,N_10807,N_11212);
and U11534 (N_11534,N_10818,N_10837);
nor U11535 (N_11535,N_10647,N_10883);
nor U11536 (N_11536,N_11027,N_11240);
or U11537 (N_11537,N_11165,N_10805);
or U11538 (N_11538,N_10703,N_11208);
nand U11539 (N_11539,N_11108,N_11008);
nand U11540 (N_11540,N_11092,N_10862);
or U11541 (N_11541,N_10542,N_10823);
nand U11542 (N_11542,N_11120,N_10768);
or U11543 (N_11543,N_10614,N_10848);
xor U11544 (N_11544,N_11191,N_11038);
or U11545 (N_11545,N_11146,N_10568);
nor U11546 (N_11546,N_10659,N_10695);
or U11547 (N_11547,N_11119,N_10930);
or U11548 (N_11548,N_10912,N_10656);
and U11549 (N_11549,N_10518,N_11236);
nand U11550 (N_11550,N_10745,N_10857);
nand U11551 (N_11551,N_10560,N_11043);
nor U11552 (N_11552,N_11126,N_10996);
xnor U11553 (N_11553,N_10972,N_10699);
nor U11554 (N_11554,N_10998,N_11085);
and U11555 (N_11555,N_10533,N_10798);
and U11556 (N_11556,N_11226,N_10523);
or U11557 (N_11557,N_10799,N_10692);
and U11558 (N_11558,N_10525,N_11179);
and U11559 (N_11559,N_11045,N_10939);
nor U11560 (N_11560,N_10554,N_10977);
and U11561 (N_11561,N_11176,N_10866);
and U11562 (N_11562,N_11113,N_10950);
or U11563 (N_11563,N_11022,N_10889);
nor U11564 (N_11564,N_11203,N_11189);
nor U11565 (N_11565,N_11060,N_10871);
and U11566 (N_11566,N_11121,N_11101);
and U11567 (N_11567,N_11075,N_10727);
nor U11568 (N_11568,N_10991,N_11145);
or U11569 (N_11569,N_10775,N_10544);
nor U11570 (N_11570,N_10522,N_10746);
or U11571 (N_11571,N_10726,N_10628);
or U11572 (N_11572,N_10979,N_10927);
or U11573 (N_11573,N_10750,N_10968);
or U11574 (N_11574,N_11159,N_10674);
or U11575 (N_11575,N_10597,N_10660);
and U11576 (N_11576,N_10771,N_10829);
nand U11577 (N_11577,N_10528,N_10973);
nand U11578 (N_11578,N_10951,N_11139);
nor U11579 (N_11579,N_10954,N_11006);
nand U11580 (N_11580,N_11019,N_10981);
nor U11581 (N_11581,N_11059,N_10685);
nor U11582 (N_11582,N_11184,N_11162);
and U11583 (N_11583,N_10537,N_10723);
or U11584 (N_11584,N_11241,N_11202);
xor U11585 (N_11585,N_10851,N_10585);
or U11586 (N_11586,N_10820,N_11182);
nand U11587 (N_11587,N_10709,N_10558);
nand U11588 (N_11588,N_11042,N_10757);
and U11589 (N_11589,N_11224,N_10579);
xor U11590 (N_11590,N_10683,N_10561);
nor U11591 (N_11591,N_11018,N_11214);
and U11592 (N_11592,N_10688,N_11071);
nand U11593 (N_11593,N_11115,N_10651);
nand U11594 (N_11594,N_10557,N_10611);
or U11595 (N_11595,N_10545,N_11091);
or U11596 (N_11596,N_11002,N_10549);
nor U11597 (N_11597,N_11206,N_10906);
nand U11598 (N_11598,N_10999,N_10854);
or U11599 (N_11599,N_10942,N_10500);
nand U11600 (N_11600,N_10594,N_10941);
nor U11601 (N_11601,N_10782,N_10591);
xnor U11602 (N_11602,N_11078,N_10758);
and U11603 (N_11603,N_11088,N_11005);
nor U11604 (N_11604,N_10872,N_10581);
or U11605 (N_11605,N_10531,N_11138);
nor U11606 (N_11606,N_11001,N_10811);
and U11607 (N_11607,N_10989,N_11199);
nand U11608 (N_11608,N_10550,N_11012);
nor U11609 (N_11609,N_11141,N_10702);
or U11610 (N_11610,N_10946,N_10535);
or U11611 (N_11611,N_11201,N_10559);
and U11612 (N_11612,N_10881,N_10516);
and U11613 (N_11613,N_11104,N_10994);
or U11614 (N_11614,N_10596,N_11107);
and U11615 (N_11615,N_10694,N_11167);
and U11616 (N_11616,N_11134,N_11041);
and U11617 (N_11617,N_11110,N_11190);
nand U11618 (N_11618,N_11172,N_10632);
nand U11619 (N_11619,N_10978,N_10809);
nand U11620 (N_11620,N_10576,N_11225);
or U11621 (N_11621,N_11057,N_11211);
nand U11622 (N_11622,N_11143,N_10960);
nor U11623 (N_11623,N_10814,N_11144);
nor U11624 (N_11624,N_10679,N_11053);
or U11625 (N_11625,N_10769,N_11078);
nor U11626 (N_11626,N_10932,N_10726);
xor U11627 (N_11627,N_10991,N_11194);
or U11628 (N_11628,N_10947,N_10934);
or U11629 (N_11629,N_10740,N_10672);
and U11630 (N_11630,N_10890,N_10840);
nand U11631 (N_11631,N_11082,N_11200);
nor U11632 (N_11632,N_10978,N_10972);
and U11633 (N_11633,N_10989,N_10611);
or U11634 (N_11634,N_11121,N_10974);
nor U11635 (N_11635,N_10923,N_10928);
nand U11636 (N_11636,N_11214,N_10676);
or U11637 (N_11637,N_11029,N_10839);
and U11638 (N_11638,N_11014,N_10645);
and U11639 (N_11639,N_10996,N_10956);
and U11640 (N_11640,N_10668,N_10844);
or U11641 (N_11641,N_10703,N_11242);
nor U11642 (N_11642,N_10505,N_10991);
and U11643 (N_11643,N_11029,N_10573);
nor U11644 (N_11644,N_11107,N_10888);
nor U11645 (N_11645,N_10740,N_10787);
nand U11646 (N_11646,N_11058,N_10753);
nor U11647 (N_11647,N_10574,N_11193);
and U11648 (N_11648,N_10503,N_10867);
nor U11649 (N_11649,N_11231,N_11191);
xnor U11650 (N_11650,N_10706,N_10998);
xnor U11651 (N_11651,N_10893,N_11245);
xnor U11652 (N_11652,N_10684,N_10886);
and U11653 (N_11653,N_11033,N_10854);
nand U11654 (N_11654,N_10723,N_10771);
nor U11655 (N_11655,N_10934,N_11032);
nor U11656 (N_11656,N_10598,N_10651);
nor U11657 (N_11657,N_11217,N_10809);
and U11658 (N_11658,N_11206,N_11184);
nand U11659 (N_11659,N_10813,N_10570);
xor U11660 (N_11660,N_10697,N_10536);
nor U11661 (N_11661,N_10847,N_10564);
and U11662 (N_11662,N_10963,N_10764);
nor U11663 (N_11663,N_10559,N_11082);
and U11664 (N_11664,N_11053,N_11056);
or U11665 (N_11665,N_11033,N_10766);
or U11666 (N_11666,N_11108,N_10739);
nor U11667 (N_11667,N_11195,N_10664);
nand U11668 (N_11668,N_10979,N_10758);
nor U11669 (N_11669,N_10620,N_10656);
and U11670 (N_11670,N_10545,N_10731);
nand U11671 (N_11671,N_11057,N_11187);
nor U11672 (N_11672,N_10983,N_10500);
or U11673 (N_11673,N_10876,N_10661);
nand U11674 (N_11674,N_10545,N_11093);
or U11675 (N_11675,N_10642,N_10501);
xnor U11676 (N_11676,N_10545,N_10569);
nand U11677 (N_11677,N_10647,N_10746);
and U11678 (N_11678,N_11133,N_10746);
and U11679 (N_11679,N_10681,N_10891);
nor U11680 (N_11680,N_10901,N_10899);
and U11681 (N_11681,N_10723,N_10604);
and U11682 (N_11682,N_10607,N_10813);
nand U11683 (N_11683,N_10894,N_11209);
xor U11684 (N_11684,N_11113,N_10756);
and U11685 (N_11685,N_10792,N_11071);
nand U11686 (N_11686,N_10871,N_11120);
or U11687 (N_11687,N_10843,N_10680);
and U11688 (N_11688,N_11231,N_11049);
or U11689 (N_11689,N_11233,N_11067);
nor U11690 (N_11690,N_10813,N_11112);
or U11691 (N_11691,N_10525,N_10807);
nand U11692 (N_11692,N_10774,N_10899);
and U11693 (N_11693,N_11066,N_11158);
and U11694 (N_11694,N_10984,N_10605);
or U11695 (N_11695,N_10949,N_10806);
nand U11696 (N_11696,N_10711,N_11201);
or U11697 (N_11697,N_11248,N_10740);
nor U11698 (N_11698,N_11085,N_11006);
nand U11699 (N_11699,N_10701,N_10621);
nor U11700 (N_11700,N_11072,N_10723);
nor U11701 (N_11701,N_10921,N_10603);
or U11702 (N_11702,N_11040,N_10545);
xnor U11703 (N_11703,N_10637,N_11105);
nor U11704 (N_11704,N_11072,N_10927);
nand U11705 (N_11705,N_11022,N_11145);
and U11706 (N_11706,N_11206,N_11081);
nand U11707 (N_11707,N_10700,N_10703);
and U11708 (N_11708,N_10924,N_10774);
xnor U11709 (N_11709,N_11188,N_10627);
and U11710 (N_11710,N_11145,N_11218);
and U11711 (N_11711,N_10924,N_10803);
and U11712 (N_11712,N_11019,N_10827);
or U11713 (N_11713,N_10604,N_11205);
nor U11714 (N_11714,N_11039,N_11005);
or U11715 (N_11715,N_10747,N_11038);
or U11716 (N_11716,N_10839,N_10622);
xor U11717 (N_11717,N_10877,N_11240);
xnor U11718 (N_11718,N_10718,N_10578);
or U11719 (N_11719,N_10976,N_10575);
and U11720 (N_11720,N_11210,N_11115);
nand U11721 (N_11721,N_10671,N_10900);
and U11722 (N_11722,N_10694,N_10770);
nor U11723 (N_11723,N_10521,N_11204);
or U11724 (N_11724,N_10576,N_10751);
nor U11725 (N_11725,N_10890,N_10607);
xnor U11726 (N_11726,N_11053,N_10622);
nand U11727 (N_11727,N_10661,N_10708);
nor U11728 (N_11728,N_11066,N_11150);
nor U11729 (N_11729,N_11073,N_10544);
nor U11730 (N_11730,N_11060,N_10906);
nor U11731 (N_11731,N_11092,N_11115);
nand U11732 (N_11732,N_10778,N_10617);
or U11733 (N_11733,N_10935,N_10781);
nor U11734 (N_11734,N_11047,N_10972);
and U11735 (N_11735,N_11044,N_10920);
nand U11736 (N_11736,N_10656,N_10992);
nor U11737 (N_11737,N_10622,N_11105);
xor U11738 (N_11738,N_11175,N_10702);
nand U11739 (N_11739,N_10797,N_10957);
and U11740 (N_11740,N_10894,N_10608);
and U11741 (N_11741,N_11191,N_10590);
and U11742 (N_11742,N_11097,N_11238);
nand U11743 (N_11743,N_11213,N_11088);
nor U11744 (N_11744,N_11073,N_10873);
nor U11745 (N_11745,N_10952,N_10882);
nand U11746 (N_11746,N_10899,N_10699);
or U11747 (N_11747,N_10936,N_10820);
or U11748 (N_11748,N_10908,N_10924);
and U11749 (N_11749,N_10562,N_10568);
nand U11750 (N_11750,N_10506,N_10987);
or U11751 (N_11751,N_11026,N_10865);
and U11752 (N_11752,N_10615,N_10536);
nor U11753 (N_11753,N_10708,N_11233);
and U11754 (N_11754,N_10771,N_11248);
and U11755 (N_11755,N_11095,N_10995);
and U11756 (N_11756,N_11042,N_11162);
or U11757 (N_11757,N_10884,N_11039);
nor U11758 (N_11758,N_10929,N_11120);
nor U11759 (N_11759,N_10601,N_10628);
nand U11760 (N_11760,N_11154,N_10749);
nor U11761 (N_11761,N_10539,N_10754);
and U11762 (N_11762,N_10881,N_10760);
xnor U11763 (N_11763,N_11080,N_11064);
or U11764 (N_11764,N_10954,N_10663);
nand U11765 (N_11765,N_10667,N_10622);
and U11766 (N_11766,N_11009,N_10528);
nor U11767 (N_11767,N_10526,N_10812);
or U11768 (N_11768,N_10526,N_11096);
and U11769 (N_11769,N_11063,N_10532);
xor U11770 (N_11770,N_11156,N_10590);
xor U11771 (N_11771,N_10958,N_11131);
xnor U11772 (N_11772,N_10525,N_10835);
and U11773 (N_11773,N_10928,N_10619);
or U11774 (N_11774,N_10761,N_10884);
and U11775 (N_11775,N_10651,N_10745);
nor U11776 (N_11776,N_10973,N_11169);
nand U11777 (N_11777,N_11117,N_10876);
and U11778 (N_11778,N_10604,N_10996);
or U11779 (N_11779,N_10652,N_10730);
nand U11780 (N_11780,N_10563,N_10763);
and U11781 (N_11781,N_11241,N_10942);
or U11782 (N_11782,N_10962,N_10585);
or U11783 (N_11783,N_10681,N_10509);
xor U11784 (N_11784,N_10566,N_11101);
xor U11785 (N_11785,N_10960,N_10879);
and U11786 (N_11786,N_11237,N_11097);
xor U11787 (N_11787,N_10977,N_11204);
xnor U11788 (N_11788,N_10542,N_11040);
nand U11789 (N_11789,N_11235,N_10825);
and U11790 (N_11790,N_11101,N_10975);
xnor U11791 (N_11791,N_10969,N_11176);
nor U11792 (N_11792,N_10846,N_10950);
nand U11793 (N_11793,N_11124,N_10517);
nor U11794 (N_11794,N_11207,N_10874);
xor U11795 (N_11795,N_10783,N_10554);
nor U11796 (N_11796,N_10931,N_10863);
nand U11797 (N_11797,N_11245,N_11044);
and U11798 (N_11798,N_10570,N_11001);
nor U11799 (N_11799,N_10794,N_10596);
and U11800 (N_11800,N_11074,N_10591);
nor U11801 (N_11801,N_10732,N_11118);
xor U11802 (N_11802,N_10913,N_11210);
nand U11803 (N_11803,N_10904,N_10533);
xnor U11804 (N_11804,N_11067,N_10814);
nand U11805 (N_11805,N_10815,N_10787);
nor U11806 (N_11806,N_10713,N_10666);
nand U11807 (N_11807,N_10987,N_10731);
nor U11808 (N_11808,N_10982,N_10502);
and U11809 (N_11809,N_11228,N_10898);
nor U11810 (N_11810,N_10782,N_11190);
nand U11811 (N_11811,N_10733,N_10941);
or U11812 (N_11812,N_11242,N_10934);
nor U11813 (N_11813,N_10828,N_10722);
nor U11814 (N_11814,N_11047,N_11129);
nor U11815 (N_11815,N_10899,N_10849);
xnor U11816 (N_11816,N_10716,N_10618);
nand U11817 (N_11817,N_10935,N_11210);
nand U11818 (N_11818,N_11068,N_10916);
nand U11819 (N_11819,N_11041,N_10981);
or U11820 (N_11820,N_10731,N_10945);
and U11821 (N_11821,N_11012,N_10793);
xnor U11822 (N_11822,N_10797,N_10816);
or U11823 (N_11823,N_11187,N_10908);
nor U11824 (N_11824,N_10848,N_10747);
or U11825 (N_11825,N_10651,N_11029);
or U11826 (N_11826,N_10681,N_10994);
nor U11827 (N_11827,N_10677,N_10888);
or U11828 (N_11828,N_10616,N_10647);
nor U11829 (N_11829,N_10903,N_10576);
nor U11830 (N_11830,N_11036,N_10806);
nor U11831 (N_11831,N_10979,N_11212);
or U11832 (N_11832,N_10820,N_10776);
nand U11833 (N_11833,N_10822,N_11222);
or U11834 (N_11834,N_10533,N_10829);
nor U11835 (N_11835,N_11036,N_11134);
nor U11836 (N_11836,N_11205,N_11024);
nand U11837 (N_11837,N_11081,N_11226);
xnor U11838 (N_11838,N_11249,N_10743);
nor U11839 (N_11839,N_10512,N_11089);
nor U11840 (N_11840,N_10822,N_10641);
nand U11841 (N_11841,N_11143,N_10892);
and U11842 (N_11842,N_10833,N_10669);
and U11843 (N_11843,N_10905,N_10910);
nand U11844 (N_11844,N_10911,N_11244);
nor U11845 (N_11845,N_10842,N_10803);
and U11846 (N_11846,N_10927,N_10649);
or U11847 (N_11847,N_11032,N_11106);
nand U11848 (N_11848,N_11221,N_10960);
or U11849 (N_11849,N_10994,N_11218);
and U11850 (N_11850,N_10766,N_10883);
or U11851 (N_11851,N_11100,N_10532);
nor U11852 (N_11852,N_11248,N_10891);
nor U11853 (N_11853,N_11040,N_11061);
or U11854 (N_11854,N_10643,N_11246);
or U11855 (N_11855,N_10558,N_10525);
and U11856 (N_11856,N_10621,N_10844);
nor U11857 (N_11857,N_10920,N_10881);
or U11858 (N_11858,N_11098,N_11076);
or U11859 (N_11859,N_10656,N_10651);
and U11860 (N_11860,N_10748,N_11031);
and U11861 (N_11861,N_10631,N_10596);
nor U11862 (N_11862,N_10828,N_10741);
xor U11863 (N_11863,N_10911,N_10775);
and U11864 (N_11864,N_11184,N_10976);
nand U11865 (N_11865,N_11194,N_11069);
nand U11866 (N_11866,N_10818,N_10915);
nor U11867 (N_11867,N_10587,N_11181);
nand U11868 (N_11868,N_10702,N_10617);
nor U11869 (N_11869,N_10855,N_11219);
and U11870 (N_11870,N_10714,N_10677);
and U11871 (N_11871,N_10826,N_10988);
nand U11872 (N_11872,N_10902,N_10743);
or U11873 (N_11873,N_11074,N_10504);
and U11874 (N_11874,N_11168,N_10891);
or U11875 (N_11875,N_10965,N_10537);
xor U11876 (N_11876,N_10501,N_11171);
xnor U11877 (N_11877,N_10817,N_11077);
and U11878 (N_11878,N_10823,N_10622);
and U11879 (N_11879,N_10654,N_11084);
nor U11880 (N_11880,N_10795,N_10891);
and U11881 (N_11881,N_10605,N_10604);
nand U11882 (N_11882,N_10987,N_11245);
or U11883 (N_11883,N_10682,N_10559);
xor U11884 (N_11884,N_10910,N_11010);
or U11885 (N_11885,N_10821,N_11086);
and U11886 (N_11886,N_11112,N_10981);
and U11887 (N_11887,N_11221,N_10697);
nor U11888 (N_11888,N_10655,N_10583);
xor U11889 (N_11889,N_11171,N_11080);
xnor U11890 (N_11890,N_10510,N_10587);
or U11891 (N_11891,N_10774,N_10895);
and U11892 (N_11892,N_11218,N_10801);
or U11893 (N_11893,N_10917,N_11087);
nor U11894 (N_11894,N_10992,N_11104);
xnor U11895 (N_11895,N_10511,N_10830);
nand U11896 (N_11896,N_10809,N_10588);
nor U11897 (N_11897,N_11077,N_10650);
nand U11898 (N_11898,N_10775,N_10681);
xnor U11899 (N_11899,N_10583,N_10613);
and U11900 (N_11900,N_10597,N_10670);
or U11901 (N_11901,N_10951,N_10799);
or U11902 (N_11902,N_10729,N_11020);
nand U11903 (N_11903,N_11230,N_10732);
nor U11904 (N_11904,N_11015,N_10778);
nand U11905 (N_11905,N_10508,N_10595);
nand U11906 (N_11906,N_10900,N_10752);
or U11907 (N_11907,N_10552,N_10844);
and U11908 (N_11908,N_10899,N_10874);
or U11909 (N_11909,N_11183,N_10637);
or U11910 (N_11910,N_10683,N_10779);
nand U11911 (N_11911,N_11235,N_11169);
nor U11912 (N_11912,N_10773,N_11029);
nand U11913 (N_11913,N_11118,N_11235);
xnor U11914 (N_11914,N_11215,N_10954);
and U11915 (N_11915,N_10950,N_10905);
nand U11916 (N_11916,N_10797,N_11045);
and U11917 (N_11917,N_11144,N_10807);
xor U11918 (N_11918,N_10839,N_10726);
and U11919 (N_11919,N_10952,N_10545);
nor U11920 (N_11920,N_10748,N_10589);
and U11921 (N_11921,N_10556,N_10859);
nand U11922 (N_11922,N_10565,N_10928);
or U11923 (N_11923,N_11140,N_10725);
xnor U11924 (N_11924,N_11193,N_11225);
xnor U11925 (N_11925,N_10500,N_10652);
nor U11926 (N_11926,N_11243,N_10813);
nand U11927 (N_11927,N_10982,N_10500);
nor U11928 (N_11928,N_11229,N_10798);
and U11929 (N_11929,N_11170,N_11200);
nor U11930 (N_11930,N_10746,N_10803);
xor U11931 (N_11931,N_10782,N_11067);
and U11932 (N_11932,N_10908,N_10946);
nor U11933 (N_11933,N_11243,N_11171);
xor U11934 (N_11934,N_11030,N_11215);
nand U11935 (N_11935,N_11008,N_10544);
nand U11936 (N_11936,N_10645,N_10928);
or U11937 (N_11937,N_10632,N_10710);
xnor U11938 (N_11938,N_10702,N_11091);
nor U11939 (N_11939,N_10805,N_11134);
nor U11940 (N_11940,N_10692,N_10607);
or U11941 (N_11941,N_10863,N_10895);
or U11942 (N_11942,N_10831,N_10633);
nor U11943 (N_11943,N_10574,N_11064);
or U11944 (N_11944,N_10913,N_10908);
nand U11945 (N_11945,N_11144,N_10879);
nor U11946 (N_11946,N_11235,N_11034);
xnor U11947 (N_11947,N_11051,N_10662);
nand U11948 (N_11948,N_10700,N_10647);
nand U11949 (N_11949,N_10825,N_10716);
or U11950 (N_11950,N_11078,N_11087);
and U11951 (N_11951,N_11204,N_10626);
and U11952 (N_11952,N_10880,N_10893);
or U11953 (N_11953,N_11113,N_11236);
nand U11954 (N_11954,N_11049,N_10662);
or U11955 (N_11955,N_10799,N_11099);
or U11956 (N_11956,N_10913,N_10958);
or U11957 (N_11957,N_10924,N_10750);
or U11958 (N_11958,N_10976,N_10835);
nor U11959 (N_11959,N_11071,N_10678);
and U11960 (N_11960,N_10663,N_10747);
and U11961 (N_11961,N_11185,N_11211);
nand U11962 (N_11962,N_10843,N_11219);
and U11963 (N_11963,N_11061,N_10856);
or U11964 (N_11964,N_11170,N_10889);
nor U11965 (N_11965,N_10776,N_10760);
nor U11966 (N_11966,N_10919,N_11228);
or U11967 (N_11967,N_10920,N_10769);
nor U11968 (N_11968,N_11247,N_10948);
xnor U11969 (N_11969,N_11128,N_10722);
nand U11970 (N_11970,N_11078,N_10961);
and U11971 (N_11971,N_11245,N_11123);
and U11972 (N_11972,N_10559,N_10732);
or U11973 (N_11973,N_10742,N_10830);
nor U11974 (N_11974,N_10776,N_10739);
and U11975 (N_11975,N_10568,N_11000);
or U11976 (N_11976,N_10527,N_10794);
and U11977 (N_11977,N_10682,N_10706);
and U11978 (N_11978,N_10844,N_10838);
nor U11979 (N_11979,N_11192,N_11110);
nor U11980 (N_11980,N_11142,N_11149);
and U11981 (N_11981,N_10773,N_11118);
xor U11982 (N_11982,N_10761,N_11187);
nand U11983 (N_11983,N_11068,N_11083);
and U11984 (N_11984,N_11203,N_10676);
nor U11985 (N_11985,N_10834,N_10958);
or U11986 (N_11986,N_10671,N_11121);
nand U11987 (N_11987,N_11249,N_11162);
or U11988 (N_11988,N_10950,N_10528);
and U11989 (N_11989,N_11105,N_10857);
and U11990 (N_11990,N_10872,N_11072);
and U11991 (N_11991,N_11194,N_10996);
or U11992 (N_11992,N_10968,N_10687);
nor U11993 (N_11993,N_10946,N_10547);
or U11994 (N_11994,N_10638,N_10928);
nand U11995 (N_11995,N_10943,N_11097);
nand U11996 (N_11996,N_10855,N_10610);
or U11997 (N_11997,N_10885,N_11016);
nor U11998 (N_11998,N_10684,N_10909);
nand U11999 (N_11999,N_11002,N_11064);
or U12000 (N_12000,N_11808,N_11685);
xor U12001 (N_12001,N_11622,N_11796);
and U12002 (N_12002,N_11312,N_11511);
nand U12003 (N_12003,N_11517,N_11754);
nor U12004 (N_12004,N_11818,N_11871);
and U12005 (N_12005,N_11355,N_11395);
nand U12006 (N_12006,N_11509,N_11743);
nor U12007 (N_12007,N_11321,N_11732);
and U12008 (N_12008,N_11368,N_11466);
or U12009 (N_12009,N_11772,N_11451);
or U12010 (N_12010,N_11566,N_11831);
nand U12011 (N_12011,N_11997,N_11946);
or U12012 (N_12012,N_11901,N_11450);
nand U12013 (N_12013,N_11474,N_11549);
xnor U12014 (N_12014,N_11801,N_11903);
or U12015 (N_12015,N_11610,N_11563);
nor U12016 (N_12016,N_11272,N_11933);
or U12017 (N_12017,N_11614,N_11583);
nand U12018 (N_12018,N_11372,N_11367);
nor U12019 (N_12019,N_11833,N_11787);
or U12020 (N_12020,N_11378,N_11364);
nand U12021 (N_12021,N_11883,N_11890);
or U12022 (N_12022,N_11740,N_11633);
nor U12023 (N_12023,N_11758,N_11483);
nand U12024 (N_12024,N_11371,N_11525);
xor U12025 (N_12025,N_11887,N_11617);
or U12026 (N_12026,N_11983,N_11965);
and U12027 (N_12027,N_11346,N_11334);
and U12028 (N_12028,N_11440,N_11287);
nor U12029 (N_12029,N_11489,N_11524);
or U12030 (N_12030,N_11710,N_11303);
nand U12031 (N_12031,N_11621,N_11435);
nor U12032 (N_12032,N_11516,N_11660);
xor U12033 (N_12033,N_11381,N_11688);
and U12034 (N_12034,N_11727,N_11313);
xnor U12035 (N_12035,N_11550,N_11891);
or U12036 (N_12036,N_11320,N_11932);
xor U12037 (N_12037,N_11845,N_11437);
nor U12038 (N_12038,N_11693,N_11264);
and U12039 (N_12039,N_11384,N_11588);
or U12040 (N_12040,N_11856,N_11971);
xor U12041 (N_12041,N_11537,N_11944);
nor U12042 (N_12042,N_11487,N_11842);
nor U12043 (N_12043,N_11734,N_11315);
nand U12044 (N_12044,N_11306,N_11806);
xnor U12045 (N_12045,N_11612,N_11514);
nor U12046 (N_12046,N_11676,N_11939);
and U12047 (N_12047,N_11812,N_11943);
or U12048 (N_12048,N_11824,N_11777);
or U12049 (N_12049,N_11492,N_11584);
and U12050 (N_12050,N_11900,N_11626);
and U12051 (N_12051,N_11804,N_11962);
xor U12052 (N_12052,N_11905,N_11724);
nor U12053 (N_12053,N_11572,N_11858);
or U12054 (N_12054,N_11714,N_11336);
nor U12055 (N_12055,N_11296,N_11337);
or U12056 (N_12056,N_11632,N_11722);
and U12057 (N_12057,N_11629,N_11847);
or U12058 (N_12058,N_11473,N_11460);
nor U12059 (N_12059,N_11565,N_11852);
nor U12060 (N_12060,N_11697,N_11426);
and U12061 (N_12061,N_11781,N_11791);
nand U12062 (N_12062,N_11659,N_11775);
nand U12063 (N_12063,N_11618,N_11674);
nand U12064 (N_12064,N_11434,N_11362);
or U12065 (N_12065,N_11874,N_11359);
xnor U12066 (N_12066,N_11653,N_11665);
or U12067 (N_12067,N_11253,N_11319);
nand U12068 (N_12068,N_11959,N_11706);
nor U12069 (N_12069,N_11508,N_11578);
nand U12070 (N_12070,N_11683,N_11580);
nor U12071 (N_12071,N_11638,N_11314);
nor U12072 (N_12072,N_11398,N_11561);
nor U12073 (N_12073,N_11627,N_11968);
nand U12074 (N_12074,N_11555,N_11488);
nand U12075 (N_12075,N_11540,N_11698);
nand U12076 (N_12076,N_11630,N_11291);
nor U12077 (N_12077,N_11351,N_11735);
nand U12078 (N_12078,N_11840,N_11338);
or U12079 (N_12079,N_11860,N_11429);
nand U12080 (N_12080,N_11803,N_11543);
nand U12081 (N_12081,N_11684,N_11530);
nand U12082 (N_12082,N_11807,N_11993);
or U12083 (N_12083,N_11298,N_11805);
xor U12084 (N_12084,N_11445,N_11832);
and U12085 (N_12085,N_11316,N_11420);
and U12086 (N_12086,N_11822,N_11654);
and U12087 (N_12087,N_11259,N_11258);
nand U12088 (N_12088,N_11780,N_11729);
and U12089 (N_12089,N_11260,N_11767);
and U12090 (N_12090,N_11708,N_11906);
nor U12091 (N_12091,N_11711,N_11385);
nor U12092 (N_12092,N_11531,N_11826);
nand U12093 (N_12093,N_11879,N_11414);
nand U12094 (N_12094,N_11407,N_11878);
or U12095 (N_12095,N_11274,N_11349);
nand U12096 (N_12096,N_11756,N_11919);
nand U12097 (N_12097,N_11476,N_11705);
nand U12098 (N_12098,N_11458,N_11495);
nor U12099 (N_12099,N_11405,N_11615);
nor U12100 (N_12100,N_11548,N_11964);
or U12101 (N_12101,N_11462,N_11394);
nor U12102 (N_12102,N_11620,N_11987);
nor U12103 (N_12103,N_11789,N_11343);
or U12104 (N_12104,N_11652,N_11585);
and U12105 (N_12105,N_11538,N_11354);
and U12106 (N_12106,N_11671,N_11744);
and U12107 (N_12107,N_11302,N_11662);
or U12108 (N_12108,N_11681,N_11342);
nor U12109 (N_12109,N_11969,N_11834);
nor U12110 (N_12110,N_11823,N_11892);
or U12111 (N_12111,N_11897,N_11886);
nand U12112 (N_12112,N_11393,N_11930);
xnor U12113 (N_12113,N_11619,N_11691);
xor U12114 (N_12114,N_11719,N_11800);
nand U12115 (N_12115,N_11976,N_11748);
nand U12116 (N_12116,N_11990,N_11573);
xnor U12117 (N_12117,N_11689,N_11816);
or U12118 (N_12118,N_11504,N_11386);
and U12119 (N_12119,N_11454,N_11733);
nor U12120 (N_12120,N_11465,N_11942);
or U12121 (N_12121,N_11938,N_11340);
nor U12122 (N_12122,N_11273,N_11898);
nand U12123 (N_12123,N_11855,N_11704);
nor U12124 (N_12124,N_11895,N_11403);
or U12125 (N_12125,N_11949,N_11650);
and U12126 (N_12126,N_11591,N_11268);
nand U12127 (N_12127,N_11482,N_11502);
xor U12128 (N_12128,N_11837,N_11920);
and U12129 (N_12129,N_11960,N_11682);
or U12130 (N_12130,N_11353,N_11271);
nand U12131 (N_12131,N_11950,N_11945);
or U12132 (N_12132,N_11283,N_11850);
nor U12133 (N_12133,N_11996,N_11738);
or U12134 (N_12134,N_11419,N_11941);
or U12135 (N_12135,N_11865,N_11739);
nand U12136 (N_12136,N_11497,N_11452);
nand U12137 (N_12137,N_11616,N_11603);
nand U12138 (N_12138,N_11762,N_11494);
and U12139 (N_12139,N_11752,N_11974);
nor U12140 (N_12140,N_11821,N_11934);
and U12141 (N_12141,N_11786,N_11776);
nand U12142 (N_12142,N_11534,N_11432);
or U12143 (N_12143,N_11276,N_11388);
or U12144 (N_12144,N_11507,N_11935);
and U12145 (N_12145,N_11383,N_11899);
nand U12146 (N_12146,N_11769,N_11637);
nand U12147 (N_12147,N_11696,N_11307);
and U12148 (N_12148,N_11764,N_11500);
nor U12149 (N_12149,N_11339,N_11422);
or U12150 (N_12150,N_11559,N_11917);
and U12151 (N_12151,N_11980,N_11973);
and U12152 (N_12152,N_11328,N_11581);
and U12153 (N_12153,N_11533,N_11810);
xnor U12154 (N_12154,N_11318,N_11267);
and U12155 (N_12155,N_11341,N_11703);
nor U12156 (N_12156,N_11408,N_11802);
or U12157 (N_12157,N_11625,N_11972);
nor U12158 (N_12158,N_11297,N_11634);
nor U12159 (N_12159,N_11503,N_11643);
or U12160 (N_12160,N_11569,N_11989);
or U12161 (N_12161,N_11373,N_11872);
nor U12162 (N_12162,N_11649,N_11423);
nor U12163 (N_12163,N_11536,N_11921);
or U12164 (N_12164,N_11811,N_11690);
nor U12165 (N_12165,N_11379,N_11606);
nor U12166 (N_12166,N_11459,N_11994);
and U12167 (N_12167,N_11468,N_11639);
and U12168 (N_12168,N_11957,N_11551);
nand U12169 (N_12169,N_11377,N_11522);
nor U12170 (N_12170,N_11457,N_11309);
and U12171 (N_12171,N_11814,N_11958);
xnor U12172 (N_12172,N_11896,N_11982);
nand U12173 (N_12173,N_11390,N_11655);
xor U12174 (N_12174,N_11501,N_11567);
nand U12175 (N_12175,N_11448,N_11322);
or U12176 (N_12176,N_11456,N_11254);
nor U12177 (N_12177,N_11783,N_11284);
and U12178 (N_12178,N_11668,N_11713);
and U12179 (N_12179,N_11392,N_11579);
xnor U12180 (N_12180,N_11925,N_11623);
nand U12181 (N_12181,N_11360,N_11988);
and U12182 (N_12182,N_11558,N_11984);
nor U12183 (N_12183,N_11765,N_11908);
nor U12184 (N_12184,N_11753,N_11527);
nor U12185 (N_12185,N_11401,N_11624);
nor U12186 (N_12186,N_11677,N_11577);
or U12187 (N_12187,N_11927,N_11396);
nor U12188 (N_12188,N_11292,N_11904);
and U12189 (N_12189,N_11888,N_11421);
nand U12190 (N_12190,N_11819,N_11279);
or U12191 (N_12191,N_11701,N_11918);
nor U12192 (N_12192,N_11771,N_11889);
xnor U12193 (N_12193,N_11709,N_11357);
and U12194 (N_12194,N_11329,N_11936);
nor U12195 (N_12195,N_11535,N_11882);
nand U12196 (N_12196,N_11726,N_11966);
and U12197 (N_12197,N_11311,N_11768);
nand U12198 (N_12198,N_11645,N_11876);
nor U12199 (N_12199,N_11479,N_11947);
or U12200 (N_12200,N_11977,N_11347);
nand U12201 (N_12201,N_11467,N_11853);
nor U12202 (N_12202,N_11409,N_11493);
nand U12203 (N_12203,N_11461,N_11692);
and U12204 (N_12204,N_11628,N_11750);
nand U12205 (N_12205,N_11557,N_11453);
or U12206 (N_12206,N_11275,N_11270);
nand U12207 (N_12207,N_11695,N_11358);
and U12208 (N_12208,N_11667,N_11412);
nand U12209 (N_12209,N_11415,N_11841);
and U12210 (N_12210,N_11374,N_11590);
and U12211 (N_12211,N_11397,N_11486);
and U12212 (N_12212,N_11499,N_11256);
nand U12213 (N_12213,N_11505,N_11931);
or U12214 (N_12214,N_11574,N_11545);
nor U12215 (N_12215,N_11277,N_11658);
or U12216 (N_12216,N_11518,N_11325);
nor U12217 (N_12217,N_11755,N_11790);
or U12218 (N_12218,N_11669,N_11387);
or U12219 (N_12219,N_11366,N_11970);
nand U12220 (N_12220,N_11375,N_11317);
xor U12221 (N_12221,N_11352,N_11675);
nor U12222 (N_12222,N_11369,N_11564);
or U12223 (N_12223,N_11736,N_11678);
nand U12224 (N_12224,N_11880,N_11289);
nand U12225 (N_12225,N_11554,N_11290);
and U12226 (N_12226,N_11417,N_11532);
nand U12227 (N_12227,N_11672,N_11849);
nand U12228 (N_12228,N_11582,N_11251);
and U12229 (N_12229,N_11348,N_11720);
nor U12230 (N_12230,N_11477,N_11828);
and U12231 (N_12231,N_11967,N_11299);
nand U12232 (N_12232,N_11700,N_11542);
xnor U12233 (N_12233,N_11361,N_11648);
or U12234 (N_12234,N_11999,N_11846);
and U12235 (N_12235,N_11922,N_11702);
nand U12236 (N_12236,N_11749,N_11282);
or U12237 (N_12237,N_11587,N_11301);
nand U12238 (N_12238,N_11609,N_11263);
nand U12239 (N_12239,N_11875,N_11449);
nor U12240 (N_12240,N_11644,N_11447);
and U12241 (N_12241,N_11571,N_11389);
or U12242 (N_12242,N_11911,N_11679);
and U12243 (N_12243,N_11952,N_11464);
or U12244 (N_12244,N_11661,N_11608);
xnor U12245 (N_12245,N_11699,N_11350);
and U12246 (N_12246,N_11295,N_11961);
and U12247 (N_12247,N_11712,N_11864);
nand U12248 (N_12248,N_11851,N_11485);
nor U12249 (N_12249,N_11664,N_11680);
nor U12250 (N_12250,N_11794,N_11912);
nand U12251 (N_12251,N_11798,N_11635);
nand U12252 (N_12252,N_11928,N_11707);
nand U12253 (N_12253,N_11280,N_11380);
nand U12254 (N_12254,N_11575,N_11718);
xor U12255 (N_12255,N_11929,N_11741);
nor U12256 (N_12256,N_11763,N_11399);
nor U12257 (N_12257,N_11835,N_11725);
nand U12258 (N_12258,N_11562,N_11416);
and U12259 (N_12259,N_11400,N_11281);
and U12260 (N_12260,N_11611,N_11586);
and U12261 (N_12261,N_11869,N_11257);
nor U12262 (N_12262,N_11469,N_11737);
nand U12263 (N_12263,N_11556,N_11376);
and U12264 (N_12264,N_11331,N_11356);
nand U12265 (N_12265,N_11528,N_11742);
and U12266 (N_12266,N_11521,N_11827);
nor U12267 (N_12267,N_11324,N_11640);
nand U12268 (N_12268,N_11365,N_11641);
or U12269 (N_12269,N_11261,N_11657);
or U12270 (N_12270,N_11478,N_11985);
nand U12271 (N_12271,N_11666,N_11867);
nor U12272 (N_12272,N_11323,N_11382);
and U12273 (N_12273,N_11940,N_11642);
or U12274 (N_12274,N_11923,N_11510);
nor U12275 (N_12275,N_11438,N_11552);
and U12276 (N_12276,N_11820,N_11975);
nor U12277 (N_12277,N_11252,N_11428);
nor U12278 (N_12278,N_11326,N_11594);
or U12279 (N_12279,N_11598,N_11817);
and U12280 (N_12280,N_11723,N_11670);
or U12281 (N_12281,N_11916,N_11907);
or U12282 (N_12282,N_11402,N_11656);
nor U12283 (N_12283,N_11496,N_11785);
or U12284 (N_12284,N_11523,N_11793);
or U12285 (N_12285,N_11784,N_11265);
xnor U12286 (N_12286,N_11915,N_11455);
nor U12287 (N_12287,N_11782,N_11859);
or U12288 (N_12288,N_11825,N_11286);
nor U12289 (N_12289,N_11986,N_11436);
nor U12290 (N_12290,N_11605,N_11269);
and U12291 (N_12291,N_11541,N_11766);
and U12292 (N_12292,N_11998,N_11278);
xnor U12293 (N_12293,N_11568,N_11751);
nand U12294 (N_12294,N_11363,N_11686);
nand U12295 (N_12295,N_11481,N_11425);
and U12296 (N_12296,N_11442,N_11333);
xnor U12297 (N_12297,N_11613,N_11861);
and U12298 (N_12298,N_11730,N_11250);
xor U12299 (N_12299,N_11547,N_11877);
or U12300 (N_12300,N_11953,N_11604);
and U12301 (N_12301,N_11868,N_11597);
xnor U12302 (N_12302,N_11570,N_11870);
xor U12303 (N_12303,N_11774,N_11539);
and U12304 (N_12304,N_11646,N_11406);
nand U12305 (N_12305,N_11813,N_11955);
xor U12306 (N_12306,N_11293,N_11717);
nor U12307 (N_12307,N_11937,N_11829);
or U12308 (N_12308,N_11963,N_11344);
and U12309 (N_12309,N_11304,N_11607);
nand U12310 (N_12310,N_11902,N_11513);
nand U12311 (N_12311,N_11600,N_11663);
nand U12312 (N_12312,N_11596,N_11761);
nand U12313 (N_12313,N_11839,N_11332);
and U12314 (N_12314,N_11439,N_11418);
or U12315 (N_12315,N_11515,N_11981);
xor U12316 (N_12316,N_11441,N_11836);
nor U12317 (N_12317,N_11431,N_11954);
or U12318 (N_12318,N_11446,N_11716);
or U12319 (N_12319,N_11843,N_11956);
and U12320 (N_12320,N_11863,N_11472);
nand U12321 (N_12321,N_11519,N_11797);
nand U12322 (N_12322,N_11471,N_11992);
nand U12323 (N_12323,N_11498,N_11924);
nor U12324 (N_12324,N_11914,N_11411);
nand U12325 (N_12325,N_11345,N_11285);
and U12326 (N_12326,N_11747,N_11391);
nand U12327 (N_12327,N_11778,N_11327);
nand U12328 (N_12328,N_11759,N_11885);
or U12329 (N_12329,N_11760,N_11520);
nand U12330 (N_12330,N_11757,N_11788);
nand U12331 (N_12331,N_11288,N_11881);
nand U12332 (N_12332,N_11770,N_11529);
or U12333 (N_12333,N_11595,N_11544);
nand U12334 (N_12334,N_11844,N_11728);
xor U12335 (N_12335,N_11255,N_11506);
xor U12336 (N_12336,N_11470,N_11978);
and U12337 (N_12337,N_11779,N_11773);
nor U12338 (N_12338,N_11443,N_11799);
nor U12339 (N_12339,N_11475,N_11909);
nor U12340 (N_12340,N_11330,N_11404);
xor U12341 (N_12341,N_11546,N_11300);
nor U12342 (N_12342,N_11673,N_11830);
and U12343 (N_12343,N_11866,N_11792);
or U12344 (N_12344,N_11305,N_11602);
xnor U12345 (N_12345,N_11512,N_11746);
nand U12346 (N_12346,N_11308,N_11926);
nor U12347 (N_12347,N_11484,N_11991);
and U12348 (N_12348,N_11592,N_11410);
xnor U12349 (N_12349,N_11294,N_11601);
nand U12350 (N_12350,N_11894,N_11413);
or U12351 (N_12351,N_11745,N_11651);
and U12352 (N_12352,N_11951,N_11636);
and U12353 (N_12353,N_11444,N_11873);
and U12354 (N_12354,N_11310,N_11593);
nand U12355 (N_12355,N_11526,N_11913);
xor U12356 (N_12356,N_11848,N_11910);
nand U12357 (N_12357,N_11370,N_11854);
and U12358 (N_12358,N_11560,N_11463);
and U12359 (N_12359,N_11335,N_11687);
nor U12360 (N_12360,N_11694,N_11862);
and U12361 (N_12361,N_11424,N_11795);
nor U12362 (N_12362,N_11995,N_11884);
and U12363 (N_12363,N_11262,N_11647);
xor U12364 (N_12364,N_11599,N_11815);
or U12365 (N_12365,N_11430,N_11715);
nand U12366 (N_12366,N_11576,N_11433);
or U12367 (N_12367,N_11589,N_11979);
nand U12368 (N_12368,N_11948,N_11266);
nor U12369 (N_12369,N_11731,N_11838);
xnor U12370 (N_12370,N_11893,N_11480);
or U12371 (N_12371,N_11721,N_11809);
and U12372 (N_12372,N_11491,N_11857);
xor U12373 (N_12373,N_11553,N_11427);
and U12374 (N_12374,N_11490,N_11631);
and U12375 (N_12375,N_11357,N_11482);
nor U12376 (N_12376,N_11513,N_11668);
nand U12377 (N_12377,N_11423,N_11814);
nor U12378 (N_12378,N_11270,N_11261);
nand U12379 (N_12379,N_11897,N_11958);
nand U12380 (N_12380,N_11529,N_11307);
nor U12381 (N_12381,N_11271,N_11352);
or U12382 (N_12382,N_11340,N_11575);
nor U12383 (N_12383,N_11692,N_11661);
nor U12384 (N_12384,N_11704,N_11722);
nand U12385 (N_12385,N_11558,N_11661);
nor U12386 (N_12386,N_11990,N_11306);
and U12387 (N_12387,N_11954,N_11619);
and U12388 (N_12388,N_11662,N_11552);
and U12389 (N_12389,N_11394,N_11519);
nor U12390 (N_12390,N_11745,N_11332);
and U12391 (N_12391,N_11782,N_11959);
nor U12392 (N_12392,N_11790,N_11853);
or U12393 (N_12393,N_11874,N_11566);
nor U12394 (N_12394,N_11532,N_11265);
nor U12395 (N_12395,N_11330,N_11703);
nor U12396 (N_12396,N_11292,N_11821);
and U12397 (N_12397,N_11290,N_11266);
and U12398 (N_12398,N_11767,N_11918);
nor U12399 (N_12399,N_11744,N_11688);
nand U12400 (N_12400,N_11643,N_11713);
nand U12401 (N_12401,N_11510,N_11384);
or U12402 (N_12402,N_11437,N_11310);
or U12403 (N_12403,N_11297,N_11583);
and U12404 (N_12404,N_11291,N_11418);
or U12405 (N_12405,N_11464,N_11655);
or U12406 (N_12406,N_11469,N_11280);
nand U12407 (N_12407,N_11774,N_11928);
or U12408 (N_12408,N_11830,N_11967);
xor U12409 (N_12409,N_11405,N_11670);
or U12410 (N_12410,N_11650,N_11723);
and U12411 (N_12411,N_11570,N_11370);
nor U12412 (N_12412,N_11885,N_11999);
or U12413 (N_12413,N_11604,N_11537);
nor U12414 (N_12414,N_11467,N_11766);
nor U12415 (N_12415,N_11411,N_11727);
or U12416 (N_12416,N_11807,N_11605);
or U12417 (N_12417,N_11262,N_11631);
nor U12418 (N_12418,N_11665,N_11383);
or U12419 (N_12419,N_11968,N_11881);
xor U12420 (N_12420,N_11820,N_11908);
nand U12421 (N_12421,N_11356,N_11450);
and U12422 (N_12422,N_11287,N_11399);
or U12423 (N_12423,N_11334,N_11691);
nand U12424 (N_12424,N_11862,N_11617);
or U12425 (N_12425,N_11654,N_11979);
nor U12426 (N_12426,N_11850,N_11925);
xor U12427 (N_12427,N_11827,N_11639);
and U12428 (N_12428,N_11780,N_11849);
or U12429 (N_12429,N_11995,N_11714);
and U12430 (N_12430,N_11564,N_11628);
and U12431 (N_12431,N_11758,N_11919);
or U12432 (N_12432,N_11690,N_11902);
nor U12433 (N_12433,N_11553,N_11974);
nand U12434 (N_12434,N_11712,N_11807);
nor U12435 (N_12435,N_11494,N_11433);
and U12436 (N_12436,N_11800,N_11570);
xnor U12437 (N_12437,N_11338,N_11786);
xnor U12438 (N_12438,N_11352,N_11993);
nor U12439 (N_12439,N_11561,N_11710);
and U12440 (N_12440,N_11279,N_11696);
or U12441 (N_12441,N_11649,N_11663);
nand U12442 (N_12442,N_11993,N_11358);
nor U12443 (N_12443,N_11646,N_11586);
nor U12444 (N_12444,N_11410,N_11713);
xnor U12445 (N_12445,N_11545,N_11570);
nand U12446 (N_12446,N_11759,N_11941);
nand U12447 (N_12447,N_11304,N_11562);
or U12448 (N_12448,N_11524,N_11821);
nor U12449 (N_12449,N_11585,N_11479);
nor U12450 (N_12450,N_11549,N_11559);
nor U12451 (N_12451,N_11819,N_11669);
nor U12452 (N_12452,N_11285,N_11456);
nand U12453 (N_12453,N_11541,N_11829);
and U12454 (N_12454,N_11363,N_11764);
or U12455 (N_12455,N_11891,N_11336);
nor U12456 (N_12456,N_11396,N_11731);
and U12457 (N_12457,N_11768,N_11540);
or U12458 (N_12458,N_11964,N_11687);
nand U12459 (N_12459,N_11334,N_11661);
and U12460 (N_12460,N_11936,N_11558);
and U12461 (N_12461,N_11251,N_11286);
or U12462 (N_12462,N_11732,N_11913);
nand U12463 (N_12463,N_11557,N_11672);
or U12464 (N_12464,N_11346,N_11856);
or U12465 (N_12465,N_11419,N_11261);
nand U12466 (N_12466,N_11629,N_11350);
nor U12467 (N_12467,N_11633,N_11809);
nor U12468 (N_12468,N_11650,N_11958);
nor U12469 (N_12469,N_11887,N_11379);
or U12470 (N_12470,N_11956,N_11701);
or U12471 (N_12471,N_11539,N_11318);
and U12472 (N_12472,N_11292,N_11888);
nor U12473 (N_12473,N_11973,N_11378);
xor U12474 (N_12474,N_11586,N_11989);
nand U12475 (N_12475,N_11893,N_11553);
xnor U12476 (N_12476,N_11276,N_11924);
nand U12477 (N_12477,N_11387,N_11550);
and U12478 (N_12478,N_11755,N_11857);
or U12479 (N_12479,N_11649,N_11264);
or U12480 (N_12480,N_11396,N_11311);
nor U12481 (N_12481,N_11670,N_11855);
or U12482 (N_12482,N_11405,N_11836);
and U12483 (N_12483,N_11795,N_11549);
nor U12484 (N_12484,N_11996,N_11344);
or U12485 (N_12485,N_11729,N_11737);
nand U12486 (N_12486,N_11748,N_11644);
and U12487 (N_12487,N_11833,N_11479);
and U12488 (N_12488,N_11299,N_11446);
nand U12489 (N_12489,N_11463,N_11976);
nor U12490 (N_12490,N_11797,N_11897);
nand U12491 (N_12491,N_11507,N_11530);
xor U12492 (N_12492,N_11321,N_11271);
and U12493 (N_12493,N_11629,N_11705);
xnor U12494 (N_12494,N_11669,N_11473);
nor U12495 (N_12495,N_11548,N_11823);
or U12496 (N_12496,N_11896,N_11331);
nand U12497 (N_12497,N_11682,N_11811);
and U12498 (N_12498,N_11448,N_11390);
nand U12499 (N_12499,N_11920,N_11838);
and U12500 (N_12500,N_11464,N_11603);
nand U12501 (N_12501,N_11889,N_11806);
nand U12502 (N_12502,N_11943,N_11256);
xor U12503 (N_12503,N_11514,N_11768);
and U12504 (N_12504,N_11964,N_11913);
nand U12505 (N_12505,N_11382,N_11708);
or U12506 (N_12506,N_11880,N_11368);
nand U12507 (N_12507,N_11778,N_11807);
or U12508 (N_12508,N_11603,N_11765);
nor U12509 (N_12509,N_11252,N_11423);
or U12510 (N_12510,N_11346,N_11830);
or U12511 (N_12511,N_11564,N_11765);
nand U12512 (N_12512,N_11625,N_11354);
nand U12513 (N_12513,N_11357,N_11965);
or U12514 (N_12514,N_11790,N_11681);
and U12515 (N_12515,N_11897,N_11424);
nand U12516 (N_12516,N_11313,N_11552);
or U12517 (N_12517,N_11956,N_11490);
nor U12518 (N_12518,N_11702,N_11463);
and U12519 (N_12519,N_11810,N_11689);
nand U12520 (N_12520,N_11962,N_11834);
nand U12521 (N_12521,N_11452,N_11639);
or U12522 (N_12522,N_11619,N_11738);
or U12523 (N_12523,N_11678,N_11543);
nor U12524 (N_12524,N_11635,N_11817);
nand U12525 (N_12525,N_11626,N_11717);
and U12526 (N_12526,N_11864,N_11735);
and U12527 (N_12527,N_11727,N_11829);
nand U12528 (N_12528,N_11781,N_11453);
xnor U12529 (N_12529,N_11552,N_11949);
and U12530 (N_12530,N_11618,N_11785);
nand U12531 (N_12531,N_11982,N_11571);
nor U12532 (N_12532,N_11718,N_11806);
nand U12533 (N_12533,N_11954,N_11413);
or U12534 (N_12534,N_11853,N_11619);
xor U12535 (N_12535,N_11343,N_11818);
nor U12536 (N_12536,N_11670,N_11412);
nor U12537 (N_12537,N_11588,N_11468);
xnor U12538 (N_12538,N_11894,N_11616);
nor U12539 (N_12539,N_11506,N_11427);
or U12540 (N_12540,N_11984,N_11749);
nand U12541 (N_12541,N_11908,N_11858);
and U12542 (N_12542,N_11449,N_11796);
xnor U12543 (N_12543,N_11623,N_11882);
and U12544 (N_12544,N_11674,N_11608);
or U12545 (N_12545,N_11576,N_11703);
or U12546 (N_12546,N_11321,N_11989);
xnor U12547 (N_12547,N_11738,N_11674);
and U12548 (N_12548,N_11531,N_11712);
or U12549 (N_12549,N_11527,N_11999);
nor U12550 (N_12550,N_11250,N_11492);
and U12551 (N_12551,N_11604,N_11554);
nor U12552 (N_12552,N_11874,N_11524);
or U12553 (N_12553,N_11985,N_11301);
or U12554 (N_12554,N_11474,N_11859);
or U12555 (N_12555,N_11525,N_11256);
xor U12556 (N_12556,N_11313,N_11643);
or U12557 (N_12557,N_11683,N_11325);
nor U12558 (N_12558,N_11355,N_11499);
and U12559 (N_12559,N_11545,N_11500);
nand U12560 (N_12560,N_11495,N_11662);
or U12561 (N_12561,N_11269,N_11917);
nor U12562 (N_12562,N_11858,N_11292);
nand U12563 (N_12563,N_11294,N_11421);
nor U12564 (N_12564,N_11451,N_11338);
or U12565 (N_12565,N_11666,N_11986);
xor U12566 (N_12566,N_11986,N_11864);
nand U12567 (N_12567,N_11260,N_11428);
nor U12568 (N_12568,N_11966,N_11594);
nand U12569 (N_12569,N_11493,N_11511);
nand U12570 (N_12570,N_11714,N_11879);
and U12571 (N_12571,N_11477,N_11893);
and U12572 (N_12572,N_11910,N_11942);
and U12573 (N_12573,N_11810,N_11463);
nor U12574 (N_12574,N_11635,N_11381);
or U12575 (N_12575,N_11767,N_11281);
or U12576 (N_12576,N_11705,N_11338);
and U12577 (N_12577,N_11535,N_11464);
nand U12578 (N_12578,N_11339,N_11533);
or U12579 (N_12579,N_11277,N_11430);
nor U12580 (N_12580,N_11889,N_11601);
and U12581 (N_12581,N_11696,N_11805);
nor U12582 (N_12582,N_11981,N_11990);
nand U12583 (N_12583,N_11991,N_11680);
or U12584 (N_12584,N_11323,N_11700);
nor U12585 (N_12585,N_11723,N_11661);
and U12586 (N_12586,N_11552,N_11629);
and U12587 (N_12587,N_11645,N_11259);
nor U12588 (N_12588,N_11435,N_11622);
and U12589 (N_12589,N_11269,N_11380);
nor U12590 (N_12590,N_11698,N_11896);
nor U12591 (N_12591,N_11511,N_11541);
nor U12592 (N_12592,N_11724,N_11427);
nor U12593 (N_12593,N_11256,N_11984);
nand U12594 (N_12594,N_11929,N_11802);
nand U12595 (N_12595,N_11706,N_11700);
or U12596 (N_12596,N_11348,N_11702);
nor U12597 (N_12597,N_11579,N_11403);
nand U12598 (N_12598,N_11656,N_11363);
nor U12599 (N_12599,N_11772,N_11897);
and U12600 (N_12600,N_11932,N_11448);
and U12601 (N_12601,N_11634,N_11432);
nor U12602 (N_12602,N_11646,N_11329);
nor U12603 (N_12603,N_11580,N_11636);
and U12604 (N_12604,N_11782,N_11929);
nor U12605 (N_12605,N_11795,N_11765);
or U12606 (N_12606,N_11351,N_11696);
nor U12607 (N_12607,N_11584,N_11285);
nand U12608 (N_12608,N_11701,N_11595);
and U12609 (N_12609,N_11628,N_11836);
and U12610 (N_12610,N_11273,N_11566);
or U12611 (N_12611,N_11296,N_11540);
or U12612 (N_12612,N_11352,N_11428);
or U12613 (N_12613,N_11484,N_11404);
or U12614 (N_12614,N_11404,N_11282);
and U12615 (N_12615,N_11378,N_11487);
and U12616 (N_12616,N_11866,N_11982);
and U12617 (N_12617,N_11607,N_11798);
nand U12618 (N_12618,N_11754,N_11607);
and U12619 (N_12619,N_11623,N_11571);
or U12620 (N_12620,N_11351,N_11517);
nor U12621 (N_12621,N_11314,N_11374);
and U12622 (N_12622,N_11974,N_11679);
nor U12623 (N_12623,N_11826,N_11507);
nor U12624 (N_12624,N_11612,N_11355);
nor U12625 (N_12625,N_11672,N_11789);
nand U12626 (N_12626,N_11322,N_11321);
and U12627 (N_12627,N_11347,N_11566);
xnor U12628 (N_12628,N_11403,N_11331);
nand U12629 (N_12629,N_11270,N_11370);
nand U12630 (N_12630,N_11540,N_11780);
xnor U12631 (N_12631,N_11780,N_11711);
or U12632 (N_12632,N_11560,N_11911);
nor U12633 (N_12633,N_11713,N_11663);
or U12634 (N_12634,N_11869,N_11640);
nor U12635 (N_12635,N_11910,N_11421);
or U12636 (N_12636,N_11889,N_11251);
nor U12637 (N_12637,N_11908,N_11865);
nor U12638 (N_12638,N_11558,N_11722);
and U12639 (N_12639,N_11966,N_11760);
nor U12640 (N_12640,N_11625,N_11664);
nand U12641 (N_12641,N_11862,N_11537);
or U12642 (N_12642,N_11596,N_11392);
nand U12643 (N_12643,N_11264,N_11267);
nor U12644 (N_12644,N_11260,N_11944);
nand U12645 (N_12645,N_11909,N_11549);
nand U12646 (N_12646,N_11749,N_11397);
and U12647 (N_12647,N_11925,N_11653);
nand U12648 (N_12648,N_11311,N_11536);
and U12649 (N_12649,N_11280,N_11927);
nand U12650 (N_12650,N_11501,N_11452);
nand U12651 (N_12651,N_11779,N_11767);
or U12652 (N_12652,N_11787,N_11968);
nand U12653 (N_12653,N_11665,N_11798);
or U12654 (N_12654,N_11387,N_11473);
or U12655 (N_12655,N_11775,N_11277);
and U12656 (N_12656,N_11313,N_11836);
nand U12657 (N_12657,N_11600,N_11261);
xnor U12658 (N_12658,N_11792,N_11304);
xnor U12659 (N_12659,N_11288,N_11961);
nor U12660 (N_12660,N_11433,N_11381);
nand U12661 (N_12661,N_11276,N_11711);
nand U12662 (N_12662,N_11640,N_11574);
nand U12663 (N_12663,N_11345,N_11971);
nand U12664 (N_12664,N_11768,N_11333);
and U12665 (N_12665,N_11907,N_11373);
xor U12666 (N_12666,N_11944,N_11660);
and U12667 (N_12667,N_11613,N_11649);
nor U12668 (N_12668,N_11832,N_11658);
or U12669 (N_12669,N_11275,N_11623);
nor U12670 (N_12670,N_11934,N_11480);
xnor U12671 (N_12671,N_11939,N_11882);
nor U12672 (N_12672,N_11434,N_11256);
nand U12673 (N_12673,N_11441,N_11463);
nor U12674 (N_12674,N_11578,N_11943);
and U12675 (N_12675,N_11694,N_11818);
and U12676 (N_12676,N_11759,N_11954);
xnor U12677 (N_12677,N_11301,N_11277);
xor U12678 (N_12678,N_11442,N_11731);
or U12679 (N_12679,N_11744,N_11530);
nand U12680 (N_12680,N_11364,N_11472);
nor U12681 (N_12681,N_11806,N_11516);
or U12682 (N_12682,N_11921,N_11320);
nand U12683 (N_12683,N_11277,N_11650);
or U12684 (N_12684,N_11784,N_11579);
and U12685 (N_12685,N_11723,N_11499);
nand U12686 (N_12686,N_11680,N_11934);
nand U12687 (N_12687,N_11694,N_11359);
or U12688 (N_12688,N_11949,N_11379);
nand U12689 (N_12689,N_11297,N_11497);
and U12690 (N_12690,N_11997,N_11399);
xor U12691 (N_12691,N_11594,N_11584);
or U12692 (N_12692,N_11552,N_11887);
nand U12693 (N_12693,N_11784,N_11745);
or U12694 (N_12694,N_11987,N_11303);
nand U12695 (N_12695,N_11642,N_11960);
or U12696 (N_12696,N_11597,N_11397);
and U12697 (N_12697,N_11652,N_11489);
nand U12698 (N_12698,N_11963,N_11781);
or U12699 (N_12699,N_11639,N_11731);
nor U12700 (N_12700,N_11843,N_11306);
or U12701 (N_12701,N_11864,N_11797);
and U12702 (N_12702,N_11830,N_11503);
nor U12703 (N_12703,N_11571,N_11991);
nor U12704 (N_12704,N_11916,N_11530);
nor U12705 (N_12705,N_11256,N_11341);
nor U12706 (N_12706,N_11355,N_11967);
and U12707 (N_12707,N_11302,N_11895);
or U12708 (N_12708,N_11281,N_11889);
nand U12709 (N_12709,N_11973,N_11889);
xnor U12710 (N_12710,N_11490,N_11582);
xnor U12711 (N_12711,N_11663,N_11786);
and U12712 (N_12712,N_11626,N_11488);
nor U12713 (N_12713,N_11977,N_11456);
and U12714 (N_12714,N_11618,N_11327);
nand U12715 (N_12715,N_11833,N_11563);
nor U12716 (N_12716,N_11488,N_11481);
and U12717 (N_12717,N_11330,N_11316);
nor U12718 (N_12718,N_11699,N_11567);
nand U12719 (N_12719,N_11713,N_11741);
nand U12720 (N_12720,N_11303,N_11988);
and U12721 (N_12721,N_11842,N_11878);
nor U12722 (N_12722,N_11510,N_11641);
nand U12723 (N_12723,N_11388,N_11319);
nor U12724 (N_12724,N_11767,N_11374);
nand U12725 (N_12725,N_11871,N_11867);
and U12726 (N_12726,N_11755,N_11957);
xor U12727 (N_12727,N_11814,N_11284);
or U12728 (N_12728,N_11694,N_11345);
or U12729 (N_12729,N_11378,N_11792);
or U12730 (N_12730,N_11570,N_11392);
and U12731 (N_12731,N_11616,N_11420);
nor U12732 (N_12732,N_11355,N_11723);
nand U12733 (N_12733,N_11838,N_11284);
nand U12734 (N_12734,N_11951,N_11350);
and U12735 (N_12735,N_11318,N_11392);
or U12736 (N_12736,N_11470,N_11981);
or U12737 (N_12737,N_11476,N_11633);
nand U12738 (N_12738,N_11922,N_11299);
or U12739 (N_12739,N_11840,N_11945);
xor U12740 (N_12740,N_11912,N_11658);
or U12741 (N_12741,N_11805,N_11460);
and U12742 (N_12742,N_11330,N_11953);
nor U12743 (N_12743,N_11843,N_11275);
or U12744 (N_12744,N_11514,N_11638);
and U12745 (N_12745,N_11661,N_11883);
and U12746 (N_12746,N_11486,N_11448);
and U12747 (N_12747,N_11471,N_11631);
xnor U12748 (N_12748,N_11945,N_11406);
and U12749 (N_12749,N_11553,N_11821);
nor U12750 (N_12750,N_12302,N_12013);
and U12751 (N_12751,N_12123,N_12599);
or U12752 (N_12752,N_12426,N_12507);
nand U12753 (N_12753,N_12186,N_12702);
nand U12754 (N_12754,N_12335,N_12205);
nand U12755 (N_12755,N_12533,N_12121);
and U12756 (N_12756,N_12556,N_12655);
and U12757 (N_12757,N_12262,N_12427);
or U12758 (N_12758,N_12707,N_12102);
xnor U12759 (N_12759,N_12404,N_12357);
nand U12760 (N_12760,N_12336,N_12004);
and U12761 (N_12761,N_12483,N_12688);
and U12762 (N_12762,N_12387,N_12429);
or U12763 (N_12763,N_12093,N_12021);
and U12764 (N_12764,N_12647,N_12201);
xnor U12765 (N_12765,N_12396,N_12215);
nor U12766 (N_12766,N_12661,N_12412);
and U12767 (N_12767,N_12731,N_12328);
nand U12768 (N_12768,N_12462,N_12699);
or U12769 (N_12769,N_12484,N_12501);
or U12770 (N_12770,N_12189,N_12146);
nand U12771 (N_12771,N_12385,N_12203);
or U12772 (N_12772,N_12468,N_12208);
nor U12773 (N_12773,N_12026,N_12683);
and U12774 (N_12774,N_12459,N_12452);
nor U12775 (N_12775,N_12508,N_12402);
or U12776 (N_12776,N_12482,N_12515);
nand U12777 (N_12777,N_12155,N_12558);
or U12778 (N_12778,N_12237,N_12517);
and U12779 (N_12779,N_12471,N_12105);
and U12780 (N_12780,N_12294,N_12691);
nand U12781 (N_12781,N_12184,N_12565);
nand U12782 (N_12782,N_12344,N_12143);
or U12783 (N_12783,N_12019,N_12368);
xor U12784 (N_12784,N_12697,N_12187);
and U12785 (N_12785,N_12183,N_12580);
nor U12786 (N_12786,N_12422,N_12420);
xor U12787 (N_12787,N_12418,N_12749);
nor U12788 (N_12788,N_12078,N_12461);
or U12789 (N_12789,N_12561,N_12159);
xor U12790 (N_12790,N_12025,N_12742);
or U12791 (N_12791,N_12126,N_12644);
nor U12792 (N_12792,N_12606,N_12322);
and U12793 (N_12793,N_12236,N_12594);
and U12794 (N_12794,N_12584,N_12235);
or U12795 (N_12795,N_12542,N_12324);
and U12796 (N_12796,N_12612,N_12129);
or U12797 (N_12797,N_12179,N_12127);
nor U12798 (N_12798,N_12704,N_12301);
and U12799 (N_12799,N_12549,N_12695);
or U12800 (N_12800,N_12052,N_12512);
or U12801 (N_12801,N_12477,N_12730);
and U12802 (N_12802,N_12364,N_12180);
and U12803 (N_12803,N_12165,N_12345);
xnor U12804 (N_12804,N_12029,N_12670);
nand U12805 (N_12805,N_12738,N_12632);
xor U12806 (N_12806,N_12496,N_12240);
and U12807 (N_12807,N_12109,N_12592);
or U12808 (N_12808,N_12510,N_12616);
and U12809 (N_12809,N_12652,N_12668);
and U12810 (N_12810,N_12503,N_12638);
nand U12811 (N_12811,N_12544,N_12272);
nand U12812 (N_12812,N_12214,N_12522);
nor U12813 (N_12813,N_12469,N_12227);
or U12814 (N_12814,N_12346,N_12254);
or U12815 (N_12815,N_12411,N_12703);
or U12816 (N_12816,N_12733,N_12329);
or U12817 (N_12817,N_12245,N_12627);
nand U12818 (N_12818,N_12623,N_12488);
nand U12819 (N_12819,N_12168,N_12534);
and U12820 (N_12820,N_12654,N_12167);
nor U12821 (N_12821,N_12048,N_12079);
and U12822 (N_12822,N_12366,N_12395);
nor U12823 (N_12823,N_12154,N_12323);
and U12824 (N_12824,N_12046,N_12247);
or U12825 (N_12825,N_12314,N_12108);
nor U12826 (N_12826,N_12091,N_12000);
nand U12827 (N_12827,N_12511,N_12628);
nor U12828 (N_12828,N_12175,N_12347);
or U12829 (N_12829,N_12225,N_12361);
nor U12830 (N_12830,N_12513,N_12028);
or U12831 (N_12831,N_12111,N_12665);
or U12832 (N_12832,N_12460,N_12113);
nor U12833 (N_12833,N_12660,N_12589);
nor U12834 (N_12834,N_12649,N_12355);
and U12835 (N_12835,N_12257,N_12125);
nor U12836 (N_12836,N_12453,N_12398);
or U12837 (N_12837,N_12475,N_12538);
nand U12838 (N_12838,N_12659,N_12309);
and U12839 (N_12839,N_12497,N_12394);
nand U12840 (N_12840,N_12288,N_12337);
nor U12841 (N_12841,N_12317,N_12626);
and U12842 (N_12842,N_12305,N_12465);
or U12843 (N_12843,N_12122,N_12074);
and U12844 (N_12844,N_12096,N_12249);
and U12845 (N_12845,N_12586,N_12082);
nor U12846 (N_12846,N_12624,N_12198);
nand U12847 (N_12847,N_12284,N_12230);
xor U12848 (N_12848,N_12621,N_12389);
or U12849 (N_12849,N_12173,N_12747);
and U12850 (N_12850,N_12350,N_12372);
or U12851 (N_12851,N_12635,N_12441);
and U12852 (N_12852,N_12409,N_12582);
nand U12853 (N_12853,N_12619,N_12748);
and U12854 (N_12854,N_12566,N_12408);
and U12855 (N_12855,N_12744,N_12149);
nand U12856 (N_12856,N_12213,N_12677);
nand U12857 (N_12857,N_12492,N_12447);
or U12858 (N_12858,N_12466,N_12645);
nand U12859 (N_12859,N_12296,N_12007);
and U12860 (N_12860,N_12015,N_12573);
or U12861 (N_12861,N_12055,N_12439);
and U12862 (N_12862,N_12546,N_12618);
nand U12863 (N_12863,N_12643,N_12410);
nand U12864 (N_12864,N_12233,N_12651);
nor U12865 (N_12865,N_12600,N_12285);
and U12866 (N_12866,N_12040,N_12370);
nor U12867 (N_12867,N_12241,N_12682);
or U12868 (N_12868,N_12119,N_12271);
and U12869 (N_12869,N_12414,N_12058);
and U12870 (N_12870,N_12630,N_12736);
and U12871 (N_12871,N_12014,N_12064);
or U12872 (N_12872,N_12070,N_12253);
xor U12873 (N_12873,N_12326,N_12724);
and U12874 (N_12874,N_12711,N_12564);
and U12875 (N_12875,N_12745,N_12527);
or U12876 (N_12876,N_12338,N_12172);
or U12877 (N_12877,N_12701,N_12110);
xnor U12878 (N_12878,N_12283,N_12428);
nor U12879 (N_12879,N_12151,N_12068);
or U12880 (N_12880,N_12547,N_12056);
nor U12881 (N_12881,N_12210,N_12648);
xnor U12882 (N_12882,N_12476,N_12479);
nor U12883 (N_12883,N_12287,N_12016);
nand U12884 (N_12884,N_12158,N_12024);
nand U12885 (N_12885,N_12552,N_12717);
nand U12886 (N_12886,N_12421,N_12219);
nand U12887 (N_12887,N_12405,N_12693);
nor U12888 (N_12888,N_12473,N_12607);
nand U12889 (N_12889,N_12188,N_12680);
nand U12890 (N_12890,N_12489,N_12737);
nand U12891 (N_12891,N_12746,N_12669);
nor U12892 (N_12892,N_12244,N_12519);
or U12893 (N_12893,N_12434,N_12560);
nor U12894 (N_12894,N_12139,N_12722);
nand U12895 (N_12895,N_12525,N_12185);
and U12896 (N_12896,N_12650,N_12057);
nand U12897 (N_12897,N_12268,N_12281);
nand U12898 (N_12898,N_12332,N_12290);
or U12899 (N_12899,N_12557,N_12521);
or U12900 (N_12900,N_12039,N_12005);
nand U12901 (N_12901,N_12112,N_12243);
and U12902 (N_12902,N_12504,N_12037);
or U12903 (N_12903,N_12279,N_12379);
xnor U12904 (N_12904,N_12231,N_12027);
or U12905 (N_12905,N_12569,N_12474);
nand U12906 (N_12906,N_12406,N_12526);
and U12907 (N_12907,N_12571,N_12339);
nor U12908 (N_12908,N_12207,N_12663);
xnor U12909 (N_12909,N_12356,N_12675);
or U12910 (N_12910,N_12164,N_12424);
nor U12911 (N_12911,N_12615,N_12502);
xnor U12912 (N_12912,N_12725,N_12330);
or U12913 (N_12913,N_12625,N_12353);
or U12914 (N_12914,N_12576,N_12666);
or U12915 (N_12915,N_12178,N_12156);
and U12916 (N_12916,N_12276,N_12059);
and U12917 (N_12917,N_12197,N_12641);
and U12918 (N_12918,N_12147,N_12255);
nand U12919 (N_12919,N_12656,N_12430);
and U12920 (N_12920,N_12587,N_12601);
nor U12921 (N_12921,N_12588,N_12274);
nand U12922 (N_12922,N_12435,N_12226);
nor U12923 (N_12923,N_12509,N_12106);
and U12924 (N_12924,N_12518,N_12516);
nor U12925 (N_12925,N_12449,N_12087);
or U12926 (N_12926,N_12009,N_12712);
or U12927 (N_12927,N_12307,N_12073);
or U12928 (N_12928,N_12354,N_12031);
nand U12929 (N_12929,N_12115,N_12676);
nor U12930 (N_12930,N_12072,N_12554);
nand U12931 (N_12931,N_12721,N_12275);
nand U12932 (N_12932,N_12472,N_12321);
nand U12933 (N_12933,N_12360,N_12690);
or U12934 (N_12934,N_12315,N_12002);
xor U12935 (N_12935,N_12499,N_12609);
nand U12936 (N_12936,N_12218,N_12083);
or U12937 (N_12937,N_12011,N_12673);
nand U12938 (N_12938,N_12559,N_12646);
or U12939 (N_12939,N_12157,N_12256);
nor U12940 (N_12940,N_12351,N_12077);
nor U12941 (N_12941,N_12191,N_12425);
nor U12942 (N_12942,N_12375,N_12708);
and U12943 (N_12943,N_12493,N_12550);
xor U12944 (N_12944,N_12136,N_12206);
and U12945 (N_12945,N_12617,N_12171);
or U12946 (N_12946,N_12685,N_12505);
and U12947 (N_12947,N_12176,N_12678);
nand U12948 (N_12948,N_12563,N_12583);
or U12949 (N_12949,N_12579,N_12034);
and U12950 (N_12950,N_12006,N_12480);
or U12951 (N_12951,N_12694,N_12306);
nand U12952 (N_12952,N_12553,N_12706);
nor U12953 (N_12953,N_12383,N_12313);
and U12954 (N_12954,N_12075,N_12363);
or U12955 (N_12955,N_12239,N_12741);
or U12956 (N_12956,N_12605,N_12597);
and U12957 (N_12957,N_12734,N_12153);
or U12958 (N_12958,N_12090,N_12470);
and U12959 (N_12959,N_12162,N_12367);
nand U12960 (N_12960,N_12388,N_12150);
or U12961 (N_12961,N_12686,N_12085);
and U12962 (N_12962,N_12629,N_12242);
nand U12963 (N_12963,N_12311,N_12467);
nand U12964 (N_12964,N_12101,N_12331);
nor U12965 (N_12965,N_12295,N_12382);
nor U12966 (N_12966,N_12248,N_12494);
and U12967 (N_12967,N_12131,N_12348);
nand U12968 (N_12968,N_12140,N_12376);
and U12969 (N_12969,N_12050,N_12739);
nand U12970 (N_12970,N_12320,N_12442);
nand U12971 (N_12971,N_12523,N_12720);
or U12972 (N_12972,N_12595,N_12174);
or U12973 (N_12973,N_12593,N_12590);
or U12974 (N_12974,N_12327,N_12152);
nand U12975 (N_12975,N_12012,N_12577);
xnor U12976 (N_12976,N_12403,N_12384);
and U12977 (N_12977,N_12018,N_12714);
nor U12978 (N_12978,N_12054,N_12719);
or U12979 (N_12979,N_12674,N_12585);
or U12980 (N_12980,N_12088,N_12228);
nand U12981 (N_12981,N_12478,N_12270);
nand U12982 (N_12982,N_12417,N_12362);
nor U12983 (N_12983,N_12041,N_12099);
nor U12984 (N_12984,N_12535,N_12065);
or U12985 (N_12985,N_12436,N_12610);
nand U12986 (N_12986,N_12551,N_12423);
nor U12987 (N_12987,N_12252,N_12263);
or U12988 (N_12988,N_12141,N_12133);
nor U12989 (N_12989,N_12743,N_12291);
and U12990 (N_12990,N_12581,N_12234);
and U12991 (N_12991,N_12407,N_12575);
and U12992 (N_12992,N_12192,N_12446);
and U12993 (N_12993,N_12092,N_12312);
nand U12994 (N_12994,N_12298,N_12705);
and U12995 (N_12995,N_12325,N_12386);
nand U12996 (N_12996,N_12204,N_12128);
and U12997 (N_12997,N_12570,N_12454);
nand U12998 (N_12998,N_12543,N_12261);
nor U12999 (N_12999,N_12299,N_12445);
and U13000 (N_13000,N_12455,N_12392);
nand U13001 (N_13001,N_12639,N_12653);
and U13002 (N_13002,N_12667,N_12138);
nor U13003 (N_13003,N_12116,N_12144);
xor U13004 (N_13004,N_12578,N_12250);
and U13005 (N_13005,N_12071,N_12698);
or U13006 (N_13006,N_12063,N_12038);
nand U13007 (N_13007,N_12166,N_12278);
and U13008 (N_13008,N_12545,N_12212);
nand U13009 (N_13009,N_12061,N_12568);
nand U13010 (N_13010,N_12642,N_12200);
nand U13011 (N_13011,N_12142,N_12437);
or U13012 (N_13012,N_12199,N_12506);
and U13013 (N_13013,N_12316,N_12319);
and U13014 (N_13014,N_12069,N_12342);
xor U13015 (N_13015,N_12486,N_12022);
nand U13016 (N_13016,N_12514,N_12740);
or U13017 (N_13017,N_12529,N_12267);
nand U13018 (N_13018,N_12491,N_12481);
nand U13019 (N_13019,N_12614,N_12400);
and U13020 (N_13020,N_12067,N_12596);
or U13021 (N_13021,N_12487,N_12051);
or U13022 (N_13022,N_12451,N_12572);
or U13023 (N_13023,N_12035,N_12130);
and U13024 (N_13024,N_12358,N_12224);
or U13025 (N_13025,N_12098,N_12042);
nor U13026 (N_13026,N_12562,N_12008);
nand U13027 (N_13027,N_12397,N_12633);
nor U13028 (N_13028,N_12163,N_12223);
nor U13029 (N_13029,N_12124,N_12097);
and U13030 (N_13030,N_12611,N_12681);
and U13031 (N_13031,N_12377,N_12490);
and U13032 (N_13032,N_12194,N_12602);
and U13033 (N_13033,N_12567,N_12148);
nor U13034 (N_13034,N_12308,N_12555);
nand U13035 (N_13035,N_12132,N_12657);
or U13036 (N_13036,N_12264,N_12293);
xnor U13037 (N_13037,N_12352,N_12463);
or U13038 (N_13038,N_12343,N_12380);
nor U13039 (N_13039,N_12732,N_12456);
or U13040 (N_13040,N_12047,N_12030);
xnor U13041 (N_13041,N_12094,N_12671);
and U13042 (N_13042,N_12443,N_12211);
nor U13043 (N_13043,N_12289,N_12217);
nor U13044 (N_13044,N_12277,N_12003);
nor U13045 (N_13045,N_12729,N_12640);
nand U13046 (N_13046,N_12114,N_12530);
or U13047 (N_13047,N_12341,N_12444);
nand U13048 (N_13048,N_12728,N_12300);
nor U13049 (N_13049,N_12696,N_12292);
nand U13050 (N_13050,N_12232,N_12591);
nor U13051 (N_13051,N_12531,N_12541);
nand U13052 (N_13052,N_12636,N_12251);
nand U13053 (N_13053,N_12726,N_12120);
and U13054 (N_13054,N_12195,N_12620);
nand U13055 (N_13055,N_12169,N_12220);
and U13056 (N_13056,N_12520,N_12723);
nor U13057 (N_13057,N_12622,N_12658);
and U13058 (N_13058,N_12598,N_12374);
and U13059 (N_13059,N_12020,N_12365);
nor U13060 (N_13060,N_12033,N_12340);
or U13061 (N_13061,N_12118,N_12727);
and U13062 (N_13062,N_12303,N_12177);
nor U13063 (N_13063,N_12679,N_12221);
nor U13064 (N_13064,N_12433,N_12349);
and U13065 (N_13065,N_12060,N_12238);
and U13066 (N_13066,N_12381,N_12333);
and U13067 (N_13067,N_12032,N_12608);
nand U13068 (N_13068,N_12161,N_12391);
nand U13069 (N_13069,N_12273,N_12664);
nor U13070 (N_13070,N_12259,N_12464);
or U13071 (N_13071,N_12672,N_12369);
and U13072 (N_13072,N_12457,N_12574);
nor U13073 (N_13073,N_12081,N_12304);
and U13074 (N_13074,N_12604,N_12448);
nor U13075 (N_13075,N_12182,N_12378);
or U13076 (N_13076,N_12202,N_12500);
or U13077 (N_13077,N_12393,N_12297);
xnor U13078 (N_13078,N_12431,N_12222);
or U13079 (N_13079,N_12045,N_12485);
nand U13080 (N_13080,N_12286,N_12181);
nand U13081 (N_13081,N_12359,N_12539);
nand U13082 (N_13082,N_12415,N_12440);
and U13083 (N_13083,N_12498,N_12170);
xnor U13084 (N_13084,N_12036,N_12334);
nor U13085 (N_13085,N_12084,N_12049);
nand U13086 (N_13086,N_12107,N_12100);
nor U13087 (N_13087,N_12246,N_12532);
xor U13088 (N_13088,N_12229,N_12137);
or U13089 (N_13089,N_12548,N_12310);
or U13090 (N_13090,N_12692,N_12715);
and U13091 (N_13091,N_12017,N_12043);
nor U13092 (N_13092,N_12528,N_12432);
nand U13093 (N_13093,N_12117,N_12637);
nor U13094 (N_13094,N_12684,N_12103);
or U13095 (N_13095,N_12689,N_12450);
nor U13096 (N_13096,N_12196,N_12160);
and U13097 (N_13097,N_12145,N_12710);
or U13098 (N_13098,N_12390,N_12023);
nor U13099 (N_13099,N_12419,N_12086);
and U13100 (N_13100,N_12413,N_12416);
nand U13101 (N_13101,N_12265,N_12001);
or U13102 (N_13102,N_12401,N_12134);
xor U13103 (N_13103,N_12318,N_12399);
xnor U13104 (N_13104,N_12631,N_12010);
nand U13105 (N_13105,N_12613,N_12062);
nor U13106 (N_13106,N_12258,N_12716);
or U13107 (N_13107,N_12193,N_12053);
nor U13108 (N_13108,N_12260,N_12718);
and U13109 (N_13109,N_12190,N_12540);
or U13110 (N_13110,N_12080,N_12709);
nand U13111 (N_13111,N_12373,N_12713);
nor U13112 (N_13112,N_12135,N_12536);
and U13113 (N_13113,N_12700,N_12216);
nand U13114 (N_13114,N_12603,N_12537);
or U13115 (N_13115,N_12095,N_12076);
nand U13116 (N_13116,N_12662,N_12269);
and U13117 (N_13117,N_12438,N_12282);
xor U13118 (N_13118,N_12735,N_12687);
xnor U13119 (N_13119,N_12634,N_12495);
nor U13120 (N_13120,N_12371,N_12066);
nor U13121 (N_13121,N_12458,N_12104);
and U13122 (N_13122,N_12524,N_12044);
nor U13123 (N_13123,N_12209,N_12280);
and U13124 (N_13124,N_12089,N_12266);
and U13125 (N_13125,N_12261,N_12110);
nor U13126 (N_13126,N_12740,N_12394);
or U13127 (N_13127,N_12725,N_12338);
xnor U13128 (N_13128,N_12090,N_12512);
or U13129 (N_13129,N_12330,N_12121);
and U13130 (N_13130,N_12590,N_12476);
and U13131 (N_13131,N_12685,N_12235);
and U13132 (N_13132,N_12053,N_12087);
or U13133 (N_13133,N_12206,N_12699);
nand U13134 (N_13134,N_12656,N_12505);
xor U13135 (N_13135,N_12393,N_12595);
or U13136 (N_13136,N_12422,N_12177);
or U13137 (N_13137,N_12138,N_12638);
and U13138 (N_13138,N_12568,N_12152);
nor U13139 (N_13139,N_12310,N_12606);
and U13140 (N_13140,N_12107,N_12118);
or U13141 (N_13141,N_12545,N_12177);
or U13142 (N_13142,N_12165,N_12640);
nor U13143 (N_13143,N_12066,N_12119);
nand U13144 (N_13144,N_12540,N_12041);
nor U13145 (N_13145,N_12327,N_12247);
nand U13146 (N_13146,N_12659,N_12131);
nand U13147 (N_13147,N_12412,N_12007);
or U13148 (N_13148,N_12276,N_12642);
or U13149 (N_13149,N_12544,N_12569);
xor U13150 (N_13150,N_12171,N_12184);
xor U13151 (N_13151,N_12140,N_12044);
and U13152 (N_13152,N_12336,N_12267);
nand U13153 (N_13153,N_12437,N_12672);
and U13154 (N_13154,N_12732,N_12523);
nand U13155 (N_13155,N_12355,N_12521);
and U13156 (N_13156,N_12122,N_12330);
and U13157 (N_13157,N_12176,N_12020);
and U13158 (N_13158,N_12706,N_12697);
nand U13159 (N_13159,N_12577,N_12070);
and U13160 (N_13160,N_12503,N_12530);
and U13161 (N_13161,N_12212,N_12683);
nand U13162 (N_13162,N_12226,N_12165);
or U13163 (N_13163,N_12035,N_12203);
xnor U13164 (N_13164,N_12491,N_12164);
and U13165 (N_13165,N_12710,N_12616);
nor U13166 (N_13166,N_12218,N_12651);
nor U13167 (N_13167,N_12207,N_12007);
and U13168 (N_13168,N_12634,N_12613);
or U13169 (N_13169,N_12534,N_12117);
nand U13170 (N_13170,N_12533,N_12743);
or U13171 (N_13171,N_12309,N_12534);
nand U13172 (N_13172,N_12697,N_12538);
or U13173 (N_13173,N_12230,N_12729);
or U13174 (N_13174,N_12561,N_12317);
and U13175 (N_13175,N_12156,N_12620);
or U13176 (N_13176,N_12211,N_12660);
nand U13177 (N_13177,N_12144,N_12030);
nand U13178 (N_13178,N_12005,N_12631);
xnor U13179 (N_13179,N_12004,N_12107);
or U13180 (N_13180,N_12397,N_12403);
or U13181 (N_13181,N_12160,N_12585);
xnor U13182 (N_13182,N_12602,N_12669);
nor U13183 (N_13183,N_12355,N_12458);
xor U13184 (N_13184,N_12504,N_12300);
or U13185 (N_13185,N_12273,N_12623);
nand U13186 (N_13186,N_12101,N_12355);
nand U13187 (N_13187,N_12444,N_12245);
nand U13188 (N_13188,N_12663,N_12203);
or U13189 (N_13189,N_12102,N_12153);
nand U13190 (N_13190,N_12297,N_12385);
nor U13191 (N_13191,N_12439,N_12192);
or U13192 (N_13192,N_12481,N_12138);
nor U13193 (N_13193,N_12715,N_12710);
nand U13194 (N_13194,N_12542,N_12001);
nand U13195 (N_13195,N_12126,N_12405);
nand U13196 (N_13196,N_12722,N_12496);
and U13197 (N_13197,N_12160,N_12501);
nor U13198 (N_13198,N_12349,N_12062);
or U13199 (N_13199,N_12099,N_12720);
nand U13200 (N_13200,N_12520,N_12659);
nor U13201 (N_13201,N_12092,N_12310);
or U13202 (N_13202,N_12286,N_12415);
nand U13203 (N_13203,N_12292,N_12016);
and U13204 (N_13204,N_12366,N_12348);
or U13205 (N_13205,N_12580,N_12207);
xor U13206 (N_13206,N_12144,N_12703);
or U13207 (N_13207,N_12677,N_12139);
or U13208 (N_13208,N_12037,N_12067);
and U13209 (N_13209,N_12444,N_12000);
nand U13210 (N_13210,N_12158,N_12002);
xor U13211 (N_13211,N_12346,N_12119);
xor U13212 (N_13212,N_12207,N_12558);
and U13213 (N_13213,N_12092,N_12734);
and U13214 (N_13214,N_12087,N_12018);
xor U13215 (N_13215,N_12478,N_12506);
and U13216 (N_13216,N_12122,N_12033);
nor U13217 (N_13217,N_12213,N_12340);
nand U13218 (N_13218,N_12726,N_12192);
nor U13219 (N_13219,N_12436,N_12447);
and U13220 (N_13220,N_12509,N_12288);
or U13221 (N_13221,N_12196,N_12464);
or U13222 (N_13222,N_12693,N_12313);
and U13223 (N_13223,N_12392,N_12677);
nand U13224 (N_13224,N_12134,N_12144);
nand U13225 (N_13225,N_12140,N_12295);
and U13226 (N_13226,N_12048,N_12015);
and U13227 (N_13227,N_12302,N_12554);
nor U13228 (N_13228,N_12586,N_12142);
or U13229 (N_13229,N_12664,N_12245);
nor U13230 (N_13230,N_12707,N_12730);
xor U13231 (N_13231,N_12360,N_12196);
nor U13232 (N_13232,N_12057,N_12149);
or U13233 (N_13233,N_12507,N_12048);
and U13234 (N_13234,N_12375,N_12743);
or U13235 (N_13235,N_12440,N_12136);
xor U13236 (N_13236,N_12006,N_12200);
nand U13237 (N_13237,N_12110,N_12398);
or U13238 (N_13238,N_12085,N_12458);
nand U13239 (N_13239,N_12118,N_12103);
xnor U13240 (N_13240,N_12496,N_12593);
or U13241 (N_13241,N_12239,N_12210);
or U13242 (N_13242,N_12222,N_12306);
nand U13243 (N_13243,N_12039,N_12084);
or U13244 (N_13244,N_12273,N_12736);
nor U13245 (N_13245,N_12250,N_12468);
nor U13246 (N_13246,N_12657,N_12111);
nand U13247 (N_13247,N_12596,N_12563);
nor U13248 (N_13248,N_12065,N_12276);
and U13249 (N_13249,N_12462,N_12292);
nor U13250 (N_13250,N_12499,N_12119);
and U13251 (N_13251,N_12380,N_12044);
nor U13252 (N_13252,N_12406,N_12288);
and U13253 (N_13253,N_12424,N_12658);
or U13254 (N_13254,N_12404,N_12155);
and U13255 (N_13255,N_12701,N_12635);
or U13256 (N_13256,N_12445,N_12114);
or U13257 (N_13257,N_12105,N_12675);
and U13258 (N_13258,N_12618,N_12630);
and U13259 (N_13259,N_12053,N_12471);
or U13260 (N_13260,N_12107,N_12311);
nor U13261 (N_13261,N_12733,N_12504);
and U13262 (N_13262,N_12391,N_12323);
nor U13263 (N_13263,N_12736,N_12472);
nor U13264 (N_13264,N_12034,N_12123);
nand U13265 (N_13265,N_12217,N_12196);
or U13266 (N_13266,N_12334,N_12556);
and U13267 (N_13267,N_12455,N_12224);
nor U13268 (N_13268,N_12488,N_12172);
nor U13269 (N_13269,N_12681,N_12070);
and U13270 (N_13270,N_12060,N_12158);
nand U13271 (N_13271,N_12612,N_12281);
nor U13272 (N_13272,N_12638,N_12352);
and U13273 (N_13273,N_12158,N_12346);
nor U13274 (N_13274,N_12239,N_12225);
nor U13275 (N_13275,N_12338,N_12096);
nor U13276 (N_13276,N_12728,N_12394);
and U13277 (N_13277,N_12415,N_12042);
or U13278 (N_13278,N_12111,N_12496);
nor U13279 (N_13279,N_12383,N_12134);
and U13280 (N_13280,N_12451,N_12641);
or U13281 (N_13281,N_12612,N_12731);
nor U13282 (N_13282,N_12592,N_12547);
xor U13283 (N_13283,N_12491,N_12008);
and U13284 (N_13284,N_12478,N_12108);
nand U13285 (N_13285,N_12055,N_12307);
nor U13286 (N_13286,N_12098,N_12029);
or U13287 (N_13287,N_12272,N_12330);
and U13288 (N_13288,N_12284,N_12058);
or U13289 (N_13289,N_12729,N_12409);
nor U13290 (N_13290,N_12726,N_12226);
nor U13291 (N_13291,N_12540,N_12402);
or U13292 (N_13292,N_12126,N_12323);
xnor U13293 (N_13293,N_12464,N_12447);
or U13294 (N_13294,N_12536,N_12518);
or U13295 (N_13295,N_12624,N_12610);
nand U13296 (N_13296,N_12635,N_12160);
xnor U13297 (N_13297,N_12282,N_12530);
or U13298 (N_13298,N_12398,N_12170);
or U13299 (N_13299,N_12079,N_12601);
nor U13300 (N_13300,N_12404,N_12419);
xnor U13301 (N_13301,N_12532,N_12651);
nand U13302 (N_13302,N_12054,N_12541);
nand U13303 (N_13303,N_12622,N_12529);
nor U13304 (N_13304,N_12613,N_12679);
or U13305 (N_13305,N_12681,N_12058);
nor U13306 (N_13306,N_12356,N_12105);
xor U13307 (N_13307,N_12598,N_12019);
or U13308 (N_13308,N_12575,N_12409);
or U13309 (N_13309,N_12200,N_12185);
nand U13310 (N_13310,N_12182,N_12533);
and U13311 (N_13311,N_12558,N_12225);
nand U13312 (N_13312,N_12162,N_12667);
or U13313 (N_13313,N_12635,N_12532);
and U13314 (N_13314,N_12022,N_12096);
and U13315 (N_13315,N_12034,N_12552);
nor U13316 (N_13316,N_12116,N_12231);
nand U13317 (N_13317,N_12270,N_12746);
and U13318 (N_13318,N_12048,N_12406);
or U13319 (N_13319,N_12699,N_12323);
and U13320 (N_13320,N_12653,N_12097);
and U13321 (N_13321,N_12512,N_12575);
or U13322 (N_13322,N_12041,N_12586);
and U13323 (N_13323,N_12505,N_12159);
and U13324 (N_13324,N_12305,N_12429);
and U13325 (N_13325,N_12529,N_12235);
xor U13326 (N_13326,N_12448,N_12345);
and U13327 (N_13327,N_12548,N_12248);
or U13328 (N_13328,N_12531,N_12230);
or U13329 (N_13329,N_12446,N_12531);
nor U13330 (N_13330,N_12745,N_12653);
nor U13331 (N_13331,N_12175,N_12440);
xnor U13332 (N_13332,N_12101,N_12271);
and U13333 (N_13333,N_12579,N_12677);
or U13334 (N_13334,N_12179,N_12332);
nand U13335 (N_13335,N_12122,N_12515);
or U13336 (N_13336,N_12384,N_12389);
or U13337 (N_13337,N_12185,N_12549);
and U13338 (N_13338,N_12107,N_12192);
or U13339 (N_13339,N_12408,N_12503);
nor U13340 (N_13340,N_12412,N_12299);
nor U13341 (N_13341,N_12497,N_12093);
and U13342 (N_13342,N_12621,N_12694);
nand U13343 (N_13343,N_12157,N_12372);
or U13344 (N_13344,N_12014,N_12112);
and U13345 (N_13345,N_12172,N_12651);
and U13346 (N_13346,N_12202,N_12673);
and U13347 (N_13347,N_12613,N_12650);
nor U13348 (N_13348,N_12014,N_12474);
nor U13349 (N_13349,N_12280,N_12661);
and U13350 (N_13350,N_12060,N_12318);
nor U13351 (N_13351,N_12009,N_12149);
or U13352 (N_13352,N_12104,N_12146);
xnor U13353 (N_13353,N_12176,N_12578);
nand U13354 (N_13354,N_12545,N_12178);
nand U13355 (N_13355,N_12130,N_12510);
and U13356 (N_13356,N_12549,N_12737);
and U13357 (N_13357,N_12629,N_12493);
nor U13358 (N_13358,N_12435,N_12736);
nor U13359 (N_13359,N_12541,N_12612);
nor U13360 (N_13360,N_12650,N_12251);
or U13361 (N_13361,N_12536,N_12579);
nor U13362 (N_13362,N_12618,N_12432);
or U13363 (N_13363,N_12069,N_12010);
nand U13364 (N_13364,N_12530,N_12115);
nand U13365 (N_13365,N_12243,N_12356);
and U13366 (N_13366,N_12347,N_12745);
nor U13367 (N_13367,N_12609,N_12551);
nor U13368 (N_13368,N_12246,N_12549);
nand U13369 (N_13369,N_12060,N_12682);
xnor U13370 (N_13370,N_12201,N_12161);
xnor U13371 (N_13371,N_12360,N_12705);
or U13372 (N_13372,N_12198,N_12340);
nor U13373 (N_13373,N_12665,N_12737);
xor U13374 (N_13374,N_12328,N_12178);
nand U13375 (N_13375,N_12744,N_12266);
xnor U13376 (N_13376,N_12386,N_12085);
and U13377 (N_13377,N_12643,N_12331);
and U13378 (N_13378,N_12705,N_12163);
nand U13379 (N_13379,N_12256,N_12045);
nor U13380 (N_13380,N_12499,N_12347);
nand U13381 (N_13381,N_12112,N_12593);
xnor U13382 (N_13382,N_12704,N_12738);
xnor U13383 (N_13383,N_12063,N_12613);
and U13384 (N_13384,N_12174,N_12050);
nor U13385 (N_13385,N_12462,N_12213);
nand U13386 (N_13386,N_12636,N_12220);
and U13387 (N_13387,N_12296,N_12569);
nor U13388 (N_13388,N_12685,N_12664);
nor U13389 (N_13389,N_12183,N_12594);
nor U13390 (N_13390,N_12260,N_12053);
and U13391 (N_13391,N_12627,N_12730);
and U13392 (N_13392,N_12310,N_12518);
or U13393 (N_13393,N_12333,N_12388);
nor U13394 (N_13394,N_12198,N_12488);
and U13395 (N_13395,N_12425,N_12289);
nand U13396 (N_13396,N_12737,N_12183);
xor U13397 (N_13397,N_12313,N_12447);
nor U13398 (N_13398,N_12254,N_12333);
nor U13399 (N_13399,N_12624,N_12292);
nor U13400 (N_13400,N_12321,N_12388);
nand U13401 (N_13401,N_12627,N_12122);
and U13402 (N_13402,N_12213,N_12599);
nor U13403 (N_13403,N_12107,N_12653);
nor U13404 (N_13404,N_12276,N_12049);
and U13405 (N_13405,N_12008,N_12264);
xor U13406 (N_13406,N_12425,N_12430);
nand U13407 (N_13407,N_12619,N_12224);
nor U13408 (N_13408,N_12075,N_12188);
nand U13409 (N_13409,N_12580,N_12730);
xor U13410 (N_13410,N_12724,N_12610);
and U13411 (N_13411,N_12112,N_12383);
nor U13412 (N_13412,N_12070,N_12573);
and U13413 (N_13413,N_12120,N_12354);
and U13414 (N_13414,N_12103,N_12405);
and U13415 (N_13415,N_12006,N_12374);
xor U13416 (N_13416,N_12688,N_12061);
nand U13417 (N_13417,N_12438,N_12310);
xor U13418 (N_13418,N_12176,N_12179);
xor U13419 (N_13419,N_12491,N_12749);
or U13420 (N_13420,N_12350,N_12050);
and U13421 (N_13421,N_12575,N_12626);
or U13422 (N_13422,N_12185,N_12456);
and U13423 (N_13423,N_12237,N_12613);
and U13424 (N_13424,N_12365,N_12241);
nor U13425 (N_13425,N_12711,N_12493);
or U13426 (N_13426,N_12721,N_12267);
xor U13427 (N_13427,N_12095,N_12279);
xor U13428 (N_13428,N_12599,N_12169);
or U13429 (N_13429,N_12529,N_12645);
or U13430 (N_13430,N_12186,N_12664);
nor U13431 (N_13431,N_12399,N_12021);
and U13432 (N_13432,N_12217,N_12233);
nand U13433 (N_13433,N_12666,N_12690);
nor U13434 (N_13434,N_12371,N_12708);
and U13435 (N_13435,N_12445,N_12449);
nor U13436 (N_13436,N_12237,N_12099);
or U13437 (N_13437,N_12560,N_12220);
nor U13438 (N_13438,N_12094,N_12432);
and U13439 (N_13439,N_12440,N_12521);
or U13440 (N_13440,N_12743,N_12139);
nor U13441 (N_13441,N_12408,N_12476);
and U13442 (N_13442,N_12527,N_12697);
nor U13443 (N_13443,N_12110,N_12038);
nand U13444 (N_13444,N_12735,N_12406);
nand U13445 (N_13445,N_12027,N_12338);
and U13446 (N_13446,N_12532,N_12693);
and U13447 (N_13447,N_12530,N_12606);
nor U13448 (N_13448,N_12210,N_12469);
nand U13449 (N_13449,N_12400,N_12390);
xnor U13450 (N_13450,N_12214,N_12241);
nor U13451 (N_13451,N_12080,N_12103);
and U13452 (N_13452,N_12585,N_12651);
xnor U13453 (N_13453,N_12326,N_12462);
xnor U13454 (N_13454,N_12062,N_12014);
nand U13455 (N_13455,N_12073,N_12690);
and U13456 (N_13456,N_12306,N_12200);
nand U13457 (N_13457,N_12418,N_12313);
nand U13458 (N_13458,N_12725,N_12243);
or U13459 (N_13459,N_12117,N_12044);
nor U13460 (N_13460,N_12529,N_12205);
and U13461 (N_13461,N_12434,N_12646);
nor U13462 (N_13462,N_12251,N_12130);
and U13463 (N_13463,N_12023,N_12455);
nand U13464 (N_13464,N_12576,N_12507);
nand U13465 (N_13465,N_12671,N_12064);
nand U13466 (N_13466,N_12418,N_12330);
nand U13467 (N_13467,N_12325,N_12686);
nand U13468 (N_13468,N_12252,N_12192);
nand U13469 (N_13469,N_12680,N_12654);
nor U13470 (N_13470,N_12592,N_12598);
nor U13471 (N_13471,N_12333,N_12173);
nor U13472 (N_13472,N_12653,N_12443);
and U13473 (N_13473,N_12722,N_12240);
nand U13474 (N_13474,N_12342,N_12084);
and U13475 (N_13475,N_12678,N_12353);
and U13476 (N_13476,N_12053,N_12586);
or U13477 (N_13477,N_12690,N_12456);
nor U13478 (N_13478,N_12479,N_12699);
and U13479 (N_13479,N_12019,N_12639);
nor U13480 (N_13480,N_12672,N_12070);
nor U13481 (N_13481,N_12464,N_12251);
nand U13482 (N_13482,N_12675,N_12107);
xor U13483 (N_13483,N_12125,N_12065);
xor U13484 (N_13484,N_12217,N_12194);
nor U13485 (N_13485,N_12460,N_12652);
and U13486 (N_13486,N_12114,N_12351);
or U13487 (N_13487,N_12132,N_12116);
nor U13488 (N_13488,N_12198,N_12715);
nor U13489 (N_13489,N_12362,N_12307);
and U13490 (N_13490,N_12565,N_12230);
and U13491 (N_13491,N_12293,N_12559);
and U13492 (N_13492,N_12067,N_12538);
nand U13493 (N_13493,N_12649,N_12477);
nor U13494 (N_13494,N_12248,N_12618);
xor U13495 (N_13495,N_12257,N_12669);
and U13496 (N_13496,N_12409,N_12299);
or U13497 (N_13497,N_12564,N_12673);
xnor U13498 (N_13498,N_12023,N_12525);
and U13499 (N_13499,N_12417,N_12621);
nand U13500 (N_13500,N_12892,N_13163);
nand U13501 (N_13501,N_12842,N_13322);
and U13502 (N_13502,N_13339,N_12979);
xor U13503 (N_13503,N_13490,N_12929);
nand U13504 (N_13504,N_12914,N_13164);
and U13505 (N_13505,N_13073,N_13055);
nand U13506 (N_13506,N_13401,N_12829);
nor U13507 (N_13507,N_13469,N_13483);
nor U13508 (N_13508,N_13039,N_13146);
nand U13509 (N_13509,N_12793,N_13109);
nor U13510 (N_13510,N_12881,N_13162);
and U13511 (N_13511,N_13279,N_13212);
nor U13512 (N_13512,N_13052,N_12805);
nor U13513 (N_13513,N_13048,N_12977);
or U13514 (N_13514,N_12893,N_13411);
and U13515 (N_13515,N_12798,N_12984);
or U13516 (N_13516,N_13463,N_13256);
and U13517 (N_13517,N_13203,N_13101);
or U13518 (N_13518,N_12757,N_13107);
xnor U13519 (N_13519,N_13333,N_13278);
or U13520 (N_13520,N_13229,N_13417);
and U13521 (N_13521,N_13042,N_13307);
nand U13522 (N_13522,N_13443,N_13481);
xnor U13523 (N_13523,N_13065,N_13239);
nand U13524 (N_13524,N_13420,N_12775);
nand U13525 (N_13525,N_13200,N_13072);
and U13526 (N_13526,N_12817,N_13398);
or U13527 (N_13527,N_12996,N_13087);
xnor U13528 (N_13528,N_13059,N_12751);
or U13529 (N_13529,N_12951,N_12788);
nand U13530 (N_13530,N_13306,N_12944);
nor U13531 (N_13531,N_12774,N_13134);
nand U13532 (N_13532,N_12916,N_13110);
nor U13533 (N_13533,N_13216,N_12981);
or U13534 (N_13534,N_13232,N_13040);
or U13535 (N_13535,N_13044,N_12867);
xnor U13536 (N_13536,N_12839,N_12763);
and U13537 (N_13537,N_12935,N_12973);
and U13538 (N_13538,N_13159,N_13319);
and U13539 (N_13539,N_12772,N_13067);
nand U13540 (N_13540,N_13453,N_12807);
nand U13541 (N_13541,N_13121,N_12771);
nor U13542 (N_13542,N_13317,N_12761);
nand U13543 (N_13543,N_13284,N_13340);
nor U13544 (N_13544,N_13103,N_12808);
and U13545 (N_13545,N_13379,N_13201);
or U13546 (N_13546,N_13427,N_13156);
nand U13547 (N_13547,N_13371,N_12803);
xnor U13548 (N_13548,N_13020,N_13428);
and U13549 (N_13549,N_13387,N_13309);
and U13550 (N_13550,N_13181,N_12928);
nor U13551 (N_13551,N_12899,N_13178);
nor U13552 (N_13552,N_13051,N_13061);
nand U13553 (N_13553,N_13118,N_13021);
and U13554 (N_13554,N_12844,N_13403);
and U13555 (N_13555,N_13258,N_13358);
and U13556 (N_13556,N_13184,N_12965);
and U13557 (N_13557,N_12989,N_12957);
nand U13558 (N_13558,N_12870,N_13288);
or U13559 (N_13559,N_13083,N_13115);
xnor U13560 (N_13560,N_13179,N_13138);
nand U13561 (N_13561,N_13347,N_12864);
nand U13562 (N_13562,N_13125,N_12851);
xor U13563 (N_13563,N_13262,N_12858);
xor U13564 (N_13564,N_12953,N_12974);
or U13565 (N_13565,N_12826,N_13384);
or U13566 (N_13566,N_13244,N_12868);
and U13567 (N_13567,N_13257,N_13252);
nor U13568 (N_13568,N_12938,N_13356);
and U13569 (N_13569,N_13094,N_13058);
xnor U13570 (N_13570,N_13374,N_13311);
or U13571 (N_13571,N_13402,N_12980);
xnor U13572 (N_13572,N_13108,N_13376);
and U13573 (N_13573,N_13189,N_13165);
nor U13574 (N_13574,N_13018,N_13167);
nor U13575 (N_13575,N_12891,N_13003);
nor U13576 (N_13576,N_13476,N_12784);
or U13577 (N_13577,N_12945,N_13260);
and U13578 (N_13578,N_13283,N_12919);
nor U13579 (N_13579,N_13082,N_13194);
xor U13580 (N_13580,N_13495,N_12838);
nor U13581 (N_13581,N_13272,N_12832);
nand U13582 (N_13582,N_12880,N_13188);
or U13583 (N_13583,N_13460,N_13173);
nor U13584 (N_13584,N_12863,N_13038);
and U13585 (N_13585,N_13360,N_12913);
and U13586 (N_13586,N_12926,N_13001);
nand U13587 (N_13587,N_12950,N_13393);
nor U13588 (N_13588,N_13486,N_12835);
and U13589 (N_13589,N_13046,N_13197);
and U13590 (N_13590,N_13015,N_13049);
xnor U13591 (N_13591,N_13350,N_13177);
xnor U13592 (N_13592,N_13354,N_12836);
and U13593 (N_13593,N_12810,N_13458);
nand U13594 (N_13594,N_13171,N_13412);
nand U13595 (N_13595,N_13474,N_13351);
or U13596 (N_13596,N_12906,N_12966);
xnor U13597 (N_13597,N_12990,N_13274);
nand U13598 (N_13598,N_12876,N_12949);
or U13599 (N_13599,N_12811,N_12831);
xnor U13600 (N_13600,N_12960,N_12964);
and U13601 (N_13601,N_13170,N_12954);
nand U13602 (N_13602,N_13445,N_12779);
and U13603 (N_13603,N_13310,N_12904);
or U13604 (N_13604,N_13142,N_13424);
nand U13605 (N_13605,N_13405,N_13346);
xnor U13606 (N_13606,N_12952,N_12959);
and U13607 (N_13607,N_13105,N_13033);
nor U13608 (N_13608,N_13377,N_13247);
or U13609 (N_13609,N_13098,N_13185);
nand U13610 (N_13610,N_13192,N_12795);
nand U13611 (N_13611,N_13468,N_12909);
and U13612 (N_13612,N_12777,N_13432);
nor U13613 (N_13613,N_12879,N_12875);
nand U13614 (N_13614,N_13023,N_12872);
or U13615 (N_13615,N_12985,N_13395);
and U13616 (N_13616,N_12902,N_13012);
and U13617 (N_13617,N_13367,N_12903);
nor U13618 (N_13618,N_13246,N_13375);
or U13619 (N_13619,N_12886,N_12961);
xnor U13620 (N_13620,N_12998,N_13030);
xnor U13621 (N_13621,N_13491,N_13263);
and U13622 (N_13622,N_13440,N_12820);
xor U13623 (N_13623,N_12895,N_13074);
nand U13624 (N_13624,N_13353,N_13066);
and U13625 (N_13625,N_12758,N_13022);
or U13626 (N_13626,N_13243,N_13352);
and U13627 (N_13627,N_13210,N_13092);
or U13628 (N_13628,N_12764,N_12806);
or U13629 (N_13629,N_13457,N_12927);
and U13630 (N_13630,N_13464,N_13472);
or U13631 (N_13631,N_13480,N_13010);
or U13632 (N_13632,N_13282,N_12991);
xor U13633 (N_13633,N_13102,N_13099);
and U13634 (N_13634,N_12994,N_12753);
and U13635 (N_13635,N_12766,N_13323);
nor U13636 (N_13636,N_13080,N_13426);
and U13637 (N_13637,N_13116,N_13295);
and U13638 (N_13638,N_13123,N_12871);
nand U13639 (N_13639,N_13315,N_13085);
xor U13640 (N_13640,N_13289,N_13029);
nor U13641 (N_13641,N_13470,N_13209);
or U13642 (N_13642,N_12920,N_13122);
and U13643 (N_13643,N_13429,N_13357);
xnor U13644 (N_13644,N_12900,N_12971);
nand U13645 (N_13645,N_12988,N_13242);
or U13646 (N_13646,N_13235,N_13435);
nor U13647 (N_13647,N_12816,N_12796);
nor U13648 (N_13648,N_13112,N_13070);
and U13649 (N_13649,N_12931,N_12941);
nand U13650 (N_13650,N_13459,N_13220);
or U13651 (N_13651,N_12780,N_13397);
or U13652 (N_13652,N_13409,N_12877);
xnor U13653 (N_13653,N_13226,N_13026);
and U13654 (N_13654,N_13245,N_12759);
nand U13655 (N_13655,N_12947,N_13349);
nand U13656 (N_13656,N_12910,N_12815);
nor U13657 (N_13657,N_13373,N_13016);
nor U13658 (N_13658,N_13413,N_13117);
nand U13659 (N_13659,N_13485,N_13191);
or U13660 (N_13660,N_13318,N_13380);
nor U13661 (N_13661,N_13293,N_13433);
nand U13662 (N_13662,N_13305,N_13314);
nor U13663 (N_13663,N_13372,N_13008);
nor U13664 (N_13664,N_13063,N_13251);
or U13665 (N_13665,N_13449,N_13407);
or U13666 (N_13666,N_13487,N_13498);
and U13667 (N_13667,N_13456,N_13136);
nor U13668 (N_13668,N_13286,N_12992);
nand U13669 (N_13669,N_12856,N_13054);
xor U13670 (N_13670,N_13215,N_13187);
xnor U13671 (N_13671,N_13013,N_12888);
or U13672 (N_13672,N_12915,N_13005);
and U13673 (N_13673,N_13439,N_13430);
and U13674 (N_13674,N_13285,N_13114);
nand U13675 (N_13675,N_12783,N_12781);
nand U13676 (N_13676,N_13205,N_13471);
and U13677 (N_13677,N_13148,N_13280);
or U13678 (N_13678,N_13275,N_12857);
and U13679 (N_13679,N_13062,N_13477);
and U13680 (N_13680,N_12969,N_12995);
nor U13681 (N_13681,N_13499,N_13277);
or U13682 (N_13682,N_13330,N_13154);
or U13683 (N_13683,N_13180,N_12855);
xnor U13684 (N_13684,N_13331,N_13291);
nand U13685 (N_13685,N_13097,N_12850);
or U13686 (N_13686,N_12978,N_13004);
or U13687 (N_13687,N_13488,N_13450);
and U13688 (N_13688,N_12897,N_13338);
nor U13689 (N_13689,N_13096,N_12801);
nand U13690 (N_13690,N_13240,N_13497);
nand U13691 (N_13691,N_12770,N_12921);
nand U13692 (N_13692,N_13287,N_13176);
xnor U13693 (N_13693,N_13128,N_13035);
or U13694 (N_13694,N_12962,N_13104);
nor U13695 (N_13695,N_13151,N_13133);
or U13696 (N_13696,N_12885,N_13382);
and U13697 (N_13697,N_13166,N_12830);
xor U13698 (N_13698,N_13423,N_12804);
nor U13699 (N_13699,N_12787,N_12976);
nand U13700 (N_13700,N_13335,N_12948);
nand U13701 (N_13701,N_13452,N_12939);
or U13702 (N_13702,N_13182,N_13190);
or U13703 (N_13703,N_12760,N_13391);
and U13704 (N_13704,N_12776,N_13392);
and U13705 (N_13705,N_12756,N_13479);
or U13706 (N_13706,N_13208,N_13320);
and U13707 (N_13707,N_13011,N_13047);
or U13708 (N_13708,N_13223,N_12861);
nand U13709 (N_13709,N_12912,N_13213);
or U13710 (N_13710,N_13196,N_12849);
and U13711 (N_13711,N_13489,N_13301);
nor U13712 (N_13712,N_12987,N_13292);
and U13713 (N_13713,N_13219,N_13045);
or U13714 (N_13714,N_13363,N_13169);
and U13715 (N_13715,N_12799,N_12778);
nor U13716 (N_13716,N_13057,N_12917);
or U13717 (N_13717,N_13365,N_13378);
nand U13718 (N_13718,N_12896,N_13345);
nor U13719 (N_13719,N_12814,N_12789);
and U13720 (N_13720,N_13294,N_12946);
and U13721 (N_13721,N_13086,N_13091);
or U13722 (N_13722,N_13172,N_12852);
nand U13723 (N_13723,N_13084,N_12866);
nand U13724 (N_13724,N_12827,N_13484);
nor U13725 (N_13725,N_13032,N_12818);
nor U13726 (N_13726,N_13462,N_13271);
xnor U13727 (N_13727,N_13264,N_13493);
and U13728 (N_13728,N_13467,N_13312);
or U13729 (N_13729,N_13473,N_13466);
and U13730 (N_13730,N_13076,N_12802);
and U13731 (N_13731,N_13144,N_13227);
or U13732 (N_13732,N_12889,N_13124);
nor U13733 (N_13733,N_13024,N_13406);
xnor U13734 (N_13734,N_13408,N_12834);
and U13735 (N_13735,N_13475,N_12873);
and U13736 (N_13736,N_13079,N_13036);
nand U13737 (N_13737,N_13233,N_13075);
nand U13738 (N_13738,N_13389,N_13451);
xnor U13739 (N_13739,N_13211,N_13043);
nand U13740 (N_13740,N_13225,N_12932);
and U13741 (N_13741,N_12792,N_13017);
or U13742 (N_13742,N_13119,N_12845);
xnor U13743 (N_13743,N_13214,N_12812);
nand U13744 (N_13744,N_13168,N_13071);
and U13745 (N_13745,N_12933,N_12983);
and U13746 (N_13746,N_13230,N_13465);
nor U13747 (N_13747,N_13081,N_13364);
xnor U13748 (N_13748,N_13217,N_13090);
nand U13749 (N_13749,N_12955,N_13361);
nor U13750 (N_13750,N_13231,N_12773);
or U13751 (N_13751,N_12821,N_13348);
or U13752 (N_13752,N_13383,N_12882);
nand U13753 (N_13753,N_13228,N_12755);
nand U13754 (N_13754,N_13496,N_13425);
xor U13755 (N_13755,N_13369,N_12970);
nand U13756 (N_13756,N_13328,N_12794);
nand U13757 (N_13757,N_12786,N_12894);
or U13758 (N_13758,N_13132,N_13069);
nand U13759 (N_13759,N_13158,N_13131);
nand U13760 (N_13760,N_13206,N_12824);
nor U13761 (N_13761,N_12828,N_13366);
or U13762 (N_13762,N_13290,N_12848);
xnor U13763 (N_13763,N_12924,N_13434);
or U13764 (N_13764,N_13334,N_12887);
and U13765 (N_13765,N_12853,N_13400);
nor U13766 (N_13766,N_12840,N_13207);
or U13767 (N_13767,N_13135,N_12769);
nor U13768 (N_13768,N_13183,N_13031);
or U13769 (N_13769,N_13325,N_12934);
and U13770 (N_13770,N_13269,N_13198);
nand U13771 (N_13771,N_13381,N_13193);
and U13772 (N_13772,N_12762,N_12767);
or U13773 (N_13773,N_12901,N_13028);
nor U13774 (N_13774,N_13053,N_13149);
or U13775 (N_13775,N_12754,N_13002);
xnor U13776 (N_13776,N_13019,N_13129);
nand U13777 (N_13777,N_13273,N_12823);
nor U13778 (N_13778,N_13009,N_13237);
and U13779 (N_13779,N_12956,N_13438);
and U13780 (N_13780,N_13140,N_13095);
and U13781 (N_13781,N_13088,N_12993);
and U13782 (N_13782,N_13419,N_13064);
nor U13783 (N_13783,N_13386,N_13414);
or U13784 (N_13784,N_13204,N_12898);
xor U13785 (N_13785,N_12943,N_12822);
and U13786 (N_13786,N_12765,N_12800);
or U13787 (N_13787,N_13308,N_13078);
nand U13788 (N_13788,N_13482,N_12874);
or U13789 (N_13789,N_12968,N_13337);
nor U13790 (N_13790,N_12813,N_13344);
nor U13791 (N_13791,N_13446,N_12847);
nand U13792 (N_13792,N_13000,N_13130);
nor U13793 (N_13793,N_12972,N_13410);
nand U13794 (N_13794,N_13153,N_13145);
or U13795 (N_13795,N_13014,N_13359);
or U13796 (N_13796,N_13316,N_13113);
and U13797 (N_13797,N_12918,N_13037);
nand U13798 (N_13798,N_12752,N_13006);
or U13799 (N_13799,N_13093,N_13368);
and U13800 (N_13800,N_12936,N_12942);
and U13801 (N_13801,N_13250,N_13416);
nor U13802 (N_13802,N_13302,N_13437);
nand U13803 (N_13803,N_13137,N_13342);
nand U13804 (N_13804,N_13089,N_13241);
or U13805 (N_13805,N_13298,N_13329);
nor U13806 (N_13806,N_13060,N_13027);
and U13807 (N_13807,N_13267,N_13303);
nor U13808 (N_13808,N_12883,N_12963);
or U13809 (N_13809,N_13396,N_12890);
nor U13810 (N_13810,N_13248,N_13254);
or U13811 (N_13811,N_13441,N_13300);
xnor U13812 (N_13812,N_13436,N_13157);
and U13813 (N_13813,N_12986,N_12999);
nor U13814 (N_13814,N_13390,N_13143);
and U13815 (N_13815,N_13195,N_13421);
xnor U13816 (N_13816,N_12825,N_12982);
nor U13817 (N_13817,N_13224,N_12750);
nor U13818 (N_13818,N_13218,N_13266);
nand U13819 (N_13819,N_12768,N_12907);
or U13820 (N_13820,N_12833,N_12908);
nand U13821 (N_13821,N_13150,N_13304);
or U13822 (N_13822,N_12862,N_12975);
nand U13823 (N_13823,N_13268,N_13399);
nor U13824 (N_13824,N_13461,N_13234);
and U13825 (N_13825,N_13186,N_13276);
nand U13826 (N_13826,N_12854,N_13404);
and U13827 (N_13827,N_13296,N_13431);
xor U13828 (N_13828,N_13341,N_12785);
nor U13829 (N_13829,N_13313,N_13050);
xnor U13830 (N_13830,N_13253,N_12967);
nor U13831 (N_13831,N_13324,N_13454);
and U13832 (N_13832,N_13068,N_13255);
xor U13833 (N_13833,N_13126,N_13388);
xor U13834 (N_13834,N_12997,N_12925);
nand U13835 (N_13835,N_13336,N_13327);
nand U13836 (N_13836,N_13261,N_13077);
nand U13837 (N_13837,N_13355,N_13385);
and U13838 (N_13838,N_13370,N_13281);
nand U13839 (N_13839,N_13299,N_13447);
xor U13840 (N_13840,N_13394,N_13147);
nand U13841 (N_13841,N_13448,N_13455);
nor U13842 (N_13842,N_13155,N_12790);
nor U13843 (N_13843,N_12797,N_13249);
nand U13844 (N_13844,N_12837,N_12911);
nor U13845 (N_13845,N_13270,N_13127);
and U13846 (N_13846,N_13343,N_12940);
xor U13847 (N_13847,N_12791,N_13265);
nor U13848 (N_13848,N_13222,N_12860);
nor U13849 (N_13849,N_13478,N_13100);
or U13850 (N_13850,N_12884,N_13175);
nand U13851 (N_13851,N_12937,N_13326);
and U13852 (N_13852,N_13141,N_13321);
xor U13853 (N_13853,N_13415,N_13007);
nor U13854 (N_13854,N_13418,N_12843);
nor U13855 (N_13855,N_12930,N_13362);
or U13856 (N_13856,N_13152,N_12958);
or U13857 (N_13857,N_13332,N_12782);
nor U13858 (N_13858,N_13492,N_13494);
nand U13859 (N_13859,N_13442,N_12923);
and U13860 (N_13860,N_12869,N_13056);
or U13861 (N_13861,N_12905,N_12809);
and U13862 (N_13862,N_13161,N_13297);
or U13863 (N_13863,N_13202,N_13236);
and U13864 (N_13864,N_13238,N_12859);
or U13865 (N_13865,N_13025,N_13221);
nor U13866 (N_13866,N_13422,N_13120);
nand U13867 (N_13867,N_12819,N_12878);
nand U13868 (N_13868,N_12841,N_12865);
xor U13869 (N_13869,N_13041,N_13034);
and U13870 (N_13870,N_13111,N_13259);
nand U13871 (N_13871,N_13139,N_12922);
nand U13872 (N_13872,N_13444,N_13174);
nor U13873 (N_13873,N_13160,N_13199);
nor U13874 (N_13874,N_13106,N_12846);
or U13875 (N_13875,N_13279,N_13228);
nor U13876 (N_13876,N_13123,N_13214);
or U13877 (N_13877,N_13089,N_13178);
nor U13878 (N_13878,N_12901,N_13332);
nand U13879 (N_13879,N_13100,N_13367);
or U13880 (N_13880,N_13024,N_12979);
xnor U13881 (N_13881,N_12795,N_12834);
or U13882 (N_13882,N_12941,N_13370);
and U13883 (N_13883,N_13158,N_12842);
nor U13884 (N_13884,N_13094,N_12870);
or U13885 (N_13885,N_12949,N_12939);
nand U13886 (N_13886,N_13407,N_13452);
nand U13887 (N_13887,N_12911,N_13323);
and U13888 (N_13888,N_13129,N_13348);
xnor U13889 (N_13889,N_13058,N_13416);
xor U13890 (N_13890,N_13168,N_13354);
xnor U13891 (N_13891,N_13233,N_13471);
nand U13892 (N_13892,N_13099,N_13153);
or U13893 (N_13893,N_13069,N_12827);
nor U13894 (N_13894,N_13493,N_12838);
nand U13895 (N_13895,N_13423,N_12983);
nor U13896 (N_13896,N_12936,N_13426);
nand U13897 (N_13897,N_12947,N_13411);
nor U13898 (N_13898,N_13400,N_12876);
nor U13899 (N_13899,N_13353,N_13025);
and U13900 (N_13900,N_13499,N_12860);
and U13901 (N_13901,N_12777,N_13244);
or U13902 (N_13902,N_13422,N_13365);
or U13903 (N_13903,N_13452,N_13256);
nor U13904 (N_13904,N_13059,N_12826);
or U13905 (N_13905,N_12844,N_13127);
nor U13906 (N_13906,N_13066,N_13198);
nand U13907 (N_13907,N_13429,N_13284);
xor U13908 (N_13908,N_12941,N_13195);
nand U13909 (N_13909,N_13327,N_12941);
or U13910 (N_13910,N_13363,N_12788);
or U13911 (N_13911,N_13227,N_12962);
or U13912 (N_13912,N_13265,N_13322);
or U13913 (N_13913,N_13195,N_13137);
nor U13914 (N_13914,N_13108,N_13030);
nand U13915 (N_13915,N_13165,N_12970);
and U13916 (N_13916,N_12821,N_13125);
or U13917 (N_13917,N_12853,N_13010);
and U13918 (N_13918,N_12982,N_12850);
nor U13919 (N_13919,N_13062,N_13099);
and U13920 (N_13920,N_13226,N_12883);
nand U13921 (N_13921,N_13249,N_13088);
nor U13922 (N_13922,N_12874,N_12818);
nor U13923 (N_13923,N_13211,N_12802);
or U13924 (N_13924,N_12789,N_12837);
xnor U13925 (N_13925,N_13224,N_13236);
or U13926 (N_13926,N_12907,N_12759);
nor U13927 (N_13927,N_13325,N_13227);
and U13928 (N_13928,N_13123,N_13454);
and U13929 (N_13929,N_13019,N_13490);
and U13930 (N_13930,N_13189,N_13172);
xor U13931 (N_13931,N_12951,N_13339);
or U13932 (N_13932,N_13003,N_13333);
nand U13933 (N_13933,N_13357,N_12876);
nand U13934 (N_13934,N_12969,N_13155);
or U13935 (N_13935,N_12783,N_12964);
nor U13936 (N_13936,N_13401,N_13339);
nand U13937 (N_13937,N_13407,N_12843);
or U13938 (N_13938,N_13290,N_12961);
and U13939 (N_13939,N_13202,N_13406);
nand U13940 (N_13940,N_13016,N_12943);
nand U13941 (N_13941,N_13250,N_13035);
or U13942 (N_13942,N_13026,N_13461);
or U13943 (N_13943,N_13050,N_13014);
nand U13944 (N_13944,N_13226,N_13255);
or U13945 (N_13945,N_13061,N_13084);
and U13946 (N_13946,N_13450,N_13473);
nor U13947 (N_13947,N_12965,N_13335);
or U13948 (N_13948,N_13084,N_13131);
nor U13949 (N_13949,N_12789,N_13026);
or U13950 (N_13950,N_13493,N_12903);
or U13951 (N_13951,N_12949,N_13026);
or U13952 (N_13952,N_13167,N_13035);
nand U13953 (N_13953,N_13466,N_12795);
nor U13954 (N_13954,N_13066,N_13456);
xor U13955 (N_13955,N_13049,N_13254);
nand U13956 (N_13956,N_12954,N_13303);
nor U13957 (N_13957,N_13292,N_13359);
nand U13958 (N_13958,N_13007,N_12868);
nand U13959 (N_13959,N_12772,N_13217);
nor U13960 (N_13960,N_13219,N_13222);
nor U13961 (N_13961,N_13447,N_13154);
or U13962 (N_13962,N_12816,N_13117);
xor U13963 (N_13963,N_13404,N_13006);
nor U13964 (N_13964,N_12815,N_12977);
and U13965 (N_13965,N_12837,N_13210);
xor U13966 (N_13966,N_12778,N_12809);
and U13967 (N_13967,N_13359,N_13160);
or U13968 (N_13968,N_12765,N_12867);
nand U13969 (N_13969,N_13436,N_12854);
and U13970 (N_13970,N_13334,N_13391);
nor U13971 (N_13971,N_13183,N_12893);
or U13972 (N_13972,N_13471,N_13262);
xnor U13973 (N_13973,N_13223,N_13066);
and U13974 (N_13974,N_13036,N_13212);
nand U13975 (N_13975,N_13043,N_12938);
xnor U13976 (N_13976,N_12762,N_12760);
nand U13977 (N_13977,N_13278,N_13166);
and U13978 (N_13978,N_13011,N_12865);
xnor U13979 (N_13979,N_13210,N_13284);
nor U13980 (N_13980,N_13241,N_12844);
and U13981 (N_13981,N_13118,N_13479);
nor U13982 (N_13982,N_13419,N_13418);
or U13983 (N_13983,N_13090,N_13376);
nand U13984 (N_13984,N_13186,N_12839);
and U13985 (N_13985,N_12973,N_12923);
nor U13986 (N_13986,N_13489,N_12830);
xnor U13987 (N_13987,N_12806,N_13246);
nor U13988 (N_13988,N_13428,N_12947);
or U13989 (N_13989,N_13215,N_12794);
or U13990 (N_13990,N_13154,N_12868);
nand U13991 (N_13991,N_13454,N_12793);
or U13992 (N_13992,N_13277,N_13422);
or U13993 (N_13993,N_13261,N_13296);
and U13994 (N_13994,N_12908,N_13454);
and U13995 (N_13995,N_13191,N_12842);
and U13996 (N_13996,N_13104,N_12895);
and U13997 (N_13997,N_12858,N_13187);
nand U13998 (N_13998,N_13409,N_12801);
and U13999 (N_13999,N_13088,N_13312);
nor U14000 (N_14000,N_13483,N_13458);
nor U14001 (N_14001,N_13452,N_12801);
nand U14002 (N_14002,N_12900,N_13420);
nor U14003 (N_14003,N_12791,N_13065);
xor U14004 (N_14004,N_13164,N_12866);
nor U14005 (N_14005,N_13217,N_13067);
and U14006 (N_14006,N_13079,N_13445);
or U14007 (N_14007,N_13459,N_13462);
or U14008 (N_14008,N_12965,N_13115);
xor U14009 (N_14009,N_13087,N_13038);
nor U14010 (N_14010,N_13253,N_13269);
nor U14011 (N_14011,N_13268,N_13001);
nor U14012 (N_14012,N_13204,N_13206);
xor U14013 (N_14013,N_13065,N_12928);
and U14014 (N_14014,N_13297,N_13270);
nor U14015 (N_14015,N_13383,N_12957);
or U14016 (N_14016,N_13225,N_13069);
or U14017 (N_14017,N_12853,N_12792);
nand U14018 (N_14018,N_13146,N_13088);
nor U14019 (N_14019,N_12819,N_13446);
nor U14020 (N_14020,N_13480,N_13280);
nand U14021 (N_14021,N_12860,N_12870);
nand U14022 (N_14022,N_13180,N_13226);
and U14023 (N_14023,N_13019,N_12861);
nor U14024 (N_14024,N_13328,N_12980);
nor U14025 (N_14025,N_12915,N_12979);
or U14026 (N_14026,N_12922,N_13370);
or U14027 (N_14027,N_13471,N_12804);
or U14028 (N_14028,N_13301,N_12853);
or U14029 (N_14029,N_12919,N_13015);
and U14030 (N_14030,N_13462,N_13093);
or U14031 (N_14031,N_13010,N_13299);
or U14032 (N_14032,N_12819,N_13352);
xnor U14033 (N_14033,N_12808,N_13481);
or U14034 (N_14034,N_13224,N_13444);
nand U14035 (N_14035,N_13205,N_13364);
nand U14036 (N_14036,N_12824,N_12884);
nand U14037 (N_14037,N_13098,N_13073);
nand U14038 (N_14038,N_12974,N_13493);
nor U14039 (N_14039,N_12875,N_13095);
nand U14040 (N_14040,N_13028,N_13478);
and U14041 (N_14041,N_13467,N_12842);
and U14042 (N_14042,N_12986,N_13474);
and U14043 (N_14043,N_13088,N_13150);
xnor U14044 (N_14044,N_12935,N_13033);
nand U14045 (N_14045,N_12842,N_13249);
or U14046 (N_14046,N_13359,N_13123);
and U14047 (N_14047,N_13029,N_13151);
xnor U14048 (N_14048,N_12972,N_13207);
or U14049 (N_14049,N_13390,N_12970);
and U14050 (N_14050,N_13268,N_13045);
nor U14051 (N_14051,N_13104,N_12810);
nand U14052 (N_14052,N_12810,N_12836);
or U14053 (N_14053,N_13050,N_13258);
xor U14054 (N_14054,N_13209,N_12985);
nand U14055 (N_14055,N_13012,N_13068);
or U14056 (N_14056,N_13320,N_12783);
nand U14057 (N_14057,N_13333,N_13269);
nand U14058 (N_14058,N_13085,N_12815);
nand U14059 (N_14059,N_13337,N_12987);
nor U14060 (N_14060,N_12925,N_13245);
nand U14061 (N_14061,N_13199,N_13440);
nand U14062 (N_14062,N_13455,N_13212);
nor U14063 (N_14063,N_12864,N_13472);
nor U14064 (N_14064,N_12867,N_12807);
and U14065 (N_14065,N_13402,N_12993);
and U14066 (N_14066,N_13282,N_12867);
xnor U14067 (N_14067,N_13369,N_12816);
and U14068 (N_14068,N_13205,N_13478);
or U14069 (N_14069,N_13039,N_13173);
nand U14070 (N_14070,N_13134,N_13266);
xnor U14071 (N_14071,N_12971,N_13053);
nor U14072 (N_14072,N_13359,N_13055);
or U14073 (N_14073,N_13002,N_13231);
and U14074 (N_14074,N_12887,N_13030);
nor U14075 (N_14075,N_13402,N_12752);
or U14076 (N_14076,N_13061,N_12793);
nand U14077 (N_14077,N_12861,N_13288);
nand U14078 (N_14078,N_13271,N_13270);
and U14079 (N_14079,N_13389,N_13347);
and U14080 (N_14080,N_13020,N_12912);
nand U14081 (N_14081,N_13329,N_12964);
xor U14082 (N_14082,N_13439,N_13428);
and U14083 (N_14083,N_13362,N_13496);
and U14084 (N_14084,N_13202,N_13232);
or U14085 (N_14085,N_12754,N_13384);
or U14086 (N_14086,N_12786,N_13293);
nand U14087 (N_14087,N_13267,N_12873);
nand U14088 (N_14088,N_12983,N_13078);
and U14089 (N_14089,N_13484,N_13212);
nand U14090 (N_14090,N_13029,N_12888);
nor U14091 (N_14091,N_12860,N_12808);
and U14092 (N_14092,N_13489,N_12885);
nand U14093 (N_14093,N_12983,N_12986);
nand U14094 (N_14094,N_12866,N_12856);
or U14095 (N_14095,N_13153,N_13108);
nor U14096 (N_14096,N_13422,N_12832);
nand U14097 (N_14097,N_12894,N_13038);
nor U14098 (N_14098,N_13230,N_13058);
nand U14099 (N_14099,N_13034,N_13491);
and U14100 (N_14100,N_13123,N_13162);
or U14101 (N_14101,N_13434,N_12980);
nand U14102 (N_14102,N_13285,N_13412);
nand U14103 (N_14103,N_13359,N_13234);
nor U14104 (N_14104,N_13189,N_13199);
and U14105 (N_14105,N_12788,N_12981);
nand U14106 (N_14106,N_13045,N_12781);
xnor U14107 (N_14107,N_13390,N_13212);
xnor U14108 (N_14108,N_13181,N_12791);
nor U14109 (N_14109,N_13053,N_12852);
nor U14110 (N_14110,N_12822,N_12988);
nand U14111 (N_14111,N_13261,N_13389);
xnor U14112 (N_14112,N_12992,N_12896);
or U14113 (N_14113,N_12807,N_13152);
and U14114 (N_14114,N_13315,N_12842);
nand U14115 (N_14115,N_13401,N_13154);
or U14116 (N_14116,N_13129,N_13175);
xnor U14117 (N_14117,N_12986,N_12853);
or U14118 (N_14118,N_12996,N_13033);
or U14119 (N_14119,N_13301,N_12778);
and U14120 (N_14120,N_12762,N_12906);
nand U14121 (N_14121,N_13228,N_13225);
xor U14122 (N_14122,N_12949,N_12776);
xnor U14123 (N_14123,N_12925,N_13233);
xor U14124 (N_14124,N_12753,N_12950);
and U14125 (N_14125,N_13235,N_13413);
or U14126 (N_14126,N_12752,N_13280);
and U14127 (N_14127,N_13422,N_13010);
nand U14128 (N_14128,N_13148,N_12955);
xnor U14129 (N_14129,N_12962,N_12861);
and U14130 (N_14130,N_12856,N_12975);
nor U14131 (N_14131,N_13123,N_12952);
and U14132 (N_14132,N_13051,N_13129);
or U14133 (N_14133,N_13432,N_13027);
and U14134 (N_14134,N_13132,N_12858);
or U14135 (N_14135,N_12974,N_12816);
and U14136 (N_14136,N_13151,N_12816);
and U14137 (N_14137,N_13374,N_13231);
and U14138 (N_14138,N_12785,N_12880);
nand U14139 (N_14139,N_13323,N_13406);
nor U14140 (N_14140,N_13445,N_13308);
xnor U14141 (N_14141,N_13298,N_12983);
nor U14142 (N_14142,N_13157,N_12752);
nand U14143 (N_14143,N_13011,N_13380);
or U14144 (N_14144,N_13057,N_13238);
xor U14145 (N_14145,N_12843,N_12854);
and U14146 (N_14146,N_12973,N_13118);
nor U14147 (N_14147,N_13026,N_13406);
xnor U14148 (N_14148,N_13470,N_13257);
nand U14149 (N_14149,N_13063,N_13026);
nand U14150 (N_14150,N_12861,N_13341);
nor U14151 (N_14151,N_12872,N_13366);
and U14152 (N_14152,N_13294,N_13107);
nor U14153 (N_14153,N_13155,N_12986);
nor U14154 (N_14154,N_13108,N_13439);
and U14155 (N_14155,N_13174,N_13165);
nor U14156 (N_14156,N_13374,N_12981);
xnor U14157 (N_14157,N_13089,N_13167);
and U14158 (N_14158,N_13084,N_13350);
nand U14159 (N_14159,N_13382,N_13315);
and U14160 (N_14160,N_12985,N_13446);
nor U14161 (N_14161,N_12750,N_13091);
nor U14162 (N_14162,N_13351,N_13364);
or U14163 (N_14163,N_13456,N_13345);
xor U14164 (N_14164,N_12999,N_12984);
and U14165 (N_14165,N_13024,N_12765);
nand U14166 (N_14166,N_13316,N_12840);
nor U14167 (N_14167,N_13451,N_13299);
and U14168 (N_14168,N_13461,N_13253);
or U14169 (N_14169,N_13039,N_12896);
nor U14170 (N_14170,N_13426,N_12946);
and U14171 (N_14171,N_13082,N_13126);
and U14172 (N_14172,N_12785,N_12928);
nand U14173 (N_14173,N_13013,N_13076);
and U14174 (N_14174,N_12917,N_12895);
or U14175 (N_14175,N_13173,N_13032);
and U14176 (N_14176,N_13030,N_13156);
xor U14177 (N_14177,N_13451,N_12785);
nand U14178 (N_14178,N_13147,N_12814);
and U14179 (N_14179,N_13254,N_12905);
or U14180 (N_14180,N_12939,N_13336);
nor U14181 (N_14181,N_13033,N_13169);
xnor U14182 (N_14182,N_12750,N_13423);
or U14183 (N_14183,N_12854,N_12752);
nor U14184 (N_14184,N_13334,N_13119);
nand U14185 (N_14185,N_13257,N_13347);
nand U14186 (N_14186,N_13462,N_12943);
nor U14187 (N_14187,N_13146,N_13127);
nor U14188 (N_14188,N_12949,N_13128);
and U14189 (N_14189,N_12815,N_13161);
xnor U14190 (N_14190,N_12888,N_13264);
or U14191 (N_14191,N_12979,N_13221);
xor U14192 (N_14192,N_12990,N_12861);
xnor U14193 (N_14193,N_13450,N_13188);
nand U14194 (N_14194,N_12862,N_13226);
or U14195 (N_14195,N_12981,N_13047);
or U14196 (N_14196,N_13284,N_13287);
nor U14197 (N_14197,N_13312,N_12993);
xnor U14198 (N_14198,N_13142,N_12761);
nor U14199 (N_14199,N_13037,N_13492);
or U14200 (N_14200,N_13380,N_13172);
nand U14201 (N_14201,N_12966,N_13038);
and U14202 (N_14202,N_13044,N_13456);
nor U14203 (N_14203,N_13007,N_13324);
nor U14204 (N_14204,N_12807,N_13359);
nor U14205 (N_14205,N_13255,N_13044);
nand U14206 (N_14206,N_13048,N_12857);
nand U14207 (N_14207,N_13184,N_13435);
or U14208 (N_14208,N_13079,N_12788);
or U14209 (N_14209,N_13325,N_13171);
nand U14210 (N_14210,N_13329,N_13383);
and U14211 (N_14211,N_13476,N_13146);
or U14212 (N_14212,N_13402,N_12794);
nand U14213 (N_14213,N_13006,N_13480);
nand U14214 (N_14214,N_12991,N_12967);
and U14215 (N_14215,N_12990,N_13266);
and U14216 (N_14216,N_13054,N_13097);
or U14217 (N_14217,N_13168,N_13131);
nor U14218 (N_14218,N_12962,N_13054);
nor U14219 (N_14219,N_12750,N_13158);
nand U14220 (N_14220,N_13304,N_13463);
and U14221 (N_14221,N_13270,N_13283);
or U14222 (N_14222,N_13405,N_13380);
or U14223 (N_14223,N_12968,N_13399);
nand U14224 (N_14224,N_12853,N_13429);
nand U14225 (N_14225,N_12808,N_12997);
nor U14226 (N_14226,N_12874,N_13002);
or U14227 (N_14227,N_12916,N_12876);
nand U14228 (N_14228,N_12823,N_12857);
and U14229 (N_14229,N_13333,N_13347);
nor U14230 (N_14230,N_13206,N_13017);
and U14231 (N_14231,N_13081,N_13393);
nor U14232 (N_14232,N_13006,N_13011);
nand U14233 (N_14233,N_12872,N_12871);
nor U14234 (N_14234,N_13456,N_13198);
and U14235 (N_14235,N_13021,N_12907);
nand U14236 (N_14236,N_13455,N_12769);
and U14237 (N_14237,N_13104,N_13338);
and U14238 (N_14238,N_13247,N_13273);
nand U14239 (N_14239,N_13041,N_13318);
nand U14240 (N_14240,N_13470,N_13398);
or U14241 (N_14241,N_12797,N_13210);
nand U14242 (N_14242,N_13008,N_13037);
and U14243 (N_14243,N_13366,N_13084);
and U14244 (N_14244,N_13086,N_12776);
nand U14245 (N_14245,N_13034,N_12824);
nor U14246 (N_14246,N_12869,N_13459);
nor U14247 (N_14247,N_13480,N_12769);
or U14248 (N_14248,N_12816,N_13354);
nor U14249 (N_14249,N_12942,N_13089);
nand U14250 (N_14250,N_13764,N_13616);
nor U14251 (N_14251,N_13856,N_13703);
nand U14252 (N_14252,N_14177,N_13805);
nand U14253 (N_14253,N_14088,N_13599);
or U14254 (N_14254,N_13697,N_13605);
or U14255 (N_14255,N_13962,N_14092);
xor U14256 (N_14256,N_13571,N_13732);
nor U14257 (N_14257,N_14182,N_14209);
nor U14258 (N_14258,N_14062,N_14167);
nand U14259 (N_14259,N_14006,N_14166);
or U14260 (N_14260,N_13928,N_13502);
xor U14261 (N_14261,N_13950,N_14127);
nand U14262 (N_14262,N_13522,N_14172);
or U14263 (N_14263,N_13613,N_13749);
nand U14264 (N_14264,N_13747,N_14032);
and U14265 (N_14265,N_13627,N_13861);
or U14266 (N_14266,N_13505,N_13809);
or U14267 (N_14267,N_14099,N_13614);
and U14268 (N_14268,N_14005,N_13816);
and U14269 (N_14269,N_13951,N_14004);
nor U14270 (N_14270,N_13968,N_13778);
nand U14271 (N_14271,N_14044,N_14247);
nor U14272 (N_14272,N_14249,N_13733);
xor U14273 (N_14273,N_14084,N_13563);
xor U14274 (N_14274,N_13716,N_13972);
nor U14275 (N_14275,N_13854,N_13783);
nand U14276 (N_14276,N_13507,N_13606);
and U14277 (N_14277,N_14055,N_13985);
nor U14278 (N_14278,N_13860,N_13779);
xor U14279 (N_14279,N_13823,N_14094);
or U14280 (N_14280,N_13902,N_13996);
nand U14281 (N_14281,N_13685,N_13899);
and U14282 (N_14282,N_14134,N_14157);
and U14283 (N_14283,N_14174,N_13953);
or U14284 (N_14284,N_14022,N_13843);
nand U14285 (N_14285,N_13837,N_13546);
nor U14286 (N_14286,N_13648,N_14171);
and U14287 (N_14287,N_13738,N_13819);
nand U14288 (N_14288,N_13775,N_13548);
or U14289 (N_14289,N_13875,N_13610);
or U14290 (N_14290,N_13913,N_13562);
and U14291 (N_14291,N_14136,N_13882);
nand U14292 (N_14292,N_13666,N_14061);
and U14293 (N_14293,N_13541,N_13516);
or U14294 (N_14294,N_14190,N_14191);
nand U14295 (N_14295,N_13900,N_13797);
nand U14296 (N_14296,N_14128,N_13592);
xor U14297 (N_14297,N_13609,N_14040);
nor U14298 (N_14298,N_13859,N_13957);
and U14299 (N_14299,N_13920,N_14104);
nor U14300 (N_14300,N_13657,N_14160);
xnor U14301 (N_14301,N_14186,N_14053);
nor U14302 (N_14302,N_13695,N_13838);
nand U14303 (N_14303,N_14144,N_14067);
nor U14304 (N_14304,N_14119,N_13892);
and U14305 (N_14305,N_13814,N_13568);
or U14306 (N_14306,N_13932,N_13940);
nand U14307 (N_14307,N_14096,N_13708);
nand U14308 (N_14308,N_14118,N_13907);
or U14309 (N_14309,N_13851,N_13628);
and U14310 (N_14310,N_13714,N_13773);
nor U14311 (N_14311,N_13622,N_13650);
nor U14312 (N_14312,N_13725,N_14154);
or U14313 (N_14313,N_14090,N_13894);
nand U14314 (N_14314,N_13791,N_14152);
or U14315 (N_14315,N_13575,N_13529);
nand U14316 (N_14316,N_14196,N_13739);
and U14317 (N_14317,N_13943,N_13848);
or U14318 (N_14318,N_13784,N_13586);
xnor U14319 (N_14319,N_13679,N_13883);
or U14320 (N_14320,N_13681,N_14208);
nor U14321 (N_14321,N_13981,N_14176);
and U14322 (N_14322,N_14031,N_14195);
nand U14323 (N_14323,N_13889,N_13821);
xnor U14324 (N_14324,N_14140,N_13873);
or U14325 (N_14325,N_14236,N_13591);
or U14326 (N_14326,N_13514,N_14016);
nor U14327 (N_14327,N_13533,N_14203);
and U14328 (N_14328,N_14057,N_13579);
nor U14329 (N_14329,N_14226,N_13970);
nand U14330 (N_14330,N_14027,N_13506);
or U14331 (N_14331,N_14000,N_14223);
or U14332 (N_14332,N_13585,N_13871);
and U14333 (N_14333,N_13788,N_13817);
nand U14334 (N_14334,N_13658,N_13511);
or U14335 (N_14335,N_13551,N_14052);
or U14336 (N_14336,N_13676,N_14151);
nor U14337 (N_14337,N_14019,N_13518);
nand U14338 (N_14338,N_13647,N_13671);
and U14339 (N_14339,N_13574,N_13852);
or U14340 (N_14340,N_14085,N_13904);
xor U14341 (N_14341,N_13526,N_13901);
or U14342 (N_14342,N_14246,N_13550);
nor U14343 (N_14343,N_13826,N_13745);
and U14344 (N_14344,N_13915,N_14066);
nor U14345 (N_14345,N_14218,N_14248);
nor U14346 (N_14346,N_13531,N_13870);
nand U14347 (N_14347,N_14064,N_13594);
nor U14348 (N_14348,N_13630,N_13960);
nor U14349 (N_14349,N_13520,N_14153);
or U14350 (N_14350,N_13555,N_13799);
or U14351 (N_14351,N_13712,N_14173);
and U14352 (N_14352,N_13631,N_13564);
or U14353 (N_14353,N_13737,N_13759);
nor U14354 (N_14354,N_13536,N_13969);
nand U14355 (N_14355,N_13834,N_13669);
nor U14356 (N_14356,N_14130,N_13527);
or U14357 (N_14357,N_13946,N_13636);
nand U14358 (N_14358,N_13980,N_13727);
nand U14359 (N_14359,N_14146,N_14237);
and U14360 (N_14360,N_13984,N_14077);
nand U14361 (N_14361,N_13992,N_13961);
nor U14362 (N_14362,N_13715,N_14222);
xnor U14363 (N_14363,N_13722,N_14220);
and U14364 (N_14364,N_13942,N_13982);
nand U14365 (N_14365,N_13668,N_13919);
or U14366 (N_14366,N_13977,N_13608);
or U14367 (N_14367,N_13909,N_13718);
and U14368 (N_14368,N_13758,N_13849);
xnor U14369 (N_14369,N_13547,N_14145);
nor U14370 (N_14370,N_14107,N_13659);
xnor U14371 (N_14371,N_14206,N_13785);
nor U14372 (N_14372,N_13895,N_13975);
or U14373 (N_14373,N_14198,N_14038);
nand U14374 (N_14374,N_13830,N_14101);
nor U14375 (N_14375,N_13807,N_13686);
nand U14376 (N_14376,N_13787,N_13641);
or U14377 (N_14377,N_13615,N_13986);
nor U14378 (N_14378,N_13661,N_13696);
nor U14379 (N_14379,N_13515,N_13963);
nand U14380 (N_14380,N_13735,N_13811);
and U14381 (N_14381,N_14193,N_14149);
nor U14382 (N_14382,N_13633,N_13927);
or U14383 (N_14383,N_14227,N_14108);
xor U14384 (N_14384,N_14213,N_13995);
nand U14385 (N_14385,N_14180,N_13748);
or U14386 (N_14386,N_14011,N_13971);
nand U14387 (N_14387,N_14243,N_14042);
nor U14388 (N_14388,N_13717,N_13517);
nand U14389 (N_14389,N_13559,N_13523);
nand U14390 (N_14390,N_13790,N_14013);
and U14391 (N_14391,N_14158,N_14161);
and U14392 (N_14392,N_14217,N_13705);
and U14393 (N_14393,N_13897,N_13554);
xnor U14394 (N_14394,N_13924,N_13908);
or U14395 (N_14395,N_14111,N_13921);
or U14396 (N_14396,N_14034,N_13690);
or U14397 (N_14397,N_13941,N_14008);
nor U14398 (N_14398,N_13626,N_14138);
and U14399 (N_14399,N_14215,N_13584);
xor U14400 (N_14400,N_14165,N_13635);
and U14401 (N_14401,N_14137,N_13624);
nor U14402 (N_14402,N_13637,N_13910);
and U14403 (N_14403,N_13741,N_13623);
or U14404 (N_14404,N_13815,N_13937);
nand U14405 (N_14405,N_13929,N_13567);
and U14406 (N_14406,N_13964,N_14116);
and U14407 (N_14407,N_14155,N_13565);
nor U14408 (N_14408,N_13954,N_14037);
and U14409 (N_14409,N_13651,N_13966);
or U14410 (N_14410,N_14010,N_13699);
or U14411 (N_14411,N_14143,N_13692);
and U14412 (N_14412,N_14081,N_14169);
nand U14413 (N_14413,N_14188,N_14002);
and U14414 (N_14414,N_14095,N_13713);
nor U14415 (N_14415,N_13639,N_13812);
nor U14416 (N_14416,N_14235,N_13833);
nor U14417 (N_14417,N_13743,N_14029);
and U14418 (N_14418,N_14048,N_14162);
or U14419 (N_14419,N_13744,N_14139);
and U14420 (N_14420,N_14023,N_13872);
or U14421 (N_14421,N_13578,N_13582);
xor U14422 (N_14422,N_13867,N_14230);
or U14423 (N_14423,N_14201,N_13543);
xnor U14424 (N_14424,N_13683,N_14123);
nor U14425 (N_14425,N_13978,N_13997);
nor U14426 (N_14426,N_14212,N_13832);
and U14427 (N_14427,N_13795,N_13673);
nand U14428 (N_14428,N_14046,N_13857);
nand U14429 (N_14429,N_13884,N_13781);
or U14430 (N_14430,N_14133,N_13914);
or U14431 (N_14431,N_13602,N_14241);
nand U14432 (N_14432,N_13770,N_13876);
nor U14433 (N_14433,N_13680,N_14098);
nand U14434 (N_14434,N_13534,N_13903);
nor U14435 (N_14435,N_13598,N_13912);
and U14436 (N_14436,N_13740,N_14229);
and U14437 (N_14437,N_14073,N_13700);
nor U14438 (N_14438,N_14021,N_14141);
xor U14439 (N_14439,N_14028,N_13508);
or U14440 (N_14440,N_13948,N_13800);
nand U14441 (N_14441,N_14184,N_13645);
nand U14442 (N_14442,N_13558,N_14074);
nand U14443 (N_14443,N_14009,N_13698);
nand U14444 (N_14444,N_13825,N_13829);
or U14445 (N_14445,N_13603,N_13893);
nand U14446 (N_14446,N_13612,N_13933);
nor U14447 (N_14447,N_13906,N_13569);
nand U14448 (N_14448,N_13760,N_13793);
and U14449 (N_14449,N_14087,N_13822);
nand U14450 (N_14450,N_13640,N_13880);
nor U14451 (N_14451,N_14200,N_13881);
nor U14452 (N_14452,N_13755,N_13600);
and U14453 (N_14453,N_13728,N_13662);
nor U14454 (N_14454,N_13580,N_13656);
nand U14455 (N_14455,N_14102,N_13844);
nor U14456 (N_14456,N_14175,N_13930);
xor U14457 (N_14457,N_13947,N_13827);
nor U14458 (N_14458,N_14179,N_13644);
or U14459 (N_14459,N_13798,N_14211);
or U14460 (N_14460,N_13752,N_13993);
or U14461 (N_14461,N_13983,N_14242);
nor U14462 (N_14462,N_13987,N_14071);
or U14463 (N_14463,N_14183,N_13878);
and U14464 (N_14464,N_13869,N_13570);
or U14465 (N_14465,N_14170,N_13596);
and U14466 (N_14466,N_13831,N_14202);
and U14467 (N_14467,N_14043,N_13707);
nor U14468 (N_14468,N_13917,N_13777);
xnor U14469 (N_14469,N_13842,N_14041);
or U14470 (N_14470,N_13839,N_14110);
nor U14471 (N_14471,N_13864,N_13802);
or U14472 (N_14472,N_13723,N_13905);
or U14473 (N_14473,N_13820,N_14219);
nor U14474 (N_14474,N_13532,N_13916);
or U14475 (N_14475,N_13588,N_14097);
nor U14476 (N_14476,N_14142,N_13835);
nor U14477 (N_14477,N_14132,N_13655);
nor U14478 (N_14478,N_13664,N_14181);
or U14479 (N_14479,N_13742,N_13756);
nor U14480 (N_14480,N_14221,N_14070);
xor U14481 (N_14481,N_13806,N_13958);
nor U14482 (N_14482,N_14225,N_13840);
or U14483 (N_14483,N_13521,N_14185);
nand U14484 (N_14484,N_13545,N_14076);
nor U14485 (N_14485,N_13763,N_13704);
nand U14486 (N_14486,N_14207,N_13710);
nand U14487 (N_14487,N_14228,N_13866);
or U14488 (N_14488,N_14080,N_14159);
nand U14489 (N_14489,N_14007,N_13935);
xnor U14490 (N_14490,N_13939,N_14148);
or U14491 (N_14491,N_13544,N_14131);
nand U14492 (N_14492,N_14168,N_13949);
and U14493 (N_14493,N_13967,N_14147);
nor U14494 (N_14494,N_13769,N_14089);
or U14495 (N_14495,N_13934,N_13796);
nand U14496 (N_14496,N_13672,N_13674);
nor U14497 (N_14497,N_13855,N_13670);
nand U14498 (N_14498,N_13865,N_14065);
nor U14499 (N_14499,N_14189,N_13885);
and U14500 (N_14500,N_14072,N_13891);
or U14501 (N_14501,N_13896,N_13772);
and U14502 (N_14502,N_14012,N_13730);
and U14503 (N_14503,N_13682,N_14122);
nand U14504 (N_14504,N_14121,N_13989);
nor U14505 (N_14505,N_14187,N_14239);
nand U14506 (N_14506,N_13539,N_13619);
xor U14507 (N_14507,N_13538,N_14079);
nand U14508 (N_14508,N_13593,N_13525);
or U14509 (N_14509,N_13553,N_13751);
nand U14510 (N_14510,N_14086,N_13999);
xor U14511 (N_14511,N_13874,N_13719);
xor U14512 (N_14512,N_14017,N_13945);
nor U14513 (N_14513,N_13706,N_13753);
nand U14514 (N_14514,N_14135,N_13590);
nand U14515 (N_14515,N_14103,N_13618);
and U14516 (N_14516,N_14069,N_13581);
xnor U14517 (N_14517,N_13702,N_14106);
or U14518 (N_14518,N_14238,N_13918);
and U14519 (N_14519,N_13786,N_13549);
nand U14520 (N_14520,N_14045,N_13938);
or U14521 (N_14521,N_13625,N_13503);
or U14522 (N_14522,N_13990,N_14205);
nand U14523 (N_14523,N_14125,N_13731);
and U14524 (N_14524,N_13530,N_14214);
xnor U14525 (N_14525,N_14063,N_14093);
nor U14526 (N_14526,N_13512,N_13801);
and U14527 (N_14527,N_14240,N_13774);
nand U14528 (N_14528,N_13956,N_13804);
nand U14529 (N_14529,N_14216,N_13890);
nor U14530 (N_14530,N_14015,N_13687);
or U14531 (N_14531,N_13762,N_13604);
and U14532 (N_14532,N_13922,N_13660);
nor U14533 (N_14533,N_13587,N_14025);
and U14534 (N_14534,N_13994,N_13955);
nand U14535 (N_14535,N_14036,N_14194);
or U14536 (N_14536,N_13677,N_13754);
nand U14537 (N_14537,N_13768,N_13643);
nor U14538 (N_14538,N_13576,N_13846);
or U14539 (N_14539,N_13684,N_13560);
nand U14540 (N_14540,N_13965,N_14068);
nand U14541 (N_14541,N_13528,N_13766);
and U14542 (N_14542,N_13726,N_13620);
xor U14543 (N_14543,N_14024,N_13836);
and U14544 (N_14544,N_13808,N_13621);
nand U14545 (N_14545,N_13776,N_13642);
or U14546 (N_14546,N_13926,N_14051);
xor U14547 (N_14547,N_13974,N_14115);
or U14548 (N_14548,N_13589,N_13654);
and U14549 (N_14549,N_13879,N_13944);
and U14550 (N_14550,N_13634,N_13583);
or U14551 (N_14551,N_13729,N_13689);
nor U14552 (N_14552,N_13794,N_13542);
nand U14553 (N_14553,N_14156,N_13675);
or U14554 (N_14554,N_13601,N_13888);
xor U14555 (N_14555,N_13510,N_13868);
nor U14556 (N_14556,N_14210,N_14124);
nand U14557 (N_14557,N_13813,N_13988);
nand U14558 (N_14558,N_13736,N_13810);
and U14559 (N_14559,N_13720,N_13652);
or U14560 (N_14560,N_13573,N_13782);
nor U14561 (N_14561,N_13519,N_14192);
or U14562 (N_14562,N_14234,N_14003);
nand U14563 (N_14563,N_13976,N_13845);
xnor U14564 (N_14564,N_14075,N_13818);
or U14565 (N_14565,N_13537,N_13617);
nand U14566 (N_14566,N_13595,N_13898);
or U14567 (N_14567,N_13663,N_13667);
nor U14568 (N_14568,N_13973,N_13646);
nor U14569 (N_14569,N_13936,N_13858);
nand U14570 (N_14570,N_14129,N_14244);
or U14571 (N_14571,N_13923,N_14058);
nor U14572 (N_14572,N_13509,N_13803);
or U14573 (N_14573,N_13931,N_14114);
nand U14574 (N_14574,N_14164,N_14078);
nor U14575 (N_14575,N_13991,N_14014);
and U14576 (N_14576,N_13691,N_14091);
nand U14577 (N_14577,N_13767,N_13862);
nand U14578 (N_14578,N_14233,N_13886);
or U14579 (N_14579,N_13500,N_14105);
xnor U14580 (N_14580,N_14163,N_13828);
or U14581 (N_14581,N_13952,N_13911);
nand U14582 (N_14582,N_13632,N_13979);
nor U14583 (N_14583,N_14035,N_13711);
nor U14584 (N_14584,N_14100,N_13877);
and U14585 (N_14585,N_13597,N_13561);
nor U14586 (N_14586,N_14026,N_14047);
or U14587 (N_14587,N_13556,N_14204);
and U14588 (N_14588,N_14231,N_14060);
and U14589 (N_14589,N_13998,N_13665);
or U14590 (N_14590,N_13765,N_14059);
nor U14591 (N_14591,N_14232,N_13535);
nor U14592 (N_14592,N_14120,N_14109);
and U14593 (N_14593,N_13552,N_13504);
nand U14594 (N_14594,N_14224,N_13853);
nand U14595 (N_14595,N_13925,N_13678);
nand U14596 (N_14596,N_14178,N_13724);
nor U14597 (N_14597,N_14113,N_13847);
or U14598 (N_14598,N_13709,N_13524);
or U14599 (N_14599,N_14199,N_13750);
nor U14600 (N_14600,N_13501,N_13701);
nor U14601 (N_14601,N_13824,N_14082);
nand U14602 (N_14602,N_13757,N_14150);
or U14603 (N_14603,N_14245,N_13629);
nor U14604 (N_14604,N_13721,N_13959);
or U14605 (N_14605,N_14112,N_14018);
xnor U14606 (N_14606,N_14050,N_14054);
and U14607 (N_14607,N_13771,N_13694);
or U14608 (N_14608,N_14126,N_13513);
xor U14609 (N_14609,N_13607,N_13863);
and U14610 (N_14610,N_13653,N_13557);
xnor U14611 (N_14611,N_13780,N_14056);
nor U14612 (N_14612,N_13789,N_13566);
nand U14613 (N_14613,N_13792,N_13761);
and U14614 (N_14614,N_13540,N_13611);
and U14615 (N_14615,N_13649,N_13887);
or U14616 (N_14616,N_14117,N_13850);
nand U14617 (N_14617,N_13577,N_13841);
and U14618 (N_14618,N_14039,N_14030);
or U14619 (N_14619,N_14020,N_13638);
nor U14620 (N_14620,N_13693,N_14083);
nor U14621 (N_14621,N_13734,N_13572);
xor U14622 (N_14622,N_14001,N_13746);
or U14623 (N_14623,N_13688,N_14049);
or U14624 (N_14624,N_14197,N_14033);
nand U14625 (N_14625,N_13841,N_14227);
and U14626 (N_14626,N_13785,N_14182);
nor U14627 (N_14627,N_13957,N_13536);
and U14628 (N_14628,N_14129,N_13583);
nor U14629 (N_14629,N_13912,N_14011);
nor U14630 (N_14630,N_13892,N_13823);
and U14631 (N_14631,N_13792,N_14129);
nand U14632 (N_14632,N_14226,N_13798);
and U14633 (N_14633,N_13889,N_13614);
and U14634 (N_14634,N_14159,N_13589);
and U14635 (N_14635,N_13725,N_13700);
or U14636 (N_14636,N_13976,N_14230);
and U14637 (N_14637,N_13750,N_13994);
xor U14638 (N_14638,N_13803,N_14004);
nor U14639 (N_14639,N_13608,N_13648);
xor U14640 (N_14640,N_14216,N_14105);
or U14641 (N_14641,N_13659,N_13929);
nand U14642 (N_14642,N_14128,N_14091);
nor U14643 (N_14643,N_13918,N_13652);
and U14644 (N_14644,N_13532,N_13737);
nand U14645 (N_14645,N_13964,N_13594);
and U14646 (N_14646,N_13907,N_13773);
and U14647 (N_14647,N_13605,N_13590);
nand U14648 (N_14648,N_13789,N_13888);
or U14649 (N_14649,N_13779,N_13824);
nand U14650 (N_14650,N_14234,N_14090);
or U14651 (N_14651,N_14054,N_13509);
or U14652 (N_14652,N_13638,N_13839);
nor U14653 (N_14653,N_13928,N_14018);
and U14654 (N_14654,N_13694,N_14089);
nor U14655 (N_14655,N_14178,N_13834);
nor U14656 (N_14656,N_14067,N_13524);
xor U14657 (N_14657,N_13820,N_13684);
nand U14658 (N_14658,N_13663,N_13693);
and U14659 (N_14659,N_14027,N_14142);
or U14660 (N_14660,N_14191,N_13797);
nand U14661 (N_14661,N_13984,N_14044);
or U14662 (N_14662,N_14017,N_13830);
xnor U14663 (N_14663,N_13866,N_13529);
nand U14664 (N_14664,N_14087,N_13978);
nor U14665 (N_14665,N_13840,N_13606);
nor U14666 (N_14666,N_13869,N_14217);
or U14667 (N_14667,N_13533,N_14222);
nand U14668 (N_14668,N_13991,N_13581);
or U14669 (N_14669,N_14158,N_13899);
and U14670 (N_14670,N_14199,N_14019);
nand U14671 (N_14671,N_13779,N_13919);
nand U14672 (N_14672,N_14219,N_13751);
or U14673 (N_14673,N_14149,N_13619);
and U14674 (N_14674,N_13768,N_13544);
nor U14675 (N_14675,N_14237,N_13658);
or U14676 (N_14676,N_14155,N_13640);
or U14677 (N_14677,N_13780,N_13670);
nand U14678 (N_14678,N_13655,N_13595);
nand U14679 (N_14679,N_13789,N_13820);
nand U14680 (N_14680,N_14014,N_13672);
or U14681 (N_14681,N_14187,N_13767);
and U14682 (N_14682,N_13528,N_14043);
or U14683 (N_14683,N_14134,N_13924);
nor U14684 (N_14684,N_13622,N_14085);
nand U14685 (N_14685,N_13820,N_13584);
nor U14686 (N_14686,N_14181,N_14175);
nor U14687 (N_14687,N_14199,N_13936);
and U14688 (N_14688,N_14051,N_13969);
nand U14689 (N_14689,N_13595,N_13642);
or U14690 (N_14690,N_13799,N_13914);
nand U14691 (N_14691,N_13619,N_13576);
nand U14692 (N_14692,N_13836,N_13617);
and U14693 (N_14693,N_14135,N_14220);
nor U14694 (N_14694,N_13618,N_13561);
nand U14695 (N_14695,N_13868,N_13831);
nand U14696 (N_14696,N_13640,N_13957);
xnor U14697 (N_14697,N_14082,N_14143);
and U14698 (N_14698,N_14182,N_13898);
nor U14699 (N_14699,N_14090,N_13924);
and U14700 (N_14700,N_14135,N_13897);
and U14701 (N_14701,N_13531,N_13970);
and U14702 (N_14702,N_13558,N_13640);
xnor U14703 (N_14703,N_13929,N_13544);
nor U14704 (N_14704,N_13621,N_14067);
nand U14705 (N_14705,N_14072,N_14099);
nand U14706 (N_14706,N_13643,N_14231);
nand U14707 (N_14707,N_13664,N_13541);
and U14708 (N_14708,N_14140,N_13766);
xnor U14709 (N_14709,N_13971,N_14239);
xor U14710 (N_14710,N_13544,N_14198);
nor U14711 (N_14711,N_13678,N_13590);
nor U14712 (N_14712,N_14102,N_13848);
or U14713 (N_14713,N_13566,N_14153);
and U14714 (N_14714,N_14167,N_13913);
or U14715 (N_14715,N_13619,N_13886);
or U14716 (N_14716,N_13666,N_13891);
or U14717 (N_14717,N_13953,N_13987);
nand U14718 (N_14718,N_13610,N_14109);
and U14719 (N_14719,N_13576,N_13703);
nor U14720 (N_14720,N_13571,N_14046);
nand U14721 (N_14721,N_14049,N_13822);
nor U14722 (N_14722,N_13926,N_13658);
or U14723 (N_14723,N_13975,N_13578);
nand U14724 (N_14724,N_13960,N_13954);
nor U14725 (N_14725,N_14141,N_13588);
or U14726 (N_14726,N_14144,N_13705);
nand U14727 (N_14727,N_14010,N_13689);
nand U14728 (N_14728,N_13644,N_14049);
nor U14729 (N_14729,N_13613,N_14067);
nor U14730 (N_14730,N_14229,N_13970);
nor U14731 (N_14731,N_13773,N_13770);
and U14732 (N_14732,N_14011,N_13525);
or U14733 (N_14733,N_14020,N_13774);
and U14734 (N_14734,N_14124,N_13725);
nand U14735 (N_14735,N_14169,N_14034);
and U14736 (N_14736,N_14056,N_14058);
xor U14737 (N_14737,N_13579,N_13676);
nand U14738 (N_14738,N_14211,N_13787);
nand U14739 (N_14739,N_13526,N_13807);
nor U14740 (N_14740,N_13500,N_13913);
nor U14741 (N_14741,N_13652,N_14224);
nand U14742 (N_14742,N_13700,N_14080);
or U14743 (N_14743,N_13552,N_13891);
xnor U14744 (N_14744,N_13580,N_13536);
or U14745 (N_14745,N_13695,N_14175);
or U14746 (N_14746,N_13570,N_13814);
nand U14747 (N_14747,N_13961,N_13917);
nor U14748 (N_14748,N_14128,N_13725);
nor U14749 (N_14749,N_14086,N_13620);
and U14750 (N_14750,N_14169,N_13767);
and U14751 (N_14751,N_14175,N_14167);
xnor U14752 (N_14752,N_13769,N_14010);
and U14753 (N_14753,N_13859,N_13927);
or U14754 (N_14754,N_14241,N_14211);
and U14755 (N_14755,N_14194,N_13565);
nor U14756 (N_14756,N_13764,N_14207);
and U14757 (N_14757,N_13508,N_13742);
nand U14758 (N_14758,N_13654,N_13668);
nor U14759 (N_14759,N_14206,N_14017);
nand U14760 (N_14760,N_14199,N_13796);
xor U14761 (N_14761,N_13958,N_14024);
and U14762 (N_14762,N_13701,N_14064);
nand U14763 (N_14763,N_14110,N_14154);
and U14764 (N_14764,N_14024,N_13943);
nor U14765 (N_14765,N_14139,N_13648);
or U14766 (N_14766,N_14019,N_13897);
xnor U14767 (N_14767,N_13801,N_14157);
and U14768 (N_14768,N_13888,N_13892);
nand U14769 (N_14769,N_14230,N_13757);
and U14770 (N_14770,N_13804,N_14206);
nor U14771 (N_14771,N_13579,N_13978);
or U14772 (N_14772,N_14018,N_14152);
and U14773 (N_14773,N_13830,N_13934);
nor U14774 (N_14774,N_14170,N_13727);
and U14775 (N_14775,N_13662,N_14229);
and U14776 (N_14776,N_13564,N_13561);
and U14777 (N_14777,N_13701,N_13881);
or U14778 (N_14778,N_14180,N_13770);
and U14779 (N_14779,N_13775,N_13518);
or U14780 (N_14780,N_13905,N_13846);
nor U14781 (N_14781,N_14216,N_13974);
xor U14782 (N_14782,N_13517,N_14066);
xor U14783 (N_14783,N_13583,N_13504);
nor U14784 (N_14784,N_13809,N_13614);
nor U14785 (N_14785,N_14208,N_13892);
xnor U14786 (N_14786,N_13594,N_13918);
and U14787 (N_14787,N_14031,N_13598);
and U14788 (N_14788,N_13909,N_13738);
nand U14789 (N_14789,N_14039,N_14049);
xor U14790 (N_14790,N_13568,N_13661);
nand U14791 (N_14791,N_14143,N_14208);
and U14792 (N_14792,N_13786,N_13816);
nand U14793 (N_14793,N_14009,N_13673);
nor U14794 (N_14794,N_13863,N_13600);
and U14795 (N_14795,N_13972,N_14141);
and U14796 (N_14796,N_13831,N_13641);
nor U14797 (N_14797,N_13841,N_14021);
and U14798 (N_14798,N_13641,N_13819);
and U14799 (N_14799,N_13901,N_13626);
or U14800 (N_14800,N_13574,N_13604);
xor U14801 (N_14801,N_13700,N_14159);
nand U14802 (N_14802,N_13619,N_13936);
and U14803 (N_14803,N_14093,N_13939);
nor U14804 (N_14804,N_14192,N_13908);
or U14805 (N_14805,N_14019,N_13764);
xor U14806 (N_14806,N_14119,N_14162);
and U14807 (N_14807,N_14092,N_14115);
nand U14808 (N_14808,N_13539,N_13908);
or U14809 (N_14809,N_14214,N_14103);
or U14810 (N_14810,N_13726,N_13707);
nand U14811 (N_14811,N_13672,N_13832);
nand U14812 (N_14812,N_14192,N_13798);
or U14813 (N_14813,N_14038,N_14212);
nand U14814 (N_14814,N_14205,N_13759);
nand U14815 (N_14815,N_13585,N_13910);
nor U14816 (N_14816,N_13994,N_14098);
and U14817 (N_14817,N_13538,N_14236);
or U14818 (N_14818,N_13743,N_14164);
or U14819 (N_14819,N_13975,N_13933);
nor U14820 (N_14820,N_13572,N_14183);
and U14821 (N_14821,N_14120,N_14125);
or U14822 (N_14822,N_14134,N_14126);
or U14823 (N_14823,N_14247,N_13621);
nand U14824 (N_14824,N_14001,N_14222);
nor U14825 (N_14825,N_14196,N_13561);
or U14826 (N_14826,N_13745,N_14211);
xor U14827 (N_14827,N_13849,N_13676);
and U14828 (N_14828,N_13532,N_13705);
and U14829 (N_14829,N_13939,N_14162);
and U14830 (N_14830,N_13782,N_13793);
nand U14831 (N_14831,N_14162,N_13961);
xnor U14832 (N_14832,N_13529,N_13846);
or U14833 (N_14833,N_14183,N_13503);
or U14834 (N_14834,N_14030,N_13663);
and U14835 (N_14835,N_13646,N_14114);
nand U14836 (N_14836,N_13751,N_14235);
and U14837 (N_14837,N_13871,N_14056);
nor U14838 (N_14838,N_13782,N_13699);
nor U14839 (N_14839,N_14237,N_13884);
and U14840 (N_14840,N_14182,N_13731);
nor U14841 (N_14841,N_13845,N_13689);
nand U14842 (N_14842,N_14152,N_13971);
and U14843 (N_14843,N_13666,N_13675);
nand U14844 (N_14844,N_13597,N_13838);
xnor U14845 (N_14845,N_13981,N_13681);
and U14846 (N_14846,N_13949,N_13675);
nor U14847 (N_14847,N_13975,N_14174);
nand U14848 (N_14848,N_13962,N_14077);
or U14849 (N_14849,N_13613,N_14106);
nand U14850 (N_14850,N_13655,N_13864);
and U14851 (N_14851,N_13899,N_14099);
nand U14852 (N_14852,N_13826,N_14091);
xor U14853 (N_14853,N_13982,N_14001);
or U14854 (N_14854,N_13748,N_14232);
and U14855 (N_14855,N_13928,N_13689);
nor U14856 (N_14856,N_13838,N_13765);
or U14857 (N_14857,N_13547,N_13814);
nor U14858 (N_14858,N_13729,N_14037);
nand U14859 (N_14859,N_14041,N_13822);
nor U14860 (N_14860,N_14137,N_13515);
and U14861 (N_14861,N_14168,N_14007);
or U14862 (N_14862,N_13562,N_13690);
or U14863 (N_14863,N_13525,N_14024);
nor U14864 (N_14864,N_13805,N_13516);
nor U14865 (N_14865,N_13592,N_14130);
or U14866 (N_14866,N_14096,N_13827);
and U14867 (N_14867,N_13843,N_14150);
nand U14868 (N_14868,N_13517,N_13952);
nor U14869 (N_14869,N_13771,N_14042);
xnor U14870 (N_14870,N_13725,N_14163);
nor U14871 (N_14871,N_14053,N_13728);
nor U14872 (N_14872,N_14191,N_14096);
nor U14873 (N_14873,N_13930,N_13706);
and U14874 (N_14874,N_13518,N_13739);
or U14875 (N_14875,N_13942,N_13951);
or U14876 (N_14876,N_13858,N_14199);
xor U14877 (N_14877,N_14133,N_14184);
or U14878 (N_14878,N_13684,N_13890);
xnor U14879 (N_14879,N_13917,N_13607);
or U14880 (N_14880,N_13886,N_13667);
nand U14881 (N_14881,N_13854,N_14164);
nand U14882 (N_14882,N_13919,N_13857);
xor U14883 (N_14883,N_13566,N_13540);
and U14884 (N_14884,N_14116,N_14007);
or U14885 (N_14885,N_14107,N_14230);
xor U14886 (N_14886,N_13623,N_14047);
xor U14887 (N_14887,N_14079,N_13942);
xor U14888 (N_14888,N_14007,N_13850);
and U14889 (N_14889,N_13632,N_13502);
or U14890 (N_14890,N_13868,N_13722);
or U14891 (N_14891,N_13900,N_13732);
nand U14892 (N_14892,N_14062,N_13841);
or U14893 (N_14893,N_13829,N_13803);
nor U14894 (N_14894,N_14018,N_13647);
and U14895 (N_14895,N_14199,N_13979);
nand U14896 (N_14896,N_13662,N_13923);
and U14897 (N_14897,N_14102,N_13804);
or U14898 (N_14898,N_13865,N_13934);
or U14899 (N_14899,N_13968,N_14034);
and U14900 (N_14900,N_13951,N_14241);
nand U14901 (N_14901,N_13653,N_14044);
or U14902 (N_14902,N_14096,N_13539);
nor U14903 (N_14903,N_13815,N_13636);
nor U14904 (N_14904,N_13600,N_14180);
and U14905 (N_14905,N_13573,N_14035);
nor U14906 (N_14906,N_14184,N_14222);
xor U14907 (N_14907,N_14067,N_13768);
and U14908 (N_14908,N_14220,N_13830);
nand U14909 (N_14909,N_13585,N_13717);
and U14910 (N_14910,N_14122,N_13782);
or U14911 (N_14911,N_13706,N_14167);
xnor U14912 (N_14912,N_13981,N_13719);
nor U14913 (N_14913,N_13592,N_14028);
or U14914 (N_14914,N_13505,N_13729);
and U14915 (N_14915,N_13593,N_13834);
nor U14916 (N_14916,N_13666,N_14025);
nand U14917 (N_14917,N_13754,N_14148);
nand U14918 (N_14918,N_13780,N_14183);
or U14919 (N_14919,N_13796,N_14187);
or U14920 (N_14920,N_13756,N_13841);
nor U14921 (N_14921,N_13883,N_13784);
nor U14922 (N_14922,N_13840,N_13903);
nor U14923 (N_14923,N_13983,N_13652);
or U14924 (N_14924,N_13932,N_13957);
xnor U14925 (N_14925,N_13506,N_13805);
or U14926 (N_14926,N_13826,N_14111);
xor U14927 (N_14927,N_13561,N_13518);
and U14928 (N_14928,N_14150,N_13663);
or U14929 (N_14929,N_13846,N_14105);
xnor U14930 (N_14930,N_13968,N_13521);
nor U14931 (N_14931,N_13922,N_14021);
xor U14932 (N_14932,N_13869,N_14049);
or U14933 (N_14933,N_14240,N_14159);
and U14934 (N_14934,N_13988,N_14114);
nor U14935 (N_14935,N_13585,N_13942);
xnor U14936 (N_14936,N_14098,N_14190);
or U14937 (N_14937,N_14064,N_13896);
nor U14938 (N_14938,N_13595,N_13873);
nand U14939 (N_14939,N_13990,N_13887);
and U14940 (N_14940,N_13715,N_14187);
nor U14941 (N_14941,N_13775,N_14196);
nand U14942 (N_14942,N_14183,N_13792);
nand U14943 (N_14943,N_14236,N_13553);
nor U14944 (N_14944,N_13632,N_13564);
nand U14945 (N_14945,N_13674,N_14244);
nand U14946 (N_14946,N_14205,N_13821);
or U14947 (N_14947,N_13599,N_14240);
xor U14948 (N_14948,N_13861,N_13940);
or U14949 (N_14949,N_13517,N_13865);
nor U14950 (N_14950,N_14230,N_13695);
and U14951 (N_14951,N_13726,N_14083);
and U14952 (N_14952,N_13686,N_13667);
nand U14953 (N_14953,N_13893,N_13703);
or U14954 (N_14954,N_13971,N_14207);
nand U14955 (N_14955,N_13508,N_13970);
nor U14956 (N_14956,N_14151,N_13515);
nor U14957 (N_14957,N_14218,N_13609);
nor U14958 (N_14958,N_14215,N_13636);
xnor U14959 (N_14959,N_14069,N_14053);
nand U14960 (N_14960,N_13892,N_14214);
and U14961 (N_14961,N_14195,N_13573);
and U14962 (N_14962,N_13960,N_14224);
xor U14963 (N_14963,N_13853,N_13705);
or U14964 (N_14964,N_13586,N_13980);
nor U14965 (N_14965,N_13691,N_13827);
nand U14966 (N_14966,N_13901,N_14089);
nand U14967 (N_14967,N_13909,N_13856);
and U14968 (N_14968,N_14107,N_14175);
nand U14969 (N_14969,N_14139,N_14023);
nand U14970 (N_14970,N_14166,N_13916);
and U14971 (N_14971,N_13583,N_13881);
or U14972 (N_14972,N_14190,N_13572);
nand U14973 (N_14973,N_13873,N_14211);
and U14974 (N_14974,N_13767,N_13673);
or U14975 (N_14975,N_13672,N_13525);
or U14976 (N_14976,N_13709,N_14028);
nor U14977 (N_14977,N_14148,N_13720);
nand U14978 (N_14978,N_14201,N_13650);
nor U14979 (N_14979,N_14043,N_13784);
xnor U14980 (N_14980,N_13794,N_13749);
and U14981 (N_14981,N_13777,N_13631);
xnor U14982 (N_14982,N_13658,N_13815);
or U14983 (N_14983,N_13866,N_13535);
or U14984 (N_14984,N_13597,N_13588);
or U14985 (N_14985,N_14220,N_14072);
nand U14986 (N_14986,N_14245,N_13616);
or U14987 (N_14987,N_13981,N_13575);
nand U14988 (N_14988,N_14143,N_13634);
nor U14989 (N_14989,N_13921,N_13756);
and U14990 (N_14990,N_14007,N_14240);
xnor U14991 (N_14991,N_14052,N_13715);
nand U14992 (N_14992,N_13700,N_14007);
nand U14993 (N_14993,N_13549,N_14203);
or U14994 (N_14994,N_13928,N_13673);
nor U14995 (N_14995,N_13530,N_14174);
and U14996 (N_14996,N_14056,N_14087);
or U14997 (N_14997,N_14001,N_13779);
and U14998 (N_14998,N_13715,N_14120);
or U14999 (N_14999,N_13713,N_13810);
nor UO_0 (O_0,N_14777,N_14591);
and UO_1 (O_1,N_14336,N_14634);
or UO_2 (O_2,N_14431,N_14364);
or UO_3 (O_3,N_14271,N_14326);
nand UO_4 (O_4,N_14656,N_14792);
and UO_5 (O_5,N_14304,N_14417);
nor UO_6 (O_6,N_14895,N_14318);
nor UO_7 (O_7,N_14558,N_14530);
nor UO_8 (O_8,N_14465,N_14801);
nand UO_9 (O_9,N_14638,N_14621);
nand UO_10 (O_10,N_14712,N_14775);
nand UO_11 (O_11,N_14316,N_14509);
nand UO_12 (O_12,N_14480,N_14323);
xnor UO_13 (O_13,N_14309,N_14719);
or UO_14 (O_14,N_14793,N_14280);
and UO_15 (O_15,N_14491,N_14628);
nor UO_16 (O_16,N_14612,N_14637);
nand UO_17 (O_17,N_14731,N_14373);
nand UO_18 (O_18,N_14305,N_14814);
nand UO_19 (O_19,N_14794,N_14698);
nand UO_20 (O_20,N_14493,N_14359);
and UO_21 (O_21,N_14481,N_14424);
or UO_22 (O_22,N_14447,N_14723);
or UO_23 (O_23,N_14541,N_14544);
nand UO_24 (O_24,N_14626,N_14702);
nor UO_25 (O_25,N_14752,N_14331);
nand UO_26 (O_26,N_14746,N_14533);
and UO_27 (O_27,N_14771,N_14349);
nand UO_28 (O_28,N_14843,N_14543);
and UO_29 (O_29,N_14337,N_14776);
or UO_30 (O_30,N_14573,N_14880);
and UO_31 (O_31,N_14958,N_14460);
and UO_32 (O_32,N_14498,N_14401);
nand UO_33 (O_33,N_14461,N_14453);
nor UO_34 (O_34,N_14837,N_14851);
or UO_35 (O_35,N_14390,N_14609);
or UO_36 (O_36,N_14984,N_14863);
and UO_37 (O_37,N_14898,N_14691);
or UO_38 (O_38,N_14583,N_14665);
nor UO_39 (O_39,N_14329,N_14919);
and UO_40 (O_40,N_14520,N_14687);
or UO_41 (O_41,N_14765,N_14388);
nand UO_42 (O_42,N_14586,N_14273);
and UO_43 (O_43,N_14299,N_14470);
and UO_44 (O_44,N_14743,N_14817);
xor UO_45 (O_45,N_14720,N_14269);
or UO_46 (O_46,N_14791,N_14615);
nor UO_47 (O_47,N_14995,N_14462);
nand UO_48 (O_48,N_14864,N_14695);
nand UO_49 (O_49,N_14866,N_14398);
and UO_50 (O_50,N_14421,N_14824);
nor UO_51 (O_51,N_14685,N_14601);
and UO_52 (O_52,N_14593,N_14550);
nor UO_53 (O_53,N_14250,N_14726);
xor UO_54 (O_54,N_14913,N_14450);
or UO_55 (O_55,N_14699,N_14799);
or UO_56 (O_56,N_14848,N_14989);
or UO_57 (O_57,N_14836,N_14857);
nand UO_58 (O_58,N_14721,N_14361);
nand UO_59 (O_59,N_14287,N_14606);
nor UO_60 (O_60,N_14713,N_14556);
and UO_61 (O_61,N_14395,N_14796);
nand UO_62 (O_62,N_14434,N_14384);
nor UO_63 (O_63,N_14839,N_14876);
nor UO_64 (O_64,N_14408,N_14522);
nor UO_65 (O_65,N_14483,N_14321);
or UO_66 (O_66,N_14734,N_14703);
nand UO_67 (O_67,N_14584,N_14741);
or UO_68 (O_68,N_14312,N_14567);
nand UO_69 (O_69,N_14887,N_14600);
nor UO_70 (O_70,N_14399,N_14875);
nor UO_71 (O_71,N_14582,N_14298);
or UO_72 (O_72,N_14565,N_14649);
and UO_73 (O_73,N_14804,N_14890);
xor UO_74 (O_74,N_14406,N_14262);
and UO_75 (O_75,N_14885,N_14708);
or UO_76 (O_76,N_14579,N_14816);
nand UO_77 (O_77,N_14983,N_14997);
or UO_78 (O_78,N_14260,N_14732);
nor UO_79 (O_79,N_14652,N_14670);
xnor UO_80 (O_80,N_14553,N_14345);
nand UO_81 (O_81,N_14275,N_14594);
or UO_82 (O_82,N_14286,N_14682);
and UO_83 (O_83,N_14371,N_14844);
nor UO_84 (O_84,N_14976,N_14631);
nor UO_85 (O_85,N_14290,N_14996);
nand UO_86 (O_86,N_14254,N_14947);
nor UO_87 (O_87,N_14500,N_14646);
nor UO_88 (O_88,N_14448,N_14454);
nand UO_89 (O_89,N_14383,N_14803);
and UO_90 (O_90,N_14639,N_14295);
or UO_91 (O_91,N_14788,N_14724);
or UO_92 (O_92,N_14856,N_14955);
or UO_93 (O_93,N_14733,N_14469);
nand UO_94 (O_94,N_14297,N_14575);
or UO_95 (O_95,N_14458,N_14907);
xnor UO_96 (O_96,N_14473,N_14671);
nor UO_97 (O_97,N_14802,N_14999);
nand UO_98 (O_98,N_14320,N_14663);
or UO_99 (O_99,N_14283,N_14915);
and UO_100 (O_100,N_14444,N_14869);
nand UO_101 (O_101,N_14756,N_14715);
nor UO_102 (O_102,N_14742,N_14909);
and UO_103 (O_103,N_14430,N_14987);
and UO_104 (O_104,N_14466,N_14605);
nand UO_105 (O_105,N_14314,N_14945);
and UO_106 (O_106,N_14954,N_14369);
nand UO_107 (O_107,N_14833,N_14459);
and UO_108 (O_108,N_14492,N_14879);
nor UO_109 (O_109,N_14753,N_14659);
nand UO_110 (O_110,N_14904,N_14402);
nand UO_111 (O_111,N_14420,N_14896);
nand UO_112 (O_112,N_14252,N_14957);
nand UO_113 (O_113,N_14868,N_14348);
or UO_114 (O_114,N_14964,N_14538);
nor UO_115 (O_115,N_14378,N_14881);
nand UO_116 (O_116,N_14767,N_14438);
and UO_117 (O_117,N_14764,N_14251);
or UO_118 (O_118,N_14668,N_14738);
nand UO_119 (O_119,N_14938,N_14974);
and UO_120 (O_120,N_14647,N_14531);
or UO_121 (O_121,N_14437,N_14784);
or UO_122 (O_122,N_14524,N_14446);
nand UO_123 (O_123,N_14820,N_14674);
xnor UO_124 (O_124,N_14324,N_14877);
or UO_125 (O_125,N_14683,N_14347);
nor UO_126 (O_126,N_14534,N_14279);
nor UO_127 (O_127,N_14405,N_14427);
or UO_128 (O_128,N_14559,N_14404);
nor UO_129 (O_129,N_14257,N_14464);
xor UO_130 (O_130,N_14570,N_14303);
nor UO_131 (O_131,N_14554,N_14797);
xor UO_132 (O_132,N_14416,N_14499);
nor UO_133 (O_133,N_14980,N_14463);
nor UO_134 (O_134,N_14903,N_14867);
and UO_135 (O_135,N_14707,N_14572);
nor UO_136 (O_136,N_14512,N_14435);
nor UO_137 (O_137,N_14255,N_14930);
or UO_138 (O_138,N_14519,N_14711);
nand UO_139 (O_139,N_14979,N_14624);
or UO_140 (O_140,N_14937,N_14315);
or UO_141 (O_141,N_14267,N_14334);
nor UO_142 (O_142,N_14479,N_14916);
nor UO_143 (O_143,N_14561,N_14672);
or UO_144 (O_144,N_14905,N_14396);
nand UO_145 (O_145,N_14566,N_14343);
nand UO_146 (O_146,N_14829,N_14942);
nor UO_147 (O_147,N_14488,N_14346);
or UO_148 (O_148,N_14988,N_14912);
nor UO_149 (O_149,N_14341,N_14823);
nor UO_150 (O_150,N_14555,N_14722);
and UO_151 (O_151,N_14736,N_14883);
nor UO_152 (O_152,N_14356,N_14840);
nand UO_153 (O_153,N_14878,N_14363);
and UO_154 (O_154,N_14889,N_14443);
nor UO_155 (O_155,N_14884,N_14353);
nor UO_156 (O_156,N_14274,N_14855);
xor UO_157 (O_157,N_14366,N_14525);
or UO_158 (O_158,N_14285,N_14832);
nor UO_159 (O_159,N_14578,N_14648);
and UO_160 (O_160,N_14658,N_14414);
nand UO_161 (O_161,N_14622,N_14679);
nor UO_162 (O_162,N_14928,N_14809);
nand UO_163 (O_163,N_14319,N_14675);
nor UO_164 (O_164,N_14783,N_14619);
and UO_165 (O_165,N_14350,N_14815);
or UO_166 (O_166,N_14908,N_14636);
and UO_167 (O_167,N_14690,N_14633);
xnor UO_168 (O_168,N_14362,N_14494);
and UO_169 (O_169,N_14412,N_14825);
nand UO_170 (O_170,N_14951,N_14476);
nor UO_171 (O_171,N_14564,N_14497);
or UO_172 (O_172,N_14900,N_14882);
or UO_173 (O_173,N_14749,N_14993);
or UO_174 (O_174,N_14986,N_14680);
or UO_175 (O_175,N_14923,N_14874);
nor UO_176 (O_176,N_14313,N_14961);
nor UO_177 (O_177,N_14360,N_14835);
xor UO_178 (O_178,N_14354,N_14693);
nor UO_179 (O_179,N_14514,N_14965);
xnor UO_180 (O_180,N_14562,N_14744);
and UO_181 (O_181,N_14689,N_14676);
or UO_182 (O_182,N_14568,N_14697);
nor UO_183 (O_183,N_14939,N_14827);
or UO_184 (O_184,N_14990,N_14985);
and UO_185 (O_185,N_14505,N_14629);
nand UO_186 (O_186,N_14375,N_14546);
nor UO_187 (O_187,N_14714,N_14892);
or UO_188 (O_188,N_14782,N_14580);
or UO_189 (O_189,N_14599,N_14261);
nand UO_190 (O_190,N_14858,N_14934);
or UO_191 (O_191,N_14760,N_14798);
and UO_192 (O_192,N_14778,N_14397);
or UO_193 (O_193,N_14620,N_14467);
xor UO_194 (O_194,N_14413,N_14376);
nand UO_195 (O_195,N_14661,N_14490);
and UO_196 (O_196,N_14651,N_14484);
xnor UO_197 (O_197,N_14841,N_14992);
nand UO_198 (O_198,N_14452,N_14681);
or UO_199 (O_199,N_14696,N_14935);
xnor UO_200 (O_200,N_14655,N_14774);
and UO_201 (O_201,N_14627,N_14577);
and UO_202 (O_202,N_14834,N_14641);
nand UO_203 (O_203,N_14901,N_14307);
or UO_204 (O_204,N_14779,N_14865);
nand UO_205 (O_205,N_14547,N_14914);
xnor UO_206 (O_206,N_14339,N_14830);
nand UO_207 (O_207,N_14969,N_14282);
or UO_208 (O_208,N_14515,N_14933);
nor UO_209 (O_209,N_14503,N_14991);
nor UO_210 (O_210,N_14924,N_14411);
nand UO_211 (O_211,N_14468,N_14560);
xnor UO_212 (O_212,N_14773,N_14894);
and UO_213 (O_213,N_14949,N_14277);
nor UO_214 (O_214,N_14664,N_14610);
or UO_215 (O_215,N_14603,N_14813);
and UO_216 (O_216,N_14539,N_14811);
and UO_217 (O_217,N_14569,N_14872);
nand UO_218 (O_218,N_14268,N_14686);
nand UO_219 (O_219,N_14739,N_14666);
nand UO_220 (O_220,N_14477,N_14852);
or UO_221 (O_221,N_14407,N_14978);
and UO_222 (O_222,N_14296,N_14367);
nand UO_223 (O_223,N_14486,N_14948);
or UO_224 (O_224,N_14998,N_14596);
or UO_225 (O_225,N_14728,N_14870);
nand UO_226 (O_226,N_14902,N_14706);
nand UO_227 (O_227,N_14625,N_14944);
or UO_228 (O_228,N_14849,N_14873);
and UO_229 (O_229,N_14755,N_14293);
and UO_230 (O_230,N_14950,N_14786);
nor UO_231 (O_231,N_14662,N_14700);
nor UO_232 (O_232,N_14781,N_14588);
nand UO_233 (O_233,N_14673,N_14403);
xnor UO_234 (O_234,N_14705,N_14335);
or UO_235 (O_235,N_14410,N_14936);
or UO_236 (O_236,N_14270,N_14385);
and UO_237 (O_237,N_14602,N_14684);
or UO_238 (O_238,N_14436,N_14451);
nor UO_239 (O_239,N_14308,N_14787);
xnor UO_240 (O_240,N_14482,N_14504);
nor UO_241 (O_241,N_14968,N_14332);
xnor UO_242 (O_242,N_14845,N_14740);
or UO_243 (O_243,N_14472,N_14807);
nand UO_244 (O_244,N_14428,N_14611);
nand UO_245 (O_245,N_14276,N_14821);
xnor UO_246 (O_246,N_14838,N_14630);
nand UO_247 (O_247,N_14501,N_14891);
nand UO_248 (O_248,N_14338,N_14392);
and UO_249 (O_249,N_14805,N_14812);
or UO_250 (O_250,N_14704,N_14517);
xnor UO_251 (O_251,N_14425,N_14644);
nand UO_252 (O_252,N_14393,N_14532);
and UO_253 (O_253,N_14943,N_14529);
nor UO_254 (O_254,N_14598,N_14946);
nand UO_255 (O_255,N_14327,N_14551);
nor UO_256 (O_256,N_14643,N_14439);
nand UO_257 (O_257,N_14545,N_14850);
nand UO_258 (O_258,N_14391,N_14495);
or UO_259 (O_259,N_14745,N_14342);
nor UO_260 (O_260,N_14351,N_14918);
xor UO_261 (O_261,N_14291,N_14677);
nor UO_262 (O_262,N_14485,N_14333);
and UO_263 (O_263,N_14374,N_14800);
and UO_264 (O_264,N_14613,N_14846);
or UO_265 (O_265,N_14853,N_14789);
nand UO_266 (O_266,N_14932,N_14737);
nor UO_267 (O_267,N_14272,N_14842);
and UO_268 (O_268,N_14906,N_14552);
nand UO_269 (O_269,N_14692,N_14502);
nor UO_270 (O_270,N_14311,N_14761);
nand UO_271 (O_271,N_14340,N_14576);
nand UO_272 (O_272,N_14859,N_14506);
or UO_273 (O_273,N_14440,N_14810);
nand UO_274 (O_274,N_14607,N_14862);
or UO_275 (O_275,N_14716,N_14288);
nor UO_276 (O_276,N_14328,N_14831);
and UO_277 (O_277,N_14614,N_14608);
and UO_278 (O_278,N_14701,N_14899);
and UO_279 (O_279,N_14527,N_14667);
and UO_280 (O_280,N_14432,N_14590);
or UO_281 (O_281,N_14478,N_14973);
nor UO_282 (O_282,N_14409,N_14292);
nand UO_283 (O_283,N_14886,N_14357);
nand UO_284 (O_284,N_14861,N_14785);
nor UO_285 (O_285,N_14618,N_14808);
nor UO_286 (O_286,N_14735,N_14927);
and UO_287 (O_287,N_14475,N_14709);
and UO_288 (O_288,N_14653,N_14289);
nor UO_289 (O_289,N_14368,N_14795);
or UO_290 (O_290,N_14557,N_14669);
and UO_291 (O_291,N_14977,N_14920);
nand UO_292 (O_292,N_14826,N_14718);
nand UO_293 (O_293,N_14370,N_14616);
and UO_294 (O_294,N_14967,N_14763);
nand UO_295 (O_295,N_14635,N_14516);
xnor UO_296 (O_296,N_14768,N_14394);
nor UO_297 (O_297,N_14489,N_14381);
and UO_298 (O_298,N_14971,N_14994);
nand UO_299 (O_299,N_14860,N_14650);
and UO_300 (O_300,N_14322,N_14278);
nor UO_301 (O_301,N_14940,N_14422);
or UO_302 (O_302,N_14387,N_14429);
nor UO_303 (O_303,N_14317,N_14926);
xnor UO_304 (O_304,N_14963,N_14352);
or UO_305 (O_305,N_14548,N_14365);
or UO_306 (O_306,N_14597,N_14748);
nor UO_307 (O_307,N_14847,N_14688);
or UO_308 (O_308,N_14623,N_14389);
and UO_309 (O_309,N_14523,N_14377);
or UO_310 (O_310,N_14344,N_14266);
or UO_311 (O_311,N_14581,N_14717);
nor UO_312 (O_312,N_14960,N_14972);
or UO_313 (O_313,N_14921,N_14474);
and UO_314 (O_314,N_14910,N_14300);
nand UO_315 (O_315,N_14540,N_14487);
nor UO_316 (O_316,N_14264,N_14981);
nand UO_317 (O_317,N_14511,N_14871);
or UO_318 (O_318,N_14507,N_14589);
xor UO_319 (O_319,N_14790,N_14710);
and UO_320 (O_320,N_14975,N_14754);
nor UO_321 (O_321,N_14526,N_14645);
nor UO_322 (O_322,N_14521,N_14772);
nor UO_323 (O_323,N_14513,N_14595);
or UO_324 (O_324,N_14694,N_14571);
and UO_325 (O_325,N_14604,N_14496);
or UO_326 (O_326,N_14982,N_14415);
nor UO_327 (O_327,N_14418,N_14654);
and UO_328 (O_328,N_14330,N_14535);
or UO_329 (O_329,N_14426,N_14657);
or UO_330 (O_330,N_14959,N_14542);
nand UO_331 (O_331,N_14727,N_14893);
or UO_332 (O_332,N_14725,N_14358);
nor UO_333 (O_333,N_14730,N_14660);
and UO_334 (O_334,N_14762,N_14751);
or UO_335 (O_335,N_14617,N_14445);
and UO_336 (O_336,N_14956,N_14750);
nor UO_337 (O_337,N_14585,N_14563);
and UO_338 (O_338,N_14766,N_14758);
nor UO_339 (O_339,N_14528,N_14953);
or UO_340 (O_340,N_14510,N_14380);
nor UO_341 (O_341,N_14549,N_14355);
nor UO_342 (O_342,N_14382,N_14302);
and UO_343 (O_343,N_14441,N_14931);
and UO_344 (O_344,N_14433,N_14423);
nand UO_345 (O_345,N_14386,N_14253);
nor UO_346 (O_346,N_14301,N_14457);
nand UO_347 (O_347,N_14537,N_14941);
or UO_348 (O_348,N_14592,N_14419);
or UO_349 (O_349,N_14455,N_14284);
xor UO_350 (O_350,N_14966,N_14379);
xnor UO_351 (O_351,N_14281,N_14897);
nor UO_352 (O_352,N_14574,N_14929);
and UO_353 (O_353,N_14632,N_14265);
nand UO_354 (O_354,N_14888,N_14449);
and UO_355 (O_355,N_14828,N_14911);
nand UO_356 (O_356,N_14922,N_14508);
xnor UO_357 (O_357,N_14471,N_14256);
and UO_358 (O_358,N_14806,N_14259);
xnor UO_359 (O_359,N_14400,N_14678);
and UO_360 (O_360,N_14640,N_14518);
or UO_361 (O_361,N_14818,N_14747);
and UO_362 (O_362,N_14442,N_14294);
and UO_363 (O_363,N_14769,N_14962);
nand UO_364 (O_364,N_14372,N_14729);
nand UO_365 (O_365,N_14325,N_14263);
nand UO_366 (O_366,N_14759,N_14536);
and UO_367 (O_367,N_14917,N_14822);
xnor UO_368 (O_368,N_14757,N_14456);
or UO_369 (O_369,N_14925,N_14306);
nor UO_370 (O_370,N_14854,N_14258);
and UO_371 (O_371,N_14952,N_14770);
nand UO_372 (O_372,N_14819,N_14642);
nor UO_373 (O_373,N_14587,N_14970);
nand UO_374 (O_374,N_14310,N_14780);
nand UO_375 (O_375,N_14989,N_14811);
and UO_376 (O_376,N_14429,N_14511);
and UO_377 (O_377,N_14751,N_14699);
xnor UO_378 (O_378,N_14783,N_14672);
and UO_379 (O_379,N_14622,N_14328);
nor UO_380 (O_380,N_14349,N_14911);
and UO_381 (O_381,N_14698,N_14394);
nand UO_382 (O_382,N_14417,N_14732);
and UO_383 (O_383,N_14252,N_14692);
or UO_384 (O_384,N_14290,N_14531);
nand UO_385 (O_385,N_14444,N_14841);
or UO_386 (O_386,N_14380,N_14535);
nor UO_387 (O_387,N_14987,N_14657);
or UO_388 (O_388,N_14395,N_14553);
nand UO_389 (O_389,N_14916,N_14360);
and UO_390 (O_390,N_14495,N_14555);
nand UO_391 (O_391,N_14603,N_14497);
and UO_392 (O_392,N_14345,N_14270);
xnor UO_393 (O_393,N_14489,N_14532);
nand UO_394 (O_394,N_14483,N_14465);
xnor UO_395 (O_395,N_14680,N_14260);
nor UO_396 (O_396,N_14969,N_14833);
nand UO_397 (O_397,N_14370,N_14945);
and UO_398 (O_398,N_14914,N_14726);
or UO_399 (O_399,N_14800,N_14729);
or UO_400 (O_400,N_14260,N_14461);
or UO_401 (O_401,N_14382,N_14377);
nand UO_402 (O_402,N_14347,N_14730);
nor UO_403 (O_403,N_14341,N_14651);
xnor UO_404 (O_404,N_14424,N_14385);
nor UO_405 (O_405,N_14476,N_14496);
xnor UO_406 (O_406,N_14886,N_14964);
or UO_407 (O_407,N_14469,N_14492);
or UO_408 (O_408,N_14800,N_14425);
and UO_409 (O_409,N_14833,N_14621);
or UO_410 (O_410,N_14813,N_14635);
nor UO_411 (O_411,N_14640,N_14617);
or UO_412 (O_412,N_14668,N_14424);
nor UO_413 (O_413,N_14426,N_14313);
and UO_414 (O_414,N_14358,N_14967);
nand UO_415 (O_415,N_14308,N_14811);
nand UO_416 (O_416,N_14437,N_14586);
nor UO_417 (O_417,N_14853,N_14296);
nand UO_418 (O_418,N_14358,N_14386);
and UO_419 (O_419,N_14722,N_14635);
nand UO_420 (O_420,N_14375,N_14279);
nor UO_421 (O_421,N_14793,N_14415);
nand UO_422 (O_422,N_14319,N_14350);
nor UO_423 (O_423,N_14316,N_14288);
nor UO_424 (O_424,N_14787,N_14872);
and UO_425 (O_425,N_14675,N_14444);
and UO_426 (O_426,N_14491,N_14541);
nor UO_427 (O_427,N_14759,N_14575);
nand UO_428 (O_428,N_14776,N_14589);
nand UO_429 (O_429,N_14640,N_14587);
nor UO_430 (O_430,N_14319,N_14397);
or UO_431 (O_431,N_14323,N_14606);
and UO_432 (O_432,N_14582,N_14402);
xor UO_433 (O_433,N_14449,N_14384);
or UO_434 (O_434,N_14813,N_14693);
and UO_435 (O_435,N_14424,N_14594);
nor UO_436 (O_436,N_14824,N_14668);
xor UO_437 (O_437,N_14322,N_14892);
nor UO_438 (O_438,N_14397,N_14725);
and UO_439 (O_439,N_14794,N_14906);
nand UO_440 (O_440,N_14729,N_14603);
and UO_441 (O_441,N_14327,N_14427);
nand UO_442 (O_442,N_14603,N_14693);
xnor UO_443 (O_443,N_14474,N_14313);
or UO_444 (O_444,N_14827,N_14837);
and UO_445 (O_445,N_14263,N_14663);
nor UO_446 (O_446,N_14355,N_14293);
nor UO_447 (O_447,N_14251,N_14979);
nand UO_448 (O_448,N_14575,N_14570);
or UO_449 (O_449,N_14257,N_14773);
or UO_450 (O_450,N_14907,N_14282);
or UO_451 (O_451,N_14647,N_14575);
nor UO_452 (O_452,N_14873,N_14840);
nor UO_453 (O_453,N_14506,N_14635);
xor UO_454 (O_454,N_14764,N_14653);
nor UO_455 (O_455,N_14293,N_14987);
or UO_456 (O_456,N_14445,N_14550);
and UO_457 (O_457,N_14417,N_14734);
and UO_458 (O_458,N_14921,N_14334);
or UO_459 (O_459,N_14823,N_14527);
and UO_460 (O_460,N_14893,N_14723);
xor UO_461 (O_461,N_14744,N_14276);
xnor UO_462 (O_462,N_14759,N_14968);
and UO_463 (O_463,N_14724,N_14453);
nand UO_464 (O_464,N_14657,N_14440);
or UO_465 (O_465,N_14877,N_14591);
nand UO_466 (O_466,N_14470,N_14464);
and UO_467 (O_467,N_14836,N_14264);
and UO_468 (O_468,N_14797,N_14448);
or UO_469 (O_469,N_14503,N_14370);
nor UO_470 (O_470,N_14784,N_14525);
and UO_471 (O_471,N_14295,N_14809);
xnor UO_472 (O_472,N_14603,N_14496);
nor UO_473 (O_473,N_14294,N_14867);
nor UO_474 (O_474,N_14340,N_14889);
and UO_475 (O_475,N_14532,N_14416);
and UO_476 (O_476,N_14348,N_14280);
or UO_477 (O_477,N_14911,N_14673);
xnor UO_478 (O_478,N_14433,N_14552);
xnor UO_479 (O_479,N_14728,N_14899);
or UO_480 (O_480,N_14796,N_14751);
and UO_481 (O_481,N_14444,N_14712);
or UO_482 (O_482,N_14810,N_14721);
nand UO_483 (O_483,N_14377,N_14390);
or UO_484 (O_484,N_14969,N_14402);
or UO_485 (O_485,N_14552,N_14846);
nor UO_486 (O_486,N_14689,N_14416);
nand UO_487 (O_487,N_14438,N_14709);
nand UO_488 (O_488,N_14491,N_14389);
xnor UO_489 (O_489,N_14641,N_14717);
nor UO_490 (O_490,N_14738,N_14306);
and UO_491 (O_491,N_14741,N_14515);
or UO_492 (O_492,N_14333,N_14432);
and UO_493 (O_493,N_14791,N_14905);
nor UO_494 (O_494,N_14630,N_14996);
xor UO_495 (O_495,N_14933,N_14610);
and UO_496 (O_496,N_14266,N_14641);
nor UO_497 (O_497,N_14940,N_14805);
and UO_498 (O_498,N_14282,N_14749);
or UO_499 (O_499,N_14418,N_14728);
nor UO_500 (O_500,N_14259,N_14400);
or UO_501 (O_501,N_14793,N_14582);
and UO_502 (O_502,N_14721,N_14475);
nand UO_503 (O_503,N_14449,N_14687);
nand UO_504 (O_504,N_14780,N_14853);
nor UO_505 (O_505,N_14350,N_14949);
nor UO_506 (O_506,N_14632,N_14899);
or UO_507 (O_507,N_14960,N_14548);
nor UO_508 (O_508,N_14387,N_14833);
and UO_509 (O_509,N_14766,N_14645);
or UO_510 (O_510,N_14544,N_14584);
nor UO_511 (O_511,N_14565,N_14584);
or UO_512 (O_512,N_14572,N_14362);
and UO_513 (O_513,N_14622,N_14904);
and UO_514 (O_514,N_14664,N_14294);
nor UO_515 (O_515,N_14855,N_14631);
and UO_516 (O_516,N_14413,N_14269);
nand UO_517 (O_517,N_14601,N_14260);
nand UO_518 (O_518,N_14572,N_14979);
xnor UO_519 (O_519,N_14872,N_14834);
nand UO_520 (O_520,N_14915,N_14849);
and UO_521 (O_521,N_14761,N_14826);
nor UO_522 (O_522,N_14914,N_14528);
or UO_523 (O_523,N_14413,N_14546);
nand UO_524 (O_524,N_14718,N_14419);
nor UO_525 (O_525,N_14679,N_14944);
xnor UO_526 (O_526,N_14293,N_14360);
and UO_527 (O_527,N_14419,N_14846);
nor UO_528 (O_528,N_14697,N_14745);
nand UO_529 (O_529,N_14412,N_14484);
or UO_530 (O_530,N_14704,N_14851);
nand UO_531 (O_531,N_14264,N_14889);
or UO_532 (O_532,N_14900,N_14447);
nand UO_533 (O_533,N_14956,N_14392);
and UO_534 (O_534,N_14990,N_14443);
and UO_535 (O_535,N_14276,N_14884);
and UO_536 (O_536,N_14638,N_14985);
or UO_537 (O_537,N_14933,N_14285);
and UO_538 (O_538,N_14649,N_14947);
nand UO_539 (O_539,N_14817,N_14448);
or UO_540 (O_540,N_14311,N_14882);
nand UO_541 (O_541,N_14704,N_14901);
and UO_542 (O_542,N_14926,N_14851);
or UO_543 (O_543,N_14798,N_14548);
or UO_544 (O_544,N_14824,N_14980);
nor UO_545 (O_545,N_14413,N_14796);
and UO_546 (O_546,N_14931,N_14744);
or UO_547 (O_547,N_14626,N_14864);
or UO_548 (O_548,N_14699,N_14702);
nor UO_549 (O_549,N_14750,N_14516);
nor UO_550 (O_550,N_14746,N_14400);
xnor UO_551 (O_551,N_14833,N_14370);
nand UO_552 (O_552,N_14486,N_14543);
nand UO_553 (O_553,N_14461,N_14265);
or UO_554 (O_554,N_14605,N_14426);
or UO_555 (O_555,N_14399,N_14869);
and UO_556 (O_556,N_14422,N_14409);
nor UO_557 (O_557,N_14582,N_14258);
xor UO_558 (O_558,N_14364,N_14548);
or UO_559 (O_559,N_14915,N_14599);
and UO_560 (O_560,N_14688,N_14493);
or UO_561 (O_561,N_14550,N_14661);
or UO_562 (O_562,N_14845,N_14376);
and UO_563 (O_563,N_14251,N_14385);
nor UO_564 (O_564,N_14259,N_14306);
and UO_565 (O_565,N_14712,N_14758);
and UO_566 (O_566,N_14867,N_14440);
and UO_567 (O_567,N_14528,N_14355);
and UO_568 (O_568,N_14399,N_14442);
or UO_569 (O_569,N_14301,N_14369);
nor UO_570 (O_570,N_14671,N_14614);
nand UO_571 (O_571,N_14275,N_14515);
or UO_572 (O_572,N_14956,N_14493);
or UO_573 (O_573,N_14546,N_14454);
nand UO_574 (O_574,N_14624,N_14492);
and UO_575 (O_575,N_14412,N_14390);
nand UO_576 (O_576,N_14555,N_14658);
xnor UO_577 (O_577,N_14713,N_14958);
or UO_578 (O_578,N_14872,N_14599);
nand UO_579 (O_579,N_14372,N_14657);
and UO_580 (O_580,N_14571,N_14485);
and UO_581 (O_581,N_14615,N_14497);
and UO_582 (O_582,N_14734,N_14402);
and UO_583 (O_583,N_14473,N_14923);
nor UO_584 (O_584,N_14392,N_14629);
nand UO_585 (O_585,N_14908,N_14982);
and UO_586 (O_586,N_14608,N_14496);
nor UO_587 (O_587,N_14383,N_14403);
nor UO_588 (O_588,N_14915,N_14893);
nor UO_589 (O_589,N_14626,N_14993);
nor UO_590 (O_590,N_14706,N_14709);
xnor UO_591 (O_591,N_14381,N_14675);
nor UO_592 (O_592,N_14926,N_14644);
and UO_593 (O_593,N_14933,N_14736);
or UO_594 (O_594,N_14434,N_14729);
and UO_595 (O_595,N_14250,N_14370);
nand UO_596 (O_596,N_14948,N_14913);
xnor UO_597 (O_597,N_14469,N_14837);
xor UO_598 (O_598,N_14438,N_14882);
or UO_599 (O_599,N_14807,N_14299);
nand UO_600 (O_600,N_14552,N_14858);
nor UO_601 (O_601,N_14405,N_14623);
and UO_602 (O_602,N_14334,N_14905);
nand UO_603 (O_603,N_14876,N_14583);
or UO_604 (O_604,N_14256,N_14466);
nor UO_605 (O_605,N_14379,N_14743);
nand UO_606 (O_606,N_14780,N_14692);
and UO_607 (O_607,N_14318,N_14552);
or UO_608 (O_608,N_14432,N_14542);
xor UO_609 (O_609,N_14393,N_14509);
nand UO_610 (O_610,N_14605,N_14757);
and UO_611 (O_611,N_14401,N_14414);
or UO_612 (O_612,N_14440,N_14272);
xor UO_613 (O_613,N_14422,N_14559);
or UO_614 (O_614,N_14624,N_14270);
and UO_615 (O_615,N_14929,N_14751);
xor UO_616 (O_616,N_14956,N_14541);
nand UO_617 (O_617,N_14394,N_14813);
or UO_618 (O_618,N_14745,N_14530);
or UO_619 (O_619,N_14786,N_14557);
nand UO_620 (O_620,N_14896,N_14626);
nand UO_621 (O_621,N_14807,N_14307);
and UO_622 (O_622,N_14871,N_14764);
or UO_623 (O_623,N_14539,N_14417);
nand UO_624 (O_624,N_14920,N_14418);
xor UO_625 (O_625,N_14772,N_14872);
and UO_626 (O_626,N_14733,N_14497);
nor UO_627 (O_627,N_14705,N_14545);
nor UO_628 (O_628,N_14424,N_14369);
nand UO_629 (O_629,N_14892,N_14372);
nor UO_630 (O_630,N_14362,N_14769);
nor UO_631 (O_631,N_14542,N_14382);
or UO_632 (O_632,N_14608,N_14588);
and UO_633 (O_633,N_14580,N_14981);
or UO_634 (O_634,N_14485,N_14543);
nand UO_635 (O_635,N_14898,N_14825);
and UO_636 (O_636,N_14325,N_14848);
xor UO_637 (O_637,N_14545,N_14972);
and UO_638 (O_638,N_14457,N_14745);
nand UO_639 (O_639,N_14773,N_14753);
or UO_640 (O_640,N_14476,N_14943);
or UO_641 (O_641,N_14880,N_14577);
and UO_642 (O_642,N_14354,N_14578);
nor UO_643 (O_643,N_14467,N_14741);
or UO_644 (O_644,N_14899,N_14824);
and UO_645 (O_645,N_14792,N_14945);
nand UO_646 (O_646,N_14481,N_14498);
or UO_647 (O_647,N_14593,N_14988);
or UO_648 (O_648,N_14799,N_14421);
nand UO_649 (O_649,N_14332,N_14668);
xnor UO_650 (O_650,N_14744,N_14457);
nand UO_651 (O_651,N_14354,N_14332);
nor UO_652 (O_652,N_14439,N_14931);
and UO_653 (O_653,N_14329,N_14699);
nor UO_654 (O_654,N_14583,N_14404);
nand UO_655 (O_655,N_14896,N_14327);
or UO_656 (O_656,N_14252,N_14745);
xnor UO_657 (O_657,N_14683,N_14308);
and UO_658 (O_658,N_14788,N_14901);
or UO_659 (O_659,N_14554,N_14759);
xnor UO_660 (O_660,N_14549,N_14856);
or UO_661 (O_661,N_14690,N_14598);
xor UO_662 (O_662,N_14262,N_14905);
and UO_663 (O_663,N_14719,N_14733);
nand UO_664 (O_664,N_14977,N_14330);
xor UO_665 (O_665,N_14779,N_14903);
nand UO_666 (O_666,N_14386,N_14925);
and UO_667 (O_667,N_14542,N_14899);
and UO_668 (O_668,N_14711,N_14815);
and UO_669 (O_669,N_14738,N_14779);
or UO_670 (O_670,N_14691,N_14872);
nand UO_671 (O_671,N_14826,N_14994);
nand UO_672 (O_672,N_14745,N_14294);
xnor UO_673 (O_673,N_14497,N_14651);
or UO_674 (O_674,N_14782,N_14649);
nor UO_675 (O_675,N_14925,N_14756);
and UO_676 (O_676,N_14481,N_14936);
nand UO_677 (O_677,N_14881,N_14458);
or UO_678 (O_678,N_14796,N_14883);
nand UO_679 (O_679,N_14617,N_14554);
nand UO_680 (O_680,N_14917,N_14373);
nor UO_681 (O_681,N_14578,N_14604);
xor UO_682 (O_682,N_14882,N_14878);
and UO_683 (O_683,N_14616,N_14849);
nor UO_684 (O_684,N_14580,N_14672);
xnor UO_685 (O_685,N_14382,N_14527);
xor UO_686 (O_686,N_14816,N_14634);
nand UO_687 (O_687,N_14467,N_14393);
nor UO_688 (O_688,N_14300,N_14692);
nor UO_689 (O_689,N_14457,N_14969);
or UO_690 (O_690,N_14582,N_14895);
xor UO_691 (O_691,N_14447,N_14697);
and UO_692 (O_692,N_14540,N_14293);
xor UO_693 (O_693,N_14789,N_14820);
nor UO_694 (O_694,N_14407,N_14896);
nand UO_695 (O_695,N_14491,N_14422);
or UO_696 (O_696,N_14648,N_14888);
xnor UO_697 (O_697,N_14956,N_14506);
xor UO_698 (O_698,N_14984,N_14785);
nor UO_699 (O_699,N_14965,N_14753);
and UO_700 (O_700,N_14535,N_14677);
nor UO_701 (O_701,N_14518,N_14845);
nor UO_702 (O_702,N_14735,N_14560);
and UO_703 (O_703,N_14599,N_14880);
nand UO_704 (O_704,N_14259,N_14250);
and UO_705 (O_705,N_14675,N_14667);
and UO_706 (O_706,N_14309,N_14800);
or UO_707 (O_707,N_14858,N_14632);
and UO_708 (O_708,N_14613,N_14576);
nor UO_709 (O_709,N_14374,N_14694);
nor UO_710 (O_710,N_14415,N_14428);
xor UO_711 (O_711,N_14480,N_14298);
nand UO_712 (O_712,N_14783,N_14559);
and UO_713 (O_713,N_14944,N_14362);
nor UO_714 (O_714,N_14708,N_14484);
nand UO_715 (O_715,N_14855,N_14760);
nor UO_716 (O_716,N_14863,N_14979);
nor UO_717 (O_717,N_14461,N_14868);
or UO_718 (O_718,N_14996,N_14743);
and UO_719 (O_719,N_14746,N_14884);
nand UO_720 (O_720,N_14834,N_14698);
and UO_721 (O_721,N_14425,N_14852);
nor UO_722 (O_722,N_14256,N_14666);
nand UO_723 (O_723,N_14444,N_14298);
nand UO_724 (O_724,N_14379,N_14562);
or UO_725 (O_725,N_14259,N_14991);
xor UO_726 (O_726,N_14683,N_14908);
and UO_727 (O_727,N_14302,N_14437);
nand UO_728 (O_728,N_14854,N_14395);
nor UO_729 (O_729,N_14951,N_14364);
or UO_730 (O_730,N_14492,N_14998);
and UO_731 (O_731,N_14396,N_14495);
or UO_732 (O_732,N_14370,N_14930);
nand UO_733 (O_733,N_14596,N_14411);
xnor UO_734 (O_734,N_14372,N_14383);
and UO_735 (O_735,N_14406,N_14823);
nor UO_736 (O_736,N_14501,N_14460);
or UO_737 (O_737,N_14419,N_14550);
nor UO_738 (O_738,N_14435,N_14941);
and UO_739 (O_739,N_14474,N_14525);
xor UO_740 (O_740,N_14556,N_14428);
nor UO_741 (O_741,N_14537,N_14519);
nand UO_742 (O_742,N_14638,N_14830);
nor UO_743 (O_743,N_14827,N_14347);
nand UO_744 (O_744,N_14762,N_14865);
or UO_745 (O_745,N_14349,N_14983);
nor UO_746 (O_746,N_14931,N_14489);
or UO_747 (O_747,N_14400,N_14670);
and UO_748 (O_748,N_14919,N_14461);
or UO_749 (O_749,N_14974,N_14574);
nand UO_750 (O_750,N_14358,N_14321);
and UO_751 (O_751,N_14934,N_14426);
or UO_752 (O_752,N_14388,N_14784);
or UO_753 (O_753,N_14864,N_14607);
and UO_754 (O_754,N_14907,N_14455);
or UO_755 (O_755,N_14480,N_14834);
nor UO_756 (O_756,N_14293,N_14415);
nand UO_757 (O_757,N_14973,N_14283);
and UO_758 (O_758,N_14286,N_14275);
nor UO_759 (O_759,N_14451,N_14368);
xnor UO_760 (O_760,N_14990,N_14587);
or UO_761 (O_761,N_14932,N_14924);
nor UO_762 (O_762,N_14933,N_14538);
nand UO_763 (O_763,N_14382,N_14543);
and UO_764 (O_764,N_14310,N_14573);
xnor UO_765 (O_765,N_14929,N_14570);
nand UO_766 (O_766,N_14998,N_14683);
xnor UO_767 (O_767,N_14723,N_14607);
nand UO_768 (O_768,N_14987,N_14629);
or UO_769 (O_769,N_14596,N_14625);
and UO_770 (O_770,N_14656,N_14614);
or UO_771 (O_771,N_14402,N_14854);
nor UO_772 (O_772,N_14323,N_14491);
nor UO_773 (O_773,N_14606,N_14839);
or UO_774 (O_774,N_14935,N_14771);
or UO_775 (O_775,N_14518,N_14794);
nor UO_776 (O_776,N_14507,N_14261);
nor UO_777 (O_777,N_14555,N_14683);
nand UO_778 (O_778,N_14390,N_14336);
nand UO_779 (O_779,N_14990,N_14740);
and UO_780 (O_780,N_14280,N_14272);
xor UO_781 (O_781,N_14533,N_14732);
or UO_782 (O_782,N_14632,N_14274);
nand UO_783 (O_783,N_14503,N_14702);
or UO_784 (O_784,N_14254,N_14466);
and UO_785 (O_785,N_14445,N_14418);
xnor UO_786 (O_786,N_14758,N_14345);
xor UO_787 (O_787,N_14562,N_14255);
and UO_788 (O_788,N_14368,N_14756);
nand UO_789 (O_789,N_14397,N_14865);
nor UO_790 (O_790,N_14264,N_14767);
and UO_791 (O_791,N_14487,N_14292);
or UO_792 (O_792,N_14966,N_14983);
nor UO_793 (O_793,N_14313,N_14552);
nand UO_794 (O_794,N_14586,N_14877);
nor UO_795 (O_795,N_14744,N_14556);
and UO_796 (O_796,N_14530,N_14500);
and UO_797 (O_797,N_14934,N_14902);
and UO_798 (O_798,N_14314,N_14929);
nor UO_799 (O_799,N_14501,N_14592);
and UO_800 (O_800,N_14693,N_14981);
and UO_801 (O_801,N_14705,N_14293);
and UO_802 (O_802,N_14304,N_14512);
or UO_803 (O_803,N_14572,N_14513);
and UO_804 (O_804,N_14656,N_14675);
nor UO_805 (O_805,N_14957,N_14911);
nand UO_806 (O_806,N_14666,N_14946);
and UO_807 (O_807,N_14709,N_14648);
or UO_808 (O_808,N_14984,N_14756);
or UO_809 (O_809,N_14824,N_14404);
nand UO_810 (O_810,N_14288,N_14873);
nor UO_811 (O_811,N_14472,N_14537);
and UO_812 (O_812,N_14587,N_14595);
nor UO_813 (O_813,N_14287,N_14678);
and UO_814 (O_814,N_14539,N_14810);
nor UO_815 (O_815,N_14636,N_14714);
or UO_816 (O_816,N_14913,N_14306);
xor UO_817 (O_817,N_14976,N_14590);
and UO_818 (O_818,N_14338,N_14470);
and UO_819 (O_819,N_14529,N_14652);
and UO_820 (O_820,N_14784,N_14771);
nand UO_821 (O_821,N_14556,N_14846);
nor UO_822 (O_822,N_14259,N_14886);
and UO_823 (O_823,N_14485,N_14857);
nor UO_824 (O_824,N_14985,N_14253);
nor UO_825 (O_825,N_14583,N_14716);
nor UO_826 (O_826,N_14620,N_14374);
or UO_827 (O_827,N_14283,N_14414);
nor UO_828 (O_828,N_14291,N_14301);
nor UO_829 (O_829,N_14679,N_14592);
nand UO_830 (O_830,N_14467,N_14420);
or UO_831 (O_831,N_14446,N_14715);
nand UO_832 (O_832,N_14559,N_14617);
nand UO_833 (O_833,N_14335,N_14956);
nor UO_834 (O_834,N_14353,N_14354);
and UO_835 (O_835,N_14959,N_14952);
and UO_836 (O_836,N_14412,N_14473);
nand UO_837 (O_837,N_14626,N_14803);
nor UO_838 (O_838,N_14600,N_14749);
nand UO_839 (O_839,N_14308,N_14617);
or UO_840 (O_840,N_14832,N_14639);
and UO_841 (O_841,N_14654,N_14683);
nor UO_842 (O_842,N_14551,N_14654);
and UO_843 (O_843,N_14708,N_14920);
and UO_844 (O_844,N_14646,N_14315);
nand UO_845 (O_845,N_14415,N_14916);
nor UO_846 (O_846,N_14581,N_14371);
xor UO_847 (O_847,N_14444,N_14628);
nand UO_848 (O_848,N_14827,N_14636);
nand UO_849 (O_849,N_14454,N_14436);
and UO_850 (O_850,N_14924,N_14630);
and UO_851 (O_851,N_14425,N_14475);
and UO_852 (O_852,N_14416,N_14727);
and UO_853 (O_853,N_14607,N_14305);
or UO_854 (O_854,N_14970,N_14603);
and UO_855 (O_855,N_14912,N_14543);
nand UO_856 (O_856,N_14501,N_14678);
xor UO_857 (O_857,N_14367,N_14420);
or UO_858 (O_858,N_14389,N_14282);
nand UO_859 (O_859,N_14372,N_14251);
nor UO_860 (O_860,N_14836,N_14921);
and UO_861 (O_861,N_14719,N_14831);
nor UO_862 (O_862,N_14658,N_14339);
or UO_863 (O_863,N_14923,N_14443);
and UO_864 (O_864,N_14555,N_14302);
nand UO_865 (O_865,N_14286,N_14661);
nor UO_866 (O_866,N_14963,N_14778);
nor UO_867 (O_867,N_14978,N_14559);
nor UO_868 (O_868,N_14375,N_14765);
and UO_869 (O_869,N_14470,N_14667);
or UO_870 (O_870,N_14919,N_14704);
or UO_871 (O_871,N_14857,N_14917);
and UO_872 (O_872,N_14604,N_14392);
and UO_873 (O_873,N_14970,N_14478);
nor UO_874 (O_874,N_14478,N_14499);
nand UO_875 (O_875,N_14398,N_14892);
nand UO_876 (O_876,N_14872,N_14833);
and UO_877 (O_877,N_14852,N_14897);
nand UO_878 (O_878,N_14849,N_14719);
nor UO_879 (O_879,N_14564,N_14965);
and UO_880 (O_880,N_14642,N_14579);
nor UO_881 (O_881,N_14948,N_14745);
and UO_882 (O_882,N_14866,N_14661);
nand UO_883 (O_883,N_14743,N_14837);
and UO_884 (O_884,N_14480,N_14605);
and UO_885 (O_885,N_14309,N_14695);
xor UO_886 (O_886,N_14860,N_14506);
and UO_887 (O_887,N_14984,N_14594);
nor UO_888 (O_888,N_14609,N_14416);
xor UO_889 (O_889,N_14379,N_14765);
or UO_890 (O_890,N_14462,N_14312);
nor UO_891 (O_891,N_14918,N_14399);
nor UO_892 (O_892,N_14588,N_14931);
and UO_893 (O_893,N_14391,N_14297);
and UO_894 (O_894,N_14468,N_14763);
or UO_895 (O_895,N_14793,N_14774);
or UO_896 (O_896,N_14618,N_14538);
nand UO_897 (O_897,N_14781,N_14443);
nand UO_898 (O_898,N_14363,N_14776);
or UO_899 (O_899,N_14349,N_14980);
nor UO_900 (O_900,N_14342,N_14339);
and UO_901 (O_901,N_14959,N_14508);
or UO_902 (O_902,N_14614,N_14869);
nand UO_903 (O_903,N_14841,N_14856);
nor UO_904 (O_904,N_14367,N_14321);
nand UO_905 (O_905,N_14600,N_14736);
nand UO_906 (O_906,N_14897,N_14371);
or UO_907 (O_907,N_14965,N_14413);
nand UO_908 (O_908,N_14708,N_14736);
nor UO_909 (O_909,N_14391,N_14590);
or UO_910 (O_910,N_14832,N_14476);
or UO_911 (O_911,N_14287,N_14618);
and UO_912 (O_912,N_14875,N_14913);
or UO_913 (O_913,N_14637,N_14456);
or UO_914 (O_914,N_14652,N_14612);
nor UO_915 (O_915,N_14877,N_14812);
and UO_916 (O_916,N_14738,N_14505);
nor UO_917 (O_917,N_14900,N_14642);
and UO_918 (O_918,N_14701,N_14719);
nor UO_919 (O_919,N_14739,N_14857);
nor UO_920 (O_920,N_14722,N_14982);
and UO_921 (O_921,N_14299,N_14999);
nor UO_922 (O_922,N_14641,N_14714);
nand UO_923 (O_923,N_14651,N_14337);
nand UO_924 (O_924,N_14723,N_14737);
or UO_925 (O_925,N_14854,N_14678);
nand UO_926 (O_926,N_14801,N_14705);
and UO_927 (O_927,N_14394,N_14861);
nor UO_928 (O_928,N_14621,N_14939);
nor UO_929 (O_929,N_14363,N_14479);
nand UO_930 (O_930,N_14324,N_14296);
nor UO_931 (O_931,N_14308,N_14822);
or UO_932 (O_932,N_14727,N_14715);
xor UO_933 (O_933,N_14751,N_14745);
nand UO_934 (O_934,N_14570,N_14484);
nand UO_935 (O_935,N_14687,N_14494);
and UO_936 (O_936,N_14720,N_14457);
nand UO_937 (O_937,N_14338,N_14658);
and UO_938 (O_938,N_14454,N_14359);
or UO_939 (O_939,N_14484,N_14873);
and UO_940 (O_940,N_14486,N_14847);
nand UO_941 (O_941,N_14423,N_14483);
and UO_942 (O_942,N_14749,N_14492);
nand UO_943 (O_943,N_14834,N_14393);
xor UO_944 (O_944,N_14292,N_14490);
and UO_945 (O_945,N_14375,N_14638);
or UO_946 (O_946,N_14868,N_14946);
or UO_947 (O_947,N_14837,N_14797);
nor UO_948 (O_948,N_14577,N_14719);
and UO_949 (O_949,N_14591,N_14669);
nand UO_950 (O_950,N_14578,N_14663);
or UO_951 (O_951,N_14896,N_14544);
and UO_952 (O_952,N_14363,N_14804);
xnor UO_953 (O_953,N_14634,N_14283);
nand UO_954 (O_954,N_14398,N_14862);
or UO_955 (O_955,N_14770,N_14428);
xnor UO_956 (O_956,N_14590,N_14294);
nor UO_957 (O_957,N_14823,N_14816);
xnor UO_958 (O_958,N_14932,N_14621);
or UO_959 (O_959,N_14340,N_14578);
and UO_960 (O_960,N_14684,N_14603);
nor UO_961 (O_961,N_14683,N_14311);
nor UO_962 (O_962,N_14260,N_14773);
nand UO_963 (O_963,N_14311,N_14766);
xor UO_964 (O_964,N_14573,N_14365);
nor UO_965 (O_965,N_14288,N_14748);
and UO_966 (O_966,N_14342,N_14871);
xnor UO_967 (O_967,N_14531,N_14689);
xor UO_968 (O_968,N_14394,N_14401);
and UO_969 (O_969,N_14410,N_14445);
and UO_970 (O_970,N_14342,N_14425);
xor UO_971 (O_971,N_14322,N_14576);
or UO_972 (O_972,N_14443,N_14949);
nor UO_973 (O_973,N_14490,N_14448);
nor UO_974 (O_974,N_14871,N_14976);
nand UO_975 (O_975,N_14470,N_14411);
xor UO_976 (O_976,N_14337,N_14267);
nand UO_977 (O_977,N_14312,N_14771);
and UO_978 (O_978,N_14726,N_14598);
or UO_979 (O_979,N_14951,N_14644);
and UO_980 (O_980,N_14881,N_14820);
xor UO_981 (O_981,N_14899,N_14801);
and UO_982 (O_982,N_14459,N_14331);
xor UO_983 (O_983,N_14811,N_14876);
nor UO_984 (O_984,N_14660,N_14348);
nand UO_985 (O_985,N_14387,N_14301);
nand UO_986 (O_986,N_14572,N_14961);
or UO_987 (O_987,N_14512,N_14268);
and UO_988 (O_988,N_14931,N_14256);
or UO_989 (O_989,N_14382,N_14447);
or UO_990 (O_990,N_14513,N_14755);
or UO_991 (O_991,N_14721,N_14354);
and UO_992 (O_992,N_14371,N_14799);
or UO_993 (O_993,N_14715,N_14726);
or UO_994 (O_994,N_14689,N_14874);
nand UO_995 (O_995,N_14449,N_14728);
or UO_996 (O_996,N_14976,N_14478);
nor UO_997 (O_997,N_14505,N_14478);
nand UO_998 (O_998,N_14559,N_14483);
nor UO_999 (O_999,N_14669,N_14705);
nor UO_1000 (O_1000,N_14982,N_14693);
nand UO_1001 (O_1001,N_14695,N_14506);
nor UO_1002 (O_1002,N_14960,N_14288);
nor UO_1003 (O_1003,N_14885,N_14415);
nand UO_1004 (O_1004,N_14389,N_14637);
or UO_1005 (O_1005,N_14425,N_14507);
xnor UO_1006 (O_1006,N_14536,N_14339);
xnor UO_1007 (O_1007,N_14957,N_14774);
and UO_1008 (O_1008,N_14652,N_14716);
xnor UO_1009 (O_1009,N_14603,N_14770);
and UO_1010 (O_1010,N_14299,N_14665);
nor UO_1011 (O_1011,N_14871,N_14490);
nand UO_1012 (O_1012,N_14718,N_14808);
or UO_1013 (O_1013,N_14443,N_14627);
or UO_1014 (O_1014,N_14775,N_14520);
and UO_1015 (O_1015,N_14627,N_14288);
nand UO_1016 (O_1016,N_14747,N_14605);
nand UO_1017 (O_1017,N_14670,N_14447);
and UO_1018 (O_1018,N_14515,N_14335);
xor UO_1019 (O_1019,N_14454,N_14937);
and UO_1020 (O_1020,N_14352,N_14453);
nor UO_1021 (O_1021,N_14620,N_14709);
and UO_1022 (O_1022,N_14338,N_14962);
and UO_1023 (O_1023,N_14930,N_14384);
nand UO_1024 (O_1024,N_14864,N_14994);
and UO_1025 (O_1025,N_14347,N_14524);
or UO_1026 (O_1026,N_14938,N_14571);
nand UO_1027 (O_1027,N_14581,N_14850);
xor UO_1028 (O_1028,N_14744,N_14508);
nor UO_1029 (O_1029,N_14851,N_14533);
or UO_1030 (O_1030,N_14686,N_14257);
or UO_1031 (O_1031,N_14556,N_14899);
nor UO_1032 (O_1032,N_14566,N_14380);
nand UO_1033 (O_1033,N_14792,N_14658);
nor UO_1034 (O_1034,N_14619,N_14292);
nand UO_1035 (O_1035,N_14720,N_14476);
or UO_1036 (O_1036,N_14780,N_14581);
and UO_1037 (O_1037,N_14447,N_14283);
or UO_1038 (O_1038,N_14438,N_14400);
and UO_1039 (O_1039,N_14575,N_14847);
nand UO_1040 (O_1040,N_14757,N_14996);
or UO_1041 (O_1041,N_14350,N_14604);
nand UO_1042 (O_1042,N_14936,N_14795);
nand UO_1043 (O_1043,N_14313,N_14989);
nor UO_1044 (O_1044,N_14932,N_14678);
and UO_1045 (O_1045,N_14803,N_14906);
and UO_1046 (O_1046,N_14500,N_14291);
xnor UO_1047 (O_1047,N_14503,N_14523);
or UO_1048 (O_1048,N_14786,N_14340);
nand UO_1049 (O_1049,N_14856,N_14941);
nor UO_1050 (O_1050,N_14958,N_14394);
nor UO_1051 (O_1051,N_14383,N_14699);
xor UO_1052 (O_1052,N_14643,N_14298);
nand UO_1053 (O_1053,N_14902,N_14973);
xor UO_1054 (O_1054,N_14841,N_14568);
xnor UO_1055 (O_1055,N_14818,N_14385);
and UO_1056 (O_1056,N_14418,N_14658);
and UO_1057 (O_1057,N_14731,N_14915);
nand UO_1058 (O_1058,N_14674,N_14900);
or UO_1059 (O_1059,N_14346,N_14261);
xnor UO_1060 (O_1060,N_14869,N_14367);
or UO_1061 (O_1061,N_14610,N_14791);
nor UO_1062 (O_1062,N_14621,N_14411);
and UO_1063 (O_1063,N_14964,N_14903);
nand UO_1064 (O_1064,N_14465,N_14406);
nor UO_1065 (O_1065,N_14826,N_14846);
and UO_1066 (O_1066,N_14816,N_14444);
or UO_1067 (O_1067,N_14658,N_14344);
and UO_1068 (O_1068,N_14939,N_14844);
and UO_1069 (O_1069,N_14705,N_14898);
nor UO_1070 (O_1070,N_14474,N_14584);
nor UO_1071 (O_1071,N_14435,N_14279);
nor UO_1072 (O_1072,N_14925,N_14656);
or UO_1073 (O_1073,N_14568,N_14294);
and UO_1074 (O_1074,N_14596,N_14725);
and UO_1075 (O_1075,N_14493,N_14406);
or UO_1076 (O_1076,N_14738,N_14474);
nand UO_1077 (O_1077,N_14999,N_14797);
nor UO_1078 (O_1078,N_14923,N_14901);
or UO_1079 (O_1079,N_14659,N_14442);
nor UO_1080 (O_1080,N_14732,N_14899);
and UO_1081 (O_1081,N_14636,N_14923);
or UO_1082 (O_1082,N_14409,N_14879);
nand UO_1083 (O_1083,N_14361,N_14846);
nand UO_1084 (O_1084,N_14269,N_14690);
nor UO_1085 (O_1085,N_14932,N_14712);
nand UO_1086 (O_1086,N_14906,N_14887);
nand UO_1087 (O_1087,N_14436,N_14690);
and UO_1088 (O_1088,N_14394,N_14680);
nor UO_1089 (O_1089,N_14955,N_14415);
nor UO_1090 (O_1090,N_14384,N_14904);
and UO_1091 (O_1091,N_14634,N_14800);
or UO_1092 (O_1092,N_14741,N_14492);
nand UO_1093 (O_1093,N_14408,N_14950);
nor UO_1094 (O_1094,N_14436,N_14481);
nor UO_1095 (O_1095,N_14845,N_14315);
and UO_1096 (O_1096,N_14883,N_14630);
xor UO_1097 (O_1097,N_14421,N_14951);
nor UO_1098 (O_1098,N_14782,N_14374);
nand UO_1099 (O_1099,N_14687,N_14528);
nor UO_1100 (O_1100,N_14773,N_14840);
nor UO_1101 (O_1101,N_14765,N_14351);
and UO_1102 (O_1102,N_14889,N_14865);
or UO_1103 (O_1103,N_14932,N_14545);
nor UO_1104 (O_1104,N_14327,N_14967);
nor UO_1105 (O_1105,N_14333,N_14555);
or UO_1106 (O_1106,N_14295,N_14798);
nor UO_1107 (O_1107,N_14260,N_14533);
nand UO_1108 (O_1108,N_14320,N_14485);
nand UO_1109 (O_1109,N_14718,N_14835);
or UO_1110 (O_1110,N_14814,N_14779);
nor UO_1111 (O_1111,N_14780,N_14910);
or UO_1112 (O_1112,N_14316,N_14841);
nand UO_1113 (O_1113,N_14495,N_14298);
or UO_1114 (O_1114,N_14250,N_14424);
or UO_1115 (O_1115,N_14339,N_14345);
nand UO_1116 (O_1116,N_14296,N_14492);
and UO_1117 (O_1117,N_14678,N_14690);
nand UO_1118 (O_1118,N_14357,N_14773);
nand UO_1119 (O_1119,N_14790,N_14484);
or UO_1120 (O_1120,N_14377,N_14920);
nor UO_1121 (O_1121,N_14990,N_14367);
and UO_1122 (O_1122,N_14772,N_14758);
nand UO_1123 (O_1123,N_14878,N_14301);
and UO_1124 (O_1124,N_14405,N_14347);
nor UO_1125 (O_1125,N_14835,N_14911);
nor UO_1126 (O_1126,N_14534,N_14621);
nand UO_1127 (O_1127,N_14650,N_14417);
or UO_1128 (O_1128,N_14946,N_14965);
or UO_1129 (O_1129,N_14942,N_14302);
xnor UO_1130 (O_1130,N_14268,N_14440);
nor UO_1131 (O_1131,N_14978,N_14641);
xnor UO_1132 (O_1132,N_14388,N_14656);
or UO_1133 (O_1133,N_14593,N_14794);
nor UO_1134 (O_1134,N_14250,N_14675);
and UO_1135 (O_1135,N_14297,N_14834);
nand UO_1136 (O_1136,N_14256,N_14941);
and UO_1137 (O_1137,N_14436,N_14748);
or UO_1138 (O_1138,N_14621,N_14460);
nor UO_1139 (O_1139,N_14456,N_14517);
nand UO_1140 (O_1140,N_14362,N_14515);
nor UO_1141 (O_1141,N_14392,N_14395);
xnor UO_1142 (O_1142,N_14650,N_14541);
and UO_1143 (O_1143,N_14948,N_14525);
and UO_1144 (O_1144,N_14448,N_14441);
or UO_1145 (O_1145,N_14258,N_14775);
nand UO_1146 (O_1146,N_14865,N_14377);
xnor UO_1147 (O_1147,N_14392,N_14616);
xor UO_1148 (O_1148,N_14529,N_14940);
and UO_1149 (O_1149,N_14931,N_14982);
xor UO_1150 (O_1150,N_14732,N_14755);
and UO_1151 (O_1151,N_14583,N_14975);
and UO_1152 (O_1152,N_14898,N_14683);
and UO_1153 (O_1153,N_14781,N_14673);
nand UO_1154 (O_1154,N_14648,N_14858);
nand UO_1155 (O_1155,N_14899,N_14655);
and UO_1156 (O_1156,N_14398,N_14363);
and UO_1157 (O_1157,N_14525,N_14854);
or UO_1158 (O_1158,N_14828,N_14913);
and UO_1159 (O_1159,N_14606,N_14501);
xor UO_1160 (O_1160,N_14791,N_14662);
xor UO_1161 (O_1161,N_14754,N_14338);
nand UO_1162 (O_1162,N_14323,N_14759);
or UO_1163 (O_1163,N_14384,N_14873);
or UO_1164 (O_1164,N_14371,N_14438);
nor UO_1165 (O_1165,N_14768,N_14595);
nor UO_1166 (O_1166,N_14379,N_14302);
nor UO_1167 (O_1167,N_14361,N_14615);
or UO_1168 (O_1168,N_14577,N_14587);
nand UO_1169 (O_1169,N_14831,N_14391);
xor UO_1170 (O_1170,N_14318,N_14321);
and UO_1171 (O_1171,N_14778,N_14511);
or UO_1172 (O_1172,N_14481,N_14953);
or UO_1173 (O_1173,N_14785,N_14445);
nor UO_1174 (O_1174,N_14490,N_14829);
and UO_1175 (O_1175,N_14771,N_14371);
nand UO_1176 (O_1176,N_14489,N_14621);
nand UO_1177 (O_1177,N_14441,N_14522);
nor UO_1178 (O_1178,N_14337,N_14881);
nor UO_1179 (O_1179,N_14267,N_14701);
or UO_1180 (O_1180,N_14525,N_14528);
and UO_1181 (O_1181,N_14583,N_14688);
nor UO_1182 (O_1182,N_14309,N_14887);
nand UO_1183 (O_1183,N_14383,N_14762);
or UO_1184 (O_1184,N_14281,N_14714);
or UO_1185 (O_1185,N_14593,N_14411);
xor UO_1186 (O_1186,N_14538,N_14963);
nor UO_1187 (O_1187,N_14259,N_14799);
or UO_1188 (O_1188,N_14553,N_14958);
or UO_1189 (O_1189,N_14963,N_14260);
nand UO_1190 (O_1190,N_14975,N_14314);
nor UO_1191 (O_1191,N_14895,N_14731);
nor UO_1192 (O_1192,N_14498,N_14514);
or UO_1193 (O_1193,N_14795,N_14959);
or UO_1194 (O_1194,N_14400,N_14493);
and UO_1195 (O_1195,N_14959,N_14307);
nand UO_1196 (O_1196,N_14793,N_14382);
nand UO_1197 (O_1197,N_14933,N_14287);
xor UO_1198 (O_1198,N_14840,N_14459);
and UO_1199 (O_1199,N_14781,N_14999);
nand UO_1200 (O_1200,N_14339,N_14582);
or UO_1201 (O_1201,N_14896,N_14648);
xnor UO_1202 (O_1202,N_14982,N_14290);
or UO_1203 (O_1203,N_14642,N_14791);
nand UO_1204 (O_1204,N_14380,N_14541);
or UO_1205 (O_1205,N_14766,N_14511);
nand UO_1206 (O_1206,N_14571,N_14782);
xor UO_1207 (O_1207,N_14525,N_14840);
nor UO_1208 (O_1208,N_14747,N_14349);
nor UO_1209 (O_1209,N_14796,N_14288);
nand UO_1210 (O_1210,N_14872,N_14803);
nor UO_1211 (O_1211,N_14860,N_14805);
and UO_1212 (O_1212,N_14466,N_14552);
nor UO_1213 (O_1213,N_14369,N_14711);
nor UO_1214 (O_1214,N_14948,N_14501);
nor UO_1215 (O_1215,N_14250,N_14271);
xnor UO_1216 (O_1216,N_14965,N_14615);
nor UO_1217 (O_1217,N_14878,N_14655);
nand UO_1218 (O_1218,N_14652,N_14373);
nor UO_1219 (O_1219,N_14700,N_14573);
xnor UO_1220 (O_1220,N_14994,N_14469);
nor UO_1221 (O_1221,N_14391,N_14439);
xor UO_1222 (O_1222,N_14636,N_14926);
nand UO_1223 (O_1223,N_14562,N_14523);
nand UO_1224 (O_1224,N_14265,N_14400);
nor UO_1225 (O_1225,N_14764,N_14837);
nor UO_1226 (O_1226,N_14427,N_14911);
or UO_1227 (O_1227,N_14352,N_14685);
and UO_1228 (O_1228,N_14420,N_14488);
nor UO_1229 (O_1229,N_14275,N_14958);
and UO_1230 (O_1230,N_14469,N_14674);
nand UO_1231 (O_1231,N_14858,N_14661);
nor UO_1232 (O_1232,N_14313,N_14309);
nand UO_1233 (O_1233,N_14275,N_14579);
or UO_1234 (O_1234,N_14855,N_14259);
nor UO_1235 (O_1235,N_14656,N_14931);
nor UO_1236 (O_1236,N_14332,N_14509);
nand UO_1237 (O_1237,N_14822,N_14492);
nand UO_1238 (O_1238,N_14959,N_14386);
nor UO_1239 (O_1239,N_14342,N_14663);
nand UO_1240 (O_1240,N_14607,N_14731);
and UO_1241 (O_1241,N_14345,N_14464);
nor UO_1242 (O_1242,N_14396,N_14619);
and UO_1243 (O_1243,N_14831,N_14325);
nand UO_1244 (O_1244,N_14934,N_14705);
or UO_1245 (O_1245,N_14670,N_14251);
nor UO_1246 (O_1246,N_14653,N_14755);
or UO_1247 (O_1247,N_14923,N_14696);
or UO_1248 (O_1248,N_14654,N_14512);
nor UO_1249 (O_1249,N_14259,N_14473);
nand UO_1250 (O_1250,N_14909,N_14590);
nor UO_1251 (O_1251,N_14355,N_14346);
nand UO_1252 (O_1252,N_14480,N_14821);
or UO_1253 (O_1253,N_14315,N_14919);
nand UO_1254 (O_1254,N_14543,N_14774);
nor UO_1255 (O_1255,N_14767,N_14701);
xnor UO_1256 (O_1256,N_14936,N_14589);
or UO_1257 (O_1257,N_14825,N_14651);
nor UO_1258 (O_1258,N_14363,N_14995);
and UO_1259 (O_1259,N_14639,N_14743);
nor UO_1260 (O_1260,N_14473,N_14374);
or UO_1261 (O_1261,N_14518,N_14281);
xnor UO_1262 (O_1262,N_14793,N_14826);
and UO_1263 (O_1263,N_14623,N_14352);
xor UO_1264 (O_1264,N_14992,N_14347);
and UO_1265 (O_1265,N_14682,N_14687);
or UO_1266 (O_1266,N_14523,N_14722);
and UO_1267 (O_1267,N_14371,N_14807);
xnor UO_1268 (O_1268,N_14480,N_14906);
nor UO_1269 (O_1269,N_14308,N_14573);
and UO_1270 (O_1270,N_14999,N_14829);
or UO_1271 (O_1271,N_14958,N_14806);
and UO_1272 (O_1272,N_14886,N_14305);
nor UO_1273 (O_1273,N_14825,N_14289);
and UO_1274 (O_1274,N_14433,N_14639);
and UO_1275 (O_1275,N_14601,N_14886);
and UO_1276 (O_1276,N_14709,N_14513);
or UO_1277 (O_1277,N_14778,N_14264);
nor UO_1278 (O_1278,N_14602,N_14617);
and UO_1279 (O_1279,N_14654,N_14391);
and UO_1280 (O_1280,N_14657,N_14877);
nor UO_1281 (O_1281,N_14633,N_14991);
nand UO_1282 (O_1282,N_14550,N_14998);
or UO_1283 (O_1283,N_14296,N_14458);
and UO_1284 (O_1284,N_14489,N_14689);
nand UO_1285 (O_1285,N_14992,N_14321);
or UO_1286 (O_1286,N_14951,N_14978);
nand UO_1287 (O_1287,N_14734,N_14439);
nor UO_1288 (O_1288,N_14584,N_14856);
nand UO_1289 (O_1289,N_14954,N_14879);
and UO_1290 (O_1290,N_14703,N_14636);
nand UO_1291 (O_1291,N_14510,N_14860);
nor UO_1292 (O_1292,N_14988,N_14255);
xor UO_1293 (O_1293,N_14369,N_14646);
or UO_1294 (O_1294,N_14363,N_14719);
xnor UO_1295 (O_1295,N_14986,N_14750);
nor UO_1296 (O_1296,N_14769,N_14850);
nand UO_1297 (O_1297,N_14927,N_14683);
and UO_1298 (O_1298,N_14829,N_14538);
and UO_1299 (O_1299,N_14541,N_14324);
nor UO_1300 (O_1300,N_14465,N_14532);
nor UO_1301 (O_1301,N_14925,N_14433);
and UO_1302 (O_1302,N_14396,N_14400);
or UO_1303 (O_1303,N_14907,N_14563);
or UO_1304 (O_1304,N_14527,N_14394);
nand UO_1305 (O_1305,N_14814,N_14687);
and UO_1306 (O_1306,N_14307,N_14605);
nor UO_1307 (O_1307,N_14530,N_14750);
nand UO_1308 (O_1308,N_14317,N_14314);
and UO_1309 (O_1309,N_14698,N_14460);
nand UO_1310 (O_1310,N_14808,N_14842);
nor UO_1311 (O_1311,N_14587,N_14727);
or UO_1312 (O_1312,N_14426,N_14900);
and UO_1313 (O_1313,N_14832,N_14655);
and UO_1314 (O_1314,N_14332,N_14381);
nand UO_1315 (O_1315,N_14723,N_14514);
nor UO_1316 (O_1316,N_14952,N_14970);
or UO_1317 (O_1317,N_14915,N_14552);
nor UO_1318 (O_1318,N_14885,N_14875);
or UO_1319 (O_1319,N_14789,N_14279);
or UO_1320 (O_1320,N_14844,N_14623);
nor UO_1321 (O_1321,N_14858,N_14468);
nand UO_1322 (O_1322,N_14888,N_14495);
and UO_1323 (O_1323,N_14454,N_14642);
nand UO_1324 (O_1324,N_14628,N_14870);
nor UO_1325 (O_1325,N_14679,N_14647);
nand UO_1326 (O_1326,N_14619,N_14938);
nor UO_1327 (O_1327,N_14496,N_14358);
and UO_1328 (O_1328,N_14632,N_14901);
or UO_1329 (O_1329,N_14402,N_14397);
and UO_1330 (O_1330,N_14400,N_14662);
nor UO_1331 (O_1331,N_14782,N_14345);
nor UO_1332 (O_1332,N_14486,N_14363);
xor UO_1333 (O_1333,N_14327,N_14695);
nand UO_1334 (O_1334,N_14798,N_14576);
nor UO_1335 (O_1335,N_14441,N_14982);
and UO_1336 (O_1336,N_14908,N_14898);
and UO_1337 (O_1337,N_14890,N_14531);
and UO_1338 (O_1338,N_14282,N_14729);
xor UO_1339 (O_1339,N_14435,N_14772);
and UO_1340 (O_1340,N_14284,N_14761);
nand UO_1341 (O_1341,N_14784,N_14606);
and UO_1342 (O_1342,N_14969,N_14601);
nand UO_1343 (O_1343,N_14363,N_14556);
nor UO_1344 (O_1344,N_14325,N_14697);
nand UO_1345 (O_1345,N_14555,N_14721);
nand UO_1346 (O_1346,N_14512,N_14835);
nand UO_1347 (O_1347,N_14417,N_14282);
nand UO_1348 (O_1348,N_14865,N_14599);
nor UO_1349 (O_1349,N_14879,N_14881);
or UO_1350 (O_1350,N_14833,N_14530);
nand UO_1351 (O_1351,N_14822,N_14339);
or UO_1352 (O_1352,N_14464,N_14368);
nor UO_1353 (O_1353,N_14873,N_14705);
nor UO_1354 (O_1354,N_14347,N_14757);
xnor UO_1355 (O_1355,N_14287,N_14386);
nor UO_1356 (O_1356,N_14912,N_14496);
and UO_1357 (O_1357,N_14664,N_14983);
nand UO_1358 (O_1358,N_14625,N_14638);
nor UO_1359 (O_1359,N_14540,N_14666);
nor UO_1360 (O_1360,N_14988,N_14418);
nand UO_1361 (O_1361,N_14538,N_14322);
nand UO_1362 (O_1362,N_14262,N_14583);
nor UO_1363 (O_1363,N_14795,N_14285);
or UO_1364 (O_1364,N_14537,N_14424);
nand UO_1365 (O_1365,N_14346,N_14796);
xor UO_1366 (O_1366,N_14985,N_14339);
nor UO_1367 (O_1367,N_14463,N_14451);
nor UO_1368 (O_1368,N_14580,N_14315);
nand UO_1369 (O_1369,N_14801,N_14906);
and UO_1370 (O_1370,N_14661,N_14704);
nand UO_1371 (O_1371,N_14690,N_14584);
or UO_1372 (O_1372,N_14412,N_14909);
or UO_1373 (O_1373,N_14835,N_14529);
or UO_1374 (O_1374,N_14647,N_14566);
nand UO_1375 (O_1375,N_14384,N_14670);
and UO_1376 (O_1376,N_14786,N_14662);
or UO_1377 (O_1377,N_14908,N_14518);
or UO_1378 (O_1378,N_14968,N_14688);
nor UO_1379 (O_1379,N_14334,N_14680);
and UO_1380 (O_1380,N_14287,N_14428);
nand UO_1381 (O_1381,N_14766,N_14267);
xor UO_1382 (O_1382,N_14972,N_14758);
nor UO_1383 (O_1383,N_14390,N_14843);
nor UO_1384 (O_1384,N_14800,N_14835);
nand UO_1385 (O_1385,N_14309,N_14819);
nand UO_1386 (O_1386,N_14788,N_14401);
xor UO_1387 (O_1387,N_14714,N_14347);
or UO_1388 (O_1388,N_14372,N_14431);
xor UO_1389 (O_1389,N_14645,N_14582);
nand UO_1390 (O_1390,N_14628,N_14409);
nor UO_1391 (O_1391,N_14794,N_14668);
nand UO_1392 (O_1392,N_14269,N_14817);
nor UO_1393 (O_1393,N_14850,N_14947);
nor UO_1394 (O_1394,N_14794,N_14257);
nor UO_1395 (O_1395,N_14633,N_14425);
or UO_1396 (O_1396,N_14810,N_14630);
and UO_1397 (O_1397,N_14807,N_14596);
or UO_1398 (O_1398,N_14278,N_14564);
and UO_1399 (O_1399,N_14344,N_14944);
xor UO_1400 (O_1400,N_14342,N_14266);
nand UO_1401 (O_1401,N_14292,N_14716);
nand UO_1402 (O_1402,N_14629,N_14766);
or UO_1403 (O_1403,N_14797,N_14922);
or UO_1404 (O_1404,N_14630,N_14588);
xnor UO_1405 (O_1405,N_14367,N_14815);
or UO_1406 (O_1406,N_14250,N_14684);
xnor UO_1407 (O_1407,N_14971,N_14645);
nand UO_1408 (O_1408,N_14853,N_14532);
and UO_1409 (O_1409,N_14639,N_14432);
nand UO_1410 (O_1410,N_14847,N_14757);
and UO_1411 (O_1411,N_14751,N_14683);
xor UO_1412 (O_1412,N_14329,N_14429);
nor UO_1413 (O_1413,N_14563,N_14298);
xor UO_1414 (O_1414,N_14337,N_14648);
nor UO_1415 (O_1415,N_14434,N_14889);
or UO_1416 (O_1416,N_14301,N_14455);
or UO_1417 (O_1417,N_14559,N_14925);
nand UO_1418 (O_1418,N_14318,N_14456);
nand UO_1419 (O_1419,N_14736,N_14927);
nor UO_1420 (O_1420,N_14424,N_14716);
nand UO_1421 (O_1421,N_14676,N_14649);
nand UO_1422 (O_1422,N_14511,N_14921);
and UO_1423 (O_1423,N_14552,N_14891);
and UO_1424 (O_1424,N_14493,N_14540);
xor UO_1425 (O_1425,N_14298,N_14899);
nor UO_1426 (O_1426,N_14333,N_14297);
or UO_1427 (O_1427,N_14361,N_14280);
or UO_1428 (O_1428,N_14793,N_14885);
xor UO_1429 (O_1429,N_14942,N_14920);
or UO_1430 (O_1430,N_14481,N_14671);
nor UO_1431 (O_1431,N_14377,N_14346);
nor UO_1432 (O_1432,N_14992,N_14286);
and UO_1433 (O_1433,N_14826,N_14448);
nand UO_1434 (O_1434,N_14873,N_14743);
nor UO_1435 (O_1435,N_14584,N_14563);
nor UO_1436 (O_1436,N_14830,N_14409);
nor UO_1437 (O_1437,N_14693,N_14850);
and UO_1438 (O_1438,N_14402,N_14678);
and UO_1439 (O_1439,N_14843,N_14846);
and UO_1440 (O_1440,N_14674,N_14633);
xor UO_1441 (O_1441,N_14729,N_14553);
xnor UO_1442 (O_1442,N_14967,N_14919);
nor UO_1443 (O_1443,N_14547,N_14753);
and UO_1444 (O_1444,N_14507,N_14514);
nor UO_1445 (O_1445,N_14854,N_14386);
or UO_1446 (O_1446,N_14536,N_14445);
nand UO_1447 (O_1447,N_14376,N_14656);
xnor UO_1448 (O_1448,N_14363,N_14275);
or UO_1449 (O_1449,N_14439,N_14657);
nand UO_1450 (O_1450,N_14596,N_14413);
nor UO_1451 (O_1451,N_14347,N_14925);
or UO_1452 (O_1452,N_14746,N_14470);
nor UO_1453 (O_1453,N_14834,N_14455);
or UO_1454 (O_1454,N_14913,N_14767);
nand UO_1455 (O_1455,N_14682,N_14323);
xnor UO_1456 (O_1456,N_14782,N_14640);
nor UO_1457 (O_1457,N_14663,N_14993);
xnor UO_1458 (O_1458,N_14880,N_14625);
xor UO_1459 (O_1459,N_14627,N_14900);
and UO_1460 (O_1460,N_14679,N_14825);
nor UO_1461 (O_1461,N_14688,N_14817);
or UO_1462 (O_1462,N_14692,N_14439);
xor UO_1463 (O_1463,N_14330,N_14311);
or UO_1464 (O_1464,N_14289,N_14995);
or UO_1465 (O_1465,N_14649,N_14314);
xor UO_1466 (O_1466,N_14936,N_14736);
nor UO_1467 (O_1467,N_14772,N_14875);
nor UO_1468 (O_1468,N_14988,N_14506);
xnor UO_1469 (O_1469,N_14736,N_14892);
nor UO_1470 (O_1470,N_14989,N_14378);
nor UO_1471 (O_1471,N_14718,N_14886);
and UO_1472 (O_1472,N_14494,N_14545);
and UO_1473 (O_1473,N_14840,N_14720);
nand UO_1474 (O_1474,N_14867,N_14597);
xnor UO_1475 (O_1475,N_14441,N_14836);
and UO_1476 (O_1476,N_14904,N_14994);
and UO_1477 (O_1477,N_14942,N_14455);
nor UO_1478 (O_1478,N_14742,N_14575);
and UO_1479 (O_1479,N_14385,N_14736);
or UO_1480 (O_1480,N_14902,N_14492);
or UO_1481 (O_1481,N_14780,N_14531);
xor UO_1482 (O_1482,N_14802,N_14953);
nor UO_1483 (O_1483,N_14475,N_14314);
nor UO_1484 (O_1484,N_14312,N_14715);
xnor UO_1485 (O_1485,N_14589,N_14346);
and UO_1486 (O_1486,N_14880,N_14859);
or UO_1487 (O_1487,N_14550,N_14390);
nor UO_1488 (O_1488,N_14973,N_14559);
nand UO_1489 (O_1489,N_14288,N_14905);
and UO_1490 (O_1490,N_14638,N_14572);
and UO_1491 (O_1491,N_14496,N_14973);
nand UO_1492 (O_1492,N_14338,N_14832);
or UO_1493 (O_1493,N_14849,N_14747);
nand UO_1494 (O_1494,N_14954,N_14837);
nand UO_1495 (O_1495,N_14938,N_14805);
nand UO_1496 (O_1496,N_14873,N_14457);
or UO_1497 (O_1497,N_14510,N_14293);
and UO_1498 (O_1498,N_14366,N_14334);
nor UO_1499 (O_1499,N_14320,N_14725);
nor UO_1500 (O_1500,N_14982,N_14739);
or UO_1501 (O_1501,N_14378,N_14284);
and UO_1502 (O_1502,N_14340,N_14326);
xnor UO_1503 (O_1503,N_14730,N_14304);
nor UO_1504 (O_1504,N_14982,N_14351);
or UO_1505 (O_1505,N_14927,N_14980);
or UO_1506 (O_1506,N_14256,N_14285);
and UO_1507 (O_1507,N_14629,N_14472);
nand UO_1508 (O_1508,N_14900,N_14704);
nand UO_1509 (O_1509,N_14530,N_14358);
and UO_1510 (O_1510,N_14280,N_14533);
or UO_1511 (O_1511,N_14932,N_14391);
and UO_1512 (O_1512,N_14911,N_14293);
or UO_1513 (O_1513,N_14624,N_14386);
and UO_1514 (O_1514,N_14627,N_14946);
and UO_1515 (O_1515,N_14553,N_14818);
or UO_1516 (O_1516,N_14679,N_14738);
nor UO_1517 (O_1517,N_14876,N_14520);
xnor UO_1518 (O_1518,N_14367,N_14594);
nand UO_1519 (O_1519,N_14781,N_14940);
nand UO_1520 (O_1520,N_14508,N_14574);
nand UO_1521 (O_1521,N_14511,N_14584);
nand UO_1522 (O_1522,N_14964,N_14677);
nor UO_1523 (O_1523,N_14781,N_14747);
and UO_1524 (O_1524,N_14378,N_14282);
nand UO_1525 (O_1525,N_14285,N_14976);
or UO_1526 (O_1526,N_14755,N_14810);
nand UO_1527 (O_1527,N_14635,N_14998);
nand UO_1528 (O_1528,N_14364,N_14837);
and UO_1529 (O_1529,N_14552,N_14547);
and UO_1530 (O_1530,N_14494,N_14278);
nor UO_1531 (O_1531,N_14278,N_14274);
xor UO_1532 (O_1532,N_14545,N_14662);
and UO_1533 (O_1533,N_14578,N_14284);
nand UO_1534 (O_1534,N_14479,N_14755);
or UO_1535 (O_1535,N_14778,N_14825);
and UO_1536 (O_1536,N_14294,N_14346);
or UO_1537 (O_1537,N_14381,N_14968);
xnor UO_1538 (O_1538,N_14841,N_14874);
and UO_1539 (O_1539,N_14317,N_14582);
or UO_1540 (O_1540,N_14684,N_14894);
and UO_1541 (O_1541,N_14854,N_14655);
nand UO_1542 (O_1542,N_14587,N_14598);
or UO_1543 (O_1543,N_14808,N_14389);
and UO_1544 (O_1544,N_14558,N_14546);
or UO_1545 (O_1545,N_14765,N_14281);
or UO_1546 (O_1546,N_14580,N_14864);
nand UO_1547 (O_1547,N_14557,N_14824);
xnor UO_1548 (O_1548,N_14533,N_14808);
and UO_1549 (O_1549,N_14525,N_14925);
and UO_1550 (O_1550,N_14589,N_14638);
or UO_1551 (O_1551,N_14850,N_14921);
or UO_1552 (O_1552,N_14870,N_14942);
nor UO_1553 (O_1553,N_14496,N_14831);
nand UO_1554 (O_1554,N_14879,N_14461);
nor UO_1555 (O_1555,N_14549,N_14780);
and UO_1556 (O_1556,N_14366,N_14924);
xor UO_1557 (O_1557,N_14353,N_14911);
and UO_1558 (O_1558,N_14693,N_14962);
nand UO_1559 (O_1559,N_14831,N_14877);
or UO_1560 (O_1560,N_14330,N_14705);
nand UO_1561 (O_1561,N_14464,N_14748);
xor UO_1562 (O_1562,N_14570,N_14646);
and UO_1563 (O_1563,N_14588,N_14265);
nand UO_1564 (O_1564,N_14441,N_14540);
and UO_1565 (O_1565,N_14752,N_14878);
and UO_1566 (O_1566,N_14742,N_14609);
nor UO_1567 (O_1567,N_14767,N_14774);
nor UO_1568 (O_1568,N_14977,N_14355);
or UO_1569 (O_1569,N_14811,N_14705);
and UO_1570 (O_1570,N_14444,N_14605);
or UO_1571 (O_1571,N_14622,N_14743);
nand UO_1572 (O_1572,N_14332,N_14385);
or UO_1573 (O_1573,N_14912,N_14505);
or UO_1574 (O_1574,N_14600,N_14368);
or UO_1575 (O_1575,N_14866,N_14423);
nand UO_1576 (O_1576,N_14736,N_14479);
and UO_1577 (O_1577,N_14327,N_14565);
nor UO_1578 (O_1578,N_14990,N_14479);
or UO_1579 (O_1579,N_14407,N_14777);
nand UO_1580 (O_1580,N_14585,N_14473);
or UO_1581 (O_1581,N_14320,N_14690);
nor UO_1582 (O_1582,N_14565,N_14977);
or UO_1583 (O_1583,N_14600,N_14422);
or UO_1584 (O_1584,N_14909,N_14682);
nor UO_1585 (O_1585,N_14751,N_14750);
or UO_1586 (O_1586,N_14976,N_14921);
and UO_1587 (O_1587,N_14589,N_14517);
and UO_1588 (O_1588,N_14815,N_14864);
and UO_1589 (O_1589,N_14429,N_14937);
nand UO_1590 (O_1590,N_14571,N_14474);
and UO_1591 (O_1591,N_14522,N_14405);
nor UO_1592 (O_1592,N_14290,N_14561);
nand UO_1593 (O_1593,N_14577,N_14776);
nor UO_1594 (O_1594,N_14727,N_14687);
nand UO_1595 (O_1595,N_14635,N_14492);
or UO_1596 (O_1596,N_14390,N_14323);
xor UO_1597 (O_1597,N_14886,N_14978);
nor UO_1598 (O_1598,N_14818,N_14878);
or UO_1599 (O_1599,N_14394,N_14279);
and UO_1600 (O_1600,N_14897,N_14329);
xor UO_1601 (O_1601,N_14667,N_14649);
and UO_1602 (O_1602,N_14771,N_14919);
or UO_1603 (O_1603,N_14777,N_14324);
nor UO_1604 (O_1604,N_14728,N_14902);
nand UO_1605 (O_1605,N_14328,N_14536);
xnor UO_1606 (O_1606,N_14590,N_14834);
nor UO_1607 (O_1607,N_14315,N_14851);
or UO_1608 (O_1608,N_14365,N_14856);
nor UO_1609 (O_1609,N_14891,N_14349);
and UO_1610 (O_1610,N_14831,N_14661);
and UO_1611 (O_1611,N_14559,N_14606);
or UO_1612 (O_1612,N_14993,N_14920);
or UO_1613 (O_1613,N_14612,N_14595);
or UO_1614 (O_1614,N_14707,N_14739);
nor UO_1615 (O_1615,N_14623,N_14749);
nand UO_1616 (O_1616,N_14957,N_14581);
and UO_1617 (O_1617,N_14972,N_14712);
nor UO_1618 (O_1618,N_14266,N_14597);
and UO_1619 (O_1619,N_14482,N_14324);
xor UO_1620 (O_1620,N_14805,N_14692);
or UO_1621 (O_1621,N_14922,N_14550);
nor UO_1622 (O_1622,N_14590,N_14891);
or UO_1623 (O_1623,N_14505,N_14670);
xor UO_1624 (O_1624,N_14315,N_14630);
or UO_1625 (O_1625,N_14937,N_14734);
nand UO_1626 (O_1626,N_14442,N_14858);
nor UO_1627 (O_1627,N_14419,N_14401);
nand UO_1628 (O_1628,N_14720,N_14342);
and UO_1629 (O_1629,N_14403,N_14535);
nor UO_1630 (O_1630,N_14629,N_14708);
nor UO_1631 (O_1631,N_14338,N_14545);
nand UO_1632 (O_1632,N_14856,N_14661);
nor UO_1633 (O_1633,N_14987,N_14253);
xnor UO_1634 (O_1634,N_14726,N_14450);
or UO_1635 (O_1635,N_14718,N_14421);
xor UO_1636 (O_1636,N_14265,N_14936);
and UO_1637 (O_1637,N_14531,N_14482);
nor UO_1638 (O_1638,N_14831,N_14771);
nand UO_1639 (O_1639,N_14737,N_14614);
or UO_1640 (O_1640,N_14484,N_14840);
nand UO_1641 (O_1641,N_14531,N_14568);
and UO_1642 (O_1642,N_14415,N_14307);
nand UO_1643 (O_1643,N_14709,N_14841);
or UO_1644 (O_1644,N_14757,N_14334);
or UO_1645 (O_1645,N_14802,N_14844);
or UO_1646 (O_1646,N_14332,N_14727);
and UO_1647 (O_1647,N_14478,N_14961);
and UO_1648 (O_1648,N_14526,N_14266);
and UO_1649 (O_1649,N_14275,N_14786);
or UO_1650 (O_1650,N_14922,N_14600);
or UO_1651 (O_1651,N_14436,N_14592);
or UO_1652 (O_1652,N_14592,N_14948);
and UO_1653 (O_1653,N_14304,N_14502);
or UO_1654 (O_1654,N_14964,N_14412);
nor UO_1655 (O_1655,N_14479,N_14863);
and UO_1656 (O_1656,N_14285,N_14327);
nor UO_1657 (O_1657,N_14822,N_14535);
or UO_1658 (O_1658,N_14275,N_14549);
nor UO_1659 (O_1659,N_14336,N_14564);
or UO_1660 (O_1660,N_14733,N_14865);
nor UO_1661 (O_1661,N_14768,N_14733);
or UO_1662 (O_1662,N_14370,N_14766);
and UO_1663 (O_1663,N_14566,N_14345);
or UO_1664 (O_1664,N_14672,N_14833);
or UO_1665 (O_1665,N_14712,N_14463);
or UO_1666 (O_1666,N_14917,N_14375);
and UO_1667 (O_1667,N_14742,N_14823);
nand UO_1668 (O_1668,N_14689,N_14388);
or UO_1669 (O_1669,N_14995,N_14766);
or UO_1670 (O_1670,N_14789,N_14835);
nand UO_1671 (O_1671,N_14860,N_14363);
xor UO_1672 (O_1672,N_14709,N_14532);
nand UO_1673 (O_1673,N_14899,N_14874);
or UO_1674 (O_1674,N_14430,N_14656);
xor UO_1675 (O_1675,N_14632,N_14829);
xor UO_1676 (O_1676,N_14492,N_14708);
nand UO_1677 (O_1677,N_14267,N_14391);
and UO_1678 (O_1678,N_14429,N_14699);
nor UO_1679 (O_1679,N_14720,N_14900);
or UO_1680 (O_1680,N_14347,N_14548);
or UO_1681 (O_1681,N_14312,N_14768);
nor UO_1682 (O_1682,N_14427,N_14305);
and UO_1683 (O_1683,N_14947,N_14496);
or UO_1684 (O_1684,N_14741,N_14620);
nand UO_1685 (O_1685,N_14547,N_14489);
nand UO_1686 (O_1686,N_14712,N_14555);
and UO_1687 (O_1687,N_14651,N_14601);
nor UO_1688 (O_1688,N_14440,N_14706);
nor UO_1689 (O_1689,N_14722,N_14490);
nand UO_1690 (O_1690,N_14406,N_14866);
nor UO_1691 (O_1691,N_14871,N_14865);
or UO_1692 (O_1692,N_14732,N_14806);
nor UO_1693 (O_1693,N_14611,N_14436);
or UO_1694 (O_1694,N_14821,N_14454);
nor UO_1695 (O_1695,N_14645,N_14688);
nor UO_1696 (O_1696,N_14665,N_14314);
nand UO_1697 (O_1697,N_14329,N_14527);
nor UO_1698 (O_1698,N_14889,N_14345);
nor UO_1699 (O_1699,N_14313,N_14863);
nand UO_1700 (O_1700,N_14973,N_14422);
nand UO_1701 (O_1701,N_14931,N_14409);
or UO_1702 (O_1702,N_14976,N_14542);
or UO_1703 (O_1703,N_14859,N_14901);
nand UO_1704 (O_1704,N_14556,N_14788);
and UO_1705 (O_1705,N_14992,N_14825);
xor UO_1706 (O_1706,N_14676,N_14426);
nor UO_1707 (O_1707,N_14566,N_14631);
nor UO_1708 (O_1708,N_14349,N_14485);
nand UO_1709 (O_1709,N_14662,N_14491);
xor UO_1710 (O_1710,N_14866,N_14898);
nand UO_1711 (O_1711,N_14628,N_14483);
nor UO_1712 (O_1712,N_14687,N_14859);
or UO_1713 (O_1713,N_14578,N_14750);
nor UO_1714 (O_1714,N_14779,N_14389);
nor UO_1715 (O_1715,N_14383,N_14930);
xnor UO_1716 (O_1716,N_14378,N_14595);
nand UO_1717 (O_1717,N_14972,N_14304);
xor UO_1718 (O_1718,N_14933,N_14600);
xor UO_1719 (O_1719,N_14402,N_14916);
nor UO_1720 (O_1720,N_14970,N_14477);
nor UO_1721 (O_1721,N_14435,N_14728);
nor UO_1722 (O_1722,N_14323,N_14788);
and UO_1723 (O_1723,N_14741,N_14293);
nor UO_1724 (O_1724,N_14908,N_14650);
and UO_1725 (O_1725,N_14666,N_14396);
xor UO_1726 (O_1726,N_14509,N_14823);
or UO_1727 (O_1727,N_14932,N_14396);
nand UO_1728 (O_1728,N_14595,N_14625);
or UO_1729 (O_1729,N_14533,N_14849);
or UO_1730 (O_1730,N_14810,N_14580);
xnor UO_1731 (O_1731,N_14521,N_14640);
or UO_1732 (O_1732,N_14805,N_14655);
nand UO_1733 (O_1733,N_14851,N_14385);
nand UO_1734 (O_1734,N_14839,N_14840);
nand UO_1735 (O_1735,N_14332,N_14503);
nand UO_1736 (O_1736,N_14315,N_14732);
or UO_1737 (O_1737,N_14809,N_14949);
or UO_1738 (O_1738,N_14966,N_14467);
or UO_1739 (O_1739,N_14310,N_14790);
and UO_1740 (O_1740,N_14745,N_14613);
and UO_1741 (O_1741,N_14687,N_14564);
nand UO_1742 (O_1742,N_14734,N_14902);
and UO_1743 (O_1743,N_14564,N_14908);
nand UO_1744 (O_1744,N_14386,N_14538);
nor UO_1745 (O_1745,N_14419,N_14535);
nand UO_1746 (O_1746,N_14725,N_14407);
or UO_1747 (O_1747,N_14405,N_14494);
or UO_1748 (O_1748,N_14698,N_14334);
or UO_1749 (O_1749,N_14433,N_14779);
nand UO_1750 (O_1750,N_14380,N_14450);
and UO_1751 (O_1751,N_14886,N_14887);
nor UO_1752 (O_1752,N_14300,N_14796);
nand UO_1753 (O_1753,N_14646,N_14980);
or UO_1754 (O_1754,N_14462,N_14882);
nor UO_1755 (O_1755,N_14667,N_14728);
nor UO_1756 (O_1756,N_14606,N_14718);
and UO_1757 (O_1757,N_14477,N_14995);
and UO_1758 (O_1758,N_14518,N_14416);
or UO_1759 (O_1759,N_14575,N_14972);
nor UO_1760 (O_1760,N_14847,N_14855);
nand UO_1761 (O_1761,N_14996,N_14568);
and UO_1762 (O_1762,N_14295,N_14846);
or UO_1763 (O_1763,N_14571,N_14361);
nor UO_1764 (O_1764,N_14496,N_14437);
nor UO_1765 (O_1765,N_14963,N_14766);
and UO_1766 (O_1766,N_14781,N_14882);
or UO_1767 (O_1767,N_14443,N_14869);
nor UO_1768 (O_1768,N_14806,N_14985);
nand UO_1769 (O_1769,N_14687,N_14332);
nor UO_1770 (O_1770,N_14797,N_14880);
and UO_1771 (O_1771,N_14311,N_14753);
nand UO_1772 (O_1772,N_14683,N_14346);
or UO_1773 (O_1773,N_14674,N_14412);
and UO_1774 (O_1774,N_14801,N_14545);
nand UO_1775 (O_1775,N_14541,N_14398);
nor UO_1776 (O_1776,N_14256,N_14891);
and UO_1777 (O_1777,N_14695,N_14394);
or UO_1778 (O_1778,N_14646,N_14549);
nor UO_1779 (O_1779,N_14842,N_14671);
and UO_1780 (O_1780,N_14950,N_14278);
xnor UO_1781 (O_1781,N_14725,N_14378);
nand UO_1782 (O_1782,N_14670,N_14887);
nor UO_1783 (O_1783,N_14590,N_14254);
nor UO_1784 (O_1784,N_14653,N_14706);
nand UO_1785 (O_1785,N_14489,N_14765);
and UO_1786 (O_1786,N_14734,N_14814);
or UO_1787 (O_1787,N_14888,N_14541);
and UO_1788 (O_1788,N_14447,N_14652);
nor UO_1789 (O_1789,N_14795,N_14544);
nand UO_1790 (O_1790,N_14862,N_14790);
xor UO_1791 (O_1791,N_14951,N_14764);
and UO_1792 (O_1792,N_14798,N_14325);
xor UO_1793 (O_1793,N_14354,N_14428);
or UO_1794 (O_1794,N_14760,N_14389);
and UO_1795 (O_1795,N_14977,N_14845);
nor UO_1796 (O_1796,N_14269,N_14803);
xor UO_1797 (O_1797,N_14606,N_14789);
xnor UO_1798 (O_1798,N_14660,N_14259);
and UO_1799 (O_1799,N_14469,N_14397);
and UO_1800 (O_1800,N_14279,N_14984);
nand UO_1801 (O_1801,N_14328,N_14270);
or UO_1802 (O_1802,N_14987,N_14434);
nand UO_1803 (O_1803,N_14869,N_14329);
and UO_1804 (O_1804,N_14387,N_14590);
nor UO_1805 (O_1805,N_14467,N_14376);
nand UO_1806 (O_1806,N_14907,N_14516);
nand UO_1807 (O_1807,N_14562,N_14358);
or UO_1808 (O_1808,N_14740,N_14386);
nand UO_1809 (O_1809,N_14333,N_14715);
and UO_1810 (O_1810,N_14340,N_14624);
nor UO_1811 (O_1811,N_14992,N_14836);
nor UO_1812 (O_1812,N_14412,N_14612);
and UO_1813 (O_1813,N_14816,N_14541);
nand UO_1814 (O_1814,N_14383,N_14251);
xnor UO_1815 (O_1815,N_14646,N_14589);
nor UO_1816 (O_1816,N_14528,N_14668);
nand UO_1817 (O_1817,N_14337,N_14919);
or UO_1818 (O_1818,N_14901,N_14448);
nor UO_1819 (O_1819,N_14793,N_14848);
and UO_1820 (O_1820,N_14556,N_14578);
and UO_1821 (O_1821,N_14951,N_14597);
nor UO_1822 (O_1822,N_14510,N_14895);
nor UO_1823 (O_1823,N_14870,N_14631);
or UO_1824 (O_1824,N_14614,N_14536);
and UO_1825 (O_1825,N_14325,N_14606);
or UO_1826 (O_1826,N_14323,N_14380);
nor UO_1827 (O_1827,N_14396,N_14665);
xnor UO_1828 (O_1828,N_14727,N_14341);
or UO_1829 (O_1829,N_14900,N_14320);
or UO_1830 (O_1830,N_14407,N_14780);
nor UO_1831 (O_1831,N_14334,N_14663);
or UO_1832 (O_1832,N_14340,N_14487);
or UO_1833 (O_1833,N_14427,N_14611);
nor UO_1834 (O_1834,N_14793,N_14312);
nand UO_1835 (O_1835,N_14265,N_14448);
nor UO_1836 (O_1836,N_14537,N_14602);
nand UO_1837 (O_1837,N_14701,N_14386);
nor UO_1838 (O_1838,N_14808,N_14597);
xnor UO_1839 (O_1839,N_14690,N_14766);
xor UO_1840 (O_1840,N_14412,N_14912);
or UO_1841 (O_1841,N_14633,N_14310);
nand UO_1842 (O_1842,N_14293,N_14332);
or UO_1843 (O_1843,N_14303,N_14609);
or UO_1844 (O_1844,N_14867,N_14492);
nor UO_1845 (O_1845,N_14793,N_14854);
nor UO_1846 (O_1846,N_14705,N_14656);
or UO_1847 (O_1847,N_14493,N_14358);
nand UO_1848 (O_1848,N_14261,N_14626);
nor UO_1849 (O_1849,N_14881,N_14577);
or UO_1850 (O_1850,N_14752,N_14687);
or UO_1851 (O_1851,N_14540,N_14424);
or UO_1852 (O_1852,N_14348,N_14288);
nand UO_1853 (O_1853,N_14962,N_14375);
or UO_1854 (O_1854,N_14436,N_14275);
nor UO_1855 (O_1855,N_14741,N_14918);
nand UO_1856 (O_1856,N_14852,N_14714);
xor UO_1857 (O_1857,N_14784,N_14993);
or UO_1858 (O_1858,N_14356,N_14695);
nand UO_1859 (O_1859,N_14734,N_14342);
or UO_1860 (O_1860,N_14370,N_14703);
nand UO_1861 (O_1861,N_14447,N_14250);
and UO_1862 (O_1862,N_14650,N_14346);
or UO_1863 (O_1863,N_14546,N_14864);
or UO_1864 (O_1864,N_14606,N_14423);
nor UO_1865 (O_1865,N_14968,N_14301);
and UO_1866 (O_1866,N_14598,N_14546);
nand UO_1867 (O_1867,N_14559,N_14305);
or UO_1868 (O_1868,N_14386,N_14377);
xor UO_1869 (O_1869,N_14847,N_14950);
nor UO_1870 (O_1870,N_14664,N_14287);
and UO_1871 (O_1871,N_14627,N_14626);
nor UO_1872 (O_1872,N_14617,N_14862);
or UO_1873 (O_1873,N_14309,N_14664);
or UO_1874 (O_1874,N_14530,N_14753);
nor UO_1875 (O_1875,N_14420,N_14507);
nor UO_1876 (O_1876,N_14521,N_14342);
nand UO_1877 (O_1877,N_14852,N_14341);
and UO_1878 (O_1878,N_14918,N_14636);
xor UO_1879 (O_1879,N_14827,N_14661);
xor UO_1880 (O_1880,N_14989,N_14287);
xor UO_1881 (O_1881,N_14267,N_14872);
nor UO_1882 (O_1882,N_14718,N_14978);
nand UO_1883 (O_1883,N_14648,N_14873);
or UO_1884 (O_1884,N_14720,N_14624);
and UO_1885 (O_1885,N_14967,N_14813);
nor UO_1886 (O_1886,N_14961,N_14957);
nand UO_1887 (O_1887,N_14756,N_14980);
or UO_1888 (O_1888,N_14946,N_14334);
nor UO_1889 (O_1889,N_14299,N_14876);
and UO_1890 (O_1890,N_14515,N_14493);
or UO_1891 (O_1891,N_14395,N_14932);
or UO_1892 (O_1892,N_14877,N_14640);
nand UO_1893 (O_1893,N_14818,N_14370);
nor UO_1894 (O_1894,N_14645,N_14979);
or UO_1895 (O_1895,N_14897,N_14780);
nand UO_1896 (O_1896,N_14890,N_14521);
nand UO_1897 (O_1897,N_14433,N_14275);
and UO_1898 (O_1898,N_14767,N_14612);
or UO_1899 (O_1899,N_14268,N_14860);
and UO_1900 (O_1900,N_14334,N_14602);
nor UO_1901 (O_1901,N_14704,N_14991);
nand UO_1902 (O_1902,N_14632,N_14334);
nand UO_1903 (O_1903,N_14359,N_14483);
or UO_1904 (O_1904,N_14848,N_14257);
nand UO_1905 (O_1905,N_14379,N_14609);
and UO_1906 (O_1906,N_14698,N_14413);
nor UO_1907 (O_1907,N_14958,N_14456);
xnor UO_1908 (O_1908,N_14859,N_14704);
and UO_1909 (O_1909,N_14433,N_14383);
nand UO_1910 (O_1910,N_14635,N_14551);
nor UO_1911 (O_1911,N_14570,N_14931);
or UO_1912 (O_1912,N_14712,N_14886);
nor UO_1913 (O_1913,N_14357,N_14502);
and UO_1914 (O_1914,N_14390,N_14651);
or UO_1915 (O_1915,N_14855,N_14986);
nand UO_1916 (O_1916,N_14662,N_14416);
and UO_1917 (O_1917,N_14589,N_14303);
nor UO_1918 (O_1918,N_14582,N_14459);
nor UO_1919 (O_1919,N_14448,N_14815);
nor UO_1920 (O_1920,N_14731,N_14535);
nor UO_1921 (O_1921,N_14679,N_14448);
or UO_1922 (O_1922,N_14623,N_14621);
and UO_1923 (O_1923,N_14966,N_14667);
nand UO_1924 (O_1924,N_14655,N_14424);
nor UO_1925 (O_1925,N_14515,N_14915);
nand UO_1926 (O_1926,N_14506,N_14920);
or UO_1927 (O_1927,N_14585,N_14673);
nor UO_1928 (O_1928,N_14637,N_14528);
and UO_1929 (O_1929,N_14910,N_14376);
and UO_1930 (O_1930,N_14874,N_14553);
xnor UO_1931 (O_1931,N_14656,N_14667);
xor UO_1932 (O_1932,N_14419,N_14791);
or UO_1933 (O_1933,N_14263,N_14267);
nor UO_1934 (O_1934,N_14311,N_14677);
nand UO_1935 (O_1935,N_14989,N_14564);
and UO_1936 (O_1936,N_14874,N_14937);
nand UO_1937 (O_1937,N_14900,N_14276);
xnor UO_1938 (O_1938,N_14612,N_14899);
and UO_1939 (O_1939,N_14860,N_14399);
nand UO_1940 (O_1940,N_14406,N_14509);
nor UO_1941 (O_1941,N_14597,N_14569);
nand UO_1942 (O_1942,N_14336,N_14326);
nor UO_1943 (O_1943,N_14516,N_14473);
nand UO_1944 (O_1944,N_14355,N_14446);
and UO_1945 (O_1945,N_14965,N_14755);
or UO_1946 (O_1946,N_14971,N_14308);
nor UO_1947 (O_1947,N_14820,N_14816);
and UO_1948 (O_1948,N_14669,N_14439);
nor UO_1949 (O_1949,N_14421,N_14656);
nor UO_1950 (O_1950,N_14836,N_14734);
and UO_1951 (O_1951,N_14370,N_14300);
nor UO_1952 (O_1952,N_14344,N_14593);
nor UO_1953 (O_1953,N_14529,N_14805);
and UO_1954 (O_1954,N_14799,N_14542);
nor UO_1955 (O_1955,N_14641,N_14785);
nand UO_1956 (O_1956,N_14465,N_14306);
and UO_1957 (O_1957,N_14597,N_14592);
nand UO_1958 (O_1958,N_14457,N_14577);
and UO_1959 (O_1959,N_14733,N_14817);
xnor UO_1960 (O_1960,N_14958,N_14440);
and UO_1961 (O_1961,N_14702,N_14768);
and UO_1962 (O_1962,N_14657,N_14331);
and UO_1963 (O_1963,N_14355,N_14519);
nor UO_1964 (O_1964,N_14405,N_14763);
or UO_1965 (O_1965,N_14517,N_14400);
xnor UO_1966 (O_1966,N_14911,N_14506);
or UO_1967 (O_1967,N_14760,N_14625);
or UO_1968 (O_1968,N_14964,N_14548);
nand UO_1969 (O_1969,N_14347,N_14744);
nand UO_1970 (O_1970,N_14972,N_14558);
nand UO_1971 (O_1971,N_14375,N_14633);
xnor UO_1972 (O_1972,N_14472,N_14750);
nor UO_1973 (O_1973,N_14708,N_14807);
nor UO_1974 (O_1974,N_14541,N_14834);
nand UO_1975 (O_1975,N_14806,N_14563);
nor UO_1976 (O_1976,N_14745,N_14628);
and UO_1977 (O_1977,N_14512,N_14594);
and UO_1978 (O_1978,N_14975,N_14346);
nand UO_1979 (O_1979,N_14386,N_14439);
or UO_1980 (O_1980,N_14426,N_14609);
nand UO_1981 (O_1981,N_14760,N_14511);
nand UO_1982 (O_1982,N_14557,N_14712);
and UO_1983 (O_1983,N_14382,N_14754);
and UO_1984 (O_1984,N_14685,N_14786);
and UO_1985 (O_1985,N_14476,N_14898);
nand UO_1986 (O_1986,N_14398,N_14428);
xor UO_1987 (O_1987,N_14687,N_14881);
nand UO_1988 (O_1988,N_14860,N_14386);
and UO_1989 (O_1989,N_14394,N_14501);
and UO_1990 (O_1990,N_14779,N_14886);
nor UO_1991 (O_1991,N_14448,N_14942);
or UO_1992 (O_1992,N_14957,N_14567);
nor UO_1993 (O_1993,N_14737,N_14799);
nand UO_1994 (O_1994,N_14796,N_14921);
nor UO_1995 (O_1995,N_14283,N_14818);
nand UO_1996 (O_1996,N_14347,N_14650);
nand UO_1997 (O_1997,N_14557,N_14928);
or UO_1998 (O_1998,N_14669,N_14927);
nor UO_1999 (O_1999,N_14857,N_14851);
endmodule