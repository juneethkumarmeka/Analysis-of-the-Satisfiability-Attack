module basic_500_3000_500_50_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xor U0 (N_0,In_139,In_168);
or U1 (N_1,In_224,In_194);
xnor U2 (N_2,In_348,In_433);
or U3 (N_3,In_22,In_101);
nor U4 (N_4,In_333,In_442);
nand U5 (N_5,In_146,In_70);
nand U6 (N_6,In_418,In_13);
xor U7 (N_7,In_327,In_371);
and U8 (N_8,In_205,In_377);
and U9 (N_9,In_459,In_378);
and U10 (N_10,In_119,In_435);
xor U11 (N_11,In_83,In_272);
nand U12 (N_12,In_249,In_282);
nand U13 (N_13,In_454,In_156);
or U14 (N_14,In_108,In_417);
or U15 (N_15,In_438,In_488);
nor U16 (N_16,In_99,In_240);
nor U17 (N_17,In_374,In_24);
xor U18 (N_18,In_117,In_40);
nand U19 (N_19,In_15,In_323);
xnor U20 (N_20,In_293,In_127);
and U21 (N_21,In_447,In_346);
nor U22 (N_22,In_299,In_344);
xnor U23 (N_23,In_50,In_495);
xnor U24 (N_24,In_18,In_120);
or U25 (N_25,In_431,In_180);
and U26 (N_26,In_265,In_430);
nor U27 (N_27,In_332,In_36);
or U28 (N_28,In_204,In_468);
or U29 (N_29,In_76,In_86);
nor U30 (N_30,In_109,In_58);
or U31 (N_31,In_392,In_362);
or U32 (N_32,In_319,In_463);
or U33 (N_33,In_111,In_302);
nand U34 (N_34,In_211,In_31);
nand U35 (N_35,In_144,In_386);
nor U36 (N_36,In_399,In_255);
nor U37 (N_37,In_421,In_169);
nor U38 (N_38,In_223,In_123);
and U39 (N_39,In_440,In_486);
and U40 (N_40,In_356,In_179);
and U41 (N_41,In_147,In_400);
nand U42 (N_42,In_263,In_242);
nand U43 (N_43,In_72,In_264);
or U44 (N_44,In_472,In_477);
or U45 (N_45,In_89,In_148);
nand U46 (N_46,In_458,In_206);
and U47 (N_47,In_260,In_30);
and U48 (N_48,In_16,In_469);
nand U49 (N_49,In_173,In_373);
or U50 (N_50,In_239,In_390);
nand U51 (N_51,In_404,In_275);
or U52 (N_52,In_107,In_256);
xor U53 (N_53,In_230,In_63);
and U54 (N_54,In_121,In_322);
nor U55 (N_55,In_286,In_296);
nor U56 (N_56,In_132,In_368);
xor U57 (N_57,In_94,In_411);
or U58 (N_58,In_443,In_301);
or U59 (N_59,In_324,In_441);
and U60 (N_60,In_217,In_163);
xnor U61 (N_61,In_175,In_184);
xor U62 (N_62,In_188,In_64);
and U63 (N_63,In_73,In_308);
or U64 (N_64,In_424,In_232);
and U65 (N_65,N_58,In_420);
nor U66 (N_66,In_383,In_406);
nand U67 (N_67,N_30,In_226);
and U68 (N_68,In_74,In_100);
nand U69 (N_69,In_492,In_314);
nor U70 (N_70,In_457,In_212);
and U71 (N_71,In_3,In_246);
nor U72 (N_72,N_6,In_353);
nand U73 (N_73,N_5,In_423);
nor U74 (N_74,In_177,In_401);
and U75 (N_75,In_485,In_251);
or U76 (N_76,In_498,N_59);
or U77 (N_77,In_408,N_37);
nor U78 (N_78,In_398,In_379);
or U79 (N_79,N_56,N_23);
nor U80 (N_80,In_25,In_416);
xor U81 (N_81,In_27,In_278);
or U82 (N_82,In_358,In_476);
and U83 (N_83,In_419,In_351);
and U84 (N_84,In_167,In_285);
or U85 (N_85,In_185,In_41);
xor U86 (N_86,In_145,In_237);
and U87 (N_87,In_65,In_381);
or U88 (N_88,In_32,In_228);
or U89 (N_89,In_234,In_466);
or U90 (N_90,In_385,In_110);
nand U91 (N_91,In_129,In_300);
xnor U92 (N_92,In_162,In_93);
nand U93 (N_93,In_59,In_269);
xor U94 (N_94,In_290,In_279);
nand U95 (N_95,In_79,In_236);
xor U96 (N_96,In_292,N_41);
or U97 (N_97,In_53,In_181);
nor U98 (N_98,In_436,In_5);
and U99 (N_99,In_48,N_22);
nor U100 (N_100,In_432,In_428);
nand U101 (N_101,In_456,In_85);
or U102 (N_102,In_387,In_200);
nand U103 (N_103,In_23,In_310);
nand U104 (N_104,N_20,In_287);
nand U105 (N_105,In_315,In_341);
or U106 (N_106,N_33,In_81);
or U107 (N_107,In_268,In_45);
or U108 (N_108,In_283,In_176);
nand U109 (N_109,In_484,In_152);
nand U110 (N_110,In_393,N_8);
or U111 (N_111,In_313,In_61);
and U112 (N_112,In_243,In_339);
nand U113 (N_113,In_170,In_75);
nor U114 (N_114,In_467,In_489);
nand U115 (N_115,In_354,N_21);
or U116 (N_116,In_222,In_49);
nand U117 (N_117,In_391,In_388);
nand U118 (N_118,In_78,In_90);
nand U119 (N_119,In_1,N_7);
and U120 (N_120,In_135,In_389);
nand U121 (N_121,In_221,In_395);
nor U122 (N_122,In_330,In_248);
or U123 (N_123,In_4,N_26);
nand U124 (N_124,N_119,In_274);
xor U125 (N_125,In_481,In_104);
nand U126 (N_126,N_2,N_18);
and U127 (N_127,In_288,N_53);
nand U128 (N_128,N_66,In_318);
nand U129 (N_129,In_210,In_191);
nor U130 (N_130,In_128,In_10);
or U131 (N_131,In_455,In_122);
nand U132 (N_132,In_462,In_271);
and U133 (N_133,N_111,N_28);
and U134 (N_134,In_158,N_63);
xor U135 (N_135,N_69,N_47);
and U136 (N_136,In_360,In_257);
xor U137 (N_137,In_67,In_483);
or U138 (N_138,In_56,N_44);
and U139 (N_139,In_241,In_62);
nand U140 (N_140,In_273,In_141);
nor U141 (N_141,N_55,In_87);
or U142 (N_142,In_337,N_14);
nor U143 (N_143,In_267,In_494);
or U144 (N_144,N_29,In_238);
xor U145 (N_145,In_247,In_326);
or U146 (N_146,In_277,In_34);
or U147 (N_147,In_172,In_231);
and U148 (N_148,In_452,N_84);
nand U149 (N_149,N_89,In_289);
nand U150 (N_150,In_215,In_20);
and U151 (N_151,In_422,N_31);
nand U152 (N_152,In_336,In_77);
nand U153 (N_153,N_113,N_115);
nand U154 (N_154,N_12,In_97);
xnor U155 (N_155,N_40,In_253);
and U156 (N_156,In_298,In_270);
xnor U157 (N_157,N_67,N_51);
nand U158 (N_158,In_198,In_195);
xor U159 (N_159,N_97,In_51);
nor U160 (N_160,In_19,In_325);
nand U161 (N_161,In_355,In_434);
nand U162 (N_162,In_493,In_92);
nand U163 (N_163,N_19,In_186);
or U164 (N_164,In_297,In_305);
or U165 (N_165,N_94,In_491);
nand U166 (N_166,In_80,In_12);
and U167 (N_167,N_27,In_44);
or U168 (N_168,In_118,In_410);
nand U169 (N_169,In_17,N_15);
xnor U170 (N_170,In_258,In_328);
nor U171 (N_171,N_36,In_312);
and U172 (N_172,In_28,In_105);
or U173 (N_173,N_62,In_439);
and U174 (N_174,N_108,In_370);
nor U175 (N_175,In_266,In_449);
or U176 (N_176,N_101,In_475);
and U177 (N_177,In_331,In_470);
or U178 (N_178,In_193,In_465);
nor U179 (N_179,N_79,In_235);
nand U180 (N_180,In_309,In_88);
nand U181 (N_181,In_66,In_153);
or U182 (N_182,N_125,In_233);
nor U183 (N_183,N_128,N_157);
nand U184 (N_184,In_403,In_219);
and U185 (N_185,In_114,N_81);
and U186 (N_186,In_39,N_3);
nor U187 (N_187,N_123,N_34);
and U188 (N_188,N_112,In_409);
or U189 (N_189,In_159,N_132);
nor U190 (N_190,In_208,In_306);
nand U191 (N_191,N_73,N_61);
and U192 (N_192,N_76,In_349);
or U193 (N_193,In_473,N_156);
xor U194 (N_194,In_142,In_124);
or U195 (N_195,In_218,In_497);
or U196 (N_196,In_451,In_499);
nor U197 (N_197,N_16,N_116);
nand U198 (N_198,In_453,In_91);
nand U199 (N_199,N_130,In_479);
nand U200 (N_200,N_126,In_480);
and U201 (N_201,In_414,In_150);
nor U202 (N_202,In_82,N_121);
xor U203 (N_203,N_91,In_164);
or U204 (N_204,N_32,N_122);
or U205 (N_205,In_149,In_376);
nand U206 (N_206,N_96,N_104);
nand U207 (N_207,In_33,In_250);
or U208 (N_208,N_154,N_98);
and U209 (N_209,In_471,In_8);
and U210 (N_210,N_78,N_48);
and U211 (N_211,In_427,N_45);
or U212 (N_212,N_93,N_117);
or U213 (N_213,N_167,In_244);
xnor U214 (N_214,N_25,In_137);
nor U215 (N_215,N_4,N_71);
and U216 (N_216,N_118,In_95);
or U217 (N_217,N_151,N_106);
nand U218 (N_218,N_95,N_50);
or U219 (N_219,In_166,N_137);
and U220 (N_220,In_369,N_145);
nor U221 (N_221,In_357,In_216);
nor U222 (N_222,In_347,N_72);
and U223 (N_223,In_199,In_155);
or U224 (N_224,In_203,In_461);
nand U225 (N_225,In_0,In_464);
xnor U226 (N_226,In_366,In_55);
and U227 (N_227,N_179,In_113);
nand U228 (N_228,In_364,In_133);
or U229 (N_229,In_316,In_307);
nor U230 (N_230,In_182,In_187);
or U231 (N_231,In_69,N_85);
or U232 (N_232,In_227,In_189);
nor U233 (N_233,In_294,In_2);
and U234 (N_234,In_57,In_397);
xnor U235 (N_235,In_54,N_90);
nor U236 (N_236,N_49,In_245);
or U237 (N_237,N_162,In_350);
or U238 (N_238,N_46,N_83);
and U239 (N_239,In_130,In_68);
nand U240 (N_240,In_437,N_223);
nor U241 (N_241,N_213,N_149);
nor U242 (N_242,In_487,In_384);
xor U243 (N_243,N_136,In_138);
xor U244 (N_244,In_157,In_84);
and U245 (N_245,N_171,In_303);
or U246 (N_246,N_212,N_215);
xor U247 (N_247,N_120,In_340);
nand U248 (N_248,In_21,N_153);
or U249 (N_249,In_214,In_412);
xor U250 (N_250,N_184,In_276);
nand U251 (N_251,N_204,N_180);
and U252 (N_252,N_86,In_343);
or U253 (N_253,N_127,In_413);
nor U254 (N_254,N_211,N_208);
xor U255 (N_255,N_39,N_54);
nand U256 (N_256,N_60,N_205);
nor U257 (N_257,In_35,N_166);
nor U258 (N_258,In_281,N_134);
nand U259 (N_259,In_284,N_177);
nand U260 (N_260,N_185,In_151);
or U261 (N_261,N_192,In_261);
nand U262 (N_262,N_82,In_375);
and U263 (N_263,N_24,N_9);
and U264 (N_264,In_96,N_77);
or U265 (N_265,N_43,N_170);
xor U266 (N_266,N_176,N_183);
or U267 (N_267,In_329,N_232);
and U268 (N_268,N_196,In_42);
xnor U269 (N_269,N_200,N_168);
and U270 (N_270,In_52,In_9);
xor U271 (N_271,In_160,N_158);
nand U272 (N_272,In_363,In_482);
and U273 (N_273,In_26,N_107);
and U274 (N_274,In_425,N_109);
or U275 (N_275,In_154,N_218);
nor U276 (N_276,In_71,In_334);
nand U277 (N_277,N_114,N_230);
or U278 (N_278,N_131,N_146);
nand U279 (N_279,N_105,In_134);
xor U280 (N_280,N_175,In_380);
and U281 (N_281,N_234,N_10);
nor U282 (N_282,N_207,In_254);
and U283 (N_283,In_382,N_237);
and U284 (N_284,N_220,In_490);
nor U285 (N_285,In_174,N_163);
or U286 (N_286,N_159,In_225);
nand U287 (N_287,In_98,N_219);
and U288 (N_288,In_38,N_225);
nor U289 (N_289,In_259,N_182);
nand U290 (N_290,N_201,N_235);
xor U291 (N_291,In_280,N_203);
nand U292 (N_292,In_396,N_138);
nand U293 (N_293,N_238,In_429);
or U294 (N_294,In_444,In_7);
or U295 (N_295,In_201,In_304);
nor U296 (N_296,N_227,In_474);
nor U297 (N_297,In_402,N_141);
nand U298 (N_298,In_207,N_217);
nand U299 (N_299,N_155,In_125);
nor U300 (N_300,N_129,N_271);
nor U301 (N_301,N_279,N_259);
nand U302 (N_302,N_268,N_216);
nor U303 (N_303,N_276,In_448);
nand U304 (N_304,N_75,N_133);
or U305 (N_305,N_261,N_296);
nor U306 (N_306,In_365,In_415);
nor U307 (N_307,N_173,In_295);
nor U308 (N_308,N_290,N_274);
nor U309 (N_309,In_445,N_257);
nand U310 (N_310,In_136,N_255);
nor U311 (N_311,N_283,N_287);
nand U312 (N_312,N_264,N_253);
nor U313 (N_313,In_37,N_202);
nor U314 (N_314,N_152,In_192);
or U315 (N_315,In_143,N_87);
nor U316 (N_316,N_236,N_252);
xnor U317 (N_317,In_446,N_240);
nor U318 (N_318,N_165,In_320);
xnor U319 (N_319,N_293,In_60);
nor U320 (N_320,N_57,N_110);
nand U321 (N_321,N_228,N_172);
nor U322 (N_322,In_178,In_126);
nand U323 (N_323,N_102,N_187);
and U324 (N_324,N_249,N_254);
and U325 (N_325,N_222,N_221);
or U326 (N_326,In_14,In_352);
or U327 (N_327,N_169,N_64);
or U328 (N_328,In_338,N_258);
nor U329 (N_329,N_281,N_35);
xor U330 (N_330,In_407,N_198);
nor U331 (N_331,In_140,In_103);
xor U332 (N_332,N_288,N_193);
or U333 (N_333,In_317,N_299);
and U334 (N_334,In_190,N_242);
or U335 (N_335,N_297,In_460);
and U336 (N_336,N_139,N_197);
and U337 (N_337,N_265,N_277);
and U338 (N_338,N_38,N_224);
nand U339 (N_339,In_478,N_239);
and U340 (N_340,N_190,N_248);
xor U341 (N_341,N_199,N_269);
or U342 (N_342,N_143,N_68);
xor U343 (N_343,N_260,N_243);
and U344 (N_344,N_285,In_372);
nor U345 (N_345,In_102,N_263);
nand U346 (N_346,N_178,N_144);
or U347 (N_347,N_17,N_289);
or U348 (N_348,N_245,In_116);
or U349 (N_349,N_92,N_181);
nor U350 (N_350,N_65,N_150);
nor U351 (N_351,N_292,In_196);
nand U352 (N_352,N_226,In_426);
nor U353 (N_353,N_266,In_359);
or U354 (N_354,N_99,N_147);
or U355 (N_355,In_183,N_209);
nand U356 (N_356,N_0,N_42);
and U357 (N_357,N_278,In_367);
xnor U358 (N_358,N_103,N_206);
and U359 (N_359,N_191,N_80);
xor U360 (N_360,N_250,N_328);
xnor U361 (N_361,N_359,N_74);
or U362 (N_362,N_194,In_47);
nand U363 (N_363,N_313,N_309);
nand U364 (N_364,N_341,N_241);
or U365 (N_365,In_335,In_321);
nand U366 (N_366,N_210,N_308);
or U367 (N_367,N_246,In_213);
xor U368 (N_368,N_339,N_352);
or U369 (N_369,N_333,N_334);
and U370 (N_370,N_124,N_302);
nor U371 (N_371,N_315,In_394);
or U372 (N_372,N_160,In_11);
or U373 (N_373,N_161,N_357);
and U374 (N_374,N_327,N_1);
nand U375 (N_375,N_353,N_195);
and U376 (N_376,N_314,N_319);
xor U377 (N_377,N_310,N_135);
xnor U378 (N_378,N_188,N_256);
xor U379 (N_379,N_262,N_70);
and U380 (N_380,N_303,N_356);
nand U381 (N_381,N_164,N_291);
nor U382 (N_382,N_11,N_300);
or U383 (N_383,N_312,N_251);
and U384 (N_384,N_358,N_140);
nand U385 (N_385,N_244,In_46);
nor U386 (N_386,N_294,N_343);
nand U387 (N_387,N_344,N_305);
or U388 (N_388,In_165,In_43);
nand U389 (N_389,N_13,N_316);
nor U390 (N_390,N_325,In_450);
nor U391 (N_391,N_186,In_291);
nor U392 (N_392,In_29,In_262);
nand U393 (N_393,In_345,N_273);
nor U394 (N_394,N_324,In_361);
xor U395 (N_395,In_252,N_337);
xor U396 (N_396,N_272,In_496);
xor U397 (N_397,N_52,N_295);
or U398 (N_398,N_286,N_329);
or U399 (N_399,N_347,N_354);
nor U400 (N_400,N_340,In_405);
and U401 (N_401,In_161,N_317);
nand U402 (N_402,In_106,N_142);
nor U403 (N_403,In_311,In_112);
nor U404 (N_404,N_321,N_306);
nand U405 (N_405,N_275,N_304);
or U406 (N_406,N_267,N_247);
or U407 (N_407,N_331,N_351);
nor U408 (N_408,N_88,N_189);
nand U409 (N_409,N_280,N_326);
xor U410 (N_410,N_349,N_270);
xnor U411 (N_411,N_348,N_301);
nor U412 (N_412,N_229,N_336);
nand U413 (N_413,In_197,In_220);
xor U414 (N_414,N_345,N_100);
nand U415 (N_415,N_338,In_6);
and U416 (N_416,In_209,In_342);
nand U417 (N_417,N_311,N_307);
nor U418 (N_418,N_342,N_233);
and U419 (N_419,N_174,In_115);
nor U420 (N_420,N_378,N_363);
nor U421 (N_421,N_400,N_346);
or U422 (N_422,N_322,N_368);
nor U423 (N_423,N_365,N_407);
nor U424 (N_424,N_391,N_214);
or U425 (N_425,N_369,N_380);
or U426 (N_426,N_397,N_298);
nand U427 (N_427,N_371,N_405);
xor U428 (N_428,N_362,In_229);
or U429 (N_429,N_381,N_379);
or U430 (N_430,N_389,N_383);
nand U431 (N_431,N_386,In_131);
nor U432 (N_432,N_402,N_387);
nor U433 (N_433,N_370,N_366);
nor U434 (N_434,N_148,N_373);
or U435 (N_435,N_355,N_374);
and U436 (N_436,N_367,N_323);
nand U437 (N_437,N_282,N_411);
xnor U438 (N_438,N_394,N_398);
nor U439 (N_439,N_408,N_418);
nand U440 (N_440,N_335,In_202);
nand U441 (N_441,N_372,N_382);
nand U442 (N_442,N_416,N_284);
nor U443 (N_443,N_388,N_413);
nand U444 (N_444,N_406,N_415);
nand U445 (N_445,N_364,N_395);
nand U446 (N_446,N_390,N_377);
nor U447 (N_447,N_404,N_332);
and U448 (N_448,N_419,N_330);
or U449 (N_449,N_231,N_376);
xnor U450 (N_450,N_385,N_412);
nor U451 (N_451,N_360,N_410);
or U452 (N_452,N_320,N_392);
nor U453 (N_453,N_318,N_375);
xor U454 (N_454,In_171,N_414);
nand U455 (N_455,N_409,N_396);
nor U456 (N_456,N_350,N_417);
or U457 (N_457,N_384,N_403);
and U458 (N_458,N_401,N_393);
or U459 (N_459,N_361,N_399);
xor U460 (N_460,N_364,N_385);
nand U461 (N_461,N_399,N_381);
and U462 (N_462,N_409,N_318);
nor U463 (N_463,N_415,N_366);
nor U464 (N_464,N_409,N_405);
and U465 (N_465,N_375,N_298);
or U466 (N_466,N_371,N_389);
and U467 (N_467,N_418,N_362);
nand U468 (N_468,N_361,N_350);
nor U469 (N_469,N_388,N_373);
or U470 (N_470,N_412,N_413);
or U471 (N_471,N_350,N_397);
or U472 (N_472,N_381,N_388);
and U473 (N_473,N_390,N_335);
nand U474 (N_474,N_369,N_282);
and U475 (N_475,N_408,N_386);
or U476 (N_476,N_411,N_388);
nor U477 (N_477,N_419,N_284);
nor U478 (N_478,N_367,N_318);
and U479 (N_479,N_405,N_369);
nand U480 (N_480,N_436,N_468);
and U481 (N_481,N_432,N_450);
nand U482 (N_482,N_465,N_444);
nand U483 (N_483,N_421,N_441);
nand U484 (N_484,N_478,N_437);
xor U485 (N_485,N_433,N_455);
xor U486 (N_486,N_431,N_438);
nand U487 (N_487,N_459,N_452);
or U488 (N_488,N_449,N_426);
or U489 (N_489,N_479,N_470);
nand U490 (N_490,N_448,N_475);
and U491 (N_491,N_476,N_440);
xnor U492 (N_492,N_451,N_453);
nand U493 (N_493,N_460,N_477);
or U494 (N_494,N_457,N_454);
xnor U495 (N_495,N_435,N_471);
nand U496 (N_496,N_430,N_467);
xor U497 (N_497,N_439,N_469);
nor U498 (N_498,N_447,N_466);
nor U499 (N_499,N_422,N_424);
xor U500 (N_500,N_420,N_423);
and U501 (N_501,N_442,N_463);
and U502 (N_502,N_446,N_474);
nor U503 (N_503,N_428,N_429);
or U504 (N_504,N_464,N_425);
or U505 (N_505,N_434,N_445);
nand U506 (N_506,N_462,N_456);
nand U507 (N_507,N_443,N_427);
xnor U508 (N_508,N_472,N_461);
xnor U509 (N_509,N_473,N_458);
nor U510 (N_510,N_461,N_459);
or U511 (N_511,N_441,N_464);
nor U512 (N_512,N_446,N_430);
and U513 (N_513,N_436,N_425);
or U514 (N_514,N_449,N_479);
and U515 (N_515,N_468,N_430);
or U516 (N_516,N_474,N_471);
and U517 (N_517,N_463,N_439);
or U518 (N_518,N_434,N_423);
or U519 (N_519,N_430,N_463);
nand U520 (N_520,N_437,N_467);
nor U521 (N_521,N_478,N_476);
and U522 (N_522,N_468,N_473);
nor U523 (N_523,N_466,N_474);
or U524 (N_524,N_434,N_470);
nand U525 (N_525,N_432,N_449);
nor U526 (N_526,N_460,N_425);
and U527 (N_527,N_468,N_435);
nor U528 (N_528,N_478,N_425);
and U529 (N_529,N_444,N_425);
xnor U530 (N_530,N_469,N_466);
or U531 (N_531,N_465,N_439);
xnor U532 (N_532,N_464,N_449);
nor U533 (N_533,N_442,N_459);
and U534 (N_534,N_473,N_470);
nor U535 (N_535,N_466,N_454);
nand U536 (N_536,N_461,N_464);
nand U537 (N_537,N_465,N_459);
xnor U538 (N_538,N_471,N_443);
and U539 (N_539,N_456,N_478);
and U540 (N_540,N_535,N_481);
or U541 (N_541,N_504,N_487);
nor U542 (N_542,N_491,N_511);
nand U543 (N_543,N_513,N_518);
or U544 (N_544,N_482,N_501);
nand U545 (N_545,N_495,N_485);
xnor U546 (N_546,N_530,N_525);
or U547 (N_547,N_522,N_538);
xnor U548 (N_548,N_503,N_534);
and U549 (N_549,N_521,N_498);
and U550 (N_550,N_502,N_488);
nand U551 (N_551,N_527,N_492);
nor U552 (N_552,N_515,N_528);
nand U553 (N_553,N_516,N_520);
nor U554 (N_554,N_537,N_507);
or U555 (N_555,N_493,N_514);
and U556 (N_556,N_505,N_529);
nand U557 (N_557,N_539,N_490);
or U558 (N_558,N_496,N_523);
xor U559 (N_559,N_536,N_494);
nor U560 (N_560,N_484,N_524);
nor U561 (N_561,N_483,N_526);
nand U562 (N_562,N_510,N_489);
nor U563 (N_563,N_512,N_533);
xnor U564 (N_564,N_497,N_500);
nor U565 (N_565,N_519,N_480);
and U566 (N_566,N_517,N_532);
and U567 (N_567,N_486,N_508);
nand U568 (N_568,N_531,N_509);
nand U569 (N_569,N_499,N_506);
or U570 (N_570,N_491,N_486);
nand U571 (N_571,N_527,N_536);
or U572 (N_572,N_490,N_499);
or U573 (N_573,N_490,N_513);
and U574 (N_574,N_537,N_492);
nor U575 (N_575,N_487,N_527);
xnor U576 (N_576,N_515,N_536);
nor U577 (N_577,N_507,N_508);
nor U578 (N_578,N_501,N_485);
nor U579 (N_579,N_529,N_539);
xor U580 (N_580,N_515,N_524);
nand U581 (N_581,N_530,N_516);
and U582 (N_582,N_493,N_490);
or U583 (N_583,N_539,N_528);
and U584 (N_584,N_510,N_490);
nor U585 (N_585,N_494,N_505);
and U586 (N_586,N_509,N_483);
or U587 (N_587,N_529,N_498);
nor U588 (N_588,N_493,N_486);
or U589 (N_589,N_508,N_527);
or U590 (N_590,N_505,N_504);
and U591 (N_591,N_516,N_535);
or U592 (N_592,N_521,N_508);
and U593 (N_593,N_513,N_506);
and U594 (N_594,N_496,N_488);
nand U595 (N_595,N_510,N_526);
nor U596 (N_596,N_502,N_503);
nand U597 (N_597,N_483,N_484);
nand U598 (N_598,N_482,N_526);
xor U599 (N_599,N_513,N_511);
xor U600 (N_600,N_551,N_555);
nor U601 (N_601,N_598,N_587);
xnor U602 (N_602,N_562,N_572);
nor U603 (N_603,N_579,N_593);
nor U604 (N_604,N_582,N_599);
or U605 (N_605,N_586,N_574);
nor U606 (N_606,N_557,N_547);
nor U607 (N_607,N_550,N_580);
nand U608 (N_608,N_540,N_556);
and U609 (N_609,N_565,N_564);
and U610 (N_610,N_576,N_573);
nand U611 (N_611,N_591,N_545);
nor U612 (N_612,N_575,N_566);
nand U613 (N_613,N_597,N_596);
and U614 (N_614,N_570,N_569);
or U615 (N_615,N_577,N_542);
nor U616 (N_616,N_541,N_548);
or U617 (N_617,N_558,N_578);
xnor U618 (N_618,N_581,N_567);
and U619 (N_619,N_560,N_595);
or U620 (N_620,N_571,N_554);
nand U621 (N_621,N_552,N_546);
or U622 (N_622,N_585,N_588);
or U623 (N_623,N_559,N_590);
nor U624 (N_624,N_592,N_583);
nand U625 (N_625,N_561,N_543);
nor U626 (N_626,N_584,N_568);
or U627 (N_627,N_544,N_553);
nor U628 (N_628,N_589,N_549);
xnor U629 (N_629,N_563,N_594);
nand U630 (N_630,N_560,N_567);
nor U631 (N_631,N_551,N_588);
nor U632 (N_632,N_549,N_573);
and U633 (N_633,N_546,N_541);
nand U634 (N_634,N_553,N_562);
nand U635 (N_635,N_561,N_558);
nor U636 (N_636,N_596,N_590);
and U637 (N_637,N_571,N_587);
or U638 (N_638,N_592,N_578);
and U639 (N_639,N_572,N_544);
and U640 (N_640,N_564,N_556);
nor U641 (N_641,N_556,N_550);
or U642 (N_642,N_546,N_587);
nand U643 (N_643,N_591,N_569);
or U644 (N_644,N_541,N_571);
and U645 (N_645,N_582,N_567);
and U646 (N_646,N_546,N_599);
or U647 (N_647,N_577,N_554);
and U648 (N_648,N_584,N_550);
or U649 (N_649,N_547,N_581);
and U650 (N_650,N_588,N_554);
and U651 (N_651,N_582,N_580);
nor U652 (N_652,N_577,N_541);
or U653 (N_653,N_544,N_548);
or U654 (N_654,N_542,N_571);
and U655 (N_655,N_599,N_542);
xnor U656 (N_656,N_585,N_546);
and U657 (N_657,N_563,N_570);
nand U658 (N_658,N_595,N_578);
xor U659 (N_659,N_540,N_583);
xor U660 (N_660,N_613,N_602);
nand U661 (N_661,N_618,N_644);
nor U662 (N_662,N_641,N_634);
nor U663 (N_663,N_649,N_629);
or U664 (N_664,N_655,N_652);
nor U665 (N_665,N_621,N_631);
xor U666 (N_666,N_651,N_646);
and U667 (N_667,N_620,N_645);
nor U668 (N_668,N_622,N_654);
xor U669 (N_669,N_657,N_656);
or U670 (N_670,N_611,N_639);
nand U671 (N_671,N_615,N_642);
nand U672 (N_672,N_605,N_647);
nand U673 (N_673,N_606,N_658);
and U674 (N_674,N_640,N_635);
or U675 (N_675,N_653,N_628);
nand U676 (N_676,N_617,N_625);
xor U677 (N_677,N_616,N_648);
nor U678 (N_678,N_604,N_636);
xor U679 (N_679,N_627,N_607);
and U680 (N_680,N_603,N_609);
nand U681 (N_681,N_623,N_608);
nor U682 (N_682,N_600,N_650);
nor U683 (N_683,N_643,N_619);
nand U684 (N_684,N_610,N_630);
and U685 (N_685,N_633,N_601);
nand U686 (N_686,N_626,N_632);
nor U687 (N_687,N_659,N_624);
nor U688 (N_688,N_638,N_612);
nor U689 (N_689,N_637,N_614);
nand U690 (N_690,N_653,N_641);
nor U691 (N_691,N_655,N_605);
and U692 (N_692,N_648,N_603);
nand U693 (N_693,N_651,N_605);
and U694 (N_694,N_607,N_652);
nor U695 (N_695,N_627,N_605);
nor U696 (N_696,N_625,N_657);
nand U697 (N_697,N_637,N_634);
xnor U698 (N_698,N_633,N_642);
or U699 (N_699,N_600,N_604);
and U700 (N_700,N_624,N_639);
and U701 (N_701,N_622,N_633);
nand U702 (N_702,N_609,N_637);
xnor U703 (N_703,N_651,N_656);
nand U704 (N_704,N_632,N_657);
and U705 (N_705,N_659,N_649);
xor U706 (N_706,N_639,N_636);
or U707 (N_707,N_630,N_608);
nand U708 (N_708,N_636,N_648);
or U709 (N_709,N_654,N_625);
nand U710 (N_710,N_610,N_618);
xor U711 (N_711,N_657,N_636);
xor U712 (N_712,N_600,N_621);
or U713 (N_713,N_644,N_633);
and U714 (N_714,N_639,N_603);
and U715 (N_715,N_618,N_608);
nor U716 (N_716,N_623,N_601);
nand U717 (N_717,N_610,N_656);
xnor U718 (N_718,N_651,N_644);
nor U719 (N_719,N_644,N_650);
and U720 (N_720,N_662,N_692);
and U721 (N_721,N_704,N_671);
and U722 (N_722,N_719,N_706);
or U723 (N_723,N_717,N_711);
nor U724 (N_724,N_707,N_665);
and U725 (N_725,N_673,N_660);
or U726 (N_726,N_674,N_712);
or U727 (N_727,N_693,N_705);
xor U728 (N_728,N_716,N_701);
or U729 (N_729,N_694,N_668);
nor U730 (N_730,N_684,N_714);
and U731 (N_731,N_715,N_679);
xor U732 (N_732,N_702,N_689);
and U733 (N_733,N_661,N_698);
nand U734 (N_734,N_699,N_680);
xnor U735 (N_735,N_663,N_664);
or U736 (N_736,N_696,N_675);
nor U737 (N_737,N_709,N_683);
nor U738 (N_738,N_672,N_667);
nand U739 (N_739,N_703,N_695);
nand U740 (N_740,N_697,N_691);
and U741 (N_741,N_682,N_677);
nor U742 (N_742,N_700,N_669);
nor U743 (N_743,N_676,N_687);
nor U744 (N_744,N_666,N_686);
xnor U745 (N_745,N_718,N_685);
and U746 (N_746,N_670,N_713);
nor U747 (N_747,N_710,N_690);
nand U748 (N_748,N_681,N_678);
and U749 (N_749,N_708,N_688);
nand U750 (N_750,N_666,N_685);
nor U751 (N_751,N_693,N_715);
and U752 (N_752,N_684,N_672);
nor U753 (N_753,N_677,N_697);
xor U754 (N_754,N_669,N_693);
or U755 (N_755,N_709,N_682);
nand U756 (N_756,N_663,N_713);
and U757 (N_757,N_708,N_664);
or U758 (N_758,N_712,N_710);
nor U759 (N_759,N_687,N_715);
or U760 (N_760,N_699,N_664);
or U761 (N_761,N_697,N_694);
nor U762 (N_762,N_671,N_719);
nor U763 (N_763,N_718,N_713);
nand U764 (N_764,N_696,N_719);
or U765 (N_765,N_714,N_665);
and U766 (N_766,N_691,N_695);
or U767 (N_767,N_706,N_717);
nand U768 (N_768,N_704,N_686);
nand U769 (N_769,N_661,N_702);
xor U770 (N_770,N_698,N_713);
nand U771 (N_771,N_704,N_662);
and U772 (N_772,N_715,N_664);
nand U773 (N_773,N_675,N_715);
and U774 (N_774,N_717,N_674);
nor U775 (N_775,N_685,N_696);
and U776 (N_776,N_694,N_675);
xnor U777 (N_777,N_717,N_661);
and U778 (N_778,N_715,N_683);
and U779 (N_779,N_679,N_717);
and U780 (N_780,N_735,N_725);
and U781 (N_781,N_758,N_763);
nand U782 (N_782,N_777,N_756);
xnor U783 (N_783,N_732,N_745);
nor U784 (N_784,N_742,N_775);
nor U785 (N_785,N_739,N_753);
or U786 (N_786,N_747,N_752);
and U787 (N_787,N_723,N_773);
nand U788 (N_788,N_761,N_743);
nand U789 (N_789,N_778,N_767);
nand U790 (N_790,N_764,N_749);
and U791 (N_791,N_754,N_731);
and U792 (N_792,N_741,N_728);
nand U793 (N_793,N_744,N_721);
nor U794 (N_794,N_730,N_760);
xnor U795 (N_795,N_727,N_755);
nor U796 (N_796,N_722,N_774);
or U797 (N_797,N_768,N_729);
nor U798 (N_798,N_733,N_772);
and U799 (N_799,N_737,N_776);
nand U800 (N_800,N_750,N_734);
or U801 (N_801,N_765,N_770);
nand U802 (N_802,N_720,N_736);
nand U803 (N_803,N_766,N_738);
or U804 (N_804,N_779,N_751);
or U805 (N_805,N_724,N_748);
nand U806 (N_806,N_740,N_726);
xnor U807 (N_807,N_746,N_757);
and U808 (N_808,N_771,N_762);
xor U809 (N_809,N_769,N_759);
and U810 (N_810,N_758,N_767);
xor U811 (N_811,N_733,N_778);
nor U812 (N_812,N_767,N_779);
nand U813 (N_813,N_725,N_779);
nand U814 (N_814,N_739,N_720);
or U815 (N_815,N_725,N_730);
and U816 (N_816,N_738,N_767);
or U817 (N_817,N_777,N_758);
or U818 (N_818,N_774,N_726);
xnor U819 (N_819,N_736,N_721);
nand U820 (N_820,N_749,N_740);
nand U821 (N_821,N_723,N_759);
or U822 (N_822,N_723,N_741);
nor U823 (N_823,N_751,N_742);
or U824 (N_824,N_772,N_755);
xor U825 (N_825,N_772,N_775);
or U826 (N_826,N_759,N_726);
xnor U827 (N_827,N_764,N_752);
nor U828 (N_828,N_726,N_775);
nand U829 (N_829,N_749,N_747);
nor U830 (N_830,N_739,N_738);
and U831 (N_831,N_761,N_728);
and U832 (N_832,N_747,N_734);
nor U833 (N_833,N_744,N_777);
nor U834 (N_834,N_742,N_767);
nor U835 (N_835,N_736,N_727);
nor U836 (N_836,N_739,N_737);
and U837 (N_837,N_736,N_760);
nand U838 (N_838,N_743,N_771);
xnor U839 (N_839,N_755,N_749);
and U840 (N_840,N_815,N_804);
nand U841 (N_841,N_798,N_839);
nand U842 (N_842,N_813,N_803);
nor U843 (N_843,N_817,N_793);
nor U844 (N_844,N_816,N_807);
and U845 (N_845,N_836,N_821);
nand U846 (N_846,N_837,N_830);
or U847 (N_847,N_799,N_824);
or U848 (N_848,N_805,N_806);
nor U849 (N_849,N_820,N_781);
nor U850 (N_850,N_838,N_818);
or U851 (N_851,N_812,N_795);
nor U852 (N_852,N_783,N_835);
nor U853 (N_853,N_789,N_810);
nor U854 (N_854,N_814,N_786);
nor U855 (N_855,N_833,N_823);
nor U856 (N_856,N_827,N_808);
nor U857 (N_857,N_819,N_829);
or U858 (N_858,N_831,N_788);
or U859 (N_859,N_826,N_834);
and U860 (N_860,N_796,N_787);
and U861 (N_861,N_785,N_801);
and U862 (N_862,N_797,N_800);
nor U863 (N_863,N_811,N_809);
nand U864 (N_864,N_794,N_790);
nor U865 (N_865,N_782,N_784);
nor U866 (N_866,N_822,N_780);
nand U867 (N_867,N_832,N_792);
nand U868 (N_868,N_802,N_825);
nand U869 (N_869,N_828,N_791);
nor U870 (N_870,N_817,N_783);
xor U871 (N_871,N_822,N_813);
nor U872 (N_872,N_815,N_780);
nand U873 (N_873,N_791,N_803);
nor U874 (N_874,N_783,N_792);
and U875 (N_875,N_783,N_834);
nor U876 (N_876,N_805,N_821);
nand U877 (N_877,N_791,N_786);
nor U878 (N_878,N_787,N_802);
and U879 (N_879,N_822,N_825);
nor U880 (N_880,N_813,N_815);
nand U881 (N_881,N_824,N_786);
and U882 (N_882,N_815,N_799);
nand U883 (N_883,N_820,N_831);
and U884 (N_884,N_807,N_805);
or U885 (N_885,N_837,N_811);
nor U886 (N_886,N_825,N_809);
nor U887 (N_887,N_797,N_827);
nand U888 (N_888,N_823,N_817);
and U889 (N_889,N_838,N_794);
and U890 (N_890,N_798,N_834);
nand U891 (N_891,N_815,N_784);
nor U892 (N_892,N_824,N_818);
and U893 (N_893,N_803,N_827);
or U894 (N_894,N_827,N_784);
and U895 (N_895,N_818,N_793);
nor U896 (N_896,N_829,N_798);
and U897 (N_897,N_838,N_783);
nand U898 (N_898,N_819,N_824);
nor U899 (N_899,N_818,N_804);
nor U900 (N_900,N_888,N_897);
and U901 (N_901,N_892,N_890);
nand U902 (N_902,N_850,N_849);
and U903 (N_903,N_841,N_894);
nor U904 (N_904,N_865,N_893);
nor U905 (N_905,N_876,N_861);
and U906 (N_906,N_870,N_868);
and U907 (N_907,N_884,N_895);
nor U908 (N_908,N_869,N_866);
nand U909 (N_909,N_856,N_889);
and U910 (N_910,N_844,N_855);
nor U911 (N_911,N_899,N_898);
and U912 (N_912,N_879,N_872);
or U913 (N_913,N_880,N_896);
nor U914 (N_914,N_886,N_843);
xor U915 (N_915,N_848,N_858);
or U916 (N_916,N_840,N_878);
xnor U917 (N_917,N_873,N_882);
or U918 (N_918,N_853,N_860);
or U919 (N_919,N_864,N_871);
nand U920 (N_920,N_854,N_847);
nand U921 (N_921,N_877,N_862);
nand U922 (N_922,N_887,N_883);
and U923 (N_923,N_875,N_845);
xor U924 (N_924,N_859,N_863);
nor U925 (N_925,N_857,N_891);
nor U926 (N_926,N_842,N_867);
nand U927 (N_927,N_846,N_885);
and U928 (N_928,N_851,N_852);
nand U929 (N_929,N_881,N_874);
or U930 (N_930,N_891,N_875);
xor U931 (N_931,N_879,N_868);
xnor U932 (N_932,N_872,N_861);
nand U933 (N_933,N_877,N_885);
nand U934 (N_934,N_844,N_847);
and U935 (N_935,N_877,N_886);
and U936 (N_936,N_880,N_841);
and U937 (N_937,N_842,N_875);
nand U938 (N_938,N_870,N_898);
nand U939 (N_939,N_859,N_894);
nor U940 (N_940,N_898,N_852);
or U941 (N_941,N_889,N_877);
and U942 (N_942,N_841,N_874);
or U943 (N_943,N_879,N_858);
nand U944 (N_944,N_893,N_847);
xnor U945 (N_945,N_869,N_879);
nand U946 (N_946,N_898,N_845);
nor U947 (N_947,N_852,N_840);
and U948 (N_948,N_892,N_851);
nand U949 (N_949,N_864,N_868);
nor U950 (N_950,N_849,N_864);
xor U951 (N_951,N_862,N_874);
nand U952 (N_952,N_881,N_847);
nor U953 (N_953,N_869,N_843);
nor U954 (N_954,N_880,N_859);
and U955 (N_955,N_867,N_843);
and U956 (N_956,N_853,N_897);
or U957 (N_957,N_889,N_876);
or U958 (N_958,N_840,N_845);
nand U959 (N_959,N_860,N_868);
or U960 (N_960,N_947,N_930);
and U961 (N_961,N_916,N_920);
nand U962 (N_962,N_942,N_908);
or U963 (N_963,N_935,N_919);
nor U964 (N_964,N_936,N_925);
nand U965 (N_965,N_938,N_949);
or U966 (N_966,N_945,N_909);
and U967 (N_967,N_957,N_950);
xor U968 (N_968,N_922,N_912);
or U969 (N_969,N_928,N_927);
nor U970 (N_970,N_929,N_933);
and U971 (N_971,N_924,N_940);
nand U972 (N_972,N_900,N_910);
or U973 (N_973,N_955,N_931);
nor U974 (N_974,N_943,N_953);
xor U975 (N_975,N_913,N_923);
nand U976 (N_976,N_952,N_956);
nor U977 (N_977,N_905,N_918);
and U978 (N_978,N_917,N_941);
nand U979 (N_979,N_903,N_948);
nand U980 (N_980,N_901,N_906);
nand U981 (N_981,N_904,N_911);
and U982 (N_982,N_939,N_946);
or U983 (N_983,N_937,N_915);
and U984 (N_984,N_951,N_902);
nand U985 (N_985,N_926,N_934);
or U986 (N_986,N_954,N_958);
and U987 (N_987,N_907,N_944);
nand U988 (N_988,N_959,N_914);
nand U989 (N_989,N_932,N_921);
nor U990 (N_990,N_942,N_943);
nor U991 (N_991,N_941,N_937);
and U992 (N_992,N_926,N_959);
or U993 (N_993,N_903,N_942);
or U994 (N_994,N_933,N_932);
nand U995 (N_995,N_934,N_908);
nor U996 (N_996,N_902,N_956);
xnor U997 (N_997,N_941,N_907);
or U998 (N_998,N_949,N_945);
or U999 (N_999,N_901,N_904);
nor U1000 (N_1000,N_936,N_949);
and U1001 (N_1001,N_944,N_959);
or U1002 (N_1002,N_947,N_939);
or U1003 (N_1003,N_929,N_935);
nand U1004 (N_1004,N_902,N_954);
or U1005 (N_1005,N_920,N_952);
xor U1006 (N_1006,N_954,N_927);
nand U1007 (N_1007,N_919,N_934);
nor U1008 (N_1008,N_956,N_938);
or U1009 (N_1009,N_936,N_902);
or U1010 (N_1010,N_912,N_953);
nand U1011 (N_1011,N_958,N_938);
or U1012 (N_1012,N_906,N_955);
nor U1013 (N_1013,N_934,N_910);
xor U1014 (N_1014,N_920,N_936);
nand U1015 (N_1015,N_943,N_957);
nor U1016 (N_1016,N_950,N_917);
nand U1017 (N_1017,N_940,N_912);
nor U1018 (N_1018,N_913,N_934);
nor U1019 (N_1019,N_912,N_927);
nand U1020 (N_1020,N_960,N_973);
xnor U1021 (N_1021,N_979,N_1016);
nand U1022 (N_1022,N_968,N_976);
and U1023 (N_1023,N_985,N_999);
nand U1024 (N_1024,N_1012,N_998);
nor U1025 (N_1025,N_1004,N_1005);
nor U1026 (N_1026,N_972,N_975);
nor U1027 (N_1027,N_1019,N_1009);
nand U1028 (N_1028,N_984,N_1018);
nand U1029 (N_1029,N_980,N_969);
or U1030 (N_1030,N_987,N_978);
or U1031 (N_1031,N_964,N_1007);
and U1032 (N_1032,N_982,N_1003);
nand U1033 (N_1033,N_1010,N_970);
nand U1034 (N_1034,N_986,N_1008);
or U1035 (N_1035,N_997,N_1002);
or U1036 (N_1036,N_992,N_962);
nand U1037 (N_1037,N_961,N_1014);
nor U1038 (N_1038,N_963,N_974);
or U1039 (N_1039,N_989,N_971);
or U1040 (N_1040,N_966,N_1011);
nor U1041 (N_1041,N_1000,N_988);
or U1042 (N_1042,N_990,N_983);
nand U1043 (N_1043,N_995,N_1013);
nand U1044 (N_1044,N_1015,N_965);
nand U1045 (N_1045,N_996,N_993);
or U1046 (N_1046,N_1017,N_981);
or U1047 (N_1047,N_1001,N_1006);
or U1048 (N_1048,N_991,N_967);
nand U1049 (N_1049,N_994,N_977);
xor U1050 (N_1050,N_982,N_994);
or U1051 (N_1051,N_1003,N_1010);
and U1052 (N_1052,N_997,N_1015);
nand U1053 (N_1053,N_975,N_1012);
nor U1054 (N_1054,N_962,N_990);
nand U1055 (N_1055,N_1018,N_967);
or U1056 (N_1056,N_985,N_969);
and U1057 (N_1057,N_972,N_1011);
nor U1058 (N_1058,N_1014,N_987);
nor U1059 (N_1059,N_991,N_1017);
or U1060 (N_1060,N_1018,N_988);
nor U1061 (N_1061,N_967,N_1017);
or U1062 (N_1062,N_971,N_987);
nor U1063 (N_1063,N_995,N_1009);
nor U1064 (N_1064,N_962,N_1007);
nor U1065 (N_1065,N_984,N_1011);
and U1066 (N_1066,N_1006,N_965);
nor U1067 (N_1067,N_1002,N_1012);
nand U1068 (N_1068,N_998,N_972);
or U1069 (N_1069,N_996,N_975);
nand U1070 (N_1070,N_968,N_1012);
and U1071 (N_1071,N_1001,N_1004);
and U1072 (N_1072,N_986,N_979);
nand U1073 (N_1073,N_966,N_1013);
or U1074 (N_1074,N_968,N_977);
nor U1075 (N_1075,N_967,N_990);
or U1076 (N_1076,N_999,N_986);
nand U1077 (N_1077,N_989,N_996);
nor U1078 (N_1078,N_1004,N_1003);
and U1079 (N_1079,N_1005,N_995);
or U1080 (N_1080,N_1070,N_1025);
and U1081 (N_1081,N_1022,N_1057);
nand U1082 (N_1082,N_1024,N_1056);
nor U1083 (N_1083,N_1058,N_1061);
and U1084 (N_1084,N_1045,N_1026);
nand U1085 (N_1085,N_1073,N_1046);
or U1086 (N_1086,N_1054,N_1069);
nor U1087 (N_1087,N_1079,N_1072);
and U1088 (N_1088,N_1030,N_1044);
nor U1089 (N_1089,N_1032,N_1075);
nor U1090 (N_1090,N_1020,N_1066);
and U1091 (N_1091,N_1071,N_1034);
or U1092 (N_1092,N_1021,N_1041);
nand U1093 (N_1093,N_1050,N_1047);
nor U1094 (N_1094,N_1076,N_1078);
nand U1095 (N_1095,N_1065,N_1059);
or U1096 (N_1096,N_1029,N_1074);
or U1097 (N_1097,N_1067,N_1028);
or U1098 (N_1098,N_1064,N_1077);
nand U1099 (N_1099,N_1033,N_1039);
nand U1100 (N_1100,N_1051,N_1031);
or U1101 (N_1101,N_1027,N_1063);
nand U1102 (N_1102,N_1042,N_1037);
nand U1103 (N_1103,N_1036,N_1052);
and U1104 (N_1104,N_1043,N_1038);
and U1105 (N_1105,N_1053,N_1049);
nor U1106 (N_1106,N_1023,N_1062);
or U1107 (N_1107,N_1035,N_1055);
nor U1108 (N_1108,N_1040,N_1048);
nor U1109 (N_1109,N_1068,N_1060);
and U1110 (N_1110,N_1034,N_1041);
and U1111 (N_1111,N_1058,N_1051);
nor U1112 (N_1112,N_1050,N_1035);
nor U1113 (N_1113,N_1067,N_1065);
or U1114 (N_1114,N_1064,N_1050);
nand U1115 (N_1115,N_1054,N_1022);
nand U1116 (N_1116,N_1040,N_1021);
nor U1117 (N_1117,N_1027,N_1057);
or U1118 (N_1118,N_1042,N_1057);
or U1119 (N_1119,N_1033,N_1063);
or U1120 (N_1120,N_1058,N_1046);
and U1121 (N_1121,N_1062,N_1077);
nand U1122 (N_1122,N_1075,N_1030);
or U1123 (N_1123,N_1076,N_1038);
nor U1124 (N_1124,N_1031,N_1076);
xor U1125 (N_1125,N_1044,N_1026);
or U1126 (N_1126,N_1041,N_1062);
nor U1127 (N_1127,N_1034,N_1069);
or U1128 (N_1128,N_1039,N_1061);
nor U1129 (N_1129,N_1059,N_1075);
nor U1130 (N_1130,N_1068,N_1053);
nor U1131 (N_1131,N_1043,N_1076);
nor U1132 (N_1132,N_1040,N_1070);
and U1133 (N_1133,N_1068,N_1073);
and U1134 (N_1134,N_1068,N_1077);
or U1135 (N_1135,N_1028,N_1078);
nor U1136 (N_1136,N_1039,N_1036);
nand U1137 (N_1137,N_1073,N_1069);
nor U1138 (N_1138,N_1053,N_1025);
and U1139 (N_1139,N_1067,N_1042);
nor U1140 (N_1140,N_1112,N_1088);
nor U1141 (N_1141,N_1083,N_1102);
nor U1142 (N_1142,N_1087,N_1110);
nand U1143 (N_1143,N_1099,N_1132);
nor U1144 (N_1144,N_1126,N_1101);
and U1145 (N_1145,N_1098,N_1127);
nand U1146 (N_1146,N_1084,N_1085);
and U1147 (N_1147,N_1111,N_1121);
and U1148 (N_1148,N_1113,N_1119);
or U1149 (N_1149,N_1138,N_1122);
nand U1150 (N_1150,N_1104,N_1134);
nand U1151 (N_1151,N_1139,N_1115);
and U1152 (N_1152,N_1089,N_1136);
and U1153 (N_1153,N_1096,N_1107);
nand U1154 (N_1154,N_1118,N_1124);
or U1155 (N_1155,N_1091,N_1128);
nand U1156 (N_1156,N_1100,N_1106);
nor U1157 (N_1157,N_1086,N_1133);
nor U1158 (N_1158,N_1109,N_1082);
or U1159 (N_1159,N_1105,N_1093);
nand U1160 (N_1160,N_1080,N_1114);
and U1161 (N_1161,N_1103,N_1125);
and U1162 (N_1162,N_1117,N_1092);
or U1163 (N_1163,N_1108,N_1120);
nor U1164 (N_1164,N_1090,N_1116);
and U1165 (N_1165,N_1081,N_1137);
and U1166 (N_1166,N_1130,N_1094);
nor U1167 (N_1167,N_1135,N_1123);
nand U1168 (N_1168,N_1095,N_1129);
nand U1169 (N_1169,N_1131,N_1097);
or U1170 (N_1170,N_1130,N_1116);
nand U1171 (N_1171,N_1087,N_1106);
nand U1172 (N_1172,N_1082,N_1137);
nand U1173 (N_1173,N_1117,N_1084);
nor U1174 (N_1174,N_1133,N_1116);
and U1175 (N_1175,N_1131,N_1104);
xnor U1176 (N_1176,N_1106,N_1137);
or U1177 (N_1177,N_1130,N_1124);
and U1178 (N_1178,N_1103,N_1129);
xnor U1179 (N_1179,N_1081,N_1112);
or U1180 (N_1180,N_1112,N_1096);
nand U1181 (N_1181,N_1119,N_1124);
nand U1182 (N_1182,N_1134,N_1118);
nor U1183 (N_1183,N_1106,N_1108);
or U1184 (N_1184,N_1100,N_1096);
xor U1185 (N_1185,N_1127,N_1093);
nand U1186 (N_1186,N_1130,N_1125);
nor U1187 (N_1187,N_1126,N_1139);
nor U1188 (N_1188,N_1093,N_1104);
or U1189 (N_1189,N_1133,N_1120);
or U1190 (N_1190,N_1096,N_1111);
or U1191 (N_1191,N_1114,N_1088);
or U1192 (N_1192,N_1090,N_1117);
or U1193 (N_1193,N_1120,N_1131);
and U1194 (N_1194,N_1117,N_1115);
nand U1195 (N_1195,N_1136,N_1080);
and U1196 (N_1196,N_1138,N_1132);
or U1197 (N_1197,N_1081,N_1095);
nor U1198 (N_1198,N_1086,N_1091);
or U1199 (N_1199,N_1117,N_1113);
and U1200 (N_1200,N_1163,N_1158);
and U1201 (N_1201,N_1186,N_1181);
or U1202 (N_1202,N_1189,N_1154);
nand U1203 (N_1203,N_1144,N_1185);
nor U1204 (N_1204,N_1182,N_1198);
and U1205 (N_1205,N_1153,N_1150);
nor U1206 (N_1206,N_1190,N_1193);
and U1207 (N_1207,N_1180,N_1177);
or U1208 (N_1208,N_1197,N_1159);
nand U1209 (N_1209,N_1142,N_1143);
xor U1210 (N_1210,N_1162,N_1191);
and U1211 (N_1211,N_1151,N_1169);
nand U1212 (N_1212,N_1161,N_1146);
and U1213 (N_1213,N_1164,N_1192);
nand U1214 (N_1214,N_1156,N_1148);
or U1215 (N_1215,N_1167,N_1178);
nand U1216 (N_1216,N_1140,N_1195);
or U1217 (N_1217,N_1196,N_1176);
xor U1218 (N_1218,N_1145,N_1149);
nor U1219 (N_1219,N_1173,N_1187);
and U1220 (N_1220,N_1184,N_1160);
or U1221 (N_1221,N_1147,N_1194);
xor U1222 (N_1222,N_1157,N_1171);
and U1223 (N_1223,N_1175,N_1174);
nand U1224 (N_1224,N_1179,N_1170);
nand U1225 (N_1225,N_1166,N_1183);
nand U1226 (N_1226,N_1188,N_1152);
nand U1227 (N_1227,N_1155,N_1141);
xor U1228 (N_1228,N_1168,N_1172);
or U1229 (N_1229,N_1165,N_1199);
or U1230 (N_1230,N_1193,N_1152);
or U1231 (N_1231,N_1185,N_1142);
and U1232 (N_1232,N_1146,N_1185);
xor U1233 (N_1233,N_1182,N_1143);
xnor U1234 (N_1234,N_1159,N_1151);
xor U1235 (N_1235,N_1194,N_1197);
and U1236 (N_1236,N_1175,N_1164);
or U1237 (N_1237,N_1181,N_1179);
nor U1238 (N_1238,N_1157,N_1149);
nor U1239 (N_1239,N_1192,N_1189);
or U1240 (N_1240,N_1177,N_1190);
and U1241 (N_1241,N_1146,N_1183);
nor U1242 (N_1242,N_1188,N_1186);
nor U1243 (N_1243,N_1165,N_1171);
or U1244 (N_1244,N_1170,N_1166);
nand U1245 (N_1245,N_1156,N_1162);
or U1246 (N_1246,N_1146,N_1173);
and U1247 (N_1247,N_1160,N_1151);
and U1248 (N_1248,N_1160,N_1150);
xor U1249 (N_1249,N_1163,N_1155);
and U1250 (N_1250,N_1152,N_1144);
nand U1251 (N_1251,N_1148,N_1188);
nand U1252 (N_1252,N_1149,N_1153);
nand U1253 (N_1253,N_1168,N_1141);
or U1254 (N_1254,N_1151,N_1158);
and U1255 (N_1255,N_1151,N_1187);
nand U1256 (N_1256,N_1154,N_1194);
nand U1257 (N_1257,N_1195,N_1163);
and U1258 (N_1258,N_1195,N_1197);
nor U1259 (N_1259,N_1198,N_1192);
nand U1260 (N_1260,N_1247,N_1216);
nor U1261 (N_1261,N_1223,N_1259);
nand U1262 (N_1262,N_1248,N_1206);
nor U1263 (N_1263,N_1200,N_1239);
nand U1264 (N_1264,N_1251,N_1249);
nor U1265 (N_1265,N_1246,N_1232);
nor U1266 (N_1266,N_1214,N_1225);
or U1267 (N_1267,N_1221,N_1213);
or U1268 (N_1268,N_1245,N_1215);
nor U1269 (N_1269,N_1231,N_1236);
or U1270 (N_1270,N_1219,N_1252);
nor U1271 (N_1271,N_1258,N_1233);
xor U1272 (N_1272,N_1241,N_1238);
or U1273 (N_1273,N_1255,N_1229);
nor U1274 (N_1274,N_1242,N_1227);
xnor U1275 (N_1275,N_1220,N_1240);
and U1276 (N_1276,N_1237,N_1234);
nand U1277 (N_1277,N_1257,N_1235);
nor U1278 (N_1278,N_1209,N_1210);
nor U1279 (N_1279,N_1212,N_1230);
and U1280 (N_1280,N_1243,N_1254);
nand U1281 (N_1281,N_1201,N_1211);
xor U1282 (N_1282,N_1250,N_1217);
or U1283 (N_1283,N_1202,N_1205);
or U1284 (N_1284,N_1222,N_1256);
or U1285 (N_1285,N_1228,N_1218);
or U1286 (N_1286,N_1224,N_1207);
nand U1287 (N_1287,N_1226,N_1253);
and U1288 (N_1288,N_1204,N_1203);
nand U1289 (N_1289,N_1208,N_1244);
nand U1290 (N_1290,N_1254,N_1241);
nor U1291 (N_1291,N_1252,N_1202);
and U1292 (N_1292,N_1218,N_1235);
or U1293 (N_1293,N_1258,N_1200);
nor U1294 (N_1294,N_1246,N_1217);
xnor U1295 (N_1295,N_1209,N_1241);
nand U1296 (N_1296,N_1243,N_1257);
nor U1297 (N_1297,N_1209,N_1213);
and U1298 (N_1298,N_1200,N_1201);
xor U1299 (N_1299,N_1255,N_1235);
nor U1300 (N_1300,N_1219,N_1254);
or U1301 (N_1301,N_1229,N_1213);
nand U1302 (N_1302,N_1219,N_1250);
and U1303 (N_1303,N_1233,N_1200);
and U1304 (N_1304,N_1239,N_1233);
and U1305 (N_1305,N_1235,N_1256);
or U1306 (N_1306,N_1220,N_1203);
nor U1307 (N_1307,N_1202,N_1251);
and U1308 (N_1308,N_1255,N_1203);
or U1309 (N_1309,N_1252,N_1251);
nand U1310 (N_1310,N_1221,N_1223);
and U1311 (N_1311,N_1214,N_1211);
or U1312 (N_1312,N_1213,N_1220);
nor U1313 (N_1313,N_1206,N_1233);
xor U1314 (N_1314,N_1226,N_1228);
nand U1315 (N_1315,N_1239,N_1215);
nand U1316 (N_1316,N_1237,N_1244);
nor U1317 (N_1317,N_1250,N_1240);
or U1318 (N_1318,N_1200,N_1203);
nor U1319 (N_1319,N_1226,N_1257);
nor U1320 (N_1320,N_1309,N_1290);
or U1321 (N_1321,N_1289,N_1285);
xnor U1322 (N_1322,N_1312,N_1276);
and U1323 (N_1323,N_1297,N_1270);
nand U1324 (N_1324,N_1306,N_1300);
nand U1325 (N_1325,N_1284,N_1286);
or U1326 (N_1326,N_1272,N_1298);
and U1327 (N_1327,N_1265,N_1269);
nor U1328 (N_1328,N_1310,N_1317);
or U1329 (N_1329,N_1274,N_1319);
and U1330 (N_1330,N_1287,N_1278);
nor U1331 (N_1331,N_1275,N_1311);
or U1332 (N_1332,N_1302,N_1308);
and U1333 (N_1333,N_1260,N_1296);
and U1334 (N_1334,N_1295,N_1261);
or U1335 (N_1335,N_1262,N_1316);
and U1336 (N_1336,N_1273,N_1283);
nor U1337 (N_1337,N_1280,N_1288);
nor U1338 (N_1338,N_1271,N_1313);
and U1339 (N_1339,N_1277,N_1282);
or U1340 (N_1340,N_1305,N_1279);
or U1341 (N_1341,N_1314,N_1266);
and U1342 (N_1342,N_1315,N_1268);
or U1343 (N_1343,N_1299,N_1293);
nor U1344 (N_1344,N_1307,N_1264);
nand U1345 (N_1345,N_1304,N_1301);
nor U1346 (N_1346,N_1263,N_1267);
or U1347 (N_1347,N_1318,N_1281);
or U1348 (N_1348,N_1303,N_1291);
nand U1349 (N_1349,N_1292,N_1294);
or U1350 (N_1350,N_1313,N_1288);
nor U1351 (N_1351,N_1270,N_1283);
and U1352 (N_1352,N_1286,N_1310);
and U1353 (N_1353,N_1294,N_1290);
nor U1354 (N_1354,N_1263,N_1262);
xnor U1355 (N_1355,N_1284,N_1290);
and U1356 (N_1356,N_1274,N_1278);
and U1357 (N_1357,N_1304,N_1292);
or U1358 (N_1358,N_1301,N_1297);
nand U1359 (N_1359,N_1267,N_1302);
or U1360 (N_1360,N_1297,N_1298);
nand U1361 (N_1361,N_1306,N_1299);
nand U1362 (N_1362,N_1307,N_1286);
xnor U1363 (N_1363,N_1284,N_1265);
and U1364 (N_1364,N_1271,N_1263);
nor U1365 (N_1365,N_1294,N_1261);
nor U1366 (N_1366,N_1313,N_1317);
and U1367 (N_1367,N_1281,N_1272);
nor U1368 (N_1368,N_1302,N_1303);
xor U1369 (N_1369,N_1305,N_1299);
nor U1370 (N_1370,N_1270,N_1281);
nand U1371 (N_1371,N_1282,N_1302);
nor U1372 (N_1372,N_1268,N_1267);
nand U1373 (N_1373,N_1309,N_1287);
xor U1374 (N_1374,N_1295,N_1316);
or U1375 (N_1375,N_1276,N_1278);
nand U1376 (N_1376,N_1280,N_1293);
nor U1377 (N_1377,N_1273,N_1278);
or U1378 (N_1378,N_1274,N_1314);
xnor U1379 (N_1379,N_1284,N_1300);
or U1380 (N_1380,N_1328,N_1376);
or U1381 (N_1381,N_1334,N_1368);
nor U1382 (N_1382,N_1340,N_1324);
xnor U1383 (N_1383,N_1350,N_1369);
xor U1384 (N_1384,N_1373,N_1338);
nor U1385 (N_1385,N_1372,N_1362);
nor U1386 (N_1386,N_1371,N_1351);
xor U1387 (N_1387,N_1370,N_1335);
and U1388 (N_1388,N_1333,N_1367);
or U1389 (N_1389,N_1323,N_1329);
or U1390 (N_1390,N_1360,N_1327);
or U1391 (N_1391,N_1375,N_1343);
and U1392 (N_1392,N_1353,N_1344);
xnor U1393 (N_1393,N_1357,N_1341);
or U1394 (N_1394,N_1363,N_1352);
or U1395 (N_1395,N_1349,N_1379);
nand U1396 (N_1396,N_1374,N_1361);
nand U1397 (N_1397,N_1345,N_1354);
or U1398 (N_1398,N_1342,N_1347);
nor U1399 (N_1399,N_1378,N_1326);
nand U1400 (N_1400,N_1331,N_1332);
nand U1401 (N_1401,N_1339,N_1356);
or U1402 (N_1402,N_1320,N_1364);
and U1403 (N_1403,N_1359,N_1348);
nand U1404 (N_1404,N_1325,N_1337);
nand U1405 (N_1405,N_1366,N_1336);
nand U1406 (N_1406,N_1377,N_1322);
nand U1407 (N_1407,N_1355,N_1330);
and U1408 (N_1408,N_1365,N_1346);
and U1409 (N_1409,N_1321,N_1358);
nand U1410 (N_1410,N_1326,N_1336);
nand U1411 (N_1411,N_1353,N_1327);
nor U1412 (N_1412,N_1322,N_1375);
nand U1413 (N_1413,N_1364,N_1373);
or U1414 (N_1414,N_1329,N_1332);
nand U1415 (N_1415,N_1378,N_1323);
nor U1416 (N_1416,N_1368,N_1379);
or U1417 (N_1417,N_1342,N_1355);
or U1418 (N_1418,N_1329,N_1339);
nor U1419 (N_1419,N_1321,N_1327);
or U1420 (N_1420,N_1348,N_1354);
nand U1421 (N_1421,N_1331,N_1344);
nand U1422 (N_1422,N_1330,N_1363);
or U1423 (N_1423,N_1326,N_1347);
nand U1424 (N_1424,N_1371,N_1320);
nor U1425 (N_1425,N_1342,N_1357);
xor U1426 (N_1426,N_1322,N_1358);
and U1427 (N_1427,N_1340,N_1344);
nor U1428 (N_1428,N_1357,N_1359);
xor U1429 (N_1429,N_1362,N_1379);
nand U1430 (N_1430,N_1362,N_1357);
or U1431 (N_1431,N_1367,N_1348);
nor U1432 (N_1432,N_1320,N_1367);
or U1433 (N_1433,N_1328,N_1377);
nand U1434 (N_1434,N_1352,N_1325);
nor U1435 (N_1435,N_1342,N_1362);
or U1436 (N_1436,N_1368,N_1357);
and U1437 (N_1437,N_1378,N_1332);
nand U1438 (N_1438,N_1354,N_1366);
and U1439 (N_1439,N_1374,N_1344);
nor U1440 (N_1440,N_1399,N_1413);
nand U1441 (N_1441,N_1419,N_1432);
or U1442 (N_1442,N_1392,N_1393);
or U1443 (N_1443,N_1404,N_1407);
or U1444 (N_1444,N_1424,N_1434);
nand U1445 (N_1445,N_1381,N_1385);
and U1446 (N_1446,N_1389,N_1402);
nand U1447 (N_1447,N_1390,N_1406);
xor U1448 (N_1448,N_1384,N_1430);
xnor U1449 (N_1449,N_1433,N_1423);
nand U1450 (N_1450,N_1435,N_1426);
nand U1451 (N_1451,N_1386,N_1400);
and U1452 (N_1452,N_1431,N_1428);
and U1453 (N_1453,N_1437,N_1417);
or U1454 (N_1454,N_1387,N_1425);
nand U1455 (N_1455,N_1411,N_1422);
nand U1456 (N_1456,N_1403,N_1401);
or U1457 (N_1457,N_1410,N_1380);
nor U1458 (N_1458,N_1412,N_1418);
and U1459 (N_1459,N_1439,N_1398);
nand U1460 (N_1460,N_1395,N_1421);
nand U1461 (N_1461,N_1415,N_1394);
nor U1462 (N_1462,N_1409,N_1388);
or U1463 (N_1463,N_1416,N_1414);
nand U1464 (N_1464,N_1383,N_1438);
nand U1465 (N_1465,N_1397,N_1405);
nand U1466 (N_1466,N_1391,N_1396);
and U1467 (N_1467,N_1436,N_1382);
and U1468 (N_1468,N_1420,N_1408);
nor U1469 (N_1469,N_1429,N_1427);
nor U1470 (N_1470,N_1432,N_1402);
nand U1471 (N_1471,N_1410,N_1385);
or U1472 (N_1472,N_1412,N_1391);
and U1473 (N_1473,N_1404,N_1416);
or U1474 (N_1474,N_1386,N_1411);
or U1475 (N_1475,N_1399,N_1398);
and U1476 (N_1476,N_1384,N_1435);
or U1477 (N_1477,N_1400,N_1430);
nand U1478 (N_1478,N_1434,N_1385);
or U1479 (N_1479,N_1392,N_1417);
or U1480 (N_1480,N_1387,N_1430);
nor U1481 (N_1481,N_1383,N_1409);
or U1482 (N_1482,N_1419,N_1381);
xnor U1483 (N_1483,N_1406,N_1401);
nor U1484 (N_1484,N_1414,N_1424);
xor U1485 (N_1485,N_1415,N_1431);
nor U1486 (N_1486,N_1383,N_1408);
or U1487 (N_1487,N_1431,N_1411);
or U1488 (N_1488,N_1420,N_1394);
nor U1489 (N_1489,N_1409,N_1424);
or U1490 (N_1490,N_1404,N_1417);
or U1491 (N_1491,N_1423,N_1429);
and U1492 (N_1492,N_1411,N_1403);
and U1493 (N_1493,N_1400,N_1385);
or U1494 (N_1494,N_1431,N_1438);
xor U1495 (N_1495,N_1439,N_1433);
and U1496 (N_1496,N_1427,N_1415);
nor U1497 (N_1497,N_1425,N_1404);
or U1498 (N_1498,N_1433,N_1381);
nand U1499 (N_1499,N_1413,N_1435);
nand U1500 (N_1500,N_1446,N_1448);
nor U1501 (N_1501,N_1454,N_1467);
nand U1502 (N_1502,N_1442,N_1485);
and U1503 (N_1503,N_1494,N_1447);
nor U1504 (N_1504,N_1498,N_1486);
xnor U1505 (N_1505,N_1455,N_1470);
or U1506 (N_1506,N_1495,N_1443);
nand U1507 (N_1507,N_1474,N_1450);
or U1508 (N_1508,N_1462,N_1461);
or U1509 (N_1509,N_1457,N_1483);
nor U1510 (N_1510,N_1466,N_1453);
or U1511 (N_1511,N_1490,N_1449);
nor U1512 (N_1512,N_1479,N_1477);
nand U1513 (N_1513,N_1460,N_1484);
nand U1514 (N_1514,N_1444,N_1459);
and U1515 (N_1515,N_1499,N_1458);
or U1516 (N_1516,N_1496,N_1497);
or U1517 (N_1517,N_1491,N_1464);
and U1518 (N_1518,N_1487,N_1451);
nor U1519 (N_1519,N_1465,N_1469);
and U1520 (N_1520,N_1478,N_1472);
nand U1521 (N_1521,N_1493,N_1463);
or U1522 (N_1522,N_1452,N_1475);
or U1523 (N_1523,N_1488,N_1440);
nor U1524 (N_1524,N_1456,N_1476);
or U1525 (N_1525,N_1482,N_1468);
or U1526 (N_1526,N_1471,N_1441);
nand U1527 (N_1527,N_1473,N_1445);
nand U1528 (N_1528,N_1480,N_1489);
nand U1529 (N_1529,N_1481,N_1492);
or U1530 (N_1530,N_1482,N_1480);
nand U1531 (N_1531,N_1462,N_1460);
nor U1532 (N_1532,N_1452,N_1454);
or U1533 (N_1533,N_1453,N_1489);
and U1534 (N_1534,N_1489,N_1456);
or U1535 (N_1535,N_1488,N_1487);
and U1536 (N_1536,N_1443,N_1445);
nand U1537 (N_1537,N_1466,N_1497);
and U1538 (N_1538,N_1455,N_1482);
nand U1539 (N_1539,N_1473,N_1495);
nand U1540 (N_1540,N_1494,N_1442);
and U1541 (N_1541,N_1448,N_1499);
and U1542 (N_1542,N_1458,N_1461);
nand U1543 (N_1543,N_1472,N_1495);
and U1544 (N_1544,N_1448,N_1455);
or U1545 (N_1545,N_1498,N_1485);
nor U1546 (N_1546,N_1448,N_1471);
nor U1547 (N_1547,N_1492,N_1483);
and U1548 (N_1548,N_1497,N_1478);
nor U1549 (N_1549,N_1461,N_1457);
nand U1550 (N_1550,N_1454,N_1461);
and U1551 (N_1551,N_1465,N_1475);
and U1552 (N_1552,N_1459,N_1495);
xor U1553 (N_1553,N_1444,N_1498);
nor U1554 (N_1554,N_1484,N_1454);
or U1555 (N_1555,N_1473,N_1472);
nand U1556 (N_1556,N_1463,N_1454);
xnor U1557 (N_1557,N_1486,N_1494);
nand U1558 (N_1558,N_1483,N_1466);
nand U1559 (N_1559,N_1478,N_1451);
or U1560 (N_1560,N_1552,N_1507);
or U1561 (N_1561,N_1515,N_1511);
nor U1562 (N_1562,N_1518,N_1537);
and U1563 (N_1563,N_1516,N_1532);
and U1564 (N_1564,N_1544,N_1557);
nor U1565 (N_1565,N_1539,N_1536);
nor U1566 (N_1566,N_1509,N_1519);
nor U1567 (N_1567,N_1505,N_1534);
and U1568 (N_1568,N_1549,N_1500);
nor U1569 (N_1569,N_1541,N_1550);
nand U1570 (N_1570,N_1521,N_1506);
xor U1571 (N_1571,N_1554,N_1502);
nor U1572 (N_1572,N_1528,N_1530);
or U1573 (N_1573,N_1526,N_1543);
xor U1574 (N_1574,N_1547,N_1546);
and U1575 (N_1575,N_1520,N_1517);
and U1576 (N_1576,N_1508,N_1538);
and U1577 (N_1577,N_1553,N_1535);
nor U1578 (N_1578,N_1551,N_1527);
nor U1579 (N_1579,N_1533,N_1531);
xnor U1580 (N_1580,N_1556,N_1513);
or U1581 (N_1581,N_1503,N_1542);
and U1582 (N_1582,N_1523,N_1559);
and U1583 (N_1583,N_1545,N_1524);
or U1584 (N_1584,N_1529,N_1522);
nand U1585 (N_1585,N_1510,N_1514);
and U1586 (N_1586,N_1501,N_1512);
nand U1587 (N_1587,N_1548,N_1540);
nor U1588 (N_1588,N_1525,N_1555);
nor U1589 (N_1589,N_1504,N_1558);
xnor U1590 (N_1590,N_1537,N_1542);
nand U1591 (N_1591,N_1534,N_1541);
nor U1592 (N_1592,N_1509,N_1549);
and U1593 (N_1593,N_1554,N_1535);
nor U1594 (N_1594,N_1525,N_1514);
or U1595 (N_1595,N_1500,N_1514);
and U1596 (N_1596,N_1536,N_1522);
or U1597 (N_1597,N_1552,N_1532);
xnor U1598 (N_1598,N_1506,N_1517);
xnor U1599 (N_1599,N_1523,N_1524);
nor U1600 (N_1600,N_1542,N_1501);
nand U1601 (N_1601,N_1520,N_1518);
or U1602 (N_1602,N_1544,N_1532);
nand U1603 (N_1603,N_1535,N_1525);
or U1604 (N_1604,N_1511,N_1549);
nand U1605 (N_1605,N_1507,N_1556);
nor U1606 (N_1606,N_1508,N_1550);
nor U1607 (N_1607,N_1512,N_1519);
or U1608 (N_1608,N_1511,N_1513);
and U1609 (N_1609,N_1514,N_1541);
nor U1610 (N_1610,N_1537,N_1557);
nor U1611 (N_1611,N_1547,N_1511);
or U1612 (N_1612,N_1532,N_1537);
nand U1613 (N_1613,N_1548,N_1552);
xor U1614 (N_1614,N_1511,N_1545);
nand U1615 (N_1615,N_1524,N_1544);
nand U1616 (N_1616,N_1551,N_1532);
xor U1617 (N_1617,N_1522,N_1542);
xor U1618 (N_1618,N_1511,N_1504);
or U1619 (N_1619,N_1539,N_1541);
or U1620 (N_1620,N_1607,N_1615);
and U1621 (N_1621,N_1606,N_1610);
and U1622 (N_1622,N_1611,N_1593);
nor U1623 (N_1623,N_1575,N_1585);
and U1624 (N_1624,N_1563,N_1590);
nor U1625 (N_1625,N_1612,N_1601);
nor U1626 (N_1626,N_1573,N_1574);
nand U1627 (N_1627,N_1614,N_1613);
nor U1628 (N_1628,N_1581,N_1595);
nor U1629 (N_1629,N_1605,N_1565);
nand U1630 (N_1630,N_1602,N_1618);
nor U1631 (N_1631,N_1584,N_1603);
nand U1632 (N_1632,N_1560,N_1566);
or U1633 (N_1633,N_1592,N_1570);
and U1634 (N_1634,N_1616,N_1567);
or U1635 (N_1635,N_1586,N_1619);
or U1636 (N_1636,N_1600,N_1578);
nor U1637 (N_1637,N_1571,N_1576);
nor U1638 (N_1638,N_1604,N_1564);
and U1639 (N_1639,N_1599,N_1582);
or U1640 (N_1640,N_1579,N_1596);
xnor U1641 (N_1641,N_1609,N_1561);
nor U1642 (N_1642,N_1617,N_1572);
nor U1643 (N_1643,N_1580,N_1569);
nor U1644 (N_1644,N_1562,N_1588);
nor U1645 (N_1645,N_1568,N_1597);
nand U1646 (N_1646,N_1608,N_1577);
nor U1647 (N_1647,N_1583,N_1598);
and U1648 (N_1648,N_1594,N_1591);
or U1649 (N_1649,N_1587,N_1589);
nor U1650 (N_1650,N_1566,N_1594);
nand U1651 (N_1651,N_1605,N_1619);
nand U1652 (N_1652,N_1564,N_1589);
and U1653 (N_1653,N_1593,N_1578);
xor U1654 (N_1654,N_1560,N_1562);
and U1655 (N_1655,N_1600,N_1581);
xnor U1656 (N_1656,N_1572,N_1584);
nand U1657 (N_1657,N_1593,N_1583);
xnor U1658 (N_1658,N_1611,N_1575);
xnor U1659 (N_1659,N_1581,N_1584);
nand U1660 (N_1660,N_1573,N_1605);
and U1661 (N_1661,N_1561,N_1582);
and U1662 (N_1662,N_1604,N_1572);
nor U1663 (N_1663,N_1573,N_1606);
or U1664 (N_1664,N_1596,N_1590);
xnor U1665 (N_1665,N_1586,N_1577);
or U1666 (N_1666,N_1571,N_1619);
or U1667 (N_1667,N_1564,N_1586);
and U1668 (N_1668,N_1577,N_1598);
nand U1669 (N_1669,N_1590,N_1560);
nor U1670 (N_1670,N_1561,N_1592);
and U1671 (N_1671,N_1595,N_1596);
or U1672 (N_1672,N_1577,N_1588);
and U1673 (N_1673,N_1588,N_1591);
and U1674 (N_1674,N_1563,N_1578);
and U1675 (N_1675,N_1580,N_1578);
and U1676 (N_1676,N_1590,N_1594);
nor U1677 (N_1677,N_1614,N_1588);
xnor U1678 (N_1678,N_1581,N_1561);
nand U1679 (N_1679,N_1604,N_1593);
or U1680 (N_1680,N_1631,N_1676);
and U1681 (N_1681,N_1630,N_1636);
nand U1682 (N_1682,N_1662,N_1668);
or U1683 (N_1683,N_1656,N_1667);
or U1684 (N_1684,N_1627,N_1665);
and U1685 (N_1685,N_1672,N_1673);
nand U1686 (N_1686,N_1640,N_1641);
or U1687 (N_1687,N_1653,N_1622);
xor U1688 (N_1688,N_1671,N_1628);
and U1689 (N_1689,N_1648,N_1674);
nor U1690 (N_1690,N_1657,N_1660);
nand U1691 (N_1691,N_1646,N_1658);
nor U1692 (N_1692,N_1675,N_1652);
xnor U1693 (N_1693,N_1677,N_1655);
or U1694 (N_1694,N_1649,N_1650);
nand U1695 (N_1695,N_1647,N_1638);
or U1696 (N_1696,N_1626,N_1639);
and U1697 (N_1697,N_1623,N_1635);
xnor U1698 (N_1698,N_1632,N_1642);
or U1699 (N_1699,N_1634,N_1654);
xor U1700 (N_1700,N_1633,N_1666);
and U1701 (N_1701,N_1678,N_1670);
nor U1702 (N_1702,N_1629,N_1679);
and U1703 (N_1703,N_1621,N_1644);
nand U1704 (N_1704,N_1625,N_1661);
nor U1705 (N_1705,N_1651,N_1624);
nor U1706 (N_1706,N_1620,N_1664);
xor U1707 (N_1707,N_1663,N_1669);
nand U1708 (N_1708,N_1643,N_1645);
nand U1709 (N_1709,N_1659,N_1637);
and U1710 (N_1710,N_1650,N_1657);
xor U1711 (N_1711,N_1623,N_1667);
and U1712 (N_1712,N_1629,N_1649);
nor U1713 (N_1713,N_1666,N_1642);
nor U1714 (N_1714,N_1637,N_1673);
nor U1715 (N_1715,N_1653,N_1667);
and U1716 (N_1716,N_1637,N_1658);
xor U1717 (N_1717,N_1660,N_1648);
and U1718 (N_1718,N_1678,N_1663);
or U1719 (N_1719,N_1664,N_1624);
xnor U1720 (N_1720,N_1675,N_1653);
or U1721 (N_1721,N_1654,N_1671);
nor U1722 (N_1722,N_1661,N_1633);
or U1723 (N_1723,N_1646,N_1636);
and U1724 (N_1724,N_1672,N_1627);
nor U1725 (N_1725,N_1675,N_1649);
and U1726 (N_1726,N_1629,N_1663);
nor U1727 (N_1727,N_1621,N_1651);
nand U1728 (N_1728,N_1654,N_1659);
nor U1729 (N_1729,N_1633,N_1658);
and U1730 (N_1730,N_1673,N_1666);
nand U1731 (N_1731,N_1667,N_1664);
or U1732 (N_1732,N_1634,N_1625);
or U1733 (N_1733,N_1664,N_1648);
or U1734 (N_1734,N_1645,N_1665);
nor U1735 (N_1735,N_1635,N_1678);
or U1736 (N_1736,N_1677,N_1654);
and U1737 (N_1737,N_1663,N_1656);
nor U1738 (N_1738,N_1639,N_1637);
nand U1739 (N_1739,N_1665,N_1667);
nor U1740 (N_1740,N_1701,N_1685);
nor U1741 (N_1741,N_1686,N_1708);
nor U1742 (N_1742,N_1725,N_1704);
nand U1743 (N_1743,N_1724,N_1709);
nor U1744 (N_1744,N_1733,N_1721);
or U1745 (N_1745,N_1731,N_1702);
xor U1746 (N_1746,N_1683,N_1728);
or U1747 (N_1747,N_1682,N_1680);
nor U1748 (N_1748,N_1694,N_1688);
nand U1749 (N_1749,N_1719,N_1696);
nor U1750 (N_1750,N_1693,N_1729);
or U1751 (N_1751,N_1735,N_1695);
xnor U1752 (N_1752,N_1737,N_1711);
or U1753 (N_1753,N_1736,N_1730);
or U1754 (N_1754,N_1717,N_1690);
and U1755 (N_1755,N_1715,N_1691);
and U1756 (N_1756,N_1684,N_1698);
nor U1757 (N_1757,N_1716,N_1681);
or U1758 (N_1758,N_1718,N_1739);
nor U1759 (N_1759,N_1710,N_1726);
nor U1760 (N_1760,N_1699,N_1732);
and U1761 (N_1761,N_1692,N_1697);
or U1762 (N_1762,N_1706,N_1705);
and U1763 (N_1763,N_1703,N_1720);
and U1764 (N_1764,N_1707,N_1734);
and U1765 (N_1765,N_1700,N_1712);
nand U1766 (N_1766,N_1727,N_1687);
and U1767 (N_1767,N_1713,N_1714);
nor U1768 (N_1768,N_1689,N_1723);
and U1769 (N_1769,N_1738,N_1722);
nor U1770 (N_1770,N_1712,N_1705);
and U1771 (N_1771,N_1700,N_1701);
xor U1772 (N_1772,N_1688,N_1708);
and U1773 (N_1773,N_1734,N_1681);
nand U1774 (N_1774,N_1711,N_1734);
or U1775 (N_1775,N_1690,N_1710);
and U1776 (N_1776,N_1701,N_1721);
and U1777 (N_1777,N_1733,N_1698);
nor U1778 (N_1778,N_1719,N_1693);
or U1779 (N_1779,N_1691,N_1713);
and U1780 (N_1780,N_1689,N_1699);
nand U1781 (N_1781,N_1705,N_1736);
or U1782 (N_1782,N_1681,N_1725);
nand U1783 (N_1783,N_1694,N_1715);
or U1784 (N_1784,N_1729,N_1709);
nor U1785 (N_1785,N_1699,N_1691);
nor U1786 (N_1786,N_1724,N_1738);
nand U1787 (N_1787,N_1714,N_1702);
or U1788 (N_1788,N_1683,N_1739);
or U1789 (N_1789,N_1739,N_1725);
nor U1790 (N_1790,N_1686,N_1725);
nor U1791 (N_1791,N_1737,N_1734);
and U1792 (N_1792,N_1689,N_1708);
nor U1793 (N_1793,N_1707,N_1688);
or U1794 (N_1794,N_1739,N_1692);
nor U1795 (N_1795,N_1687,N_1691);
xor U1796 (N_1796,N_1729,N_1683);
and U1797 (N_1797,N_1714,N_1726);
or U1798 (N_1798,N_1707,N_1708);
or U1799 (N_1799,N_1697,N_1712);
or U1800 (N_1800,N_1776,N_1755);
nor U1801 (N_1801,N_1768,N_1762);
nand U1802 (N_1802,N_1797,N_1760);
or U1803 (N_1803,N_1761,N_1749);
or U1804 (N_1804,N_1778,N_1744);
nand U1805 (N_1805,N_1771,N_1782);
nand U1806 (N_1806,N_1759,N_1772);
nor U1807 (N_1807,N_1795,N_1788);
or U1808 (N_1808,N_1769,N_1796);
and U1809 (N_1809,N_1765,N_1742);
nor U1810 (N_1810,N_1774,N_1750);
or U1811 (N_1811,N_1741,N_1756);
and U1812 (N_1812,N_1783,N_1770);
or U1813 (N_1813,N_1763,N_1745);
nor U1814 (N_1814,N_1787,N_1754);
xor U1815 (N_1815,N_1784,N_1799);
nor U1816 (N_1816,N_1793,N_1775);
or U1817 (N_1817,N_1789,N_1794);
nor U1818 (N_1818,N_1777,N_1758);
nor U1819 (N_1819,N_1773,N_1786);
or U1820 (N_1820,N_1766,N_1753);
nand U1821 (N_1821,N_1752,N_1746);
xnor U1822 (N_1822,N_1747,N_1798);
and U1823 (N_1823,N_1743,N_1767);
nand U1824 (N_1824,N_1757,N_1781);
and U1825 (N_1825,N_1748,N_1792);
and U1826 (N_1826,N_1785,N_1791);
or U1827 (N_1827,N_1780,N_1740);
nor U1828 (N_1828,N_1751,N_1764);
nor U1829 (N_1829,N_1790,N_1779);
nor U1830 (N_1830,N_1772,N_1793);
nor U1831 (N_1831,N_1754,N_1788);
nand U1832 (N_1832,N_1784,N_1753);
or U1833 (N_1833,N_1755,N_1789);
or U1834 (N_1834,N_1783,N_1798);
and U1835 (N_1835,N_1752,N_1761);
xor U1836 (N_1836,N_1776,N_1783);
nor U1837 (N_1837,N_1764,N_1742);
and U1838 (N_1838,N_1777,N_1764);
nand U1839 (N_1839,N_1778,N_1787);
xor U1840 (N_1840,N_1751,N_1757);
nor U1841 (N_1841,N_1746,N_1788);
nor U1842 (N_1842,N_1793,N_1786);
nor U1843 (N_1843,N_1744,N_1793);
or U1844 (N_1844,N_1754,N_1758);
nand U1845 (N_1845,N_1796,N_1788);
nand U1846 (N_1846,N_1756,N_1785);
nand U1847 (N_1847,N_1790,N_1791);
nand U1848 (N_1848,N_1792,N_1772);
and U1849 (N_1849,N_1740,N_1760);
nand U1850 (N_1850,N_1763,N_1788);
and U1851 (N_1851,N_1769,N_1779);
or U1852 (N_1852,N_1790,N_1781);
nor U1853 (N_1853,N_1798,N_1797);
and U1854 (N_1854,N_1774,N_1741);
nor U1855 (N_1855,N_1751,N_1745);
and U1856 (N_1856,N_1766,N_1765);
nor U1857 (N_1857,N_1788,N_1782);
nand U1858 (N_1858,N_1756,N_1751);
xor U1859 (N_1859,N_1768,N_1753);
and U1860 (N_1860,N_1834,N_1820);
nand U1861 (N_1861,N_1821,N_1808);
and U1862 (N_1862,N_1824,N_1800);
and U1863 (N_1863,N_1853,N_1827);
nand U1864 (N_1864,N_1829,N_1801);
and U1865 (N_1865,N_1825,N_1812);
nor U1866 (N_1866,N_1836,N_1856);
and U1867 (N_1867,N_1823,N_1850);
or U1868 (N_1868,N_1852,N_1818);
or U1869 (N_1869,N_1838,N_1833);
or U1870 (N_1870,N_1844,N_1807);
nand U1871 (N_1871,N_1859,N_1809);
and U1872 (N_1872,N_1813,N_1846);
and U1873 (N_1873,N_1851,N_1830);
nand U1874 (N_1874,N_1817,N_1847);
or U1875 (N_1875,N_1819,N_1815);
or U1876 (N_1876,N_1806,N_1855);
or U1877 (N_1877,N_1837,N_1857);
or U1878 (N_1878,N_1843,N_1826);
or U1879 (N_1879,N_1804,N_1810);
nand U1880 (N_1880,N_1802,N_1803);
nor U1881 (N_1881,N_1840,N_1822);
and U1882 (N_1882,N_1854,N_1845);
nand U1883 (N_1883,N_1814,N_1811);
or U1884 (N_1884,N_1831,N_1816);
and U1885 (N_1885,N_1839,N_1805);
and U1886 (N_1886,N_1835,N_1832);
and U1887 (N_1887,N_1858,N_1848);
or U1888 (N_1888,N_1842,N_1849);
or U1889 (N_1889,N_1828,N_1841);
xnor U1890 (N_1890,N_1845,N_1800);
nor U1891 (N_1891,N_1806,N_1802);
xor U1892 (N_1892,N_1840,N_1802);
nand U1893 (N_1893,N_1853,N_1826);
or U1894 (N_1894,N_1856,N_1809);
nand U1895 (N_1895,N_1835,N_1805);
or U1896 (N_1896,N_1847,N_1801);
nand U1897 (N_1897,N_1827,N_1816);
nor U1898 (N_1898,N_1838,N_1813);
nor U1899 (N_1899,N_1812,N_1844);
and U1900 (N_1900,N_1839,N_1813);
or U1901 (N_1901,N_1839,N_1808);
nand U1902 (N_1902,N_1803,N_1841);
or U1903 (N_1903,N_1831,N_1807);
or U1904 (N_1904,N_1829,N_1814);
nor U1905 (N_1905,N_1842,N_1846);
xnor U1906 (N_1906,N_1843,N_1836);
nor U1907 (N_1907,N_1825,N_1835);
nor U1908 (N_1908,N_1848,N_1847);
nand U1909 (N_1909,N_1854,N_1846);
nand U1910 (N_1910,N_1805,N_1820);
or U1911 (N_1911,N_1824,N_1806);
or U1912 (N_1912,N_1840,N_1818);
nand U1913 (N_1913,N_1838,N_1806);
xnor U1914 (N_1914,N_1839,N_1831);
xnor U1915 (N_1915,N_1848,N_1810);
nor U1916 (N_1916,N_1850,N_1844);
or U1917 (N_1917,N_1826,N_1852);
xor U1918 (N_1918,N_1823,N_1838);
and U1919 (N_1919,N_1830,N_1810);
nand U1920 (N_1920,N_1894,N_1865);
nand U1921 (N_1921,N_1916,N_1907);
xor U1922 (N_1922,N_1884,N_1877);
nor U1923 (N_1923,N_1892,N_1899);
nor U1924 (N_1924,N_1889,N_1896);
nor U1925 (N_1925,N_1862,N_1898);
nand U1926 (N_1926,N_1906,N_1885);
xnor U1927 (N_1927,N_1912,N_1913);
or U1928 (N_1928,N_1911,N_1871);
nor U1929 (N_1929,N_1869,N_1868);
nand U1930 (N_1930,N_1890,N_1886);
xnor U1931 (N_1931,N_1897,N_1883);
nor U1932 (N_1932,N_1915,N_1902);
nand U1933 (N_1933,N_1872,N_1880);
and U1934 (N_1934,N_1873,N_1914);
nand U1935 (N_1935,N_1878,N_1910);
and U1936 (N_1936,N_1864,N_1860);
nor U1937 (N_1937,N_1866,N_1861);
nor U1938 (N_1938,N_1904,N_1909);
or U1939 (N_1939,N_1876,N_1870);
nand U1940 (N_1940,N_1901,N_1895);
nor U1941 (N_1941,N_1919,N_1882);
and U1942 (N_1942,N_1893,N_1888);
or U1943 (N_1943,N_1918,N_1900);
or U1944 (N_1944,N_1881,N_1891);
nand U1945 (N_1945,N_1863,N_1903);
xnor U1946 (N_1946,N_1874,N_1905);
nand U1947 (N_1947,N_1917,N_1879);
nor U1948 (N_1948,N_1867,N_1908);
or U1949 (N_1949,N_1875,N_1887);
or U1950 (N_1950,N_1881,N_1912);
and U1951 (N_1951,N_1892,N_1869);
nor U1952 (N_1952,N_1902,N_1887);
nand U1953 (N_1953,N_1904,N_1869);
nand U1954 (N_1954,N_1888,N_1866);
nor U1955 (N_1955,N_1881,N_1875);
or U1956 (N_1956,N_1867,N_1893);
nor U1957 (N_1957,N_1902,N_1904);
nor U1958 (N_1958,N_1872,N_1891);
nor U1959 (N_1959,N_1899,N_1905);
or U1960 (N_1960,N_1887,N_1903);
nor U1961 (N_1961,N_1909,N_1914);
nand U1962 (N_1962,N_1865,N_1874);
or U1963 (N_1963,N_1866,N_1886);
xnor U1964 (N_1964,N_1913,N_1882);
xnor U1965 (N_1965,N_1915,N_1899);
nor U1966 (N_1966,N_1906,N_1890);
nor U1967 (N_1967,N_1875,N_1870);
or U1968 (N_1968,N_1910,N_1880);
or U1969 (N_1969,N_1914,N_1874);
and U1970 (N_1970,N_1911,N_1900);
xnor U1971 (N_1971,N_1864,N_1903);
and U1972 (N_1972,N_1910,N_1864);
nor U1973 (N_1973,N_1866,N_1902);
or U1974 (N_1974,N_1895,N_1892);
and U1975 (N_1975,N_1881,N_1890);
nor U1976 (N_1976,N_1860,N_1906);
nor U1977 (N_1977,N_1883,N_1867);
and U1978 (N_1978,N_1875,N_1892);
nor U1979 (N_1979,N_1868,N_1883);
nor U1980 (N_1980,N_1928,N_1973);
nor U1981 (N_1981,N_1941,N_1978);
nand U1982 (N_1982,N_1957,N_1970);
or U1983 (N_1983,N_1968,N_1944);
nor U1984 (N_1984,N_1931,N_1950);
nor U1985 (N_1985,N_1937,N_1976);
xnor U1986 (N_1986,N_1954,N_1934);
and U1987 (N_1987,N_1924,N_1930);
nor U1988 (N_1988,N_1947,N_1964);
nand U1989 (N_1989,N_1958,N_1966);
or U1990 (N_1990,N_1972,N_1923);
and U1991 (N_1991,N_1969,N_1960);
nor U1992 (N_1992,N_1967,N_1940);
nor U1993 (N_1993,N_1920,N_1961);
nor U1994 (N_1994,N_1956,N_1922);
or U1995 (N_1995,N_1953,N_1927);
xnor U1996 (N_1996,N_1932,N_1925);
and U1997 (N_1997,N_1951,N_1942);
nand U1998 (N_1998,N_1936,N_1938);
or U1999 (N_1999,N_1977,N_1975);
or U2000 (N_2000,N_1974,N_1955);
xor U2001 (N_2001,N_1971,N_1933);
or U2002 (N_2002,N_1945,N_1921);
nand U2003 (N_2003,N_1935,N_1939);
and U2004 (N_2004,N_1929,N_1979);
or U2005 (N_2005,N_1962,N_1959);
nor U2006 (N_2006,N_1946,N_1963);
xor U2007 (N_2007,N_1949,N_1943);
nand U2008 (N_2008,N_1965,N_1952);
or U2009 (N_2009,N_1948,N_1926);
nand U2010 (N_2010,N_1958,N_1932);
xnor U2011 (N_2011,N_1968,N_1956);
and U2012 (N_2012,N_1959,N_1955);
or U2013 (N_2013,N_1961,N_1948);
or U2014 (N_2014,N_1968,N_1933);
or U2015 (N_2015,N_1971,N_1951);
and U2016 (N_2016,N_1969,N_1966);
and U2017 (N_2017,N_1975,N_1973);
nand U2018 (N_2018,N_1974,N_1954);
and U2019 (N_2019,N_1927,N_1961);
nor U2020 (N_2020,N_1948,N_1950);
or U2021 (N_2021,N_1925,N_1923);
nand U2022 (N_2022,N_1941,N_1975);
and U2023 (N_2023,N_1920,N_1930);
or U2024 (N_2024,N_1963,N_1923);
nor U2025 (N_2025,N_1931,N_1964);
and U2026 (N_2026,N_1961,N_1932);
or U2027 (N_2027,N_1956,N_1937);
or U2028 (N_2028,N_1967,N_1942);
nand U2029 (N_2029,N_1950,N_1940);
and U2030 (N_2030,N_1947,N_1958);
and U2031 (N_2031,N_1926,N_1952);
and U2032 (N_2032,N_1947,N_1951);
and U2033 (N_2033,N_1924,N_1922);
or U2034 (N_2034,N_1940,N_1962);
or U2035 (N_2035,N_1964,N_1923);
xor U2036 (N_2036,N_1961,N_1963);
and U2037 (N_2037,N_1942,N_1962);
and U2038 (N_2038,N_1951,N_1963);
or U2039 (N_2039,N_1943,N_1963);
xnor U2040 (N_2040,N_2025,N_1980);
xnor U2041 (N_2041,N_1986,N_2035);
nand U2042 (N_2042,N_2006,N_2003);
and U2043 (N_2043,N_2032,N_1981);
nor U2044 (N_2044,N_2010,N_2011);
nand U2045 (N_2045,N_1990,N_2027);
nor U2046 (N_2046,N_1999,N_2024);
nor U2047 (N_2047,N_2021,N_2014);
or U2048 (N_2048,N_2001,N_2031);
nor U2049 (N_2049,N_2018,N_2037);
and U2050 (N_2050,N_2038,N_1987);
xnor U2051 (N_2051,N_1994,N_2019);
nand U2052 (N_2052,N_2036,N_1988);
and U2053 (N_2053,N_2017,N_2000);
and U2054 (N_2054,N_2007,N_2028);
or U2055 (N_2055,N_2022,N_2002);
xnor U2056 (N_2056,N_1983,N_2013);
and U2057 (N_2057,N_2039,N_1997);
nor U2058 (N_2058,N_1996,N_1995);
and U2059 (N_2059,N_2033,N_2023);
xor U2060 (N_2060,N_2009,N_1998);
nor U2061 (N_2061,N_2020,N_1992);
nand U2062 (N_2062,N_2012,N_2026);
or U2063 (N_2063,N_1991,N_2015);
nor U2064 (N_2064,N_2016,N_2030);
nand U2065 (N_2065,N_1985,N_1993);
and U2066 (N_2066,N_2029,N_2005);
nor U2067 (N_2067,N_1982,N_2008);
and U2068 (N_2068,N_1984,N_2034);
and U2069 (N_2069,N_1989,N_2004);
or U2070 (N_2070,N_2016,N_1981);
and U2071 (N_2071,N_2034,N_2031);
and U2072 (N_2072,N_1991,N_1996);
xnor U2073 (N_2073,N_2000,N_2013);
xor U2074 (N_2074,N_1980,N_2007);
nor U2075 (N_2075,N_1994,N_2014);
nor U2076 (N_2076,N_2003,N_1991);
or U2077 (N_2077,N_2006,N_2010);
and U2078 (N_2078,N_2015,N_2009);
nor U2079 (N_2079,N_1999,N_2011);
nor U2080 (N_2080,N_2030,N_1998);
and U2081 (N_2081,N_2028,N_2029);
or U2082 (N_2082,N_1991,N_2036);
and U2083 (N_2083,N_2009,N_2019);
or U2084 (N_2084,N_2008,N_1981);
or U2085 (N_2085,N_2022,N_1980);
nor U2086 (N_2086,N_2007,N_1988);
nor U2087 (N_2087,N_2009,N_1981);
nor U2088 (N_2088,N_1994,N_1986);
nor U2089 (N_2089,N_2015,N_2013);
nand U2090 (N_2090,N_2004,N_2015);
nor U2091 (N_2091,N_1983,N_2023);
nor U2092 (N_2092,N_2012,N_1999);
nand U2093 (N_2093,N_1998,N_2024);
xnor U2094 (N_2094,N_2008,N_2000);
or U2095 (N_2095,N_2003,N_2023);
and U2096 (N_2096,N_2032,N_1992);
nor U2097 (N_2097,N_2001,N_2024);
xor U2098 (N_2098,N_2035,N_2032);
and U2099 (N_2099,N_2026,N_2003);
or U2100 (N_2100,N_2099,N_2073);
or U2101 (N_2101,N_2047,N_2070);
nor U2102 (N_2102,N_2097,N_2044);
nor U2103 (N_2103,N_2096,N_2078);
and U2104 (N_2104,N_2085,N_2095);
or U2105 (N_2105,N_2046,N_2065);
or U2106 (N_2106,N_2068,N_2089);
and U2107 (N_2107,N_2080,N_2043);
nand U2108 (N_2108,N_2040,N_2059);
xnor U2109 (N_2109,N_2087,N_2041);
xnor U2110 (N_2110,N_2090,N_2053);
and U2111 (N_2111,N_2091,N_2064);
nor U2112 (N_2112,N_2093,N_2058);
nor U2113 (N_2113,N_2076,N_2081);
and U2114 (N_2114,N_2051,N_2056);
or U2115 (N_2115,N_2062,N_2063);
and U2116 (N_2116,N_2071,N_2088);
nand U2117 (N_2117,N_2086,N_2079);
or U2118 (N_2118,N_2067,N_2077);
and U2119 (N_2119,N_2084,N_2042);
or U2120 (N_2120,N_2069,N_2094);
or U2121 (N_2121,N_2061,N_2082);
and U2122 (N_2122,N_2050,N_2098);
xnor U2123 (N_2123,N_2092,N_2074);
nor U2124 (N_2124,N_2048,N_2049);
nor U2125 (N_2125,N_2054,N_2052);
and U2126 (N_2126,N_2057,N_2060);
or U2127 (N_2127,N_2083,N_2045);
nand U2128 (N_2128,N_2075,N_2072);
nand U2129 (N_2129,N_2055,N_2066);
nand U2130 (N_2130,N_2067,N_2085);
or U2131 (N_2131,N_2092,N_2083);
and U2132 (N_2132,N_2097,N_2089);
xor U2133 (N_2133,N_2070,N_2065);
nor U2134 (N_2134,N_2052,N_2085);
or U2135 (N_2135,N_2097,N_2082);
xor U2136 (N_2136,N_2078,N_2049);
and U2137 (N_2137,N_2055,N_2080);
xor U2138 (N_2138,N_2080,N_2079);
or U2139 (N_2139,N_2086,N_2090);
nor U2140 (N_2140,N_2045,N_2069);
nand U2141 (N_2141,N_2049,N_2054);
and U2142 (N_2142,N_2067,N_2060);
nand U2143 (N_2143,N_2042,N_2078);
and U2144 (N_2144,N_2086,N_2095);
nand U2145 (N_2145,N_2043,N_2062);
nand U2146 (N_2146,N_2052,N_2073);
nor U2147 (N_2147,N_2069,N_2059);
or U2148 (N_2148,N_2063,N_2098);
or U2149 (N_2149,N_2062,N_2041);
nor U2150 (N_2150,N_2058,N_2077);
and U2151 (N_2151,N_2054,N_2088);
or U2152 (N_2152,N_2078,N_2071);
nand U2153 (N_2153,N_2055,N_2046);
nand U2154 (N_2154,N_2057,N_2052);
xor U2155 (N_2155,N_2077,N_2071);
nor U2156 (N_2156,N_2082,N_2079);
and U2157 (N_2157,N_2063,N_2043);
nand U2158 (N_2158,N_2060,N_2097);
nor U2159 (N_2159,N_2099,N_2052);
and U2160 (N_2160,N_2137,N_2135);
or U2161 (N_2161,N_2117,N_2106);
nand U2162 (N_2162,N_2126,N_2144);
nor U2163 (N_2163,N_2139,N_2111);
or U2164 (N_2164,N_2102,N_2128);
nand U2165 (N_2165,N_2110,N_2153);
nor U2166 (N_2166,N_2114,N_2100);
and U2167 (N_2167,N_2143,N_2157);
nor U2168 (N_2168,N_2146,N_2159);
or U2169 (N_2169,N_2154,N_2119);
nor U2170 (N_2170,N_2136,N_2141);
or U2171 (N_2171,N_2145,N_2127);
nor U2172 (N_2172,N_2140,N_2104);
nor U2173 (N_2173,N_2142,N_2134);
nor U2174 (N_2174,N_2107,N_2118);
nor U2175 (N_2175,N_2123,N_2150);
and U2176 (N_2176,N_2129,N_2131);
or U2177 (N_2177,N_2103,N_2148);
or U2178 (N_2178,N_2101,N_2152);
nand U2179 (N_2179,N_2125,N_2109);
and U2180 (N_2180,N_2105,N_2158);
xnor U2181 (N_2181,N_2156,N_2113);
nor U2182 (N_2182,N_2120,N_2151);
nor U2183 (N_2183,N_2116,N_2149);
or U2184 (N_2184,N_2121,N_2108);
nand U2185 (N_2185,N_2133,N_2155);
xor U2186 (N_2186,N_2112,N_2124);
and U2187 (N_2187,N_2122,N_2147);
and U2188 (N_2188,N_2130,N_2132);
and U2189 (N_2189,N_2138,N_2115);
nand U2190 (N_2190,N_2136,N_2132);
nand U2191 (N_2191,N_2113,N_2116);
xor U2192 (N_2192,N_2100,N_2151);
nor U2193 (N_2193,N_2110,N_2158);
nand U2194 (N_2194,N_2157,N_2121);
and U2195 (N_2195,N_2117,N_2102);
nor U2196 (N_2196,N_2132,N_2131);
xor U2197 (N_2197,N_2113,N_2134);
nor U2198 (N_2198,N_2110,N_2103);
or U2199 (N_2199,N_2151,N_2110);
and U2200 (N_2200,N_2118,N_2128);
nand U2201 (N_2201,N_2131,N_2147);
and U2202 (N_2202,N_2143,N_2148);
or U2203 (N_2203,N_2152,N_2128);
nor U2204 (N_2204,N_2108,N_2135);
xor U2205 (N_2205,N_2132,N_2121);
and U2206 (N_2206,N_2152,N_2111);
nor U2207 (N_2207,N_2146,N_2157);
nand U2208 (N_2208,N_2149,N_2155);
nand U2209 (N_2209,N_2123,N_2113);
or U2210 (N_2210,N_2140,N_2121);
and U2211 (N_2211,N_2153,N_2115);
or U2212 (N_2212,N_2114,N_2130);
nor U2213 (N_2213,N_2100,N_2130);
or U2214 (N_2214,N_2154,N_2106);
nand U2215 (N_2215,N_2133,N_2126);
nor U2216 (N_2216,N_2158,N_2136);
xor U2217 (N_2217,N_2152,N_2154);
nand U2218 (N_2218,N_2122,N_2124);
or U2219 (N_2219,N_2138,N_2125);
xor U2220 (N_2220,N_2169,N_2180);
or U2221 (N_2221,N_2212,N_2175);
nand U2222 (N_2222,N_2185,N_2168);
nand U2223 (N_2223,N_2201,N_2186);
or U2224 (N_2224,N_2163,N_2203);
nand U2225 (N_2225,N_2204,N_2191);
nor U2226 (N_2226,N_2215,N_2167);
nor U2227 (N_2227,N_2173,N_2207);
nand U2228 (N_2228,N_2182,N_2205);
nand U2229 (N_2229,N_2174,N_2200);
or U2230 (N_2230,N_2184,N_2161);
nor U2231 (N_2231,N_2162,N_2188);
nor U2232 (N_2232,N_2165,N_2193);
or U2233 (N_2233,N_2192,N_2211);
or U2234 (N_2234,N_2195,N_2183);
nand U2235 (N_2235,N_2206,N_2196);
nand U2236 (N_2236,N_2214,N_2160);
and U2237 (N_2237,N_2219,N_2164);
nand U2238 (N_2238,N_2202,N_2189);
nand U2239 (N_2239,N_2208,N_2178);
and U2240 (N_2240,N_2198,N_2172);
or U2241 (N_2241,N_2170,N_2217);
or U2242 (N_2242,N_2194,N_2176);
or U2243 (N_2243,N_2209,N_2210);
nor U2244 (N_2244,N_2187,N_2181);
and U2245 (N_2245,N_2177,N_2216);
or U2246 (N_2246,N_2190,N_2199);
nor U2247 (N_2247,N_2197,N_2166);
and U2248 (N_2248,N_2218,N_2171);
nand U2249 (N_2249,N_2179,N_2213);
xor U2250 (N_2250,N_2211,N_2207);
xnor U2251 (N_2251,N_2176,N_2182);
or U2252 (N_2252,N_2212,N_2203);
and U2253 (N_2253,N_2199,N_2179);
or U2254 (N_2254,N_2182,N_2178);
nand U2255 (N_2255,N_2198,N_2207);
nand U2256 (N_2256,N_2170,N_2177);
nand U2257 (N_2257,N_2185,N_2169);
or U2258 (N_2258,N_2182,N_2166);
and U2259 (N_2259,N_2194,N_2162);
xor U2260 (N_2260,N_2165,N_2194);
xnor U2261 (N_2261,N_2214,N_2201);
or U2262 (N_2262,N_2160,N_2189);
nand U2263 (N_2263,N_2187,N_2208);
nor U2264 (N_2264,N_2179,N_2171);
nand U2265 (N_2265,N_2185,N_2217);
nor U2266 (N_2266,N_2193,N_2206);
nand U2267 (N_2267,N_2176,N_2193);
and U2268 (N_2268,N_2197,N_2211);
or U2269 (N_2269,N_2171,N_2212);
and U2270 (N_2270,N_2175,N_2167);
and U2271 (N_2271,N_2172,N_2160);
xor U2272 (N_2272,N_2179,N_2184);
and U2273 (N_2273,N_2162,N_2197);
nor U2274 (N_2274,N_2204,N_2212);
and U2275 (N_2275,N_2168,N_2194);
xnor U2276 (N_2276,N_2184,N_2187);
or U2277 (N_2277,N_2184,N_2205);
or U2278 (N_2278,N_2186,N_2168);
xnor U2279 (N_2279,N_2170,N_2196);
and U2280 (N_2280,N_2271,N_2254);
or U2281 (N_2281,N_2245,N_2259);
and U2282 (N_2282,N_2233,N_2274);
nand U2283 (N_2283,N_2230,N_2267);
nor U2284 (N_2284,N_2229,N_2257);
nand U2285 (N_2285,N_2240,N_2239);
nor U2286 (N_2286,N_2237,N_2224);
nor U2287 (N_2287,N_2252,N_2236);
xor U2288 (N_2288,N_2263,N_2273);
or U2289 (N_2289,N_2265,N_2256);
xor U2290 (N_2290,N_2248,N_2228);
or U2291 (N_2291,N_2242,N_2234);
and U2292 (N_2292,N_2255,N_2220);
and U2293 (N_2293,N_2226,N_2264);
or U2294 (N_2294,N_2244,N_2268);
nand U2295 (N_2295,N_2247,N_2253);
and U2296 (N_2296,N_2227,N_2269);
nor U2297 (N_2297,N_2262,N_2225);
xor U2298 (N_2298,N_2258,N_2221);
and U2299 (N_2299,N_2223,N_2238);
nor U2300 (N_2300,N_2270,N_2260);
nor U2301 (N_2301,N_2250,N_2278);
nor U2302 (N_2302,N_2266,N_2251);
nor U2303 (N_2303,N_2275,N_2246);
or U2304 (N_2304,N_2272,N_2277);
and U2305 (N_2305,N_2231,N_2279);
nand U2306 (N_2306,N_2232,N_2249);
and U2307 (N_2307,N_2222,N_2261);
and U2308 (N_2308,N_2243,N_2276);
or U2309 (N_2309,N_2241,N_2235);
nand U2310 (N_2310,N_2269,N_2279);
and U2311 (N_2311,N_2258,N_2241);
nand U2312 (N_2312,N_2272,N_2244);
or U2313 (N_2313,N_2250,N_2266);
nor U2314 (N_2314,N_2279,N_2235);
nor U2315 (N_2315,N_2223,N_2268);
nor U2316 (N_2316,N_2274,N_2272);
and U2317 (N_2317,N_2226,N_2274);
or U2318 (N_2318,N_2241,N_2240);
nor U2319 (N_2319,N_2236,N_2239);
and U2320 (N_2320,N_2248,N_2235);
nor U2321 (N_2321,N_2273,N_2252);
xor U2322 (N_2322,N_2234,N_2245);
or U2323 (N_2323,N_2260,N_2268);
or U2324 (N_2324,N_2253,N_2230);
nand U2325 (N_2325,N_2227,N_2229);
nor U2326 (N_2326,N_2225,N_2228);
or U2327 (N_2327,N_2243,N_2230);
or U2328 (N_2328,N_2224,N_2275);
and U2329 (N_2329,N_2243,N_2258);
nand U2330 (N_2330,N_2253,N_2277);
nand U2331 (N_2331,N_2256,N_2260);
nand U2332 (N_2332,N_2241,N_2269);
nor U2333 (N_2333,N_2269,N_2222);
and U2334 (N_2334,N_2221,N_2238);
or U2335 (N_2335,N_2223,N_2255);
nor U2336 (N_2336,N_2258,N_2220);
nand U2337 (N_2337,N_2237,N_2231);
nor U2338 (N_2338,N_2259,N_2241);
or U2339 (N_2339,N_2258,N_2246);
or U2340 (N_2340,N_2297,N_2287);
nand U2341 (N_2341,N_2337,N_2334);
and U2342 (N_2342,N_2335,N_2321);
or U2343 (N_2343,N_2336,N_2283);
and U2344 (N_2344,N_2339,N_2301);
nand U2345 (N_2345,N_2330,N_2303);
and U2346 (N_2346,N_2305,N_2322);
and U2347 (N_2347,N_2294,N_2309);
nor U2348 (N_2348,N_2299,N_2291);
nand U2349 (N_2349,N_2326,N_2325);
nand U2350 (N_2350,N_2338,N_2319);
and U2351 (N_2351,N_2328,N_2308);
nor U2352 (N_2352,N_2296,N_2315);
nand U2353 (N_2353,N_2289,N_2285);
nor U2354 (N_2354,N_2286,N_2288);
or U2355 (N_2355,N_2304,N_2314);
and U2356 (N_2356,N_2312,N_2293);
nand U2357 (N_2357,N_2298,N_2292);
xnor U2358 (N_2358,N_2331,N_2300);
nand U2359 (N_2359,N_2324,N_2310);
or U2360 (N_2360,N_2316,N_2329);
nor U2361 (N_2361,N_2323,N_2332);
nor U2362 (N_2362,N_2295,N_2320);
or U2363 (N_2363,N_2306,N_2307);
nor U2364 (N_2364,N_2282,N_2302);
nand U2365 (N_2365,N_2311,N_2333);
nand U2366 (N_2366,N_2317,N_2284);
nand U2367 (N_2367,N_2327,N_2281);
nor U2368 (N_2368,N_2290,N_2313);
or U2369 (N_2369,N_2318,N_2280);
or U2370 (N_2370,N_2318,N_2328);
and U2371 (N_2371,N_2289,N_2296);
nand U2372 (N_2372,N_2310,N_2322);
or U2373 (N_2373,N_2338,N_2337);
or U2374 (N_2374,N_2327,N_2336);
nor U2375 (N_2375,N_2294,N_2282);
nand U2376 (N_2376,N_2304,N_2300);
nor U2377 (N_2377,N_2296,N_2324);
nor U2378 (N_2378,N_2320,N_2313);
and U2379 (N_2379,N_2291,N_2308);
nand U2380 (N_2380,N_2311,N_2286);
or U2381 (N_2381,N_2326,N_2316);
xnor U2382 (N_2382,N_2333,N_2295);
nor U2383 (N_2383,N_2325,N_2313);
nand U2384 (N_2384,N_2336,N_2330);
xnor U2385 (N_2385,N_2289,N_2306);
nor U2386 (N_2386,N_2335,N_2330);
or U2387 (N_2387,N_2334,N_2320);
nor U2388 (N_2388,N_2339,N_2319);
nand U2389 (N_2389,N_2311,N_2336);
or U2390 (N_2390,N_2326,N_2329);
nor U2391 (N_2391,N_2318,N_2339);
nand U2392 (N_2392,N_2293,N_2335);
nand U2393 (N_2393,N_2301,N_2331);
nor U2394 (N_2394,N_2313,N_2307);
nand U2395 (N_2395,N_2304,N_2317);
nor U2396 (N_2396,N_2302,N_2306);
or U2397 (N_2397,N_2295,N_2293);
nor U2398 (N_2398,N_2294,N_2316);
nor U2399 (N_2399,N_2327,N_2293);
and U2400 (N_2400,N_2381,N_2358);
and U2401 (N_2401,N_2360,N_2379);
and U2402 (N_2402,N_2384,N_2366);
or U2403 (N_2403,N_2359,N_2369);
and U2404 (N_2404,N_2350,N_2365);
nand U2405 (N_2405,N_2390,N_2356);
nand U2406 (N_2406,N_2348,N_2351);
xnor U2407 (N_2407,N_2373,N_2364);
xnor U2408 (N_2408,N_2355,N_2353);
xor U2409 (N_2409,N_2382,N_2344);
nand U2410 (N_2410,N_2354,N_2394);
xor U2411 (N_2411,N_2340,N_2357);
or U2412 (N_2412,N_2397,N_2375);
and U2413 (N_2413,N_2378,N_2383);
nand U2414 (N_2414,N_2387,N_2398);
or U2415 (N_2415,N_2376,N_2341);
nand U2416 (N_2416,N_2347,N_2367);
xnor U2417 (N_2417,N_2346,N_2345);
and U2418 (N_2418,N_2380,N_2363);
or U2419 (N_2419,N_2370,N_2374);
or U2420 (N_2420,N_2352,N_2377);
or U2421 (N_2421,N_2385,N_2393);
nand U2422 (N_2422,N_2368,N_2349);
and U2423 (N_2423,N_2388,N_2399);
or U2424 (N_2424,N_2395,N_2392);
nor U2425 (N_2425,N_2386,N_2342);
or U2426 (N_2426,N_2391,N_2362);
nand U2427 (N_2427,N_2389,N_2371);
nor U2428 (N_2428,N_2396,N_2372);
nor U2429 (N_2429,N_2361,N_2343);
or U2430 (N_2430,N_2390,N_2365);
and U2431 (N_2431,N_2381,N_2341);
and U2432 (N_2432,N_2349,N_2355);
nor U2433 (N_2433,N_2342,N_2388);
nand U2434 (N_2434,N_2372,N_2374);
or U2435 (N_2435,N_2340,N_2394);
nand U2436 (N_2436,N_2387,N_2346);
nor U2437 (N_2437,N_2381,N_2364);
and U2438 (N_2438,N_2342,N_2344);
nor U2439 (N_2439,N_2345,N_2353);
or U2440 (N_2440,N_2340,N_2374);
or U2441 (N_2441,N_2350,N_2354);
nand U2442 (N_2442,N_2398,N_2362);
nor U2443 (N_2443,N_2392,N_2379);
xnor U2444 (N_2444,N_2389,N_2391);
nor U2445 (N_2445,N_2381,N_2380);
nor U2446 (N_2446,N_2340,N_2349);
nor U2447 (N_2447,N_2353,N_2360);
or U2448 (N_2448,N_2379,N_2395);
nor U2449 (N_2449,N_2372,N_2356);
and U2450 (N_2450,N_2384,N_2373);
xor U2451 (N_2451,N_2386,N_2362);
nor U2452 (N_2452,N_2342,N_2382);
nand U2453 (N_2453,N_2347,N_2358);
nor U2454 (N_2454,N_2382,N_2383);
or U2455 (N_2455,N_2351,N_2391);
or U2456 (N_2456,N_2362,N_2392);
xnor U2457 (N_2457,N_2343,N_2363);
nand U2458 (N_2458,N_2364,N_2396);
and U2459 (N_2459,N_2376,N_2389);
nor U2460 (N_2460,N_2445,N_2412);
nor U2461 (N_2461,N_2415,N_2425);
nor U2462 (N_2462,N_2413,N_2434);
nand U2463 (N_2463,N_2420,N_2424);
nor U2464 (N_2464,N_2444,N_2442);
nand U2465 (N_2465,N_2429,N_2450);
xnor U2466 (N_2466,N_2416,N_2418);
or U2467 (N_2467,N_2454,N_2432);
nor U2468 (N_2468,N_2403,N_2437);
and U2469 (N_2469,N_2439,N_2406);
nand U2470 (N_2470,N_2401,N_2443);
xnor U2471 (N_2471,N_2448,N_2456);
nor U2472 (N_2472,N_2447,N_2457);
nor U2473 (N_2473,N_2421,N_2410);
xor U2474 (N_2474,N_2407,N_2449);
xnor U2475 (N_2475,N_2419,N_2414);
nand U2476 (N_2476,N_2411,N_2431);
nand U2477 (N_2477,N_2408,N_2428);
xnor U2478 (N_2478,N_2451,N_2427);
and U2479 (N_2479,N_2458,N_2438);
nand U2480 (N_2480,N_2452,N_2422);
nor U2481 (N_2481,N_2430,N_2459);
or U2482 (N_2482,N_2435,N_2404);
nor U2483 (N_2483,N_2441,N_2446);
nand U2484 (N_2484,N_2440,N_2400);
nand U2485 (N_2485,N_2433,N_2455);
or U2486 (N_2486,N_2423,N_2405);
nor U2487 (N_2487,N_2436,N_2402);
and U2488 (N_2488,N_2453,N_2426);
or U2489 (N_2489,N_2417,N_2409);
and U2490 (N_2490,N_2457,N_2433);
nor U2491 (N_2491,N_2435,N_2414);
nand U2492 (N_2492,N_2439,N_2447);
nor U2493 (N_2493,N_2422,N_2439);
nor U2494 (N_2494,N_2452,N_2432);
nor U2495 (N_2495,N_2449,N_2419);
xnor U2496 (N_2496,N_2441,N_2458);
nor U2497 (N_2497,N_2440,N_2449);
nor U2498 (N_2498,N_2408,N_2425);
and U2499 (N_2499,N_2433,N_2445);
or U2500 (N_2500,N_2413,N_2417);
and U2501 (N_2501,N_2433,N_2414);
nand U2502 (N_2502,N_2402,N_2400);
and U2503 (N_2503,N_2426,N_2429);
and U2504 (N_2504,N_2447,N_2453);
or U2505 (N_2505,N_2423,N_2429);
nand U2506 (N_2506,N_2444,N_2449);
nand U2507 (N_2507,N_2453,N_2408);
and U2508 (N_2508,N_2457,N_2437);
and U2509 (N_2509,N_2438,N_2401);
nand U2510 (N_2510,N_2418,N_2433);
xnor U2511 (N_2511,N_2433,N_2426);
or U2512 (N_2512,N_2441,N_2459);
and U2513 (N_2513,N_2410,N_2453);
nand U2514 (N_2514,N_2430,N_2421);
nor U2515 (N_2515,N_2442,N_2456);
xnor U2516 (N_2516,N_2452,N_2447);
nor U2517 (N_2517,N_2450,N_2407);
and U2518 (N_2518,N_2458,N_2423);
xnor U2519 (N_2519,N_2401,N_2432);
or U2520 (N_2520,N_2511,N_2514);
nor U2521 (N_2521,N_2484,N_2508);
nand U2522 (N_2522,N_2515,N_2497);
nand U2523 (N_2523,N_2466,N_2502);
or U2524 (N_2524,N_2476,N_2460);
xor U2525 (N_2525,N_2483,N_2498);
nor U2526 (N_2526,N_2462,N_2503);
or U2527 (N_2527,N_2491,N_2482);
or U2528 (N_2528,N_2494,N_2500);
and U2529 (N_2529,N_2464,N_2501);
nor U2530 (N_2530,N_2465,N_2485);
or U2531 (N_2531,N_2499,N_2467);
nand U2532 (N_2532,N_2475,N_2507);
and U2533 (N_2533,N_2469,N_2489);
xor U2534 (N_2534,N_2477,N_2470);
nand U2535 (N_2535,N_2510,N_2481);
or U2536 (N_2536,N_2488,N_2471);
or U2537 (N_2537,N_2479,N_2504);
or U2538 (N_2538,N_2461,N_2505);
nand U2539 (N_2539,N_2495,N_2517);
nand U2540 (N_2540,N_2480,N_2519);
and U2541 (N_2541,N_2486,N_2473);
or U2542 (N_2542,N_2472,N_2516);
nor U2543 (N_2543,N_2496,N_2474);
nand U2544 (N_2544,N_2512,N_2468);
nand U2545 (N_2545,N_2518,N_2492);
xnor U2546 (N_2546,N_2463,N_2490);
or U2547 (N_2547,N_2478,N_2506);
xor U2548 (N_2548,N_2487,N_2493);
or U2549 (N_2549,N_2509,N_2513);
and U2550 (N_2550,N_2475,N_2461);
or U2551 (N_2551,N_2490,N_2493);
nand U2552 (N_2552,N_2513,N_2489);
or U2553 (N_2553,N_2503,N_2508);
or U2554 (N_2554,N_2479,N_2469);
or U2555 (N_2555,N_2494,N_2462);
xnor U2556 (N_2556,N_2506,N_2495);
nor U2557 (N_2557,N_2513,N_2510);
and U2558 (N_2558,N_2460,N_2473);
xnor U2559 (N_2559,N_2497,N_2496);
nand U2560 (N_2560,N_2490,N_2502);
nor U2561 (N_2561,N_2497,N_2462);
nand U2562 (N_2562,N_2500,N_2482);
or U2563 (N_2563,N_2495,N_2493);
xor U2564 (N_2564,N_2504,N_2509);
nor U2565 (N_2565,N_2508,N_2476);
or U2566 (N_2566,N_2462,N_2498);
nand U2567 (N_2567,N_2504,N_2516);
or U2568 (N_2568,N_2510,N_2471);
nand U2569 (N_2569,N_2501,N_2473);
or U2570 (N_2570,N_2464,N_2477);
nor U2571 (N_2571,N_2491,N_2518);
nor U2572 (N_2572,N_2517,N_2477);
or U2573 (N_2573,N_2479,N_2516);
xor U2574 (N_2574,N_2470,N_2473);
and U2575 (N_2575,N_2470,N_2495);
or U2576 (N_2576,N_2463,N_2469);
xnor U2577 (N_2577,N_2511,N_2482);
nor U2578 (N_2578,N_2470,N_2503);
and U2579 (N_2579,N_2499,N_2487);
and U2580 (N_2580,N_2540,N_2544);
and U2581 (N_2581,N_2554,N_2539);
or U2582 (N_2582,N_2564,N_2528);
nand U2583 (N_2583,N_2521,N_2555);
or U2584 (N_2584,N_2548,N_2547);
nand U2585 (N_2585,N_2573,N_2557);
nand U2586 (N_2586,N_2527,N_2569);
nor U2587 (N_2587,N_2537,N_2561);
xnor U2588 (N_2588,N_2549,N_2568);
or U2589 (N_2589,N_2520,N_2526);
and U2590 (N_2590,N_2536,N_2535);
xnor U2591 (N_2591,N_2534,N_2524);
and U2592 (N_2592,N_2579,N_2530);
nor U2593 (N_2593,N_2577,N_2522);
or U2594 (N_2594,N_2566,N_2543);
xnor U2595 (N_2595,N_2571,N_2572);
and U2596 (N_2596,N_2523,N_2542);
nand U2597 (N_2597,N_2525,N_2532);
xor U2598 (N_2598,N_2550,N_2563);
and U2599 (N_2599,N_2552,N_2565);
xor U2600 (N_2600,N_2529,N_2556);
or U2601 (N_2601,N_2541,N_2551);
or U2602 (N_2602,N_2576,N_2578);
xnor U2603 (N_2603,N_2562,N_2533);
or U2604 (N_2604,N_2574,N_2545);
nor U2605 (N_2605,N_2538,N_2567);
or U2606 (N_2606,N_2559,N_2553);
and U2607 (N_2607,N_2558,N_2560);
and U2608 (N_2608,N_2546,N_2575);
and U2609 (N_2609,N_2570,N_2531);
nor U2610 (N_2610,N_2553,N_2522);
or U2611 (N_2611,N_2526,N_2534);
and U2612 (N_2612,N_2528,N_2521);
xor U2613 (N_2613,N_2523,N_2557);
or U2614 (N_2614,N_2557,N_2535);
or U2615 (N_2615,N_2531,N_2524);
or U2616 (N_2616,N_2522,N_2547);
nand U2617 (N_2617,N_2537,N_2565);
or U2618 (N_2618,N_2550,N_2574);
nor U2619 (N_2619,N_2574,N_2521);
nor U2620 (N_2620,N_2535,N_2551);
and U2621 (N_2621,N_2564,N_2571);
nor U2622 (N_2622,N_2578,N_2570);
and U2623 (N_2623,N_2559,N_2565);
or U2624 (N_2624,N_2574,N_2547);
xnor U2625 (N_2625,N_2542,N_2565);
nor U2626 (N_2626,N_2528,N_2556);
and U2627 (N_2627,N_2552,N_2579);
nand U2628 (N_2628,N_2547,N_2525);
nor U2629 (N_2629,N_2563,N_2526);
and U2630 (N_2630,N_2535,N_2540);
nand U2631 (N_2631,N_2551,N_2528);
and U2632 (N_2632,N_2555,N_2527);
nor U2633 (N_2633,N_2537,N_2578);
and U2634 (N_2634,N_2574,N_2530);
or U2635 (N_2635,N_2572,N_2579);
nand U2636 (N_2636,N_2526,N_2553);
nor U2637 (N_2637,N_2535,N_2530);
and U2638 (N_2638,N_2562,N_2555);
or U2639 (N_2639,N_2576,N_2545);
and U2640 (N_2640,N_2629,N_2590);
or U2641 (N_2641,N_2638,N_2635);
nor U2642 (N_2642,N_2597,N_2585);
and U2643 (N_2643,N_2599,N_2598);
and U2644 (N_2644,N_2587,N_2621);
nor U2645 (N_2645,N_2595,N_2600);
or U2646 (N_2646,N_2619,N_2603);
or U2647 (N_2647,N_2586,N_2620);
xor U2648 (N_2648,N_2612,N_2616);
or U2649 (N_2649,N_2606,N_2580);
or U2650 (N_2650,N_2596,N_2602);
nand U2651 (N_2651,N_2632,N_2634);
and U2652 (N_2652,N_2604,N_2631);
nand U2653 (N_2653,N_2624,N_2614);
or U2654 (N_2654,N_2601,N_2636);
nor U2655 (N_2655,N_2589,N_2610);
nand U2656 (N_2656,N_2615,N_2618);
xnor U2657 (N_2657,N_2583,N_2605);
and U2658 (N_2658,N_2607,N_2639);
nor U2659 (N_2659,N_2581,N_2591);
nand U2660 (N_2660,N_2628,N_2584);
nor U2661 (N_2661,N_2637,N_2630);
nand U2662 (N_2662,N_2611,N_2623);
nor U2663 (N_2663,N_2622,N_2627);
nor U2664 (N_2664,N_2625,N_2582);
nand U2665 (N_2665,N_2613,N_2626);
xnor U2666 (N_2666,N_2594,N_2588);
or U2667 (N_2667,N_2593,N_2633);
nor U2668 (N_2668,N_2617,N_2609);
nor U2669 (N_2669,N_2608,N_2592);
nand U2670 (N_2670,N_2613,N_2602);
or U2671 (N_2671,N_2612,N_2635);
or U2672 (N_2672,N_2581,N_2615);
or U2673 (N_2673,N_2613,N_2624);
and U2674 (N_2674,N_2594,N_2622);
and U2675 (N_2675,N_2605,N_2589);
or U2676 (N_2676,N_2589,N_2599);
nor U2677 (N_2677,N_2613,N_2590);
nand U2678 (N_2678,N_2580,N_2595);
nor U2679 (N_2679,N_2597,N_2632);
xor U2680 (N_2680,N_2597,N_2616);
and U2681 (N_2681,N_2620,N_2613);
nor U2682 (N_2682,N_2594,N_2614);
nor U2683 (N_2683,N_2587,N_2588);
and U2684 (N_2684,N_2597,N_2599);
or U2685 (N_2685,N_2635,N_2625);
nor U2686 (N_2686,N_2611,N_2617);
xnor U2687 (N_2687,N_2625,N_2624);
nand U2688 (N_2688,N_2611,N_2589);
and U2689 (N_2689,N_2606,N_2596);
or U2690 (N_2690,N_2631,N_2591);
xor U2691 (N_2691,N_2584,N_2588);
nand U2692 (N_2692,N_2625,N_2584);
nor U2693 (N_2693,N_2581,N_2584);
and U2694 (N_2694,N_2620,N_2593);
nand U2695 (N_2695,N_2616,N_2624);
and U2696 (N_2696,N_2626,N_2606);
or U2697 (N_2697,N_2634,N_2628);
and U2698 (N_2698,N_2622,N_2628);
nand U2699 (N_2699,N_2602,N_2637);
nor U2700 (N_2700,N_2656,N_2681);
and U2701 (N_2701,N_2658,N_2660);
xor U2702 (N_2702,N_2688,N_2699);
nor U2703 (N_2703,N_2651,N_2669);
and U2704 (N_2704,N_2650,N_2659);
nor U2705 (N_2705,N_2647,N_2646);
nor U2706 (N_2706,N_2640,N_2684);
or U2707 (N_2707,N_2670,N_2666);
nor U2708 (N_2708,N_2678,N_2676);
nand U2709 (N_2709,N_2689,N_2698);
and U2710 (N_2710,N_2655,N_2696);
nor U2711 (N_2711,N_2672,N_2662);
and U2712 (N_2712,N_2641,N_2674);
and U2713 (N_2713,N_2690,N_2673);
nor U2714 (N_2714,N_2675,N_2694);
xor U2715 (N_2715,N_2642,N_2665);
xor U2716 (N_2716,N_2695,N_2677);
nand U2717 (N_2717,N_2671,N_2680);
or U2718 (N_2718,N_2664,N_2654);
or U2719 (N_2719,N_2697,N_2648);
and U2720 (N_2720,N_2686,N_2693);
and U2721 (N_2721,N_2657,N_2663);
nand U2722 (N_2722,N_2645,N_2679);
or U2723 (N_2723,N_2687,N_2644);
nand U2724 (N_2724,N_2692,N_2683);
xor U2725 (N_2725,N_2649,N_2667);
and U2726 (N_2726,N_2652,N_2691);
and U2727 (N_2727,N_2682,N_2685);
nand U2728 (N_2728,N_2668,N_2661);
nor U2729 (N_2729,N_2653,N_2643);
nand U2730 (N_2730,N_2642,N_2685);
xnor U2731 (N_2731,N_2695,N_2670);
and U2732 (N_2732,N_2683,N_2684);
and U2733 (N_2733,N_2648,N_2658);
nand U2734 (N_2734,N_2668,N_2647);
nor U2735 (N_2735,N_2660,N_2648);
nor U2736 (N_2736,N_2671,N_2661);
nand U2737 (N_2737,N_2653,N_2677);
nor U2738 (N_2738,N_2678,N_2694);
and U2739 (N_2739,N_2654,N_2645);
and U2740 (N_2740,N_2648,N_2644);
xnor U2741 (N_2741,N_2648,N_2664);
and U2742 (N_2742,N_2669,N_2644);
and U2743 (N_2743,N_2699,N_2665);
nor U2744 (N_2744,N_2689,N_2660);
nand U2745 (N_2745,N_2685,N_2658);
nand U2746 (N_2746,N_2671,N_2659);
nor U2747 (N_2747,N_2698,N_2674);
nor U2748 (N_2748,N_2694,N_2652);
or U2749 (N_2749,N_2659,N_2645);
and U2750 (N_2750,N_2684,N_2656);
or U2751 (N_2751,N_2663,N_2699);
nor U2752 (N_2752,N_2649,N_2654);
and U2753 (N_2753,N_2661,N_2693);
nor U2754 (N_2754,N_2666,N_2643);
nand U2755 (N_2755,N_2697,N_2658);
nor U2756 (N_2756,N_2675,N_2643);
nor U2757 (N_2757,N_2657,N_2652);
nor U2758 (N_2758,N_2653,N_2693);
nor U2759 (N_2759,N_2682,N_2665);
xor U2760 (N_2760,N_2701,N_2702);
nor U2761 (N_2761,N_2759,N_2730);
xor U2762 (N_2762,N_2725,N_2707);
nor U2763 (N_2763,N_2737,N_2726);
xor U2764 (N_2764,N_2757,N_2749);
and U2765 (N_2765,N_2745,N_2755);
nor U2766 (N_2766,N_2708,N_2742);
nand U2767 (N_2767,N_2716,N_2711);
and U2768 (N_2768,N_2732,N_2743);
nor U2769 (N_2769,N_2719,N_2753);
nor U2770 (N_2770,N_2741,N_2703);
or U2771 (N_2771,N_2712,N_2700);
xnor U2772 (N_2772,N_2724,N_2728);
nor U2773 (N_2773,N_2748,N_2735);
nand U2774 (N_2774,N_2720,N_2739);
nand U2775 (N_2775,N_2709,N_2750);
xnor U2776 (N_2776,N_2722,N_2736);
or U2777 (N_2777,N_2704,N_2733);
and U2778 (N_2778,N_2706,N_2713);
and U2779 (N_2779,N_2731,N_2705);
nor U2780 (N_2780,N_2747,N_2729);
nor U2781 (N_2781,N_2758,N_2718);
nand U2782 (N_2782,N_2717,N_2714);
nand U2783 (N_2783,N_2710,N_2734);
nand U2784 (N_2784,N_2740,N_2723);
nor U2785 (N_2785,N_2738,N_2754);
nor U2786 (N_2786,N_2721,N_2727);
or U2787 (N_2787,N_2715,N_2746);
nor U2788 (N_2788,N_2756,N_2744);
nor U2789 (N_2789,N_2752,N_2751);
and U2790 (N_2790,N_2712,N_2724);
nor U2791 (N_2791,N_2725,N_2708);
nand U2792 (N_2792,N_2718,N_2704);
nand U2793 (N_2793,N_2745,N_2750);
nor U2794 (N_2794,N_2742,N_2753);
or U2795 (N_2795,N_2734,N_2726);
nor U2796 (N_2796,N_2713,N_2710);
nor U2797 (N_2797,N_2750,N_2703);
and U2798 (N_2798,N_2741,N_2752);
nor U2799 (N_2799,N_2716,N_2714);
or U2800 (N_2800,N_2726,N_2751);
or U2801 (N_2801,N_2745,N_2743);
or U2802 (N_2802,N_2716,N_2738);
nor U2803 (N_2803,N_2736,N_2728);
and U2804 (N_2804,N_2711,N_2701);
and U2805 (N_2805,N_2723,N_2722);
or U2806 (N_2806,N_2730,N_2732);
nand U2807 (N_2807,N_2732,N_2736);
or U2808 (N_2808,N_2735,N_2739);
nor U2809 (N_2809,N_2735,N_2740);
and U2810 (N_2810,N_2736,N_2700);
nand U2811 (N_2811,N_2759,N_2755);
or U2812 (N_2812,N_2710,N_2733);
nand U2813 (N_2813,N_2747,N_2759);
or U2814 (N_2814,N_2714,N_2730);
or U2815 (N_2815,N_2758,N_2704);
or U2816 (N_2816,N_2705,N_2710);
nor U2817 (N_2817,N_2746,N_2724);
or U2818 (N_2818,N_2713,N_2721);
nand U2819 (N_2819,N_2752,N_2755);
or U2820 (N_2820,N_2775,N_2781);
nor U2821 (N_2821,N_2800,N_2778);
or U2822 (N_2822,N_2814,N_2787);
nand U2823 (N_2823,N_2799,N_2818);
and U2824 (N_2824,N_2772,N_2807);
xnor U2825 (N_2825,N_2813,N_2768);
nor U2826 (N_2826,N_2760,N_2816);
nand U2827 (N_2827,N_2783,N_2806);
nand U2828 (N_2828,N_2798,N_2802);
and U2829 (N_2829,N_2789,N_2762);
nor U2830 (N_2830,N_2801,N_2808);
nand U2831 (N_2831,N_2780,N_2767);
xor U2832 (N_2832,N_2815,N_2765);
or U2833 (N_2833,N_2786,N_2774);
nor U2834 (N_2834,N_2804,N_2790);
nor U2835 (N_2835,N_2788,N_2764);
nor U2836 (N_2836,N_2817,N_2776);
nor U2837 (N_2837,N_2777,N_2794);
or U2838 (N_2838,N_2770,N_2810);
or U2839 (N_2839,N_2809,N_2784);
nand U2840 (N_2840,N_2812,N_2805);
nor U2841 (N_2841,N_2779,N_2769);
and U2842 (N_2842,N_2763,N_2796);
and U2843 (N_2843,N_2811,N_2797);
nand U2844 (N_2844,N_2785,N_2795);
nor U2845 (N_2845,N_2803,N_2792);
or U2846 (N_2846,N_2773,N_2782);
nor U2847 (N_2847,N_2793,N_2791);
nand U2848 (N_2848,N_2771,N_2761);
or U2849 (N_2849,N_2766,N_2819);
and U2850 (N_2850,N_2790,N_2760);
and U2851 (N_2851,N_2790,N_2788);
and U2852 (N_2852,N_2802,N_2800);
or U2853 (N_2853,N_2802,N_2814);
and U2854 (N_2854,N_2790,N_2786);
or U2855 (N_2855,N_2773,N_2785);
and U2856 (N_2856,N_2795,N_2767);
xnor U2857 (N_2857,N_2798,N_2812);
or U2858 (N_2858,N_2785,N_2799);
nor U2859 (N_2859,N_2812,N_2801);
xor U2860 (N_2860,N_2806,N_2791);
nand U2861 (N_2861,N_2772,N_2780);
or U2862 (N_2862,N_2798,N_2804);
and U2863 (N_2863,N_2805,N_2779);
nand U2864 (N_2864,N_2760,N_2794);
nand U2865 (N_2865,N_2781,N_2760);
and U2866 (N_2866,N_2803,N_2791);
nor U2867 (N_2867,N_2805,N_2819);
and U2868 (N_2868,N_2776,N_2815);
or U2869 (N_2869,N_2809,N_2781);
and U2870 (N_2870,N_2787,N_2799);
nand U2871 (N_2871,N_2796,N_2767);
nor U2872 (N_2872,N_2761,N_2787);
and U2873 (N_2873,N_2810,N_2783);
nand U2874 (N_2874,N_2787,N_2783);
or U2875 (N_2875,N_2817,N_2793);
or U2876 (N_2876,N_2762,N_2791);
nand U2877 (N_2877,N_2806,N_2792);
nand U2878 (N_2878,N_2775,N_2796);
or U2879 (N_2879,N_2793,N_2795);
nand U2880 (N_2880,N_2864,N_2841);
xor U2881 (N_2881,N_2825,N_2822);
nand U2882 (N_2882,N_2859,N_2868);
nand U2883 (N_2883,N_2857,N_2829);
and U2884 (N_2884,N_2858,N_2875);
xnor U2885 (N_2885,N_2834,N_2878);
or U2886 (N_2886,N_2874,N_2836);
nor U2887 (N_2887,N_2837,N_2879);
nand U2888 (N_2888,N_2839,N_2830);
nand U2889 (N_2889,N_2828,N_2851);
nor U2890 (N_2890,N_2850,N_2824);
nand U2891 (N_2891,N_2849,N_2842);
or U2892 (N_2892,N_2826,N_2833);
nand U2893 (N_2893,N_2840,N_2821);
and U2894 (N_2894,N_2867,N_2852);
and U2895 (N_2895,N_2863,N_2847);
or U2896 (N_2896,N_2845,N_2823);
nand U2897 (N_2897,N_2838,N_2848);
or U2898 (N_2898,N_2844,N_2832);
or U2899 (N_2899,N_2827,N_2860);
or U2900 (N_2900,N_2855,N_2831);
nand U2901 (N_2901,N_2843,N_2856);
or U2902 (N_2902,N_2835,N_2820);
nand U2903 (N_2903,N_2853,N_2865);
nor U2904 (N_2904,N_2870,N_2866);
nand U2905 (N_2905,N_2876,N_2861);
or U2906 (N_2906,N_2854,N_2877);
xor U2907 (N_2907,N_2869,N_2873);
and U2908 (N_2908,N_2846,N_2862);
xnor U2909 (N_2909,N_2871,N_2872);
and U2910 (N_2910,N_2848,N_2867);
and U2911 (N_2911,N_2839,N_2841);
nor U2912 (N_2912,N_2874,N_2854);
xor U2913 (N_2913,N_2837,N_2840);
nand U2914 (N_2914,N_2833,N_2842);
and U2915 (N_2915,N_2874,N_2879);
or U2916 (N_2916,N_2857,N_2877);
and U2917 (N_2917,N_2829,N_2860);
nand U2918 (N_2918,N_2833,N_2835);
nor U2919 (N_2919,N_2821,N_2852);
or U2920 (N_2920,N_2869,N_2824);
and U2921 (N_2921,N_2840,N_2879);
and U2922 (N_2922,N_2879,N_2852);
or U2923 (N_2923,N_2864,N_2846);
nor U2924 (N_2924,N_2852,N_2854);
xor U2925 (N_2925,N_2865,N_2846);
and U2926 (N_2926,N_2866,N_2838);
or U2927 (N_2927,N_2869,N_2867);
nor U2928 (N_2928,N_2850,N_2822);
and U2929 (N_2929,N_2833,N_2867);
nor U2930 (N_2930,N_2821,N_2824);
nand U2931 (N_2931,N_2837,N_2833);
or U2932 (N_2932,N_2857,N_2875);
xnor U2933 (N_2933,N_2853,N_2829);
xnor U2934 (N_2934,N_2822,N_2878);
or U2935 (N_2935,N_2863,N_2852);
and U2936 (N_2936,N_2833,N_2852);
and U2937 (N_2937,N_2863,N_2874);
and U2938 (N_2938,N_2823,N_2829);
nand U2939 (N_2939,N_2845,N_2855);
nand U2940 (N_2940,N_2906,N_2891);
nor U2941 (N_2941,N_2925,N_2928);
nor U2942 (N_2942,N_2919,N_2887);
or U2943 (N_2943,N_2911,N_2937);
nand U2944 (N_2944,N_2900,N_2921);
nand U2945 (N_2945,N_2897,N_2924);
and U2946 (N_2946,N_2895,N_2886);
nor U2947 (N_2947,N_2913,N_2883);
nor U2948 (N_2948,N_2894,N_2902);
xor U2949 (N_2949,N_2889,N_2927);
xor U2950 (N_2950,N_2939,N_2916);
nor U2951 (N_2951,N_2930,N_2905);
or U2952 (N_2952,N_2931,N_2885);
nor U2953 (N_2953,N_2932,N_2899);
and U2954 (N_2954,N_2890,N_2907);
nand U2955 (N_2955,N_2920,N_2904);
nor U2956 (N_2956,N_2896,N_2898);
or U2957 (N_2957,N_2908,N_2933);
xnor U2958 (N_2958,N_2912,N_2914);
nand U2959 (N_2959,N_2881,N_2892);
or U2960 (N_2960,N_2903,N_2884);
and U2961 (N_2961,N_2882,N_2918);
nor U2962 (N_2962,N_2917,N_2888);
and U2963 (N_2963,N_2936,N_2909);
and U2964 (N_2964,N_2910,N_2935);
nand U2965 (N_2965,N_2934,N_2893);
nand U2966 (N_2966,N_2901,N_2915);
nand U2967 (N_2967,N_2929,N_2880);
nand U2968 (N_2968,N_2938,N_2923);
and U2969 (N_2969,N_2926,N_2922);
or U2970 (N_2970,N_2933,N_2936);
xnor U2971 (N_2971,N_2894,N_2904);
or U2972 (N_2972,N_2926,N_2933);
or U2973 (N_2973,N_2931,N_2933);
or U2974 (N_2974,N_2881,N_2909);
nor U2975 (N_2975,N_2923,N_2882);
nor U2976 (N_2976,N_2915,N_2917);
xor U2977 (N_2977,N_2917,N_2901);
or U2978 (N_2978,N_2891,N_2923);
nand U2979 (N_2979,N_2880,N_2911);
nor U2980 (N_2980,N_2895,N_2901);
and U2981 (N_2981,N_2925,N_2904);
nand U2982 (N_2982,N_2917,N_2882);
nand U2983 (N_2983,N_2915,N_2911);
and U2984 (N_2984,N_2900,N_2885);
nand U2985 (N_2985,N_2926,N_2916);
and U2986 (N_2986,N_2934,N_2920);
or U2987 (N_2987,N_2919,N_2888);
xor U2988 (N_2988,N_2939,N_2886);
and U2989 (N_2989,N_2887,N_2890);
nand U2990 (N_2990,N_2913,N_2925);
nand U2991 (N_2991,N_2907,N_2886);
nand U2992 (N_2992,N_2901,N_2916);
xnor U2993 (N_2993,N_2927,N_2886);
and U2994 (N_2994,N_2935,N_2889);
or U2995 (N_2995,N_2908,N_2899);
nor U2996 (N_2996,N_2933,N_2906);
xnor U2997 (N_2997,N_2882,N_2884);
or U2998 (N_2998,N_2907,N_2927);
and U2999 (N_2999,N_2920,N_2927);
nor UO_0 (O_0,N_2989,N_2943);
and UO_1 (O_1,N_2941,N_2978);
or UO_2 (O_2,N_2960,N_2991);
nor UO_3 (O_3,N_2948,N_2959);
nand UO_4 (O_4,N_2973,N_2997);
nor UO_5 (O_5,N_2947,N_2969);
nand UO_6 (O_6,N_2988,N_2979);
nand UO_7 (O_7,N_2981,N_2990);
nor UO_8 (O_8,N_2994,N_2985);
and UO_9 (O_9,N_2992,N_2951);
nand UO_10 (O_10,N_2957,N_2964);
or UO_11 (O_11,N_2975,N_2970);
and UO_12 (O_12,N_2955,N_2966);
nand UO_13 (O_13,N_2993,N_2995);
or UO_14 (O_14,N_2956,N_2958);
and UO_15 (O_15,N_2952,N_2977);
nand UO_16 (O_16,N_2963,N_2998);
and UO_17 (O_17,N_2974,N_2949);
and UO_18 (O_18,N_2945,N_2987);
nand UO_19 (O_19,N_2986,N_2982);
and UO_20 (O_20,N_2962,N_2942);
nor UO_21 (O_21,N_2950,N_2983);
and UO_22 (O_22,N_2980,N_2961);
or UO_23 (O_23,N_2946,N_2984);
nor UO_24 (O_24,N_2954,N_2971);
xor UO_25 (O_25,N_2953,N_2976);
or UO_26 (O_26,N_2968,N_2965);
or UO_27 (O_27,N_2972,N_2999);
or UO_28 (O_28,N_2944,N_2996);
xnor UO_29 (O_29,N_2940,N_2967);
nor UO_30 (O_30,N_2955,N_2991);
nand UO_31 (O_31,N_2941,N_2952);
nor UO_32 (O_32,N_2952,N_2975);
xnor UO_33 (O_33,N_2984,N_2959);
or UO_34 (O_34,N_2997,N_2971);
nand UO_35 (O_35,N_2960,N_2949);
nand UO_36 (O_36,N_2993,N_2964);
and UO_37 (O_37,N_2962,N_2989);
and UO_38 (O_38,N_2952,N_2966);
nor UO_39 (O_39,N_2981,N_2942);
nand UO_40 (O_40,N_2965,N_2964);
nand UO_41 (O_41,N_2961,N_2978);
xor UO_42 (O_42,N_2959,N_2994);
and UO_43 (O_43,N_2966,N_2963);
and UO_44 (O_44,N_2985,N_2969);
nor UO_45 (O_45,N_2976,N_2986);
nand UO_46 (O_46,N_2974,N_2942);
or UO_47 (O_47,N_2972,N_2955);
nor UO_48 (O_48,N_2976,N_2969);
nor UO_49 (O_49,N_2953,N_2981);
xor UO_50 (O_50,N_2960,N_2976);
and UO_51 (O_51,N_2963,N_2945);
and UO_52 (O_52,N_2981,N_2943);
nand UO_53 (O_53,N_2940,N_2977);
or UO_54 (O_54,N_2990,N_2966);
nand UO_55 (O_55,N_2958,N_2986);
nor UO_56 (O_56,N_2973,N_2986);
and UO_57 (O_57,N_2999,N_2942);
nor UO_58 (O_58,N_2999,N_2977);
nor UO_59 (O_59,N_2979,N_2941);
xnor UO_60 (O_60,N_2940,N_2956);
and UO_61 (O_61,N_2954,N_2962);
or UO_62 (O_62,N_2952,N_2980);
and UO_63 (O_63,N_2988,N_2984);
and UO_64 (O_64,N_2956,N_2941);
and UO_65 (O_65,N_2966,N_2999);
or UO_66 (O_66,N_2967,N_2957);
nor UO_67 (O_67,N_2968,N_2997);
nand UO_68 (O_68,N_2953,N_2947);
and UO_69 (O_69,N_2978,N_2957);
nand UO_70 (O_70,N_2954,N_2987);
or UO_71 (O_71,N_2972,N_2970);
and UO_72 (O_72,N_2957,N_2947);
xor UO_73 (O_73,N_2994,N_2984);
nor UO_74 (O_74,N_2972,N_2941);
nor UO_75 (O_75,N_2963,N_2962);
or UO_76 (O_76,N_2982,N_2974);
or UO_77 (O_77,N_2981,N_2966);
or UO_78 (O_78,N_2944,N_2988);
and UO_79 (O_79,N_2992,N_2947);
nor UO_80 (O_80,N_2947,N_2998);
and UO_81 (O_81,N_2956,N_2972);
nand UO_82 (O_82,N_2998,N_2976);
nor UO_83 (O_83,N_2957,N_2971);
and UO_84 (O_84,N_2953,N_2970);
nor UO_85 (O_85,N_2973,N_2943);
nand UO_86 (O_86,N_2995,N_2947);
nor UO_87 (O_87,N_2983,N_2973);
and UO_88 (O_88,N_2942,N_2949);
or UO_89 (O_89,N_2969,N_2952);
nand UO_90 (O_90,N_2971,N_2963);
and UO_91 (O_91,N_2958,N_2984);
and UO_92 (O_92,N_2979,N_2975);
and UO_93 (O_93,N_2956,N_2955);
nor UO_94 (O_94,N_2957,N_2987);
nand UO_95 (O_95,N_2955,N_2993);
nor UO_96 (O_96,N_2953,N_2946);
and UO_97 (O_97,N_2963,N_2948);
and UO_98 (O_98,N_2944,N_2984);
nor UO_99 (O_99,N_2956,N_2953);
nand UO_100 (O_100,N_2974,N_2984);
xor UO_101 (O_101,N_2995,N_2944);
nor UO_102 (O_102,N_2966,N_2958);
nor UO_103 (O_103,N_2965,N_2966);
and UO_104 (O_104,N_2985,N_2991);
nor UO_105 (O_105,N_2994,N_2992);
and UO_106 (O_106,N_2961,N_2952);
and UO_107 (O_107,N_2964,N_2952);
nand UO_108 (O_108,N_2967,N_2976);
nor UO_109 (O_109,N_2948,N_2965);
and UO_110 (O_110,N_2947,N_2978);
nand UO_111 (O_111,N_2973,N_2951);
nand UO_112 (O_112,N_2962,N_2970);
nand UO_113 (O_113,N_2958,N_2979);
nand UO_114 (O_114,N_2965,N_2945);
xor UO_115 (O_115,N_2940,N_2958);
or UO_116 (O_116,N_2948,N_2991);
and UO_117 (O_117,N_2956,N_2963);
nor UO_118 (O_118,N_2999,N_2981);
nand UO_119 (O_119,N_2959,N_2947);
nand UO_120 (O_120,N_2965,N_2957);
or UO_121 (O_121,N_2958,N_2996);
or UO_122 (O_122,N_2983,N_2993);
or UO_123 (O_123,N_2966,N_2992);
or UO_124 (O_124,N_2967,N_2942);
nand UO_125 (O_125,N_2970,N_2959);
nor UO_126 (O_126,N_2985,N_2956);
and UO_127 (O_127,N_2964,N_2979);
nand UO_128 (O_128,N_2967,N_2954);
and UO_129 (O_129,N_2983,N_2967);
or UO_130 (O_130,N_2953,N_2975);
or UO_131 (O_131,N_2994,N_2986);
and UO_132 (O_132,N_2980,N_2985);
xnor UO_133 (O_133,N_2981,N_2987);
xor UO_134 (O_134,N_2941,N_2953);
nand UO_135 (O_135,N_2979,N_2967);
nor UO_136 (O_136,N_2974,N_2964);
nor UO_137 (O_137,N_2985,N_2960);
nand UO_138 (O_138,N_2940,N_2994);
or UO_139 (O_139,N_2949,N_2968);
nor UO_140 (O_140,N_2956,N_2990);
or UO_141 (O_141,N_2944,N_2979);
xnor UO_142 (O_142,N_2976,N_2941);
xor UO_143 (O_143,N_2965,N_2974);
nor UO_144 (O_144,N_2978,N_2988);
or UO_145 (O_145,N_2972,N_2973);
nor UO_146 (O_146,N_2997,N_2975);
xor UO_147 (O_147,N_2956,N_2996);
and UO_148 (O_148,N_2961,N_2975);
nand UO_149 (O_149,N_2960,N_2963);
and UO_150 (O_150,N_2950,N_2988);
nor UO_151 (O_151,N_2973,N_2977);
nor UO_152 (O_152,N_2964,N_2950);
xnor UO_153 (O_153,N_2990,N_2971);
nand UO_154 (O_154,N_2946,N_2985);
or UO_155 (O_155,N_2975,N_2966);
and UO_156 (O_156,N_2999,N_2944);
and UO_157 (O_157,N_2965,N_2944);
nor UO_158 (O_158,N_2966,N_2991);
nor UO_159 (O_159,N_2959,N_2991);
nor UO_160 (O_160,N_2977,N_2976);
and UO_161 (O_161,N_2943,N_2945);
nand UO_162 (O_162,N_2989,N_2994);
nor UO_163 (O_163,N_2945,N_2946);
nor UO_164 (O_164,N_2951,N_2977);
nor UO_165 (O_165,N_2978,N_2948);
or UO_166 (O_166,N_2954,N_2975);
and UO_167 (O_167,N_2960,N_2986);
or UO_168 (O_168,N_2980,N_2962);
nor UO_169 (O_169,N_2981,N_2985);
or UO_170 (O_170,N_2996,N_2946);
nand UO_171 (O_171,N_2944,N_2986);
nor UO_172 (O_172,N_2967,N_2994);
or UO_173 (O_173,N_2999,N_2971);
nor UO_174 (O_174,N_2948,N_2979);
nor UO_175 (O_175,N_2942,N_2978);
or UO_176 (O_176,N_2952,N_2949);
and UO_177 (O_177,N_2959,N_2999);
nand UO_178 (O_178,N_2973,N_2980);
and UO_179 (O_179,N_2965,N_2956);
nor UO_180 (O_180,N_2988,N_2976);
or UO_181 (O_181,N_2980,N_2965);
nand UO_182 (O_182,N_2977,N_2974);
and UO_183 (O_183,N_2978,N_2981);
or UO_184 (O_184,N_2975,N_2980);
nor UO_185 (O_185,N_2963,N_2999);
and UO_186 (O_186,N_2998,N_2991);
nand UO_187 (O_187,N_2951,N_2945);
xor UO_188 (O_188,N_2957,N_2980);
nor UO_189 (O_189,N_2946,N_2980);
nor UO_190 (O_190,N_2953,N_2948);
nand UO_191 (O_191,N_2999,N_2948);
nor UO_192 (O_192,N_2984,N_2950);
nand UO_193 (O_193,N_2954,N_2945);
xor UO_194 (O_194,N_2998,N_2944);
or UO_195 (O_195,N_2971,N_2994);
nor UO_196 (O_196,N_2979,N_2953);
nor UO_197 (O_197,N_2953,N_2959);
and UO_198 (O_198,N_2965,N_2962);
or UO_199 (O_199,N_2982,N_2941);
or UO_200 (O_200,N_2962,N_2951);
or UO_201 (O_201,N_2988,N_2954);
or UO_202 (O_202,N_2971,N_2995);
nor UO_203 (O_203,N_2994,N_2969);
nand UO_204 (O_204,N_2950,N_2948);
or UO_205 (O_205,N_2972,N_2992);
and UO_206 (O_206,N_2966,N_2988);
nor UO_207 (O_207,N_2991,N_2942);
or UO_208 (O_208,N_2964,N_2975);
or UO_209 (O_209,N_2975,N_2960);
nor UO_210 (O_210,N_2949,N_2982);
and UO_211 (O_211,N_2957,N_2983);
or UO_212 (O_212,N_2974,N_2952);
nor UO_213 (O_213,N_2949,N_2954);
and UO_214 (O_214,N_2985,N_2982);
nor UO_215 (O_215,N_2994,N_2993);
nand UO_216 (O_216,N_2941,N_2960);
or UO_217 (O_217,N_2969,N_2960);
nand UO_218 (O_218,N_2948,N_2974);
and UO_219 (O_219,N_2941,N_2966);
nor UO_220 (O_220,N_2992,N_2941);
nor UO_221 (O_221,N_2983,N_2990);
and UO_222 (O_222,N_2965,N_2947);
nand UO_223 (O_223,N_2963,N_2967);
nor UO_224 (O_224,N_2948,N_2941);
or UO_225 (O_225,N_2991,N_2970);
nor UO_226 (O_226,N_2952,N_2963);
nand UO_227 (O_227,N_2978,N_2968);
or UO_228 (O_228,N_2993,N_2962);
nor UO_229 (O_229,N_2953,N_2978);
and UO_230 (O_230,N_2959,N_2997);
nand UO_231 (O_231,N_2986,N_2954);
nand UO_232 (O_232,N_2962,N_2957);
xor UO_233 (O_233,N_2943,N_2986);
or UO_234 (O_234,N_2983,N_2970);
or UO_235 (O_235,N_2951,N_2986);
nor UO_236 (O_236,N_2992,N_2957);
nand UO_237 (O_237,N_2941,N_2989);
nand UO_238 (O_238,N_2978,N_2997);
nand UO_239 (O_239,N_2953,N_2989);
and UO_240 (O_240,N_2972,N_2943);
nand UO_241 (O_241,N_2966,N_2961);
nor UO_242 (O_242,N_2999,N_2969);
or UO_243 (O_243,N_2980,N_2995);
and UO_244 (O_244,N_2999,N_2983);
or UO_245 (O_245,N_2984,N_2956);
nand UO_246 (O_246,N_2988,N_2982);
nor UO_247 (O_247,N_2951,N_2979);
and UO_248 (O_248,N_2990,N_2993);
or UO_249 (O_249,N_2963,N_2951);
or UO_250 (O_250,N_2952,N_2998);
nor UO_251 (O_251,N_2965,N_2993);
and UO_252 (O_252,N_2946,N_2975);
or UO_253 (O_253,N_2953,N_2940);
and UO_254 (O_254,N_2942,N_2989);
nand UO_255 (O_255,N_2962,N_2982);
nand UO_256 (O_256,N_2968,N_2996);
or UO_257 (O_257,N_2942,N_2990);
nor UO_258 (O_258,N_2940,N_2970);
nand UO_259 (O_259,N_2992,N_2960);
nand UO_260 (O_260,N_2947,N_2945);
nand UO_261 (O_261,N_2941,N_2957);
nand UO_262 (O_262,N_2958,N_2960);
nand UO_263 (O_263,N_2993,N_2943);
xnor UO_264 (O_264,N_2959,N_2998);
nor UO_265 (O_265,N_2955,N_2951);
nand UO_266 (O_266,N_2965,N_2982);
or UO_267 (O_267,N_2994,N_2976);
or UO_268 (O_268,N_2961,N_2951);
or UO_269 (O_269,N_2963,N_2978);
or UO_270 (O_270,N_2946,N_2993);
and UO_271 (O_271,N_2992,N_2953);
or UO_272 (O_272,N_2963,N_2969);
nand UO_273 (O_273,N_2975,N_2996);
xor UO_274 (O_274,N_2953,N_2943);
and UO_275 (O_275,N_2982,N_2990);
nor UO_276 (O_276,N_2957,N_2942);
nand UO_277 (O_277,N_2991,N_2990);
nand UO_278 (O_278,N_2962,N_2956);
and UO_279 (O_279,N_2969,N_2987);
nor UO_280 (O_280,N_2993,N_2984);
xnor UO_281 (O_281,N_2955,N_2975);
nand UO_282 (O_282,N_2965,N_2953);
nand UO_283 (O_283,N_2960,N_2971);
nand UO_284 (O_284,N_2977,N_2944);
nand UO_285 (O_285,N_2962,N_2985);
nand UO_286 (O_286,N_2978,N_2977);
and UO_287 (O_287,N_2968,N_2974);
or UO_288 (O_288,N_2996,N_2969);
nor UO_289 (O_289,N_2951,N_2987);
or UO_290 (O_290,N_2961,N_2981);
and UO_291 (O_291,N_2956,N_2986);
nor UO_292 (O_292,N_2975,N_2977);
nor UO_293 (O_293,N_2941,N_2959);
and UO_294 (O_294,N_2997,N_2993);
and UO_295 (O_295,N_2951,N_2952);
xnor UO_296 (O_296,N_2967,N_2988);
or UO_297 (O_297,N_2946,N_2983);
nor UO_298 (O_298,N_2992,N_2949);
nand UO_299 (O_299,N_2949,N_2989);
and UO_300 (O_300,N_2992,N_2975);
and UO_301 (O_301,N_2951,N_2975);
and UO_302 (O_302,N_2942,N_2940);
nor UO_303 (O_303,N_2941,N_2996);
or UO_304 (O_304,N_2967,N_2980);
nor UO_305 (O_305,N_2957,N_2999);
nor UO_306 (O_306,N_2968,N_2986);
or UO_307 (O_307,N_2942,N_2956);
nand UO_308 (O_308,N_2970,N_2954);
or UO_309 (O_309,N_2984,N_2952);
nand UO_310 (O_310,N_2958,N_2949);
nor UO_311 (O_311,N_2959,N_2966);
or UO_312 (O_312,N_2942,N_2984);
nand UO_313 (O_313,N_2982,N_2989);
nor UO_314 (O_314,N_2975,N_2957);
and UO_315 (O_315,N_2982,N_2975);
nor UO_316 (O_316,N_2997,N_2944);
nand UO_317 (O_317,N_2995,N_2942);
or UO_318 (O_318,N_2987,N_2948);
and UO_319 (O_319,N_2949,N_2953);
nand UO_320 (O_320,N_2948,N_2967);
nor UO_321 (O_321,N_2957,N_2954);
nand UO_322 (O_322,N_2959,N_2957);
or UO_323 (O_323,N_2994,N_2968);
and UO_324 (O_324,N_2990,N_2961);
or UO_325 (O_325,N_2955,N_2980);
xor UO_326 (O_326,N_2956,N_2997);
nand UO_327 (O_327,N_2999,N_2984);
and UO_328 (O_328,N_2958,N_2981);
or UO_329 (O_329,N_2968,N_2971);
nor UO_330 (O_330,N_2962,N_2967);
nand UO_331 (O_331,N_2941,N_2993);
or UO_332 (O_332,N_2975,N_2985);
nor UO_333 (O_333,N_2995,N_2998);
xor UO_334 (O_334,N_2947,N_2990);
or UO_335 (O_335,N_2998,N_2992);
or UO_336 (O_336,N_2945,N_2969);
nand UO_337 (O_337,N_2983,N_2980);
and UO_338 (O_338,N_2946,N_2971);
or UO_339 (O_339,N_2948,N_2992);
or UO_340 (O_340,N_2989,N_2957);
nor UO_341 (O_341,N_2982,N_2964);
xnor UO_342 (O_342,N_2999,N_2976);
xnor UO_343 (O_343,N_2976,N_2995);
nand UO_344 (O_344,N_2962,N_2988);
and UO_345 (O_345,N_2998,N_2946);
nand UO_346 (O_346,N_2994,N_2978);
or UO_347 (O_347,N_2979,N_2985);
xor UO_348 (O_348,N_2977,N_2960);
xnor UO_349 (O_349,N_2981,N_2993);
and UO_350 (O_350,N_2990,N_2970);
or UO_351 (O_351,N_2977,N_2957);
or UO_352 (O_352,N_2956,N_2957);
nor UO_353 (O_353,N_2989,N_2961);
nand UO_354 (O_354,N_2966,N_2967);
nand UO_355 (O_355,N_2990,N_2962);
and UO_356 (O_356,N_2979,N_2970);
and UO_357 (O_357,N_2980,N_2972);
nand UO_358 (O_358,N_2993,N_2986);
or UO_359 (O_359,N_2983,N_2966);
nand UO_360 (O_360,N_2962,N_2973);
and UO_361 (O_361,N_2997,N_2995);
nor UO_362 (O_362,N_2971,N_2992);
nand UO_363 (O_363,N_2981,N_2976);
nor UO_364 (O_364,N_2941,N_2964);
or UO_365 (O_365,N_2971,N_2976);
and UO_366 (O_366,N_2975,N_2976);
nand UO_367 (O_367,N_2976,N_2962);
and UO_368 (O_368,N_2942,N_2960);
xor UO_369 (O_369,N_2964,N_2971);
and UO_370 (O_370,N_2953,N_2995);
nand UO_371 (O_371,N_2985,N_2948);
nand UO_372 (O_372,N_2948,N_2962);
nand UO_373 (O_373,N_2980,N_2976);
or UO_374 (O_374,N_2971,N_2986);
nand UO_375 (O_375,N_2946,N_2955);
nand UO_376 (O_376,N_2986,N_2974);
nand UO_377 (O_377,N_2971,N_2947);
nor UO_378 (O_378,N_2952,N_2991);
xnor UO_379 (O_379,N_2995,N_2967);
nand UO_380 (O_380,N_2951,N_2954);
xor UO_381 (O_381,N_2960,N_2967);
nor UO_382 (O_382,N_2963,N_2944);
nor UO_383 (O_383,N_2989,N_2998);
nand UO_384 (O_384,N_2972,N_2979);
or UO_385 (O_385,N_2947,N_2940);
nand UO_386 (O_386,N_2979,N_2945);
nand UO_387 (O_387,N_2951,N_2947);
xor UO_388 (O_388,N_2986,N_2942);
or UO_389 (O_389,N_2992,N_2976);
nand UO_390 (O_390,N_2960,N_2996);
and UO_391 (O_391,N_2950,N_2990);
or UO_392 (O_392,N_2957,N_2945);
nor UO_393 (O_393,N_2989,N_2952);
nor UO_394 (O_394,N_2982,N_2946);
nand UO_395 (O_395,N_2968,N_2987);
and UO_396 (O_396,N_2974,N_2976);
and UO_397 (O_397,N_2964,N_2999);
nor UO_398 (O_398,N_2972,N_2984);
or UO_399 (O_399,N_2955,N_2997);
or UO_400 (O_400,N_2999,N_2946);
nand UO_401 (O_401,N_2953,N_2991);
and UO_402 (O_402,N_2996,N_2985);
nor UO_403 (O_403,N_2946,N_2972);
and UO_404 (O_404,N_2971,N_2969);
nor UO_405 (O_405,N_2999,N_2941);
or UO_406 (O_406,N_2971,N_2940);
nand UO_407 (O_407,N_2948,N_2986);
and UO_408 (O_408,N_2950,N_2940);
or UO_409 (O_409,N_2977,N_2958);
and UO_410 (O_410,N_2991,N_2993);
and UO_411 (O_411,N_2970,N_2969);
or UO_412 (O_412,N_2984,N_2947);
or UO_413 (O_413,N_2962,N_2974);
nor UO_414 (O_414,N_2962,N_2964);
and UO_415 (O_415,N_2996,N_2999);
xor UO_416 (O_416,N_2962,N_2972);
nand UO_417 (O_417,N_2987,N_2978);
xor UO_418 (O_418,N_2954,N_2969);
nor UO_419 (O_419,N_2947,N_2989);
nand UO_420 (O_420,N_2943,N_2940);
nand UO_421 (O_421,N_2989,N_2974);
nand UO_422 (O_422,N_2998,N_2954);
nor UO_423 (O_423,N_2968,N_2960);
or UO_424 (O_424,N_2958,N_2963);
nand UO_425 (O_425,N_2975,N_2941);
nor UO_426 (O_426,N_2967,N_2990);
nand UO_427 (O_427,N_2972,N_2944);
and UO_428 (O_428,N_2975,N_2988);
nor UO_429 (O_429,N_2998,N_2957);
nand UO_430 (O_430,N_2989,N_2997);
and UO_431 (O_431,N_2970,N_2981);
nor UO_432 (O_432,N_2993,N_2953);
nand UO_433 (O_433,N_2971,N_2989);
and UO_434 (O_434,N_2993,N_2958);
nor UO_435 (O_435,N_2992,N_2990);
nor UO_436 (O_436,N_2981,N_2960);
nor UO_437 (O_437,N_2989,N_2954);
or UO_438 (O_438,N_2977,N_2985);
and UO_439 (O_439,N_2961,N_2987);
or UO_440 (O_440,N_2993,N_2960);
nand UO_441 (O_441,N_2985,N_2951);
nor UO_442 (O_442,N_2940,N_2976);
nor UO_443 (O_443,N_2977,N_2969);
and UO_444 (O_444,N_2948,N_2952);
or UO_445 (O_445,N_2976,N_2970);
and UO_446 (O_446,N_2960,N_2946);
or UO_447 (O_447,N_2977,N_2964);
or UO_448 (O_448,N_2967,N_2953);
or UO_449 (O_449,N_2992,N_2961);
nand UO_450 (O_450,N_2972,N_2994);
and UO_451 (O_451,N_2960,N_2974);
or UO_452 (O_452,N_2996,N_2986);
nand UO_453 (O_453,N_2952,N_2978);
or UO_454 (O_454,N_2995,N_2970);
nor UO_455 (O_455,N_2988,N_2968);
nor UO_456 (O_456,N_2940,N_2974);
and UO_457 (O_457,N_2997,N_2964);
nor UO_458 (O_458,N_2989,N_2948);
nand UO_459 (O_459,N_2951,N_2941);
xor UO_460 (O_460,N_2972,N_2997);
xnor UO_461 (O_461,N_2956,N_2946);
nor UO_462 (O_462,N_2957,N_2984);
xnor UO_463 (O_463,N_2997,N_2994);
or UO_464 (O_464,N_2980,N_2994);
nand UO_465 (O_465,N_2978,N_2999);
nand UO_466 (O_466,N_2990,N_2954);
nor UO_467 (O_467,N_2944,N_2955);
and UO_468 (O_468,N_2947,N_2960);
nand UO_469 (O_469,N_2983,N_2992);
and UO_470 (O_470,N_2950,N_2996);
or UO_471 (O_471,N_2985,N_2989);
or UO_472 (O_472,N_2979,N_2965);
nor UO_473 (O_473,N_2959,N_2976);
nor UO_474 (O_474,N_2963,N_2973);
xnor UO_475 (O_475,N_2991,N_2962);
or UO_476 (O_476,N_2986,N_2997);
nand UO_477 (O_477,N_2965,N_2958);
or UO_478 (O_478,N_2962,N_2961);
nor UO_479 (O_479,N_2982,N_2943);
and UO_480 (O_480,N_2997,N_2996);
and UO_481 (O_481,N_2989,N_2973);
nor UO_482 (O_482,N_2962,N_2943);
or UO_483 (O_483,N_2978,N_2998);
and UO_484 (O_484,N_2943,N_2999);
xor UO_485 (O_485,N_2943,N_2963);
nand UO_486 (O_486,N_2990,N_2969);
nor UO_487 (O_487,N_2940,N_2946);
and UO_488 (O_488,N_2946,N_2941);
and UO_489 (O_489,N_2945,N_2970);
xnor UO_490 (O_490,N_2972,N_2974);
or UO_491 (O_491,N_2966,N_2948);
and UO_492 (O_492,N_2991,N_2983);
and UO_493 (O_493,N_2964,N_2988);
and UO_494 (O_494,N_2940,N_2993);
nor UO_495 (O_495,N_2987,N_2994);
or UO_496 (O_496,N_2951,N_2966);
nor UO_497 (O_497,N_2953,N_2997);
or UO_498 (O_498,N_2982,N_2972);
or UO_499 (O_499,N_2983,N_2996);
endmodule