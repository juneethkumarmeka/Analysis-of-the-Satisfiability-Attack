module basic_2000_20000_2500_4_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_1977,In_690);
nor U1 (N_1,In_1197,In_852);
and U2 (N_2,In_337,In_1524);
nor U3 (N_3,In_1292,In_1113);
or U4 (N_4,In_1559,In_181);
and U5 (N_5,In_282,In_1152);
nand U6 (N_6,In_727,In_360);
or U7 (N_7,In_890,In_7);
or U8 (N_8,In_1675,In_1624);
and U9 (N_9,In_18,In_1746);
or U10 (N_10,In_80,In_233);
or U11 (N_11,In_31,In_914);
nor U12 (N_12,In_1264,In_1852);
nor U13 (N_13,In_630,In_1778);
and U14 (N_14,In_1328,In_757);
nand U15 (N_15,In_920,In_1057);
or U16 (N_16,In_759,In_715);
nor U17 (N_17,In_1375,In_626);
nor U18 (N_18,In_1296,In_1828);
and U19 (N_19,In_332,In_32);
and U20 (N_20,In_45,In_1698);
and U21 (N_21,In_1514,In_202);
or U22 (N_22,In_216,In_1003);
or U23 (N_23,In_604,In_53);
nor U24 (N_24,In_717,In_389);
or U25 (N_25,In_1859,In_1067);
nand U26 (N_26,In_450,In_1616);
nor U27 (N_27,In_1034,In_1135);
or U28 (N_28,In_427,In_1918);
nand U29 (N_29,In_64,In_83);
and U30 (N_30,In_811,In_721);
and U31 (N_31,In_818,In_873);
and U32 (N_32,In_409,In_1081);
or U33 (N_33,In_1826,In_1767);
nor U34 (N_34,In_1325,In_240);
nand U35 (N_35,In_290,In_194);
nor U36 (N_36,In_1434,In_1192);
and U37 (N_37,In_997,In_1405);
and U38 (N_38,In_959,In_1769);
or U39 (N_39,In_203,In_1992);
or U40 (N_40,In_613,In_1509);
nand U41 (N_41,In_1127,In_1409);
or U42 (N_42,In_590,In_1215);
or U43 (N_43,In_99,In_636);
nor U44 (N_44,In_1044,In_1773);
or U45 (N_45,In_1202,In_658);
nor U46 (N_46,In_243,In_1100);
and U47 (N_47,In_505,In_131);
and U48 (N_48,In_769,In_909);
or U49 (N_49,In_230,In_605);
nand U50 (N_50,In_1586,In_860);
and U51 (N_51,In_583,In_1048);
nand U52 (N_52,In_1390,In_783);
and U53 (N_53,In_264,In_1200);
nand U54 (N_54,In_795,In_758);
or U55 (N_55,In_1936,In_1742);
or U56 (N_56,In_536,In_1686);
nor U57 (N_57,In_1201,In_1695);
nand U58 (N_58,In_1145,In_1752);
or U59 (N_59,In_1950,In_1275);
nor U60 (N_60,In_1897,In_513);
and U61 (N_61,In_159,In_1149);
nand U62 (N_62,In_534,In_654);
and U63 (N_63,In_1761,In_1782);
nand U64 (N_64,In_382,In_1133);
nand U65 (N_65,In_1089,In_29);
or U66 (N_66,In_415,In_241);
nor U67 (N_67,In_1819,In_761);
nand U68 (N_68,In_963,In_1534);
nand U69 (N_69,In_51,In_455);
nor U70 (N_70,In_888,In_842);
and U71 (N_71,In_1199,In_1435);
nor U72 (N_72,In_1234,In_350);
nor U73 (N_73,In_1533,In_1723);
nor U74 (N_74,In_1455,In_1472);
or U75 (N_75,In_1013,In_220);
or U76 (N_76,In_1531,In_82);
or U77 (N_77,In_516,In_1049);
nand U78 (N_78,In_796,In_1912);
nor U79 (N_79,In_1810,In_1353);
and U80 (N_80,In_1261,In_1357);
nand U81 (N_81,In_1453,In_958);
nand U82 (N_82,In_1942,In_1254);
nand U83 (N_83,In_1232,In_40);
and U84 (N_84,In_591,In_74);
and U85 (N_85,In_416,In_1456);
and U86 (N_86,In_1310,In_1799);
and U87 (N_87,In_1317,In_1573);
nor U88 (N_88,In_856,In_140);
nor U89 (N_89,In_88,In_1816);
nor U90 (N_90,In_195,In_84);
nand U91 (N_91,In_487,In_1344);
nor U92 (N_92,In_1653,In_1278);
and U93 (N_93,In_610,In_479);
nor U94 (N_94,In_933,In_1667);
or U95 (N_95,In_169,In_1106);
and U96 (N_96,In_770,In_1258);
nor U97 (N_97,In_1737,In_1471);
nand U98 (N_98,In_1934,In_1512);
nand U99 (N_99,In_1743,In_1022);
or U100 (N_100,In_1063,In_1439);
and U101 (N_101,In_1478,In_1703);
nand U102 (N_102,In_907,In_547);
nand U103 (N_103,In_1958,In_1403);
nand U104 (N_104,In_1733,In_42);
nand U105 (N_105,In_1907,In_1715);
or U106 (N_106,In_270,In_541);
nor U107 (N_107,In_1558,In_805);
and U108 (N_108,In_582,In_296);
nand U109 (N_109,In_452,In_1447);
or U110 (N_110,In_647,In_947);
or U111 (N_111,In_1805,In_47);
or U112 (N_112,In_261,In_1727);
and U113 (N_113,In_1792,In_787);
nor U114 (N_114,In_932,In_369);
or U115 (N_115,In_135,In_1652);
and U116 (N_116,In_968,In_639);
or U117 (N_117,In_388,In_1881);
or U118 (N_118,In_1648,In_120);
nand U119 (N_119,In_1763,In_408);
nor U120 (N_120,In_85,In_1047);
or U121 (N_121,In_27,In_407);
nand U122 (N_122,In_186,In_735);
nor U123 (N_123,In_1917,In_661);
and U124 (N_124,In_1143,In_372);
nand U125 (N_125,In_1502,In_1130);
nor U126 (N_126,In_98,In_112);
and U127 (N_127,In_437,In_979);
nor U128 (N_128,In_1785,In_297);
and U129 (N_129,In_1422,In_1158);
or U130 (N_130,In_293,In_697);
or U131 (N_131,In_1326,In_329);
and U132 (N_132,In_859,In_1822);
nand U133 (N_133,In_1346,In_574);
nand U134 (N_134,In_865,In_1104);
and U135 (N_135,In_1968,In_1380);
nand U136 (N_136,In_231,In_4);
or U137 (N_137,In_1015,In_1736);
and U138 (N_138,In_1486,In_1361);
nand U139 (N_139,In_786,In_916);
nand U140 (N_140,In_1632,In_1233);
and U141 (N_141,In_1775,In_1645);
nor U142 (N_142,In_1592,In_1026);
or U143 (N_143,In_726,In_1869);
xor U144 (N_144,In_1076,In_866);
or U145 (N_145,In_1321,In_70);
nand U146 (N_146,In_995,In_503);
or U147 (N_147,In_1208,In_1914);
nand U148 (N_148,In_941,In_899);
and U149 (N_149,In_791,In_820);
and U150 (N_150,In_1239,In_1451);
and U151 (N_151,In_724,In_280);
nor U152 (N_152,In_1381,In_309);
nor U153 (N_153,In_105,In_1838);
and U154 (N_154,In_1561,In_746);
nand U155 (N_155,In_1322,In_43);
and U156 (N_156,In_1760,In_922);
nor U157 (N_157,In_964,In_921);
or U158 (N_158,In_1285,In_77);
nand U159 (N_159,In_592,In_1072);
nand U160 (N_160,In_21,In_1904);
nor U161 (N_161,In_570,In_1448);
and U162 (N_162,In_872,In_1011);
and U163 (N_163,In_227,In_609);
and U164 (N_164,In_133,In_566);
nor U165 (N_165,In_1943,In_1386);
nor U166 (N_166,In_1873,In_1277);
nand U167 (N_167,In_138,In_1610);
or U168 (N_168,In_573,In_1609);
nand U169 (N_169,In_1488,In_1498);
nor U170 (N_170,In_716,In_784);
and U171 (N_171,In_1101,In_723);
or U172 (N_172,In_1755,In_1295);
nor U173 (N_173,In_734,In_560);
and U174 (N_174,In_1781,In_1622);
nor U175 (N_175,In_700,In_1569);
and U176 (N_176,In_1438,In_468);
and U177 (N_177,In_238,In_720);
nor U178 (N_178,In_355,In_1832);
nand U179 (N_179,In_1814,In_1466);
nand U180 (N_180,In_1168,In_550);
nand U181 (N_181,In_641,In_540);
and U182 (N_182,In_1287,In_575);
and U183 (N_183,In_126,In_1696);
or U184 (N_184,In_1906,In_1383);
and U185 (N_185,In_1801,In_1568);
nand U186 (N_186,In_1867,In_1139);
nand U187 (N_187,In_1378,In_586);
and U188 (N_188,In_823,In_1046);
and U189 (N_189,In_1465,In_1181);
nand U190 (N_190,In_1148,In_1399);
nor U191 (N_191,In_1180,In_308);
nor U192 (N_192,In_363,In_67);
or U193 (N_193,In_300,In_1855);
nor U194 (N_194,In_59,In_1087);
and U195 (N_195,In_1679,In_1583);
and U196 (N_196,In_1175,In_508);
or U197 (N_197,In_917,In_197);
or U198 (N_198,In_136,In_1210);
or U199 (N_199,In_1817,In_1074);
and U200 (N_200,In_1613,In_793);
and U201 (N_201,In_1699,In_587);
and U202 (N_202,In_1646,In_165);
and U203 (N_203,In_1019,In_666);
and U204 (N_204,In_502,In_563);
nor U205 (N_205,In_391,In_1999);
or U206 (N_206,In_49,In_1473);
nor U207 (N_207,In_901,In_1213);
nor U208 (N_208,In_785,In_274);
or U209 (N_209,In_497,In_63);
and U210 (N_210,In_1997,In_1820);
or U211 (N_211,In_306,In_310);
nand U212 (N_212,In_434,In_1896);
nor U213 (N_213,In_928,In_714);
and U214 (N_214,In_1341,In_1915);
and U215 (N_215,In_210,In_777);
nand U216 (N_216,In_361,In_910);
nand U217 (N_217,In_1280,In_1260);
and U218 (N_218,In_1706,In_753);
nor U219 (N_219,In_188,In_1387);
or U220 (N_220,In_827,In_1132);
and U221 (N_221,In_638,In_1187);
nand U222 (N_222,In_1824,In_413);
nor U223 (N_223,In_1732,In_289);
nor U224 (N_224,In_1449,In_1605);
nor U225 (N_225,In_285,In_1627);
or U226 (N_226,In_1982,In_196);
nor U227 (N_227,In_473,In_1614);
nor U228 (N_228,In_1097,In_26);
nor U229 (N_229,In_421,In_453);
nor U230 (N_230,In_527,In_1602);
nor U231 (N_231,In_464,In_1415);
nand U232 (N_232,In_1579,In_1671);
or U233 (N_233,In_1861,In_1229);
nand U234 (N_234,In_66,In_529);
and U235 (N_235,In_1137,In_1880);
nand U236 (N_236,In_960,In_1482);
nand U237 (N_237,In_564,In_1198);
nor U238 (N_238,In_1410,In_1928);
nor U239 (N_239,In_295,In_376);
or U240 (N_240,In_1414,In_162);
or U241 (N_241,In_1521,In_358);
and U242 (N_242,In_632,In_668);
or U243 (N_243,In_1241,In_1253);
nand U244 (N_244,In_810,In_1617);
nand U245 (N_245,In_606,In_1166);
xnor U246 (N_246,In_1582,In_1659);
nor U247 (N_247,In_1900,In_885);
and U248 (N_248,In_1281,In_1837);
and U249 (N_249,In_1790,In_1697);
or U250 (N_250,In_1297,In_1885);
nand U251 (N_251,In_1165,In_36);
nor U252 (N_252,In_903,In_871);
nand U253 (N_253,In_850,In_199);
or U254 (N_254,In_30,In_713);
nand U255 (N_255,In_1980,In_837);
nand U256 (N_256,In_118,In_849);
nor U257 (N_257,In_366,In_1910);
or U258 (N_258,In_139,In_1476);
or U259 (N_259,In_620,In_1227);
or U260 (N_260,In_596,In_906);
or U261 (N_261,In_3,In_33);
nand U262 (N_262,In_478,In_443);
nand U263 (N_263,In_1384,In_1772);
nand U264 (N_264,In_184,In_1464);
and U265 (N_265,In_1669,In_1660);
nor U266 (N_266,In_480,In_1474);
and U267 (N_267,In_870,In_1511);
nor U268 (N_268,In_1901,In_1331);
or U269 (N_269,In_1176,In_1847);
nor U270 (N_270,In_1726,In_1445);
nand U271 (N_271,In_1560,In_1195);
and U272 (N_272,In_1062,In_1787);
and U273 (N_273,In_167,In_1487);
or U274 (N_274,In_891,In_103);
nor U275 (N_275,In_262,In_631);
or U276 (N_276,In_803,In_340);
and U277 (N_277,In_749,In_333);
nand U278 (N_278,In_384,In_245);
and U279 (N_279,In_652,In_1043);
nand U280 (N_280,In_648,In_213);
and U281 (N_281,In_545,In_904);
nand U282 (N_282,In_380,In_1017);
nor U283 (N_283,In_678,In_1189);
nor U284 (N_284,In_371,In_1251);
and U285 (N_285,In_78,In_940);
nand U286 (N_286,In_1944,In_313);
nand U287 (N_287,In_535,In_1834);
nand U288 (N_288,In_23,In_318);
or U289 (N_289,In_108,In_304);
nand U290 (N_290,In_130,In_562);
nor U291 (N_291,In_403,In_284);
nor U292 (N_292,In_1758,In_322);
and U293 (N_293,In_1956,In_1762);
or U294 (N_294,In_250,In_1348);
or U295 (N_295,In_945,In_331);
and U296 (N_296,In_599,In_552);
and U297 (N_297,In_1818,In_1557);
and U298 (N_298,In_429,In_68);
nand U299 (N_299,In_1364,In_211);
or U300 (N_300,In_1507,In_578);
nand U301 (N_301,In_1739,In_38);
or U302 (N_302,In_1985,In_1981);
nand U303 (N_303,In_1173,In_279);
or U304 (N_304,In_1032,In_905);
nor U305 (N_305,In_303,In_488);
nor U306 (N_306,In_19,In_1593);
and U307 (N_307,In_1946,In_191);
or U308 (N_308,In_1940,In_92);
nor U309 (N_309,In_1935,In_1400);
or U310 (N_310,In_1116,In_1150);
nand U311 (N_311,In_396,In_1721);
nor U312 (N_312,In_368,In_1874);
or U313 (N_313,In_1536,In_160);
nor U314 (N_314,In_1108,In_1857);
and U315 (N_315,In_1407,In_344);
nor U316 (N_316,In_1007,In_671);
or U317 (N_317,In_973,In_1725);
nand U318 (N_318,In_462,In_204);
and U319 (N_319,In_1843,In_39);
nand U320 (N_320,In_1257,In_1349);
or U321 (N_321,In_686,In_778);
nand U322 (N_322,In_209,In_1294);
nor U323 (N_323,In_1099,In_1962);
nand U324 (N_324,In_1941,In_1329);
and U325 (N_325,In_1903,In_37);
and U326 (N_326,In_822,In_76);
or U327 (N_327,In_834,In_1242);
or U328 (N_328,In_25,In_1244);
nor U329 (N_329,In_315,In_1355);
and U330 (N_330,In_1225,In_1978);
or U331 (N_331,In_766,In_1182);
nand U332 (N_332,In_1418,In_383);
nand U333 (N_333,In_266,In_1926);
and U334 (N_334,In_660,In_1938);
nor U335 (N_335,In_1639,In_1491);
or U336 (N_336,In_519,In_1800);
nand U337 (N_337,In_861,In_1895);
nor U338 (N_338,In_1061,In_773);
and U339 (N_339,In_1996,In_1649);
and U340 (N_340,In_998,In_347);
or U341 (N_341,In_1423,In_373);
nor U342 (N_342,In_397,In_1306);
and U343 (N_343,In_9,In_615);
and U344 (N_344,In_1892,In_386);
or U345 (N_345,In_176,In_674);
or U346 (N_346,In_673,In_732);
nor U347 (N_347,In_755,In_1821);
nand U348 (N_348,In_980,In_1735);
nor U349 (N_349,In_433,In_524);
nand U350 (N_350,In_565,In_225);
nand U351 (N_351,In_1126,In_526);
or U352 (N_352,In_1630,In_1028);
and U353 (N_353,In_460,In_1332);
nor U354 (N_354,In_628,In_1879);
nor U355 (N_355,In_426,In_588);
and U356 (N_356,In_431,In_1899);
nand U357 (N_357,In_1898,In_1641);
nand U358 (N_358,In_1179,In_679);
and U359 (N_359,In_1095,In_1394);
or U360 (N_360,In_926,In_708);
nand U361 (N_361,In_161,In_1663);
or U362 (N_362,In_212,In_1309);
nand U363 (N_363,In_1483,In_50);
or U364 (N_364,In_249,In_612);
or U365 (N_365,In_463,In_692);
and U366 (N_366,In_694,In_1690);
or U367 (N_367,In_1428,In_1395);
or U368 (N_368,In_477,In_1077);
nand U369 (N_369,In_28,In_869);
nor U370 (N_370,In_493,In_1995);
and U371 (N_371,In_1856,In_15);
and U372 (N_372,In_1604,In_1922);
nand U373 (N_373,In_1052,In_966);
nor U374 (N_374,In_857,In_1849);
and U375 (N_375,In_1111,In_1413);
nand U376 (N_376,In_934,In_1658);
nand U377 (N_377,In_342,In_22);
and U378 (N_378,In_1780,In_1256);
or U379 (N_379,In_754,In_878);
nor U380 (N_380,In_1994,In_874);
nor U381 (N_381,In_1685,In_1759);
nor U382 (N_382,In_1594,In_771);
nor U383 (N_383,In_1267,In_614);
nand U384 (N_384,In_1987,In_772);
nand U385 (N_385,In_762,In_494);
and U386 (N_386,In_518,In_515);
nor U387 (N_387,In_1655,In_1636);
or U388 (N_388,In_908,In_466);
and U389 (N_389,In_1041,In_406);
and U390 (N_390,In_307,In_137);
and U391 (N_391,In_1584,In_619);
and U392 (N_392,In_1872,In_10);
or U393 (N_393,In_804,In_830);
nand U394 (N_394,In_931,In_634);
nand U395 (N_395,In_1114,In_1998);
nor U396 (N_396,In_1038,In_1957);
or U397 (N_397,In_1556,In_110);
nand U398 (N_398,In_589,In_1450);
or U399 (N_399,In_1845,In_242);
or U400 (N_400,In_799,In_1206);
and U401 (N_401,In_467,In_1530);
and U402 (N_402,In_115,In_1091);
nor U403 (N_403,In_894,In_672);
nor U404 (N_404,In_1343,In_236);
nor U405 (N_405,In_1515,In_1420);
and U406 (N_406,In_1283,In_1719);
nor U407 (N_407,In_846,In_1083);
nor U408 (N_408,In_442,In_1298);
or U409 (N_409,In_430,In_353);
nor U410 (N_410,In_577,In_767);
nand U411 (N_411,In_1628,In_999);
nor U412 (N_412,In_269,In_247);
nand U413 (N_413,In_1866,In_509);
or U414 (N_414,In_61,In_1314);
nor U415 (N_415,In_978,In_445);
or U416 (N_416,In_1036,In_258);
and U417 (N_417,In_760,In_316);
or U418 (N_418,In_1598,In_168);
nor U419 (N_419,In_663,In_1868);
nor U420 (N_420,In_1815,In_207);
or U421 (N_421,In_1337,In_1651);
nor U422 (N_422,In_221,In_967);
nor U423 (N_423,In_292,In_1554);
nand U424 (N_424,In_1124,In_1220);
nand U425 (N_425,In_600,In_379);
and U426 (N_426,In_1286,In_1608);
nor U427 (N_427,In_736,In_288);
nor U428 (N_428,In_1147,In_670);
nor U429 (N_429,In_1537,In_312);
and U430 (N_430,In_1027,In_375);
and U431 (N_431,In_1211,In_496);
or U432 (N_432,In_1118,In_1002);
nand U433 (N_433,In_879,In_323);
or U434 (N_434,In_35,In_1754);
or U435 (N_435,In_1004,In_395);
and U436 (N_436,In_733,In_449);
nor U437 (N_437,In_1372,In_1983);
nor U438 (N_438,In_1446,In_788);
or U439 (N_439,In_1831,In_1960);
or U440 (N_440,In_677,In_1071);
nand U441 (N_441,In_265,In_1427);
nor U442 (N_442,In_1416,In_1272);
nand U443 (N_443,In_977,In_1209);
and U444 (N_444,In_1676,In_1722);
xnor U445 (N_445,In_1268,In_553);
nand U446 (N_446,In_601,In_511);
nor U447 (N_447,In_2,In_402);
or U448 (N_448,In_1082,In_370);
nand U449 (N_449,In_438,In_929);
or U450 (N_450,In_393,In_46);
nand U451 (N_451,In_1237,In_341);
nor U452 (N_452,In_1990,In_401);
and U453 (N_453,In_1745,In_75);
nand U454 (N_454,In_228,In_1094);
nor U455 (N_455,In_1485,In_798);
and U456 (N_456,In_171,In_1633);
nand U457 (N_457,In_1389,In_1597);
nor U458 (N_458,In_1040,In_1545);
nand U459 (N_459,In_1231,In_1882);
nor U460 (N_460,In_593,In_1704);
and U461 (N_461,In_259,In_179);
or U462 (N_462,In_1039,In_157);
or U463 (N_463,In_569,In_1001);
and U464 (N_464,In_1562,In_1);
nand U465 (N_465,In_1905,In_1481);
nor U466 (N_466,In_1734,In_198);
and U467 (N_467,In_1005,In_1884);
nor U468 (N_468,In_1406,In_1964);
and U469 (N_469,In_554,In_832);
nor U470 (N_470,In_504,In_1248);
nand U471 (N_471,In_166,In_79);
or U472 (N_472,In_436,In_1069);
and U473 (N_473,In_1316,In_1029);
and U474 (N_474,In_1933,In_868);
and U475 (N_475,In_208,In_1647);
nand U476 (N_476,In_471,In_1526);
or U477 (N_477,In_1334,In_1952);
nor U478 (N_478,In_1894,In_706);
nand U479 (N_479,In_522,In_1305);
nor U480 (N_480,In_1783,In_528);
and U481 (N_481,In_1365,In_1454);
and U482 (N_482,In_399,In_1771);
or U483 (N_483,In_1975,In_1469);
and U484 (N_484,In_1984,In_1269);
nor U485 (N_485,In_1270,In_1382);
and U486 (N_486,In_768,In_1496);
nor U487 (N_487,In_1953,In_546);
nand U488 (N_488,In_1080,In_498);
nand U489 (N_489,In_1188,In_918);
and U490 (N_490,In_338,In_988);
nor U491 (N_491,In_52,In_913);
nand U492 (N_492,In_655,In_17);
and U493 (N_493,In_603,In_1535);
or U494 (N_494,In_1924,In_1596);
or U495 (N_495,In_561,In_656);
or U496 (N_496,In_1865,In_1327);
and U497 (N_497,In_1738,In_792);
nor U498 (N_498,In_1065,In_1571);
or U499 (N_499,In_1419,In_440);
or U500 (N_500,In_1932,In_702);
nor U501 (N_501,In_993,In_1342);
nand U502 (N_502,In_5,In_1490);
nand U503 (N_503,In_1190,In_567);
or U504 (N_504,In_495,In_930);
nand U505 (N_505,In_117,In_183);
and U506 (N_506,In_1204,In_1988);
and U507 (N_507,In_177,In_483);
or U508 (N_508,In_1105,In_1177);
nand U509 (N_509,In_622,In_1131);
nor U510 (N_510,In_283,In_886);
and U511 (N_511,In_1276,In_1479);
and U512 (N_512,In_1740,In_150);
nand U513 (N_513,In_537,In_273);
nand U514 (N_514,In_972,In_954);
nor U515 (N_515,In_863,In_847);
and U516 (N_516,In_1833,In_1073);
nor U517 (N_517,In_1844,In_481);
nand U518 (N_518,In_1461,In_1523);
and U519 (N_519,In_1169,In_1250);
nand U520 (N_520,In_1058,In_1525);
nor U521 (N_521,In_1347,In_1290);
or U522 (N_522,In_1666,In_1713);
and U523 (N_523,In_824,In_938);
and U524 (N_524,In_517,In_902);
nand U525 (N_525,In_398,In_145);
or U526 (N_526,In_836,In_114);
and U527 (N_527,In_1923,In_1452);
nor U528 (N_528,In_974,In_1302);
nor U529 (N_529,In_689,In_356);
xnor U530 (N_530,In_812,In_629);
or U531 (N_531,In_1979,In_829);
nand U532 (N_532,In_1858,In_1408);
nor U533 (N_533,In_643,In_946);
nor U534 (N_534,In_1635,In_1689);
and U535 (N_535,In_1566,In_1803);
or U536 (N_536,In_1282,In_1494);
nand U537 (N_537,In_965,In_1522);
nand U538 (N_538,In_625,In_328);
nor U539 (N_539,In_953,In_800);
nor U540 (N_540,In_113,In_1037);
nand U541 (N_541,In_132,In_1018);
or U542 (N_542,In_214,In_255);
nor U543 (N_543,In_555,In_205);
and U544 (N_544,In_1330,In_835);
nor U545 (N_545,In_394,In_143);
and U546 (N_546,In_659,In_925);
or U547 (N_547,In_164,In_111);
nor U548 (N_548,In_982,In_844);
xnor U549 (N_549,In_1807,In_525);
and U550 (N_550,In_69,In_173);
nor U551 (N_551,In_1788,In_201);
nand U552 (N_552,In_1110,In_1945);
and U553 (N_553,In_531,In_1708);
and U554 (N_554,In_1350,In_608);
nor U555 (N_555,In_1437,In_1541);
or U556 (N_556,In_542,In_1318);
nor U557 (N_557,In_144,In_994);
nand U558 (N_558,In_301,In_1644);
nand U559 (N_559,In_1768,In_1710);
nor U560 (N_560,In_1020,In_252);
nor U561 (N_561,In_699,In_1966);
and U562 (N_562,In_1576,In_1141);
and U563 (N_563,In_633,In_490);
nand U564 (N_564,In_48,In_1460);
nor U565 (N_565,In_1623,In_877);
nor U566 (N_566,In_731,In_549);
and U567 (N_567,In_1731,In_971);
and U568 (N_568,In_653,In_1489);
nand U569 (N_569,In_175,In_937);
and U570 (N_570,In_1823,In_1379);
nor U571 (N_571,In_1546,In_667);
or U572 (N_572,In_1714,In_1430);
nand U573 (N_573,In_825,In_275);
nand U574 (N_574,In_148,In_1010);
nor U575 (N_575,In_662,In_1115);
nand U576 (N_576,In_1811,In_153);
or U577 (N_577,In_1528,In_246);
and U578 (N_578,In_1969,In_983);
nor U579 (N_579,In_244,In_428);
and U580 (N_580,In_680,In_1508);
nor U581 (N_581,In_801,In_1552);
nor U582 (N_582,In_691,In_345);
or U583 (N_583,In_883,In_665);
or U584 (N_584,In_302,In_1911);
and U585 (N_585,In_1307,In_1841);
nor U586 (N_586,In_1955,In_1581);
nor U587 (N_587,In_14,In_501);
and U588 (N_588,In_234,In_1404);
and U589 (N_589,In_1068,In_875);
or U590 (N_590,In_1516,In_1757);
nand U591 (N_591,In_54,In_743);
and U592 (N_592,In_1411,In_1219);
nand U593 (N_593,In_1851,In_750);
nor U594 (N_594,In_390,In_335);
or U595 (N_595,In_1519,In_927);
nor U596 (N_596,In_645,In_1889);
nor U597 (N_597,In_617,In_1477);
nand U598 (N_598,In_1230,In_1398);
or U599 (N_599,In_459,In_119);
and U600 (N_600,In_1023,In_1886);
nand U601 (N_601,In_34,In_1377);
nand U602 (N_602,In_1064,In_712);
nor U603 (N_603,In_1796,In_1376);
nand U604 (N_604,In_124,In_97);
or U605 (N_605,In_155,In_1144);
and U606 (N_606,In_1919,In_1207);
nor U607 (N_607,In_675,In_400);
nor U608 (N_608,In_1262,In_1876);
and U609 (N_609,In_1304,In_1517);
and U610 (N_610,In_984,In_95);
nand U611 (N_611,In_1595,In_0);
nor U612 (N_612,In_597,In_1888);
and U613 (N_613,In_802,In_89);
or U614 (N_614,In_1544,In_1354);
or U615 (N_615,In_20,In_752);
or U616 (N_616,In_81,In_1954);
or U617 (N_617,In_486,In_1112);
nor U618 (N_618,In_1504,In_1656);
and U619 (N_619,In_1591,In_192);
and U620 (N_620,In_412,In_991);
nand U621 (N_621,In_55,In_1678);
or U622 (N_622,In_738,In_319);
nor U623 (N_623,In_1025,In_1436);
or U624 (N_624,In_414,In_419);
nor U625 (N_625,In_684,In_949);
and U626 (N_626,In_172,In_405);
or U627 (N_627,In_441,In_816);
and U628 (N_628,In_327,In_90);
nor U629 (N_629,In_330,In_1939);
nor U630 (N_630,In_1887,In_1682);
nor U631 (N_631,In_808,In_944);
or U632 (N_632,In_1243,In_651);
and U633 (N_633,In_1902,In_8);
and U634 (N_634,In_544,In_1315);
nand U635 (N_635,In_719,In_521);
nor U636 (N_636,In_1059,In_41);
and U637 (N_637,In_1585,In_789);
or U638 (N_638,In_271,In_1967);
and U639 (N_639,In_701,In_1860);
nand U640 (N_640,In_896,In_1850);
and U641 (N_641,In_476,In_568);
and U642 (N_642,In_1812,In_410);
nand U643 (N_643,In_1443,In_1288);
nor U644 (N_644,In_1520,In_739);
nand U645 (N_645,In_475,In_1532);
or U646 (N_646,In_900,In_1716);
or U647 (N_647,In_737,In_1640);
and U648 (N_648,In_1756,In_657);
or U649 (N_649,In_951,In_882);
nand U650 (N_650,In_1564,In_623);
and U651 (N_651,In_1134,In_1335);
or U652 (N_652,In_1086,In_1748);
or U653 (N_653,In_1893,In_1674);
nand U654 (N_654,In_1661,In_1078);
and U655 (N_655,In_334,In_1673);
nor U656 (N_656,In_354,In_1683);
nor U657 (N_657,In_1273,In_1947);
nand U658 (N_658,In_100,In_1770);
or U659 (N_659,In_1146,In_1301);
xor U660 (N_660,In_611,In_532);
and U661 (N_661,In_1122,In_1601);
nand U662 (N_662,In_1016,In_461);
or U663 (N_663,In_87,In_1421);
nor U664 (N_664,In_745,In_1138);
nor U665 (N_665,In_147,In_1553);
nor U666 (N_666,In_189,In_650);
and U667 (N_667,In_1631,In_248);
nor U668 (N_668,In_321,In_1412);
nand U669 (N_669,In_294,In_1589);
nand U670 (N_670,In_851,In_1223);
nor U671 (N_671,In_1170,In_742);
or U672 (N_672,In_484,In_1587);
xor U673 (N_673,In_833,In_359);
nor U674 (N_674,In_239,In_491);
or U675 (N_675,In_897,In_765);
nor U676 (N_676,In_1970,In_13);
nor U677 (N_677,In_1650,In_728);
and U678 (N_678,In_580,In_1747);
or U679 (N_679,In_447,In_1749);
nor U680 (N_680,In_598,In_1864);
and U681 (N_681,In_1468,In_1929);
or U682 (N_682,In_1777,In_1707);
and U683 (N_683,In_952,In_813);
nor U684 (N_684,In_1371,In_1961);
or U685 (N_685,In_418,In_1266);
nand U686 (N_686,In_1324,In_365);
nand U687 (N_687,In_1129,In_1462);
nor U688 (N_688,In_705,In_1991);
nor U689 (N_689,In_1396,In_1538);
or U690 (N_690,In_451,In_1366);
nor U691 (N_691,In_1654,In_1429);
nand U692 (N_692,In_1240,In_1764);
or U693 (N_693,In_1670,In_1164);
nand U694 (N_694,In_1042,In_1840);
or U695 (N_695,In_424,In_392);
nor U696 (N_696,In_985,In_158);
or U697 (N_697,In_385,In_956);
or U698 (N_698,In_1701,In_780);
and U699 (N_699,In_506,In_709);
nor U700 (N_700,In_1878,In_1320);
or U701 (N_701,In_336,In_992);
nor U702 (N_702,In_190,In_936);
or U703 (N_703,In_439,In_747);
or U704 (N_704,In_1174,In_1615);
or U705 (N_705,In_1931,In_1927);
nor U706 (N_706,In_1031,In_814);
nor U707 (N_707,In_1259,In_725);
nor U708 (N_708,In_180,In_128);
nor U709 (N_709,In_1588,In_1090);
nand U710 (N_710,In_343,In_1637);
and U711 (N_711,In_1388,In_1795);
nand U712 (N_712,In_91,In_1128);
nand U713 (N_713,In_1830,In_1352);
nor U714 (N_714,In_807,In_235);
and U715 (N_715,In_718,In_1774);
or U716 (N_716,In_579,In_1684);
and U717 (N_717,In_423,In_698);
xor U718 (N_718,In_326,In_1600);
nand U719 (N_719,In_1070,In_1513);
nor U720 (N_720,In_311,In_1779);
nand U721 (N_721,In_1662,In_1440);
nand U722 (N_722,In_123,In_1643);
nand U723 (N_723,In_122,In_1629);
and U724 (N_724,In_1875,In_935);
and U725 (N_725,In_1093,In_815);
and U726 (N_726,In_790,In_219);
or U727 (N_727,In_57,In_848);
or U728 (N_728,In_520,In_1319);
and U729 (N_729,In_1555,In_1724);
and U730 (N_730,In_915,In_710);
nand U731 (N_731,In_538,In_1096);
nand U732 (N_732,In_895,In_1625);
and U733 (N_733,In_1235,In_1103);
nor U734 (N_734,In_149,In_425);
nor U735 (N_735,In_939,In_1311);
nand U736 (N_736,In_581,In_551);
nand U737 (N_737,In_1373,In_756);
and U738 (N_738,In_912,In_1539);
nor U739 (N_739,In_1730,In_1501);
nand U740 (N_740,In_602,In_1107);
nand U741 (N_741,In_1236,In_1360);
or U742 (N_742,In_1527,In_1368);
nor U743 (N_743,In_1842,In_256);
nand U744 (N_744,In_1692,In_986);
nor U745 (N_745,In_156,In_1060);
and U746 (N_746,In_11,In_585);
nor U747 (N_747,In_106,In_1603);
or U748 (N_748,In_1853,In_683);
and U749 (N_749,In_1299,In_1444);
nand U750 (N_750,In_1391,In_298);
and U751 (N_751,In_253,In_1565);
nor U752 (N_752,In_1274,In_305);
or U753 (N_753,In_1681,In_187);
nor U754 (N_754,In_996,In_387);
and U755 (N_755,In_73,In_748);
and U756 (N_756,In_685,In_1336);
nand U757 (N_757,In_1580,In_222);
nor U758 (N_758,In_1493,In_1045);
nand U759 (N_759,In_107,In_775);
or U760 (N_760,In_446,In_1621);
nand U761 (N_761,In_1687,In_854);
and U762 (N_762,In_1863,In_499);
and U763 (N_763,In_1224,In_1765);
or U764 (N_764,In_1247,In_955);
nor U765 (N_765,In_1829,In_840);
and U766 (N_766,In_1442,In_1351);
nor U767 (N_767,In_741,In_16);
nor U768 (N_768,In_981,In_1323);
or U769 (N_769,In_6,In_989);
nor U770 (N_770,In_1374,In_1949);
nor U771 (N_771,In_1217,In_1463);
nor U772 (N_772,In_1252,In_558);
nand U773 (N_773,In_893,In_146);
and U774 (N_774,In_530,In_1634);
nor U775 (N_775,In_969,In_1599);
nor U776 (N_776,In_272,In_1951);
and U777 (N_777,In_1289,In_1255);
nand U778 (N_778,In_1221,In_1618);
nor U779 (N_779,In_1218,In_1030);
and U780 (N_780,In_1789,In_200);
or U781 (N_781,In_1680,In_1672);
nor U782 (N_782,In_843,In_1203);
or U783 (N_783,In_1154,In_1470);
nand U784 (N_784,In_223,In_1467);
or U785 (N_785,In_740,In_1393);
nor U786 (N_786,In_1839,In_1156);
or U787 (N_787,In_559,In_1974);
or U788 (N_788,In_1121,In_1109);
nor U789 (N_789,In_217,In_12);
and U790 (N_790,In_1877,In_1212);
nand U791 (N_791,In_1191,In_1709);
nand U792 (N_792,In_1854,In_1424);
nor U793 (N_793,In_1657,In_1677);
and U794 (N_794,In_1033,In_377);
or U795 (N_795,In_1009,In_1161);
nand U796 (N_796,In_1798,In_276);
or U797 (N_797,In_1973,In_1510);
and U798 (N_798,In_1125,In_1356);
nand U799 (N_799,In_182,In_1426);
nor U800 (N_800,In_828,In_422);
or U801 (N_801,In_96,In_1862);
nor U802 (N_802,In_696,In_1367);
or U803 (N_803,In_1171,In_942);
nor U804 (N_804,In_1809,In_1293);
or U805 (N_805,In_571,In_364);
nor U806 (N_806,In_1620,In_267);
nor U807 (N_807,In_1055,In_1920);
or U808 (N_808,In_1162,In_432);
or U809 (N_809,In_711,In_1263);
and U810 (N_810,In_474,In_1540);
or U811 (N_811,In_510,In_1908);
nand U812 (N_812,In_1155,In_1808);
nor U813 (N_813,In_693,In_839);
and U814 (N_814,In_1542,In_961);
nor U815 (N_815,In_892,In_987);
and U816 (N_816,In_1729,In_635);
and U817 (N_817,In_1612,In_60);
nand U818 (N_818,In_1417,In_1786);
nor U819 (N_819,In_1205,In_729);
and U820 (N_820,In_287,In_251);
nor U821 (N_821,In_1891,In_1385);
and U822 (N_822,In_1702,In_1784);
or U823 (N_823,In_1157,In_821);
nor U824 (N_824,In_806,In_1500);
nor U825 (N_825,In_224,In_470);
nand U826 (N_826,In_1806,In_1228);
and U827 (N_827,In_1433,In_781);
xnor U828 (N_828,In_776,In_1153);
nand U829 (N_829,In_794,In_193);
nor U830 (N_830,In_1606,In_1216);
nand U831 (N_831,In_142,In_154);
nand U832 (N_832,In_1567,In_378);
nand U833 (N_833,In_970,In_444);
nor U834 (N_834,In_676,In_819);
nand U835 (N_835,In_1303,In_456);
nor U836 (N_836,In_817,In_1345);
nor U837 (N_837,In_512,In_924);
nand U838 (N_838,In_174,In_637);
or U839 (N_839,In_1976,In_62);
or U840 (N_840,In_1948,In_232);
and U841 (N_841,In_838,In_576);
nor U842 (N_842,In_72,In_1728);
or U843 (N_843,In_86,In_492);
nor U844 (N_844,In_1549,In_352);
nor U845 (N_845,In_1214,In_1120);
nor U846 (N_846,In_1163,In_1459);
nand U847 (N_847,In_1271,In_1827);
nor U848 (N_848,In_1705,In_1457);
or U849 (N_849,In_1505,In_642);
and U850 (N_850,In_1123,In_1397);
and U851 (N_851,In_557,In_109);
nor U852 (N_852,In_898,In_1959);
and U853 (N_853,In_595,In_1265);
nor U854 (N_854,In_948,In_411);
and U855 (N_855,In_71,In_1021);
nor U856 (N_856,In_349,In_257);
nor U857 (N_857,In_357,In_703);
nand U858 (N_858,In_514,In_975);
or U859 (N_859,In_624,In_1720);
and U860 (N_860,In_572,In_1909);
or U861 (N_861,In_314,In_1117);
or U862 (N_862,In_889,In_1401);
and U863 (N_863,In_1186,In_24);
or U864 (N_864,In_93,In_845);
nor U865 (N_865,In_779,In_1506);
and U866 (N_866,In_58,In_646);
nand U867 (N_867,In_1054,In_1804);
or U868 (N_868,In_1547,In_695);
or U869 (N_869,In_1313,In_320);
and U870 (N_870,In_1921,In_1712);
and U871 (N_871,In_435,In_1503);
or U872 (N_872,In_621,In_881);
nand U873 (N_873,In_1751,In_1193);
nor U874 (N_874,In_482,In_163);
nand U875 (N_875,In_454,In_1196);
nand U876 (N_876,In_730,In_911);
and U877 (N_877,In_260,In_887);
or U878 (N_878,In_1590,In_764);
nor U879 (N_879,In_1151,In_1750);
nand U880 (N_880,In_1245,In_485);
and U881 (N_881,In_1766,In_226);
nor U882 (N_882,In_797,In_500);
nor U883 (N_883,In_1965,In_1551);
nor U884 (N_884,In_1392,In_1136);
nand U885 (N_885,In_1238,In_325);
nor U886 (N_886,In_1333,In_1084);
and U887 (N_887,In_1989,In_465);
nand U888 (N_888,In_826,In_127);
and U889 (N_889,In_864,In_351);
nor U890 (N_890,In_1279,In_1871);
or U891 (N_891,In_858,In_1711);
or U892 (N_892,In_1012,In_1870);
and U893 (N_893,In_374,In_1363);
and U894 (N_894,In_1492,In_649);
or U895 (N_895,In_417,In_281);
nand U896 (N_896,In_134,In_681);
nor U897 (N_897,In_867,In_1339);
or U898 (N_898,In_1053,In_1548);
nor U899 (N_899,In_1300,In_65);
nand U900 (N_900,In_1194,In_1688);
or U901 (N_901,In_704,In_277);
nor U902 (N_902,In_1358,In_121);
or U903 (N_903,In_616,In_556);
or U904 (N_904,In_1008,In_1066);
and U905 (N_905,In_215,In_774);
nor U906 (N_906,In_1529,In_254);
nor U907 (N_907,In_862,In_339);
nand U908 (N_908,In_751,In_129);
or U909 (N_909,In_1668,In_94);
nand U910 (N_910,In_1495,In_152);
nor U911 (N_911,In_627,In_1518);
or U912 (N_912,In_1665,In_1085);
nand U913 (N_913,In_185,In_1051);
nand U914 (N_914,In_1890,In_489);
nand U915 (N_915,In_1431,In_880);
or U916 (N_916,In_218,In_404);
or U917 (N_917,In_141,In_278);
nor U918 (N_918,In_782,In_1993);
and U919 (N_919,In_1693,In_1226);
and U920 (N_920,In_607,In_957);
and U921 (N_921,In_1575,In_1543);
nand U922 (N_922,In_1425,In_1813);
nor U923 (N_923,In_44,In_853);
and U924 (N_924,In_1338,In_299);
nor U925 (N_925,In_1611,In_170);
or U926 (N_926,In_1184,In_286);
nand U927 (N_927,In_1572,In_809);
nand U928 (N_928,In_990,In_1183);
nand U929 (N_929,In_1312,In_1370);
nand U930 (N_930,In_229,In_458);
nor U931 (N_931,In_1835,In_543);
or U932 (N_932,In_1846,In_687);
or U933 (N_933,In_1972,In_640);
nand U934 (N_934,In_104,In_1480);
nand U935 (N_935,In_457,In_263);
and U936 (N_936,In_1802,In_1000);
or U937 (N_937,In_1432,In_1578);
nand U938 (N_938,In_1797,In_1475);
nand U939 (N_939,In_101,In_1291);
nor U940 (N_940,In_1717,In_664);
nand U941 (N_941,In_1402,In_1925);
nand U942 (N_942,In_317,In_539);
or U943 (N_943,In_1718,In_1056);
nor U944 (N_944,In_1497,In_1550);
nor U945 (N_945,In_707,In_56);
nand U946 (N_946,In_876,In_644);
nand U947 (N_947,In_1642,In_831);
or U948 (N_948,In_1744,In_125);
and U949 (N_949,In_682,In_923);
nor U950 (N_950,In_1916,In_1913);
nand U951 (N_951,In_1222,In_1638);
nor U952 (N_952,In_1119,In_548);
or U953 (N_953,In_1793,In_1574);
or U954 (N_954,In_1825,In_1249);
nand U955 (N_955,In_523,In_1626);
nor U956 (N_956,In_943,In_1741);
nor U957 (N_957,In_584,In_1092);
or U958 (N_958,In_618,In_976);
and U959 (N_959,In_722,In_1050);
nand U960 (N_960,In_116,In_1178);
nor U961 (N_961,In_1185,In_1691);
nand U962 (N_962,In_1340,In_919);
nor U963 (N_963,In_1577,In_1006);
nor U964 (N_964,In_1458,In_1499);
nand U965 (N_965,In_1563,In_950);
or U966 (N_966,In_1484,In_1986);
and U967 (N_967,In_962,In_324);
nor U968 (N_968,In_1791,In_1308);
nand U969 (N_969,In_884,In_268);
and U970 (N_970,In_472,In_469);
or U971 (N_971,In_1963,In_1883);
or U972 (N_972,In_420,In_206);
nand U973 (N_973,In_1014,In_669);
nor U974 (N_974,In_1088,In_367);
nor U975 (N_975,In_102,In_1619);
nor U976 (N_976,In_237,In_291);
and U977 (N_977,In_1776,In_151);
nor U978 (N_978,In_1930,In_1359);
nand U979 (N_979,In_1098,In_1024);
nand U980 (N_980,In_1441,In_533);
or U981 (N_981,In_841,In_1836);
nand U982 (N_982,In_1246,In_1035);
and U983 (N_983,In_1694,In_763);
or U984 (N_984,In_1167,In_744);
nor U985 (N_985,In_1664,In_1753);
nor U986 (N_986,In_1369,In_507);
nor U987 (N_987,In_1159,In_362);
or U988 (N_988,In_1362,In_1794);
nand U989 (N_989,In_348,In_688);
or U990 (N_990,In_178,In_346);
or U991 (N_991,In_1570,In_1140);
or U992 (N_992,In_1142,In_1102);
and U993 (N_993,In_448,In_1848);
nand U994 (N_994,In_1160,In_1700);
nand U995 (N_995,In_1607,In_1937);
nand U996 (N_996,In_1079,In_1284);
nor U997 (N_997,In_1075,In_1172);
nand U998 (N_998,In_855,In_381);
nand U999 (N_999,In_1971,In_594);
nand U1000 (N_1000,In_1327,In_1298);
or U1001 (N_1001,In_191,In_1166);
nor U1002 (N_1002,In_1227,In_1765);
nor U1003 (N_1003,In_1205,In_1671);
or U1004 (N_1004,In_575,In_914);
nand U1005 (N_1005,In_1113,In_911);
or U1006 (N_1006,In_1749,In_166);
nand U1007 (N_1007,In_861,In_243);
nand U1008 (N_1008,In_240,In_1998);
nand U1009 (N_1009,In_1078,In_1961);
nor U1010 (N_1010,In_964,In_698);
or U1011 (N_1011,In_1899,In_854);
and U1012 (N_1012,In_1994,In_883);
nand U1013 (N_1013,In_1390,In_1149);
nor U1014 (N_1014,In_1439,In_927);
and U1015 (N_1015,In_623,In_1366);
nand U1016 (N_1016,In_1792,In_662);
nand U1017 (N_1017,In_821,In_1026);
nand U1018 (N_1018,In_1093,In_694);
and U1019 (N_1019,In_1449,In_253);
nand U1020 (N_1020,In_537,In_1862);
and U1021 (N_1021,In_406,In_477);
or U1022 (N_1022,In_1471,In_1947);
nor U1023 (N_1023,In_439,In_1189);
nand U1024 (N_1024,In_604,In_272);
nor U1025 (N_1025,In_220,In_1316);
and U1026 (N_1026,In_1027,In_246);
nand U1027 (N_1027,In_989,In_1603);
nand U1028 (N_1028,In_392,In_25);
nand U1029 (N_1029,In_626,In_1872);
or U1030 (N_1030,In_686,In_1504);
and U1031 (N_1031,In_629,In_695);
nand U1032 (N_1032,In_893,In_644);
or U1033 (N_1033,In_712,In_1700);
or U1034 (N_1034,In_1800,In_204);
and U1035 (N_1035,In_1277,In_1863);
nand U1036 (N_1036,In_271,In_566);
nand U1037 (N_1037,In_153,In_499);
nor U1038 (N_1038,In_989,In_258);
nand U1039 (N_1039,In_882,In_979);
nor U1040 (N_1040,In_354,In_1917);
nor U1041 (N_1041,In_1827,In_719);
nand U1042 (N_1042,In_1712,In_567);
or U1043 (N_1043,In_944,In_1836);
and U1044 (N_1044,In_1136,In_57);
or U1045 (N_1045,In_1560,In_801);
or U1046 (N_1046,In_1377,In_4);
or U1047 (N_1047,In_1379,In_748);
and U1048 (N_1048,In_498,In_1031);
and U1049 (N_1049,In_1447,In_1543);
nor U1050 (N_1050,In_1125,In_1556);
or U1051 (N_1051,In_1965,In_1711);
nand U1052 (N_1052,In_1469,In_1904);
nand U1053 (N_1053,In_1870,In_345);
xnor U1054 (N_1054,In_36,In_616);
and U1055 (N_1055,In_262,In_24);
or U1056 (N_1056,In_282,In_1951);
and U1057 (N_1057,In_1428,In_1150);
and U1058 (N_1058,In_1128,In_271);
or U1059 (N_1059,In_309,In_1041);
or U1060 (N_1060,In_1798,In_245);
nor U1061 (N_1061,In_998,In_1501);
and U1062 (N_1062,In_1048,In_1477);
or U1063 (N_1063,In_494,In_350);
nand U1064 (N_1064,In_291,In_317);
nand U1065 (N_1065,In_1076,In_1208);
or U1066 (N_1066,In_1769,In_1928);
xor U1067 (N_1067,In_1538,In_196);
nand U1068 (N_1068,In_951,In_1541);
or U1069 (N_1069,In_472,In_1777);
nor U1070 (N_1070,In_1861,In_63);
nor U1071 (N_1071,In_1832,In_168);
and U1072 (N_1072,In_1111,In_529);
nand U1073 (N_1073,In_1595,In_765);
and U1074 (N_1074,In_1312,In_1216);
or U1075 (N_1075,In_1211,In_1761);
or U1076 (N_1076,In_86,In_1228);
and U1077 (N_1077,In_34,In_766);
nor U1078 (N_1078,In_1027,In_1196);
nor U1079 (N_1079,In_880,In_1753);
and U1080 (N_1080,In_545,In_945);
nor U1081 (N_1081,In_1335,In_1515);
or U1082 (N_1082,In_1208,In_1163);
nor U1083 (N_1083,In_630,In_1814);
nor U1084 (N_1084,In_1610,In_1387);
or U1085 (N_1085,In_1484,In_1366);
nand U1086 (N_1086,In_140,In_252);
or U1087 (N_1087,In_42,In_325);
nor U1088 (N_1088,In_551,In_1868);
and U1089 (N_1089,In_1653,In_1133);
nand U1090 (N_1090,In_1854,In_204);
nand U1091 (N_1091,In_1111,In_216);
nand U1092 (N_1092,In_146,In_854);
nand U1093 (N_1093,In_1844,In_155);
nand U1094 (N_1094,In_669,In_1264);
nor U1095 (N_1095,In_428,In_200);
and U1096 (N_1096,In_1171,In_699);
nor U1097 (N_1097,In_1758,In_501);
nand U1098 (N_1098,In_1725,In_660);
nand U1099 (N_1099,In_381,In_1134);
nand U1100 (N_1100,In_1996,In_367);
nor U1101 (N_1101,In_760,In_166);
and U1102 (N_1102,In_1203,In_1880);
nor U1103 (N_1103,In_187,In_433);
nor U1104 (N_1104,In_1200,In_1508);
nand U1105 (N_1105,In_687,In_1978);
nor U1106 (N_1106,In_536,In_362);
or U1107 (N_1107,In_1917,In_1887);
nor U1108 (N_1108,In_1295,In_40);
nand U1109 (N_1109,In_1491,In_969);
nor U1110 (N_1110,In_601,In_67);
nor U1111 (N_1111,In_106,In_1167);
nor U1112 (N_1112,In_1796,In_1201);
nand U1113 (N_1113,In_1284,In_309);
and U1114 (N_1114,In_1620,In_1936);
and U1115 (N_1115,In_1662,In_1371);
and U1116 (N_1116,In_1858,In_903);
and U1117 (N_1117,In_1086,In_1512);
and U1118 (N_1118,In_1135,In_722);
nand U1119 (N_1119,In_328,In_794);
nand U1120 (N_1120,In_1857,In_64);
or U1121 (N_1121,In_439,In_1395);
or U1122 (N_1122,In_672,In_1170);
nor U1123 (N_1123,In_1297,In_456);
nor U1124 (N_1124,In_794,In_736);
and U1125 (N_1125,In_917,In_383);
nor U1126 (N_1126,In_172,In_1432);
nor U1127 (N_1127,In_480,In_1661);
and U1128 (N_1128,In_1862,In_1242);
xor U1129 (N_1129,In_952,In_1434);
and U1130 (N_1130,In_1579,In_337);
nor U1131 (N_1131,In_1545,In_351);
and U1132 (N_1132,In_265,In_1057);
nand U1133 (N_1133,In_1672,In_66);
nand U1134 (N_1134,In_1880,In_1279);
nor U1135 (N_1135,In_1125,In_479);
nand U1136 (N_1136,In_732,In_1236);
and U1137 (N_1137,In_1755,In_1574);
and U1138 (N_1138,In_758,In_452);
and U1139 (N_1139,In_1001,In_919);
and U1140 (N_1140,In_1582,In_1199);
nand U1141 (N_1141,In_146,In_1963);
or U1142 (N_1142,In_1173,In_79);
nor U1143 (N_1143,In_686,In_501);
or U1144 (N_1144,In_580,In_741);
or U1145 (N_1145,In_494,In_1178);
and U1146 (N_1146,In_144,In_1030);
or U1147 (N_1147,In_1649,In_104);
or U1148 (N_1148,In_99,In_1334);
nand U1149 (N_1149,In_63,In_520);
nor U1150 (N_1150,In_629,In_1757);
nand U1151 (N_1151,In_879,In_1446);
or U1152 (N_1152,In_1778,In_1432);
nand U1153 (N_1153,In_367,In_101);
nor U1154 (N_1154,In_1346,In_572);
or U1155 (N_1155,In_1189,In_1717);
nand U1156 (N_1156,In_1161,In_1011);
nor U1157 (N_1157,In_1388,In_715);
or U1158 (N_1158,In_136,In_1557);
nand U1159 (N_1159,In_1728,In_4);
nand U1160 (N_1160,In_1853,In_142);
or U1161 (N_1161,In_1055,In_1125);
nand U1162 (N_1162,In_1252,In_1680);
or U1163 (N_1163,In_845,In_1578);
and U1164 (N_1164,In_1980,In_443);
or U1165 (N_1165,In_133,In_50);
or U1166 (N_1166,In_1941,In_1529);
and U1167 (N_1167,In_492,In_1117);
and U1168 (N_1168,In_1953,In_1243);
or U1169 (N_1169,In_850,In_62);
and U1170 (N_1170,In_403,In_142);
and U1171 (N_1171,In_546,In_833);
nand U1172 (N_1172,In_1621,In_405);
nand U1173 (N_1173,In_104,In_1707);
nor U1174 (N_1174,In_947,In_1492);
nor U1175 (N_1175,In_354,In_1703);
nor U1176 (N_1176,In_292,In_21);
nor U1177 (N_1177,In_425,In_52);
and U1178 (N_1178,In_352,In_1624);
or U1179 (N_1179,In_1006,In_1559);
nand U1180 (N_1180,In_1242,In_990);
nand U1181 (N_1181,In_1907,In_1362);
nand U1182 (N_1182,In_1288,In_166);
or U1183 (N_1183,In_999,In_1627);
nand U1184 (N_1184,In_1583,In_1302);
nand U1185 (N_1185,In_233,In_1913);
and U1186 (N_1186,In_1042,In_392);
nor U1187 (N_1187,In_1118,In_1810);
and U1188 (N_1188,In_138,In_522);
nand U1189 (N_1189,In_191,In_1919);
or U1190 (N_1190,In_1581,In_1400);
and U1191 (N_1191,In_1081,In_1420);
or U1192 (N_1192,In_1780,In_1721);
and U1193 (N_1193,In_1108,In_566);
nand U1194 (N_1194,In_1159,In_9);
or U1195 (N_1195,In_986,In_1225);
nand U1196 (N_1196,In_1616,In_1318);
or U1197 (N_1197,In_5,In_66);
and U1198 (N_1198,In_549,In_760);
nand U1199 (N_1199,In_1596,In_316);
nand U1200 (N_1200,In_1776,In_238);
or U1201 (N_1201,In_1815,In_788);
or U1202 (N_1202,In_728,In_1318);
nor U1203 (N_1203,In_1162,In_114);
nor U1204 (N_1204,In_301,In_829);
nor U1205 (N_1205,In_1583,In_1282);
or U1206 (N_1206,In_1731,In_303);
and U1207 (N_1207,In_735,In_625);
nor U1208 (N_1208,In_1062,In_843);
or U1209 (N_1209,In_1867,In_1833);
nand U1210 (N_1210,In_1504,In_782);
nor U1211 (N_1211,In_1830,In_1413);
and U1212 (N_1212,In_977,In_493);
or U1213 (N_1213,In_1392,In_829);
nor U1214 (N_1214,In_1120,In_411);
nor U1215 (N_1215,In_1011,In_497);
or U1216 (N_1216,In_26,In_537);
xnor U1217 (N_1217,In_827,In_408);
nand U1218 (N_1218,In_702,In_1809);
and U1219 (N_1219,In_1827,In_1431);
nand U1220 (N_1220,In_688,In_877);
or U1221 (N_1221,In_1585,In_1778);
nor U1222 (N_1222,In_1032,In_746);
or U1223 (N_1223,In_1444,In_276);
nor U1224 (N_1224,In_918,In_1033);
nor U1225 (N_1225,In_1137,In_228);
and U1226 (N_1226,In_718,In_81);
nand U1227 (N_1227,In_1868,In_1538);
and U1228 (N_1228,In_209,In_1205);
nor U1229 (N_1229,In_1526,In_1170);
nand U1230 (N_1230,In_993,In_265);
nand U1231 (N_1231,In_322,In_997);
and U1232 (N_1232,In_716,In_1441);
and U1233 (N_1233,In_482,In_377);
or U1234 (N_1234,In_725,In_1203);
and U1235 (N_1235,In_1329,In_1318);
nand U1236 (N_1236,In_1410,In_1247);
or U1237 (N_1237,In_993,In_1278);
nor U1238 (N_1238,In_226,In_1007);
nand U1239 (N_1239,In_482,In_933);
or U1240 (N_1240,In_1584,In_1875);
and U1241 (N_1241,In_1449,In_1840);
or U1242 (N_1242,In_1481,In_1326);
or U1243 (N_1243,In_813,In_96);
nor U1244 (N_1244,In_399,In_340);
or U1245 (N_1245,In_1195,In_966);
nand U1246 (N_1246,In_1885,In_1872);
and U1247 (N_1247,In_1216,In_1166);
and U1248 (N_1248,In_1118,In_83);
or U1249 (N_1249,In_1865,In_765);
nand U1250 (N_1250,In_844,In_698);
nand U1251 (N_1251,In_176,In_423);
and U1252 (N_1252,In_816,In_844);
and U1253 (N_1253,In_588,In_731);
or U1254 (N_1254,In_1216,In_15);
nor U1255 (N_1255,In_1600,In_1580);
nor U1256 (N_1256,In_817,In_1857);
nor U1257 (N_1257,In_931,In_1914);
nor U1258 (N_1258,In_549,In_732);
nor U1259 (N_1259,In_7,In_1631);
nand U1260 (N_1260,In_847,In_952);
and U1261 (N_1261,In_853,In_1244);
and U1262 (N_1262,In_1245,In_1265);
nor U1263 (N_1263,In_1266,In_1021);
nor U1264 (N_1264,In_603,In_1820);
nand U1265 (N_1265,In_103,In_1325);
nand U1266 (N_1266,In_205,In_436);
xnor U1267 (N_1267,In_761,In_463);
and U1268 (N_1268,In_112,In_692);
nor U1269 (N_1269,In_897,In_112);
and U1270 (N_1270,In_621,In_1019);
and U1271 (N_1271,In_628,In_816);
nand U1272 (N_1272,In_501,In_664);
and U1273 (N_1273,In_1246,In_1015);
and U1274 (N_1274,In_1785,In_948);
nor U1275 (N_1275,In_640,In_1839);
nor U1276 (N_1276,In_502,In_1522);
nor U1277 (N_1277,In_218,In_409);
nor U1278 (N_1278,In_1778,In_879);
nor U1279 (N_1279,In_1260,In_685);
or U1280 (N_1280,In_1513,In_844);
nor U1281 (N_1281,In_530,In_996);
nor U1282 (N_1282,In_1783,In_1520);
nor U1283 (N_1283,In_1815,In_768);
nand U1284 (N_1284,In_824,In_1978);
or U1285 (N_1285,In_580,In_255);
or U1286 (N_1286,In_798,In_96);
nor U1287 (N_1287,In_729,In_898);
or U1288 (N_1288,In_1224,In_495);
nand U1289 (N_1289,In_1567,In_831);
nor U1290 (N_1290,In_998,In_1235);
or U1291 (N_1291,In_462,In_313);
and U1292 (N_1292,In_955,In_1119);
nand U1293 (N_1293,In_1395,In_1404);
and U1294 (N_1294,In_1031,In_396);
nand U1295 (N_1295,In_895,In_1541);
nor U1296 (N_1296,In_909,In_340);
xnor U1297 (N_1297,In_1701,In_794);
or U1298 (N_1298,In_1017,In_1674);
nor U1299 (N_1299,In_1376,In_1735);
nor U1300 (N_1300,In_415,In_1506);
or U1301 (N_1301,In_771,In_1690);
and U1302 (N_1302,In_1520,In_217);
nand U1303 (N_1303,In_1481,In_584);
or U1304 (N_1304,In_1354,In_445);
and U1305 (N_1305,In_861,In_426);
and U1306 (N_1306,In_1480,In_497);
nor U1307 (N_1307,In_1065,In_210);
nand U1308 (N_1308,In_1188,In_630);
nand U1309 (N_1309,In_1178,In_405);
or U1310 (N_1310,In_897,In_1504);
nor U1311 (N_1311,In_1125,In_401);
nand U1312 (N_1312,In_229,In_1670);
and U1313 (N_1313,In_1010,In_1494);
nand U1314 (N_1314,In_790,In_1382);
nand U1315 (N_1315,In_401,In_927);
and U1316 (N_1316,In_1184,In_1790);
or U1317 (N_1317,In_1169,In_1129);
nor U1318 (N_1318,In_235,In_922);
or U1319 (N_1319,In_359,In_239);
and U1320 (N_1320,In_1753,In_151);
nor U1321 (N_1321,In_155,In_1099);
nor U1322 (N_1322,In_807,In_483);
or U1323 (N_1323,In_261,In_505);
nand U1324 (N_1324,In_1177,In_318);
nor U1325 (N_1325,In_1876,In_1371);
nor U1326 (N_1326,In_1070,In_409);
or U1327 (N_1327,In_1872,In_796);
or U1328 (N_1328,In_1689,In_1224);
nand U1329 (N_1329,In_1765,In_1101);
or U1330 (N_1330,In_1202,In_1656);
or U1331 (N_1331,In_540,In_289);
and U1332 (N_1332,In_1522,In_758);
and U1333 (N_1333,In_310,In_1151);
and U1334 (N_1334,In_1063,In_1540);
xor U1335 (N_1335,In_1925,In_1499);
and U1336 (N_1336,In_1527,In_1591);
nand U1337 (N_1337,In_1327,In_386);
nor U1338 (N_1338,In_1192,In_728);
or U1339 (N_1339,In_1272,In_1985);
or U1340 (N_1340,In_592,In_683);
nand U1341 (N_1341,In_1077,In_1344);
and U1342 (N_1342,In_1011,In_385);
nor U1343 (N_1343,In_1012,In_402);
or U1344 (N_1344,In_1008,In_1437);
nor U1345 (N_1345,In_1348,In_1931);
nor U1346 (N_1346,In_398,In_425);
nand U1347 (N_1347,In_1970,In_1848);
nor U1348 (N_1348,In_1329,In_616);
and U1349 (N_1349,In_972,In_1456);
nor U1350 (N_1350,In_846,In_1178);
nor U1351 (N_1351,In_1160,In_1697);
nor U1352 (N_1352,In_661,In_127);
nand U1353 (N_1353,In_1220,In_663);
nor U1354 (N_1354,In_744,In_615);
nand U1355 (N_1355,In_390,In_1655);
nand U1356 (N_1356,In_1630,In_751);
or U1357 (N_1357,In_619,In_1564);
and U1358 (N_1358,In_974,In_653);
or U1359 (N_1359,In_424,In_1924);
nand U1360 (N_1360,In_1230,In_41);
nand U1361 (N_1361,In_102,In_1533);
or U1362 (N_1362,In_472,In_767);
nand U1363 (N_1363,In_1822,In_557);
nor U1364 (N_1364,In_1084,In_827);
nor U1365 (N_1365,In_1256,In_750);
nor U1366 (N_1366,In_1151,In_971);
nor U1367 (N_1367,In_446,In_1602);
or U1368 (N_1368,In_875,In_1455);
and U1369 (N_1369,In_456,In_1427);
nand U1370 (N_1370,In_566,In_1254);
nor U1371 (N_1371,In_497,In_1611);
or U1372 (N_1372,In_297,In_696);
or U1373 (N_1373,In_230,In_388);
nor U1374 (N_1374,In_1282,In_969);
nand U1375 (N_1375,In_997,In_522);
nor U1376 (N_1376,In_262,In_643);
or U1377 (N_1377,In_1875,In_1897);
and U1378 (N_1378,In_88,In_1895);
nor U1379 (N_1379,In_1319,In_1508);
nor U1380 (N_1380,In_845,In_279);
or U1381 (N_1381,In_443,In_355);
nand U1382 (N_1382,In_1301,In_996);
nand U1383 (N_1383,In_1600,In_1953);
or U1384 (N_1384,In_1123,In_1071);
and U1385 (N_1385,In_1551,In_1547);
nor U1386 (N_1386,In_531,In_623);
nor U1387 (N_1387,In_1127,In_304);
or U1388 (N_1388,In_1212,In_772);
and U1389 (N_1389,In_1773,In_1423);
nor U1390 (N_1390,In_1902,In_1188);
and U1391 (N_1391,In_1003,In_334);
or U1392 (N_1392,In_1640,In_987);
and U1393 (N_1393,In_1904,In_533);
and U1394 (N_1394,In_1045,In_1176);
and U1395 (N_1395,In_1619,In_1360);
and U1396 (N_1396,In_1819,In_577);
nor U1397 (N_1397,In_1502,In_1802);
or U1398 (N_1398,In_392,In_291);
nand U1399 (N_1399,In_564,In_135);
and U1400 (N_1400,In_1323,In_1320);
xnor U1401 (N_1401,In_1100,In_1998);
or U1402 (N_1402,In_515,In_1158);
or U1403 (N_1403,In_637,In_823);
nor U1404 (N_1404,In_1123,In_586);
or U1405 (N_1405,In_1043,In_549);
or U1406 (N_1406,In_435,In_1875);
and U1407 (N_1407,In_387,In_59);
and U1408 (N_1408,In_1579,In_1908);
and U1409 (N_1409,In_410,In_1476);
and U1410 (N_1410,In_250,In_1072);
xor U1411 (N_1411,In_863,In_377);
and U1412 (N_1412,In_1436,In_985);
nor U1413 (N_1413,In_796,In_292);
and U1414 (N_1414,In_727,In_1388);
or U1415 (N_1415,In_1137,In_1470);
or U1416 (N_1416,In_1780,In_364);
nor U1417 (N_1417,In_650,In_1613);
and U1418 (N_1418,In_1436,In_63);
nand U1419 (N_1419,In_914,In_1509);
or U1420 (N_1420,In_1643,In_1731);
and U1421 (N_1421,In_1638,In_1032);
nand U1422 (N_1422,In_590,In_1713);
nor U1423 (N_1423,In_843,In_1402);
nand U1424 (N_1424,In_816,In_376);
or U1425 (N_1425,In_1258,In_940);
nor U1426 (N_1426,In_1594,In_481);
and U1427 (N_1427,In_673,In_1430);
and U1428 (N_1428,In_1856,In_1667);
nand U1429 (N_1429,In_742,In_498);
nor U1430 (N_1430,In_1727,In_457);
or U1431 (N_1431,In_1568,In_807);
nor U1432 (N_1432,In_1665,In_987);
or U1433 (N_1433,In_1515,In_394);
nand U1434 (N_1434,In_864,In_1904);
nor U1435 (N_1435,In_112,In_10);
nand U1436 (N_1436,In_1104,In_1699);
nor U1437 (N_1437,In_813,In_1131);
and U1438 (N_1438,In_1603,In_693);
and U1439 (N_1439,In_1749,In_1677);
nor U1440 (N_1440,In_73,In_245);
and U1441 (N_1441,In_1415,In_593);
or U1442 (N_1442,In_1406,In_821);
nand U1443 (N_1443,In_1201,In_3);
and U1444 (N_1444,In_762,In_615);
or U1445 (N_1445,In_482,In_239);
or U1446 (N_1446,In_1345,In_977);
nor U1447 (N_1447,In_1426,In_417);
nor U1448 (N_1448,In_678,In_267);
and U1449 (N_1449,In_732,In_1351);
and U1450 (N_1450,In_1762,In_511);
nand U1451 (N_1451,In_1864,In_1970);
nor U1452 (N_1452,In_565,In_775);
nor U1453 (N_1453,In_948,In_1034);
nand U1454 (N_1454,In_67,In_398);
or U1455 (N_1455,In_1725,In_859);
or U1456 (N_1456,In_431,In_805);
or U1457 (N_1457,In_467,In_1844);
nor U1458 (N_1458,In_518,In_1377);
or U1459 (N_1459,In_300,In_951);
or U1460 (N_1460,In_681,In_295);
nor U1461 (N_1461,In_1880,In_1007);
nand U1462 (N_1462,In_1071,In_1282);
and U1463 (N_1463,In_1177,In_1229);
and U1464 (N_1464,In_425,In_915);
or U1465 (N_1465,In_975,In_663);
nand U1466 (N_1466,In_616,In_1252);
nand U1467 (N_1467,In_1137,In_1602);
nor U1468 (N_1468,In_112,In_1635);
or U1469 (N_1469,In_1648,In_219);
nand U1470 (N_1470,In_1359,In_935);
or U1471 (N_1471,In_921,In_343);
nor U1472 (N_1472,In_809,In_253);
or U1473 (N_1473,In_1785,In_830);
and U1474 (N_1474,In_1559,In_1416);
nand U1475 (N_1475,In_1186,In_1856);
nor U1476 (N_1476,In_88,In_1258);
nor U1477 (N_1477,In_742,In_1874);
and U1478 (N_1478,In_68,In_1617);
and U1479 (N_1479,In_1373,In_1189);
nand U1480 (N_1480,In_727,In_910);
and U1481 (N_1481,In_950,In_836);
and U1482 (N_1482,In_1440,In_383);
nand U1483 (N_1483,In_1520,In_1856);
or U1484 (N_1484,In_520,In_635);
and U1485 (N_1485,In_208,In_1730);
nand U1486 (N_1486,In_943,In_494);
and U1487 (N_1487,In_137,In_1383);
or U1488 (N_1488,In_811,In_476);
and U1489 (N_1489,In_1085,In_1459);
and U1490 (N_1490,In_1750,In_1947);
nand U1491 (N_1491,In_890,In_656);
nand U1492 (N_1492,In_1592,In_997);
nand U1493 (N_1493,In_541,In_1308);
or U1494 (N_1494,In_295,In_1027);
nor U1495 (N_1495,In_190,In_1170);
and U1496 (N_1496,In_1925,In_153);
nor U1497 (N_1497,In_100,In_1315);
or U1498 (N_1498,In_1251,In_1257);
nand U1499 (N_1499,In_1051,In_1699);
nor U1500 (N_1500,In_203,In_1092);
nand U1501 (N_1501,In_21,In_780);
and U1502 (N_1502,In_1295,In_311);
or U1503 (N_1503,In_1707,In_1588);
and U1504 (N_1504,In_972,In_1714);
nand U1505 (N_1505,In_1938,In_1289);
nor U1506 (N_1506,In_686,In_1944);
and U1507 (N_1507,In_63,In_794);
and U1508 (N_1508,In_819,In_1361);
and U1509 (N_1509,In_1248,In_446);
and U1510 (N_1510,In_1395,In_1958);
and U1511 (N_1511,In_881,In_851);
and U1512 (N_1512,In_1919,In_38);
or U1513 (N_1513,In_760,In_1687);
nor U1514 (N_1514,In_66,In_762);
nand U1515 (N_1515,In_987,In_767);
or U1516 (N_1516,In_1423,In_430);
nor U1517 (N_1517,In_1145,In_1616);
nand U1518 (N_1518,In_780,In_1954);
nand U1519 (N_1519,In_299,In_735);
and U1520 (N_1520,In_458,In_1028);
or U1521 (N_1521,In_91,In_245);
and U1522 (N_1522,In_491,In_1084);
nand U1523 (N_1523,In_790,In_1433);
and U1524 (N_1524,In_663,In_531);
or U1525 (N_1525,In_212,In_55);
or U1526 (N_1526,In_668,In_549);
nor U1527 (N_1527,In_1121,In_406);
or U1528 (N_1528,In_1114,In_1977);
nor U1529 (N_1529,In_1286,In_588);
nand U1530 (N_1530,In_1857,In_1803);
nor U1531 (N_1531,In_1077,In_1563);
or U1532 (N_1532,In_1898,In_1466);
nand U1533 (N_1533,In_1230,In_1440);
nand U1534 (N_1534,In_834,In_357);
nand U1535 (N_1535,In_1084,In_1963);
nor U1536 (N_1536,In_1007,In_1782);
nand U1537 (N_1537,In_313,In_1009);
nor U1538 (N_1538,In_1607,In_1198);
or U1539 (N_1539,In_410,In_1522);
nor U1540 (N_1540,In_1058,In_1932);
or U1541 (N_1541,In_1014,In_873);
nor U1542 (N_1542,In_377,In_1194);
or U1543 (N_1543,In_1402,In_1493);
and U1544 (N_1544,In_1793,In_1156);
and U1545 (N_1545,In_1101,In_1095);
nor U1546 (N_1546,In_711,In_148);
or U1547 (N_1547,In_1775,In_1718);
and U1548 (N_1548,In_1894,In_1356);
nand U1549 (N_1549,In_1846,In_1046);
and U1550 (N_1550,In_1895,In_1884);
and U1551 (N_1551,In_579,In_197);
and U1552 (N_1552,In_23,In_1153);
or U1553 (N_1553,In_1685,In_284);
or U1554 (N_1554,In_1370,In_787);
and U1555 (N_1555,In_1290,In_863);
nor U1556 (N_1556,In_1848,In_1350);
nor U1557 (N_1557,In_516,In_659);
nor U1558 (N_1558,In_1689,In_1472);
xnor U1559 (N_1559,In_1298,In_515);
nand U1560 (N_1560,In_1778,In_876);
nor U1561 (N_1561,In_1173,In_1752);
or U1562 (N_1562,In_1559,In_931);
nor U1563 (N_1563,In_480,In_1213);
and U1564 (N_1564,In_1840,In_572);
nor U1565 (N_1565,In_1688,In_191);
nand U1566 (N_1566,In_304,In_1270);
and U1567 (N_1567,In_1841,In_1321);
nand U1568 (N_1568,In_1575,In_1713);
or U1569 (N_1569,In_737,In_832);
nand U1570 (N_1570,In_1872,In_602);
nor U1571 (N_1571,In_469,In_756);
nand U1572 (N_1572,In_1124,In_36);
nand U1573 (N_1573,In_1316,In_1611);
or U1574 (N_1574,In_192,In_498);
nand U1575 (N_1575,In_1206,In_190);
nor U1576 (N_1576,In_499,In_1290);
nor U1577 (N_1577,In_1773,In_558);
or U1578 (N_1578,In_985,In_1340);
and U1579 (N_1579,In_1553,In_1302);
and U1580 (N_1580,In_1208,In_289);
nand U1581 (N_1581,In_1835,In_216);
and U1582 (N_1582,In_1531,In_1483);
nor U1583 (N_1583,In_649,In_205);
nand U1584 (N_1584,In_1396,In_1029);
or U1585 (N_1585,In_1941,In_718);
nor U1586 (N_1586,In_1411,In_238);
and U1587 (N_1587,In_1928,In_1454);
nand U1588 (N_1588,In_667,In_71);
or U1589 (N_1589,In_1676,In_63);
or U1590 (N_1590,In_296,In_1961);
nor U1591 (N_1591,In_1955,In_673);
nor U1592 (N_1592,In_1305,In_1872);
or U1593 (N_1593,In_658,In_50);
nand U1594 (N_1594,In_1976,In_1526);
and U1595 (N_1595,In_506,In_1446);
and U1596 (N_1596,In_409,In_1533);
xor U1597 (N_1597,In_669,In_1843);
nand U1598 (N_1598,In_1072,In_29);
nand U1599 (N_1599,In_1831,In_886);
nand U1600 (N_1600,In_419,In_224);
and U1601 (N_1601,In_1394,In_1484);
and U1602 (N_1602,In_621,In_87);
or U1603 (N_1603,In_258,In_1389);
and U1604 (N_1604,In_1320,In_667);
and U1605 (N_1605,In_533,In_1170);
nand U1606 (N_1606,In_888,In_1980);
or U1607 (N_1607,In_697,In_102);
nand U1608 (N_1608,In_511,In_425);
and U1609 (N_1609,In_709,In_895);
nand U1610 (N_1610,In_324,In_1431);
nand U1611 (N_1611,In_1173,In_49);
nor U1612 (N_1612,In_924,In_1872);
xor U1613 (N_1613,In_1183,In_1485);
or U1614 (N_1614,In_1593,In_303);
nand U1615 (N_1615,In_725,In_46);
or U1616 (N_1616,In_1367,In_550);
nand U1617 (N_1617,In_971,In_584);
and U1618 (N_1618,In_55,In_1637);
and U1619 (N_1619,In_1086,In_1115);
nor U1620 (N_1620,In_974,In_1486);
and U1621 (N_1621,In_965,In_500);
and U1622 (N_1622,In_366,In_1676);
nand U1623 (N_1623,In_1436,In_73);
nor U1624 (N_1624,In_1826,In_1286);
or U1625 (N_1625,In_1214,In_453);
and U1626 (N_1626,In_762,In_660);
or U1627 (N_1627,In_1683,In_1611);
nand U1628 (N_1628,In_1157,In_1380);
nand U1629 (N_1629,In_758,In_1288);
or U1630 (N_1630,In_730,In_440);
or U1631 (N_1631,In_236,In_1954);
nand U1632 (N_1632,In_1485,In_158);
nand U1633 (N_1633,In_340,In_1657);
or U1634 (N_1634,In_1066,In_161);
and U1635 (N_1635,In_622,In_244);
or U1636 (N_1636,In_1650,In_1996);
or U1637 (N_1637,In_280,In_46);
or U1638 (N_1638,In_625,In_336);
nand U1639 (N_1639,In_1365,In_576);
nand U1640 (N_1640,In_954,In_787);
or U1641 (N_1641,In_291,In_718);
or U1642 (N_1642,In_1655,In_1188);
and U1643 (N_1643,In_539,In_261);
and U1644 (N_1644,In_4,In_1561);
nor U1645 (N_1645,In_326,In_710);
nor U1646 (N_1646,In_1789,In_1754);
nand U1647 (N_1647,In_660,In_1205);
nand U1648 (N_1648,In_300,In_638);
nor U1649 (N_1649,In_954,In_535);
nand U1650 (N_1650,In_1544,In_1674);
or U1651 (N_1651,In_93,In_1419);
nor U1652 (N_1652,In_1011,In_754);
and U1653 (N_1653,In_715,In_120);
nor U1654 (N_1654,In_86,In_1522);
nor U1655 (N_1655,In_186,In_901);
or U1656 (N_1656,In_1789,In_1792);
and U1657 (N_1657,In_166,In_1077);
or U1658 (N_1658,In_1197,In_25);
nor U1659 (N_1659,In_1814,In_818);
and U1660 (N_1660,In_736,In_1371);
nand U1661 (N_1661,In_355,In_554);
nor U1662 (N_1662,In_1306,In_1595);
and U1663 (N_1663,In_1001,In_183);
or U1664 (N_1664,In_1653,In_470);
nor U1665 (N_1665,In_1889,In_1840);
or U1666 (N_1666,In_734,In_600);
and U1667 (N_1667,In_185,In_594);
nand U1668 (N_1668,In_408,In_1675);
and U1669 (N_1669,In_253,In_757);
or U1670 (N_1670,In_1207,In_324);
or U1671 (N_1671,In_39,In_993);
or U1672 (N_1672,In_534,In_329);
nand U1673 (N_1673,In_1530,In_1914);
nor U1674 (N_1674,In_52,In_565);
or U1675 (N_1675,In_308,In_87);
nand U1676 (N_1676,In_623,In_1434);
nor U1677 (N_1677,In_27,In_1381);
nand U1678 (N_1678,In_1568,In_496);
and U1679 (N_1679,In_763,In_403);
and U1680 (N_1680,In_1843,In_1924);
nand U1681 (N_1681,In_1401,In_1612);
nor U1682 (N_1682,In_1744,In_1833);
nor U1683 (N_1683,In_1781,In_1791);
nor U1684 (N_1684,In_872,In_1872);
and U1685 (N_1685,In_475,In_1557);
or U1686 (N_1686,In_1410,In_494);
and U1687 (N_1687,In_763,In_1870);
or U1688 (N_1688,In_1947,In_32);
nor U1689 (N_1689,In_1954,In_549);
and U1690 (N_1690,In_841,In_639);
nand U1691 (N_1691,In_1496,In_1519);
nand U1692 (N_1692,In_911,In_91);
or U1693 (N_1693,In_1381,In_67);
nand U1694 (N_1694,In_415,In_1044);
or U1695 (N_1695,In_1084,In_884);
and U1696 (N_1696,In_913,In_845);
or U1697 (N_1697,In_1236,In_86);
nand U1698 (N_1698,In_773,In_1610);
and U1699 (N_1699,In_144,In_743);
nand U1700 (N_1700,In_1085,In_511);
or U1701 (N_1701,In_1175,In_892);
and U1702 (N_1702,In_724,In_1665);
nor U1703 (N_1703,In_1515,In_576);
nand U1704 (N_1704,In_43,In_1585);
nand U1705 (N_1705,In_549,In_1872);
nor U1706 (N_1706,In_800,In_110);
nor U1707 (N_1707,In_1218,In_1535);
nand U1708 (N_1708,In_548,In_13);
and U1709 (N_1709,In_746,In_1102);
nor U1710 (N_1710,In_104,In_1959);
and U1711 (N_1711,In_844,In_514);
and U1712 (N_1712,In_926,In_1320);
nand U1713 (N_1713,In_944,In_570);
and U1714 (N_1714,In_179,In_923);
nor U1715 (N_1715,In_487,In_1992);
nor U1716 (N_1716,In_356,In_730);
nand U1717 (N_1717,In_1885,In_1916);
nor U1718 (N_1718,In_1391,In_456);
and U1719 (N_1719,In_85,In_628);
nor U1720 (N_1720,In_1878,In_17);
nor U1721 (N_1721,In_448,In_58);
or U1722 (N_1722,In_1545,In_1112);
nor U1723 (N_1723,In_1216,In_914);
or U1724 (N_1724,In_628,In_676);
nor U1725 (N_1725,In_377,In_151);
or U1726 (N_1726,In_1841,In_394);
and U1727 (N_1727,In_298,In_278);
nand U1728 (N_1728,In_542,In_1680);
nand U1729 (N_1729,In_663,In_1223);
and U1730 (N_1730,In_301,In_266);
or U1731 (N_1731,In_1687,In_758);
and U1732 (N_1732,In_1686,In_1062);
nand U1733 (N_1733,In_963,In_612);
or U1734 (N_1734,In_1284,In_632);
nor U1735 (N_1735,In_941,In_1390);
and U1736 (N_1736,In_729,In_605);
or U1737 (N_1737,In_503,In_1602);
or U1738 (N_1738,In_1408,In_1732);
and U1739 (N_1739,In_396,In_1053);
nor U1740 (N_1740,In_1331,In_1923);
and U1741 (N_1741,In_376,In_1445);
or U1742 (N_1742,In_77,In_957);
nor U1743 (N_1743,In_968,In_1579);
nand U1744 (N_1744,In_1415,In_1692);
nor U1745 (N_1745,In_361,In_585);
nand U1746 (N_1746,In_998,In_410);
and U1747 (N_1747,In_1357,In_677);
nand U1748 (N_1748,In_384,In_1255);
nor U1749 (N_1749,In_961,In_1834);
or U1750 (N_1750,In_1934,In_363);
nand U1751 (N_1751,In_985,In_1424);
or U1752 (N_1752,In_1804,In_1024);
nand U1753 (N_1753,In_1287,In_669);
and U1754 (N_1754,In_1020,In_1351);
and U1755 (N_1755,In_417,In_568);
or U1756 (N_1756,In_1645,In_1850);
or U1757 (N_1757,In_946,In_52);
and U1758 (N_1758,In_353,In_1647);
or U1759 (N_1759,In_963,In_449);
nor U1760 (N_1760,In_804,In_778);
xnor U1761 (N_1761,In_147,In_151);
nor U1762 (N_1762,In_11,In_770);
xnor U1763 (N_1763,In_569,In_1988);
nor U1764 (N_1764,In_1298,In_115);
or U1765 (N_1765,In_62,In_517);
and U1766 (N_1766,In_571,In_655);
nand U1767 (N_1767,In_499,In_726);
or U1768 (N_1768,In_1510,In_405);
and U1769 (N_1769,In_1642,In_956);
nor U1770 (N_1770,In_1676,In_1741);
and U1771 (N_1771,In_1774,In_1633);
nand U1772 (N_1772,In_524,In_91);
nand U1773 (N_1773,In_71,In_895);
nor U1774 (N_1774,In_91,In_1755);
or U1775 (N_1775,In_303,In_1566);
and U1776 (N_1776,In_1472,In_183);
xnor U1777 (N_1777,In_848,In_223);
and U1778 (N_1778,In_276,In_85);
nand U1779 (N_1779,In_302,In_1711);
nor U1780 (N_1780,In_329,In_936);
or U1781 (N_1781,In_840,In_764);
nor U1782 (N_1782,In_274,In_1579);
and U1783 (N_1783,In_1889,In_1693);
nand U1784 (N_1784,In_126,In_637);
nor U1785 (N_1785,In_1360,In_599);
and U1786 (N_1786,In_1161,In_954);
nand U1787 (N_1787,In_1188,In_1373);
and U1788 (N_1788,In_952,In_617);
nand U1789 (N_1789,In_1278,In_807);
nand U1790 (N_1790,In_1836,In_776);
nand U1791 (N_1791,In_1235,In_1435);
or U1792 (N_1792,In_786,In_1320);
and U1793 (N_1793,In_998,In_618);
or U1794 (N_1794,In_14,In_1251);
nor U1795 (N_1795,In_1386,In_979);
nand U1796 (N_1796,In_1760,In_1675);
nor U1797 (N_1797,In_231,In_791);
nand U1798 (N_1798,In_1566,In_953);
nor U1799 (N_1799,In_1800,In_432);
nand U1800 (N_1800,In_249,In_261);
nor U1801 (N_1801,In_1650,In_134);
nor U1802 (N_1802,In_2,In_1530);
and U1803 (N_1803,In_1297,In_1737);
and U1804 (N_1804,In_1133,In_809);
or U1805 (N_1805,In_469,In_1649);
nor U1806 (N_1806,In_968,In_1478);
nor U1807 (N_1807,In_934,In_1372);
and U1808 (N_1808,In_1990,In_654);
nor U1809 (N_1809,In_1021,In_214);
or U1810 (N_1810,In_1786,In_148);
and U1811 (N_1811,In_1665,In_752);
nor U1812 (N_1812,In_1022,In_1020);
or U1813 (N_1813,In_1087,In_479);
nor U1814 (N_1814,In_1362,In_1682);
and U1815 (N_1815,In_1416,In_1972);
nor U1816 (N_1816,In_134,In_1154);
or U1817 (N_1817,In_86,In_1224);
and U1818 (N_1818,In_932,In_475);
nand U1819 (N_1819,In_602,In_152);
and U1820 (N_1820,In_809,In_1888);
nand U1821 (N_1821,In_429,In_109);
nand U1822 (N_1822,In_1917,In_173);
nand U1823 (N_1823,In_423,In_1726);
nand U1824 (N_1824,In_838,In_1336);
nor U1825 (N_1825,In_1267,In_852);
nand U1826 (N_1826,In_995,In_1975);
nand U1827 (N_1827,In_105,In_1285);
nand U1828 (N_1828,In_712,In_1957);
nor U1829 (N_1829,In_1309,In_1907);
nand U1830 (N_1830,In_354,In_1044);
nand U1831 (N_1831,In_7,In_1445);
nand U1832 (N_1832,In_963,In_652);
or U1833 (N_1833,In_1203,In_728);
and U1834 (N_1834,In_1770,In_304);
and U1835 (N_1835,In_1626,In_1789);
and U1836 (N_1836,In_1268,In_1862);
and U1837 (N_1837,In_717,In_1909);
nor U1838 (N_1838,In_61,In_1822);
nor U1839 (N_1839,In_1238,In_855);
nor U1840 (N_1840,In_443,In_1979);
nand U1841 (N_1841,In_1230,In_892);
nor U1842 (N_1842,In_557,In_1427);
and U1843 (N_1843,In_337,In_1131);
nand U1844 (N_1844,In_497,In_183);
or U1845 (N_1845,In_867,In_555);
or U1846 (N_1846,In_1374,In_1827);
and U1847 (N_1847,In_1777,In_379);
nor U1848 (N_1848,In_1637,In_1552);
nor U1849 (N_1849,In_764,In_1249);
nand U1850 (N_1850,In_1660,In_1759);
nand U1851 (N_1851,In_881,In_118);
and U1852 (N_1852,In_231,In_1693);
or U1853 (N_1853,In_58,In_761);
nor U1854 (N_1854,In_223,In_1345);
nor U1855 (N_1855,In_1250,In_13);
and U1856 (N_1856,In_1112,In_607);
and U1857 (N_1857,In_1248,In_697);
or U1858 (N_1858,In_592,In_1317);
nor U1859 (N_1859,In_851,In_848);
nand U1860 (N_1860,In_847,In_720);
and U1861 (N_1861,In_402,In_459);
or U1862 (N_1862,In_24,In_4);
nor U1863 (N_1863,In_1136,In_675);
or U1864 (N_1864,In_94,In_164);
nand U1865 (N_1865,In_1143,In_60);
and U1866 (N_1866,In_952,In_48);
and U1867 (N_1867,In_1447,In_153);
or U1868 (N_1868,In_435,In_433);
nand U1869 (N_1869,In_1157,In_1065);
xor U1870 (N_1870,In_1588,In_1542);
nand U1871 (N_1871,In_776,In_1333);
or U1872 (N_1872,In_1383,In_210);
or U1873 (N_1873,In_455,In_743);
nand U1874 (N_1874,In_169,In_677);
and U1875 (N_1875,In_286,In_1641);
nor U1876 (N_1876,In_1644,In_370);
and U1877 (N_1877,In_174,In_1022);
nor U1878 (N_1878,In_16,In_1868);
or U1879 (N_1879,In_531,In_1036);
and U1880 (N_1880,In_310,In_1192);
nor U1881 (N_1881,In_1958,In_655);
nand U1882 (N_1882,In_1392,In_1322);
or U1883 (N_1883,In_1253,In_916);
nor U1884 (N_1884,In_344,In_614);
or U1885 (N_1885,In_1024,In_1595);
nor U1886 (N_1886,In_757,In_1836);
nor U1887 (N_1887,In_550,In_898);
nor U1888 (N_1888,In_164,In_417);
nand U1889 (N_1889,In_1877,In_1215);
or U1890 (N_1890,In_1387,In_1557);
nor U1891 (N_1891,In_1643,In_1156);
or U1892 (N_1892,In_271,In_1426);
and U1893 (N_1893,In_1209,In_644);
or U1894 (N_1894,In_1926,In_674);
and U1895 (N_1895,In_143,In_770);
nor U1896 (N_1896,In_647,In_909);
nand U1897 (N_1897,In_27,In_1010);
and U1898 (N_1898,In_842,In_425);
nor U1899 (N_1899,In_1524,In_41);
and U1900 (N_1900,In_1259,In_665);
nor U1901 (N_1901,In_361,In_1622);
nand U1902 (N_1902,In_1117,In_322);
and U1903 (N_1903,In_827,In_1695);
and U1904 (N_1904,In_1972,In_1714);
nor U1905 (N_1905,In_1530,In_700);
or U1906 (N_1906,In_1270,In_1807);
nor U1907 (N_1907,In_1973,In_1793);
nor U1908 (N_1908,In_735,In_1784);
nor U1909 (N_1909,In_531,In_1897);
or U1910 (N_1910,In_1522,In_243);
and U1911 (N_1911,In_966,In_1406);
nor U1912 (N_1912,In_84,In_331);
nor U1913 (N_1913,In_899,In_1281);
and U1914 (N_1914,In_548,In_1458);
nand U1915 (N_1915,In_732,In_866);
nor U1916 (N_1916,In_963,In_337);
nand U1917 (N_1917,In_1065,In_1591);
nand U1918 (N_1918,In_558,In_1262);
nor U1919 (N_1919,In_209,In_1654);
nor U1920 (N_1920,In_826,In_1749);
or U1921 (N_1921,In_1546,In_294);
nand U1922 (N_1922,In_1100,In_553);
nand U1923 (N_1923,In_401,In_1163);
nor U1924 (N_1924,In_277,In_1676);
or U1925 (N_1925,In_226,In_948);
and U1926 (N_1926,In_575,In_40);
nand U1927 (N_1927,In_2,In_1651);
or U1928 (N_1928,In_1876,In_1879);
or U1929 (N_1929,In_1849,In_668);
or U1930 (N_1930,In_1441,In_1718);
or U1931 (N_1931,In_205,In_1670);
nor U1932 (N_1932,In_56,In_1118);
and U1933 (N_1933,In_813,In_645);
nor U1934 (N_1934,In_340,In_90);
and U1935 (N_1935,In_751,In_1351);
nor U1936 (N_1936,In_1751,In_723);
nor U1937 (N_1937,In_1668,In_531);
nor U1938 (N_1938,In_1796,In_453);
and U1939 (N_1939,In_824,In_417);
nor U1940 (N_1940,In_557,In_1686);
nand U1941 (N_1941,In_361,In_1255);
nor U1942 (N_1942,In_778,In_484);
or U1943 (N_1943,In_1514,In_1368);
and U1944 (N_1944,In_1205,In_1093);
and U1945 (N_1945,In_1450,In_1912);
nand U1946 (N_1946,In_594,In_155);
and U1947 (N_1947,In_1224,In_1913);
nor U1948 (N_1948,In_1831,In_1971);
and U1949 (N_1949,In_621,In_107);
nand U1950 (N_1950,In_1691,In_1069);
nand U1951 (N_1951,In_1216,In_1429);
nand U1952 (N_1952,In_1544,In_1494);
nand U1953 (N_1953,In_1741,In_271);
and U1954 (N_1954,In_1832,In_1677);
or U1955 (N_1955,In_92,In_1952);
or U1956 (N_1956,In_591,In_331);
nand U1957 (N_1957,In_691,In_339);
and U1958 (N_1958,In_906,In_248);
nor U1959 (N_1959,In_802,In_1698);
and U1960 (N_1960,In_1521,In_1087);
or U1961 (N_1961,In_1400,In_359);
nor U1962 (N_1962,In_1935,In_1749);
and U1963 (N_1963,In_1806,In_1053);
nand U1964 (N_1964,In_288,In_1990);
nand U1965 (N_1965,In_81,In_1254);
nor U1966 (N_1966,In_1796,In_369);
and U1967 (N_1967,In_781,In_331);
nor U1968 (N_1968,In_1679,In_1874);
and U1969 (N_1969,In_455,In_16);
nor U1970 (N_1970,In_1424,In_712);
or U1971 (N_1971,In_180,In_862);
nand U1972 (N_1972,In_116,In_35);
nor U1973 (N_1973,In_1057,In_1511);
nand U1974 (N_1974,In_1887,In_944);
nor U1975 (N_1975,In_341,In_554);
or U1976 (N_1976,In_413,In_401);
nand U1977 (N_1977,In_220,In_714);
nor U1978 (N_1978,In_708,In_11);
and U1979 (N_1979,In_998,In_1925);
and U1980 (N_1980,In_1650,In_1890);
nand U1981 (N_1981,In_734,In_585);
nor U1982 (N_1982,In_1562,In_732);
nor U1983 (N_1983,In_1745,In_1651);
or U1984 (N_1984,In_922,In_1226);
or U1985 (N_1985,In_901,In_801);
nor U1986 (N_1986,In_1746,In_555);
or U1987 (N_1987,In_923,In_1446);
and U1988 (N_1988,In_639,In_679);
and U1989 (N_1989,In_118,In_1684);
or U1990 (N_1990,In_946,In_218);
or U1991 (N_1991,In_290,In_285);
nor U1992 (N_1992,In_396,In_181);
and U1993 (N_1993,In_1982,In_357);
or U1994 (N_1994,In_774,In_683);
nor U1995 (N_1995,In_11,In_1656);
nand U1996 (N_1996,In_1346,In_1646);
nor U1997 (N_1997,In_1151,In_1005);
and U1998 (N_1998,In_1935,In_1561);
or U1999 (N_1999,In_323,In_585);
nor U2000 (N_2000,In_278,In_45);
and U2001 (N_2001,In_1973,In_1604);
and U2002 (N_2002,In_971,In_1595);
and U2003 (N_2003,In_515,In_365);
nand U2004 (N_2004,In_198,In_971);
and U2005 (N_2005,In_232,In_913);
nand U2006 (N_2006,In_1026,In_1044);
nand U2007 (N_2007,In_1781,In_1006);
nor U2008 (N_2008,In_1868,In_1128);
nor U2009 (N_2009,In_1662,In_1354);
or U2010 (N_2010,In_1229,In_1593);
and U2011 (N_2011,In_1818,In_1707);
nand U2012 (N_2012,In_1182,In_214);
and U2013 (N_2013,In_1802,In_1275);
nor U2014 (N_2014,In_1442,In_1054);
nand U2015 (N_2015,In_324,In_1290);
nor U2016 (N_2016,In_941,In_981);
or U2017 (N_2017,In_1555,In_252);
or U2018 (N_2018,In_338,In_24);
or U2019 (N_2019,In_1749,In_1189);
nand U2020 (N_2020,In_1844,In_175);
nand U2021 (N_2021,In_1150,In_1725);
nor U2022 (N_2022,In_735,In_823);
nor U2023 (N_2023,In_703,In_691);
nand U2024 (N_2024,In_1772,In_1204);
or U2025 (N_2025,In_547,In_405);
or U2026 (N_2026,In_639,In_433);
nand U2027 (N_2027,In_350,In_289);
or U2028 (N_2028,In_1682,In_1164);
or U2029 (N_2029,In_642,In_937);
or U2030 (N_2030,In_1219,In_1832);
and U2031 (N_2031,In_103,In_315);
nor U2032 (N_2032,In_1313,In_1509);
or U2033 (N_2033,In_1573,In_100);
or U2034 (N_2034,In_938,In_393);
and U2035 (N_2035,In_560,In_1589);
nand U2036 (N_2036,In_235,In_1154);
nor U2037 (N_2037,In_335,In_1637);
nor U2038 (N_2038,In_841,In_192);
nor U2039 (N_2039,In_548,In_1152);
nand U2040 (N_2040,In_1907,In_720);
nand U2041 (N_2041,In_210,In_373);
or U2042 (N_2042,In_455,In_1315);
nor U2043 (N_2043,In_1892,In_1624);
nand U2044 (N_2044,In_1683,In_1754);
nand U2045 (N_2045,In_1493,In_1338);
nor U2046 (N_2046,In_64,In_478);
or U2047 (N_2047,In_90,In_785);
nand U2048 (N_2048,In_1389,In_1984);
and U2049 (N_2049,In_456,In_1850);
nand U2050 (N_2050,In_1352,In_910);
nor U2051 (N_2051,In_593,In_1348);
or U2052 (N_2052,In_1401,In_354);
nor U2053 (N_2053,In_1056,In_1743);
and U2054 (N_2054,In_1924,In_344);
and U2055 (N_2055,In_770,In_1669);
and U2056 (N_2056,In_853,In_916);
and U2057 (N_2057,In_1447,In_184);
or U2058 (N_2058,In_1043,In_1488);
nor U2059 (N_2059,In_1895,In_454);
and U2060 (N_2060,In_778,In_1150);
and U2061 (N_2061,In_694,In_1892);
and U2062 (N_2062,In_1530,In_209);
or U2063 (N_2063,In_817,In_235);
nor U2064 (N_2064,In_1903,In_1617);
and U2065 (N_2065,In_838,In_679);
nor U2066 (N_2066,In_1904,In_1410);
nand U2067 (N_2067,In_427,In_822);
nand U2068 (N_2068,In_583,In_894);
or U2069 (N_2069,In_15,In_1556);
nand U2070 (N_2070,In_889,In_1798);
nor U2071 (N_2071,In_1123,In_1244);
nand U2072 (N_2072,In_1217,In_1847);
nand U2073 (N_2073,In_669,In_638);
and U2074 (N_2074,In_1761,In_1647);
or U2075 (N_2075,In_762,In_502);
or U2076 (N_2076,In_793,In_481);
or U2077 (N_2077,In_1551,In_1727);
nor U2078 (N_2078,In_177,In_713);
nor U2079 (N_2079,In_1256,In_434);
and U2080 (N_2080,In_632,In_851);
and U2081 (N_2081,In_1039,In_379);
nor U2082 (N_2082,In_229,In_38);
nand U2083 (N_2083,In_1034,In_1476);
and U2084 (N_2084,In_302,In_1360);
nor U2085 (N_2085,In_117,In_1206);
nor U2086 (N_2086,In_1866,In_1839);
nor U2087 (N_2087,In_1885,In_812);
and U2088 (N_2088,In_1355,In_687);
nor U2089 (N_2089,In_1604,In_1702);
nor U2090 (N_2090,In_197,In_508);
nor U2091 (N_2091,In_1950,In_1819);
nand U2092 (N_2092,In_234,In_1906);
and U2093 (N_2093,In_536,In_230);
nand U2094 (N_2094,In_729,In_1320);
or U2095 (N_2095,In_693,In_813);
nor U2096 (N_2096,In_1564,In_885);
nor U2097 (N_2097,In_646,In_405);
and U2098 (N_2098,In_140,In_1080);
nand U2099 (N_2099,In_1789,In_266);
and U2100 (N_2100,In_220,In_419);
or U2101 (N_2101,In_1907,In_1216);
nor U2102 (N_2102,In_1381,In_933);
nand U2103 (N_2103,In_44,In_971);
or U2104 (N_2104,In_1859,In_176);
nor U2105 (N_2105,In_333,In_801);
nor U2106 (N_2106,In_1314,In_891);
nand U2107 (N_2107,In_491,In_231);
nor U2108 (N_2108,In_165,In_447);
nand U2109 (N_2109,In_158,In_1036);
and U2110 (N_2110,In_1254,In_539);
or U2111 (N_2111,In_778,In_1754);
and U2112 (N_2112,In_1764,In_1500);
and U2113 (N_2113,In_90,In_1085);
nor U2114 (N_2114,In_1869,In_84);
or U2115 (N_2115,In_956,In_642);
nand U2116 (N_2116,In_1734,In_15);
or U2117 (N_2117,In_1326,In_1721);
or U2118 (N_2118,In_1534,In_1122);
nand U2119 (N_2119,In_1780,In_1668);
nand U2120 (N_2120,In_1933,In_37);
nand U2121 (N_2121,In_823,In_1054);
nor U2122 (N_2122,In_1181,In_901);
or U2123 (N_2123,In_630,In_1561);
or U2124 (N_2124,In_81,In_1064);
and U2125 (N_2125,In_1365,In_1316);
and U2126 (N_2126,In_122,In_1653);
nor U2127 (N_2127,In_1485,In_1595);
or U2128 (N_2128,In_866,In_567);
nand U2129 (N_2129,In_1651,In_66);
nor U2130 (N_2130,In_533,In_1950);
and U2131 (N_2131,In_1706,In_988);
nor U2132 (N_2132,In_1598,In_433);
nand U2133 (N_2133,In_373,In_273);
nand U2134 (N_2134,In_1652,In_1070);
and U2135 (N_2135,In_1460,In_358);
nor U2136 (N_2136,In_663,In_190);
nor U2137 (N_2137,In_1349,In_868);
nand U2138 (N_2138,In_1548,In_257);
or U2139 (N_2139,In_1160,In_520);
nand U2140 (N_2140,In_948,In_88);
and U2141 (N_2141,In_1537,In_1539);
and U2142 (N_2142,In_994,In_1895);
or U2143 (N_2143,In_792,In_1682);
nand U2144 (N_2144,In_1516,In_1695);
nor U2145 (N_2145,In_156,In_1036);
and U2146 (N_2146,In_440,In_1997);
or U2147 (N_2147,In_1112,In_720);
nand U2148 (N_2148,In_526,In_1007);
and U2149 (N_2149,In_1762,In_30);
nor U2150 (N_2150,In_563,In_1172);
or U2151 (N_2151,In_1632,In_1914);
and U2152 (N_2152,In_764,In_105);
and U2153 (N_2153,In_952,In_1296);
or U2154 (N_2154,In_405,In_834);
or U2155 (N_2155,In_49,In_726);
nor U2156 (N_2156,In_1456,In_1880);
or U2157 (N_2157,In_972,In_261);
nand U2158 (N_2158,In_985,In_566);
nor U2159 (N_2159,In_71,In_1506);
and U2160 (N_2160,In_156,In_1649);
nand U2161 (N_2161,In_1558,In_1545);
nand U2162 (N_2162,In_252,In_148);
nand U2163 (N_2163,In_343,In_916);
nand U2164 (N_2164,In_1610,In_1596);
xor U2165 (N_2165,In_1151,In_1920);
or U2166 (N_2166,In_1152,In_1169);
nor U2167 (N_2167,In_128,In_1492);
xnor U2168 (N_2168,In_823,In_1392);
or U2169 (N_2169,In_498,In_1788);
nor U2170 (N_2170,In_493,In_357);
and U2171 (N_2171,In_1230,In_396);
nor U2172 (N_2172,In_7,In_1535);
or U2173 (N_2173,In_696,In_456);
nand U2174 (N_2174,In_529,In_1579);
and U2175 (N_2175,In_1466,In_472);
nand U2176 (N_2176,In_405,In_1119);
xor U2177 (N_2177,In_1996,In_436);
and U2178 (N_2178,In_1707,In_771);
nor U2179 (N_2179,In_1164,In_1747);
and U2180 (N_2180,In_67,In_1942);
or U2181 (N_2181,In_1673,In_1490);
and U2182 (N_2182,In_1546,In_664);
nor U2183 (N_2183,In_16,In_1941);
nor U2184 (N_2184,In_1129,In_367);
and U2185 (N_2185,In_1917,In_1970);
nor U2186 (N_2186,In_452,In_591);
or U2187 (N_2187,In_337,In_620);
and U2188 (N_2188,In_369,In_391);
nand U2189 (N_2189,In_1931,In_1299);
and U2190 (N_2190,In_214,In_247);
or U2191 (N_2191,In_86,In_60);
and U2192 (N_2192,In_628,In_661);
nor U2193 (N_2193,In_556,In_1050);
nand U2194 (N_2194,In_1338,In_1548);
nand U2195 (N_2195,In_536,In_1218);
and U2196 (N_2196,In_1513,In_1609);
nor U2197 (N_2197,In_1430,In_322);
and U2198 (N_2198,In_1623,In_291);
nor U2199 (N_2199,In_1120,In_710);
nand U2200 (N_2200,In_1323,In_330);
or U2201 (N_2201,In_1687,In_820);
nand U2202 (N_2202,In_1012,In_1356);
nor U2203 (N_2203,In_1005,In_333);
and U2204 (N_2204,In_785,In_504);
or U2205 (N_2205,In_1885,In_671);
or U2206 (N_2206,In_903,In_259);
nand U2207 (N_2207,In_900,In_552);
nor U2208 (N_2208,In_1546,In_105);
nor U2209 (N_2209,In_1702,In_1856);
and U2210 (N_2210,In_1098,In_535);
nor U2211 (N_2211,In_479,In_1961);
and U2212 (N_2212,In_956,In_572);
and U2213 (N_2213,In_337,In_298);
nor U2214 (N_2214,In_1829,In_604);
nand U2215 (N_2215,In_1675,In_1942);
and U2216 (N_2216,In_988,In_1709);
and U2217 (N_2217,In_666,In_553);
nor U2218 (N_2218,In_623,In_593);
or U2219 (N_2219,In_1105,In_1552);
and U2220 (N_2220,In_904,In_209);
or U2221 (N_2221,In_1921,In_1389);
nor U2222 (N_2222,In_700,In_456);
nand U2223 (N_2223,In_983,In_472);
nand U2224 (N_2224,In_18,In_1878);
nand U2225 (N_2225,In_1971,In_1216);
and U2226 (N_2226,In_1170,In_948);
nor U2227 (N_2227,In_287,In_225);
and U2228 (N_2228,In_1641,In_578);
nor U2229 (N_2229,In_1157,In_283);
and U2230 (N_2230,In_243,In_1710);
nor U2231 (N_2231,In_1295,In_1718);
or U2232 (N_2232,In_1730,In_720);
and U2233 (N_2233,In_1502,In_941);
nor U2234 (N_2234,In_190,In_62);
nor U2235 (N_2235,In_1630,In_610);
nand U2236 (N_2236,In_1525,In_1067);
nand U2237 (N_2237,In_539,In_1470);
nor U2238 (N_2238,In_1818,In_555);
and U2239 (N_2239,In_1234,In_83);
nand U2240 (N_2240,In_1561,In_866);
or U2241 (N_2241,In_416,In_1522);
nand U2242 (N_2242,In_284,In_131);
and U2243 (N_2243,In_943,In_947);
or U2244 (N_2244,In_88,In_611);
and U2245 (N_2245,In_1501,In_1419);
nor U2246 (N_2246,In_106,In_1415);
nor U2247 (N_2247,In_1866,In_486);
or U2248 (N_2248,In_1806,In_765);
or U2249 (N_2249,In_134,In_1657);
nand U2250 (N_2250,In_657,In_436);
and U2251 (N_2251,In_1844,In_452);
nor U2252 (N_2252,In_1771,In_1595);
or U2253 (N_2253,In_55,In_1243);
nand U2254 (N_2254,In_1491,In_1372);
nor U2255 (N_2255,In_827,In_526);
or U2256 (N_2256,In_1924,In_1550);
nand U2257 (N_2257,In_1590,In_1805);
nor U2258 (N_2258,In_1688,In_650);
and U2259 (N_2259,In_0,In_1070);
and U2260 (N_2260,In_551,In_1604);
nor U2261 (N_2261,In_1527,In_1837);
nand U2262 (N_2262,In_1347,In_401);
or U2263 (N_2263,In_98,In_1841);
and U2264 (N_2264,In_189,In_1759);
nand U2265 (N_2265,In_499,In_1148);
and U2266 (N_2266,In_1045,In_1695);
nand U2267 (N_2267,In_1860,In_419);
or U2268 (N_2268,In_403,In_762);
and U2269 (N_2269,In_183,In_1855);
nand U2270 (N_2270,In_629,In_610);
or U2271 (N_2271,In_549,In_7);
nand U2272 (N_2272,In_645,In_1780);
nor U2273 (N_2273,In_1140,In_1110);
nor U2274 (N_2274,In_1271,In_252);
xnor U2275 (N_2275,In_25,In_522);
and U2276 (N_2276,In_1132,In_219);
nand U2277 (N_2277,In_1348,In_1590);
nor U2278 (N_2278,In_1155,In_451);
or U2279 (N_2279,In_1575,In_1288);
nor U2280 (N_2280,In_1444,In_1147);
or U2281 (N_2281,In_1305,In_1856);
or U2282 (N_2282,In_1165,In_1879);
nand U2283 (N_2283,In_447,In_604);
or U2284 (N_2284,In_1076,In_1055);
xor U2285 (N_2285,In_237,In_851);
and U2286 (N_2286,In_1606,In_1819);
and U2287 (N_2287,In_985,In_1185);
nand U2288 (N_2288,In_403,In_628);
or U2289 (N_2289,In_1357,In_1331);
nand U2290 (N_2290,In_359,In_115);
nand U2291 (N_2291,In_9,In_325);
nand U2292 (N_2292,In_1946,In_1754);
and U2293 (N_2293,In_1770,In_212);
nor U2294 (N_2294,In_1928,In_1263);
and U2295 (N_2295,In_318,In_1231);
or U2296 (N_2296,In_1782,In_1942);
or U2297 (N_2297,In_564,In_712);
nand U2298 (N_2298,In_1169,In_744);
nor U2299 (N_2299,In_766,In_800);
nand U2300 (N_2300,In_76,In_228);
or U2301 (N_2301,In_1805,In_285);
or U2302 (N_2302,In_516,In_468);
and U2303 (N_2303,In_236,In_1721);
and U2304 (N_2304,In_1270,In_1402);
and U2305 (N_2305,In_902,In_261);
or U2306 (N_2306,In_1592,In_1327);
and U2307 (N_2307,In_53,In_1450);
or U2308 (N_2308,In_948,In_1310);
or U2309 (N_2309,In_780,In_82);
nor U2310 (N_2310,In_572,In_249);
or U2311 (N_2311,In_586,In_1299);
nor U2312 (N_2312,In_437,In_455);
and U2313 (N_2313,In_490,In_906);
nand U2314 (N_2314,In_1884,In_1739);
nand U2315 (N_2315,In_932,In_1361);
or U2316 (N_2316,In_395,In_464);
nor U2317 (N_2317,In_729,In_992);
or U2318 (N_2318,In_1742,In_241);
or U2319 (N_2319,In_1443,In_260);
and U2320 (N_2320,In_480,In_1281);
or U2321 (N_2321,In_295,In_1063);
and U2322 (N_2322,In_82,In_422);
nor U2323 (N_2323,In_1999,In_1958);
and U2324 (N_2324,In_35,In_1458);
nand U2325 (N_2325,In_869,In_1630);
nor U2326 (N_2326,In_188,In_416);
nor U2327 (N_2327,In_1295,In_1914);
or U2328 (N_2328,In_881,In_19);
or U2329 (N_2329,In_420,In_31);
and U2330 (N_2330,In_1819,In_526);
and U2331 (N_2331,In_773,In_868);
nand U2332 (N_2332,In_16,In_336);
xor U2333 (N_2333,In_1212,In_1884);
and U2334 (N_2334,In_1367,In_1488);
nand U2335 (N_2335,In_1258,In_1033);
and U2336 (N_2336,In_280,In_563);
and U2337 (N_2337,In_1645,In_1158);
or U2338 (N_2338,In_1787,In_741);
nand U2339 (N_2339,In_1029,In_1710);
and U2340 (N_2340,In_458,In_820);
and U2341 (N_2341,In_732,In_1825);
nand U2342 (N_2342,In_1786,In_956);
and U2343 (N_2343,In_538,In_817);
or U2344 (N_2344,In_179,In_485);
nor U2345 (N_2345,In_509,In_580);
nor U2346 (N_2346,In_582,In_1196);
and U2347 (N_2347,In_560,In_964);
and U2348 (N_2348,In_1512,In_1434);
nor U2349 (N_2349,In_627,In_338);
and U2350 (N_2350,In_1704,In_1365);
nand U2351 (N_2351,In_92,In_303);
xnor U2352 (N_2352,In_1639,In_897);
nand U2353 (N_2353,In_10,In_882);
nand U2354 (N_2354,In_41,In_1207);
nor U2355 (N_2355,In_139,In_319);
and U2356 (N_2356,In_1056,In_1949);
or U2357 (N_2357,In_1885,In_1717);
nand U2358 (N_2358,In_1171,In_1118);
nor U2359 (N_2359,In_1912,In_1388);
and U2360 (N_2360,In_834,In_1071);
or U2361 (N_2361,In_1263,In_500);
and U2362 (N_2362,In_703,In_1372);
and U2363 (N_2363,In_1624,In_950);
nand U2364 (N_2364,In_855,In_554);
nand U2365 (N_2365,In_762,In_1291);
or U2366 (N_2366,In_508,In_1305);
and U2367 (N_2367,In_287,In_1353);
nor U2368 (N_2368,In_323,In_329);
or U2369 (N_2369,In_1358,In_729);
nor U2370 (N_2370,In_802,In_1787);
and U2371 (N_2371,In_1018,In_690);
or U2372 (N_2372,In_866,In_824);
or U2373 (N_2373,In_1145,In_1226);
nor U2374 (N_2374,In_808,In_124);
nor U2375 (N_2375,In_55,In_229);
and U2376 (N_2376,In_102,In_1289);
nor U2377 (N_2377,In_1697,In_1001);
or U2378 (N_2378,In_1307,In_1014);
nand U2379 (N_2379,In_1923,In_1663);
nand U2380 (N_2380,In_1722,In_744);
or U2381 (N_2381,In_1395,In_1358);
nand U2382 (N_2382,In_1863,In_1540);
nor U2383 (N_2383,In_518,In_898);
nor U2384 (N_2384,In_1382,In_1053);
and U2385 (N_2385,In_865,In_768);
or U2386 (N_2386,In_1720,In_225);
or U2387 (N_2387,In_1025,In_1903);
nor U2388 (N_2388,In_910,In_1807);
or U2389 (N_2389,In_1119,In_1380);
or U2390 (N_2390,In_1157,In_280);
nand U2391 (N_2391,In_771,In_219);
nand U2392 (N_2392,In_25,In_1339);
nand U2393 (N_2393,In_180,In_916);
nand U2394 (N_2394,In_1101,In_1307);
or U2395 (N_2395,In_1651,In_1205);
and U2396 (N_2396,In_1245,In_1532);
and U2397 (N_2397,In_109,In_1025);
nand U2398 (N_2398,In_607,In_635);
nand U2399 (N_2399,In_1944,In_931);
nand U2400 (N_2400,In_1127,In_1987);
and U2401 (N_2401,In_1185,In_1284);
or U2402 (N_2402,In_1631,In_944);
and U2403 (N_2403,In_1437,In_735);
or U2404 (N_2404,In_1743,In_518);
nor U2405 (N_2405,In_314,In_706);
xor U2406 (N_2406,In_1472,In_1354);
or U2407 (N_2407,In_1058,In_508);
nand U2408 (N_2408,In_991,In_1538);
or U2409 (N_2409,In_607,In_1457);
or U2410 (N_2410,In_1569,In_1380);
or U2411 (N_2411,In_942,In_172);
and U2412 (N_2412,In_1355,In_1207);
or U2413 (N_2413,In_349,In_34);
and U2414 (N_2414,In_455,In_413);
nor U2415 (N_2415,In_1954,In_906);
and U2416 (N_2416,In_354,In_314);
nor U2417 (N_2417,In_1166,In_965);
nand U2418 (N_2418,In_254,In_1321);
or U2419 (N_2419,In_493,In_550);
nor U2420 (N_2420,In_1058,In_1646);
or U2421 (N_2421,In_972,In_1436);
and U2422 (N_2422,In_371,In_469);
and U2423 (N_2423,In_217,In_836);
or U2424 (N_2424,In_123,In_1386);
and U2425 (N_2425,In_479,In_1073);
or U2426 (N_2426,In_1235,In_392);
nand U2427 (N_2427,In_307,In_868);
nor U2428 (N_2428,In_1826,In_719);
nor U2429 (N_2429,In_529,In_551);
nor U2430 (N_2430,In_1221,In_1755);
xnor U2431 (N_2431,In_1987,In_293);
or U2432 (N_2432,In_603,In_1958);
nor U2433 (N_2433,In_25,In_1476);
nand U2434 (N_2434,In_1455,In_902);
nand U2435 (N_2435,In_1011,In_1426);
or U2436 (N_2436,In_943,In_1930);
nor U2437 (N_2437,In_1203,In_1778);
or U2438 (N_2438,In_1144,In_1841);
nor U2439 (N_2439,In_1973,In_1824);
nand U2440 (N_2440,In_855,In_1900);
and U2441 (N_2441,In_202,In_1641);
nand U2442 (N_2442,In_362,In_126);
nor U2443 (N_2443,In_1210,In_384);
nor U2444 (N_2444,In_1684,In_1836);
nor U2445 (N_2445,In_1696,In_1817);
nand U2446 (N_2446,In_1620,In_824);
nor U2447 (N_2447,In_351,In_1318);
nor U2448 (N_2448,In_1610,In_77);
nand U2449 (N_2449,In_642,In_271);
nor U2450 (N_2450,In_1383,In_814);
nor U2451 (N_2451,In_1660,In_851);
nor U2452 (N_2452,In_1479,In_139);
nor U2453 (N_2453,In_1123,In_1564);
or U2454 (N_2454,In_231,In_922);
nor U2455 (N_2455,In_1131,In_239);
nor U2456 (N_2456,In_1343,In_783);
or U2457 (N_2457,In_1104,In_679);
nor U2458 (N_2458,In_340,In_1108);
nor U2459 (N_2459,In_1574,In_248);
nand U2460 (N_2460,In_47,In_436);
or U2461 (N_2461,In_587,In_301);
nor U2462 (N_2462,In_1536,In_1164);
nand U2463 (N_2463,In_126,In_911);
and U2464 (N_2464,In_956,In_651);
or U2465 (N_2465,In_816,In_1487);
and U2466 (N_2466,In_1543,In_65);
nand U2467 (N_2467,In_1943,In_20);
and U2468 (N_2468,In_546,In_862);
and U2469 (N_2469,In_209,In_769);
or U2470 (N_2470,In_686,In_840);
nor U2471 (N_2471,In_1964,In_1034);
and U2472 (N_2472,In_1199,In_1957);
nand U2473 (N_2473,In_999,In_1411);
or U2474 (N_2474,In_1250,In_1184);
nor U2475 (N_2475,In_178,In_659);
nand U2476 (N_2476,In_1278,In_1041);
and U2477 (N_2477,In_231,In_1248);
nor U2478 (N_2478,In_342,In_1942);
or U2479 (N_2479,In_1731,In_369);
and U2480 (N_2480,In_1932,In_844);
nor U2481 (N_2481,In_480,In_1332);
nand U2482 (N_2482,In_443,In_1514);
or U2483 (N_2483,In_1152,In_683);
nor U2484 (N_2484,In_333,In_1836);
nor U2485 (N_2485,In_1108,In_774);
nor U2486 (N_2486,In_1852,In_1247);
nor U2487 (N_2487,In_225,In_1742);
xor U2488 (N_2488,In_1327,In_572);
nand U2489 (N_2489,In_998,In_80);
nand U2490 (N_2490,In_660,In_1718);
or U2491 (N_2491,In_1535,In_378);
or U2492 (N_2492,In_138,In_477);
nand U2493 (N_2493,In_422,In_376);
nand U2494 (N_2494,In_326,In_756);
xnor U2495 (N_2495,In_853,In_654);
and U2496 (N_2496,In_357,In_175);
and U2497 (N_2497,In_1395,In_1272);
or U2498 (N_2498,In_1307,In_224);
nor U2499 (N_2499,In_122,In_1273);
nor U2500 (N_2500,In_1468,In_1309);
nand U2501 (N_2501,In_431,In_283);
nor U2502 (N_2502,In_1728,In_1321);
or U2503 (N_2503,In_1400,In_669);
nand U2504 (N_2504,In_958,In_452);
and U2505 (N_2505,In_810,In_1797);
nor U2506 (N_2506,In_361,In_207);
or U2507 (N_2507,In_250,In_697);
and U2508 (N_2508,In_19,In_1238);
xnor U2509 (N_2509,In_386,In_740);
or U2510 (N_2510,In_684,In_231);
and U2511 (N_2511,In_122,In_1312);
and U2512 (N_2512,In_510,In_322);
or U2513 (N_2513,In_1168,In_531);
and U2514 (N_2514,In_632,In_442);
nor U2515 (N_2515,In_838,In_1450);
and U2516 (N_2516,In_625,In_264);
or U2517 (N_2517,In_362,In_209);
nor U2518 (N_2518,In_1482,In_1588);
nand U2519 (N_2519,In_1043,In_941);
nor U2520 (N_2520,In_1005,In_1160);
or U2521 (N_2521,In_6,In_87);
and U2522 (N_2522,In_1943,In_1480);
and U2523 (N_2523,In_307,In_1182);
and U2524 (N_2524,In_1613,In_1359);
nand U2525 (N_2525,In_444,In_1471);
nor U2526 (N_2526,In_1976,In_164);
and U2527 (N_2527,In_1328,In_1070);
and U2528 (N_2528,In_1188,In_1060);
and U2529 (N_2529,In_166,In_629);
nand U2530 (N_2530,In_778,In_675);
and U2531 (N_2531,In_568,In_735);
nor U2532 (N_2532,In_1731,In_1187);
and U2533 (N_2533,In_1208,In_1702);
or U2534 (N_2534,In_1748,In_1986);
and U2535 (N_2535,In_775,In_1588);
or U2536 (N_2536,In_1187,In_317);
nor U2537 (N_2537,In_757,In_416);
or U2538 (N_2538,In_982,In_533);
and U2539 (N_2539,In_717,In_52);
and U2540 (N_2540,In_795,In_1460);
or U2541 (N_2541,In_441,In_110);
nand U2542 (N_2542,In_1350,In_1264);
and U2543 (N_2543,In_857,In_1091);
nand U2544 (N_2544,In_1105,In_1993);
and U2545 (N_2545,In_1341,In_713);
and U2546 (N_2546,In_1732,In_1741);
nand U2547 (N_2547,In_1261,In_1258);
nor U2548 (N_2548,In_1096,In_687);
and U2549 (N_2549,In_54,In_1181);
and U2550 (N_2550,In_538,In_1536);
nor U2551 (N_2551,In_1078,In_564);
nand U2552 (N_2552,In_776,In_1547);
or U2553 (N_2553,In_93,In_1945);
or U2554 (N_2554,In_1903,In_1590);
nand U2555 (N_2555,In_322,In_1245);
nor U2556 (N_2556,In_95,In_685);
and U2557 (N_2557,In_1925,In_107);
or U2558 (N_2558,In_396,In_373);
and U2559 (N_2559,In_524,In_1513);
or U2560 (N_2560,In_743,In_1701);
nor U2561 (N_2561,In_1052,In_500);
nand U2562 (N_2562,In_1259,In_1122);
nand U2563 (N_2563,In_350,In_1984);
nand U2564 (N_2564,In_727,In_986);
nand U2565 (N_2565,In_221,In_174);
or U2566 (N_2566,In_1099,In_147);
and U2567 (N_2567,In_1148,In_633);
nand U2568 (N_2568,In_1888,In_919);
nor U2569 (N_2569,In_533,In_123);
or U2570 (N_2570,In_1358,In_979);
or U2571 (N_2571,In_568,In_683);
nor U2572 (N_2572,In_1961,In_554);
nand U2573 (N_2573,In_290,In_199);
nor U2574 (N_2574,In_544,In_1054);
or U2575 (N_2575,In_1003,In_1533);
and U2576 (N_2576,In_1576,In_1159);
nor U2577 (N_2577,In_937,In_1915);
nor U2578 (N_2578,In_1716,In_637);
or U2579 (N_2579,In_655,In_356);
nand U2580 (N_2580,In_890,In_398);
and U2581 (N_2581,In_1447,In_905);
or U2582 (N_2582,In_1852,In_258);
nor U2583 (N_2583,In_1684,In_114);
and U2584 (N_2584,In_890,In_354);
nand U2585 (N_2585,In_987,In_1829);
and U2586 (N_2586,In_440,In_1840);
nor U2587 (N_2587,In_1231,In_724);
nor U2588 (N_2588,In_1576,In_20);
nand U2589 (N_2589,In_926,In_1226);
or U2590 (N_2590,In_1955,In_1076);
or U2591 (N_2591,In_1644,In_628);
and U2592 (N_2592,In_1139,In_1254);
nand U2593 (N_2593,In_39,In_1183);
nand U2594 (N_2594,In_820,In_1205);
and U2595 (N_2595,In_1400,In_1488);
or U2596 (N_2596,In_1036,In_278);
nand U2597 (N_2597,In_981,In_1694);
and U2598 (N_2598,In_1325,In_1390);
nand U2599 (N_2599,In_621,In_654);
and U2600 (N_2600,In_1238,In_582);
and U2601 (N_2601,In_1255,In_1978);
and U2602 (N_2602,In_1182,In_1714);
or U2603 (N_2603,In_806,In_1744);
nor U2604 (N_2604,In_325,In_1173);
and U2605 (N_2605,In_760,In_173);
and U2606 (N_2606,In_1554,In_1125);
nor U2607 (N_2607,In_813,In_146);
or U2608 (N_2608,In_934,In_903);
nand U2609 (N_2609,In_866,In_1130);
nand U2610 (N_2610,In_1174,In_496);
or U2611 (N_2611,In_615,In_337);
or U2612 (N_2612,In_1891,In_1079);
and U2613 (N_2613,In_1417,In_1075);
or U2614 (N_2614,In_1879,In_1657);
or U2615 (N_2615,In_1739,In_1988);
and U2616 (N_2616,In_1686,In_1074);
or U2617 (N_2617,In_1398,In_1172);
and U2618 (N_2618,In_80,In_385);
nor U2619 (N_2619,In_1616,In_1571);
nor U2620 (N_2620,In_1922,In_324);
or U2621 (N_2621,In_1681,In_75);
or U2622 (N_2622,In_756,In_887);
nor U2623 (N_2623,In_306,In_806);
nor U2624 (N_2624,In_364,In_398);
or U2625 (N_2625,In_541,In_811);
nand U2626 (N_2626,In_409,In_1945);
or U2627 (N_2627,In_407,In_635);
and U2628 (N_2628,In_51,In_979);
or U2629 (N_2629,In_1720,In_1385);
nor U2630 (N_2630,In_205,In_270);
nor U2631 (N_2631,In_432,In_11);
nand U2632 (N_2632,In_466,In_1646);
or U2633 (N_2633,In_469,In_1116);
nor U2634 (N_2634,In_578,In_1935);
nor U2635 (N_2635,In_31,In_1828);
nor U2636 (N_2636,In_881,In_1462);
nor U2637 (N_2637,In_633,In_424);
or U2638 (N_2638,In_1074,In_305);
nand U2639 (N_2639,In_725,In_1450);
nor U2640 (N_2640,In_448,In_1440);
and U2641 (N_2641,In_311,In_49);
nand U2642 (N_2642,In_1139,In_1918);
nand U2643 (N_2643,In_772,In_1520);
or U2644 (N_2644,In_1756,In_257);
nor U2645 (N_2645,In_1543,In_1353);
or U2646 (N_2646,In_364,In_1041);
and U2647 (N_2647,In_468,In_845);
nor U2648 (N_2648,In_104,In_707);
nand U2649 (N_2649,In_682,In_1996);
or U2650 (N_2650,In_1335,In_267);
and U2651 (N_2651,In_1415,In_1425);
or U2652 (N_2652,In_365,In_1489);
nand U2653 (N_2653,In_1694,In_654);
nand U2654 (N_2654,In_1918,In_770);
nand U2655 (N_2655,In_126,In_642);
nor U2656 (N_2656,In_1496,In_1551);
nand U2657 (N_2657,In_1049,In_1779);
nand U2658 (N_2658,In_536,In_711);
nand U2659 (N_2659,In_881,In_478);
or U2660 (N_2660,In_1929,In_1956);
or U2661 (N_2661,In_1124,In_380);
or U2662 (N_2662,In_701,In_1158);
and U2663 (N_2663,In_1116,In_852);
and U2664 (N_2664,In_901,In_1056);
and U2665 (N_2665,In_799,In_1084);
or U2666 (N_2666,In_1870,In_1937);
and U2667 (N_2667,In_1648,In_154);
nor U2668 (N_2668,In_611,In_1034);
nand U2669 (N_2669,In_861,In_945);
or U2670 (N_2670,In_115,In_147);
nor U2671 (N_2671,In_1375,In_557);
and U2672 (N_2672,In_251,In_1592);
nand U2673 (N_2673,In_1104,In_34);
and U2674 (N_2674,In_1438,In_1321);
nor U2675 (N_2675,In_1730,In_1382);
or U2676 (N_2676,In_1978,In_810);
or U2677 (N_2677,In_857,In_117);
or U2678 (N_2678,In_264,In_185);
nand U2679 (N_2679,In_236,In_984);
nor U2680 (N_2680,In_1751,In_1399);
and U2681 (N_2681,In_594,In_1622);
nand U2682 (N_2682,In_199,In_979);
nand U2683 (N_2683,In_1723,In_1938);
and U2684 (N_2684,In_1264,In_349);
nand U2685 (N_2685,In_392,In_1146);
nor U2686 (N_2686,In_635,In_1940);
or U2687 (N_2687,In_49,In_843);
and U2688 (N_2688,In_1408,In_377);
or U2689 (N_2689,In_171,In_973);
nand U2690 (N_2690,In_825,In_1246);
and U2691 (N_2691,In_1881,In_1420);
xor U2692 (N_2692,In_293,In_1685);
nand U2693 (N_2693,In_1102,In_31);
or U2694 (N_2694,In_1840,In_1087);
and U2695 (N_2695,In_1943,In_410);
or U2696 (N_2696,In_984,In_1104);
and U2697 (N_2697,In_941,In_133);
nor U2698 (N_2698,In_256,In_1681);
nor U2699 (N_2699,In_30,In_1055);
nor U2700 (N_2700,In_200,In_1123);
nand U2701 (N_2701,In_345,In_546);
nor U2702 (N_2702,In_1494,In_472);
or U2703 (N_2703,In_148,In_1229);
nor U2704 (N_2704,In_472,In_1605);
nand U2705 (N_2705,In_1893,In_774);
nor U2706 (N_2706,In_1027,In_1457);
or U2707 (N_2707,In_1838,In_472);
and U2708 (N_2708,In_1710,In_169);
and U2709 (N_2709,In_146,In_671);
and U2710 (N_2710,In_1138,In_231);
and U2711 (N_2711,In_1250,In_654);
nor U2712 (N_2712,In_227,In_1139);
and U2713 (N_2713,In_533,In_1000);
nor U2714 (N_2714,In_1376,In_1809);
or U2715 (N_2715,In_1312,In_125);
nor U2716 (N_2716,In_1857,In_1463);
or U2717 (N_2717,In_908,In_1307);
and U2718 (N_2718,In_434,In_1515);
and U2719 (N_2719,In_47,In_1421);
and U2720 (N_2720,In_1583,In_911);
nand U2721 (N_2721,In_1732,In_838);
or U2722 (N_2722,In_1916,In_543);
nor U2723 (N_2723,In_1028,In_1454);
nor U2724 (N_2724,In_1240,In_1820);
nand U2725 (N_2725,In_212,In_1087);
and U2726 (N_2726,In_494,In_816);
and U2727 (N_2727,In_853,In_1414);
and U2728 (N_2728,In_1526,In_1513);
or U2729 (N_2729,In_84,In_20);
nor U2730 (N_2730,In_1448,In_1800);
nor U2731 (N_2731,In_1593,In_745);
or U2732 (N_2732,In_341,In_917);
nor U2733 (N_2733,In_1052,In_705);
nand U2734 (N_2734,In_1646,In_1070);
nand U2735 (N_2735,In_401,In_326);
nor U2736 (N_2736,In_790,In_918);
nand U2737 (N_2737,In_540,In_1067);
nand U2738 (N_2738,In_1300,In_270);
or U2739 (N_2739,In_121,In_442);
nor U2740 (N_2740,In_920,In_1779);
xor U2741 (N_2741,In_445,In_535);
and U2742 (N_2742,In_427,In_173);
or U2743 (N_2743,In_1752,In_1476);
or U2744 (N_2744,In_40,In_1676);
and U2745 (N_2745,In_1784,In_767);
nor U2746 (N_2746,In_1139,In_1056);
nor U2747 (N_2747,In_1273,In_682);
nand U2748 (N_2748,In_998,In_99);
or U2749 (N_2749,In_596,In_737);
or U2750 (N_2750,In_368,In_1312);
nand U2751 (N_2751,In_526,In_295);
or U2752 (N_2752,In_653,In_1021);
nor U2753 (N_2753,In_845,In_350);
or U2754 (N_2754,In_1290,In_132);
nand U2755 (N_2755,In_280,In_1008);
or U2756 (N_2756,In_794,In_1113);
and U2757 (N_2757,In_1036,In_1386);
nand U2758 (N_2758,In_1341,In_1008);
and U2759 (N_2759,In_1147,In_467);
or U2760 (N_2760,In_1154,In_622);
nand U2761 (N_2761,In_1809,In_675);
nand U2762 (N_2762,In_1027,In_1038);
nor U2763 (N_2763,In_1885,In_1709);
nor U2764 (N_2764,In_1037,In_1077);
or U2765 (N_2765,In_1919,In_1322);
nor U2766 (N_2766,In_390,In_546);
or U2767 (N_2767,In_809,In_1999);
nor U2768 (N_2768,In_607,In_900);
nor U2769 (N_2769,In_451,In_806);
and U2770 (N_2770,In_1686,In_1090);
and U2771 (N_2771,In_1866,In_1816);
nor U2772 (N_2772,In_224,In_530);
nand U2773 (N_2773,In_643,In_1959);
or U2774 (N_2774,In_176,In_501);
nor U2775 (N_2775,In_1830,In_228);
or U2776 (N_2776,In_941,In_1578);
nand U2777 (N_2777,In_1663,In_992);
xor U2778 (N_2778,In_521,In_1024);
nand U2779 (N_2779,In_1541,In_105);
nor U2780 (N_2780,In_1655,In_583);
and U2781 (N_2781,In_185,In_1590);
and U2782 (N_2782,In_1769,In_1518);
nor U2783 (N_2783,In_901,In_1791);
nand U2784 (N_2784,In_1739,In_136);
or U2785 (N_2785,In_1599,In_1240);
nand U2786 (N_2786,In_1539,In_1906);
nand U2787 (N_2787,In_1186,In_1538);
and U2788 (N_2788,In_276,In_1622);
or U2789 (N_2789,In_586,In_33);
xor U2790 (N_2790,In_244,In_573);
nor U2791 (N_2791,In_671,In_385);
nand U2792 (N_2792,In_218,In_1198);
nor U2793 (N_2793,In_1254,In_1346);
and U2794 (N_2794,In_1857,In_97);
nor U2795 (N_2795,In_665,In_244);
and U2796 (N_2796,In_698,In_940);
nor U2797 (N_2797,In_122,In_1057);
nor U2798 (N_2798,In_1617,In_1727);
nand U2799 (N_2799,In_1968,In_1658);
and U2800 (N_2800,In_1835,In_1685);
or U2801 (N_2801,In_862,In_1060);
or U2802 (N_2802,In_831,In_982);
nand U2803 (N_2803,In_1562,In_1322);
or U2804 (N_2804,In_1565,In_1421);
and U2805 (N_2805,In_201,In_730);
nor U2806 (N_2806,In_880,In_639);
nor U2807 (N_2807,In_264,In_960);
or U2808 (N_2808,In_1129,In_659);
and U2809 (N_2809,In_863,In_703);
nor U2810 (N_2810,In_766,In_1894);
nand U2811 (N_2811,In_1973,In_999);
nand U2812 (N_2812,In_1329,In_1427);
or U2813 (N_2813,In_385,In_1153);
and U2814 (N_2814,In_1687,In_1784);
and U2815 (N_2815,In_981,In_845);
or U2816 (N_2816,In_850,In_1538);
nor U2817 (N_2817,In_1068,In_1704);
nor U2818 (N_2818,In_1286,In_1388);
or U2819 (N_2819,In_1304,In_486);
nor U2820 (N_2820,In_1528,In_1445);
and U2821 (N_2821,In_1207,In_964);
nor U2822 (N_2822,In_578,In_1877);
nor U2823 (N_2823,In_331,In_1704);
nor U2824 (N_2824,In_787,In_424);
nand U2825 (N_2825,In_710,In_508);
nor U2826 (N_2826,In_469,In_1741);
nor U2827 (N_2827,In_1870,In_584);
or U2828 (N_2828,In_663,In_428);
nor U2829 (N_2829,In_947,In_7);
nand U2830 (N_2830,In_1255,In_171);
or U2831 (N_2831,In_1379,In_127);
or U2832 (N_2832,In_619,In_1531);
nand U2833 (N_2833,In_636,In_1363);
nand U2834 (N_2834,In_300,In_1174);
or U2835 (N_2835,In_1536,In_1535);
nand U2836 (N_2836,In_1732,In_891);
nor U2837 (N_2837,In_152,In_845);
xnor U2838 (N_2838,In_254,In_909);
and U2839 (N_2839,In_1379,In_627);
nand U2840 (N_2840,In_789,In_567);
nand U2841 (N_2841,In_1303,In_1439);
nor U2842 (N_2842,In_76,In_666);
or U2843 (N_2843,In_270,In_274);
or U2844 (N_2844,In_950,In_1792);
nand U2845 (N_2845,In_1009,In_650);
nor U2846 (N_2846,In_1474,In_758);
nor U2847 (N_2847,In_1104,In_1071);
or U2848 (N_2848,In_1723,In_390);
and U2849 (N_2849,In_399,In_688);
nor U2850 (N_2850,In_425,In_1410);
and U2851 (N_2851,In_1533,In_869);
xnor U2852 (N_2852,In_1562,In_1206);
and U2853 (N_2853,In_1088,In_1140);
nor U2854 (N_2854,In_1483,In_1067);
or U2855 (N_2855,In_1290,In_1372);
and U2856 (N_2856,In_1128,In_1078);
or U2857 (N_2857,In_1039,In_314);
or U2858 (N_2858,In_201,In_312);
nand U2859 (N_2859,In_281,In_1555);
and U2860 (N_2860,In_85,In_509);
nand U2861 (N_2861,In_828,In_411);
and U2862 (N_2862,In_115,In_1090);
and U2863 (N_2863,In_1121,In_126);
or U2864 (N_2864,In_1643,In_672);
and U2865 (N_2865,In_1824,In_1407);
nor U2866 (N_2866,In_921,In_655);
and U2867 (N_2867,In_1085,In_345);
nor U2868 (N_2868,In_416,In_1496);
xnor U2869 (N_2869,In_1011,In_1215);
or U2870 (N_2870,In_1701,In_1091);
nor U2871 (N_2871,In_700,In_586);
and U2872 (N_2872,In_615,In_1160);
nor U2873 (N_2873,In_1887,In_194);
nor U2874 (N_2874,In_296,In_361);
nand U2875 (N_2875,In_721,In_1414);
nor U2876 (N_2876,In_1931,In_1759);
and U2877 (N_2877,In_1047,In_763);
or U2878 (N_2878,In_1716,In_1563);
and U2879 (N_2879,In_382,In_1194);
and U2880 (N_2880,In_171,In_483);
nand U2881 (N_2881,In_697,In_666);
or U2882 (N_2882,In_1,In_774);
and U2883 (N_2883,In_1621,In_1956);
or U2884 (N_2884,In_980,In_380);
and U2885 (N_2885,In_354,In_253);
or U2886 (N_2886,In_1963,In_1456);
nand U2887 (N_2887,In_1443,In_1149);
and U2888 (N_2888,In_636,In_402);
or U2889 (N_2889,In_526,In_602);
nand U2890 (N_2890,In_1656,In_127);
or U2891 (N_2891,In_1941,In_1194);
or U2892 (N_2892,In_1809,In_463);
and U2893 (N_2893,In_669,In_1978);
or U2894 (N_2894,In_396,In_770);
or U2895 (N_2895,In_368,In_448);
nand U2896 (N_2896,In_2,In_180);
and U2897 (N_2897,In_937,In_1549);
nor U2898 (N_2898,In_738,In_767);
or U2899 (N_2899,In_1845,In_578);
or U2900 (N_2900,In_389,In_831);
and U2901 (N_2901,In_1588,In_1857);
and U2902 (N_2902,In_488,In_1263);
or U2903 (N_2903,In_1855,In_1244);
nand U2904 (N_2904,In_629,In_1585);
and U2905 (N_2905,In_517,In_1300);
and U2906 (N_2906,In_953,In_1541);
or U2907 (N_2907,In_1922,In_32);
nor U2908 (N_2908,In_1393,In_1206);
nor U2909 (N_2909,In_753,In_563);
nor U2910 (N_2910,In_987,In_1072);
nand U2911 (N_2911,In_825,In_595);
nor U2912 (N_2912,In_433,In_1345);
and U2913 (N_2913,In_497,In_472);
and U2914 (N_2914,In_0,In_1417);
or U2915 (N_2915,In_1829,In_206);
nor U2916 (N_2916,In_881,In_1130);
and U2917 (N_2917,In_785,In_941);
nand U2918 (N_2918,In_1627,In_303);
nor U2919 (N_2919,In_159,In_734);
or U2920 (N_2920,In_499,In_417);
nand U2921 (N_2921,In_213,In_3);
nand U2922 (N_2922,In_1011,In_529);
and U2923 (N_2923,In_149,In_96);
nor U2924 (N_2924,In_1832,In_1232);
and U2925 (N_2925,In_227,In_1909);
and U2926 (N_2926,In_1879,In_648);
nand U2927 (N_2927,In_1335,In_1667);
nand U2928 (N_2928,In_613,In_889);
or U2929 (N_2929,In_828,In_544);
and U2930 (N_2930,In_367,In_1276);
or U2931 (N_2931,In_1727,In_332);
and U2932 (N_2932,In_81,In_644);
and U2933 (N_2933,In_1723,In_109);
nor U2934 (N_2934,In_1192,In_1511);
and U2935 (N_2935,In_1703,In_1670);
nand U2936 (N_2936,In_503,In_1003);
nor U2937 (N_2937,In_438,In_1474);
nor U2938 (N_2938,In_1033,In_1665);
and U2939 (N_2939,In_236,In_143);
nor U2940 (N_2940,In_697,In_122);
nand U2941 (N_2941,In_1662,In_1039);
nand U2942 (N_2942,In_981,In_1711);
nand U2943 (N_2943,In_1380,In_912);
nand U2944 (N_2944,In_1755,In_369);
and U2945 (N_2945,In_1624,In_1426);
nand U2946 (N_2946,In_426,In_1732);
nor U2947 (N_2947,In_519,In_146);
or U2948 (N_2948,In_99,In_1793);
or U2949 (N_2949,In_9,In_1915);
and U2950 (N_2950,In_594,In_1354);
nand U2951 (N_2951,In_703,In_318);
or U2952 (N_2952,In_1818,In_1002);
nor U2953 (N_2953,In_835,In_187);
nor U2954 (N_2954,In_499,In_1536);
nor U2955 (N_2955,In_1252,In_568);
nor U2956 (N_2956,In_1280,In_1885);
nor U2957 (N_2957,In_1260,In_851);
or U2958 (N_2958,In_183,In_452);
nand U2959 (N_2959,In_1153,In_1187);
nor U2960 (N_2960,In_274,In_1994);
nor U2961 (N_2961,In_1567,In_606);
and U2962 (N_2962,In_536,In_1701);
or U2963 (N_2963,In_451,In_270);
and U2964 (N_2964,In_976,In_854);
or U2965 (N_2965,In_1723,In_818);
nor U2966 (N_2966,In_1948,In_950);
or U2967 (N_2967,In_509,In_1208);
nand U2968 (N_2968,In_1965,In_213);
nor U2969 (N_2969,In_1135,In_1982);
and U2970 (N_2970,In_1198,In_1307);
nor U2971 (N_2971,In_1980,In_259);
or U2972 (N_2972,In_667,In_1223);
nand U2973 (N_2973,In_862,In_1909);
nor U2974 (N_2974,In_148,In_154);
nand U2975 (N_2975,In_1220,In_1981);
nor U2976 (N_2976,In_1002,In_1188);
nand U2977 (N_2977,In_1692,In_1148);
and U2978 (N_2978,In_366,In_595);
nand U2979 (N_2979,In_1353,In_1742);
or U2980 (N_2980,In_39,In_891);
nand U2981 (N_2981,In_747,In_656);
nand U2982 (N_2982,In_1971,In_1146);
nand U2983 (N_2983,In_1543,In_1521);
and U2984 (N_2984,In_49,In_1650);
or U2985 (N_2985,In_284,In_330);
nor U2986 (N_2986,In_675,In_1716);
nor U2987 (N_2987,In_1780,In_275);
or U2988 (N_2988,In_972,In_1012);
nor U2989 (N_2989,In_267,In_757);
and U2990 (N_2990,In_125,In_1015);
or U2991 (N_2991,In_1146,In_951);
nor U2992 (N_2992,In_129,In_1999);
nand U2993 (N_2993,In_1666,In_1799);
nand U2994 (N_2994,In_1218,In_429);
nor U2995 (N_2995,In_1187,In_1533);
and U2996 (N_2996,In_1545,In_1190);
and U2997 (N_2997,In_1133,In_191);
nor U2998 (N_2998,In_49,In_214);
and U2999 (N_2999,In_719,In_1957);
nand U3000 (N_3000,In_103,In_1045);
nand U3001 (N_3001,In_929,In_371);
and U3002 (N_3002,In_120,In_425);
nand U3003 (N_3003,In_1012,In_327);
nand U3004 (N_3004,In_1256,In_1738);
and U3005 (N_3005,In_1096,In_1328);
nor U3006 (N_3006,In_1668,In_1604);
nor U3007 (N_3007,In_1634,In_710);
and U3008 (N_3008,In_147,In_637);
and U3009 (N_3009,In_1659,In_50);
and U3010 (N_3010,In_94,In_239);
nand U3011 (N_3011,In_1736,In_888);
nor U3012 (N_3012,In_1649,In_492);
nor U3013 (N_3013,In_1692,In_1759);
nor U3014 (N_3014,In_1664,In_296);
and U3015 (N_3015,In_1040,In_12);
nand U3016 (N_3016,In_1721,In_1402);
nor U3017 (N_3017,In_973,In_493);
and U3018 (N_3018,In_1902,In_162);
nand U3019 (N_3019,In_416,In_1378);
and U3020 (N_3020,In_1038,In_400);
nor U3021 (N_3021,In_654,In_968);
nor U3022 (N_3022,In_1777,In_225);
nand U3023 (N_3023,In_257,In_244);
nor U3024 (N_3024,In_670,In_874);
and U3025 (N_3025,In_1266,In_307);
or U3026 (N_3026,In_931,In_339);
and U3027 (N_3027,In_736,In_864);
and U3028 (N_3028,In_736,In_522);
nor U3029 (N_3029,In_153,In_674);
and U3030 (N_3030,In_1072,In_790);
or U3031 (N_3031,In_1029,In_1830);
and U3032 (N_3032,In_1324,In_1270);
or U3033 (N_3033,In_462,In_1568);
or U3034 (N_3034,In_874,In_1497);
or U3035 (N_3035,In_46,In_1650);
nor U3036 (N_3036,In_1865,In_999);
and U3037 (N_3037,In_1237,In_641);
nand U3038 (N_3038,In_1993,In_1789);
or U3039 (N_3039,In_352,In_1810);
or U3040 (N_3040,In_159,In_361);
and U3041 (N_3041,In_1607,In_1604);
nand U3042 (N_3042,In_1759,In_39);
nand U3043 (N_3043,In_966,In_67);
nand U3044 (N_3044,In_1748,In_574);
and U3045 (N_3045,In_1236,In_691);
nand U3046 (N_3046,In_1559,In_377);
nor U3047 (N_3047,In_269,In_1633);
nand U3048 (N_3048,In_833,In_505);
nand U3049 (N_3049,In_184,In_929);
nand U3050 (N_3050,In_970,In_1124);
nor U3051 (N_3051,In_1058,In_1338);
nor U3052 (N_3052,In_1962,In_339);
or U3053 (N_3053,In_1566,In_933);
nand U3054 (N_3054,In_1277,In_559);
and U3055 (N_3055,In_1541,In_260);
nor U3056 (N_3056,In_1557,In_976);
and U3057 (N_3057,In_938,In_1154);
nand U3058 (N_3058,In_203,In_746);
nor U3059 (N_3059,In_1479,In_1389);
or U3060 (N_3060,In_974,In_131);
and U3061 (N_3061,In_80,In_311);
xor U3062 (N_3062,In_1788,In_91);
nand U3063 (N_3063,In_1506,In_224);
and U3064 (N_3064,In_338,In_1275);
nor U3065 (N_3065,In_388,In_151);
nand U3066 (N_3066,In_553,In_1491);
or U3067 (N_3067,In_1024,In_1183);
and U3068 (N_3068,In_682,In_1402);
and U3069 (N_3069,In_1061,In_1405);
nand U3070 (N_3070,In_1021,In_1896);
nor U3071 (N_3071,In_152,In_1811);
nor U3072 (N_3072,In_349,In_1786);
nand U3073 (N_3073,In_1335,In_540);
nor U3074 (N_3074,In_822,In_909);
nand U3075 (N_3075,In_1258,In_995);
nand U3076 (N_3076,In_1699,In_221);
or U3077 (N_3077,In_1640,In_964);
nand U3078 (N_3078,In_1398,In_1519);
and U3079 (N_3079,In_1665,In_1023);
nor U3080 (N_3080,In_209,In_1652);
or U3081 (N_3081,In_4,In_1073);
and U3082 (N_3082,In_81,In_97);
xor U3083 (N_3083,In_475,In_1054);
or U3084 (N_3084,In_650,In_661);
nor U3085 (N_3085,In_504,In_141);
nor U3086 (N_3086,In_366,In_809);
nor U3087 (N_3087,In_812,In_1197);
and U3088 (N_3088,In_184,In_1043);
nand U3089 (N_3089,In_1223,In_1210);
and U3090 (N_3090,In_792,In_239);
and U3091 (N_3091,In_1638,In_891);
or U3092 (N_3092,In_1066,In_3);
or U3093 (N_3093,In_1878,In_1179);
nor U3094 (N_3094,In_1271,In_881);
and U3095 (N_3095,In_695,In_472);
xnor U3096 (N_3096,In_371,In_214);
nor U3097 (N_3097,In_606,In_975);
nand U3098 (N_3098,In_43,In_1580);
and U3099 (N_3099,In_1269,In_893);
and U3100 (N_3100,In_909,In_207);
or U3101 (N_3101,In_1120,In_1391);
or U3102 (N_3102,In_1110,In_914);
nor U3103 (N_3103,In_1079,In_1463);
and U3104 (N_3104,In_50,In_40);
nor U3105 (N_3105,In_984,In_1570);
xor U3106 (N_3106,In_1070,In_575);
nand U3107 (N_3107,In_1342,In_600);
nor U3108 (N_3108,In_565,In_1437);
nor U3109 (N_3109,In_1743,In_1454);
or U3110 (N_3110,In_1606,In_868);
nor U3111 (N_3111,In_348,In_169);
nor U3112 (N_3112,In_1615,In_1104);
nor U3113 (N_3113,In_146,In_342);
nand U3114 (N_3114,In_1670,In_904);
nor U3115 (N_3115,In_1199,In_1799);
and U3116 (N_3116,In_1519,In_1195);
or U3117 (N_3117,In_1596,In_762);
or U3118 (N_3118,In_579,In_1036);
and U3119 (N_3119,In_484,In_1352);
and U3120 (N_3120,In_292,In_426);
or U3121 (N_3121,In_1504,In_3);
and U3122 (N_3122,In_242,In_1602);
nor U3123 (N_3123,In_195,In_1877);
and U3124 (N_3124,In_392,In_765);
nand U3125 (N_3125,In_1537,In_467);
nand U3126 (N_3126,In_1990,In_1977);
nand U3127 (N_3127,In_871,In_1930);
nand U3128 (N_3128,In_1889,In_3);
or U3129 (N_3129,In_1747,In_175);
or U3130 (N_3130,In_1090,In_1505);
nand U3131 (N_3131,In_450,In_873);
nand U3132 (N_3132,In_1432,In_1292);
nand U3133 (N_3133,In_1969,In_1301);
nand U3134 (N_3134,In_1173,In_1369);
or U3135 (N_3135,In_220,In_1495);
and U3136 (N_3136,In_581,In_1281);
or U3137 (N_3137,In_1255,In_790);
and U3138 (N_3138,In_1006,In_1942);
or U3139 (N_3139,In_288,In_203);
and U3140 (N_3140,In_1572,In_513);
nor U3141 (N_3141,In_1272,In_1994);
and U3142 (N_3142,In_312,In_1354);
or U3143 (N_3143,In_1527,In_794);
nand U3144 (N_3144,In_1691,In_1901);
nand U3145 (N_3145,In_308,In_1233);
and U3146 (N_3146,In_1213,In_1544);
nand U3147 (N_3147,In_722,In_847);
nand U3148 (N_3148,In_1941,In_593);
and U3149 (N_3149,In_424,In_1406);
or U3150 (N_3150,In_296,In_1314);
nor U3151 (N_3151,In_1340,In_1385);
nand U3152 (N_3152,In_1493,In_1068);
or U3153 (N_3153,In_1349,In_775);
nor U3154 (N_3154,In_154,In_235);
and U3155 (N_3155,In_437,In_1920);
or U3156 (N_3156,In_56,In_530);
nand U3157 (N_3157,In_490,In_1702);
nand U3158 (N_3158,In_935,In_1933);
nand U3159 (N_3159,In_72,In_746);
nand U3160 (N_3160,In_457,In_1380);
nor U3161 (N_3161,In_119,In_1364);
or U3162 (N_3162,In_360,In_602);
nand U3163 (N_3163,In_678,In_1423);
nand U3164 (N_3164,In_856,In_233);
and U3165 (N_3165,In_1445,In_88);
or U3166 (N_3166,In_1341,In_65);
nor U3167 (N_3167,In_15,In_383);
nor U3168 (N_3168,In_1508,In_1115);
nand U3169 (N_3169,In_690,In_286);
nand U3170 (N_3170,In_1017,In_1965);
and U3171 (N_3171,In_1840,In_718);
nand U3172 (N_3172,In_1918,In_1875);
nand U3173 (N_3173,In_1081,In_349);
nand U3174 (N_3174,In_925,In_40);
and U3175 (N_3175,In_822,In_1038);
or U3176 (N_3176,In_1358,In_1586);
or U3177 (N_3177,In_1736,In_1900);
nand U3178 (N_3178,In_542,In_100);
xor U3179 (N_3179,In_279,In_246);
or U3180 (N_3180,In_1785,In_899);
nand U3181 (N_3181,In_1095,In_1278);
nand U3182 (N_3182,In_310,In_1232);
nand U3183 (N_3183,In_1564,In_1387);
nor U3184 (N_3184,In_1366,In_1834);
nand U3185 (N_3185,In_1953,In_1156);
and U3186 (N_3186,In_960,In_33);
nand U3187 (N_3187,In_1797,In_1626);
nand U3188 (N_3188,In_1712,In_1101);
xor U3189 (N_3189,In_157,In_493);
and U3190 (N_3190,In_18,In_1711);
nor U3191 (N_3191,In_1165,In_767);
and U3192 (N_3192,In_616,In_1000);
nand U3193 (N_3193,In_258,In_348);
and U3194 (N_3194,In_1940,In_1279);
nor U3195 (N_3195,In_218,In_1481);
xnor U3196 (N_3196,In_278,In_1509);
or U3197 (N_3197,In_876,In_1406);
or U3198 (N_3198,In_320,In_1751);
or U3199 (N_3199,In_1202,In_1888);
nand U3200 (N_3200,In_410,In_665);
or U3201 (N_3201,In_1463,In_286);
or U3202 (N_3202,In_538,In_634);
nand U3203 (N_3203,In_1450,In_1428);
nor U3204 (N_3204,In_1073,In_936);
and U3205 (N_3205,In_798,In_187);
or U3206 (N_3206,In_823,In_1932);
or U3207 (N_3207,In_783,In_1426);
nor U3208 (N_3208,In_1708,In_1221);
xnor U3209 (N_3209,In_829,In_1841);
nor U3210 (N_3210,In_1159,In_766);
and U3211 (N_3211,In_1070,In_233);
nand U3212 (N_3212,In_1353,In_876);
and U3213 (N_3213,In_1729,In_949);
nor U3214 (N_3214,In_1131,In_123);
or U3215 (N_3215,In_1718,In_378);
or U3216 (N_3216,In_666,In_953);
xnor U3217 (N_3217,In_75,In_1726);
nand U3218 (N_3218,In_342,In_302);
or U3219 (N_3219,In_934,In_385);
nor U3220 (N_3220,In_1530,In_752);
or U3221 (N_3221,In_1256,In_657);
and U3222 (N_3222,In_637,In_1086);
nor U3223 (N_3223,In_674,In_891);
xor U3224 (N_3224,In_1063,In_418);
nand U3225 (N_3225,In_1246,In_448);
and U3226 (N_3226,In_1316,In_882);
nor U3227 (N_3227,In_1479,In_1156);
nor U3228 (N_3228,In_1579,In_493);
nand U3229 (N_3229,In_650,In_725);
nor U3230 (N_3230,In_47,In_155);
nor U3231 (N_3231,In_1713,In_283);
nand U3232 (N_3232,In_1164,In_637);
or U3233 (N_3233,In_420,In_1000);
nor U3234 (N_3234,In_602,In_1593);
nor U3235 (N_3235,In_1878,In_470);
and U3236 (N_3236,In_1322,In_705);
and U3237 (N_3237,In_291,In_1158);
nor U3238 (N_3238,In_1153,In_1718);
or U3239 (N_3239,In_1716,In_1867);
xor U3240 (N_3240,In_1901,In_830);
nor U3241 (N_3241,In_1876,In_440);
nand U3242 (N_3242,In_21,In_1921);
or U3243 (N_3243,In_28,In_974);
nor U3244 (N_3244,In_1792,In_1206);
nand U3245 (N_3245,In_1277,In_1459);
or U3246 (N_3246,In_141,In_932);
nor U3247 (N_3247,In_617,In_1467);
nor U3248 (N_3248,In_321,In_1921);
nand U3249 (N_3249,In_1052,In_1554);
nor U3250 (N_3250,In_316,In_808);
nand U3251 (N_3251,In_524,In_1915);
nor U3252 (N_3252,In_1710,In_393);
nand U3253 (N_3253,In_1732,In_602);
nand U3254 (N_3254,In_1367,In_1684);
nor U3255 (N_3255,In_1563,In_234);
or U3256 (N_3256,In_615,In_1045);
nor U3257 (N_3257,In_1405,In_434);
and U3258 (N_3258,In_1522,In_895);
nor U3259 (N_3259,In_1829,In_1131);
or U3260 (N_3260,In_44,In_408);
nand U3261 (N_3261,In_1562,In_1756);
nor U3262 (N_3262,In_245,In_286);
and U3263 (N_3263,In_536,In_1981);
or U3264 (N_3264,In_1113,In_226);
and U3265 (N_3265,In_431,In_1361);
or U3266 (N_3266,In_1552,In_906);
or U3267 (N_3267,In_1180,In_306);
and U3268 (N_3268,In_596,In_40);
or U3269 (N_3269,In_1274,In_1312);
nor U3270 (N_3270,In_1738,In_542);
and U3271 (N_3271,In_298,In_17);
nand U3272 (N_3272,In_1077,In_251);
nand U3273 (N_3273,In_1151,In_483);
nor U3274 (N_3274,In_1751,In_1840);
and U3275 (N_3275,In_1058,In_468);
nand U3276 (N_3276,In_784,In_857);
nor U3277 (N_3277,In_1061,In_1818);
nor U3278 (N_3278,In_1256,In_1852);
and U3279 (N_3279,In_888,In_1418);
nand U3280 (N_3280,In_365,In_684);
nor U3281 (N_3281,In_1450,In_255);
and U3282 (N_3282,In_976,In_928);
and U3283 (N_3283,In_548,In_770);
or U3284 (N_3284,In_1143,In_417);
or U3285 (N_3285,In_952,In_1261);
and U3286 (N_3286,In_1288,In_630);
or U3287 (N_3287,In_1166,In_294);
and U3288 (N_3288,In_1630,In_817);
nand U3289 (N_3289,In_1638,In_1061);
and U3290 (N_3290,In_789,In_1990);
and U3291 (N_3291,In_170,In_370);
and U3292 (N_3292,In_1562,In_860);
nor U3293 (N_3293,In_469,In_1958);
and U3294 (N_3294,In_144,In_349);
nand U3295 (N_3295,In_294,In_1992);
nand U3296 (N_3296,In_695,In_1298);
nor U3297 (N_3297,In_1820,In_275);
and U3298 (N_3298,In_1710,In_1711);
or U3299 (N_3299,In_637,In_769);
nand U3300 (N_3300,In_1291,In_857);
nand U3301 (N_3301,In_1618,In_480);
or U3302 (N_3302,In_1053,In_616);
nor U3303 (N_3303,In_1039,In_494);
nand U3304 (N_3304,In_722,In_1824);
nand U3305 (N_3305,In_1127,In_1205);
and U3306 (N_3306,In_1295,In_1957);
nor U3307 (N_3307,In_469,In_1174);
nand U3308 (N_3308,In_1359,In_83);
nand U3309 (N_3309,In_943,In_599);
and U3310 (N_3310,In_1756,In_118);
or U3311 (N_3311,In_1932,In_1419);
and U3312 (N_3312,In_622,In_1999);
nor U3313 (N_3313,In_1417,In_1052);
or U3314 (N_3314,In_1523,In_982);
nor U3315 (N_3315,In_307,In_270);
and U3316 (N_3316,In_36,In_1535);
or U3317 (N_3317,In_391,In_1838);
and U3318 (N_3318,In_357,In_45);
and U3319 (N_3319,In_126,In_1497);
or U3320 (N_3320,In_776,In_1350);
or U3321 (N_3321,In_701,In_1498);
nor U3322 (N_3322,In_475,In_427);
nand U3323 (N_3323,In_287,In_1313);
nor U3324 (N_3324,In_896,In_408);
nand U3325 (N_3325,In_1860,In_714);
nand U3326 (N_3326,In_313,In_1964);
nand U3327 (N_3327,In_753,In_1401);
and U3328 (N_3328,In_1182,In_834);
nand U3329 (N_3329,In_335,In_1063);
nand U3330 (N_3330,In_805,In_222);
and U3331 (N_3331,In_373,In_1156);
nand U3332 (N_3332,In_1159,In_964);
or U3333 (N_3333,In_1761,In_1701);
nor U3334 (N_3334,In_401,In_1360);
nand U3335 (N_3335,In_898,In_485);
nand U3336 (N_3336,In_1417,In_1547);
nand U3337 (N_3337,In_517,In_1681);
or U3338 (N_3338,In_1334,In_1271);
and U3339 (N_3339,In_1574,In_559);
nand U3340 (N_3340,In_1630,In_1000);
and U3341 (N_3341,In_877,In_316);
and U3342 (N_3342,In_1971,In_760);
or U3343 (N_3343,In_701,In_1516);
and U3344 (N_3344,In_1756,In_1717);
and U3345 (N_3345,In_958,In_1250);
nand U3346 (N_3346,In_825,In_1436);
nand U3347 (N_3347,In_1532,In_26);
nor U3348 (N_3348,In_1570,In_1925);
nor U3349 (N_3349,In_1946,In_560);
or U3350 (N_3350,In_333,In_1439);
or U3351 (N_3351,In_14,In_146);
nand U3352 (N_3352,In_30,In_1297);
nor U3353 (N_3353,In_1112,In_811);
nand U3354 (N_3354,In_1357,In_1822);
or U3355 (N_3355,In_691,In_39);
nor U3356 (N_3356,In_1137,In_516);
nor U3357 (N_3357,In_1450,In_428);
nand U3358 (N_3358,In_483,In_104);
nor U3359 (N_3359,In_971,In_1686);
nor U3360 (N_3360,In_1356,In_1166);
and U3361 (N_3361,In_1350,In_429);
nand U3362 (N_3362,In_1945,In_1963);
nand U3363 (N_3363,In_1287,In_1479);
xor U3364 (N_3364,In_1723,In_1402);
nand U3365 (N_3365,In_1587,In_1721);
and U3366 (N_3366,In_1454,In_1039);
nor U3367 (N_3367,In_1068,In_447);
nor U3368 (N_3368,In_101,In_1001);
or U3369 (N_3369,In_483,In_1815);
nor U3370 (N_3370,In_292,In_211);
xor U3371 (N_3371,In_1090,In_156);
or U3372 (N_3372,In_704,In_218);
nand U3373 (N_3373,In_1989,In_1873);
nand U3374 (N_3374,In_154,In_255);
or U3375 (N_3375,In_1853,In_1335);
and U3376 (N_3376,In_1266,In_239);
or U3377 (N_3377,In_997,In_1108);
and U3378 (N_3378,In_1785,In_1212);
nand U3379 (N_3379,In_192,In_1560);
xor U3380 (N_3380,In_909,In_1204);
or U3381 (N_3381,In_35,In_1470);
nand U3382 (N_3382,In_595,In_1144);
nand U3383 (N_3383,In_263,In_371);
and U3384 (N_3384,In_1592,In_46);
nand U3385 (N_3385,In_111,In_132);
and U3386 (N_3386,In_1820,In_1182);
or U3387 (N_3387,In_724,In_1409);
nor U3388 (N_3388,In_1814,In_967);
and U3389 (N_3389,In_929,In_172);
and U3390 (N_3390,In_1654,In_1857);
or U3391 (N_3391,In_514,In_1062);
and U3392 (N_3392,In_1753,In_1233);
or U3393 (N_3393,In_230,In_1596);
or U3394 (N_3394,In_719,In_1556);
nand U3395 (N_3395,In_446,In_792);
nor U3396 (N_3396,In_138,In_873);
and U3397 (N_3397,In_177,In_50);
and U3398 (N_3398,In_849,In_1658);
and U3399 (N_3399,In_1796,In_1316);
nor U3400 (N_3400,In_126,In_598);
nor U3401 (N_3401,In_1922,In_1527);
nand U3402 (N_3402,In_473,In_1671);
and U3403 (N_3403,In_1237,In_1024);
nor U3404 (N_3404,In_452,In_421);
and U3405 (N_3405,In_467,In_1670);
nor U3406 (N_3406,In_44,In_949);
and U3407 (N_3407,In_990,In_820);
and U3408 (N_3408,In_550,In_1288);
nor U3409 (N_3409,In_279,In_820);
and U3410 (N_3410,In_1758,In_370);
nand U3411 (N_3411,In_1622,In_1701);
nor U3412 (N_3412,In_1488,In_674);
and U3413 (N_3413,In_1891,In_426);
or U3414 (N_3414,In_104,In_1229);
nand U3415 (N_3415,In_129,In_1929);
and U3416 (N_3416,In_154,In_445);
and U3417 (N_3417,In_207,In_1355);
nor U3418 (N_3418,In_1224,In_737);
nand U3419 (N_3419,In_1977,In_1772);
and U3420 (N_3420,In_218,In_338);
nor U3421 (N_3421,In_1103,In_164);
and U3422 (N_3422,In_676,In_590);
or U3423 (N_3423,In_1557,In_1707);
or U3424 (N_3424,In_1545,In_617);
nand U3425 (N_3425,In_793,In_1546);
nand U3426 (N_3426,In_52,In_818);
xor U3427 (N_3427,In_352,In_1509);
nand U3428 (N_3428,In_764,In_34);
or U3429 (N_3429,In_1103,In_573);
nor U3430 (N_3430,In_655,In_564);
and U3431 (N_3431,In_1206,In_834);
or U3432 (N_3432,In_718,In_771);
and U3433 (N_3433,In_238,In_127);
nand U3434 (N_3434,In_388,In_1956);
xnor U3435 (N_3435,In_1721,In_79);
nor U3436 (N_3436,In_1586,In_336);
nand U3437 (N_3437,In_1306,In_1381);
xnor U3438 (N_3438,In_526,In_843);
or U3439 (N_3439,In_639,In_1296);
and U3440 (N_3440,In_830,In_30);
and U3441 (N_3441,In_1466,In_1375);
nand U3442 (N_3442,In_691,In_251);
nand U3443 (N_3443,In_1354,In_735);
nand U3444 (N_3444,In_79,In_976);
or U3445 (N_3445,In_933,In_1209);
nand U3446 (N_3446,In_274,In_15);
and U3447 (N_3447,In_1468,In_1325);
nor U3448 (N_3448,In_784,In_295);
nand U3449 (N_3449,In_1815,In_1990);
or U3450 (N_3450,In_763,In_1842);
and U3451 (N_3451,In_1823,In_1186);
or U3452 (N_3452,In_1265,In_1007);
nand U3453 (N_3453,In_1011,In_1967);
and U3454 (N_3454,In_1636,In_365);
nor U3455 (N_3455,In_1306,In_1488);
or U3456 (N_3456,In_782,In_803);
and U3457 (N_3457,In_1113,In_22);
nand U3458 (N_3458,In_561,In_898);
and U3459 (N_3459,In_1394,In_1818);
or U3460 (N_3460,In_484,In_565);
and U3461 (N_3461,In_98,In_878);
nor U3462 (N_3462,In_748,In_1869);
and U3463 (N_3463,In_532,In_1237);
nand U3464 (N_3464,In_170,In_1702);
and U3465 (N_3465,In_442,In_217);
nor U3466 (N_3466,In_1897,In_1452);
nor U3467 (N_3467,In_1484,In_883);
and U3468 (N_3468,In_1367,In_391);
and U3469 (N_3469,In_1915,In_1844);
nor U3470 (N_3470,In_801,In_946);
nand U3471 (N_3471,In_674,In_1088);
nand U3472 (N_3472,In_1508,In_1479);
or U3473 (N_3473,In_1470,In_1945);
or U3474 (N_3474,In_1230,In_529);
nor U3475 (N_3475,In_114,In_1393);
or U3476 (N_3476,In_1539,In_1550);
nand U3477 (N_3477,In_927,In_1484);
nor U3478 (N_3478,In_1646,In_56);
and U3479 (N_3479,In_305,In_1258);
or U3480 (N_3480,In_1178,In_305);
nor U3481 (N_3481,In_1257,In_618);
and U3482 (N_3482,In_392,In_1715);
or U3483 (N_3483,In_165,In_1870);
and U3484 (N_3484,In_1951,In_1971);
nand U3485 (N_3485,In_486,In_511);
or U3486 (N_3486,In_1711,In_362);
and U3487 (N_3487,In_250,In_764);
nand U3488 (N_3488,In_1982,In_1778);
nor U3489 (N_3489,In_1396,In_1547);
nand U3490 (N_3490,In_993,In_1224);
nand U3491 (N_3491,In_919,In_1664);
and U3492 (N_3492,In_1587,In_268);
nand U3493 (N_3493,In_257,In_677);
nor U3494 (N_3494,In_102,In_1244);
and U3495 (N_3495,In_824,In_510);
or U3496 (N_3496,In_638,In_149);
nor U3497 (N_3497,In_1284,In_1583);
or U3498 (N_3498,In_643,In_488);
and U3499 (N_3499,In_468,In_1684);
or U3500 (N_3500,In_177,In_1195);
or U3501 (N_3501,In_1841,In_156);
nand U3502 (N_3502,In_1535,In_1235);
nor U3503 (N_3503,In_1052,In_1370);
or U3504 (N_3504,In_1579,In_172);
or U3505 (N_3505,In_912,In_409);
or U3506 (N_3506,In_1157,In_452);
or U3507 (N_3507,In_558,In_62);
and U3508 (N_3508,In_304,In_1203);
or U3509 (N_3509,In_507,In_1971);
or U3510 (N_3510,In_1512,In_946);
nor U3511 (N_3511,In_1605,In_1883);
and U3512 (N_3512,In_1928,In_1725);
and U3513 (N_3513,In_245,In_1226);
and U3514 (N_3514,In_528,In_1400);
nand U3515 (N_3515,In_1344,In_344);
and U3516 (N_3516,In_566,In_228);
nand U3517 (N_3517,In_27,In_951);
nand U3518 (N_3518,In_785,In_1753);
nor U3519 (N_3519,In_925,In_1918);
and U3520 (N_3520,In_332,In_1750);
nand U3521 (N_3521,In_1044,In_1766);
nand U3522 (N_3522,In_1094,In_512);
and U3523 (N_3523,In_797,In_1196);
nor U3524 (N_3524,In_1099,In_1188);
or U3525 (N_3525,In_650,In_1146);
or U3526 (N_3526,In_1215,In_564);
and U3527 (N_3527,In_1310,In_363);
and U3528 (N_3528,In_1660,In_258);
and U3529 (N_3529,In_1264,In_170);
nor U3530 (N_3530,In_987,In_657);
and U3531 (N_3531,In_1287,In_1247);
or U3532 (N_3532,In_1707,In_743);
and U3533 (N_3533,In_1689,In_307);
nand U3534 (N_3534,In_1914,In_1773);
or U3535 (N_3535,In_1438,In_39);
nor U3536 (N_3536,In_1916,In_573);
nor U3537 (N_3537,In_367,In_805);
nand U3538 (N_3538,In_1285,In_569);
nand U3539 (N_3539,In_444,In_206);
or U3540 (N_3540,In_1788,In_1989);
or U3541 (N_3541,In_777,In_882);
nor U3542 (N_3542,In_126,In_775);
and U3543 (N_3543,In_685,In_1994);
nor U3544 (N_3544,In_286,In_1081);
nor U3545 (N_3545,In_1106,In_1484);
nand U3546 (N_3546,In_770,In_679);
nand U3547 (N_3547,In_1353,In_302);
or U3548 (N_3548,In_1591,In_258);
nor U3549 (N_3549,In_1017,In_1962);
nand U3550 (N_3550,In_812,In_1308);
or U3551 (N_3551,In_667,In_1429);
and U3552 (N_3552,In_1948,In_1350);
nor U3553 (N_3553,In_1274,In_1708);
nand U3554 (N_3554,In_574,In_1167);
nand U3555 (N_3555,In_380,In_331);
nand U3556 (N_3556,In_298,In_1808);
nand U3557 (N_3557,In_1103,In_578);
and U3558 (N_3558,In_1884,In_1045);
nor U3559 (N_3559,In_1749,In_1387);
nand U3560 (N_3560,In_1593,In_910);
and U3561 (N_3561,In_1628,In_1185);
nand U3562 (N_3562,In_1537,In_1459);
or U3563 (N_3563,In_815,In_635);
nor U3564 (N_3564,In_1947,In_1170);
nand U3565 (N_3565,In_1198,In_1863);
nand U3566 (N_3566,In_291,In_295);
and U3567 (N_3567,In_302,In_155);
and U3568 (N_3568,In_1123,In_1789);
and U3569 (N_3569,In_892,In_725);
nor U3570 (N_3570,In_1824,In_1135);
nor U3571 (N_3571,In_1177,In_1219);
nor U3572 (N_3572,In_1734,In_776);
or U3573 (N_3573,In_1090,In_113);
and U3574 (N_3574,In_1885,In_1452);
nor U3575 (N_3575,In_1738,In_593);
nand U3576 (N_3576,In_1264,In_895);
nand U3577 (N_3577,In_917,In_1469);
nor U3578 (N_3578,In_1824,In_1597);
nor U3579 (N_3579,In_284,In_395);
nor U3580 (N_3580,In_1723,In_69);
and U3581 (N_3581,In_1467,In_778);
nand U3582 (N_3582,In_329,In_269);
nor U3583 (N_3583,In_1878,In_1302);
and U3584 (N_3584,In_979,In_602);
or U3585 (N_3585,In_1635,In_1549);
nand U3586 (N_3586,In_309,In_228);
nand U3587 (N_3587,In_791,In_818);
and U3588 (N_3588,In_1407,In_4);
nor U3589 (N_3589,In_1340,In_734);
nand U3590 (N_3590,In_517,In_606);
nand U3591 (N_3591,In_1436,In_987);
nand U3592 (N_3592,In_848,In_1986);
nor U3593 (N_3593,In_322,In_1564);
and U3594 (N_3594,In_444,In_1901);
and U3595 (N_3595,In_1112,In_1795);
nand U3596 (N_3596,In_1345,In_906);
nand U3597 (N_3597,In_1627,In_1118);
and U3598 (N_3598,In_1530,In_271);
nor U3599 (N_3599,In_1467,In_120);
and U3600 (N_3600,In_1688,In_1098);
nand U3601 (N_3601,In_42,In_1471);
nand U3602 (N_3602,In_1090,In_453);
or U3603 (N_3603,In_347,In_1137);
or U3604 (N_3604,In_562,In_1704);
nand U3605 (N_3605,In_672,In_860);
and U3606 (N_3606,In_461,In_1207);
nor U3607 (N_3607,In_1146,In_1580);
nor U3608 (N_3608,In_1397,In_1528);
and U3609 (N_3609,In_1390,In_1997);
nor U3610 (N_3610,In_1346,In_1794);
nand U3611 (N_3611,In_933,In_744);
or U3612 (N_3612,In_64,In_1216);
and U3613 (N_3613,In_1095,In_850);
and U3614 (N_3614,In_1158,In_1026);
nor U3615 (N_3615,In_1572,In_478);
or U3616 (N_3616,In_323,In_1775);
and U3617 (N_3617,In_571,In_76);
nand U3618 (N_3618,In_902,In_838);
nor U3619 (N_3619,In_1332,In_1209);
nand U3620 (N_3620,In_701,In_1527);
nand U3621 (N_3621,In_725,In_658);
nand U3622 (N_3622,In_1247,In_1932);
nand U3623 (N_3623,In_718,In_1640);
and U3624 (N_3624,In_1431,In_1850);
nor U3625 (N_3625,In_1302,In_418);
nand U3626 (N_3626,In_1384,In_1125);
xor U3627 (N_3627,In_1047,In_928);
nor U3628 (N_3628,In_1466,In_461);
or U3629 (N_3629,In_495,In_620);
nor U3630 (N_3630,In_412,In_1338);
and U3631 (N_3631,In_753,In_469);
nand U3632 (N_3632,In_481,In_83);
and U3633 (N_3633,In_1425,In_1019);
nor U3634 (N_3634,In_1514,In_648);
nor U3635 (N_3635,In_522,In_27);
or U3636 (N_3636,In_1606,In_1618);
or U3637 (N_3637,In_146,In_279);
and U3638 (N_3638,In_30,In_1326);
nand U3639 (N_3639,In_1815,In_990);
and U3640 (N_3640,In_797,In_2);
nor U3641 (N_3641,In_1104,In_656);
nand U3642 (N_3642,In_166,In_1034);
nor U3643 (N_3643,In_1830,In_1463);
nor U3644 (N_3644,In_1214,In_1775);
or U3645 (N_3645,In_525,In_1956);
nand U3646 (N_3646,In_1932,In_1906);
nor U3647 (N_3647,In_808,In_1181);
nor U3648 (N_3648,In_230,In_734);
nand U3649 (N_3649,In_1237,In_1300);
nor U3650 (N_3650,In_1229,In_1070);
nand U3651 (N_3651,In_355,In_1746);
nand U3652 (N_3652,In_1222,In_1433);
nand U3653 (N_3653,In_1508,In_116);
or U3654 (N_3654,In_545,In_1613);
nand U3655 (N_3655,In_1468,In_1007);
nor U3656 (N_3656,In_736,In_1934);
and U3657 (N_3657,In_732,In_284);
or U3658 (N_3658,In_1067,In_1734);
and U3659 (N_3659,In_1586,In_1708);
nand U3660 (N_3660,In_1844,In_1609);
and U3661 (N_3661,In_407,In_428);
and U3662 (N_3662,In_192,In_1014);
nand U3663 (N_3663,In_1826,In_1197);
nor U3664 (N_3664,In_1380,In_223);
nand U3665 (N_3665,In_258,In_1075);
and U3666 (N_3666,In_1489,In_57);
and U3667 (N_3667,In_346,In_1805);
and U3668 (N_3668,In_131,In_656);
nand U3669 (N_3669,In_691,In_1023);
and U3670 (N_3670,In_135,In_1419);
nor U3671 (N_3671,In_1504,In_1010);
and U3672 (N_3672,In_119,In_1493);
and U3673 (N_3673,In_758,In_1573);
nor U3674 (N_3674,In_412,In_439);
nor U3675 (N_3675,In_351,In_1916);
xnor U3676 (N_3676,In_1879,In_185);
and U3677 (N_3677,In_880,In_335);
nand U3678 (N_3678,In_1700,In_1620);
or U3679 (N_3679,In_1857,In_1553);
or U3680 (N_3680,In_1587,In_352);
and U3681 (N_3681,In_409,In_1310);
or U3682 (N_3682,In_820,In_255);
nand U3683 (N_3683,In_1755,In_651);
and U3684 (N_3684,In_1438,In_1765);
and U3685 (N_3685,In_800,In_944);
nor U3686 (N_3686,In_1919,In_1735);
or U3687 (N_3687,In_175,In_1472);
or U3688 (N_3688,In_271,In_1533);
nand U3689 (N_3689,In_419,In_25);
nor U3690 (N_3690,In_51,In_494);
nor U3691 (N_3691,In_14,In_609);
nor U3692 (N_3692,In_23,In_461);
nand U3693 (N_3693,In_1992,In_1386);
and U3694 (N_3694,In_663,In_648);
or U3695 (N_3695,In_1593,In_1598);
nand U3696 (N_3696,In_1031,In_755);
or U3697 (N_3697,In_1444,In_55);
and U3698 (N_3698,In_815,In_939);
nor U3699 (N_3699,In_824,In_525);
or U3700 (N_3700,In_1627,In_1102);
and U3701 (N_3701,In_1870,In_1665);
nand U3702 (N_3702,In_501,In_1263);
nor U3703 (N_3703,In_922,In_1796);
and U3704 (N_3704,In_1666,In_1933);
nand U3705 (N_3705,In_1036,In_797);
and U3706 (N_3706,In_494,In_97);
nor U3707 (N_3707,In_1560,In_825);
nor U3708 (N_3708,In_985,In_64);
or U3709 (N_3709,In_1008,In_1269);
or U3710 (N_3710,In_734,In_1813);
or U3711 (N_3711,In_310,In_1866);
nand U3712 (N_3712,In_1601,In_1351);
or U3713 (N_3713,In_585,In_448);
nand U3714 (N_3714,In_1319,In_434);
or U3715 (N_3715,In_1883,In_1187);
or U3716 (N_3716,In_686,In_1380);
and U3717 (N_3717,In_212,In_604);
or U3718 (N_3718,In_402,In_1675);
nand U3719 (N_3719,In_1014,In_831);
nand U3720 (N_3720,In_1712,In_710);
nand U3721 (N_3721,In_1952,In_460);
nor U3722 (N_3722,In_845,In_1315);
nor U3723 (N_3723,In_1470,In_1216);
and U3724 (N_3724,In_71,In_573);
nor U3725 (N_3725,In_1971,In_1154);
nor U3726 (N_3726,In_932,In_676);
nand U3727 (N_3727,In_440,In_723);
and U3728 (N_3728,In_627,In_712);
and U3729 (N_3729,In_1199,In_136);
nand U3730 (N_3730,In_79,In_458);
nand U3731 (N_3731,In_1496,In_607);
nand U3732 (N_3732,In_124,In_812);
or U3733 (N_3733,In_187,In_1304);
xnor U3734 (N_3734,In_400,In_1094);
and U3735 (N_3735,In_1204,In_1901);
nand U3736 (N_3736,In_1938,In_1466);
and U3737 (N_3737,In_99,In_1228);
nor U3738 (N_3738,In_440,In_92);
nor U3739 (N_3739,In_1580,In_17);
or U3740 (N_3740,In_1474,In_1212);
nor U3741 (N_3741,In_461,In_729);
nor U3742 (N_3742,In_1992,In_1525);
nand U3743 (N_3743,In_485,In_1456);
and U3744 (N_3744,In_1719,In_928);
nand U3745 (N_3745,In_1569,In_296);
nand U3746 (N_3746,In_590,In_1721);
or U3747 (N_3747,In_1477,In_1739);
and U3748 (N_3748,In_624,In_596);
nand U3749 (N_3749,In_1179,In_1574);
or U3750 (N_3750,In_843,In_250);
and U3751 (N_3751,In_1724,In_768);
or U3752 (N_3752,In_1677,In_1864);
nor U3753 (N_3753,In_377,In_620);
and U3754 (N_3754,In_1273,In_222);
and U3755 (N_3755,In_1514,In_351);
and U3756 (N_3756,In_1350,In_315);
nor U3757 (N_3757,In_1813,In_1602);
nand U3758 (N_3758,In_1333,In_955);
and U3759 (N_3759,In_1814,In_1253);
nor U3760 (N_3760,In_1919,In_1125);
or U3761 (N_3761,In_1048,In_36);
or U3762 (N_3762,In_858,In_1817);
nor U3763 (N_3763,In_160,In_1399);
and U3764 (N_3764,In_1818,In_900);
nor U3765 (N_3765,In_1472,In_1707);
or U3766 (N_3766,In_315,In_820);
or U3767 (N_3767,In_1268,In_845);
or U3768 (N_3768,In_983,In_498);
nand U3769 (N_3769,In_1655,In_1688);
nor U3770 (N_3770,In_496,In_1016);
or U3771 (N_3771,In_1384,In_631);
nand U3772 (N_3772,In_1604,In_571);
nor U3773 (N_3773,In_773,In_1488);
and U3774 (N_3774,In_874,In_582);
or U3775 (N_3775,In_1285,In_1081);
nor U3776 (N_3776,In_1016,In_105);
nand U3777 (N_3777,In_1481,In_918);
nor U3778 (N_3778,In_1795,In_910);
or U3779 (N_3779,In_991,In_1884);
nor U3780 (N_3780,In_1742,In_394);
nand U3781 (N_3781,In_585,In_1380);
nor U3782 (N_3782,In_425,In_1951);
nor U3783 (N_3783,In_1436,In_941);
nor U3784 (N_3784,In_1588,In_1340);
or U3785 (N_3785,In_1326,In_1392);
and U3786 (N_3786,In_112,In_1433);
and U3787 (N_3787,In_777,In_1426);
nand U3788 (N_3788,In_49,In_334);
nand U3789 (N_3789,In_1774,In_1176);
nor U3790 (N_3790,In_1795,In_1733);
and U3791 (N_3791,In_831,In_1050);
or U3792 (N_3792,In_1846,In_762);
xnor U3793 (N_3793,In_633,In_519);
nand U3794 (N_3794,In_599,In_1642);
nand U3795 (N_3795,In_505,In_1176);
and U3796 (N_3796,In_7,In_120);
nand U3797 (N_3797,In_1021,In_1068);
and U3798 (N_3798,In_1401,In_1302);
or U3799 (N_3799,In_1396,In_45);
or U3800 (N_3800,In_1703,In_803);
or U3801 (N_3801,In_404,In_610);
nand U3802 (N_3802,In_595,In_1622);
or U3803 (N_3803,In_694,In_540);
or U3804 (N_3804,In_7,In_153);
nor U3805 (N_3805,In_453,In_933);
nand U3806 (N_3806,In_585,In_1664);
nand U3807 (N_3807,In_557,In_502);
nand U3808 (N_3808,In_1803,In_629);
and U3809 (N_3809,In_1901,In_1825);
nor U3810 (N_3810,In_91,In_1801);
nand U3811 (N_3811,In_480,In_116);
or U3812 (N_3812,In_1531,In_1154);
or U3813 (N_3813,In_1961,In_1860);
or U3814 (N_3814,In_1007,In_1871);
nor U3815 (N_3815,In_1588,In_1902);
or U3816 (N_3816,In_641,In_635);
nand U3817 (N_3817,In_248,In_1294);
nor U3818 (N_3818,In_776,In_123);
and U3819 (N_3819,In_1156,In_1390);
nor U3820 (N_3820,In_794,In_1293);
nand U3821 (N_3821,In_822,In_1214);
nor U3822 (N_3822,In_207,In_1069);
and U3823 (N_3823,In_641,In_1831);
and U3824 (N_3824,In_528,In_302);
nand U3825 (N_3825,In_408,In_479);
or U3826 (N_3826,In_1333,In_85);
or U3827 (N_3827,In_42,In_889);
nor U3828 (N_3828,In_1037,In_1501);
or U3829 (N_3829,In_397,In_420);
or U3830 (N_3830,In_1396,In_1035);
nand U3831 (N_3831,In_1745,In_1729);
or U3832 (N_3832,In_660,In_526);
nand U3833 (N_3833,In_1942,In_1718);
and U3834 (N_3834,In_513,In_1189);
and U3835 (N_3835,In_1999,In_880);
or U3836 (N_3836,In_1109,In_1478);
or U3837 (N_3837,In_1590,In_1639);
and U3838 (N_3838,In_1376,In_1351);
nand U3839 (N_3839,In_1973,In_1085);
and U3840 (N_3840,In_1040,In_688);
nor U3841 (N_3841,In_1980,In_1688);
nand U3842 (N_3842,In_775,In_22);
or U3843 (N_3843,In_445,In_134);
nand U3844 (N_3844,In_1592,In_717);
and U3845 (N_3845,In_765,In_1720);
nand U3846 (N_3846,In_1933,In_1885);
nor U3847 (N_3847,In_1785,In_1546);
and U3848 (N_3848,In_986,In_1140);
and U3849 (N_3849,In_1366,In_1798);
or U3850 (N_3850,In_1466,In_1996);
nor U3851 (N_3851,In_315,In_1338);
nor U3852 (N_3852,In_247,In_1311);
or U3853 (N_3853,In_1176,In_389);
nor U3854 (N_3854,In_1213,In_454);
and U3855 (N_3855,In_320,In_801);
or U3856 (N_3856,In_317,In_902);
nor U3857 (N_3857,In_1227,In_725);
nand U3858 (N_3858,In_1504,In_1832);
nor U3859 (N_3859,In_1972,In_463);
or U3860 (N_3860,In_1766,In_464);
nand U3861 (N_3861,In_902,In_1171);
and U3862 (N_3862,In_24,In_529);
and U3863 (N_3863,In_1829,In_329);
and U3864 (N_3864,In_1134,In_1133);
or U3865 (N_3865,In_521,In_576);
or U3866 (N_3866,In_199,In_623);
and U3867 (N_3867,In_224,In_1916);
xnor U3868 (N_3868,In_808,In_826);
or U3869 (N_3869,In_647,In_1728);
nand U3870 (N_3870,In_411,In_1316);
or U3871 (N_3871,In_1719,In_57);
nand U3872 (N_3872,In_713,In_227);
nor U3873 (N_3873,In_990,In_267);
nor U3874 (N_3874,In_497,In_366);
nand U3875 (N_3875,In_418,In_1611);
nor U3876 (N_3876,In_909,In_209);
or U3877 (N_3877,In_683,In_708);
nor U3878 (N_3878,In_701,In_917);
nand U3879 (N_3879,In_997,In_580);
or U3880 (N_3880,In_1692,In_998);
or U3881 (N_3881,In_1386,In_508);
nor U3882 (N_3882,In_1891,In_1890);
nand U3883 (N_3883,In_1889,In_1170);
nor U3884 (N_3884,In_119,In_967);
and U3885 (N_3885,In_17,In_1029);
nor U3886 (N_3886,In_1158,In_1393);
nor U3887 (N_3887,In_1088,In_930);
nor U3888 (N_3888,In_1229,In_1979);
xnor U3889 (N_3889,In_1141,In_1759);
and U3890 (N_3890,In_779,In_940);
or U3891 (N_3891,In_996,In_216);
nand U3892 (N_3892,In_1086,In_391);
nor U3893 (N_3893,In_1766,In_1675);
nor U3894 (N_3894,In_126,In_53);
and U3895 (N_3895,In_1013,In_184);
or U3896 (N_3896,In_1609,In_1648);
nand U3897 (N_3897,In_1693,In_1408);
and U3898 (N_3898,In_251,In_1296);
nor U3899 (N_3899,In_148,In_1744);
nand U3900 (N_3900,In_915,In_290);
and U3901 (N_3901,In_215,In_1785);
xor U3902 (N_3902,In_851,In_1132);
and U3903 (N_3903,In_1169,In_1917);
or U3904 (N_3904,In_479,In_817);
or U3905 (N_3905,In_208,In_1759);
nor U3906 (N_3906,In_277,In_757);
nor U3907 (N_3907,In_1594,In_797);
or U3908 (N_3908,In_726,In_230);
nand U3909 (N_3909,In_948,In_1359);
and U3910 (N_3910,In_292,In_665);
and U3911 (N_3911,In_1625,In_324);
nor U3912 (N_3912,In_1645,In_1397);
nand U3913 (N_3913,In_388,In_227);
xor U3914 (N_3914,In_93,In_1669);
nor U3915 (N_3915,In_1729,In_870);
or U3916 (N_3916,In_780,In_622);
nand U3917 (N_3917,In_1782,In_1466);
nand U3918 (N_3918,In_1966,In_858);
nand U3919 (N_3919,In_788,In_1713);
nor U3920 (N_3920,In_1008,In_1560);
nand U3921 (N_3921,In_1459,In_1051);
nor U3922 (N_3922,In_1296,In_372);
nand U3923 (N_3923,In_958,In_388);
and U3924 (N_3924,In_529,In_61);
and U3925 (N_3925,In_932,In_904);
nand U3926 (N_3926,In_1380,In_524);
nor U3927 (N_3927,In_727,In_234);
nor U3928 (N_3928,In_451,In_659);
or U3929 (N_3929,In_290,In_374);
nand U3930 (N_3930,In_812,In_854);
nor U3931 (N_3931,In_143,In_866);
nand U3932 (N_3932,In_1818,In_1331);
nor U3933 (N_3933,In_431,In_1251);
or U3934 (N_3934,In_1635,In_1170);
nand U3935 (N_3935,In_921,In_531);
xor U3936 (N_3936,In_1751,In_1047);
or U3937 (N_3937,In_926,In_180);
and U3938 (N_3938,In_335,In_437);
nor U3939 (N_3939,In_1630,In_1126);
and U3940 (N_3940,In_1945,In_1884);
nand U3941 (N_3941,In_496,In_1411);
and U3942 (N_3942,In_963,In_1379);
and U3943 (N_3943,In_1148,In_542);
and U3944 (N_3944,In_1549,In_895);
nand U3945 (N_3945,In_319,In_75);
nor U3946 (N_3946,In_1786,In_354);
nand U3947 (N_3947,In_1792,In_1793);
or U3948 (N_3948,In_1708,In_1311);
xor U3949 (N_3949,In_1778,In_1269);
nor U3950 (N_3950,In_1324,In_1239);
and U3951 (N_3951,In_1376,In_818);
nor U3952 (N_3952,In_809,In_730);
nor U3953 (N_3953,In_1650,In_386);
nand U3954 (N_3954,In_513,In_1418);
nor U3955 (N_3955,In_1177,In_1133);
nand U3956 (N_3956,In_1052,In_627);
or U3957 (N_3957,In_1403,In_853);
nand U3958 (N_3958,In_1403,In_1248);
and U3959 (N_3959,In_1329,In_331);
and U3960 (N_3960,In_518,In_757);
and U3961 (N_3961,In_1657,In_65);
or U3962 (N_3962,In_1647,In_985);
and U3963 (N_3963,In_1989,In_1378);
and U3964 (N_3964,In_472,In_803);
or U3965 (N_3965,In_187,In_893);
and U3966 (N_3966,In_471,In_1203);
nand U3967 (N_3967,In_898,In_1333);
and U3968 (N_3968,In_1302,In_77);
nor U3969 (N_3969,In_772,In_234);
xnor U3970 (N_3970,In_1182,In_1645);
nor U3971 (N_3971,In_1512,In_1083);
nor U3972 (N_3972,In_124,In_136);
nor U3973 (N_3973,In_442,In_780);
and U3974 (N_3974,In_1144,In_1072);
and U3975 (N_3975,In_1213,In_491);
and U3976 (N_3976,In_204,In_542);
nor U3977 (N_3977,In_1485,In_1688);
nor U3978 (N_3978,In_1494,In_1689);
and U3979 (N_3979,In_981,In_310);
nor U3980 (N_3980,In_1642,In_488);
nand U3981 (N_3981,In_776,In_1875);
and U3982 (N_3982,In_876,In_1906);
nor U3983 (N_3983,In_1679,In_1510);
nand U3984 (N_3984,In_1712,In_1635);
nand U3985 (N_3985,In_1871,In_1442);
and U3986 (N_3986,In_814,In_1740);
nor U3987 (N_3987,In_73,In_1276);
or U3988 (N_3988,In_644,In_1304);
nand U3989 (N_3989,In_808,In_676);
or U3990 (N_3990,In_979,In_121);
nand U3991 (N_3991,In_325,In_12);
or U3992 (N_3992,In_1379,In_1302);
nor U3993 (N_3993,In_1406,In_475);
or U3994 (N_3994,In_510,In_90);
or U3995 (N_3995,In_1758,In_831);
and U3996 (N_3996,In_508,In_1490);
nand U3997 (N_3997,In_1481,In_231);
and U3998 (N_3998,In_1394,In_1009);
and U3999 (N_3999,In_320,In_1532);
nand U4000 (N_4000,In_240,In_112);
or U4001 (N_4001,In_183,In_681);
nand U4002 (N_4002,In_1080,In_839);
and U4003 (N_4003,In_874,In_187);
and U4004 (N_4004,In_1439,In_615);
nand U4005 (N_4005,In_728,In_72);
nand U4006 (N_4006,In_1913,In_976);
nor U4007 (N_4007,In_658,In_1140);
nor U4008 (N_4008,In_292,In_1745);
and U4009 (N_4009,In_1296,In_802);
nand U4010 (N_4010,In_1194,In_333);
nand U4011 (N_4011,In_1741,In_1643);
and U4012 (N_4012,In_749,In_1923);
and U4013 (N_4013,In_1976,In_495);
or U4014 (N_4014,In_1291,In_431);
nor U4015 (N_4015,In_1660,In_237);
or U4016 (N_4016,In_211,In_441);
nand U4017 (N_4017,In_144,In_872);
or U4018 (N_4018,In_1050,In_1652);
nor U4019 (N_4019,In_22,In_437);
nor U4020 (N_4020,In_1347,In_1644);
nor U4021 (N_4021,In_648,In_1511);
nor U4022 (N_4022,In_1585,In_1539);
nor U4023 (N_4023,In_1512,In_1938);
nand U4024 (N_4024,In_428,In_692);
nor U4025 (N_4025,In_878,In_1439);
or U4026 (N_4026,In_906,In_1643);
and U4027 (N_4027,In_1821,In_1436);
nor U4028 (N_4028,In_1920,In_1590);
or U4029 (N_4029,In_1366,In_711);
nor U4030 (N_4030,In_879,In_1133);
nand U4031 (N_4031,In_1544,In_1240);
nand U4032 (N_4032,In_1152,In_1094);
or U4033 (N_4033,In_1020,In_983);
nor U4034 (N_4034,In_1904,In_1638);
nor U4035 (N_4035,In_1154,In_1331);
or U4036 (N_4036,In_1141,In_465);
nor U4037 (N_4037,In_926,In_920);
nand U4038 (N_4038,In_31,In_1627);
or U4039 (N_4039,In_1936,In_1354);
and U4040 (N_4040,In_1952,In_1532);
and U4041 (N_4041,In_1986,In_1419);
or U4042 (N_4042,In_1890,In_847);
nand U4043 (N_4043,In_943,In_57);
and U4044 (N_4044,In_174,In_67);
nand U4045 (N_4045,In_996,In_1016);
nand U4046 (N_4046,In_712,In_1609);
or U4047 (N_4047,In_1232,In_632);
or U4048 (N_4048,In_500,In_224);
and U4049 (N_4049,In_1721,In_826);
and U4050 (N_4050,In_194,In_305);
and U4051 (N_4051,In_804,In_1652);
and U4052 (N_4052,In_1413,In_228);
and U4053 (N_4053,In_1030,In_1770);
and U4054 (N_4054,In_1049,In_1726);
and U4055 (N_4055,In_333,In_238);
and U4056 (N_4056,In_224,In_1147);
nor U4057 (N_4057,In_466,In_744);
and U4058 (N_4058,In_1421,In_911);
or U4059 (N_4059,In_426,In_1718);
and U4060 (N_4060,In_609,In_1494);
nor U4061 (N_4061,In_1602,In_198);
or U4062 (N_4062,In_1109,In_1960);
and U4063 (N_4063,In_962,In_1403);
and U4064 (N_4064,In_638,In_1702);
and U4065 (N_4065,In_534,In_1327);
nand U4066 (N_4066,In_598,In_1792);
and U4067 (N_4067,In_1125,In_247);
nor U4068 (N_4068,In_405,In_253);
and U4069 (N_4069,In_1544,In_59);
xor U4070 (N_4070,In_79,In_1240);
and U4071 (N_4071,In_1668,In_825);
nand U4072 (N_4072,In_436,In_282);
or U4073 (N_4073,In_573,In_1576);
nand U4074 (N_4074,In_575,In_1788);
or U4075 (N_4075,In_655,In_1926);
and U4076 (N_4076,In_1938,In_709);
and U4077 (N_4077,In_1200,In_605);
nand U4078 (N_4078,In_1226,In_36);
nor U4079 (N_4079,In_509,In_948);
nand U4080 (N_4080,In_489,In_983);
and U4081 (N_4081,In_1271,In_1998);
nor U4082 (N_4082,In_1426,In_1676);
and U4083 (N_4083,In_705,In_701);
and U4084 (N_4084,In_1732,In_593);
nand U4085 (N_4085,In_1075,In_204);
nand U4086 (N_4086,In_552,In_1557);
and U4087 (N_4087,In_1078,In_961);
or U4088 (N_4088,In_1864,In_1780);
nor U4089 (N_4089,In_1987,In_1637);
or U4090 (N_4090,In_1932,In_1801);
or U4091 (N_4091,In_88,In_416);
nor U4092 (N_4092,In_1345,In_1118);
and U4093 (N_4093,In_1034,In_990);
nor U4094 (N_4094,In_1074,In_444);
and U4095 (N_4095,In_633,In_1576);
or U4096 (N_4096,In_1214,In_902);
nand U4097 (N_4097,In_1284,In_240);
or U4098 (N_4098,In_646,In_1443);
and U4099 (N_4099,In_848,In_488);
or U4100 (N_4100,In_1942,In_1193);
or U4101 (N_4101,In_647,In_1867);
or U4102 (N_4102,In_755,In_176);
nand U4103 (N_4103,In_660,In_1767);
nand U4104 (N_4104,In_676,In_1065);
nor U4105 (N_4105,In_1670,In_1248);
nor U4106 (N_4106,In_1522,In_223);
or U4107 (N_4107,In_1694,In_1577);
nor U4108 (N_4108,In_101,In_589);
or U4109 (N_4109,In_1353,In_932);
or U4110 (N_4110,In_552,In_1588);
nand U4111 (N_4111,In_1235,In_76);
nor U4112 (N_4112,In_1972,In_229);
nand U4113 (N_4113,In_828,In_1679);
and U4114 (N_4114,In_1989,In_290);
nand U4115 (N_4115,In_946,In_818);
nor U4116 (N_4116,In_135,In_74);
and U4117 (N_4117,In_1020,In_1375);
nand U4118 (N_4118,In_1123,In_1319);
or U4119 (N_4119,In_1804,In_701);
nand U4120 (N_4120,In_265,In_780);
or U4121 (N_4121,In_994,In_877);
nand U4122 (N_4122,In_36,In_1800);
or U4123 (N_4123,In_918,In_1474);
or U4124 (N_4124,In_422,In_255);
nor U4125 (N_4125,In_1149,In_1184);
nor U4126 (N_4126,In_66,In_1990);
xnor U4127 (N_4127,In_957,In_1614);
or U4128 (N_4128,In_1602,In_1774);
or U4129 (N_4129,In_1085,In_1856);
nor U4130 (N_4130,In_158,In_1125);
and U4131 (N_4131,In_1658,In_1495);
nor U4132 (N_4132,In_248,In_1048);
nor U4133 (N_4133,In_717,In_1260);
nand U4134 (N_4134,In_610,In_212);
nand U4135 (N_4135,In_1449,In_707);
or U4136 (N_4136,In_573,In_584);
and U4137 (N_4137,In_151,In_1284);
nand U4138 (N_4138,In_344,In_463);
or U4139 (N_4139,In_1540,In_1071);
nor U4140 (N_4140,In_1875,In_1134);
and U4141 (N_4141,In_242,In_90);
or U4142 (N_4142,In_1639,In_1487);
nor U4143 (N_4143,In_959,In_248);
nand U4144 (N_4144,In_1601,In_1874);
and U4145 (N_4145,In_236,In_1353);
nor U4146 (N_4146,In_1732,In_1133);
or U4147 (N_4147,In_659,In_1754);
nor U4148 (N_4148,In_676,In_389);
nor U4149 (N_4149,In_1316,In_1632);
and U4150 (N_4150,In_1536,In_336);
nor U4151 (N_4151,In_1837,In_498);
or U4152 (N_4152,In_1818,In_1737);
or U4153 (N_4153,In_1233,In_1578);
or U4154 (N_4154,In_628,In_538);
nor U4155 (N_4155,In_1346,In_1014);
and U4156 (N_4156,In_1687,In_303);
and U4157 (N_4157,In_1629,In_1757);
nor U4158 (N_4158,In_1655,In_1854);
nor U4159 (N_4159,In_1754,In_1334);
and U4160 (N_4160,In_103,In_1621);
and U4161 (N_4161,In_1479,In_1756);
nand U4162 (N_4162,In_351,In_1445);
and U4163 (N_4163,In_618,In_277);
nor U4164 (N_4164,In_240,In_1887);
nor U4165 (N_4165,In_714,In_1450);
and U4166 (N_4166,In_1218,In_1195);
and U4167 (N_4167,In_965,In_694);
nor U4168 (N_4168,In_1229,In_753);
and U4169 (N_4169,In_894,In_163);
or U4170 (N_4170,In_534,In_1359);
xnor U4171 (N_4171,In_376,In_1604);
nor U4172 (N_4172,In_1807,In_1022);
nand U4173 (N_4173,In_1439,In_932);
or U4174 (N_4174,In_1911,In_1221);
nor U4175 (N_4175,In_234,In_1421);
nor U4176 (N_4176,In_1987,In_743);
nand U4177 (N_4177,In_650,In_954);
and U4178 (N_4178,In_1641,In_1805);
nand U4179 (N_4179,In_802,In_727);
nor U4180 (N_4180,In_803,In_161);
nor U4181 (N_4181,In_234,In_1794);
and U4182 (N_4182,In_787,In_993);
nor U4183 (N_4183,In_1320,In_1504);
nand U4184 (N_4184,In_698,In_534);
nand U4185 (N_4185,In_705,In_1426);
nand U4186 (N_4186,In_6,In_1387);
and U4187 (N_4187,In_306,In_1996);
nor U4188 (N_4188,In_1183,In_480);
nor U4189 (N_4189,In_1877,In_1453);
or U4190 (N_4190,In_1612,In_1322);
nor U4191 (N_4191,In_187,In_1539);
nor U4192 (N_4192,In_1033,In_667);
and U4193 (N_4193,In_527,In_631);
nor U4194 (N_4194,In_1163,In_1702);
or U4195 (N_4195,In_1633,In_1360);
nor U4196 (N_4196,In_898,In_574);
and U4197 (N_4197,In_1577,In_1278);
xnor U4198 (N_4198,In_275,In_1426);
nor U4199 (N_4199,In_950,In_38);
or U4200 (N_4200,In_1816,In_344);
nand U4201 (N_4201,In_1282,In_734);
and U4202 (N_4202,In_831,In_1824);
xnor U4203 (N_4203,In_369,In_173);
nand U4204 (N_4204,In_144,In_207);
and U4205 (N_4205,In_934,In_974);
xor U4206 (N_4206,In_1559,In_919);
or U4207 (N_4207,In_1250,In_1728);
nand U4208 (N_4208,In_1889,In_273);
or U4209 (N_4209,In_1842,In_567);
nor U4210 (N_4210,In_404,In_1748);
or U4211 (N_4211,In_1085,In_1299);
or U4212 (N_4212,In_745,In_671);
or U4213 (N_4213,In_857,In_106);
nor U4214 (N_4214,In_1289,In_827);
nand U4215 (N_4215,In_779,In_1452);
or U4216 (N_4216,In_1359,In_1591);
and U4217 (N_4217,In_1792,In_331);
or U4218 (N_4218,In_1513,In_1464);
nor U4219 (N_4219,In_382,In_1057);
and U4220 (N_4220,In_853,In_1700);
and U4221 (N_4221,In_1830,In_1032);
nor U4222 (N_4222,In_1277,In_1112);
nand U4223 (N_4223,In_1275,In_14);
and U4224 (N_4224,In_1337,In_1528);
or U4225 (N_4225,In_142,In_1990);
or U4226 (N_4226,In_105,In_1335);
nand U4227 (N_4227,In_1473,In_904);
nand U4228 (N_4228,In_147,In_265);
nor U4229 (N_4229,In_1046,In_1081);
nand U4230 (N_4230,In_272,In_1187);
xnor U4231 (N_4231,In_1316,In_1941);
or U4232 (N_4232,In_1214,In_504);
and U4233 (N_4233,In_1326,In_576);
or U4234 (N_4234,In_1309,In_605);
or U4235 (N_4235,In_312,In_1823);
or U4236 (N_4236,In_87,In_1222);
nor U4237 (N_4237,In_422,In_1486);
and U4238 (N_4238,In_1037,In_772);
nand U4239 (N_4239,In_484,In_712);
and U4240 (N_4240,In_1201,In_410);
nor U4241 (N_4241,In_702,In_169);
or U4242 (N_4242,In_367,In_1067);
and U4243 (N_4243,In_521,In_531);
or U4244 (N_4244,In_868,In_8);
nor U4245 (N_4245,In_146,In_1593);
nand U4246 (N_4246,In_1172,In_708);
or U4247 (N_4247,In_1703,In_169);
and U4248 (N_4248,In_1278,In_1033);
nor U4249 (N_4249,In_1963,In_967);
nor U4250 (N_4250,In_1007,In_221);
nor U4251 (N_4251,In_455,In_1025);
nand U4252 (N_4252,In_1556,In_860);
nor U4253 (N_4253,In_372,In_455);
and U4254 (N_4254,In_1604,In_1899);
nand U4255 (N_4255,In_458,In_1789);
xor U4256 (N_4256,In_20,In_270);
and U4257 (N_4257,In_1505,In_94);
nand U4258 (N_4258,In_851,In_224);
or U4259 (N_4259,In_705,In_1267);
nor U4260 (N_4260,In_1566,In_175);
nand U4261 (N_4261,In_1700,In_444);
nand U4262 (N_4262,In_1796,In_795);
or U4263 (N_4263,In_1144,In_511);
xnor U4264 (N_4264,In_582,In_1787);
nor U4265 (N_4265,In_822,In_1292);
or U4266 (N_4266,In_1479,In_105);
nor U4267 (N_4267,In_1561,In_288);
or U4268 (N_4268,In_300,In_450);
nor U4269 (N_4269,In_622,In_947);
nand U4270 (N_4270,In_1621,In_1833);
nor U4271 (N_4271,In_1393,In_1571);
nor U4272 (N_4272,In_1007,In_277);
nor U4273 (N_4273,In_1696,In_1188);
nor U4274 (N_4274,In_103,In_275);
and U4275 (N_4275,In_1953,In_1814);
or U4276 (N_4276,In_116,In_147);
nor U4277 (N_4277,In_1213,In_1526);
or U4278 (N_4278,In_774,In_558);
and U4279 (N_4279,In_231,In_1915);
nor U4280 (N_4280,In_288,In_1306);
and U4281 (N_4281,In_0,In_643);
or U4282 (N_4282,In_659,In_1925);
nand U4283 (N_4283,In_844,In_1790);
and U4284 (N_4284,In_1909,In_1802);
nand U4285 (N_4285,In_647,In_815);
nand U4286 (N_4286,In_415,In_360);
and U4287 (N_4287,In_204,In_519);
nand U4288 (N_4288,In_984,In_129);
or U4289 (N_4289,In_1811,In_209);
and U4290 (N_4290,In_1758,In_1415);
nand U4291 (N_4291,In_1993,In_1146);
nor U4292 (N_4292,In_356,In_330);
or U4293 (N_4293,In_1171,In_1993);
or U4294 (N_4294,In_334,In_1216);
and U4295 (N_4295,In_1197,In_1605);
nor U4296 (N_4296,In_1900,In_1862);
nand U4297 (N_4297,In_1136,In_1432);
nand U4298 (N_4298,In_1711,In_373);
nor U4299 (N_4299,In_1517,In_15);
and U4300 (N_4300,In_1374,In_1484);
nand U4301 (N_4301,In_866,In_1581);
or U4302 (N_4302,In_1003,In_142);
nand U4303 (N_4303,In_865,In_1376);
nand U4304 (N_4304,In_1840,In_1894);
and U4305 (N_4305,In_1705,In_320);
or U4306 (N_4306,In_1009,In_1248);
nand U4307 (N_4307,In_504,In_1181);
nor U4308 (N_4308,In_1819,In_1706);
or U4309 (N_4309,In_1382,In_786);
xnor U4310 (N_4310,In_1519,In_1353);
or U4311 (N_4311,In_373,In_1182);
nor U4312 (N_4312,In_1484,In_453);
or U4313 (N_4313,In_1085,In_1591);
nor U4314 (N_4314,In_1364,In_1356);
or U4315 (N_4315,In_1070,In_599);
nand U4316 (N_4316,In_1987,In_1747);
nor U4317 (N_4317,In_1993,In_1416);
nand U4318 (N_4318,In_1226,In_1863);
nor U4319 (N_4319,In_883,In_1381);
or U4320 (N_4320,In_1244,In_536);
nand U4321 (N_4321,In_853,In_603);
nand U4322 (N_4322,In_223,In_1978);
and U4323 (N_4323,In_9,In_956);
or U4324 (N_4324,In_1634,In_1830);
xor U4325 (N_4325,In_1622,In_1101);
and U4326 (N_4326,In_1013,In_1103);
or U4327 (N_4327,In_1875,In_482);
and U4328 (N_4328,In_1189,In_782);
nand U4329 (N_4329,In_700,In_692);
and U4330 (N_4330,In_1242,In_81);
or U4331 (N_4331,In_1785,In_1865);
nor U4332 (N_4332,In_695,In_414);
nand U4333 (N_4333,In_1749,In_1299);
or U4334 (N_4334,In_786,In_1577);
or U4335 (N_4335,In_1678,In_1120);
or U4336 (N_4336,In_1909,In_1906);
nor U4337 (N_4337,In_1997,In_899);
nor U4338 (N_4338,In_1680,In_1724);
or U4339 (N_4339,In_145,In_199);
or U4340 (N_4340,In_579,In_58);
nand U4341 (N_4341,In_1383,In_973);
and U4342 (N_4342,In_873,In_1309);
or U4343 (N_4343,In_658,In_554);
nor U4344 (N_4344,In_1521,In_1657);
nor U4345 (N_4345,In_1888,In_1170);
nor U4346 (N_4346,In_1057,In_1615);
nand U4347 (N_4347,In_243,In_1099);
nor U4348 (N_4348,In_1011,In_203);
nor U4349 (N_4349,In_512,In_598);
nor U4350 (N_4350,In_1292,In_255);
nand U4351 (N_4351,In_1276,In_362);
nor U4352 (N_4352,In_158,In_1732);
or U4353 (N_4353,In_1728,In_139);
and U4354 (N_4354,In_1600,In_369);
nand U4355 (N_4355,In_109,In_1949);
and U4356 (N_4356,In_1340,In_1626);
nor U4357 (N_4357,In_1134,In_1111);
and U4358 (N_4358,In_531,In_1461);
nor U4359 (N_4359,In_1976,In_71);
nand U4360 (N_4360,In_880,In_1262);
and U4361 (N_4361,In_1368,In_1825);
nand U4362 (N_4362,In_673,In_1687);
or U4363 (N_4363,In_1186,In_73);
nand U4364 (N_4364,In_1952,In_154);
nand U4365 (N_4365,In_181,In_1761);
nand U4366 (N_4366,In_927,In_72);
or U4367 (N_4367,In_287,In_1474);
nor U4368 (N_4368,In_1068,In_683);
nand U4369 (N_4369,In_558,In_517);
and U4370 (N_4370,In_1945,In_1703);
or U4371 (N_4371,In_1196,In_1592);
nor U4372 (N_4372,In_1734,In_1200);
nand U4373 (N_4373,In_1606,In_1373);
or U4374 (N_4374,In_1730,In_77);
nor U4375 (N_4375,In_613,In_1168);
or U4376 (N_4376,In_1446,In_1669);
or U4377 (N_4377,In_497,In_750);
and U4378 (N_4378,In_1624,In_1473);
or U4379 (N_4379,In_1542,In_1833);
or U4380 (N_4380,In_1590,In_1696);
nand U4381 (N_4381,In_1739,In_438);
nand U4382 (N_4382,In_331,In_1392);
nand U4383 (N_4383,In_1883,In_336);
nor U4384 (N_4384,In_1985,In_1170);
or U4385 (N_4385,In_1061,In_433);
and U4386 (N_4386,In_385,In_886);
nor U4387 (N_4387,In_1765,In_1945);
or U4388 (N_4388,In_1321,In_640);
nor U4389 (N_4389,In_860,In_1160);
nand U4390 (N_4390,In_592,In_1758);
nor U4391 (N_4391,In_1908,In_109);
nand U4392 (N_4392,In_1976,In_1827);
nand U4393 (N_4393,In_1435,In_7);
nor U4394 (N_4394,In_843,In_119);
nand U4395 (N_4395,In_431,In_594);
nand U4396 (N_4396,In_1441,In_1997);
or U4397 (N_4397,In_950,In_1507);
or U4398 (N_4398,In_1048,In_269);
and U4399 (N_4399,In_1213,In_1664);
xnor U4400 (N_4400,In_167,In_1505);
or U4401 (N_4401,In_1964,In_728);
or U4402 (N_4402,In_1651,In_502);
and U4403 (N_4403,In_57,In_152);
or U4404 (N_4404,In_1926,In_137);
or U4405 (N_4405,In_835,In_404);
nand U4406 (N_4406,In_339,In_1140);
nor U4407 (N_4407,In_768,In_293);
and U4408 (N_4408,In_1623,In_736);
nand U4409 (N_4409,In_1338,In_395);
or U4410 (N_4410,In_737,In_645);
or U4411 (N_4411,In_1303,In_1340);
nand U4412 (N_4412,In_1218,In_1237);
nor U4413 (N_4413,In_656,In_481);
xnor U4414 (N_4414,In_499,In_1055);
nor U4415 (N_4415,In_379,In_386);
nand U4416 (N_4416,In_176,In_824);
nor U4417 (N_4417,In_951,In_443);
or U4418 (N_4418,In_559,In_1987);
nor U4419 (N_4419,In_444,In_1304);
nand U4420 (N_4420,In_1415,In_1166);
or U4421 (N_4421,In_984,In_348);
and U4422 (N_4422,In_624,In_705);
nand U4423 (N_4423,In_83,In_1022);
and U4424 (N_4424,In_1847,In_1925);
and U4425 (N_4425,In_855,In_1920);
nand U4426 (N_4426,In_1534,In_324);
and U4427 (N_4427,In_1237,In_1497);
nor U4428 (N_4428,In_564,In_1321);
or U4429 (N_4429,In_369,In_425);
nor U4430 (N_4430,In_737,In_1772);
or U4431 (N_4431,In_1071,In_1445);
or U4432 (N_4432,In_1766,In_517);
and U4433 (N_4433,In_25,In_1873);
nor U4434 (N_4434,In_1748,In_1832);
nor U4435 (N_4435,In_79,In_997);
or U4436 (N_4436,In_1217,In_1442);
xnor U4437 (N_4437,In_1125,In_1086);
and U4438 (N_4438,In_1093,In_555);
or U4439 (N_4439,In_51,In_778);
and U4440 (N_4440,In_643,In_1400);
nor U4441 (N_4441,In_1197,In_1633);
and U4442 (N_4442,In_1373,In_1738);
nand U4443 (N_4443,In_1233,In_1919);
nand U4444 (N_4444,In_124,In_421);
nor U4445 (N_4445,In_1561,In_320);
and U4446 (N_4446,In_685,In_683);
and U4447 (N_4447,In_392,In_719);
nor U4448 (N_4448,In_1926,In_678);
nand U4449 (N_4449,In_171,In_603);
nand U4450 (N_4450,In_481,In_1339);
nor U4451 (N_4451,In_1877,In_1081);
nor U4452 (N_4452,In_8,In_374);
nand U4453 (N_4453,In_1001,In_728);
and U4454 (N_4454,In_579,In_986);
nor U4455 (N_4455,In_475,In_1451);
or U4456 (N_4456,In_1319,In_437);
or U4457 (N_4457,In_496,In_1257);
nand U4458 (N_4458,In_321,In_1631);
and U4459 (N_4459,In_1768,In_1411);
nor U4460 (N_4460,In_414,In_281);
nand U4461 (N_4461,In_1739,In_1338);
nor U4462 (N_4462,In_515,In_829);
nand U4463 (N_4463,In_1186,In_6);
or U4464 (N_4464,In_689,In_1097);
or U4465 (N_4465,In_1007,In_1166);
nor U4466 (N_4466,In_923,In_1559);
and U4467 (N_4467,In_1824,In_503);
nand U4468 (N_4468,In_179,In_387);
nor U4469 (N_4469,In_765,In_1368);
nor U4470 (N_4470,In_1056,In_941);
nor U4471 (N_4471,In_1519,In_109);
or U4472 (N_4472,In_1752,In_583);
and U4473 (N_4473,In_626,In_913);
or U4474 (N_4474,In_1859,In_188);
or U4475 (N_4475,In_1385,In_1423);
or U4476 (N_4476,In_1275,In_609);
nand U4477 (N_4477,In_1036,In_1390);
nand U4478 (N_4478,In_144,In_1695);
nand U4479 (N_4479,In_955,In_528);
nand U4480 (N_4480,In_880,In_1179);
and U4481 (N_4481,In_151,In_180);
nor U4482 (N_4482,In_1429,In_555);
nor U4483 (N_4483,In_500,In_615);
and U4484 (N_4484,In_999,In_1790);
nand U4485 (N_4485,In_1559,In_956);
or U4486 (N_4486,In_475,In_513);
or U4487 (N_4487,In_856,In_1616);
xor U4488 (N_4488,In_837,In_1419);
and U4489 (N_4489,In_617,In_334);
nor U4490 (N_4490,In_240,In_548);
and U4491 (N_4491,In_460,In_1493);
nor U4492 (N_4492,In_614,In_1847);
nor U4493 (N_4493,In_1577,In_95);
or U4494 (N_4494,In_663,In_283);
nor U4495 (N_4495,In_1896,In_1903);
and U4496 (N_4496,In_344,In_572);
and U4497 (N_4497,In_1428,In_658);
or U4498 (N_4498,In_879,In_499);
and U4499 (N_4499,In_1504,In_989);
or U4500 (N_4500,In_929,In_280);
and U4501 (N_4501,In_298,In_372);
nand U4502 (N_4502,In_199,In_29);
nor U4503 (N_4503,In_762,In_1924);
nor U4504 (N_4504,In_59,In_1484);
or U4505 (N_4505,In_1508,In_1220);
nand U4506 (N_4506,In_1408,In_1583);
nor U4507 (N_4507,In_1277,In_431);
or U4508 (N_4508,In_201,In_1435);
nor U4509 (N_4509,In_1911,In_1104);
nor U4510 (N_4510,In_1274,In_587);
nand U4511 (N_4511,In_665,In_123);
and U4512 (N_4512,In_213,In_1777);
and U4513 (N_4513,In_389,In_506);
nand U4514 (N_4514,In_1944,In_1603);
nor U4515 (N_4515,In_1600,In_340);
nor U4516 (N_4516,In_1147,In_1436);
and U4517 (N_4517,In_1097,In_390);
or U4518 (N_4518,In_1998,In_1771);
nand U4519 (N_4519,In_1949,In_147);
or U4520 (N_4520,In_1522,In_975);
and U4521 (N_4521,In_320,In_1385);
or U4522 (N_4522,In_1329,In_160);
or U4523 (N_4523,In_696,In_1332);
or U4524 (N_4524,In_412,In_629);
nand U4525 (N_4525,In_416,In_406);
and U4526 (N_4526,In_1886,In_273);
or U4527 (N_4527,In_1001,In_1306);
or U4528 (N_4528,In_174,In_527);
and U4529 (N_4529,In_1908,In_756);
nor U4530 (N_4530,In_1249,In_547);
and U4531 (N_4531,In_1408,In_1226);
nor U4532 (N_4532,In_440,In_966);
nand U4533 (N_4533,In_1709,In_567);
or U4534 (N_4534,In_616,In_337);
nand U4535 (N_4535,In_1756,In_1317);
nor U4536 (N_4536,In_94,In_66);
or U4537 (N_4537,In_1445,In_222);
nand U4538 (N_4538,In_430,In_924);
nand U4539 (N_4539,In_966,In_1781);
nor U4540 (N_4540,In_687,In_1879);
nand U4541 (N_4541,In_239,In_199);
nand U4542 (N_4542,In_840,In_225);
and U4543 (N_4543,In_1317,In_74);
nor U4544 (N_4544,In_522,In_1531);
nor U4545 (N_4545,In_1212,In_265);
and U4546 (N_4546,In_1181,In_538);
nand U4547 (N_4547,In_1137,In_11);
nor U4548 (N_4548,In_1729,In_175);
or U4549 (N_4549,In_1273,In_1820);
or U4550 (N_4550,In_1813,In_1774);
nor U4551 (N_4551,In_49,In_1980);
nand U4552 (N_4552,In_384,In_331);
or U4553 (N_4553,In_545,In_746);
or U4554 (N_4554,In_155,In_172);
or U4555 (N_4555,In_30,In_1402);
or U4556 (N_4556,In_388,In_1387);
nor U4557 (N_4557,In_1334,In_792);
nand U4558 (N_4558,In_172,In_1914);
or U4559 (N_4559,In_1866,In_257);
nand U4560 (N_4560,In_1390,In_190);
and U4561 (N_4561,In_758,In_604);
or U4562 (N_4562,In_885,In_351);
and U4563 (N_4563,In_303,In_554);
or U4564 (N_4564,In_427,In_876);
nor U4565 (N_4565,In_1168,In_464);
xnor U4566 (N_4566,In_1926,In_1565);
nand U4567 (N_4567,In_1181,In_1734);
and U4568 (N_4568,In_672,In_793);
or U4569 (N_4569,In_307,In_1600);
nand U4570 (N_4570,In_1106,In_1445);
nor U4571 (N_4571,In_588,In_1498);
nand U4572 (N_4572,In_213,In_316);
and U4573 (N_4573,In_1654,In_1408);
or U4574 (N_4574,In_1312,In_81);
nand U4575 (N_4575,In_556,In_761);
nand U4576 (N_4576,In_439,In_1745);
nor U4577 (N_4577,In_781,In_811);
and U4578 (N_4578,In_1839,In_1935);
nor U4579 (N_4579,In_711,In_1553);
and U4580 (N_4580,In_1660,In_1985);
nand U4581 (N_4581,In_1691,In_1545);
and U4582 (N_4582,In_369,In_1484);
nand U4583 (N_4583,In_979,In_1550);
nor U4584 (N_4584,In_1434,In_930);
and U4585 (N_4585,In_340,In_1235);
nor U4586 (N_4586,In_1961,In_270);
nand U4587 (N_4587,In_1101,In_772);
or U4588 (N_4588,In_287,In_1254);
nor U4589 (N_4589,In_1728,In_519);
or U4590 (N_4590,In_1475,In_1886);
nand U4591 (N_4591,In_538,In_59);
nor U4592 (N_4592,In_418,In_295);
nor U4593 (N_4593,In_831,In_1029);
or U4594 (N_4594,In_876,In_1101);
or U4595 (N_4595,In_5,In_413);
nand U4596 (N_4596,In_1317,In_1937);
or U4597 (N_4597,In_859,In_178);
or U4598 (N_4598,In_1878,In_290);
and U4599 (N_4599,In_515,In_1324);
nand U4600 (N_4600,In_1519,In_1751);
nand U4601 (N_4601,In_1337,In_1353);
and U4602 (N_4602,In_793,In_302);
and U4603 (N_4603,In_142,In_1663);
or U4604 (N_4604,In_869,In_305);
nor U4605 (N_4605,In_502,In_706);
nor U4606 (N_4606,In_1020,In_1332);
nor U4607 (N_4607,In_1300,In_1366);
nor U4608 (N_4608,In_747,In_255);
nand U4609 (N_4609,In_184,In_1993);
or U4610 (N_4610,In_655,In_810);
nor U4611 (N_4611,In_222,In_1545);
nor U4612 (N_4612,In_445,In_1949);
nand U4613 (N_4613,In_1171,In_1860);
nand U4614 (N_4614,In_1029,In_854);
nor U4615 (N_4615,In_2,In_465);
and U4616 (N_4616,In_1722,In_536);
and U4617 (N_4617,In_215,In_1103);
nand U4618 (N_4618,In_1211,In_1939);
and U4619 (N_4619,In_1100,In_478);
or U4620 (N_4620,In_860,In_1772);
or U4621 (N_4621,In_183,In_1393);
or U4622 (N_4622,In_1867,In_1847);
nor U4623 (N_4623,In_958,In_742);
nor U4624 (N_4624,In_1829,In_1255);
nor U4625 (N_4625,In_1965,In_75);
or U4626 (N_4626,In_1030,In_283);
nand U4627 (N_4627,In_517,In_1659);
nand U4628 (N_4628,In_1617,In_1995);
or U4629 (N_4629,In_1153,In_433);
nand U4630 (N_4630,In_651,In_125);
or U4631 (N_4631,In_412,In_50);
xor U4632 (N_4632,In_549,In_508);
nand U4633 (N_4633,In_33,In_582);
and U4634 (N_4634,In_1134,In_781);
nor U4635 (N_4635,In_563,In_1038);
nand U4636 (N_4636,In_190,In_742);
and U4637 (N_4637,In_1252,In_1668);
nor U4638 (N_4638,In_1138,In_1287);
nand U4639 (N_4639,In_1118,In_124);
and U4640 (N_4640,In_586,In_1735);
or U4641 (N_4641,In_89,In_239);
or U4642 (N_4642,In_1780,In_1681);
nor U4643 (N_4643,In_913,In_1284);
nor U4644 (N_4644,In_52,In_1931);
or U4645 (N_4645,In_1942,In_1535);
nor U4646 (N_4646,In_1177,In_1048);
nor U4647 (N_4647,In_1413,In_1592);
and U4648 (N_4648,In_294,In_1705);
or U4649 (N_4649,In_782,In_1176);
and U4650 (N_4650,In_70,In_627);
nand U4651 (N_4651,In_157,In_658);
and U4652 (N_4652,In_274,In_165);
and U4653 (N_4653,In_787,In_21);
xnor U4654 (N_4654,In_1273,In_1925);
and U4655 (N_4655,In_1023,In_111);
or U4656 (N_4656,In_1691,In_778);
or U4657 (N_4657,In_1575,In_638);
and U4658 (N_4658,In_1528,In_1785);
nor U4659 (N_4659,In_645,In_1445);
nand U4660 (N_4660,In_483,In_210);
nand U4661 (N_4661,In_1341,In_34);
nand U4662 (N_4662,In_213,In_1961);
nor U4663 (N_4663,In_1503,In_937);
nor U4664 (N_4664,In_1574,In_610);
xnor U4665 (N_4665,In_185,In_28);
nand U4666 (N_4666,In_173,In_888);
or U4667 (N_4667,In_1606,In_333);
and U4668 (N_4668,In_1676,In_819);
or U4669 (N_4669,In_648,In_303);
nand U4670 (N_4670,In_370,In_1376);
or U4671 (N_4671,In_215,In_1645);
and U4672 (N_4672,In_558,In_254);
nor U4673 (N_4673,In_1957,In_306);
or U4674 (N_4674,In_1743,In_1476);
or U4675 (N_4675,In_239,In_940);
and U4676 (N_4676,In_1984,In_1962);
and U4677 (N_4677,In_201,In_1394);
nor U4678 (N_4678,In_364,In_270);
and U4679 (N_4679,In_1701,In_1205);
and U4680 (N_4680,In_1664,In_1812);
and U4681 (N_4681,In_1041,In_357);
and U4682 (N_4682,In_1,In_862);
or U4683 (N_4683,In_746,In_1233);
and U4684 (N_4684,In_1073,In_559);
nand U4685 (N_4685,In_1938,In_835);
or U4686 (N_4686,In_1060,In_1013);
and U4687 (N_4687,In_228,In_1424);
nor U4688 (N_4688,In_638,In_1953);
nand U4689 (N_4689,In_333,In_1813);
or U4690 (N_4690,In_1298,In_677);
nand U4691 (N_4691,In_592,In_1834);
or U4692 (N_4692,In_1971,In_1597);
and U4693 (N_4693,In_476,In_1553);
or U4694 (N_4694,In_167,In_771);
nand U4695 (N_4695,In_372,In_1682);
nor U4696 (N_4696,In_395,In_1752);
nand U4697 (N_4697,In_1466,In_802);
nor U4698 (N_4698,In_320,In_1572);
or U4699 (N_4699,In_707,In_958);
nor U4700 (N_4700,In_1026,In_1728);
nand U4701 (N_4701,In_1767,In_1476);
or U4702 (N_4702,In_1318,In_811);
nand U4703 (N_4703,In_829,In_1008);
xnor U4704 (N_4704,In_449,In_266);
nor U4705 (N_4705,In_786,In_825);
or U4706 (N_4706,In_1939,In_639);
nand U4707 (N_4707,In_869,In_434);
nor U4708 (N_4708,In_1447,In_1780);
nor U4709 (N_4709,In_95,In_906);
and U4710 (N_4710,In_897,In_495);
and U4711 (N_4711,In_260,In_553);
nand U4712 (N_4712,In_925,In_246);
nor U4713 (N_4713,In_614,In_322);
and U4714 (N_4714,In_1970,In_498);
nand U4715 (N_4715,In_300,In_1437);
nor U4716 (N_4716,In_578,In_242);
nand U4717 (N_4717,In_1305,In_1350);
or U4718 (N_4718,In_1576,In_398);
nor U4719 (N_4719,In_1962,In_1161);
or U4720 (N_4720,In_738,In_60);
or U4721 (N_4721,In_177,In_1348);
nor U4722 (N_4722,In_804,In_1784);
nor U4723 (N_4723,In_1789,In_397);
nor U4724 (N_4724,In_71,In_1954);
nand U4725 (N_4725,In_142,In_983);
and U4726 (N_4726,In_1117,In_139);
xor U4727 (N_4727,In_1463,In_1205);
and U4728 (N_4728,In_1730,In_645);
or U4729 (N_4729,In_1344,In_778);
or U4730 (N_4730,In_501,In_1053);
and U4731 (N_4731,In_1659,In_388);
nor U4732 (N_4732,In_465,In_1043);
nand U4733 (N_4733,In_1952,In_1902);
and U4734 (N_4734,In_648,In_1423);
and U4735 (N_4735,In_1645,In_528);
nor U4736 (N_4736,In_967,In_278);
and U4737 (N_4737,In_500,In_682);
or U4738 (N_4738,In_698,In_1834);
nor U4739 (N_4739,In_765,In_1321);
and U4740 (N_4740,In_812,In_409);
or U4741 (N_4741,In_1564,In_660);
or U4742 (N_4742,In_675,In_852);
nand U4743 (N_4743,In_901,In_1091);
and U4744 (N_4744,In_978,In_1670);
nand U4745 (N_4745,In_1359,In_664);
and U4746 (N_4746,In_1652,In_681);
or U4747 (N_4747,In_888,In_867);
or U4748 (N_4748,In_1079,In_714);
nand U4749 (N_4749,In_309,In_1486);
nor U4750 (N_4750,In_1530,In_1067);
and U4751 (N_4751,In_798,In_1930);
and U4752 (N_4752,In_51,In_38);
or U4753 (N_4753,In_556,In_1680);
nor U4754 (N_4754,In_708,In_475);
nand U4755 (N_4755,In_1411,In_1724);
nand U4756 (N_4756,In_1372,In_728);
nor U4757 (N_4757,In_1960,In_1163);
nor U4758 (N_4758,In_1105,In_1367);
or U4759 (N_4759,In_159,In_611);
or U4760 (N_4760,In_113,In_333);
or U4761 (N_4761,In_57,In_1223);
nor U4762 (N_4762,In_883,In_1526);
nand U4763 (N_4763,In_1058,In_1670);
and U4764 (N_4764,In_523,In_1819);
nor U4765 (N_4765,In_1755,In_389);
and U4766 (N_4766,In_1881,In_712);
nand U4767 (N_4767,In_191,In_110);
and U4768 (N_4768,In_1481,In_1706);
nand U4769 (N_4769,In_384,In_576);
and U4770 (N_4770,In_1710,In_222);
or U4771 (N_4771,In_94,In_1456);
xnor U4772 (N_4772,In_1768,In_1662);
nor U4773 (N_4773,In_493,In_1450);
nand U4774 (N_4774,In_1928,In_1093);
nand U4775 (N_4775,In_1160,In_1979);
and U4776 (N_4776,In_1861,In_1433);
nand U4777 (N_4777,In_482,In_455);
nor U4778 (N_4778,In_1364,In_96);
or U4779 (N_4779,In_1052,In_429);
or U4780 (N_4780,In_1014,In_477);
and U4781 (N_4781,In_933,In_1010);
and U4782 (N_4782,In_1868,In_882);
and U4783 (N_4783,In_1095,In_438);
nor U4784 (N_4784,In_1977,In_796);
or U4785 (N_4785,In_763,In_1599);
nand U4786 (N_4786,In_1791,In_252);
nand U4787 (N_4787,In_698,In_1556);
and U4788 (N_4788,In_1320,In_921);
nand U4789 (N_4789,In_235,In_1624);
nor U4790 (N_4790,In_457,In_123);
nand U4791 (N_4791,In_112,In_1755);
nor U4792 (N_4792,In_416,In_832);
nand U4793 (N_4793,In_1753,In_1868);
and U4794 (N_4794,In_1304,In_1029);
nand U4795 (N_4795,In_1509,In_948);
nor U4796 (N_4796,In_951,In_1871);
and U4797 (N_4797,In_1418,In_885);
and U4798 (N_4798,In_1041,In_1662);
nor U4799 (N_4799,In_78,In_1167);
nand U4800 (N_4800,In_586,In_1399);
or U4801 (N_4801,In_64,In_1430);
or U4802 (N_4802,In_464,In_757);
nand U4803 (N_4803,In_142,In_1643);
nor U4804 (N_4804,In_1443,In_1138);
nor U4805 (N_4805,In_532,In_196);
nor U4806 (N_4806,In_383,In_439);
and U4807 (N_4807,In_1371,In_1693);
or U4808 (N_4808,In_739,In_1988);
and U4809 (N_4809,In_771,In_1416);
nor U4810 (N_4810,In_1113,In_1428);
or U4811 (N_4811,In_1571,In_1911);
and U4812 (N_4812,In_1169,In_144);
nor U4813 (N_4813,In_1132,In_327);
nor U4814 (N_4814,In_281,In_1337);
nor U4815 (N_4815,In_237,In_281);
nor U4816 (N_4816,In_788,In_768);
nor U4817 (N_4817,In_681,In_899);
nand U4818 (N_4818,In_1659,In_1669);
nand U4819 (N_4819,In_1492,In_237);
nand U4820 (N_4820,In_1878,In_783);
and U4821 (N_4821,In_1139,In_970);
nor U4822 (N_4822,In_1080,In_1355);
or U4823 (N_4823,In_216,In_1533);
nor U4824 (N_4824,In_467,In_411);
or U4825 (N_4825,In_180,In_1260);
and U4826 (N_4826,In_991,In_17);
nor U4827 (N_4827,In_1903,In_1981);
nand U4828 (N_4828,In_352,In_10);
and U4829 (N_4829,In_626,In_1620);
nand U4830 (N_4830,In_305,In_409);
nor U4831 (N_4831,In_785,In_176);
nor U4832 (N_4832,In_535,In_513);
nor U4833 (N_4833,In_1479,In_281);
or U4834 (N_4834,In_243,In_762);
nand U4835 (N_4835,In_544,In_585);
nand U4836 (N_4836,In_1105,In_1467);
or U4837 (N_4837,In_1317,In_200);
nand U4838 (N_4838,In_957,In_1432);
or U4839 (N_4839,In_274,In_1605);
nor U4840 (N_4840,In_772,In_552);
nand U4841 (N_4841,In_1787,In_839);
nand U4842 (N_4842,In_1445,In_1317);
nor U4843 (N_4843,In_507,In_1328);
and U4844 (N_4844,In_978,In_762);
and U4845 (N_4845,In_0,In_1971);
nor U4846 (N_4846,In_1147,In_49);
nor U4847 (N_4847,In_821,In_602);
or U4848 (N_4848,In_1043,In_588);
or U4849 (N_4849,In_127,In_1764);
and U4850 (N_4850,In_1351,In_1454);
and U4851 (N_4851,In_1152,In_1775);
and U4852 (N_4852,In_1476,In_253);
nor U4853 (N_4853,In_1193,In_365);
or U4854 (N_4854,In_1454,In_532);
nand U4855 (N_4855,In_860,In_786);
nor U4856 (N_4856,In_887,In_1042);
and U4857 (N_4857,In_1784,In_261);
nor U4858 (N_4858,In_1143,In_1586);
nor U4859 (N_4859,In_1923,In_1327);
nor U4860 (N_4860,In_58,In_1618);
or U4861 (N_4861,In_1685,In_526);
nand U4862 (N_4862,In_1039,In_1424);
and U4863 (N_4863,In_1186,In_1254);
nor U4864 (N_4864,In_577,In_1878);
and U4865 (N_4865,In_95,In_1489);
and U4866 (N_4866,In_1702,In_1501);
and U4867 (N_4867,In_1440,In_1499);
nand U4868 (N_4868,In_684,In_528);
and U4869 (N_4869,In_1455,In_135);
or U4870 (N_4870,In_1161,In_427);
and U4871 (N_4871,In_791,In_770);
and U4872 (N_4872,In_14,In_973);
nand U4873 (N_4873,In_130,In_568);
nor U4874 (N_4874,In_787,In_892);
and U4875 (N_4875,In_451,In_1098);
and U4876 (N_4876,In_1245,In_1071);
nand U4877 (N_4877,In_1573,In_691);
and U4878 (N_4878,In_619,In_1245);
nand U4879 (N_4879,In_48,In_1191);
nor U4880 (N_4880,In_1701,In_53);
or U4881 (N_4881,In_1312,In_657);
nor U4882 (N_4882,In_1137,In_531);
nand U4883 (N_4883,In_1583,In_1080);
nor U4884 (N_4884,In_1593,In_1417);
or U4885 (N_4885,In_1044,In_881);
nand U4886 (N_4886,In_1106,In_1713);
or U4887 (N_4887,In_181,In_308);
or U4888 (N_4888,In_1343,In_325);
nand U4889 (N_4889,In_448,In_1618);
nand U4890 (N_4890,In_476,In_1861);
and U4891 (N_4891,In_161,In_209);
or U4892 (N_4892,In_984,In_1957);
nand U4893 (N_4893,In_1599,In_348);
nor U4894 (N_4894,In_423,In_1584);
nand U4895 (N_4895,In_1198,In_196);
or U4896 (N_4896,In_709,In_353);
nor U4897 (N_4897,In_975,In_34);
or U4898 (N_4898,In_1928,In_307);
and U4899 (N_4899,In_1013,In_87);
nor U4900 (N_4900,In_1537,In_527);
nand U4901 (N_4901,In_1025,In_237);
and U4902 (N_4902,In_1524,In_1988);
nor U4903 (N_4903,In_971,In_1117);
and U4904 (N_4904,In_1901,In_638);
nand U4905 (N_4905,In_240,In_1536);
and U4906 (N_4906,In_1011,In_439);
or U4907 (N_4907,In_1168,In_783);
nor U4908 (N_4908,In_989,In_332);
or U4909 (N_4909,In_825,In_698);
or U4910 (N_4910,In_90,In_1471);
nor U4911 (N_4911,In_590,In_1198);
and U4912 (N_4912,In_14,In_181);
nor U4913 (N_4913,In_680,In_812);
or U4914 (N_4914,In_1147,In_679);
nand U4915 (N_4915,In_1297,In_1488);
nand U4916 (N_4916,In_231,In_1148);
nand U4917 (N_4917,In_700,In_863);
nand U4918 (N_4918,In_593,In_336);
or U4919 (N_4919,In_38,In_838);
and U4920 (N_4920,In_921,In_1539);
nor U4921 (N_4921,In_725,In_643);
nand U4922 (N_4922,In_1452,In_1839);
nor U4923 (N_4923,In_1985,In_1367);
and U4924 (N_4924,In_350,In_135);
nor U4925 (N_4925,In_1256,In_802);
or U4926 (N_4926,In_1969,In_721);
nor U4927 (N_4927,In_1958,In_746);
nand U4928 (N_4928,In_1143,In_260);
nand U4929 (N_4929,In_408,In_1808);
and U4930 (N_4930,In_185,In_633);
or U4931 (N_4931,In_815,In_343);
nand U4932 (N_4932,In_425,In_580);
nand U4933 (N_4933,In_1221,In_1434);
or U4934 (N_4934,In_1214,In_268);
nor U4935 (N_4935,In_1659,In_1270);
or U4936 (N_4936,In_470,In_99);
nor U4937 (N_4937,In_366,In_318);
nand U4938 (N_4938,In_880,In_863);
or U4939 (N_4939,In_1005,In_1624);
and U4940 (N_4940,In_397,In_1713);
and U4941 (N_4941,In_1069,In_1669);
and U4942 (N_4942,In_1626,In_839);
or U4943 (N_4943,In_201,In_1880);
or U4944 (N_4944,In_570,In_810);
or U4945 (N_4945,In_402,In_1893);
nor U4946 (N_4946,In_1839,In_1612);
or U4947 (N_4947,In_947,In_1270);
or U4948 (N_4948,In_1884,In_1384);
and U4949 (N_4949,In_345,In_194);
or U4950 (N_4950,In_801,In_35);
and U4951 (N_4951,In_613,In_1841);
nor U4952 (N_4952,In_477,In_1104);
and U4953 (N_4953,In_1226,In_583);
and U4954 (N_4954,In_461,In_1682);
nand U4955 (N_4955,In_1055,In_451);
or U4956 (N_4956,In_782,In_1385);
or U4957 (N_4957,In_1496,In_929);
and U4958 (N_4958,In_428,In_109);
or U4959 (N_4959,In_755,In_1970);
nor U4960 (N_4960,In_83,In_651);
nand U4961 (N_4961,In_1706,In_783);
nand U4962 (N_4962,In_1403,In_494);
and U4963 (N_4963,In_11,In_776);
nand U4964 (N_4964,In_1513,In_260);
or U4965 (N_4965,In_1007,In_1868);
nor U4966 (N_4966,In_1063,In_1710);
and U4967 (N_4967,In_610,In_1153);
or U4968 (N_4968,In_1759,In_86);
or U4969 (N_4969,In_1169,In_762);
xnor U4970 (N_4970,In_593,In_1989);
or U4971 (N_4971,In_290,In_1915);
and U4972 (N_4972,In_1918,In_877);
and U4973 (N_4973,In_1167,In_1457);
nor U4974 (N_4974,In_1693,In_25);
or U4975 (N_4975,In_312,In_930);
xor U4976 (N_4976,In_743,In_1944);
or U4977 (N_4977,In_1231,In_425);
nand U4978 (N_4978,In_1562,In_1338);
nand U4979 (N_4979,In_1815,In_163);
and U4980 (N_4980,In_474,In_575);
nor U4981 (N_4981,In_1649,In_675);
and U4982 (N_4982,In_494,In_1816);
nand U4983 (N_4983,In_1318,In_1905);
or U4984 (N_4984,In_1754,In_1244);
nand U4985 (N_4985,In_574,In_1913);
nor U4986 (N_4986,In_113,In_1031);
nand U4987 (N_4987,In_798,In_590);
nor U4988 (N_4988,In_419,In_151);
nor U4989 (N_4989,In_854,In_1937);
and U4990 (N_4990,In_271,In_306);
and U4991 (N_4991,In_788,In_1);
nand U4992 (N_4992,In_596,In_173);
nor U4993 (N_4993,In_139,In_1203);
nor U4994 (N_4994,In_1741,In_1177);
or U4995 (N_4995,In_298,In_1124);
or U4996 (N_4996,In_753,In_819);
and U4997 (N_4997,In_266,In_1759);
and U4998 (N_4998,In_1327,In_971);
and U4999 (N_4999,In_1074,In_691);
and U5000 (N_5000,N_568,N_3984);
or U5001 (N_5001,N_4783,N_2988);
nand U5002 (N_5002,N_2024,N_2642);
or U5003 (N_5003,N_2569,N_2644);
and U5004 (N_5004,N_4049,N_2512);
nand U5005 (N_5005,N_4058,N_2810);
nor U5006 (N_5006,N_3558,N_2052);
and U5007 (N_5007,N_240,N_2539);
and U5008 (N_5008,N_3274,N_1142);
or U5009 (N_5009,N_4556,N_3905);
and U5010 (N_5010,N_3157,N_3396);
and U5011 (N_5011,N_1014,N_4247);
nand U5012 (N_5012,N_305,N_3115);
nand U5013 (N_5013,N_1514,N_849);
and U5014 (N_5014,N_4963,N_838);
and U5015 (N_5015,N_2541,N_4747);
nor U5016 (N_5016,N_2470,N_736);
and U5017 (N_5017,N_3304,N_1256);
nor U5018 (N_5018,N_1577,N_1333);
and U5019 (N_5019,N_2974,N_4444);
nor U5020 (N_5020,N_463,N_2911);
and U5021 (N_5021,N_388,N_3895);
or U5022 (N_5022,N_3767,N_2095);
and U5023 (N_5023,N_4347,N_3764);
or U5024 (N_5024,N_1557,N_258);
nor U5025 (N_5025,N_991,N_3956);
or U5026 (N_5026,N_3281,N_2181);
or U5027 (N_5027,N_1175,N_3441);
nor U5028 (N_5028,N_3527,N_3769);
nand U5029 (N_5029,N_1075,N_577);
and U5030 (N_5030,N_1431,N_2110);
and U5031 (N_5031,N_3900,N_4284);
and U5032 (N_5032,N_3692,N_1642);
or U5033 (N_5033,N_4136,N_3319);
or U5034 (N_5034,N_4588,N_1796);
or U5035 (N_5035,N_92,N_3091);
or U5036 (N_5036,N_3418,N_3989);
or U5037 (N_5037,N_2792,N_1835);
and U5038 (N_5038,N_1461,N_1071);
or U5039 (N_5039,N_5,N_937);
nand U5040 (N_5040,N_1424,N_2838);
or U5041 (N_5041,N_2937,N_4786);
nand U5042 (N_5042,N_4387,N_2383);
and U5043 (N_5043,N_1073,N_978);
and U5044 (N_5044,N_4709,N_4408);
nand U5045 (N_5045,N_4238,N_1053);
or U5046 (N_5046,N_3676,N_3585);
and U5047 (N_5047,N_2057,N_2578);
or U5048 (N_5048,N_3272,N_3716);
nand U5049 (N_5049,N_3062,N_1485);
and U5050 (N_5050,N_98,N_4380);
nand U5051 (N_5051,N_606,N_4397);
and U5052 (N_5052,N_1715,N_3361);
nand U5053 (N_5053,N_4517,N_830);
nand U5054 (N_5054,N_3871,N_4606);
nand U5055 (N_5055,N_1049,N_3647);
nor U5056 (N_5056,N_2670,N_2674);
and U5057 (N_5057,N_94,N_468);
nand U5058 (N_5058,N_4390,N_1327);
or U5059 (N_5059,N_4946,N_4642);
nor U5060 (N_5060,N_2149,N_1566);
and U5061 (N_5061,N_4314,N_3011);
or U5062 (N_5062,N_3301,N_1776);
and U5063 (N_5063,N_4173,N_3000);
nor U5064 (N_5064,N_3753,N_1900);
nor U5065 (N_5065,N_1916,N_4596);
and U5066 (N_5066,N_4940,N_4042);
and U5067 (N_5067,N_89,N_903);
nor U5068 (N_5068,N_1180,N_821);
or U5069 (N_5069,N_3076,N_2069);
nor U5070 (N_5070,N_3582,N_3508);
and U5071 (N_5071,N_3873,N_928);
nand U5072 (N_5072,N_4743,N_3089);
nor U5073 (N_5073,N_3284,N_3721);
and U5074 (N_5074,N_4666,N_1598);
or U5075 (N_5075,N_4643,N_1027);
and U5076 (N_5076,N_1126,N_1940);
or U5077 (N_5077,N_3228,N_340);
xor U5078 (N_5078,N_1948,N_4644);
nand U5079 (N_5079,N_2289,N_4610);
nor U5080 (N_5080,N_3183,N_2272);
nor U5081 (N_5081,N_706,N_4865);
nand U5082 (N_5082,N_646,N_3487);
xor U5083 (N_5083,N_106,N_3724);
or U5084 (N_5084,N_1058,N_2604);
nor U5085 (N_5085,N_4029,N_4857);
nand U5086 (N_5086,N_4075,N_1910);
or U5087 (N_5087,N_2793,N_3636);
or U5088 (N_5088,N_1930,N_1280);
and U5089 (N_5089,N_3077,N_1960);
nand U5090 (N_5090,N_2517,N_3860);
and U5091 (N_5091,N_2100,N_1774);
and U5092 (N_5092,N_1119,N_3863);
xor U5093 (N_5093,N_4785,N_1045);
nor U5094 (N_5094,N_134,N_1618);
or U5095 (N_5095,N_1068,N_3739);
or U5096 (N_5096,N_1095,N_1330);
or U5097 (N_5097,N_197,N_2285);
and U5098 (N_5098,N_20,N_4132);
nand U5099 (N_5099,N_4420,N_3291);
nor U5100 (N_5100,N_1007,N_1161);
and U5101 (N_5101,N_1662,N_4683);
nor U5102 (N_5102,N_1989,N_2653);
nor U5103 (N_5103,N_1301,N_4030);
nor U5104 (N_5104,N_4595,N_2135);
nor U5105 (N_5105,N_1286,N_822);
or U5106 (N_5106,N_3188,N_4613);
nand U5107 (N_5107,N_2909,N_2115);
and U5108 (N_5108,N_2805,N_2431);
nor U5109 (N_5109,N_3922,N_853);
or U5110 (N_5110,N_1714,N_1993);
nand U5111 (N_5111,N_1483,N_4543);
nand U5112 (N_5112,N_3293,N_3914);
and U5113 (N_5113,N_515,N_1754);
nor U5114 (N_5114,N_4125,N_3203);
nor U5115 (N_5115,N_2331,N_1460);
or U5116 (N_5116,N_2968,N_4482);
or U5117 (N_5117,N_1229,N_1310);
and U5118 (N_5118,N_2048,N_4922);
nor U5119 (N_5119,N_2593,N_895);
nand U5120 (N_5120,N_4591,N_3757);
or U5121 (N_5121,N_2926,N_2319);
nor U5122 (N_5122,N_694,N_3014);
nand U5123 (N_5123,N_656,N_4685);
and U5124 (N_5124,N_3916,N_1607);
nor U5125 (N_5125,N_4676,N_2628);
nand U5126 (N_5126,N_4241,N_4013);
nor U5127 (N_5127,N_101,N_3363);
nand U5128 (N_5128,N_3273,N_145);
nor U5129 (N_5129,N_3229,N_4102);
and U5130 (N_5130,N_1364,N_4593);
nand U5131 (N_5131,N_803,N_3933);
and U5132 (N_5132,N_2071,N_1169);
nor U5133 (N_5133,N_3479,N_4586);
and U5134 (N_5134,N_4501,N_363);
nand U5135 (N_5135,N_3019,N_1628);
and U5136 (N_5136,N_3109,N_715);
or U5137 (N_5137,N_3731,N_3384);
or U5138 (N_5138,N_3619,N_3867);
and U5139 (N_5139,N_1140,N_4536);
nor U5140 (N_5140,N_41,N_4693);
and U5141 (N_5141,N_875,N_1672);
nand U5142 (N_5142,N_4359,N_4008);
and U5143 (N_5143,N_971,N_4090);
and U5144 (N_5144,N_1663,N_4291);
nor U5145 (N_5145,N_2086,N_720);
and U5146 (N_5146,N_808,N_4781);
or U5147 (N_5147,N_2066,N_3249);
nand U5148 (N_5148,N_1089,N_3897);
nor U5149 (N_5149,N_1845,N_2065);
nor U5150 (N_5150,N_176,N_2671);
nand U5151 (N_5151,N_4761,N_2932);
nand U5152 (N_5152,N_1625,N_3199);
or U5153 (N_5153,N_1814,N_1291);
nor U5154 (N_5154,N_2186,N_2298);
and U5155 (N_5155,N_2236,N_2006);
nand U5156 (N_5156,N_2162,N_2627);
nor U5157 (N_5157,N_1030,N_374);
and U5158 (N_5158,N_3518,N_1329);
nand U5159 (N_5159,N_1252,N_1970);
xnor U5160 (N_5160,N_3110,N_4389);
nor U5161 (N_5161,N_1187,N_4634);
and U5162 (N_5162,N_4858,N_1455);
and U5163 (N_5163,N_3821,N_3126);
nor U5164 (N_5164,N_2336,N_2238);
or U5165 (N_5165,N_864,N_3775);
nand U5166 (N_5166,N_2920,N_4934);
xnor U5167 (N_5167,N_3413,N_1253);
or U5168 (N_5168,N_2786,N_2630);
and U5169 (N_5169,N_2324,N_1885);
nand U5170 (N_5170,N_4778,N_890);
or U5171 (N_5171,N_1406,N_3697);
or U5172 (N_5172,N_4776,N_2905);
nor U5173 (N_5173,N_2606,N_934);
and U5174 (N_5174,N_3197,N_3111);
or U5175 (N_5175,N_3950,N_188);
or U5176 (N_5176,N_933,N_1235);
and U5177 (N_5177,N_329,N_4849);
and U5178 (N_5178,N_3499,N_3377);
and U5179 (N_5179,N_4711,N_1454);
or U5180 (N_5180,N_1047,N_1304);
nor U5181 (N_5181,N_233,N_393);
nor U5182 (N_5182,N_2405,N_2170);
nand U5183 (N_5183,N_1933,N_2465);
and U5184 (N_5184,N_4334,N_508);
nand U5185 (N_5185,N_1387,N_4718);
or U5186 (N_5186,N_3358,N_4060);
or U5187 (N_5187,N_2344,N_4765);
nand U5188 (N_5188,N_1323,N_1318);
or U5189 (N_5189,N_1787,N_2664);
nand U5190 (N_5190,N_4128,N_1317);
nor U5191 (N_5191,N_732,N_4686);
nand U5192 (N_5192,N_1353,N_462);
nor U5193 (N_5193,N_4253,N_4119);
nand U5194 (N_5194,N_2146,N_2801);
nor U5195 (N_5195,N_2998,N_2143);
nor U5196 (N_5196,N_4897,N_4520);
nor U5197 (N_5197,N_1171,N_4821);
and U5198 (N_5198,N_3806,N_396);
or U5199 (N_5199,N_1769,N_4364);
or U5200 (N_5200,N_8,N_1349);
or U5201 (N_5201,N_2037,N_2242);
and U5202 (N_5202,N_2262,N_4590);
and U5203 (N_5203,N_4848,N_2680);
nand U5204 (N_5204,N_200,N_1464);
or U5205 (N_5205,N_1024,N_4016);
nand U5206 (N_5206,N_1004,N_3569);
and U5207 (N_5207,N_4037,N_744);
nor U5208 (N_5208,N_2827,N_251);
nor U5209 (N_5209,N_4023,N_1467);
or U5210 (N_5210,N_3432,N_4887);
and U5211 (N_5211,N_1409,N_1328);
and U5212 (N_5212,N_4679,N_4218);
nor U5213 (N_5213,N_2546,N_1549);
and U5214 (N_5214,N_813,N_31);
nand U5215 (N_5215,N_1442,N_3161);
nand U5216 (N_5216,N_4758,N_2545);
or U5217 (N_5217,N_2661,N_686);
nor U5218 (N_5218,N_3024,N_629);
nor U5219 (N_5219,N_3113,N_3788);
or U5220 (N_5220,N_973,N_3765);
and U5221 (N_5221,N_1636,N_3064);
nor U5222 (N_5222,N_2172,N_4001);
nand U5223 (N_5223,N_23,N_3918);
and U5224 (N_5224,N_461,N_4196);
and U5225 (N_5225,N_3285,N_2798);
and U5226 (N_5226,N_1553,N_3594);
and U5227 (N_5227,N_2113,N_2097);
and U5228 (N_5228,N_385,N_311);
or U5229 (N_5229,N_2073,N_817);
nor U5230 (N_5230,N_2053,N_2976);
or U5231 (N_5231,N_1121,N_2111);
or U5232 (N_5232,N_2326,N_2585);
and U5233 (N_5233,N_4026,N_3093);
nand U5234 (N_5234,N_3350,N_1360);
and U5235 (N_5235,N_758,N_3618);
nand U5236 (N_5236,N_2571,N_2273);
nand U5237 (N_5237,N_4235,N_4830);
nor U5238 (N_5238,N_2466,N_3470);
nor U5239 (N_5239,N_35,N_3190);
and U5240 (N_5240,N_3565,N_4394);
nor U5241 (N_5241,N_2624,N_668);
nand U5242 (N_5242,N_2449,N_2646);
or U5243 (N_5243,N_584,N_1770);
nand U5244 (N_5244,N_219,N_2865);
nand U5245 (N_5245,N_905,N_1655);
nor U5246 (N_5246,N_1762,N_2590);
nand U5247 (N_5247,N_2257,N_4532);
or U5248 (N_5248,N_2244,N_4752);
nand U5249 (N_5249,N_4583,N_2581);
and U5250 (N_5250,N_512,N_1249);
or U5251 (N_5251,N_157,N_3294);
nor U5252 (N_5252,N_4257,N_2775);
or U5253 (N_5253,N_1673,N_4975);
nand U5254 (N_5254,N_2315,N_1681);
and U5255 (N_5255,N_1730,N_286);
nand U5256 (N_5256,N_3845,N_2212);
nand U5257 (N_5257,N_4920,N_625);
or U5258 (N_5258,N_2211,N_1222);
nand U5259 (N_5259,N_392,N_4348);
or U5260 (N_5260,N_1477,N_77);
nor U5261 (N_5261,N_1279,N_1240);
and U5262 (N_5262,N_2046,N_892);
nor U5263 (N_5263,N_1688,N_3898);
or U5264 (N_5264,N_4872,N_173);
nand U5265 (N_5265,N_659,N_3887);
and U5266 (N_5266,N_1895,N_1810);
and U5267 (N_5267,N_189,N_2643);
nand U5268 (N_5268,N_3768,N_4764);
and U5269 (N_5269,N_1021,N_3399);
or U5270 (N_5270,N_1729,N_1778);
nand U5271 (N_5271,N_2364,N_2044);
nand U5272 (N_5272,N_4689,N_1670);
and U5273 (N_5273,N_3392,N_246);
or U5274 (N_5274,N_3570,N_3810);
and U5275 (N_5275,N_3118,N_2879);
nand U5276 (N_5276,N_919,N_3861);
and U5277 (N_5277,N_2663,N_4889);
and U5278 (N_5278,N_1182,N_1141);
nand U5279 (N_5279,N_2791,N_2996);
nor U5280 (N_5280,N_2462,N_1443);
or U5281 (N_5281,N_2596,N_4112);
nand U5282 (N_5282,N_801,N_1669);
or U5283 (N_5283,N_1435,N_3991);
and U5284 (N_5284,N_2999,N_3778);
nand U5285 (N_5285,N_3711,N_467);
nor U5286 (N_5286,N_4627,N_1639);
nand U5287 (N_5287,N_4386,N_525);
or U5288 (N_5288,N_4289,N_1504);
and U5289 (N_5289,N_3774,N_1338);
nor U5290 (N_5290,N_3114,N_3187);
and U5291 (N_5291,N_1649,N_2860);
or U5292 (N_5292,N_1255,N_1659);
xnor U5293 (N_5293,N_4856,N_105);
nor U5294 (N_5294,N_3397,N_436);
nor U5295 (N_5295,N_3435,N_1275);
nor U5296 (N_5296,N_3206,N_4991);
nor U5297 (N_5297,N_2304,N_1740);
and U5298 (N_5298,N_2036,N_1055);
and U5299 (N_5299,N_676,N_3543);
and U5300 (N_5300,N_526,N_4398);
nor U5301 (N_5301,N_2544,N_3428);
and U5302 (N_5302,N_3815,N_2963);
or U5303 (N_5303,N_4226,N_3101);
and U5304 (N_5304,N_2339,N_3560);
or U5305 (N_5305,N_4742,N_4913);
nor U5306 (N_5306,N_4053,N_2766);
or U5307 (N_5307,N_1959,N_4962);
nor U5308 (N_5308,N_669,N_1159);
or U5309 (N_5309,N_519,N_4101);
and U5310 (N_5310,N_1491,N_2455);
nor U5311 (N_5311,N_3278,N_4714);
or U5312 (N_5312,N_4004,N_1147);
and U5313 (N_5313,N_2514,N_947);
or U5314 (N_5314,N_2558,N_1154);
and U5315 (N_5315,N_3255,N_2323);
nor U5316 (N_5316,N_1416,N_4937);
or U5317 (N_5317,N_643,N_3971);
and U5318 (N_5318,N_38,N_636);
and U5319 (N_5319,N_221,N_2338);
and U5320 (N_5320,N_4371,N_3528);
nor U5321 (N_5321,N_2270,N_1368);
nor U5322 (N_5322,N_762,N_4771);
and U5323 (N_5323,N_3877,N_4234);
nor U5324 (N_5324,N_4094,N_2842);
or U5325 (N_5325,N_2609,N_4483);
or U5326 (N_5326,N_3364,N_2283);
or U5327 (N_5327,N_2369,N_3913);
nand U5328 (N_5328,N_3927,N_2467);
nor U5329 (N_5329,N_3885,N_306);
or U5330 (N_5330,N_218,N_1979);
xnor U5331 (N_5331,N_1295,N_170);
and U5332 (N_5332,N_1674,N_2045);
nand U5333 (N_5333,N_109,N_2991);
nand U5334 (N_5334,N_769,N_1379);
nand U5335 (N_5335,N_418,N_824);
nor U5336 (N_5336,N_1798,N_3705);
and U5337 (N_5337,N_1597,N_2787);
nand U5338 (N_5338,N_399,N_1032);
or U5339 (N_5339,N_2278,N_351);
or U5340 (N_5340,N_4375,N_4938);
or U5341 (N_5341,N_2328,N_551);
nand U5342 (N_5342,N_4510,N_2524);
and U5343 (N_5343,N_2249,N_2830);
and U5344 (N_5344,N_548,N_4189);
nand U5345 (N_5345,N_3303,N_4722);
nor U5346 (N_5346,N_4108,N_865);
and U5347 (N_5347,N_786,N_4274);
nor U5348 (N_5348,N_2009,N_2707);
and U5349 (N_5349,N_4808,N_2521);
nor U5350 (N_5350,N_842,N_415);
or U5351 (N_5351,N_3082,N_1965);
nand U5352 (N_5352,N_3696,N_360);
nor U5353 (N_5353,N_495,N_3473);
or U5354 (N_5354,N_4999,N_4163);
and U5355 (N_5355,N_2892,N_2358);
and U5356 (N_5356,N_1228,N_0);
or U5357 (N_5357,N_1727,N_3953);
nand U5358 (N_5358,N_3192,N_2333);
nand U5359 (N_5359,N_836,N_214);
or U5360 (N_5360,N_4989,N_602);
and U5361 (N_5361,N_215,N_299);
nand U5362 (N_5362,N_4870,N_1980);
nor U5363 (N_5363,N_829,N_3912);
nand U5364 (N_5364,N_3974,N_4955);
and U5365 (N_5365,N_2373,N_2828);
nand U5366 (N_5366,N_1535,N_1191);
nor U5367 (N_5367,N_2101,N_3864);
or U5368 (N_5368,N_2231,N_4124);
or U5369 (N_5369,N_2028,N_1111);
or U5370 (N_5370,N_1808,N_480);
or U5371 (N_5371,N_2003,N_82);
nor U5372 (N_5372,N_649,N_550);
nor U5373 (N_5373,N_4010,N_3853);
and U5374 (N_5374,N_1498,N_3872);
nand U5375 (N_5375,N_293,N_2964);
nand U5376 (N_5376,N_3265,N_1366);
nor U5377 (N_5377,N_3084,N_3575);
nor U5378 (N_5378,N_4076,N_4592);
or U5379 (N_5379,N_3153,N_2499);
or U5380 (N_5380,N_2396,N_490);
and U5381 (N_5381,N_1302,N_2796);
nor U5382 (N_5382,N_1167,N_4696);
and U5383 (N_5383,N_3207,N_66);
nor U5384 (N_5384,N_1847,N_2757);
or U5385 (N_5385,N_3866,N_988);
or U5386 (N_5386,N_2492,N_304);
and U5387 (N_5387,N_1487,N_2380);
and U5388 (N_5388,N_1105,N_1543);
and U5389 (N_5389,N_3529,N_2423);
or U5390 (N_5390,N_4288,N_4635);
nor U5391 (N_5391,N_1201,N_2351);
or U5392 (N_5392,N_1325,N_1102);
xnor U5393 (N_5393,N_2694,N_1997);
nand U5394 (N_5394,N_2265,N_3638);
nor U5395 (N_5395,N_1319,N_67);
nor U5396 (N_5396,N_4019,N_3010);
nand U5397 (N_5397,N_4712,N_1897);
nand U5398 (N_5398,N_1365,N_4706);
nand U5399 (N_5399,N_3745,N_2923);
and U5400 (N_5400,N_3218,N_746);
nor U5401 (N_5401,N_69,N_1921);
nand U5402 (N_5402,N_2738,N_1133);
or U5403 (N_5403,N_3073,N_1698);
and U5404 (N_5404,N_4249,N_4576);
and U5405 (N_5405,N_2934,N_53);
and U5406 (N_5406,N_3931,N_185);
nor U5407 (N_5407,N_2607,N_4154);
nand U5408 (N_5408,N_402,N_1062);
and U5409 (N_5409,N_1041,N_4067);
nand U5410 (N_5410,N_3411,N_1528);
or U5411 (N_5411,N_2193,N_1974);
or U5412 (N_5412,N_3379,N_347);
nand U5413 (N_5413,N_1195,N_4307);
nor U5414 (N_5414,N_4749,N_1995);
and U5415 (N_5415,N_4732,N_1724);
nor U5416 (N_5416,N_132,N_1377);
or U5417 (N_5417,N_380,N_3258);
and U5418 (N_5418,N_3362,N_3020);
and U5419 (N_5419,N_1227,N_2128);
nand U5420 (N_5420,N_1110,N_1703);
xor U5421 (N_5421,N_1101,N_4162);
or U5422 (N_5422,N_3590,N_3040);
and U5423 (N_5423,N_4555,N_1010);
and U5424 (N_5424,N_4259,N_2033);
and U5425 (N_5425,N_3820,N_2978);
nor U5426 (N_5426,N_1029,N_3577);
nor U5427 (N_5427,N_3576,N_1254);
nand U5428 (N_5428,N_4986,N_4947);
and U5429 (N_5429,N_2439,N_1436);
nor U5430 (N_5430,N_3300,N_691);
and U5431 (N_5431,N_3983,N_1116);
xnor U5432 (N_5432,N_2799,N_465);
and U5433 (N_5433,N_751,N_2759);
and U5434 (N_5434,N_2132,N_4020);
nand U5435 (N_5435,N_263,N_549);
nor U5436 (N_5436,N_255,N_3253);
nand U5437 (N_5437,N_1516,N_1257);
nor U5438 (N_5438,N_1173,N_3925);
nand U5439 (N_5439,N_767,N_1135);
nand U5440 (N_5440,N_4031,N_2844);
and U5441 (N_5441,N_2200,N_4737);
nor U5442 (N_5442,N_4188,N_1592);
nor U5443 (N_5443,N_4292,N_4505);
nor U5444 (N_5444,N_3029,N_1766);
nor U5445 (N_5445,N_4330,N_4539);
or U5446 (N_5446,N_509,N_79);
nand U5447 (N_5447,N_1745,N_976);
nand U5448 (N_5448,N_2726,N_4403);
or U5449 (N_5449,N_2705,N_520);
and U5450 (N_5450,N_3458,N_3641);
nand U5451 (N_5451,N_3424,N_274);
and U5452 (N_5452,N_4977,N_3087);
nor U5453 (N_5453,N_2912,N_4011);
nor U5454 (N_5454,N_3390,N_2279);
nor U5455 (N_5455,N_3168,N_1217);
nor U5456 (N_5456,N_2247,N_802);
nor U5457 (N_5457,N_757,N_737);
or U5458 (N_5458,N_3223,N_3476);
nand U5459 (N_5459,N_1694,N_1156);
nand U5460 (N_5460,N_2150,N_1371);
nand U5461 (N_5461,N_2124,N_1051);
or U5462 (N_5462,N_3988,N_943);
or U5463 (N_5463,N_2800,N_1671);
and U5464 (N_5464,N_721,N_965);
nor U5465 (N_5465,N_1421,N_195);
or U5466 (N_5466,N_3259,N_3750);
nor U5467 (N_5467,N_4611,N_719);
or U5468 (N_5468,N_920,N_4337);
or U5469 (N_5469,N_4702,N_3893);
nor U5470 (N_5470,N_2239,N_2735);
nand U5471 (N_5471,N_3232,N_3770);
xor U5472 (N_5472,N_321,N_3256);
nor U5473 (N_5473,N_545,N_308);
and U5474 (N_5474,N_1691,N_4768);
nand U5475 (N_5475,N_3682,N_834);
or U5476 (N_5476,N_640,N_2263);
and U5477 (N_5477,N_2325,N_3456);
or U5478 (N_5478,N_2429,N_196);
and U5479 (N_5479,N_3143,N_3483);
nand U5480 (N_5480,N_3314,N_1719);
nor U5481 (N_5481,N_682,N_1028);
nor U5482 (N_5482,N_3661,N_40);
and U5483 (N_5483,N_1937,N_3858);
or U5484 (N_5484,N_3648,N_3846);
nand U5485 (N_5485,N_444,N_3052);
and U5486 (N_5486,N_968,N_4041);
and U5487 (N_5487,N_2134,N_1548);
nand U5488 (N_5488,N_323,N_4636);
nand U5489 (N_5489,N_2352,N_142);
and U5490 (N_5490,N_1812,N_2254);
or U5491 (N_5491,N_3485,N_2971);
or U5492 (N_5492,N_4825,N_724);
nor U5493 (N_5493,N_2075,N_2294);
or U5494 (N_5494,N_710,N_4598);
and U5495 (N_5495,N_3910,N_3184);
nor U5496 (N_5496,N_383,N_3308);
nor U5497 (N_5497,N_2498,N_3280);
nor U5498 (N_5498,N_1925,N_4179);
nor U5499 (N_5499,N_1233,N_4096);
and U5500 (N_5500,N_315,N_4881);
and U5501 (N_5501,N_3043,N_1244);
and U5502 (N_5502,N_357,N_3320);
nor U5503 (N_5503,N_4974,N_2210);
and U5504 (N_5504,N_302,N_1865);
or U5505 (N_5505,N_25,N_1376);
and U5506 (N_5506,N_2602,N_3078);
or U5507 (N_5507,N_2902,N_3501);
nand U5508 (N_5508,N_3117,N_1050);
and U5509 (N_5509,N_1608,N_322);
and U5510 (N_5510,N_975,N_2708);
or U5511 (N_5511,N_696,N_4);
and U5512 (N_5512,N_1011,N_4987);
and U5513 (N_5513,N_1947,N_479);
and U5514 (N_5514,N_4993,N_404);
or U5515 (N_5515,N_726,N_2950);
and U5516 (N_5516,N_3584,N_1247);
nand U5517 (N_5517,N_76,N_2523);
nand U5518 (N_5518,N_3964,N_4303);
or U5519 (N_5519,N_314,N_3706);
and U5520 (N_5520,N_591,N_1085);
xor U5521 (N_5521,N_348,N_2107);
or U5522 (N_5522,N_1200,N_4419);
and U5523 (N_5523,N_4028,N_386);
nor U5524 (N_5524,N_3804,N_1828);
and U5525 (N_5525,N_422,N_1412);
nand U5526 (N_5526,N_2561,N_2496);
and U5527 (N_5527,N_1710,N_3631);
nand U5528 (N_5528,N_3694,N_2615);
nand U5529 (N_5529,N_180,N_4942);
nor U5530 (N_5530,N_476,N_2486);
and U5531 (N_5531,N_1840,N_110);
nor U5532 (N_5532,N_1524,N_675);
nand U5533 (N_5533,N_328,N_1706);
or U5534 (N_5534,N_3718,N_1343);
and U5535 (N_5535,N_1206,N_994);
nand U5536 (N_5536,N_2577,N_2381);
or U5537 (N_5537,N_2355,N_1760);
nor U5538 (N_5538,N_3807,N_3474);
and U5539 (N_5539,N_1130,N_4077);
nand U5540 (N_5540,N_734,N_4431);
and U5541 (N_5541,N_4430,N_1869);
nand U5542 (N_5542,N_1036,N_2566);
and U5543 (N_5543,N_4981,N_1137);
and U5544 (N_5544,N_914,N_2774);
and U5545 (N_5545,N_1456,N_1680);
nor U5546 (N_5546,N_1849,N_2675);
nor U5547 (N_5547,N_3651,N_198);
and U5548 (N_5548,N_3493,N_3098);
or U5549 (N_5549,N_1112,N_252);
nand U5550 (N_5550,N_2990,N_1518);
or U5551 (N_5551,N_4086,N_429);
nand U5552 (N_5552,N_1305,N_4385);
nand U5553 (N_5553,N_3240,N_4577);
or U5554 (N_5554,N_2921,N_2074);
and U5555 (N_5555,N_783,N_2948);
or U5556 (N_5556,N_957,N_1693);
or U5557 (N_5557,N_4192,N_1186);
nand U5558 (N_5558,N_4767,N_2576);
and U5559 (N_5559,N_713,N_1400);
or U5560 (N_5560,N_2430,N_795);
or U5561 (N_5561,N_4772,N_1837);
nand U5562 (N_5562,N_868,N_2637);
nand U5563 (N_5563,N_3678,N_2245);
and U5564 (N_5564,N_641,N_3382);
or U5565 (N_5565,N_4186,N_569);
nor U5566 (N_5566,N_887,N_2625);
nor U5567 (N_5567,N_3595,N_2120);
nor U5568 (N_5568,N_4628,N_530);
nor U5569 (N_5569,N_3323,N_3650);
and U5570 (N_5570,N_3195,N_3579);
and U5571 (N_5571,N_2297,N_1733);
nand U5572 (N_5572,N_2977,N_2724);
and U5573 (N_5573,N_2614,N_2010);
nor U5574 (N_5574,N_2483,N_2507);
nor U5575 (N_5575,N_647,N_3262);
nand U5576 (N_5576,N_4757,N_2400);
and U5577 (N_5577,N_1576,N_3247);
or U5578 (N_5578,N_4932,N_4639);
or U5579 (N_5579,N_1347,N_2858);
nand U5580 (N_5580,N_4658,N_15);
and U5581 (N_5581,N_3522,N_615);
and U5582 (N_5582,N_431,N_4734);
nor U5583 (N_5583,N_3475,N_1689);
nand U5584 (N_5584,N_3511,N_494);
and U5585 (N_5585,N_192,N_1282);
and U5586 (N_5586,N_1272,N_847);
or U5587 (N_5587,N_3979,N_3505);
nand U5588 (N_5588,N_1391,N_1374);
or U5589 (N_5589,N_2015,N_3345);
and U5590 (N_5590,N_1811,N_1707);
nand U5591 (N_5591,N_1,N_1493);
and U5592 (N_5592,N_2391,N_33);
xor U5593 (N_5593,N_4516,N_2397);
nand U5594 (N_5594,N_1386,N_4123);
nand U5595 (N_5595,N_442,N_4262);
or U5596 (N_5596,N_1093,N_4861);
or U5597 (N_5597,N_1108,N_1894);
nor U5598 (N_5598,N_151,N_2755);
nor U5599 (N_5599,N_4632,N_2234);
nand U5600 (N_5600,N_1824,N_4057);
nor U5601 (N_5601,N_3385,N_3427);
nand U5602 (N_5602,N_2823,N_368);
nor U5603 (N_5603,N_2070,N_908);
nor U5604 (N_5604,N_3904,N_4038);
nor U5605 (N_5605,N_3567,N_1582);
and U5606 (N_5606,N_820,N_460);
or U5607 (N_5607,N_394,N_2291);
or U5608 (N_5608,N_1134,N_4869);
nor U5609 (N_5609,N_1914,N_3026);
or U5610 (N_5610,N_456,N_4953);
or U5611 (N_5611,N_446,N_4282);
or U5612 (N_5612,N_4522,N_4388);
and U5613 (N_5613,N_223,N_18);
nand U5614 (N_5614,N_3046,N_1370);
nor U5615 (N_5615,N_278,N_1118);
or U5616 (N_5616,N_4850,N_178);
nor U5617 (N_5617,N_3354,N_4766);
and U5618 (N_5618,N_1590,N_2667);
or U5619 (N_5619,N_3535,N_4804);
and U5620 (N_5620,N_772,N_1153);
nor U5621 (N_5621,N_1005,N_4418);
and U5622 (N_5622,N_2859,N_1850);
or U5623 (N_5623,N_199,N_3972);
nand U5624 (N_5624,N_2712,N_4528);
nand U5625 (N_5625,N_3202,N_3513);
or U5626 (N_5626,N_2224,N_2307);
nand U5627 (N_5627,N_1857,N_2094);
and U5628 (N_5628,N_2139,N_4640);
or U5629 (N_5629,N_3690,N_723);
and U5630 (N_5630,N_504,N_4473);
or U5631 (N_5631,N_1932,N_4298);
nor U5632 (N_5632,N_1678,N_499);
nor U5633 (N_5633,N_1190,N_3882);
nand U5634 (N_5634,N_4369,N_4748);
or U5635 (N_5635,N_1158,N_4275);
nand U5636 (N_5636,N_3238,N_1615);
nand U5637 (N_5637,N_4280,N_4823);
and U5638 (N_5638,N_3924,N_4176);
or U5639 (N_5639,N_1984,N_3680);
nand U5640 (N_5640,N_1722,N_2444);
nor U5641 (N_5641,N_3626,N_2946);
nor U5642 (N_5642,N_4838,N_3321);
xor U5643 (N_5643,N_1350,N_2020);
and U5644 (N_5644,N_658,N_1983);
or U5645 (N_5645,N_4061,N_373);
and U5646 (N_5646,N_2411,N_951);
or U5647 (N_5647,N_4297,N_1422);
and U5648 (N_5648,N_3150,N_3586);
or U5649 (N_5649,N_4368,N_2634);
nand U5650 (N_5650,N_1237,N_2727);
nand U5651 (N_5651,N_2770,N_2221);
nor U5652 (N_5652,N_4678,N_432);
nor U5653 (N_5653,N_4571,N_2218);
nand U5654 (N_5654,N_3786,N_2692);
nand U5655 (N_5655,N_1781,N_4251);
nand U5656 (N_5656,N_4971,N_3523);
or U5657 (N_5657,N_1773,N_1103);
nand U5658 (N_5658,N_2583,N_397);
or U5659 (N_5659,N_1196,N_1293);
nand U5660 (N_5660,N_806,N_3338);
nand U5661 (N_5661,N_4815,N_4172);
xnor U5662 (N_5662,N_1749,N_4996);
and U5663 (N_5663,N_1941,N_3938);
nor U5664 (N_5664,N_167,N_3099);
or U5665 (N_5665,N_529,N_1266);
or U5666 (N_5666,N_2131,N_1872);
nor U5667 (N_5667,N_3667,N_2804);
and U5668 (N_5668,N_2989,N_3674);
nand U5669 (N_5669,N_2725,N_1128);
or U5670 (N_5670,N_2750,N_24);
nand U5671 (N_5671,N_2821,N_964);
xor U5672 (N_5672,N_275,N_4286);
nor U5673 (N_5673,N_990,N_4811);
nor U5674 (N_5674,N_4441,N_1568);
nand U5675 (N_5675,N_1311,N_4225);
and U5676 (N_5676,N_2886,N_871);
nand U5677 (N_5677,N_4618,N_2617);
nand U5678 (N_5678,N_2361,N_2479);
or U5679 (N_5679,N_4336,N_924);
nand U5680 (N_5680,N_46,N_71);
or U5681 (N_5681,N_1610,N_2880);
and U5682 (N_5682,N_1711,N_1026);
nor U5683 (N_5683,N_1448,N_85);
nor U5684 (N_5684,N_1189,N_1742);
nand U5685 (N_5685,N_1231,N_2760);
xor U5686 (N_5686,N_3186,N_1643);
nand U5687 (N_5687,N_789,N_3208);
and U5688 (N_5688,N_2877,N_837);
nor U5689 (N_5689,N_2510,N_1417);
and U5690 (N_5690,N_370,N_3837);
and U5691 (N_5691,N_1297,N_3681);
and U5692 (N_5692,N_1451,N_2480);
and U5693 (N_5693,N_3758,N_1429);
or U5694 (N_5694,N_2406,N_708);
nand U5695 (N_5695,N_3656,N_2043);
nor U5696 (N_5696,N_2154,N_1076);
or U5697 (N_5697,N_123,N_1596);
nor U5698 (N_5698,N_3198,N_4695);
and U5699 (N_5699,N_2296,N_350);
and U5700 (N_5700,N_1019,N_2440);
nand U5701 (N_5701,N_3935,N_3654);
nor U5702 (N_5702,N_1458,N_4131);
nor U5703 (N_5703,N_1825,N_4694);
or U5704 (N_5704,N_4973,N_4198);
and U5705 (N_5705,N_1219,N_57);
nand U5706 (N_5706,N_2360,N_2169);
nand U5707 (N_5707,N_1623,N_2951);
nor U5708 (N_5708,N_2408,N_1411);
xor U5709 (N_5709,N_2311,N_4335);
nand U5710 (N_5710,N_3295,N_1757);
or U5711 (N_5711,N_872,N_1359);
xnor U5712 (N_5712,N_1777,N_3236);
and U5713 (N_5713,N_1425,N_3222);
nand U5714 (N_5714,N_1551,N_4447);
and U5715 (N_5715,N_1717,N_3336);
nor U5716 (N_5716,N_913,N_3124);
or U5717 (N_5717,N_4672,N_4381);
nor U5718 (N_5718,N_1564,N_2437);
nor U5719 (N_5719,N_3175,N_209);
and U5720 (N_5720,N_4952,N_4477);
and U5721 (N_5721,N_2269,N_4508);
or U5722 (N_5722,N_3865,N_4719);
and U5723 (N_5723,N_2876,N_693);
nand U5724 (N_5724,N_4845,N_1542);
nand U5725 (N_5725,N_4421,N_4574);
nand U5726 (N_5726,N_4374,N_4175);
nor U5727 (N_5727,N_4662,N_3142);
and U5728 (N_5728,N_4106,N_2092);
and U5729 (N_5729,N_4453,N_3264);
and U5730 (N_5730,N_4304,N_1991);
nand U5731 (N_5731,N_73,N_2795);
and U5732 (N_5732,N_680,N_4399);
nand U5733 (N_5733,N_1973,N_229);
and U5734 (N_5734,N_4142,N_1709);
nand U5735 (N_5735,N_1685,N_3917);
or U5736 (N_5736,N_2919,N_1405);
or U5737 (N_5737,N_3717,N_1539);
and U5738 (N_5738,N_4667,N_4151);
and U5739 (N_5739,N_2309,N_4843);
nor U5740 (N_5740,N_3604,N_3177);
or U5741 (N_5741,N_2824,N_2428);
or U5742 (N_5742,N_3103,N_1994);
nor U5743 (N_5743,N_2478,N_4305);
nand U5744 (N_5744,N_4828,N_292);
or U5745 (N_5745,N_3270,N_3730);
nand U5746 (N_5746,N_1918,N_2895);
nor U5747 (N_5747,N_600,N_4497);
nand U5748 (N_5748,N_4554,N_2145);
and U5749 (N_5749,N_2117,N_3796);
nand U5750 (N_5750,N_894,N_727);
or U5751 (N_5751,N_2370,N_3932);
nand U5752 (N_5752,N_1851,N_1225);
and U5753 (N_5753,N_862,N_247);
or U5754 (N_5754,N_2412,N_3776);
nor U5755 (N_5755,N_3683,N_773);
xnor U5756 (N_5756,N_2461,N_4818);
nand U5757 (N_5757,N_2061,N_1942);
and U5758 (N_5758,N_2472,N_1432);
and U5759 (N_5759,N_2870,N_3693);
and U5760 (N_5760,N_4378,N_2573);
nand U5761 (N_5761,N_4460,N_3862);
or U5762 (N_5762,N_4156,N_3532);
nor U5763 (N_5763,N_3571,N_483);
nor U5764 (N_5764,N_3937,N_1321);
nor U5765 (N_5765,N_2749,N_4071);
nor U5766 (N_5766,N_3756,N_1462);
nor U5767 (N_5767,N_1226,N_2717);
and U5768 (N_5768,N_4594,N_3843);
nor U5769 (N_5769,N_935,N_4500);
or U5770 (N_5770,N_521,N_1818);
nand U5771 (N_5771,N_10,N_880);
nor U5772 (N_5772,N_2049,N_2589);
xnor U5773 (N_5773,N_3340,N_1534);
and U5774 (N_5774,N_3002,N_437);
or U5775 (N_5775,N_3663,N_2651);
nand U5776 (N_5776,N_2840,N_3426);
and U5777 (N_5777,N_2209,N_2890);
and U5778 (N_5778,N_51,N_3226);
and U5779 (N_5779,N_2217,N_1939);
nand U5780 (N_5780,N_4509,N_1896);
xor U5781 (N_5781,N_4868,N_2022);
xor U5782 (N_5782,N_537,N_372);
nor U5783 (N_5783,N_896,N_367);
or U5784 (N_5784,N_3225,N_2385);
or U5785 (N_5785,N_3415,N_4032);
or U5786 (N_5786,N_1780,N_4174);
or U5787 (N_5787,N_3611,N_4990);
or U5788 (N_5788,N_4095,N_4629);
nor U5789 (N_5789,N_4540,N_1139);
or U5790 (N_5790,N_582,N_3923);
nor U5791 (N_5791,N_518,N_4988);
nor U5792 (N_5792,N_248,N_3790);
and U5793 (N_5793,N_1384,N_3902);
xnor U5794 (N_5794,N_4802,N_1519);
nor U5795 (N_5795,N_4948,N_3545);
and U5796 (N_5796,N_4538,N_1888);
nand U5797 (N_5797,N_2513,N_2849);
or U5798 (N_5798,N_2109,N_3635);
nand U5799 (N_5799,N_1526,N_2631);
nor U5800 (N_5800,N_1591,N_484);
nand U5801 (N_5801,N_3334,N_3085);
or U5802 (N_5802,N_1913,N_1150);
or U5803 (N_5803,N_2185,N_3987);
nand U5804 (N_5804,N_4504,N_1043);
or U5805 (N_5805,N_2197,N_242);
or U5806 (N_5806,N_4494,N_1000);
nor U5807 (N_5807,N_3708,N_4553);
and U5808 (N_5808,N_2767,N_3617);
or U5809 (N_5809,N_49,N_488);
and U5810 (N_5810,N_850,N_1113);
nand U5811 (N_5811,N_4703,N_4281);
nand U5812 (N_5812,N_277,N_4542);
nor U5813 (N_5813,N_3341,N_3534);
and U5814 (N_5814,N_3856,N_469);
or U5815 (N_5815,N_4214,N_4065);
or U5816 (N_5816,N_4034,N_4559);
or U5817 (N_5817,N_4340,N_440);
and U5818 (N_5818,N_4894,N_3803);
xnor U5819 (N_5819,N_4548,N_714);
and U5820 (N_5820,N_835,N_4463);
nor U5821 (N_5821,N_3307,N_1250);
nand U5822 (N_5822,N_177,N_1270);
nand U5823 (N_5823,N_4361,N_1866);
nand U5824 (N_5824,N_2864,N_2235);
nor U5825 (N_5825,N_140,N_2158);
nor U5826 (N_5826,N_4796,N_4260);
nand U5827 (N_5827,N_949,N_4191);
and U5828 (N_5828,N_3946,N_901);
or U5829 (N_5829,N_1802,N_1816);
nand U5830 (N_5830,N_4242,N_2700);
or U5831 (N_5831,N_2443,N_3224);
or U5832 (N_5832,N_3044,N_3241);
or U5833 (N_5833,N_2756,N_4885);
and U5834 (N_5834,N_3782,N_1605);
and U5835 (N_5835,N_377,N_1839);
nand U5836 (N_5836,N_4917,N_2863);
nor U5837 (N_5837,N_4180,N_2967);
nor U5838 (N_5838,N_3154,N_3355);
nor U5839 (N_5839,N_4582,N_1541);
or U5840 (N_5840,N_1527,N_2636);
or U5841 (N_5841,N_740,N_3830);
nand U5842 (N_5842,N_4564,N_13);
and U5843 (N_5843,N_2426,N_554);
nor U5844 (N_5844,N_4829,N_1269);
or U5845 (N_5845,N_1123,N_3357);
nor U5846 (N_5846,N_3205,N_2746);
nand U5847 (N_5847,N_1683,N_2587);
or U5848 (N_5848,N_4197,N_4898);
or U5849 (N_5849,N_1520,N_4022);
and U5850 (N_5850,N_4212,N_3652);
nor U5851 (N_5851,N_2340,N_2267);
nand U5852 (N_5852,N_1170,N_2350);
nor U5853 (N_5853,N_3075,N_2754);
nor U5854 (N_5854,N_2747,N_2374);
nand U5855 (N_5855,N_1248,N_1624);
or U5856 (N_5856,N_206,N_2178);
and U5857 (N_5857,N_4914,N_4707);
or U5858 (N_5858,N_3921,N_1695);
or U5859 (N_5859,N_1967,N_3639);
or U5860 (N_5860,N_3550,N_4750);
nor U5861 (N_5861,N_4392,N_1234);
nor U5862 (N_5862,N_4333,N_307);
nor U5863 (N_5863,N_1759,N_2215);
nor U5864 (N_5864,N_2812,N_4153);
or U5865 (N_5865,N_4464,N_1957);
nand U5866 (N_5866,N_2040,N_4411);
nor U5867 (N_5867,N_4912,N_3140);
nor U5868 (N_5868,N_4492,N_3670);
or U5869 (N_5869,N_4137,N_3814);
or U5870 (N_5870,N_4435,N_3985);
and U5871 (N_5871,N_3530,N_4994);
or U5872 (N_5872,N_3773,N_1619);
nor U5873 (N_5873,N_3387,N_4690);
nor U5874 (N_5874,N_3297,N_1120);
or U5875 (N_5875,N_2330,N_3737);
and U5876 (N_5876,N_267,N_4243);
nand U5877 (N_5877,N_2055,N_2119);
or U5878 (N_5878,N_313,N_1806);
and U5879 (N_5879,N_2206,N_2062);
nand U5880 (N_5880,N_4118,N_3368);
nor U5881 (N_5881,N_3045,N_2782);
or U5882 (N_5882,N_1362,N_666);
nand U5883 (N_5883,N_1595,N_1909);
nand U5884 (N_5884,N_2138,N_1986);
nand U5885 (N_5885,N_165,N_2762);
nor U5886 (N_5886,N_1638,N_2697);
nand U5887 (N_5887,N_316,N_2303);
and U5888 (N_5888,N_4417,N_4700);
and U5889 (N_5889,N_276,N_96);
and U5890 (N_5890,N_4614,N_1779);
nor U5891 (N_5891,N_624,N_3176);
nor U5892 (N_5892,N_4003,N_4759);
and U5893 (N_5893,N_2686,N_4888);
or U5894 (N_5894,N_272,N_1558);
and U5895 (N_5895,N_1203,N_2761);
nor U5896 (N_5896,N_2659,N_2456);
nand U5897 (N_5897,N_4992,N_3655);
nand U5898 (N_5898,N_4687,N_996);
nor U5899 (N_5899,N_923,N_27);
nor U5900 (N_5900,N_4079,N_1646);
or U5901 (N_5901,N_2856,N_208);
nand U5902 (N_5902,N_4144,N_581);
or U5903 (N_5903,N_1492,N_2647);
nand U5904 (N_5904,N_2310,N_3780);
or U5905 (N_5905,N_2730,N_4401);
or U5906 (N_5906,N_453,N_2813);
nor U5907 (N_5907,N_4819,N_130);
or U5908 (N_5908,N_169,N_3630);
nor U5909 (N_5909,N_2039,N_2367);
and U5910 (N_5910,N_1522,N_4817);
nand U5911 (N_5911,N_1438,N_3128);
nor U5912 (N_5912,N_3139,N_2349);
and U5913 (N_5913,N_2687,N_542);
nand U5914 (N_5914,N_2819,N_1132);
nand U5915 (N_5915,N_174,N_3146);
nand U5916 (N_5916,N_3468,N_4455);
nand U5917 (N_5917,N_269,N_2807);
or U5918 (N_5918,N_4793,N_697);
and U5919 (N_5919,N_3995,N_1723);
or U5920 (N_5920,N_2171,N_1437);
or U5921 (N_5921,N_4600,N_4139);
and U5922 (N_5922,N_4353,N_2416);
or U5923 (N_5923,N_1361,N_2563);
nor U5924 (N_5924,N_1300,N_4048);
or U5925 (N_5925,N_1686,N_3404);
nand U5926 (N_5926,N_3959,N_3144);
and U5927 (N_5927,N_770,N_359);
and U5928 (N_5928,N_4466,N_296);
or U5929 (N_5929,N_4213,N_1466);
nor U5930 (N_5930,N_2772,N_1408);
or U5931 (N_5931,N_4921,N_1741);
nor U5932 (N_5932,N_4884,N_4351);
nor U5933 (N_5933,N_2096,N_879);
nand U5934 (N_5934,N_204,N_3489);
and U5935 (N_5935,N_1369,N_4813);
nand U5936 (N_5936,N_361,N_592);
and U5937 (N_5937,N_11,N_4146);
or U5938 (N_5938,N_4265,N_1912);
or U5939 (N_5939,N_3325,N_4462);
nand U5940 (N_5940,N_4088,N_4788);
nand U5941 (N_5941,N_2468,N_4486);
nor U5942 (N_5942,N_65,N_2940);
nand U5943 (N_5943,N_279,N_3460);
or U5944 (N_5944,N_4127,N_1192);
or U5945 (N_5945,N_2276,N_3919);
nand U5946 (N_5946,N_416,N_2862);
or U5947 (N_5947,N_907,N_4239);
nand U5948 (N_5948,N_1906,N_4294);
and U5949 (N_5949,N_763,N_621);
nor U5950 (N_5950,N_939,N_523);
nand U5951 (N_5951,N_1890,N_2112);
or U5952 (N_5952,N_4533,N_270);
nand U5953 (N_5953,N_1853,N_4487);
and U5954 (N_5954,N_560,N_2781);
and U5955 (N_5955,N_2387,N_2685);
nand U5956 (N_5956,N_1164,N_493);
nand U5957 (N_5957,N_962,N_3785);
or U5958 (N_5958,N_3699,N_4910);
nor U5959 (N_5959,N_93,N_2958);
and U5960 (N_5960,N_3378,N_4451);
nor U5961 (N_5961,N_2993,N_4923);
nor U5962 (N_5962,N_4668,N_2108);
or U5963 (N_5963,N_794,N_637);
and U5964 (N_5964,N_379,N_398);
xor U5965 (N_5965,N_4995,N_888);
nand U5966 (N_5966,N_3841,N_1020);
nand U5967 (N_5967,N_3331,N_3999);
and U5968 (N_5968,N_3907,N_2230);
nor U5969 (N_5969,N_1469,N_3875);
nand U5970 (N_5970,N_408,N_1523);
or U5971 (N_5971,N_423,N_395);
or U5972 (N_5972,N_160,N_449);
and U5973 (N_5973,N_3105,N_497);
or U5974 (N_5974,N_60,N_522);
nor U5975 (N_5975,N_532,N_4082);
and U5976 (N_5976,N_4688,N_1922);
nand U5977 (N_5977,N_2564,N_3055);
nand U5978 (N_5978,N_4860,N_1107);
and U5979 (N_5979,N_4148,N_4316);
nor U5980 (N_5980,N_3982,N_4909);
nor U5981 (N_5981,N_1578,N_2463);
nand U5982 (N_5982,N_3941,N_3625);
and U5983 (N_5983,N_4452,N_3679);
nor U5984 (N_5984,N_987,N_4114);
nor U5985 (N_5985,N_4836,N_3243);
nand U5986 (N_5986,N_1772,N_80);
nand U5987 (N_5987,N_1517,N_3193);
or U5988 (N_5988,N_4183,N_2012);
and U5989 (N_5989,N_4256,N_2025);
nand U5990 (N_5990,N_3047,N_3819);
and U5991 (N_5991,N_3324,N_2929);
nor U5992 (N_5992,N_1002,N_3313);
or U5993 (N_5993,N_2451,N_4511);
nand U5994 (N_5994,N_3242,N_3145);
and U5995 (N_5995,N_3729,N_64);
or U5996 (N_5996,N_2222,N_2180);
and U5997 (N_5997,N_1968,N_4795);
and U5998 (N_5998,N_2834,N_4892);
or U5999 (N_5999,N_2935,N_748);
nor U6000 (N_6000,N_3180,N_4875);
nor U6001 (N_6001,N_4620,N_674);
nand U6002 (N_6002,N_3665,N_2829);
or U6003 (N_6003,N_4040,N_3832);
nor U6004 (N_6004,N_1484,N_1513);
or U6005 (N_6005,N_531,N_3509);
and U6006 (N_6006,N_4208,N_301);
or U6007 (N_6007,N_3032,N_63);
nand U6008 (N_6008,N_1086,N_2076);
nand U6009 (N_6009,N_915,N_4223);
and U6010 (N_6010,N_3713,N_4203);
nand U6011 (N_6011,N_4006,N_3732);
nand U6012 (N_6012,N_738,N_4446);
and U6013 (N_6013,N_609,N_3138);
or U6014 (N_6014,N_19,N_4774);
or U6015 (N_6015,N_2500,N_1031);
and U6016 (N_6016,N_1985,N_4471);
or U6017 (N_6017,N_3276,N_147);
and U6018 (N_6018,N_2050,N_4631);
nor U6019 (N_6019,N_926,N_1804);
or U6020 (N_6020,N_3001,N_2005);
nand U6021 (N_6021,N_1439,N_1490);
nand U6022 (N_6022,N_1908,N_4727);
nand U6023 (N_6023,N_4943,N_3416);
nor U6024 (N_6024,N_4269,N_2388);
and U6025 (N_6025,N_1856,N_3502);
or U6026 (N_6026,N_1637,N_4847);
or U6027 (N_6027,N_3498,N_4601);
nand U6028 (N_6028,N_2487,N_3878);
nor U6029 (N_6029,N_3936,N_3299);
or U6030 (N_6030,N_4358,N_44);
or U6031 (N_6031,N_1211,N_365);
nor U6032 (N_6032,N_4479,N_4220);
xor U6033 (N_6033,N_172,N_657);
nand U6034 (N_6034,N_1367,N_3417);
nor U6035 (N_6035,N_1611,N_910);
nor U6036 (N_6036,N_1622,N_245);
and U6037 (N_6037,N_3848,N_424);
nor U6038 (N_6038,N_1537,N_1813);
nand U6039 (N_6039,N_163,N_4755);
and U6040 (N_6040,N_4459,N_1732);
nor U6041 (N_6041,N_1276,N_2873);
and U6042 (N_6042,N_271,N_3443);
and U6043 (N_6043,N_4194,N_1768);
nor U6044 (N_6044,N_4215,N_1944);
nand U6045 (N_6045,N_1788,N_312);
xnor U6046 (N_6046,N_2560,N_141);
nor U6047 (N_6047,N_3722,N_3343);
nand U6048 (N_6048,N_2632,N_3137);
nand U6049 (N_6049,N_445,N_2314);
nand U6050 (N_6050,N_2201,N_1278);
nor U6051 (N_6051,N_4141,N_4519);
or U6052 (N_6052,N_4740,N_3478);
nand U6053 (N_6053,N_3649,N_1271);
nor U6054 (N_6054,N_725,N_2994);
and U6055 (N_6055,N_2869,N_547);
nor U6056 (N_6056,N_1264,N_3836);
or U6057 (N_6057,N_3388,N_2359);
and U6058 (N_6058,N_1860,N_2526);
nor U6059 (N_6059,N_3261,N_809);
nor U6060 (N_6060,N_1716,N_2284);
nand U6061 (N_6061,N_159,N_2835);
and U6062 (N_6062,N_2715,N_1081);
and U6063 (N_6063,N_1791,N_1390);
or U6064 (N_6064,N_1929,N_893);
xnor U6065 (N_6065,N_426,N_2395);
nor U6066 (N_6066,N_698,N_2925);
nand U6067 (N_6067,N_1160,N_3437);
nor U6068 (N_6068,N_3503,N_2928);
and U6069 (N_6069,N_2601,N_4204);
or U6070 (N_6070,N_1826,N_4891);
or U6071 (N_6071,N_2136,N_664);
or U6072 (N_6072,N_104,N_4078);
or U6073 (N_6073,N_3288,N_3620);
nand U6074 (N_6074,N_4122,N_2662);
and U6075 (N_6075,N_632,N_1125);
or U6076 (N_6076,N_3899,N_3801);
nor U6077 (N_6077,N_3213,N_3578);
nand U6078 (N_6078,N_4524,N_3870);
and U6079 (N_6079,N_295,N_191);
nand U6080 (N_6080,N_1033,N_1322);
xor U6081 (N_6081,N_4866,N_4954);
nor U6082 (N_6082,N_4960,N_3149);
or U6083 (N_6083,N_3668,N_133);
and U6084 (N_6084,N_688,N_4780);
nand U6085 (N_6085,N_1212,N_4854);
or U6086 (N_6086,N_611,N_2972);
nor U6087 (N_6087,N_203,N_4018);
or U6088 (N_6088,N_3645,N_2626);
nand U6089 (N_6089,N_3521,N_2184);
nor U6090 (N_6090,N_3003,N_4025);
nor U6091 (N_6091,N_2790,N_931);
nand U6092 (N_6092,N_4797,N_1827);
nor U6093 (N_6093,N_2995,N_4052);
and U6094 (N_6094,N_4373,N_1911);
nand U6095 (N_6095,N_627,N_3539);
or U6096 (N_6096,N_3486,N_3556);
and U6097 (N_6097,N_2207,N_4824);
nor U6098 (N_6098,N_3452,N_1648);
and U6099 (N_6099,N_4299,N_3152);
nand U6100 (N_6100,N_3621,N_1069);
and U6101 (N_6101,N_3080,N_2295);
and U6102 (N_6102,N_1838,N_2794);
and U6103 (N_6103,N_2161,N_1634);
or U6104 (N_6104,N_3204,N_544);
and U6105 (N_6105,N_1335,N_2219);
and U6106 (N_6106,N_119,N_902);
or U6107 (N_6107,N_175,N_4177);
or U6108 (N_6108,N_3185,N_3346);
nand U6109 (N_6109,N_4902,N_4998);
nand U6110 (N_6110,N_960,N_1880);
or U6111 (N_6111,N_3191,N_3201);
or U6112 (N_6112,N_4822,N_21);
and U6113 (N_6113,N_614,N_4107);
or U6114 (N_6114,N_4352,N_4240);
and U6115 (N_6115,N_236,N_2551);
or U6116 (N_6116,N_2586,N_4903);
nand U6117 (N_6117,N_3450,N_1148);
and U6118 (N_6118,N_3463,N_689);
or U6119 (N_6119,N_3494,N_4609);
nand U6120 (N_6120,N_2153,N_1094);
and U6121 (N_6121,N_1565,N_2274);
nor U6122 (N_6122,N_4450,N_1497);
nor U6123 (N_6123,N_2907,N_280);
or U6124 (N_6124,N_2458,N_1761);
or U6125 (N_6125,N_4728,N_2343);
nand U6126 (N_6126,N_362,N_3419);
and U6127 (N_6127,N_679,N_3170);
nand U6128 (N_6128,N_2445,N_2372);
or U6129 (N_6129,N_4731,N_349);
and U6130 (N_6130,N_1952,N_4730);
nor U6131 (N_6131,N_2130,N_4169);
nor U6132 (N_6132,N_563,N_3653);
or U6133 (N_6133,N_2753,N_55);
nand U6134 (N_6134,N_4134,N_899);
nand U6135 (N_6135,N_2348,N_238);
nand U6136 (N_6136,N_1855,N_4587);
or U6137 (N_6137,N_1481,N_1640);
nand U6138 (N_6138,N_1794,N_2981);
and U6139 (N_6139,N_4621,N_590);
nand U6140 (N_6140,N_3497,N_3901);
nand U6141 (N_6141,N_2904,N_2857);
nand U6142 (N_6142,N_927,N_4393);
nand U6143 (N_6143,N_1127,N_1953);
and U6144 (N_6144,N_819,N_1955);
nor U6145 (N_6145,N_4365,N_4363);
nor U6146 (N_6146,N_4211,N_1599);
nor U6147 (N_6147,N_1829,N_2016);
and U6148 (N_6148,N_1499,N_1882);
nor U6149 (N_6149,N_2030,N_2522);
nand U6150 (N_6150,N_1987,N_3);
or U6151 (N_6151,N_2945,N_4193);
nor U6152 (N_6152,N_941,N_3167);
nor U6153 (N_6153,N_999,N_4043);
nor U6154 (N_6154,N_3194,N_701);
nor U6155 (N_6155,N_421,N_2106);
nand U6156 (N_6156,N_298,N_2228);
or U6157 (N_6157,N_1312,N_438);
nand U6158 (N_6158,N_4874,N_3822);
nand U6159 (N_6159,N_4207,N_3182);
or U6160 (N_6160,N_1016,N_843);
nor U6161 (N_6161,N_1221,N_4007);
nor U6162 (N_6162,N_556,N_4293);
and U6163 (N_6163,N_485,N_2357);
and U6164 (N_6164,N_4246,N_1044);
or U6165 (N_6165,N_1585,N_1265);
or U6166 (N_6166,N_2872,N_4790);
or U6167 (N_6167,N_2719,N_3061);
or U6168 (N_6168,N_3840,N_4321);
nand U6169 (N_6169,N_2419,N_4081);
nand U6170 (N_6170,N_588,N_4457);
nor U6171 (N_6171,N_3189,N_3892);
and U6172 (N_6172,N_2182,N_205);
nor U6173 (N_6173,N_2771,N_1392);
nand U6174 (N_6174,N_1751,N_107);
and U6175 (N_6175,N_4047,N_540);
nand U6176 (N_6176,N_409,N_781);
nand U6177 (N_6177,N_112,N_1059);
and U6178 (N_6178,N_3789,N_4936);
nor U6179 (N_6179,N_4698,N_1342);
nor U6180 (N_6180,N_3329,N_2327);
or U6181 (N_6181,N_3316,N_2924);
nand U6182 (N_6182,N_1844,N_4653);
xor U6183 (N_6183,N_2875,N_3121);
and U6184 (N_6184,N_1166,N_2888);
or U6185 (N_6185,N_2542,N_4415);
and U6186 (N_6186,N_291,N_1380);
nand U6187 (N_6187,N_4070,N_4597);
nand U6188 (N_6188,N_1383,N_1496);
and U6189 (N_6189,N_3488,N_3797);
nand U6190 (N_6190,N_3886,N_3598);
or U6191 (N_6191,N_950,N_3322);
or U6192 (N_6192,N_4287,N_287);
or U6193 (N_6193,N_4495,N_2833);
nand U6194 (N_6194,N_2943,N_718);
nor U6195 (N_6195,N_1399,N_3122);
or U6196 (N_6196,N_4366,N_4699);
xnor U6197 (N_6197,N_3009,N_2346);
or U6198 (N_6198,N_2598,N_2316);
or U6199 (N_6199,N_1945,N_4147);
and U6200 (N_6200,N_4315,N_2668);
nand U6201 (N_6201,N_4982,N_417);
or U6202 (N_6202,N_1373,N_2477);
nand U6203 (N_6203,N_143,N_1863);
nor U6204 (N_6204,N_566,N_3957);
nand U6205 (N_6205,N_3136,N_3311);
nor U6206 (N_6206,N_541,N_256);
and U6207 (N_6207,N_2392,N_4671);
nand U6208 (N_6208,N_2758,N_4270);
or U6209 (N_6209,N_840,N_4531);
nor U6210 (N_6210,N_330,N_4880);
nand U6211 (N_6211,N_3978,N_4426);
nor U6212 (N_6212,N_2280,N_3277);
nand U6213 (N_6213,N_3420,N_1891);
nor U6214 (N_6214,N_1533,N_327);
or U6215 (N_6215,N_3591,N_36);
or U6216 (N_6216,N_765,N_1954);
or U6217 (N_6217,N_2457,N_355);
nand U6218 (N_6218,N_4150,N_3200);
or U6219 (N_6219,N_4616,N_319);
nand U6220 (N_6220,N_1503,N_3615);
nor U6221 (N_6221,N_3051,N_598);
nor U6222 (N_6222,N_2784,N_234);
or U6223 (N_6223,N_2947,N_4878);
nor U6224 (N_6224,N_535,N_3454);
nor U6225 (N_6225,N_4480,N_3794);
or U6226 (N_6226,N_3888,N_478);
and U6227 (N_6227,N_3691,N_2874);
or U6228 (N_6228,N_346,N_4468);
or U6229 (N_6229,N_4372,N_2122);
or U6230 (N_6230,N_135,N_2474);
or U6231 (N_6231,N_1038,N_1594);
or U6232 (N_6232,N_2629,N_498);
and U6233 (N_6233,N_1799,N_4798);
nand U6234 (N_6234,N_1433,N_3421);
or U6235 (N_6235,N_634,N_29);
xnor U6236 (N_6236,N_814,N_427);
and U6237 (N_6237,N_3781,N_505);
or U6238 (N_6238,N_3504,N_597);
or U6239 (N_6239,N_1284,N_1259);
or U6240 (N_6240,N_1962,N_1982);
nand U6241 (N_6241,N_2090,N_4327);
nor U6242 (N_6242,N_2410,N_239);
and U6243 (N_6243,N_253,N_72);
or U6244 (N_6244,N_2699,N_4178);
nand U6245 (N_6245,N_2382,N_2778);
and U6246 (N_6246,N_1756,N_2537);
and U6247 (N_6247,N_854,N_4541);
nor U6248 (N_6248,N_1563,N_1509);
nand U6249 (N_6249,N_4930,N_1470);
or U6250 (N_6250,N_1705,N_3868);
and U6251 (N_6251,N_2378,N_533);
nand U6252 (N_6252,N_220,N_4663);
nor U6253 (N_6253,N_4354,N_3564);
nand U6254 (N_6254,N_1771,N_534);
nor U6255 (N_6255,N_4656,N_4754);
or U6256 (N_6256,N_2871,N_2788);
or U6257 (N_6257,N_52,N_2417);
and U6258 (N_6258,N_626,N_3573);
or U6259 (N_6259,N_477,N_1951);
nor U6260 (N_6260,N_703,N_2806);
or U6261 (N_6261,N_1290,N_4814);
or U6262 (N_6262,N_1966,N_474);
nand U6263 (N_6263,N_2232,N_1486);
or U6264 (N_6264,N_2949,N_1747);
nor U6265 (N_6265,N_4302,N_1696);
nand U6266 (N_6266,N_1878,N_1216);
and U6267 (N_6267,N_3027,N_2195);
or U6268 (N_6268,N_1631,N_2822);
or U6269 (N_6269,N_4449,N_524);
nor U6270 (N_6270,N_2365,N_3028);
nor U6271 (N_6271,N_2952,N_3562);
nand U6272 (N_6272,N_1905,N_1168);
or U6273 (N_6273,N_1285,N_1281);
or U6274 (N_6274,N_4782,N_2420);
and U6275 (N_6275,N_778,N_3703);
nor U6276 (N_6276,N_1540,N_1731);
and U6277 (N_6277,N_3506,N_3962);
and U6278 (N_6278,N_1205,N_4309);
and U6279 (N_6279,N_2620,N_1468);
nor U6280 (N_6280,N_4296,N_2026);
nor U6281 (N_6281,N_4879,N_4929);
nand U6282 (N_6282,N_2691,N_4831);
nand U6283 (N_6283,N_193,N_3057);
nand U6284 (N_6284,N_2669,N_3948);
nand U6285 (N_6285,N_337,N_1656);
and U6286 (N_6286,N_3335,N_2640);
nand U6287 (N_6287,N_2312,N_2501);
nand U6288 (N_6288,N_217,N_2803);
nand U6289 (N_6289,N_1074,N_528);
nand U6290 (N_6290,N_3409,N_3034);
nand U6291 (N_6291,N_2191,N_1473);
xor U6292 (N_6292,N_3096,N_616);
and U6293 (N_6293,N_916,N_716);
nand U6294 (N_6294,N_858,N_4182);
nand U6295 (N_6295,N_712,N_4465);
or U6296 (N_6296,N_2167,N_454);
or U6297 (N_6297,N_2588,N_839);
nand U6298 (N_6298,N_4723,N_707);
or U6299 (N_6299,N_3549,N_2944);
or U6300 (N_6300,N_4130,N_4530);
and U6301 (N_6301,N_1630,N_3053);
nand U6302 (N_6302,N_564,N_2018);
nand U6303 (N_6303,N_4717,N_984);
or U6304 (N_6304,N_1258,N_4165);
nand U6305 (N_6305,N_376,N_3715);
nand U6306 (N_6306,N_1819,N_2434);
nor U6307 (N_6307,N_4805,N_4862);
or U6308 (N_6308,N_1924,N_3169);
nand U6309 (N_6309,N_2884,N_2300);
nand U6310 (N_6310,N_760,N_1013);
or U6311 (N_6311,N_3482,N_3162);
nand U6312 (N_6312,N_4735,N_2176);
nor U6313 (N_6313,N_3544,N_3771);
or U6314 (N_6314,N_628,N_1677);
nand U6315 (N_6315,N_4158,N_3824);
or U6316 (N_6316,N_4306,N_1274);
nor U6317 (N_6317,N_3855,N_150);
or U6318 (N_6318,N_1332,N_3747);
nor U6319 (N_6319,N_1194,N_2237);
nor U6320 (N_6320,N_2703,N_3944);
and U6321 (N_6321,N_4978,N_1066);
nor U6322 (N_6322,N_860,N_3116);
and U6323 (N_6323,N_81,N_4886);
and U6324 (N_6324,N_1067,N_4493);
nor U6325 (N_6325,N_594,N_3623);
nor U6326 (N_6326,N_2356,N_2550);
nand U6327 (N_6327,N_1820,N_4502);
nor U6328 (N_6328,N_2538,N_1099);
and U6329 (N_6329,N_1396,N_4896);
nand U6330 (N_6330,N_237,N_4651);
nand U6331 (N_6331,N_2773,N_844);
and U6332 (N_6332,N_1447,N_2931);
or U6333 (N_6333,N_2308,N_364);
nand U6334 (N_6334,N_4072,N_3461);
nor U6335 (N_6335,N_3975,N_3980);
or U6336 (N_6336,N_695,N_1144);
nand U6337 (N_6337,N_2292,N_1034);
nand U6338 (N_6338,N_791,N_4615);
and U6339 (N_6339,N_1471,N_2347);
and U6340 (N_6340,N_3230,N_4607);
or U6341 (N_6341,N_1232,N_2058);
nand U6342 (N_6342,N_50,N_3465);
and U6343 (N_6343,N_574,N_268);
nand U6344 (N_6344,N_2105,N_3616);
and U6345 (N_6345,N_2104,N_43);
or U6346 (N_6346,N_489,N_4526);
or U6347 (N_6347,N_4789,N_2572);
nand U6348 (N_6348,N_148,N_3760);
nor U6349 (N_6349,N_1588,N_4669);
and U6350 (N_6350,N_3267,N_3086);
nor U6351 (N_6351,N_587,N_4605);
or U6352 (N_6352,N_909,N_759);
nand U6353 (N_6353,N_3120,N_3687);
nand U6354 (N_6354,N_3072,N_2910);
and U6355 (N_6355,N_3561,N_2484);
or U6356 (N_6356,N_798,N_1602);
or U6357 (N_6357,N_2293,N_661);
nand U6358 (N_6358,N_3728,N_99);
xnor U6359 (N_6359,N_343,N_2490);
xnor U6360 (N_6360,N_2190,N_1104);
nand U6361 (N_6361,N_4680,N_4458);
and U6362 (N_6362,N_1617,N_320);
nor U6363 (N_6363,N_125,N_2682);
or U6364 (N_6364,N_1867,N_2047);
nand U6365 (N_6365,N_1087,N_4036);
and U6366 (N_6366,N_1676,N_2818);
or U6367 (N_6367,N_1080,N_1394);
nor U6368 (N_6368,N_1202,N_1183);
nor U6369 (N_6369,N_3339,N_3531);
or U6370 (N_6370,N_3445,N_4697);
and U6371 (N_6371,N_2448,N_4376);
or U6372 (N_6372,N_3849,N_2404);
nor U6373 (N_6373,N_4331,N_3640);
or U6374 (N_6374,N_1241,N_3634);
and U6375 (N_6375,N_833,N_4655);
nand U6376 (N_6376,N_873,N_3266);
or U6377 (N_6377,N_1326,N_2533);
or U6378 (N_6378,N_4054,N_4893);
nor U6379 (N_6379,N_516,N_832);
or U6380 (N_6380,N_232,N_1767);
nand U6381 (N_6381,N_2832,N_2666);
nand U6382 (N_6382,N_2742,N_3583);
nor U6383 (N_6383,N_904,N_882);
nand U6384 (N_6384,N_3131,N_2525);
nor U6385 (N_6385,N_4839,N_741);
or U6386 (N_6386,N_121,N_3723);
xor U6387 (N_6387,N_2390,N_1627);
and U6388 (N_6388,N_3106,N_353);
or U6389 (N_6389,N_997,N_1626);
nand U6390 (N_6390,N_2809,N_3608);
and U6391 (N_6391,N_2531,N_3951);
nand U6392 (N_6392,N_3067,N_2494);
nand U6393 (N_6393,N_244,N_390);
nor U6394 (N_6394,N_2611,N_622);
nand U6395 (N_6395,N_2720,N_4427);
or U6396 (N_6396,N_1988,N_995);
and U6397 (N_6397,N_1652,N_117);
nor U6398 (N_6398,N_4951,N_1292);
or U6399 (N_6399,N_4472,N_4810);
and U6400 (N_6400,N_2187,N_161);
or U6401 (N_6401,N_4945,N_262);
nand U6402 (N_6402,N_4637,N_2418);
nor U6403 (N_6403,N_3662,N_3763);
nor U6404 (N_6404,N_3318,N_6);
nand U6405 (N_6405,N_3554,N_2706);
and U6406 (N_6406,N_4066,N_3943);
nor U6407 (N_6407,N_3977,N_2597);
and U6408 (N_6408,N_3772,N_4187);
nand U6409 (N_6409,N_1174,N_4779);
nand U6410 (N_6410,N_4129,N_1363);
and U6411 (N_6411,N_4326,N_1223);
or U6412 (N_6412,N_2175,N_2497);
or U6413 (N_6413,N_3251,N_511);
or U6414 (N_6414,N_3381,N_617);
or U6415 (N_6415,N_2797,N_7);
or U6416 (N_6416,N_4496,N_1268);
or U6417 (N_6417,N_1277,N_26);
xor U6418 (N_6418,N_1488,N_764);
nand U6419 (N_6419,N_1556,N_3402);
or U6420 (N_6420,N_3961,N_487);
nand U6421 (N_6421,N_2612,N_974);
and U6422 (N_6422,N_1958,N_4190);
nand U6423 (N_6423,N_3784,N_623);
nor U6424 (N_6424,N_317,N_3940);
nor U6425 (N_6425,N_543,N_3881);
nand U6426 (N_6426,N_3367,N_2282);
nor U6427 (N_6427,N_884,N_84);
and U6428 (N_6428,N_3282,N_3380);
nor U6429 (N_6429,N_3353,N_1864);
and U6430 (N_6430,N_2549,N_3042);
and U6431 (N_6431,N_2845,N_4882);
or U6432 (N_6432,N_4877,N_4424);
nor U6433 (N_6433,N_3453,N_1708);
nand U6434 (N_6434,N_2927,N_3436);
xor U6435 (N_6435,N_1971,N_4402);
nand U6436 (N_6436,N_4833,N_4578);
or U6437 (N_6437,N_2695,N_4097);
nor U6438 (N_6438,N_2518,N_1633);
or U6439 (N_6439,N_846,N_2173);
nand U6440 (N_6440,N_1972,N_2689);
nand U6441 (N_6441,N_925,N_2594);
nand U6442 (N_6442,N_963,N_705);
or U6443 (N_6443,N_2763,N_2748);
nor U6444 (N_6444,N_1220,N_4250);
nor U6445 (N_6445,N_2454,N_3263);
nor U6446 (N_6446,N_4046,N_906);
nand U6447 (N_6447,N_1395,N_254);
or U6448 (N_6448,N_1589,N_667);
xnor U6449 (N_6449,N_3876,N_1136);
or U6450 (N_6450,N_87,N_785);
and U6451 (N_6451,N_2547,N_3102);
nor U6452 (N_6452,N_3592,N_4201);
nor U6453 (N_6453,N_3609,N_3896);
nor U6454 (N_6454,N_2082,N_1750);
nor U6455 (N_6455,N_1039,N_4724);
or U6456 (N_6456,N_870,N_3572);
nor U6457 (N_6457,N_1657,N_575);
nand U6458 (N_6458,N_1403,N_1430);
or U6459 (N_6459,N_3889,N_3787);
nor U6460 (N_6460,N_2906,N_45);
xnor U6461 (N_6461,N_2266,N_4009);
nand U6462 (N_6462,N_2489,N_4599);
or U6463 (N_6463,N_3412,N_2363);
nor U6464 (N_6464,N_1450,N_1352);
nand U6465 (N_6465,N_2672,N_333);
or U6466 (N_6466,N_3828,N_608);
or U6467 (N_6467,N_3669,N_565);
or U6468 (N_6468,N_1720,N_4641);
nor U6469 (N_6469,N_1441,N_1899);
nor U6470 (N_6470,N_443,N_4851);
and U6471 (N_6471,N_3094,N_1976);
or U6472 (N_6472,N_4626,N_1789);
nor U6473 (N_6473,N_4904,N_4873);
and U6474 (N_6474,N_4222,N_1309);
nand U6475 (N_6475,N_1091,N_619);
nand U6476 (N_6476,N_3720,N_4770);
nand U6477 (N_6477,N_3701,N_4012);
nor U6478 (N_6478,N_3779,N_3599);
or U6479 (N_6479,N_4121,N_1923);
nor U6480 (N_6480,N_1613,N_2565);
nor U6481 (N_6481,N_3471,N_75);
or U6482 (N_6482,N_4835,N_2320);
nor U6483 (N_6483,N_4603,N_492);
nor U6484 (N_6484,N_1870,N_156);
nor U6485 (N_6485,N_1331,N_2306);
and U6486 (N_6486,N_579,N_3833);
or U6487 (N_6487,N_4645,N_4266);
or U6488 (N_6488,N_4083,N_411);
and U6489 (N_6489,N_2938,N_2893);
and U6490 (N_6490,N_900,N_3869);
nor U6491 (N_6491,N_4283,N_4950);
nand U6492 (N_6492,N_2702,N_2216);
nor U6493 (N_6493,N_4499,N_681);
or U6494 (N_6494,N_1500,N_2765);
nor U6495 (N_6495,N_2709,N_3519);
and U6496 (N_6496,N_3605,N_16);
nand U6497 (N_6497,N_4552,N_3507);
nand U6498 (N_6498,N_690,N_3227);
nor U6499 (N_6499,N_1904,N_4406);
and U6500 (N_6500,N_536,N_406);
nor U6501 (N_6501,N_4428,N_227);
xnor U6502 (N_6502,N_553,N_3219);
or U6503 (N_6503,N_4143,N_2189);
or U6504 (N_6504,N_2488,N_3949);
nand U6505 (N_6505,N_685,N_2056);
or U6506 (N_6506,N_4229,N_2530);
nand U6507 (N_6507,N_4098,N_1736);
or U6508 (N_6508,N_3632,N_4059);
nor U6509 (N_6509,N_3472,N_2305);
and U6510 (N_6510,N_4716,N_3269);
and U6511 (N_6511,N_4736,N_3123);
nor U6512 (N_6512,N_294,N_86);
nand U6513 (N_6513,N_774,N_2591);
and U6514 (N_6514,N_1213,N_665);
and U6515 (N_6515,N_61,N_1538);
nor U6516 (N_6516,N_2379,N_179);
or U6517 (N_6517,N_3525,N_4313);
and U6518 (N_6518,N_3969,N_3677);
nand U6519 (N_6519,N_502,N_952);
nor U6520 (N_6520,N_4454,N_1056);
nand U6521 (N_6521,N_2867,N_3271);
or U6522 (N_6522,N_4073,N_2246);
nor U6523 (N_6523,N_1515,N_3851);
or U6524 (N_6524,N_2959,N_335);
and U6525 (N_6525,N_1621,N_3799);
xor U6526 (N_6526,N_1428,N_3613);
or U6527 (N_6527,N_78,N_4278);
and U6528 (N_6528,N_1679,N_1950);
or U6529 (N_6529,N_250,N_4956);
and U6530 (N_6530,N_731,N_266);
nor U6531 (N_6531,N_2839,N_83);
and U6532 (N_6532,N_2127,N_4760);
or U6533 (N_6533,N_1919,N_3793);
or U6534 (N_6534,N_1700,N_2137);
or U6535 (N_6535,N_2253,N_2681);
or U6536 (N_6536,N_2183,N_4310);
nor U6537 (N_6537,N_4612,N_4859);
nor U6538 (N_6538,N_555,N_2736);
and U6539 (N_6539,N_3891,N_1783);
and U6540 (N_6540,N_2366,N_3134);
and U6541 (N_6541,N_2192,N_1687);
nor U6542 (N_6542,N_4549,N_2679);
and U6543 (N_6543,N_1832,N_1792);
or U6544 (N_6544,N_1419,N_2684);
nor U6545 (N_6545,N_2091,N_2027);
or U6546 (N_6546,N_2000,N_2019);
or U6547 (N_6547,N_752,N_2362);
nor U6548 (N_6548,N_735,N_3826);
or U6549 (N_6549,N_1752,N_62);
or U6550 (N_6550,N_3684,N_3250);
nor U6551 (N_6551,N_3741,N_4478);
or U6552 (N_6552,N_225,N_1131);
nor U6553 (N_6553,N_4708,N_4422);
and U6554 (N_6554,N_4852,N_4589);
nand U6555 (N_6555,N_3593,N_4565);
and U6556 (N_6556,N_3065,N_216);
nand U6557 (N_6557,N_2710,N_3838);
nor U6558 (N_6558,N_1666,N_341);
nand U6559 (N_6559,N_1251,N_3491);
nand U6560 (N_6560,N_3614,N_4512);
and U6561 (N_6561,N_1427,N_2277);
nor U6562 (N_6562,N_3244,N_940);
or U6563 (N_6563,N_1040,N_2960);
or U6564 (N_6564,N_378,N_4649);
nor U6565 (N_6565,N_4604,N_4660);
and U6566 (N_6566,N_144,N_2853);
nand U6567 (N_6567,N_4237,N_441);
and U6568 (N_6568,N_4966,N_1915);
or U6569 (N_6569,N_2345,N_14);
and U6570 (N_6570,N_2389,N_3906);
nand U6571 (N_6571,N_2371,N_4899);
nor U6572 (N_6572,N_4701,N_4979);
nor U6573 (N_6573,N_3023,N_3212);
nand U6574 (N_6574,N_1887,N_2847);
nand U6575 (N_6575,N_3351,N_4939);
nor U6576 (N_6576,N_2878,N_153);
or U6577 (N_6577,N_2579,N_2922);
nor U6578 (N_6578,N_4140,N_1199);
and U6579 (N_6579,N_743,N_260);
nand U6580 (N_6580,N_1476,N_4692);
nor U6581 (N_6581,N_800,N_3423);
or U6582 (N_6582,N_2913,N_1505);
nand U6583 (N_6583,N_1109,N_4329);
or U6584 (N_6584,N_3119,N_4219);
nand U6585 (N_6585,N_70,N_2554);
or U6586 (N_6586,N_1334,N_2121);
nand U6587 (N_6587,N_1560,N_3021);
or U6588 (N_6588,N_3400,N_2248);
or U6589 (N_6589,N_3439,N_332);
nor U6590 (N_6590,N_3816,N_2102);
nor U6591 (N_6591,N_3069,N_921);
xnor U6592 (N_6592,N_793,N_4855);
nor U6593 (N_6593,N_4944,N_1735);
or U6594 (N_6594,N_2421,N_2067);
and U6595 (N_6595,N_3459,N_4763);
and U6596 (N_6596,N_2008,N_3097);
xor U6597 (N_6597,N_4585,N_1315);
or U6598 (N_6598,N_956,N_2435);
nor U6599 (N_6599,N_2891,N_3624);
or U6600 (N_6600,N_120,N_1927);
nand U6601 (N_6601,N_434,N_1583);
nand U6602 (N_6602,N_1472,N_4045);
or U6603 (N_6603,N_405,N_2970);
nand U6604 (N_6604,N_4715,N_955);
nor U6605 (N_6605,N_2077,N_2004);
or U6606 (N_6606,N_1393,N_2889);
nor U6607 (N_6607,N_1340,N_1398);
and U6608 (N_6608,N_4546,N_3071);
nand U6609 (N_6609,N_4276,N_1042);
or U6610 (N_6610,N_2271,N_3657);
or U6611 (N_6611,N_538,N_4812);
nor U6612 (N_6612,N_3496,N_784);
or U6613 (N_6613,N_344,N_155);
and U6614 (N_6614,N_2649,N_4513);
nor U6615 (N_6615,N_4005,N_3540);
nor U6616 (N_6616,N_1378,N_1188);
nor U6617 (N_6617,N_810,N_4584);
or U6618 (N_6618,N_1701,N_4775);
or U6619 (N_6619,N_2548,N_2982);
and U6620 (N_6620,N_1482,N_3386);
and U6621 (N_6621,N_816,N_3761);
nor U6622 (N_6622,N_3965,N_4051);
nand U6623 (N_6623,N_1879,N_2503);
and U6624 (N_6624,N_2442,N_1149);
nor U6625 (N_6625,N_2635,N_2337);
and U6626 (N_6626,N_1114,N_4489);
and U6627 (N_6627,N_3217,N_1283);
xnor U6628 (N_6628,N_4210,N_3013);
nor U6629 (N_6629,N_3246,N_3602);
nand U6630 (N_6630,N_2223,N_1848);
or U6631 (N_6631,N_28,N_3660);
nor U6632 (N_6632,N_1197,N_644);
or U6633 (N_6633,N_1434,N_922);
nor U6634 (N_6634,N_1410,N_4514);
or U6635 (N_6635,N_3642,N_12);
nor U6636 (N_6636,N_633,N_3719);
or U6637 (N_6637,N_2042,N_4972);
nand U6638 (N_6638,N_1805,N_603);
or U6639 (N_6639,N_1079,N_1009);
and U6640 (N_6640,N_3551,N_3036);
nor U6641 (N_6641,N_3279,N_3490);
nor U6642 (N_6642,N_4933,N_2701);
nor U6643 (N_6643,N_2633,N_2711);
nand U6644 (N_6644,N_4674,N_168);
and U6645 (N_6645,N_4328,N_4841);
or U6646 (N_6646,N_4915,N_2506);
nand U6647 (N_6647,N_4021,N_2281);
and U6648 (N_6648,N_1726,N_1580);
nand U6649 (N_6649,N_4290,N_273);
and U6650 (N_6650,N_2168,N_648);
and U6651 (N_6651,N_1084,N_4602);
nand U6652 (N_6652,N_3079,N_4544);
nor U6653 (N_6653,N_1146,N_1926);
or U6654 (N_6654,N_4377,N_2031);
nand U6655 (N_6655,N_1298,N_42);
nand U6656 (N_6656,N_938,N_4924);
or U6657 (N_6657,N_4439,N_2014);
and U6658 (N_6658,N_4407,N_2716);
and U6659 (N_6659,N_4518,N_4799);
or U6660 (N_6660,N_4133,N_138);
nor U6661 (N_6661,N_2038,N_2259);
or U6662 (N_6662,N_2987,N_4063);
nor U6663 (N_6663,N_4230,N_1506);
nand U6664 (N_6664,N_2126,N_4807);
or U6665 (N_6665,N_3580,N_3108);
and U6666 (N_6666,N_4014,N_473);
or U6667 (N_6667,N_389,N_2621);
and U6668 (N_6668,N_455,N_2251);
and U6669 (N_6669,N_4227,N_1579);
or U6670 (N_6670,N_2011,N_2353);
nand U6671 (N_6671,N_2261,N_3041);
and U6672 (N_6672,N_1609,N_3008);
nand U6673 (N_6673,N_4410,N_1243);
xor U6674 (N_6674,N_3671,N_4343);
or U6675 (N_6675,N_2741,N_2220);
nand U6676 (N_6676,N_2152,N_4648);
nor U6677 (N_6677,N_1308,N_930);
or U6678 (N_6678,N_3857,N_2393);
or U6679 (N_6679,N_4681,N_1239);
nor U6680 (N_6680,N_3376,N_2718);
and U6681 (N_6681,N_2084,N_585);
nand U6682 (N_6682,N_660,N_3248);
and U6683 (N_6683,N_3966,N_3512);
or U6684 (N_6684,N_22,N_2409);
or U6685 (N_6685,N_4344,N_4957);
and U6686 (N_6686,N_1357,N_2502);
and U6687 (N_6687,N_711,N_3375);
and U6688 (N_6688,N_3464,N_3880);
nand U6689 (N_6689,N_4842,N_1339);
nand U6690 (N_6690,N_3165,N_2469);
nor U6691 (N_6691,N_4787,N_56);
nor U6692 (N_6692,N_692,N_32);
nor U6693 (N_6693,N_3920,N_2657);
or U6694 (N_6694,N_1704,N_4529);
nand U6695 (N_6695,N_407,N_3360);
or U6696 (N_6696,N_1833,N_4573);
and U6697 (N_6697,N_500,N_2973);
and U6698 (N_6698,N_3477,N_1737);
and U6699 (N_6699,N_4744,N_1198);
nand U6700 (N_6700,N_1354,N_1728);
and U6701 (N_6701,N_4557,N_1692);
nor U6702 (N_6702,N_942,N_825);
and U6703 (N_6703,N_2815,N_654);
or U6704 (N_6704,N_2638,N_2079);
or U6705 (N_6705,N_3125,N_2250);
nand U6706 (N_6706,N_1117,N_102);
nand U6707 (N_6707,N_1184,N_2855);
or U6708 (N_6708,N_645,N_704);
or U6709 (N_6709,N_1632,N_187);
nand U6710 (N_6710,N_4103,N_1587);
nor U6711 (N_6711,N_982,N_1822);
and U6712 (N_6712,N_2673,N_1521);
or U6713 (N_6713,N_4216,N_95);
nand U6714 (N_6714,N_3107,N_4560);
nor U6715 (N_6715,N_2683,N_4498);
nor U6716 (N_6716,N_3818,N_2088);
or U6717 (N_6717,N_596,N_756);
and U6718 (N_6718,N_2529,N_281);
nor U6719 (N_6719,N_2433,N_4166);
or U6720 (N_6720,N_4675,N_2785);
nor U6721 (N_6721,N_1006,N_805);
or U6722 (N_6722,N_959,N_3607);
and U6723 (N_6723,N_3727,N_2897);
and U6724 (N_6724,N_2081,N_4900);
nor U6725 (N_6725,N_113,N_2);
nand U6726 (N_6726,N_673,N_4918);
nor U6727 (N_6727,N_4832,N_1593);
and U6728 (N_6728,N_3606,N_1178);
and U6729 (N_6729,N_382,N_954);
nand U6730 (N_6730,N_3393,N_4976);
nand U6731 (N_6731,N_4720,N_261);
nand U6732 (N_6732,N_3231,N_3050);
nand U6733 (N_6733,N_381,N_1889);
nor U6734 (N_6734,N_558,N_2054);
or U6735 (N_6735,N_2557,N_1641);
and U6736 (N_6736,N_39,N_4820);
or U6737 (N_6737,N_1746,N_4200);
nand U6738 (N_6738,N_2164,N_3054);
nor U6739 (N_6739,N_1209,N_3754);
nand U6740 (N_6740,N_1423,N_517);
nand U6741 (N_6741,N_2511,N_3347);
nand U6742 (N_6742,N_137,N_108);
nand U6743 (N_6743,N_3196,N_1289);
nand U6744 (N_6744,N_3389,N_211);
and U6745 (N_6745,N_288,N_284);
or U6746 (N_6746,N_4906,N_1511);
nand U6747 (N_6747,N_1418,N_3209);
and U6748 (N_6748,N_3783,N_3970);
or U6749 (N_6749,N_867,N_3016);
and U6750 (N_6750,N_1415,N_3148);
and U6751 (N_6751,N_2985,N_969);
nor U6752 (N_6752,N_54,N_4367);
nand U6753 (N_6753,N_4503,N_1846);
or U6754 (N_6754,N_1088,N_3714);
nand U6755 (N_6755,N_90,N_2290);
nand U6756 (N_6756,N_2652,N_352);
nor U6757 (N_6757,N_457,N_400);
or U6758 (N_6758,N_3448,N_980);
and U6759 (N_6759,N_3568,N_4624);
nand U6760 (N_6760,N_1907,N_4338);
and U6761 (N_6761,N_164,N_4341);
or U6762 (N_6762,N_3659,N_290);
nor U6763 (N_6763,N_989,N_856);
nor U6764 (N_6764,N_3934,N_1898);
and U6765 (N_6765,N_2243,N_1946);
nor U6766 (N_6766,N_3005,N_3986);
and U6767 (N_6767,N_655,N_1404);
or U6768 (N_6768,N_4445,N_886);
nand U6769 (N_6769,N_2789,N_2515);
nand U6770 (N_6770,N_1713,N_2894);
nor U6771 (N_6771,N_1561,N_1288);
and U6772 (N_6772,N_1862,N_1975);
and U6773 (N_6773,N_4157,N_4149);
nand U6774 (N_6774,N_796,N_3939);
nor U6775 (N_6775,N_4738,N_4762);
nor U6776 (N_6776,N_4116,N_182);
nand U6777 (N_6777,N_1445,N_571);
or U6778 (N_6778,N_3305,N_3237);
nand U6779 (N_6779,N_1324,N_4181);
nor U6780 (N_6780,N_3298,N_2962);
and U6781 (N_6781,N_4349,N_1245);
or U6782 (N_6782,N_945,N_3883);
nand U6783 (N_6783,N_2302,N_3517);
nor U6784 (N_6784,N_391,N_1782);
nand U6785 (N_6785,N_452,N_2831);
nor U6786 (N_6786,N_610,N_4476);
xor U6787 (N_6787,N_4425,N_1106);
nor U6788 (N_6788,N_2966,N_3286);
or U6789 (N_6789,N_37,N_1647);
nand U6790 (N_6790,N_827,N_3566);
nand U6791 (N_6791,N_3095,N_2177);
nand U6792 (N_6792,N_4245,N_3132);
or U6793 (N_6793,N_334,N_4751);
or U6794 (N_6794,N_2739,N_985);
nand U6795 (N_6795,N_2881,N_3612);
nand U6796 (N_6796,N_2645,N_2979);
or U6797 (N_6797,N_4085,N_2318);
or U6798 (N_6798,N_642,N_2450);
nor U6799 (N_6799,N_3546,N_2475);
or U6800 (N_6800,N_4927,N_3017);
nand U6801 (N_6801,N_604,N_4654);
and U6802 (N_6802,N_2883,N_4652);
or U6803 (N_6803,N_1381,N_2743);
nor U6804 (N_6804,N_3942,N_1876);
and U6805 (N_6805,N_4890,N_2194);
or U6806 (N_6806,N_2592,N_74);
or U6807 (N_6807,N_4301,N_1413);
and U6808 (N_6808,N_881,N_3622);
or U6809 (N_6809,N_4404,N_259);
nand U6810 (N_6810,N_3812,N_2955);
and U6811 (N_6811,N_4254,N_3163);
nor U6812 (N_6812,N_4853,N_2574);
nor U6813 (N_6813,N_586,N_59);
and U6814 (N_6814,N_1303,N_4000);
and U6815 (N_6815,N_1115,N_3081);
and U6816 (N_6816,N_2064,N_3356);
nand U6817 (N_6817,N_3510,N_3835);
or U6818 (N_6818,N_4370,N_2852);
nor U6819 (N_6819,N_3433,N_1559);
nand U6820 (N_6820,N_2808,N_4726);
nor U6821 (N_6821,N_2072,N_683);
and U6822 (N_6822,N_4846,N_4039);
nand U6823 (N_6823,N_3287,N_1479);
nand U6824 (N_6824,N_570,N_3557);
nand U6825 (N_6825,N_2713,N_4113);
nand U6826 (N_6826,N_4104,N_788);
and U6827 (N_6827,N_4608,N_4115);
or U6828 (N_6828,N_3689,N_3798);
or U6829 (N_6829,N_3344,N_1892);
nor U6830 (N_6830,N_1157,N_3831);
xnor U6831 (N_6831,N_1510,N_2432);
and U6832 (N_6832,N_561,N_2202);
nand U6833 (N_6833,N_792,N_2208);
nand U6834 (N_6834,N_4834,N_3707);
and U6835 (N_6835,N_4195,N_3429);
and U6836 (N_6836,N_2471,N_2464);
or U6837 (N_6837,N_186,N_1316);
and U6838 (N_6838,N_4469,N_3968);
and U6839 (N_6839,N_2802,N_2334);
and U6840 (N_6840,N_4360,N_3726);
nand U6841 (N_6841,N_797,N_2957);
nand U6842 (N_6842,N_2407,N_3216);
or U6843 (N_6843,N_4809,N_2452);
or U6844 (N_6844,N_282,N_826);
nor U6845 (N_6845,N_4570,N_2068);
and U6846 (N_6846,N_3908,N_559);
or U6847 (N_6847,N_3997,N_410);
nor U6848 (N_6848,N_4630,N_638);
nor U6849 (N_6849,N_1480,N_2140);
and U6850 (N_6850,N_2394,N_546);
or U6851 (N_6851,N_2575,N_1969);
or U6852 (N_6852,N_4547,N_4308);
nor U6853 (N_6853,N_4622,N_3166);
nor U6854 (N_6854,N_4908,N_3160);
and U6855 (N_6855,N_4935,N_1397);
or U6856 (N_6856,N_2562,N_918);
and U6857 (N_6857,N_3791,N_4117);
nand U6858 (N_6858,N_1236,N_779);
nand U6859 (N_6859,N_3960,N_958);
nor U6860 (N_6860,N_3104,N_3365);
xnor U6861 (N_6861,N_2752,N_2552);
nand U6862 (N_6862,N_4409,N_48);
and U6863 (N_6863,N_413,N_4958);
nor U6864 (N_6864,N_3903,N_2427);
xnor U6865 (N_6865,N_552,N_1935);
or U6866 (N_6866,N_799,N_2199);
and U6867 (N_6867,N_671,N_127);
and U6868 (N_6868,N_912,N_1682);
or U6869 (N_6869,N_2814,N_310);
or U6870 (N_6870,N_2536,N_2969);
nor U6871 (N_6871,N_1003,N_4248);
or U6872 (N_6872,N_181,N_3795);
nand U6873 (N_6873,N_4355,N_3809);
nor U6874 (N_6874,N_2896,N_451);
and U6875 (N_6875,N_4423,N_4261);
and U6876 (N_6876,N_1886,N_1803);
or U6877 (N_6877,N_3440,N_2255);
nand U6878 (N_6878,N_3100,N_728);
and U6879 (N_6879,N_3733,N_1388);
nand U6880 (N_6880,N_841,N_818);
or U6881 (N_6881,N_2165,N_747);
and U6882 (N_6882,N_4126,N_4267);
or U6883 (N_6883,N_3007,N_1874);
nor U6884 (N_6884,N_599,N_607);
nand U6885 (N_6885,N_2229,N_4959);
nor U6886 (N_6886,N_1238,N_1934);
or U6887 (N_6887,N_2286,N_4184);
and U6888 (N_6888,N_2690,N_4580);
and U6889 (N_6889,N_1314,N_1990);
or U6890 (N_6890,N_3181,N_230);
nand U6891 (N_6891,N_3037,N_354);
or U6892 (N_6892,N_4984,N_2035);
and U6893 (N_6893,N_1793,N_4876);
nor U6894 (N_6894,N_3068,N_342);
and U6895 (N_6895,N_1836,N_3646);
and U6896 (N_6896,N_771,N_1841);
or U6897 (N_6897,N_3526,N_2887);
nand U6898 (N_6898,N_4657,N_2986);
nand U6899 (N_6899,N_2505,N_4002);
nor U6900 (N_6900,N_2495,N_4318);
nand U6901 (N_6901,N_2903,N_3688);
and U6902 (N_6902,N_4109,N_3686);
or U6903 (N_6903,N_3059,N_2732);
and U6904 (N_6904,N_1529,N_3438);
nor U6905 (N_6905,N_593,N_128);
or U6906 (N_6906,N_387,N_4258);
nand U6907 (N_6907,N_4356,N_2868);
and U6908 (N_6908,N_3369,N_639);
and U6909 (N_6909,N_2240,N_3283);
and U6910 (N_6910,N_1341,N_303);
and U6911 (N_6911,N_2728,N_2745);
nand U6912 (N_6912,N_1718,N_4581);
and U6913 (N_6913,N_3643,N_1459);
nor U6914 (N_6914,N_3533,N_3147);
nor U6915 (N_6915,N_1821,N_146);
nand U6916 (N_6916,N_4434,N_3395);
nor U6917 (N_6917,N_1145,N_2776);
nor U6918 (N_6918,N_768,N_983);
and U6919 (N_6919,N_2384,N_2954);
or U6920 (N_6920,N_4068,N_1530);
nor U6921 (N_6921,N_3310,N_58);
or U6922 (N_6922,N_2083,N_1917);
and U6923 (N_6923,N_1260,N_3637);
nand U6924 (N_6924,N_2459,N_2941);
nand U6925 (N_6925,N_3245,N_1193);
and U6926 (N_6926,N_2453,N_1463);
nand U6927 (N_6927,N_2553,N_2213);
xor U6928 (N_6928,N_4967,N_1858);
nand U6929 (N_6929,N_1001,N_3675);
nor U6930 (N_6930,N_2540,N_1964);
and U6931 (N_6931,N_3332,N_3022);
xnor U6932 (N_6932,N_4745,N_4753);
and U6933 (N_6933,N_612,N_3215);
or U6934 (N_6934,N_2089,N_1017);
or U6935 (N_6935,N_2619,N_557);
and U6936 (N_6936,N_1070,N_2508);
or U6937 (N_6937,N_3268,N_1660);
nand U6938 (N_6938,N_1977,N_1151);
nand U6939 (N_6939,N_3317,N_1152);
nand U6940 (N_6940,N_3751,N_3628);
nor U6941 (N_6941,N_3915,N_3746);
and U6942 (N_6942,N_2321,N_501);
or U6943 (N_6943,N_3430,N_1868);
and U6944 (N_6944,N_1474,N_4481);
nand U6945 (N_6945,N_1344,N_4545);
nand U6946 (N_6946,N_1861,N_3736);
and U6947 (N_6947,N_966,N_3135);
and U6948 (N_6948,N_4895,N_2196);
nor U6949 (N_6949,N_3839,N_3515);
nor U6950 (N_6950,N_1532,N_1207);
nor U6951 (N_6951,N_4342,N_1507);
and U6952 (N_6952,N_1998,N_4691);
or U6953 (N_6953,N_3695,N_4506);
nor U6954 (N_6954,N_2198,N_1875);
and U6955 (N_6955,N_2377,N_1242);
nand U6956 (N_6956,N_2078,N_2103);
nand U6957 (N_6957,N_3537,N_3151);
or U6958 (N_6958,N_848,N_3327);
nand U6959 (N_6959,N_1961,N_4414);
nor U6960 (N_6960,N_3179,N_986);
nor U6961 (N_6961,N_2698,N_1920);
and U6962 (N_6962,N_3372,N_2256);
nor U6963 (N_6963,N_3048,N_2696);
and U6964 (N_6964,N_2731,N_1382);
and U6965 (N_6965,N_3030,N_2580);
and U6966 (N_6966,N_1389,N_136);
and U6967 (N_6967,N_4416,N_3112);
or U6968 (N_6968,N_2543,N_573);
nor U6969 (N_6969,N_4383,N_2460);
and U6970 (N_6970,N_4561,N_2556);
and U6971 (N_6971,N_2779,N_2080);
or U6972 (N_6972,N_4562,N_1453);
or U6973 (N_6973,N_1163,N_4803);
nand U6974 (N_6974,N_4684,N_869);
nand U6975 (N_6975,N_3401,N_1620);
or U6976 (N_6976,N_1815,N_2029);
nand U6977 (N_6977,N_1702,N_2438);
nand U6978 (N_6978,N_4961,N_897);
nand U6979 (N_6979,N_4568,N_2174);
or U6980 (N_6980,N_4677,N_210);
nand U6981 (N_6981,N_2528,N_1124);
and U6982 (N_6982,N_491,N_3766);
nor U6983 (N_6983,N_3130,N_2841);
nor U6984 (N_6984,N_3825,N_3909);
or U6985 (N_6985,N_4713,N_1210);
or U6986 (N_6986,N_2144,N_2142);
nand U6987 (N_6987,N_1348,N_4647);
and U6988 (N_6988,N_1508,N_152);
or U6989 (N_6989,N_1606,N_631);
nor U6990 (N_6990,N_4317,N_775);
nor U6991 (N_6991,N_4325,N_1684);
and U6992 (N_6992,N_1570,N_471);
nand U6993 (N_6993,N_3257,N_3742);
nand U6994 (N_6994,N_129,N_2734);
and U6995 (N_6995,N_618,N_1385);
nand U6996 (N_6996,N_4100,N_3817);
and U6997 (N_6997,N_2983,N_1978);
or U6998 (N_6998,N_4575,N_576);
or U6999 (N_6999,N_4985,N_4670);
or U7000 (N_7000,N_1358,N_3802);
or U7001 (N_7001,N_2157,N_1097);
nor U7002 (N_7002,N_2570,N_2166);
or U7003 (N_7003,N_1931,N_2918);
or U7004 (N_7004,N_572,N_3328);
or U7005 (N_7005,N_30,N_4515);
nand U7006 (N_7006,N_433,N_2063);
and U7007 (N_7007,N_2159,N_2975);
nand U7008 (N_7008,N_3039,N_605);
nor U7009 (N_7009,N_3973,N_2516);
nor U7010 (N_7010,N_1763,N_4429);
nand U7011 (N_7011,N_183,N_4905);
nand U7012 (N_7012,N_1562,N_2402);
or U7013 (N_7013,N_1654,N_4791);
nor U7014 (N_7014,N_2322,N_2933);
or U7015 (N_7015,N_3252,N_403);
and U7016 (N_7016,N_766,N_4928);
or U7017 (N_7017,N_1600,N_2151);
nand U7018 (N_7018,N_790,N_3058);
nand U7019 (N_7019,N_1721,N_948);
and U7020 (N_7020,N_1739,N_264);
and U7021 (N_7021,N_4964,N_1785);
nand U7022 (N_7022,N_4324,N_2608);
or U7023 (N_7023,N_4659,N_2613);
or U7024 (N_7024,N_2129,N_4623);
and U7025 (N_7025,N_583,N_1653);
nor U7026 (N_7026,N_1501,N_4152);
nor U7027 (N_7027,N_420,N_2882);
and U7028 (N_7028,N_428,N_804);
or U7029 (N_7029,N_687,N_929);
nor U7030 (N_7030,N_1246,N_3449);
and U7031 (N_7031,N_439,N_4285);
nand U7032 (N_7032,N_2777,N_1928);
nand U7033 (N_7033,N_2087,N_3451);
or U7034 (N_7034,N_3006,N_3603);
and U7035 (N_7035,N_2059,N_265);
nor U7036 (N_7036,N_510,N_4069);
or U7037 (N_7037,N_1098,N_4916);
nor U7038 (N_7038,N_4801,N_4300);
and U7039 (N_7039,N_1287,N_1573);
or U7040 (N_7040,N_2676,N_2639);
and U7041 (N_7041,N_745,N_2233);
and U7042 (N_7042,N_3541,N_1603);
nor U7043 (N_7043,N_4800,N_4756);
nor U7044 (N_7044,N_3374,N_3038);
or U7045 (N_7045,N_1531,N_122);
nand U7046 (N_7046,N_2768,N_325);
or U7047 (N_7047,N_4405,N_458);
nor U7048 (N_7048,N_503,N_3018);
nor U7049 (N_7049,N_1575,N_202);
and U7050 (N_7050,N_1809,N_4244);
and U7051 (N_7051,N_470,N_2595);
nor U7052 (N_7052,N_1823,N_4362);
nor U7053 (N_7053,N_4074,N_1346);
nand U7054 (N_7054,N_1753,N_1320);
nand U7055 (N_7055,N_2399,N_88);
nand U7056 (N_7056,N_1854,N_866);
nand U7057 (N_7057,N_1738,N_2398);
and U7058 (N_7058,N_4110,N_993);
and U7059 (N_7059,N_3457,N_4572);
xor U7060 (N_7060,N_567,N_2415);
or U7061 (N_7061,N_3015,N_1936);
nand U7062 (N_7062,N_2401,N_3359);
nor U7063 (N_7063,N_3410,N_475);
nor U7064 (N_7064,N_4883,N_2413);
nor U7065 (N_7065,N_2848,N_4015);
nor U7066 (N_7066,N_1873,N_4925);
and U7067 (N_7067,N_2227,N_722);
nor U7068 (N_7068,N_1877,N_620);
and U7069 (N_7069,N_2916,N_1584);
and U7070 (N_7070,N_3083,N_2446);
nand U7071 (N_7071,N_2723,N_4558);
nand U7072 (N_7072,N_753,N_4794);
nor U7073 (N_7073,N_1645,N_4228);
or U7074 (N_7074,N_4092,N_481);
or U7075 (N_7075,N_4185,N_807);
and U7076 (N_7076,N_1313,N_4475);
nand U7077 (N_7077,N_3874,N_4205);
and U7078 (N_7078,N_4442,N_1658);
or U7079 (N_7079,N_4035,N_482);
nand U7080 (N_7080,N_2603,N_4440);
nor U7081 (N_7081,N_1817,N_3481);
nand U7082 (N_7082,N_384,N_1402);
and U7083 (N_7083,N_2509,N_2414);
nand U7084 (N_7084,N_4432,N_435);
and U7085 (N_7085,N_2917,N_309);
nor U7086 (N_7086,N_4412,N_4826);
nor U7087 (N_7087,N_300,N_3462);
and U7088 (N_7088,N_3542,N_2332);
and U7089 (N_7089,N_936,N_4384);
and U7090 (N_7090,N_3290,N_3740);
nand U7091 (N_7091,N_1008,N_1943);
nand U7092 (N_7092,N_3133,N_3792);
and U7093 (N_7093,N_3469,N_3049);
nand U7094 (N_7094,N_4739,N_2568);
nor U7095 (N_7095,N_1401,N_1635);
nand U7096 (N_7096,N_3455,N_1177);
and U7097 (N_7097,N_1629,N_4433);
and U7098 (N_7098,N_1064,N_1092);
and U7099 (N_7099,N_2826,N_2118);
and U7100 (N_7100,N_3155,N_630);
and U7101 (N_7101,N_4579,N_4056);
nor U7102 (N_7102,N_970,N_4111);
or U7103 (N_7103,N_9,N_1035);
and U7104 (N_7104,N_2900,N_1790);
nand U7105 (N_7105,N_2205,N_3447);
nor U7106 (N_7106,N_4490,N_283);
nor U7107 (N_7107,N_3954,N_1902);
or U7108 (N_7108,N_3963,N_2125);
nor U7109 (N_7109,N_447,N_2836);
or U7110 (N_7110,N_4024,N_3239);
nand U7111 (N_7111,N_4233,N_2899);
or U7112 (N_7112,N_224,N_4816);
and U7113 (N_7113,N_2204,N_730);
and U7114 (N_7114,N_4777,N_2980);
and U7115 (N_7115,N_812,N_2001);
and U7116 (N_7116,N_4027,N_3596);
or U7117 (N_7117,N_1204,N_338);
or U7118 (N_7118,N_3829,N_4217);
nand U7119 (N_7119,N_2447,N_662);
or U7120 (N_7120,N_1786,N_3852);
and U7121 (N_7121,N_2485,N_2942);
nor U7122 (N_7122,N_1550,N_2733);
and U7123 (N_7123,N_2693,N_811);
or U7124 (N_7124,N_3859,N_3879);
or U7125 (N_7125,N_2751,N_1525);
and U7126 (N_7126,N_1999,N_2704);
nand U7127 (N_7127,N_672,N_358);
nor U7128 (N_7128,N_2820,N_855);
and U7129 (N_7129,N_3434,N_4710);
nand U7130 (N_7130,N_1082,N_2618);
or U7131 (N_7131,N_2002,N_2354);
nor U7132 (N_7132,N_2287,N_4970);
and U7133 (N_7133,N_3538,N_3805);
or U7134 (N_7134,N_3823,N_2301);
nor U7135 (N_7135,N_241,N_3800);
and U7136 (N_7136,N_3074,N_4980);
or U7137 (N_7137,N_4279,N_1801);
nand U7138 (N_7138,N_2605,N_3672);
nor U7139 (N_7139,N_2317,N_1544);
or U7140 (N_7140,N_2600,N_139);
or U7141 (N_7141,N_1023,N_589);
and U7142 (N_7142,N_3066,N_578);
and U7143 (N_7143,N_3466,N_527);
nor U7144 (N_7144,N_2688,N_3156);
and U7145 (N_7145,N_2658,N_2425);
nor U7146 (N_7146,N_3600,N_3735);
nand U7147 (N_7147,N_1465,N_750);
nand U7148 (N_7148,N_2034,N_3254);
nand U7149 (N_7149,N_324,N_4443);
and U7150 (N_7150,N_496,N_651);
nor U7151 (N_7151,N_2721,N_2616);
nand U7152 (N_7152,N_1495,N_2491);
nor U7153 (N_7153,N_506,N_3349);
and U7154 (N_7154,N_3025,N_4650);
nor U7155 (N_7155,N_1048,N_1475);
or U7156 (N_7156,N_2148,N_782);
xor U7157 (N_7157,N_1061,N_4272);
nand U7158 (N_7158,N_2599,N_4837);
nor U7159 (N_7159,N_4461,N_1552);
nand U7160 (N_7160,N_401,N_4138);
and U7161 (N_7161,N_1831,N_2313);
or U7162 (N_7162,N_777,N_3004);
nand U7163 (N_7163,N_3850,N_1446);
nor U7164 (N_7164,N_2481,N_3403);
nand U7165 (N_7165,N_1176,N_3398);
nand U7166 (N_7166,N_1616,N_932);
and U7167 (N_7167,N_3842,N_3383);
and U7168 (N_7168,N_2623,N_2141);
nor U7169 (N_7169,N_2584,N_2961);
nand U7170 (N_7170,N_1644,N_3847);
nand U7171 (N_7171,N_4231,N_3589);
or U7172 (N_7172,N_3990,N_1764);
xnor U7173 (N_7173,N_3333,N_3309);
nand U7174 (N_7174,N_1581,N_3088);
or U7175 (N_7175,N_652,N_3748);
nand U7176 (N_7176,N_2386,N_3422);
nand U7177 (N_7177,N_1444,N_4844);
nand U7178 (N_7178,N_2914,N_4320);
nor U7179 (N_7179,N_2965,N_3993);
nand U7180 (N_7180,N_2226,N_2817);
nor U7181 (N_7181,N_4277,N_124);
nor U7182 (N_7182,N_3056,N_2368);
and U7183 (N_7183,N_776,N_2610);
nand U7184 (N_7184,N_2816,N_4202);
and U7185 (N_7185,N_103,N_2885);
nor U7186 (N_7186,N_754,N_787);
nor U7187 (N_7187,N_717,N_1060);
nor U7188 (N_7188,N_3408,N_4969);
or U7189 (N_7189,N_2225,N_3644);
nand U7190 (N_7190,N_3658,N_2342);
and U7191 (N_7191,N_2021,N_1830);
and U7192 (N_7192,N_3425,N_3930);
nor U7193 (N_7193,N_2017,N_2375);
nor U7194 (N_7194,N_3520,N_2436);
and U7195 (N_7195,N_91,N_2441);
nand U7196 (N_7196,N_2534,N_2846);
and U7197 (N_7197,N_2422,N_1072);
or U7198 (N_7198,N_430,N_4345);
and U7199 (N_7199,N_4323,N_4507);
nor U7200 (N_7200,N_1843,N_1208);
nand U7201 (N_7201,N_1734,N_4145);
xor U7202 (N_7202,N_2655,N_851);
and U7203 (N_7203,N_1690,N_1651);
nor U7204 (N_7204,N_3296,N_3221);
or U7205 (N_7205,N_2214,N_4907);
or U7206 (N_7206,N_2740,N_2252);
nand U7207 (N_7207,N_2866,N_4155);
nor U7208 (N_7208,N_3070,N_3012);
nand U7209 (N_7209,N_4391,N_4055);
nor U7210 (N_7210,N_1744,N_1834);
nor U7211 (N_7211,N_1555,N_1078);
nand U7212 (N_7212,N_2268,N_2953);
and U7213 (N_7213,N_2648,N_1155);
and U7214 (N_7214,N_3164,N_4273);
or U7215 (N_7215,N_4160,N_1129);
nor U7216 (N_7216,N_3063,N_3738);
nor U7217 (N_7217,N_154,N_709);
nor U7218 (N_7218,N_874,N_2051);
or U7219 (N_7219,N_2085,N_4534);
nor U7220 (N_7220,N_4159,N_3548);
and U7221 (N_7221,N_4379,N_2329);
and U7222 (N_7222,N_4488,N_1122);
nor U7223 (N_7223,N_4550,N_1263);
nor U7224 (N_7224,N_3158,N_2123);
nand U7225 (N_7225,N_3926,N_4382);
and U7226 (N_7226,N_1665,N_3210);
nor U7227 (N_7227,N_917,N_4525);
or U7228 (N_7228,N_111,N_3994);
nand U7229 (N_7229,N_226,N_3370);
or U7230 (N_7230,N_4168,N_166);
or U7231 (N_7231,N_4926,N_249);
nor U7232 (N_7232,N_1725,N_3414);
nor U7233 (N_7233,N_2567,N_2041);
nor U7234 (N_7234,N_371,N_2532);
nor U7235 (N_7235,N_4949,N_4569);
nand U7236 (N_7236,N_4087,N_2861);
nor U7237 (N_7237,N_678,N_1963);
and U7238 (N_7238,N_859,N_1996);
nor U7239 (N_7239,N_3627,N_4784);
xor U7240 (N_7240,N_4725,N_3234);
or U7241 (N_7241,N_3890,N_1172);
or U7242 (N_7242,N_507,N_852);
nand U7243 (N_7243,N_4080,N_3813);
and U7244 (N_7244,N_889,N_2837);
nand U7245 (N_7245,N_4983,N_911);
nand U7246 (N_7246,N_1572,N_2258);
nand U7247 (N_7247,N_339,N_898);
or U7248 (N_7248,N_2744,N_118);
or U7249 (N_7249,N_1420,N_3235);
and U7250 (N_7250,N_2527,N_1586);
nand U7251 (N_7251,N_944,N_2555);
nor U7252 (N_7252,N_4968,N_412);
or U7253 (N_7253,N_891,N_3629);
and U7254 (N_7254,N_4099,N_3173);
nor U7255 (N_7255,N_4661,N_702);
and U7256 (N_7256,N_3894,N_222);
nand U7257 (N_7257,N_3031,N_2764);
or U7258 (N_7258,N_1218,N_1903);
nor U7259 (N_7259,N_3685,N_3834);
or U7260 (N_7260,N_2783,N_3911);
nor U7261 (N_7261,N_4312,N_2060);
nor U7262 (N_7262,N_4867,N_4396);
nor U7263 (N_7263,N_3552,N_3709);
nor U7264 (N_7264,N_4646,N_2656);
nor U7265 (N_7265,N_1852,N_2504);
and U7266 (N_7266,N_1181,N_3947);
and U7267 (N_7267,N_459,N_2288);
and U7268 (N_7268,N_3275,N_977);
or U7269 (N_7269,N_4448,N_4209);
nor U7270 (N_7270,N_1022,N_4523);
or U7271 (N_7271,N_3444,N_4792);
nor U7272 (N_7272,N_2908,N_3827);
nand U7273 (N_7273,N_2275,N_4232);
and U7274 (N_7274,N_4619,N_1949);
nand U7275 (N_7275,N_2403,N_1065);
or U7276 (N_7276,N_2714,N_3371);
nor U7277 (N_7277,N_2482,N_514);
nand U7278 (N_7278,N_755,N_2677);
nand U7279 (N_7279,N_3588,N_3998);
nand U7280 (N_7280,N_1185,N_861);
or U7281 (N_7281,N_885,N_1775);
or U7282 (N_7282,N_3514,N_171);
nor U7283 (N_7283,N_663,N_2099);
and U7284 (N_7284,N_3214,N_4084);
or U7285 (N_7285,N_2811,N_1601);
or U7286 (N_7286,N_1057,N_1449);
and U7287 (N_7287,N_2007,N_3159);
or U7288 (N_7288,N_2093,N_4350);
and U7289 (N_7289,N_700,N_47);
nor U7290 (N_7290,N_3844,N_158);
nor U7291 (N_7291,N_1883,N_562);
nor U7292 (N_7292,N_4566,N_414);
or U7293 (N_7293,N_2203,N_2930);
nand U7294 (N_7294,N_3233,N_4319);
and U7295 (N_7295,N_1536,N_3467);
or U7296 (N_7296,N_1881,N_4704);
nand U7297 (N_7297,N_2493,N_212);
nor U7298 (N_7298,N_4965,N_3759);
and U7299 (N_7299,N_450,N_1307);
nand U7300 (N_7300,N_1046,N_1037);
nor U7301 (N_7301,N_3092,N_297);
nand U7302 (N_7302,N_184,N_1261);
and U7303 (N_7303,N_1956,N_1457);
nor U7304 (N_7304,N_3633,N_3174);
or U7305 (N_7305,N_3127,N_4827);
nor U7306 (N_7306,N_4033,N_3673);
and U7307 (N_7307,N_4567,N_194);
and U7308 (N_7308,N_4467,N_3712);
nand U7309 (N_7309,N_3292,N_3597);
nand U7310 (N_7310,N_815,N_3743);
nand U7311 (N_7311,N_1795,N_1306);
or U7312 (N_7312,N_1554,N_2160);
nand U7313 (N_7313,N_2147,N_1179);
nor U7314 (N_7314,N_3664,N_4625);
and U7315 (N_7315,N_4997,N_1712);
nor U7316 (N_7316,N_97,N_3484);
or U7317 (N_7317,N_4456,N_4535);
nand U7318 (N_7318,N_1015,N_684);
nand U7319 (N_7319,N_1784,N_1807);
or U7320 (N_7320,N_4199,N_1675);
or U7321 (N_7321,N_3500,N_3407);
and U7322 (N_7322,N_3302,N_1567);
nor U7323 (N_7323,N_3698,N_729);
or U7324 (N_7324,N_4919,N_3563);
nand U7325 (N_7325,N_366,N_4901);
or U7326 (N_7326,N_4733,N_2665);
nor U7327 (N_7327,N_1375,N_336);
nor U7328 (N_7328,N_190,N_972);
or U7329 (N_7329,N_3406,N_4806);
nand U7330 (N_7330,N_1267,N_2622);
or U7331 (N_7331,N_4769,N_4268);
or U7332 (N_7332,N_4474,N_2660);
or U7333 (N_7333,N_1650,N_289);
or U7334 (N_7334,N_742,N_1667);
and U7335 (N_7335,N_1614,N_2098);
nor U7336 (N_7336,N_749,N_4357);
or U7337 (N_7337,N_2188,N_1096);
nand U7338 (N_7338,N_2678,N_1165);
nor U7339 (N_7339,N_2133,N_4773);
nor U7340 (N_7340,N_1571,N_1489);
nor U7341 (N_7341,N_4093,N_4491);
and U7342 (N_7342,N_1083,N_318);
and U7343 (N_7343,N_4161,N_3744);
or U7344 (N_7344,N_1893,N_2769);
nor U7345 (N_7345,N_4062,N_2939);
or U7346 (N_7346,N_739,N_1871);
nor U7347 (N_7347,N_3172,N_4485);
nand U7348 (N_7348,N_3559,N_2341);
or U7349 (N_7349,N_1426,N_876);
or U7350 (N_7350,N_828,N_4864);
nor U7351 (N_7351,N_3431,N_34);
nand U7352 (N_7352,N_3391,N_3342);
or U7353 (N_7353,N_967,N_3553);
and U7354 (N_7354,N_979,N_3220);
and U7355 (N_7355,N_4527,N_1938);
or U7356 (N_7356,N_345,N_4252);
nor U7357 (N_7357,N_3178,N_17);
and U7358 (N_7358,N_1414,N_4551);
nor U7359 (N_7359,N_1294,N_149);
nand U7360 (N_7360,N_4064,N_4741);
and U7361 (N_7361,N_2729,N_1355);
or U7362 (N_7362,N_3702,N_2956);
or U7363 (N_7363,N_2424,N_2641);
and U7364 (N_7364,N_4236,N_2476);
or U7365 (N_7365,N_1901,N_3446);
nand U7366 (N_7366,N_1372,N_257);
and U7367 (N_7367,N_3492,N_3574);
and U7368 (N_7368,N_3405,N_2850);
nor U7369 (N_7369,N_448,N_3306);
and U7370 (N_7370,N_2654,N_115);
nor U7371 (N_7371,N_2825,N_3811);
nand U7372 (N_7372,N_4563,N_2992);
nor U7373 (N_7373,N_699,N_3967);
xor U7374 (N_7374,N_4050,N_3601);
and U7375 (N_7375,N_1138,N_3610);
and U7376 (N_7376,N_4017,N_4120);
nor U7377 (N_7377,N_4332,N_3710);
or U7378 (N_7378,N_3929,N_1407);
or U7379 (N_7379,N_4664,N_1296);
or U7380 (N_7380,N_1090,N_228);
or U7381 (N_7381,N_3090,N_3755);
nor U7382 (N_7382,N_3555,N_1502);
nor U7383 (N_7383,N_4840,N_1604);
nor U7384 (N_7384,N_2032,N_4436);
nand U7385 (N_7385,N_4673,N_3326);
or U7386 (N_7386,N_3033,N_4413);
or U7387 (N_7387,N_1440,N_823);
and U7388 (N_7388,N_877,N_4171);
nor U7389 (N_7389,N_2843,N_4264);
and U7390 (N_7390,N_1336,N_2156);
nand U7391 (N_7391,N_2163,N_946);
and U7392 (N_7392,N_100,N_878);
or U7393 (N_7393,N_3524,N_1992);
or U7394 (N_7394,N_1100,N_331);
nand U7395 (N_7395,N_3337,N_126);
nand U7396 (N_7396,N_4224,N_419);
or U7397 (N_7397,N_1697,N_1478);
nor U7398 (N_7398,N_1337,N_2264);
nand U7399 (N_7399,N_2854,N_635);
nand U7400 (N_7400,N_2519,N_3035);
nor U7401 (N_7401,N_114,N_4091);
nor U7402 (N_7402,N_4339,N_4271);
and U7403 (N_7403,N_1054,N_3700);
nand U7404 (N_7404,N_2520,N_3996);
or U7405 (N_7405,N_1345,N_1800);
and U7406 (N_7406,N_3992,N_2473);
or U7407 (N_7407,N_3442,N_992);
nor U7408 (N_7408,N_4617,N_3955);
and U7409 (N_7409,N_4170,N_1214);
or U7410 (N_7410,N_2535,N_2241);
nand U7411 (N_7411,N_3547,N_3315);
and U7412 (N_7412,N_4484,N_1797);
and U7413 (N_7413,N_1842,N_3958);
or U7414 (N_7414,N_1224,N_4470);
or U7415 (N_7415,N_3725,N_486);
and U7416 (N_7416,N_845,N_1612);
or U7417 (N_7417,N_1547,N_1452);
nand U7418 (N_7418,N_2023,N_4044);
or U7419 (N_7419,N_2260,N_3352);
or U7420 (N_7420,N_1018,N_464);
nor U7421 (N_7421,N_3587,N_513);
and U7422 (N_7422,N_2376,N_425);
nand U7423 (N_7423,N_2114,N_1351);
and U7424 (N_7424,N_883,N_3976);
or U7425 (N_7425,N_4255,N_4537);
nor U7426 (N_7426,N_326,N_3516);
nand U7427 (N_7427,N_601,N_3581);
nor U7428 (N_7428,N_3289,N_375);
or U7429 (N_7429,N_4395,N_2851);
nor U7430 (N_7430,N_2915,N_3752);
and U7431 (N_7431,N_3330,N_981);
nor U7432 (N_7432,N_1230,N_207);
or U7433 (N_7433,N_2582,N_116);
or U7434 (N_7434,N_953,N_2936);
or U7435 (N_7435,N_4135,N_1668);
and U7436 (N_7436,N_3777,N_595);
nor U7437 (N_7437,N_4089,N_4295);
and U7438 (N_7438,N_857,N_4263);
nor U7439 (N_7439,N_1143,N_4221);
and U7440 (N_7440,N_863,N_2650);
nor U7441 (N_7441,N_1299,N_4322);
nor U7442 (N_7442,N_4167,N_472);
nor U7443 (N_7443,N_733,N_3129);
and U7444 (N_7444,N_1494,N_1574);
nor U7445 (N_7445,N_1356,N_1162);
nor U7446 (N_7446,N_2179,N_68);
and U7447 (N_7447,N_285,N_3394);
nor U7448 (N_7448,N_2155,N_4746);
nand U7449 (N_7449,N_3734,N_4633);
nor U7450 (N_7450,N_162,N_4105);
and U7451 (N_7451,N_2299,N_3666);
and U7452 (N_7452,N_1012,N_1546);
and U7453 (N_7453,N_4437,N_670);
or U7454 (N_7454,N_653,N_3749);
and U7455 (N_7455,N_3536,N_2898);
and U7456 (N_7456,N_1758,N_201);
nor U7457 (N_7457,N_4665,N_3952);
nor U7458 (N_7458,N_2722,N_1884);
nand U7459 (N_7459,N_4931,N_4682);
or U7460 (N_7460,N_4521,N_3312);
or U7461 (N_7461,N_998,N_2737);
or U7462 (N_7462,N_2559,N_3211);
nand U7463 (N_7463,N_3141,N_231);
nand U7464 (N_7464,N_1569,N_1755);
or U7465 (N_7465,N_580,N_2013);
and U7466 (N_7466,N_2984,N_3260);
or U7467 (N_7467,N_4705,N_3480);
and U7468 (N_7468,N_4346,N_131);
and U7469 (N_7469,N_3981,N_4941);
nand U7470 (N_7470,N_1699,N_831);
or U7471 (N_7471,N_3854,N_3348);
or U7472 (N_7472,N_4729,N_1215);
and U7473 (N_7473,N_4311,N_4638);
and U7474 (N_7474,N_1512,N_4164);
nand U7475 (N_7475,N_613,N_539);
nand U7476 (N_7476,N_961,N_1664);
nor U7477 (N_7477,N_4871,N_1025);
and U7478 (N_7478,N_3373,N_1077);
or U7479 (N_7479,N_3060,N_677);
nor U7480 (N_7480,N_235,N_2780);
and U7481 (N_7481,N_369,N_1063);
and U7482 (N_7482,N_3171,N_2335);
and U7483 (N_7483,N_3928,N_1765);
or U7484 (N_7484,N_2116,N_761);
or U7485 (N_7485,N_4438,N_1743);
and U7486 (N_7486,N_3366,N_1748);
nor U7487 (N_7487,N_1859,N_3808);
or U7488 (N_7488,N_1545,N_3704);
or U7489 (N_7489,N_4911,N_4863);
nand U7490 (N_7490,N_213,N_4206);
or U7491 (N_7491,N_1273,N_3495);
and U7492 (N_7492,N_356,N_3884);
and U7493 (N_7493,N_650,N_3762);
or U7494 (N_7494,N_1661,N_2901);
and U7495 (N_7495,N_1981,N_4721);
nor U7496 (N_7496,N_4400,N_3945);
and U7497 (N_7497,N_2997,N_466);
nand U7498 (N_7498,N_1262,N_1052);
nor U7499 (N_7499,N_243,N_780);
or U7500 (N_7500,N_4996,N_1098);
nor U7501 (N_7501,N_4911,N_4246);
nor U7502 (N_7502,N_3605,N_3924);
nand U7503 (N_7503,N_4109,N_307);
and U7504 (N_7504,N_4599,N_1991);
nor U7505 (N_7505,N_4710,N_2979);
or U7506 (N_7506,N_602,N_1542);
or U7507 (N_7507,N_3721,N_910);
or U7508 (N_7508,N_1284,N_2618);
or U7509 (N_7509,N_2087,N_4515);
or U7510 (N_7510,N_1778,N_10);
nor U7511 (N_7511,N_87,N_2900);
nor U7512 (N_7512,N_4584,N_1314);
and U7513 (N_7513,N_1157,N_2097);
nor U7514 (N_7514,N_2173,N_4310);
nand U7515 (N_7515,N_2013,N_984);
and U7516 (N_7516,N_2038,N_4129);
nor U7517 (N_7517,N_4390,N_3717);
nand U7518 (N_7518,N_2725,N_1898);
or U7519 (N_7519,N_1576,N_1744);
or U7520 (N_7520,N_2002,N_3885);
nor U7521 (N_7521,N_1719,N_2961);
nor U7522 (N_7522,N_1736,N_3183);
and U7523 (N_7523,N_4950,N_1076);
and U7524 (N_7524,N_2252,N_4767);
or U7525 (N_7525,N_2134,N_3390);
or U7526 (N_7526,N_4062,N_179);
and U7527 (N_7527,N_4295,N_2231);
nand U7528 (N_7528,N_2884,N_315);
nand U7529 (N_7529,N_4099,N_4349);
nor U7530 (N_7530,N_1662,N_4446);
and U7531 (N_7531,N_48,N_1171);
and U7532 (N_7532,N_3466,N_3784);
nand U7533 (N_7533,N_1393,N_282);
and U7534 (N_7534,N_2381,N_324);
nand U7535 (N_7535,N_1419,N_3969);
or U7536 (N_7536,N_4117,N_3028);
or U7537 (N_7537,N_3047,N_823);
or U7538 (N_7538,N_3939,N_469);
nor U7539 (N_7539,N_2165,N_1829);
nor U7540 (N_7540,N_3880,N_4419);
and U7541 (N_7541,N_3451,N_1719);
nor U7542 (N_7542,N_2436,N_1823);
and U7543 (N_7543,N_2812,N_1113);
or U7544 (N_7544,N_2918,N_2025);
and U7545 (N_7545,N_2851,N_1501);
or U7546 (N_7546,N_4058,N_331);
and U7547 (N_7547,N_204,N_2130);
or U7548 (N_7548,N_1906,N_2093);
nand U7549 (N_7549,N_3927,N_4089);
nand U7550 (N_7550,N_4594,N_4212);
nand U7551 (N_7551,N_4646,N_1203);
and U7552 (N_7552,N_2106,N_574);
and U7553 (N_7553,N_3567,N_906);
nand U7554 (N_7554,N_2038,N_1613);
nor U7555 (N_7555,N_935,N_1401);
and U7556 (N_7556,N_3088,N_2928);
nand U7557 (N_7557,N_3641,N_83);
and U7558 (N_7558,N_308,N_186);
and U7559 (N_7559,N_4425,N_4972);
nor U7560 (N_7560,N_1104,N_4521);
and U7561 (N_7561,N_4437,N_4907);
or U7562 (N_7562,N_2754,N_4018);
and U7563 (N_7563,N_1637,N_4688);
nand U7564 (N_7564,N_1394,N_629);
nand U7565 (N_7565,N_680,N_2743);
nand U7566 (N_7566,N_3730,N_4682);
nand U7567 (N_7567,N_4148,N_1129);
or U7568 (N_7568,N_1537,N_2812);
and U7569 (N_7569,N_2477,N_3735);
and U7570 (N_7570,N_2059,N_345);
nand U7571 (N_7571,N_731,N_4162);
and U7572 (N_7572,N_3216,N_419);
nand U7573 (N_7573,N_2157,N_3943);
nand U7574 (N_7574,N_899,N_4050);
nor U7575 (N_7575,N_3500,N_138);
nand U7576 (N_7576,N_2259,N_4477);
or U7577 (N_7577,N_713,N_1559);
and U7578 (N_7578,N_1034,N_3390);
or U7579 (N_7579,N_1946,N_3853);
nand U7580 (N_7580,N_1772,N_811);
nand U7581 (N_7581,N_2090,N_1872);
and U7582 (N_7582,N_1822,N_1837);
or U7583 (N_7583,N_2533,N_3707);
nor U7584 (N_7584,N_4351,N_118);
nand U7585 (N_7585,N_2095,N_3835);
and U7586 (N_7586,N_1443,N_2907);
nor U7587 (N_7587,N_3519,N_306);
or U7588 (N_7588,N_2530,N_3704);
nor U7589 (N_7589,N_3129,N_4320);
and U7590 (N_7590,N_2711,N_4840);
and U7591 (N_7591,N_595,N_2517);
nor U7592 (N_7592,N_4993,N_2891);
or U7593 (N_7593,N_4719,N_1332);
and U7594 (N_7594,N_1885,N_520);
and U7595 (N_7595,N_2876,N_1596);
or U7596 (N_7596,N_1206,N_4806);
nor U7597 (N_7597,N_1761,N_4556);
nor U7598 (N_7598,N_1805,N_4979);
nand U7599 (N_7599,N_3303,N_3793);
and U7600 (N_7600,N_1609,N_173);
nor U7601 (N_7601,N_2672,N_3817);
nand U7602 (N_7602,N_3236,N_4220);
or U7603 (N_7603,N_2320,N_3884);
nand U7604 (N_7604,N_708,N_3338);
and U7605 (N_7605,N_2351,N_2933);
or U7606 (N_7606,N_1109,N_4110);
and U7607 (N_7607,N_2521,N_348);
nand U7608 (N_7608,N_777,N_3549);
and U7609 (N_7609,N_2469,N_3897);
nor U7610 (N_7610,N_1960,N_1941);
or U7611 (N_7611,N_2664,N_1794);
nand U7612 (N_7612,N_1346,N_3339);
nor U7613 (N_7613,N_295,N_237);
and U7614 (N_7614,N_3722,N_4658);
or U7615 (N_7615,N_2301,N_1462);
or U7616 (N_7616,N_1236,N_473);
nand U7617 (N_7617,N_4016,N_2570);
nor U7618 (N_7618,N_182,N_813);
and U7619 (N_7619,N_2212,N_4360);
nor U7620 (N_7620,N_525,N_2458);
and U7621 (N_7621,N_1682,N_1727);
and U7622 (N_7622,N_721,N_4327);
or U7623 (N_7623,N_4819,N_1842);
or U7624 (N_7624,N_696,N_4439);
nor U7625 (N_7625,N_2934,N_4406);
or U7626 (N_7626,N_4867,N_3036);
and U7627 (N_7627,N_876,N_2767);
and U7628 (N_7628,N_3243,N_1552);
nand U7629 (N_7629,N_3690,N_2496);
or U7630 (N_7630,N_3755,N_4193);
or U7631 (N_7631,N_2317,N_2548);
or U7632 (N_7632,N_3562,N_135);
nor U7633 (N_7633,N_2733,N_2830);
nor U7634 (N_7634,N_3599,N_4462);
nor U7635 (N_7635,N_4465,N_4157);
nor U7636 (N_7636,N_4346,N_1446);
nand U7637 (N_7637,N_3404,N_1012);
xnor U7638 (N_7638,N_1868,N_1243);
nand U7639 (N_7639,N_464,N_1197);
nand U7640 (N_7640,N_3416,N_1656);
nor U7641 (N_7641,N_4606,N_3063);
and U7642 (N_7642,N_2231,N_4850);
nand U7643 (N_7643,N_965,N_151);
nor U7644 (N_7644,N_4789,N_3005);
and U7645 (N_7645,N_4724,N_659);
nand U7646 (N_7646,N_4966,N_3092);
or U7647 (N_7647,N_2524,N_3745);
nand U7648 (N_7648,N_4861,N_2702);
or U7649 (N_7649,N_4282,N_21);
nand U7650 (N_7650,N_4755,N_2900);
and U7651 (N_7651,N_3016,N_2582);
or U7652 (N_7652,N_2112,N_4488);
or U7653 (N_7653,N_2275,N_3471);
nor U7654 (N_7654,N_2270,N_4248);
or U7655 (N_7655,N_1148,N_777);
and U7656 (N_7656,N_2054,N_3797);
and U7657 (N_7657,N_3356,N_668);
nand U7658 (N_7658,N_1424,N_2798);
xor U7659 (N_7659,N_3585,N_3537);
and U7660 (N_7660,N_541,N_2394);
and U7661 (N_7661,N_2523,N_4731);
or U7662 (N_7662,N_3012,N_2604);
or U7663 (N_7663,N_3868,N_2438);
nand U7664 (N_7664,N_1450,N_2239);
and U7665 (N_7665,N_2242,N_1603);
nand U7666 (N_7666,N_1764,N_3703);
nor U7667 (N_7667,N_4720,N_3600);
nor U7668 (N_7668,N_2842,N_1129);
nand U7669 (N_7669,N_1048,N_4556);
nor U7670 (N_7670,N_2120,N_4503);
and U7671 (N_7671,N_2209,N_551);
nor U7672 (N_7672,N_1339,N_4909);
or U7673 (N_7673,N_1148,N_3339);
and U7674 (N_7674,N_1505,N_4264);
nor U7675 (N_7675,N_3922,N_3017);
nand U7676 (N_7676,N_2961,N_2685);
nor U7677 (N_7677,N_3611,N_624);
or U7678 (N_7678,N_3946,N_4747);
nor U7679 (N_7679,N_3896,N_4489);
nor U7680 (N_7680,N_2853,N_2226);
nand U7681 (N_7681,N_3583,N_4384);
nor U7682 (N_7682,N_698,N_3012);
nor U7683 (N_7683,N_1170,N_4120);
and U7684 (N_7684,N_4077,N_3712);
or U7685 (N_7685,N_3594,N_1663);
nand U7686 (N_7686,N_2927,N_3685);
nand U7687 (N_7687,N_934,N_2758);
nor U7688 (N_7688,N_367,N_1840);
or U7689 (N_7689,N_1989,N_2514);
or U7690 (N_7690,N_2899,N_455);
nor U7691 (N_7691,N_2774,N_2008);
or U7692 (N_7692,N_3767,N_3684);
and U7693 (N_7693,N_3956,N_3933);
nor U7694 (N_7694,N_4951,N_1616);
or U7695 (N_7695,N_2757,N_2667);
nand U7696 (N_7696,N_3098,N_1251);
and U7697 (N_7697,N_1050,N_1372);
or U7698 (N_7698,N_288,N_2435);
or U7699 (N_7699,N_3209,N_1584);
or U7700 (N_7700,N_4105,N_2769);
and U7701 (N_7701,N_3001,N_378);
nand U7702 (N_7702,N_3797,N_4644);
and U7703 (N_7703,N_4975,N_1968);
or U7704 (N_7704,N_1046,N_162);
nor U7705 (N_7705,N_1767,N_1395);
nor U7706 (N_7706,N_4097,N_4340);
nand U7707 (N_7707,N_2970,N_547);
nand U7708 (N_7708,N_784,N_499);
and U7709 (N_7709,N_4743,N_37);
or U7710 (N_7710,N_336,N_3027);
or U7711 (N_7711,N_1325,N_179);
nand U7712 (N_7712,N_857,N_4638);
or U7713 (N_7713,N_1759,N_4725);
and U7714 (N_7714,N_1715,N_523);
and U7715 (N_7715,N_2258,N_4035);
and U7716 (N_7716,N_2480,N_63);
and U7717 (N_7717,N_927,N_706);
nor U7718 (N_7718,N_876,N_1143);
nor U7719 (N_7719,N_2811,N_2076);
nor U7720 (N_7720,N_2006,N_1204);
nor U7721 (N_7721,N_3052,N_4300);
and U7722 (N_7722,N_1768,N_2301);
or U7723 (N_7723,N_369,N_1820);
or U7724 (N_7724,N_1760,N_3359);
nand U7725 (N_7725,N_1875,N_3645);
or U7726 (N_7726,N_3792,N_3587);
and U7727 (N_7727,N_4824,N_2413);
and U7728 (N_7728,N_4696,N_3424);
nand U7729 (N_7729,N_570,N_3935);
or U7730 (N_7730,N_2088,N_3983);
nand U7731 (N_7731,N_35,N_3766);
or U7732 (N_7732,N_4003,N_3446);
nand U7733 (N_7733,N_2413,N_4894);
nand U7734 (N_7734,N_3490,N_1028);
or U7735 (N_7735,N_2443,N_3084);
and U7736 (N_7736,N_4873,N_1341);
nor U7737 (N_7737,N_1273,N_4615);
nor U7738 (N_7738,N_42,N_4522);
and U7739 (N_7739,N_4328,N_1313);
and U7740 (N_7740,N_3183,N_1092);
nand U7741 (N_7741,N_3557,N_3040);
nand U7742 (N_7742,N_3635,N_710);
or U7743 (N_7743,N_32,N_1057);
or U7744 (N_7744,N_2414,N_3962);
or U7745 (N_7745,N_1784,N_3033);
nor U7746 (N_7746,N_2319,N_3372);
nand U7747 (N_7747,N_1833,N_4611);
nor U7748 (N_7748,N_282,N_710);
and U7749 (N_7749,N_541,N_1412);
nand U7750 (N_7750,N_1134,N_4811);
or U7751 (N_7751,N_1789,N_2477);
nand U7752 (N_7752,N_4280,N_1803);
nand U7753 (N_7753,N_4068,N_4903);
nand U7754 (N_7754,N_4459,N_1314);
nor U7755 (N_7755,N_823,N_4769);
nand U7756 (N_7756,N_4908,N_4784);
nor U7757 (N_7757,N_4138,N_4410);
or U7758 (N_7758,N_3182,N_3413);
nand U7759 (N_7759,N_4144,N_3005);
or U7760 (N_7760,N_4205,N_243);
nor U7761 (N_7761,N_811,N_444);
nand U7762 (N_7762,N_2732,N_3775);
or U7763 (N_7763,N_1347,N_3377);
and U7764 (N_7764,N_1716,N_917);
nor U7765 (N_7765,N_3820,N_3075);
and U7766 (N_7766,N_2543,N_922);
nor U7767 (N_7767,N_1591,N_4383);
xnor U7768 (N_7768,N_335,N_4339);
nor U7769 (N_7769,N_3617,N_4397);
or U7770 (N_7770,N_417,N_3769);
nand U7771 (N_7771,N_790,N_1726);
nor U7772 (N_7772,N_1552,N_3081);
nand U7773 (N_7773,N_2031,N_1448);
xor U7774 (N_7774,N_143,N_3945);
nor U7775 (N_7775,N_98,N_4077);
or U7776 (N_7776,N_605,N_2296);
nor U7777 (N_7777,N_2348,N_347);
nor U7778 (N_7778,N_381,N_4077);
nand U7779 (N_7779,N_586,N_1776);
or U7780 (N_7780,N_1974,N_2267);
or U7781 (N_7781,N_339,N_2784);
and U7782 (N_7782,N_3866,N_1364);
nor U7783 (N_7783,N_4343,N_2555);
nand U7784 (N_7784,N_4821,N_3532);
or U7785 (N_7785,N_2426,N_316);
and U7786 (N_7786,N_1070,N_4956);
and U7787 (N_7787,N_3595,N_2986);
or U7788 (N_7788,N_828,N_1563);
or U7789 (N_7789,N_3017,N_4446);
nor U7790 (N_7790,N_4090,N_4569);
and U7791 (N_7791,N_4647,N_1268);
nor U7792 (N_7792,N_1503,N_1075);
nor U7793 (N_7793,N_230,N_1738);
and U7794 (N_7794,N_3397,N_2417);
nor U7795 (N_7795,N_3332,N_4179);
nor U7796 (N_7796,N_4243,N_2714);
nor U7797 (N_7797,N_658,N_299);
nor U7798 (N_7798,N_4900,N_163);
and U7799 (N_7799,N_3808,N_4717);
and U7800 (N_7800,N_4390,N_2871);
nor U7801 (N_7801,N_2765,N_207);
or U7802 (N_7802,N_2309,N_2655);
nand U7803 (N_7803,N_3273,N_4622);
nor U7804 (N_7804,N_81,N_4566);
or U7805 (N_7805,N_4269,N_353);
and U7806 (N_7806,N_4305,N_4844);
nand U7807 (N_7807,N_1713,N_4144);
nor U7808 (N_7808,N_2217,N_3941);
or U7809 (N_7809,N_794,N_1567);
nand U7810 (N_7810,N_4080,N_4915);
or U7811 (N_7811,N_180,N_4454);
nor U7812 (N_7812,N_2599,N_2356);
or U7813 (N_7813,N_4356,N_2761);
nand U7814 (N_7814,N_3190,N_3573);
nor U7815 (N_7815,N_1583,N_706);
and U7816 (N_7816,N_485,N_1229);
and U7817 (N_7817,N_3198,N_1378);
nand U7818 (N_7818,N_241,N_4904);
and U7819 (N_7819,N_4894,N_4913);
or U7820 (N_7820,N_4675,N_4588);
nand U7821 (N_7821,N_4948,N_886);
nor U7822 (N_7822,N_4224,N_1413);
nor U7823 (N_7823,N_3186,N_3742);
or U7824 (N_7824,N_3145,N_2298);
or U7825 (N_7825,N_1524,N_3913);
nor U7826 (N_7826,N_1190,N_491);
nand U7827 (N_7827,N_2416,N_3612);
or U7828 (N_7828,N_4882,N_2759);
or U7829 (N_7829,N_4144,N_3948);
or U7830 (N_7830,N_4376,N_2921);
nor U7831 (N_7831,N_4495,N_756);
or U7832 (N_7832,N_1185,N_66);
nor U7833 (N_7833,N_2608,N_551);
nor U7834 (N_7834,N_3925,N_105);
nand U7835 (N_7835,N_3411,N_1488);
nand U7836 (N_7836,N_2184,N_436);
or U7837 (N_7837,N_174,N_4528);
or U7838 (N_7838,N_309,N_1244);
and U7839 (N_7839,N_3765,N_337);
and U7840 (N_7840,N_1110,N_2999);
or U7841 (N_7841,N_3517,N_3273);
nand U7842 (N_7842,N_4595,N_3137);
nand U7843 (N_7843,N_4842,N_296);
nand U7844 (N_7844,N_4697,N_3757);
or U7845 (N_7845,N_2309,N_1364);
or U7846 (N_7846,N_1220,N_1931);
nor U7847 (N_7847,N_4456,N_4528);
nand U7848 (N_7848,N_812,N_1587);
and U7849 (N_7849,N_3765,N_3795);
and U7850 (N_7850,N_2176,N_4054);
nand U7851 (N_7851,N_4317,N_2258);
nand U7852 (N_7852,N_1736,N_3506);
nand U7853 (N_7853,N_139,N_2376);
nand U7854 (N_7854,N_4659,N_4760);
nor U7855 (N_7855,N_2567,N_1972);
nor U7856 (N_7856,N_2570,N_1284);
nor U7857 (N_7857,N_1678,N_503);
nand U7858 (N_7858,N_2208,N_4672);
xor U7859 (N_7859,N_4164,N_2408);
or U7860 (N_7860,N_1650,N_3839);
nor U7861 (N_7861,N_1723,N_1425);
nand U7862 (N_7862,N_2357,N_2727);
and U7863 (N_7863,N_402,N_4453);
and U7864 (N_7864,N_3972,N_2734);
nand U7865 (N_7865,N_586,N_4362);
and U7866 (N_7866,N_3511,N_3913);
nand U7867 (N_7867,N_3411,N_4847);
and U7868 (N_7868,N_4270,N_4707);
and U7869 (N_7869,N_221,N_2529);
nand U7870 (N_7870,N_3204,N_4885);
or U7871 (N_7871,N_603,N_4409);
or U7872 (N_7872,N_2458,N_401);
nor U7873 (N_7873,N_3385,N_4224);
and U7874 (N_7874,N_4859,N_759);
nor U7875 (N_7875,N_3862,N_2523);
or U7876 (N_7876,N_864,N_97);
and U7877 (N_7877,N_1924,N_3609);
and U7878 (N_7878,N_4482,N_702);
or U7879 (N_7879,N_3670,N_1853);
nand U7880 (N_7880,N_1778,N_4981);
nand U7881 (N_7881,N_4641,N_3301);
nand U7882 (N_7882,N_4580,N_892);
and U7883 (N_7883,N_3457,N_1550);
nand U7884 (N_7884,N_2844,N_508);
and U7885 (N_7885,N_611,N_4502);
nor U7886 (N_7886,N_1516,N_792);
nor U7887 (N_7887,N_2613,N_263);
or U7888 (N_7888,N_2883,N_4083);
nand U7889 (N_7889,N_3331,N_2498);
nor U7890 (N_7890,N_4146,N_2064);
and U7891 (N_7891,N_3688,N_3279);
or U7892 (N_7892,N_1989,N_3292);
nand U7893 (N_7893,N_4754,N_2783);
or U7894 (N_7894,N_744,N_3163);
and U7895 (N_7895,N_3450,N_406);
and U7896 (N_7896,N_1228,N_4769);
or U7897 (N_7897,N_3401,N_1366);
and U7898 (N_7898,N_1494,N_3585);
and U7899 (N_7899,N_1244,N_2624);
and U7900 (N_7900,N_3427,N_303);
nand U7901 (N_7901,N_623,N_2501);
or U7902 (N_7902,N_1252,N_3300);
nand U7903 (N_7903,N_2992,N_4818);
or U7904 (N_7904,N_81,N_501);
nand U7905 (N_7905,N_3526,N_439);
nor U7906 (N_7906,N_1049,N_2442);
and U7907 (N_7907,N_872,N_780);
or U7908 (N_7908,N_4390,N_428);
nand U7909 (N_7909,N_2107,N_4508);
or U7910 (N_7910,N_2641,N_839);
nand U7911 (N_7911,N_4802,N_1925);
or U7912 (N_7912,N_255,N_3468);
and U7913 (N_7913,N_1844,N_4060);
and U7914 (N_7914,N_4591,N_508);
and U7915 (N_7915,N_780,N_2643);
and U7916 (N_7916,N_1561,N_211);
nand U7917 (N_7917,N_3340,N_3254);
or U7918 (N_7918,N_4713,N_4744);
nor U7919 (N_7919,N_852,N_1018);
or U7920 (N_7920,N_3708,N_1732);
nand U7921 (N_7921,N_4531,N_3935);
nand U7922 (N_7922,N_3669,N_2862);
nand U7923 (N_7923,N_1684,N_459);
nor U7924 (N_7924,N_3754,N_470);
nor U7925 (N_7925,N_3847,N_219);
nand U7926 (N_7926,N_3815,N_2889);
and U7927 (N_7927,N_3924,N_1759);
nand U7928 (N_7928,N_3762,N_3165);
nand U7929 (N_7929,N_4701,N_4713);
or U7930 (N_7930,N_3330,N_1698);
nor U7931 (N_7931,N_1298,N_550);
nor U7932 (N_7932,N_4389,N_4959);
or U7933 (N_7933,N_2328,N_580);
or U7934 (N_7934,N_2178,N_305);
nand U7935 (N_7935,N_1286,N_1435);
nand U7936 (N_7936,N_1340,N_2276);
and U7937 (N_7937,N_1710,N_4917);
and U7938 (N_7938,N_543,N_1048);
and U7939 (N_7939,N_1616,N_1698);
or U7940 (N_7940,N_2646,N_3500);
and U7941 (N_7941,N_1669,N_4222);
or U7942 (N_7942,N_3510,N_3797);
nor U7943 (N_7943,N_3064,N_940);
nor U7944 (N_7944,N_3208,N_2342);
nor U7945 (N_7945,N_3194,N_4182);
nand U7946 (N_7946,N_4779,N_2009);
nand U7947 (N_7947,N_4585,N_713);
nand U7948 (N_7948,N_2091,N_248);
nor U7949 (N_7949,N_695,N_878);
nand U7950 (N_7950,N_3496,N_4268);
nor U7951 (N_7951,N_2561,N_3781);
nor U7952 (N_7952,N_782,N_4760);
and U7953 (N_7953,N_4005,N_4125);
nor U7954 (N_7954,N_121,N_580);
nand U7955 (N_7955,N_1826,N_3903);
nand U7956 (N_7956,N_2096,N_4300);
or U7957 (N_7957,N_2910,N_2877);
nand U7958 (N_7958,N_132,N_4302);
or U7959 (N_7959,N_2517,N_2126);
and U7960 (N_7960,N_1021,N_4111);
and U7961 (N_7961,N_4384,N_1273);
or U7962 (N_7962,N_4126,N_485);
and U7963 (N_7963,N_1046,N_4997);
or U7964 (N_7964,N_3814,N_1399);
nor U7965 (N_7965,N_3088,N_2360);
nor U7966 (N_7966,N_4904,N_1295);
nand U7967 (N_7967,N_2718,N_1432);
nor U7968 (N_7968,N_539,N_562);
nor U7969 (N_7969,N_4118,N_3733);
nor U7970 (N_7970,N_1977,N_611);
or U7971 (N_7971,N_4940,N_4221);
and U7972 (N_7972,N_4706,N_835);
nor U7973 (N_7973,N_4324,N_429);
and U7974 (N_7974,N_1434,N_4308);
and U7975 (N_7975,N_1429,N_3772);
and U7976 (N_7976,N_2620,N_1911);
and U7977 (N_7977,N_914,N_164);
nor U7978 (N_7978,N_1900,N_2629);
or U7979 (N_7979,N_2200,N_885);
nand U7980 (N_7980,N_4863,N_2271);
nand U7981 (N_7981,N_1992,N_2792);
nand U7982 (N_7982,N_973,N_1049);
or U7983 (N_7983,N_2224,N_412);
nor U7984 (N_7984,N_839,N_4734);
nor U7985 (N_7985,N_1613,N_241);
nand U7986 (N_7986,N_4632,N_3371);
nor U7987 (N_7987,N_1645,N_2940);
or U7988 (N_7988,N_3423,N_3741);
nand U7989 (N_7989,N_2996,N_2754);
or U7990 (N_7990,N_3543,N_3619);
or U7991 (N_7991,N_3889,N_899);
or U7992 (N_7992,N_810,N_1229);
and U7993 (N_7993,N_4507,N_4754);
nand U7994 (N_7994,N_2722,N_3019);
nor U7995 (N_7995,N_3662,N_357);
or U7996 (N_7996,N_1209,N_4074);
nor U7997 (N_7997,N_2321,N_4345);
nor U7998 (N_7998,N_3324,N_4507);
nand U7999 (N_7999,N_3736,N_1603);
nor U8000 (N_8000,N_3106,N_3390);
and U8001 (N_8001,N_250,N_2072);
or U8002 (N_8002,N_2666,N_1162);
and U8003 (N_8003,N_3899,N_2813);
nor U8004 (N_8004,N_2494,N_3043);
or U8005 (N_8005,N_3304,N_2903);
nand U8006 (N_8006,N_2842,N_2702);
and U8007 (N_8007,N_4890,N_2227);
or U8008 (N_8008,N_2186,N_4179);
or U8009 (N_8009,N_3577,N_3044);
nor U8010 (N_8010,N_4603,N_4099);
or U8011 (N_8011,N_743,N_2740);
nand U8012 (N_8012,N_2132,N_1185);
and U8013 (N_8013,N_718,N_1021);
nand U8014 (N_8014,N_199,N_4223);
and U8015 (N_8015,N_4199,N_4274);
nand U8016 (N_8016,N_4984,N_3440);
or U8017 (N_8017,N_825,N_1692);
or U8018 (N_8018,N_902,N_3646);
or U8019 (N_8019,N_1482,N_4194);
and U8020 (N_8020,N_2281,N_2316);
nor U8021 (N_8021,N_2521,N_3535);
nand U8022 (N_8022,N_260,N_4900);
nor U8023 (N_8023,N_3446,N_3931);
and U8024 (N_8024,N_623,N_965);
nor U8025 (N_8025,N_1397,N_2175);
nand U8026 (N_8026,N_4954,N_2097);
nand U8027 (N_8027,N_4496,N_872);
nand U8028 (N_8028,N_1393,N_2977);
or U8029 (N_8029,N_2280,N_3207);
and U8030 (N_8030,N_2252,N_52);
nor U8031 (N_8031,N_712,N_993);
or U8032 (N_8032,N_2764,N_4077);
and U8033 (N_8033,N_483,N_3319);
nand U8034 (N_8034,N_930,N_2447);
nor U8035 (N_8035,N_4173,N_274);
nand U8036 (N_8036,N_4468,N_313);
or U8037 (N_8037,N_4799,N_2076);
nor U8038 (N_8038,N_2826,N_1135);
or U8039 (N_8039,N_3287,N_1421);
and U8040 (N_8040,N_4282,N_4210);
or U8041 (N_8041,N_783,N_275);
nand U8042 (N_8042,N_341,N_3091);
or U8043 (N_8043,N_1643,N_3903);
nand U8044 (N_8044,N_3283,N_4815);
or U8045 (N_8045,N_2166,N_1342);
or U8046 (N_8046,N_3453,N_633);
or U8047 (N_8047,N_1599,N_4109);
nand U8048 (N_8048,N_2771,N_591);
or U8049 (N_8049,N_1586,N_774);
or U8050 (N_8050,N_2409,N_235);
nor U8051 (N_8051,N_244,N_1064);
nor U8052 (N_8052,N_4354,N_3699);
or U8053 (N_8053,N_2559,N_4039);
nor U8054 (N_8054,N_3302,N_2924);
nand U8055 (N_8055,N_252,N_1272);
and U8056 (N_8056,N_2884,N_4964);
nor U8057 (N_8057,N_1139,N_451);
nand U8058 (N_8058,N_1839,N_3354);
or U8059 (N_8059,N_2941,N_3561);
and U8060 (N_8060,N_4914,N_2536);
and U8061 (N_8061,N_2440,N_525);
or U8062 (N_8062,N_3585,N_4474);
and U8063 (N_8063,N_336,N_3925);
nand U8064 (N_8064,N_2979,N_1119);
nand U8065 (N_8065,N_3004,N_4697);
nand U8066 (N_8066,N_2001,N_2666);
or U8067 (N_8067,N_2474,N_1247);
nand U8068 (N_8068,N_4578,N_3515);
nand U8069 (N_8069,N_3072,N_2336);
or U8070 (N_8070,N_3377,N_477);
or U8071 (N_8071,N_4518,N_2089);
nor U8072 (N_8072,N_4708,N_1226);
or U8073 (N_8073,N_4279,N_4362);
nor U8074 (N_8074,N_2458,N_1529);
or U8075 (N_8075,N_1639,N_1243);
or U8076 (N_8076,N_3719,N_1821);
or U8077 (N_8077,N_4764,N_564);
nand U8078 (N_8078,N_461,N_4111);
nor U8079 (N_8079,N_2316,N_2994);
nor U8080 (N_8080,N_4928,N_301);
or U8081 (N_8081,N_2720,N_1185);
nor U8082 (N_8082,N_3018,N_723);
nand U8083 (N_8083,N_4830,N_3854);
nand U8084 (N_8084,N_2359,N_4549);
and U8085 (N_8085,N_3120,N_4201);
nand U8086 (N_8086,N_3311,N_3967);
and U8087 (N_8087,N_1109,N_4835);
nand U8088 (N_8088,N_1541,N_4898);
or U8089 (N_8089,N_764,N_4178);
nand U8090 (N_8090,N_681,N_3511);
nand U8091 (N_8091,N_1531,N_106);
nand U8092 (N_8092,N_3090,N_2335);
nor U8093 (N_8093,N_4465,N_2767);
nor U8094 (N_8094,N_2680,N_2027);
and U8095 (N_8095,N_3925,N_1493);
and U8096 (N_8096,N_4112,N_896);
or U8097 (N_8097,N_4156,N_4423);
or U8098 (N_8098,N_1189,N_1590);
nand U8099 (N_8099,N_2436,N_4442);
or U8100 (N_8100,N_167,N_295);
or U8101 (N_8101,N_1671,N_1629);
and U8102 (N_8102,N_1587,N_3092);
and U8103 (N_8103,N_2248,N_3629);
or U8104 (N_8104,N_928,N_2537);
nor U8105 (N_8105,N_2417,N_4076);
and U8106 (N_8106,N_1155,N_1087);
nor U8107 (N_8107,N_2471,N_256);
nor U8108 (N_8108,N_3480,N_2147);
nand U8109 (N_8109,N_4634,N_2136);
nor U8110 (N_8110,N_4367,N_81);
or U8111 (N_8111,N_3008,N_1413);
or U8112 (N_8112,N_2469,N_970);
and U8113 (N_8113,N_3294,N_1192);
nor U8114 (N_8114,N_1117,N_190);
or U8115 (N_8115,N_3527,N_2669);
or U8116 (N_8116,N_2159,N_2925);
nor U8117 (N_8117,N_4940,N_4489);
or U8118 (N_8118,N_4878,N_2772);
nand U8119 (N_8119,N_4054,N_1957);
or U8120 (N_8120,N_1064,N_1483);
or U8121 (N_8121,N_606,N_4205);
and U8122 (N_8122,N_4640,N_419);
and U8123 (N_8123,N_666,N_4334);
nor U8124 (N_8124,N_4719,N_338);
nor U8125 (N_8125,N_1104,N_1307);
xnor U8126 (N_8126,N_4501,N_3493);
and U8127 (N_8127,N_871,N_3240);
or U8128 (N_8128,N_4079,N_4602);
nor U8129 (N_8129,N_1941,N_1177);
nor U8130 (N_8130,N_3478,N_2469);
and U8131 (N_8131,N_2115,N_101);
or U8132 (N_8132,N_4408,N_250);
and U8133 (N_8133,N_2107,N_3729);
nand U8134 (N_8134,N_1802,N_1645);
nand U8135 (N_8135,N_3883,N_1760);
or U8136 (N_8136,N_1849,N_156);
nor U8137 (N_8137,N_646,N_2430);
nor U8138 (N_8138,N_3130,N_1219);
nand U8139 (N_8139,N_4809,N_2970);
or U8140 (N_8140,N_1000,N_1119);
nand U8141 (N_8141,N_471,N_4992);
and U8142 (N_8142,N_536,N_2424);
or U8143 (N_8143,N_986,N_2799);
or U8144 (N_8144,N_4809,N_641);
and U8145 (N_8145,N_313,N_4970);
or U8146 (N_8146,N_1564,N_318);
or U8147 (N_8147,N_2884,N_1902);
nor U8148 (N_8148,N_850,N_973);
nand U8149 (N_8149,N_4975,N_3986);
or U8150 (N_8150,N_671,N_3642);
and U8151 (N_8151,N_4970,N_487);
and U8152 (N_8152,N_524,N_480);
nand U8153 (N_8153,N_1253,N_863);
nand U8154 (N_8154,N_747,N_3499);
nand U8155 (N_8155,N_3109,N_4127);
nor U8156 (N_8156,N_40,N_2351);
nor U8157 (N_8157,N_1637,N_1374);
nand U8158 (N_8158,N_4052,N_1332);
nor U8159 (N_8159,N_4174,N_118);
and U8160 (N_8160,N_815,N_752);
or U8161 (N_8161,N_3186,N_175);
or U8162 (N_8162,N_2968,N_4162);
nand U8163 (N_8163,N_1930,N_1065);
nand U8164 (N_8164,N_3107,N_2810);
or U8165 (N_8165,N_2627,N_164);
nor U8166 (N_8166,N_2820,N_2653);
nor U8167 (N_8167,N_87,N_2603);
nor U8168 (N_8168,N_3422,N_2366);
and U8169 (N_8169,N_1457,N_4007);
and U8170 (N_8170,N_184,N_4104);
and U8171 (N_8171,N_1857,N_3418);
nor U8172 (N_8172,N_778,N_2169);
nor U8173 (N_8173,N_831,N_1079);
and U8174 (N_8174,N_641,N_4104);
nor U8175 (N_8175,N_4628,N_1952);
nand U8176 (N_8176,N_3895,N_2868);
nor U8177 (N_8177,N_3717,N_1314);
and U8178 (N_8178,N_1833,N_82);
and U8179 (N_8179,N_3518,N_2555);
and U8180 (N_8180,N_3361,N_2677);
nand U8181 (N_8181,N_2020,N_1871);
and U8182 (N_8182,N_3174,N_4525);
nor U8183 (N_8183,N_175,N_4035);
or U8184 (N_8184,N_3700,N_1878);
and U8185 (N_8185,N_1203,N_1982);
or U8186 (N_8186,N_4492,N_1547);
nor U8187 (N_8187,N_154,N_3299);
nand U8188 (N_8188,N_53,N_1957);
and U8189 (N_8189,N_2425,N_173);
nand U8190 (N_8190,N_1980,N_3591);
and U8191 (N_8191,N_2717,N_4462);
or U8192 (N_8192,N_1422,N_3707);
nor U8193 (N_8193,N_778,N_1546);
nand U8194 (N_8194,N_2522,N_4441);
or U8195 (N_8195,N_252,N_1391);
nand U8196 (N_8196,N_3017,N_259);
and U8197 (N_8197,N_1167,N_1138);
nand U8198 (N_8198,N_803,N_4314);
or U8199 (N_8199,N_4324,N_2912);
nand U8200 (N_8200,N_4796,N_3550);
and U8201 (N_8201,N_605,N_1947);
and U8202 (N_8202,N_4516,N_4694);
nor U8203 (N_8203,N_4506,N_1887);
nor U8204 (N_8204,N_3247,N_1360);
nand U8205 (N_8205,N_3868,N_4567);
and U8206 (N_8206,N_307,N_4605);
nand U8207 (N_8207,N_2706,N_3966);
nand U8208 (N_8208,N_58,N_1659);
or U8209 (N_8209,N_3491,N_1250);
or U8210 (N_8210,N_3201,N_0);
or U8211 (N_8211,N_968,N_4679);
nor U8212 (N_8212,N_149,N_4579);
or U8213 (N_8213,N_1118,N_2403);
or U8214 (N_8214,N_4402,N_3544);
and U8215 (N_8215,N_4306,N_1136);
and U8216 (N_8216,N_1381,N_4987);
nor U8217 (N_8217,N_3787,N_2928);
or U8218 (N_8218,N_2720,N_3928);
and U8219 (N_8219,N_2857,N_1653);
and U8220 (N_8220,N_4280,N_715);
and U8221 (N_8221,N_1631,N_1739);
and U8222 (N_8222,N_1411,N_3078);
and U8223 (N_8223,N_2238,N_2538);
or U8224 (N_8224,N_4817,N_4363);
nor U8225 (N_8225,N_4924,N_2816);
or U8226 (N_8226,N_157,N_4574);
nor U8227 (N_8227,N_4236,N_2535);
or U8228 (N_8228,N_2550,N_2078);
or U8229 (N_8229,N_2757,N_994);
nand U8230 (N_8230,N_842,N_3105);
and U8231 (N_8231,N_693,N_3195);
nand U8232 (N_8232,N_2881,N_4386);
nand U8233 (N_8233,N_2899,N_496);
or U8234 (N_8234,N_3447,N_2633);
or U8235 (N_8235,N_4420,N_3453);
and U8236 (N_8236,N_2030,N_3038);
and U8237 (N_8237,N_4907,N_1224);
and U8238 (N_8238,N_2336,N_734);
nor U8239 (N_8239,N_1260,N_4351);
or U8240 (N_8240,N_4828,N_3993);
nor U8241 (N_8241,N_3805,N_4165);
or U8242 (N_8242,N_3495,N_1796);
or U8243 (N_8243,N_2451,N_294);
nand U8244 (N_8244,N_4498,N_140);
nor U8245 (N_8245,N_3506,N_4490);
nor U8246 (N_8246,N_1188,N_3800);
nand U8247 (N_8247,N_3408,N_1773);
nor U8248 (N_8248,N_4410,N_1741);
nand U8249 (N_8249,N_3811,N_2623);
or U8250 (N_8250,N_2896,N_4563);
nor U8251 (N_8251,N_2713,N_127);
and U8252 (N_8252,N_2411,N_1068);
nor U8253 (N_8253,N_1529,N_1110);
nand U8254 (N_8254,N_3798,N_2703);
or U8255 (N_8255,N_2565,N_1216);
nor U8256 (N_8256,N_2790,N_1708);
and U8257 (N_8257,N_344,N_4632);
xnor U8258 (N_8258,N_1146,N_2756);
or U8259 (N_8259,N_4507,N_2731);
or U8260 (N_8260,N_3394,N_3795);
nor U8261 (N_8261,N_4772,N_1537);
nand U8262 (N_8262,N_1969,N_1266);
nand U8263 (N_8263,N_3544,N_696);
nand U8264 (N_8264,N_4710,N_4232);
and U8265 (N_8265,N_1629,N_2501);
nor U8266 (N_8266,N_1757,N_246);
and U8267 (N_8267,N_3056,N_3851);
nor U8268 (N_8268,N_4358,N_771);
nand U8269 (N_8269,N_967,N_1881);
nand U8270 (N_8270,N_2855,N_3529);
nor U8271 (N_8271,N_2713,N_160);
and U8272 (N_8272,N_319,N_1503);
nand U8273 (N_8273,N_1508,N_4318);
nor U8274 (N_8274,N_4214,N_1007);
or U8275 (N_8275,N_2204,N_2979);
and U8276 (N_8276,N_3756,N_4870);
nor U8277 (N_8277,N_2197,N_4024);
and U8278 (N_8278,N_3294,N_3332);
nand U8279 (N_8279,N_3449,N_3727);
or U8280 (N_8280,N_763,N_706);
nand U8281 (N_8281,N_4229,N_3949);
and U8282 (N_8282,N_2685,N_2969);
or U8283 (N_8283,N_2945,N_3926);
nand U8284 (N_8284,N_2043,N_1040);
or U8285 (N_8285,N_638,N_326);
nor U8286 (N_8286,N_273,N_3687);
nor U8287 (N_8287,N_2139,N_3991);
or U8288 (N_8288,N_1133,N_2553);
nand U8289 (N_8289,N_2774,N_2748);
or U8290 (N_8290,N_3032,N_2265);
or U8291 (N_8291,N_2971,N_3842);
and U8292 (N_8292,N_177,N_791);
nand U8293 (N_8293,N_2025,N_3972);
and U8294 (N_8294,N_3456,N_2439);
nor U8295 (N_8295,N_3082,N_2739);
nor U8296 (N_8296,N_2684,N_4586);
nor U8297 (N_8297,N_2212,N_1884);
and U8298 (N_8298,N_2420,N_3324);
nand U8299 (N_8299,N_3132,N_3303);
or U8300 (N_8300,N_4874,N_3592);
and U8301 (N_8301,N_724,N_2101);
or U8302 (N_8302,N_3540,N_101);
nor U8303 (N_8303,N_3704,N_412);
and U8304 (N_8304,N_3842,N_3951);
or U8305 (N_8305,N_3983,N_4141);
nand U8306 (N_8306,N_2527,N_2639);
nor U8307 (N_8307,N_1026,N_2720);
or U8308 (N_8308,N_2940,N_341);
nand U8309 (N_8309,N_2715,N_4345);
and U8310 (N_8310,N_662,N_2370);
nand U8311 (N_8311,N_1475,N_4466);
or U8312 (N_8312,N_2074,N_1218);
or U8313 (N_8313,N_2811,N_1671);
and U8314 (N_8314,N_2623,N_4722);
nand U8315 (N_8315,N_1743,N_1911);
nor U8316 (N_8316,N_3316,N_1070);
nor U8317 (N_8317,N_1332,N_4323);
nor U8318 (N_8318,N_3085,N_3059);
and U8319 (N_8319,N_4595,N_896);
nor U8320 (N_8320,N_3905,N_4078);
nor U8321 (N_8321,N_3425,N_3302);
nor U8322 (N_8322,N_3733,N_2346);
or U8323 (N_8323,N_4911,N_2383);
or U8324 (N_8324,N_1337,N_3238);
nor U8325 (N_8325,N_4893,N_4813);
nor U8326 (N_8326,N_851,N_4292);
nand U8327 (N_8327,N_822,N_2318);
nand U8328 (N_8328,N_3257,N_1798);
nand U8329 (N_8329,N_4465,N_3832);
nand U8330 (N_8330,N_4612,N_3388);
or U8331 (N_8331,N_984,N_2816);
nor U8332 (N_8332,N_2938,N_2904);
nand U8333 (N_8333,N_3251,N_2036);
or U8334 (N_8334,N_4253,N_3443);
or U8335 (N_8335,N_2832,N_1218);
nor U8336 (N_8336,N_1229,N_1668);
nand U8337 (N_8337,N_2512,N_4164);
nor U8338 (N_8338,N_133,N_3125);
or U8339 (N_8339,N_1484,N_3400);
nor U8340 (N_8340,N_3467,N_1813);
nand U8341 (N_8341,N_552,N_2408);
nand U8342 (N_8342,N_638,N_3483);
nor U8343 (N_8343,N_4633,N_2465);
and U8344 (N_8344,N_1522,N_4747);
or U8345 (N_8345,N_2618,N_4398);
nor U8346 (N_8346,N_3029,N_3487);
or U8347 (N_8347,N_1406,N_1656);
or U8348 (N_8348,N_1409,N_1690);
or U8349 (N_8349,N_26,N_4691);
and U8350 (N_8350,N_301,N_3422);
or U8351 (N_8351,N_489,N_4238);
nand U8352 (N_8352,N_1566,N_1334);
and U8353 (N_8353,N_650,N_4752);
nor U8354 (N_8354,N_1055,N_421);
and U8355 (N_8355,N_1941,N_2180);
nor U8356 (N_8356,N_4629,N_3565);
nor U8357 (N_8357,N_1026,N_868);
nor U8358 (N_8358,N_3614,N_3353);
nand U8359 (N_8359,N_2268,N_154);
nor U8360 (N_8360,N_2454,N_2923);
or U8361 (N_8361,N_4113,N_770);
or U8362 (N_8362,N_1613,N_4550);
and U8363 (N_8363,N_4726,N_3135);
or U8364 (N_8364,N_4165,N_3496);
nor U8365 (N_8365,N_762,N_2558);
or U8366 (N_8366,N_3392,N_4190);
and U8367 (N_8367,N_4625,N_2730);
and U8368 (N_8368,N_4722,N_4320);
nor U8369 (N_8369,N_3016,N_54);
and U8370 (N_8370,N_3598,N_1999);
nor U8371 (N_8371,N_2331,N_3299);
nor U8372 (N_8372,N_3852,N_4401);
and U8373 (N_8373,N_258,N_3964);
nor U8374 (N_8374,N_140,N_562);
and U8375 (N_8375,N_2292,N_650);
nand U8376 (N_8376,N_3053,N_4136);
nand U8377 (N_8377,N_4673,N_1843);
nor U8378 (N_8378,N_1130,N_3342);
or U8379 (N_8379,N_1032,N_4428);
or U8380 (N_8380,N_1710,N_1134);
nand U8381 (N_8381,N_1262,N_3398);
or U8382 (N_8382,N_1387,N_3896);
and U8383 (N_8383,N_2510,N_2222);
and U8384 (N_8384,N_4119,N_1030);
nor U8385 (N_8385,N_3145,N_2873);
and U8386 (N_8386,N_3166,N_3652);
nor U8387 (N_8387,N_4172,N_4954);
nand U8388 (N_8388,N_284,N_3407);
or U8389 (N_8389,N_3561,N_702);
nor U8390 (N_8390,N_222,N_3190);
nor U8391 (N_8391,N_1099,N_2002);
and U8392 (N_8392,N_2809,N_3419);
xnor U8393 (N_8393,N_3790,N_1049);
and U8394 (N_8394,N_1673,N_3821);
nand U8395 (N_8395,N_4778,N_1666);
and U8396 (N_8396,N_563,N_1791);
or U8397 (N_8397,N_601,N_3874);
nand U8398 (N_8398,N_4255,N_154);
and U8399 (N_8399,N_4286,N_2524);
nand U8400 (N_8400,N_4955,N_1221);
nor U8401 (N_8401,N_4846,N_3683);
nand U8402 (N_8402,N_1031,N_4401);
nand U8403 (N_8403,N_455,N_2441);
nand U8404 (N_8404,N_2944,N_3693);
nor U8405 (N_8405,N_2085,N_536);
nand U8406 (N_8406,N_4342,N_1298);
nor U8407 (N_8407,N_1203,N_3594);
or U8408 (N_8408,N_2086,N_2145);
nor U8409 (N_8409,N_3360,N_1414);
or U8410 (N_8410,N_3436,N_1079);
nor U8411 (N_8411,N_3178,N_4934);
nor U8412 (N_8412,N_2916,N_2472);
and U8413 (N_8413,N_2821,N_1738);
and U8414 (N_8414,N_4509,N_1786);
or U8415 (N_8415,N_1044,N_4937);
and U8416 (N_8416,N_4880,N_3957);
nor U8417 (N_8417,N_2178,N_4571);
nand U8418 (N_8418,N_1594,N_2375);
nor U8419 (N_8419,N_4320,N_3195);
nor U8420 (N_8420,N_2003,N_3848);
or U8421 (N_8421,N_2702,N_3973);
and U8422 (N_8422,N_3333,N_4205);
nor U8423 (N_8423,N_3218,N_4612);
or U8424 (N_8424,N_3042,N_4632);
nand U8425 (N_8425,N_1855,N_4430);
and U8426 (N_8426,N_4081,N_2051);
nand U8427 (N_8427,N_4656,N_4662);
or U8428 (N_8428,N_1404,N_1174);
or U8429 (N_8429,N_4047,N_4073);
or U8430 (N_8430,N_4991,N_2393);
nand U8431 (N_8431,N_3895,N_4988);
or U8432 (N_8432,N_1976,N_1137);
or U8433 (N_8433,N_3037,N_3654);
nand U8434 (N_8434,N_2945,N_1257);
or U8435 (N_8435,N_2218,N_4251);
and U8436 (N_8436,N_1718,N_3837);
nand U8437 (N_8437,N_784,N_1321);
nand U8438 (N_8438,N_2742,N_4877);
or U8439 (N_8439,N_2502,N_2393);
and U8440 (N_8440,N_4940,N_4164);
nand U8441 (N_8441,N_3775,N_3389);
nor U8442 (N_8442,N_4030,N_1840);
nand U8443 (N_8443,N_4104,N_3177);
nand U8444 (N_8444,N_3626,N_1514);
nand U8445 (N_8445,N_544,N_2054);
and U8446 (N_8446,N_1414,N_3463);
and U8447 (N_8447,N_1261,N_4401);
nor U8448 (N_8448,N_1738,N_4756);
nand U8449 (N_8449,N_949,N_3108);
and U8450 (N_8450,N_3298,N_1910);
or U8451 (N_8451,N_481,N_4195);
nor U8452 (N_8452,N_468,N_4272);
nand U8453 (N_8453,N_2144,N_2312);
and U8454 (N_8454,N_2396,N_3689);
and U8455 (N_8455,N_2397,N_70);
nand U8456 (N_8456,N_836,N_1776);
nor U8457 (N_8457,N_2197,N_1462);
nor U8458 (N_8458,N_3409,N_3313);
nand U8459 (N_8459,N_1604,N_4102);
or U8460 (N_8460,N_4823,N_616);
and U8461 (N_8461,N_4074,N_3622);
and U8462 (N_8462,N_2511,N_3086);
nor U8463 (N_8463,N_3249,N_549);
nor U8464 (N_8464,N_1149,N_914);
nand U8465 (N_8465,N_4700,N_820);
and U8466 (N_8466,N_251,N_1951);
nand U8467 (N_8467,N_3426,N_120);
and U8468 (N_8468,N_2286,N_1870);
and U8469 (N_8469,N_2234,N_4936);
nand U8470 (N_8470,N_4426,N_1861);
nor U8471 (N_8471,N_4234,N_899);
and U8472 (N_8472,N_3729,N_1048);
or U8473 (N_8473,N_4954,N_2983);
nand U8474 (N_8474,N_392,N_995);
nand U8475 (N_8475,N_2801,N_928);
nor U8476 (N_8476,N_2482,N_3218);
or U8477 (N_8477,N_1878,N_4161);
and U8478 (N_8478,N_4457,N_342);
nor U8479 (N_8479,N_4149,N_22);
xor U8480 (N_8480,N_4733,N_177);
nor U8481 (N_8481,N_1153,N_3539);
and U8482 (N_8482,N_2516,N_3618);
nor U8483 (N_8483,N_1538,N_3409);
or U8484 (N_8484,N_2130,N_2394);
xor U8485 (N_8485,N_4536,N_427);
nor U8486 (N_8486,N_4117,N_2150);
or U8487 (N_8487,N_1651,N_2347);
nand U8488 (N_8488,N_3672,N_4228);
or U8489 (N_8489,N_3834,N_4667);
and U8490 (N_8490,N_3967,N_2638);
nor U8491 (N_8491,N_2013,N_3942);
nand U8492 (N_8492,N_1827,N_3508);
nor U8493 (N_8493,N_3665,N_1234);
nor U8494 (N_8494,N_322,N_2734);
or U8495 (N_8495,N_78,N_2631);
or U8496 (N_8496,N_3463,N_4086);
nand U8497 (N_8497,N_1749,N_1410);
or U8498 (N_8498,N_4228,N_2197);
or U8499 (N_8499,N_380,N_1156);
or U8500 (N_8500,N_1125,N_1723);
or U8501 (N_8501,N_3856,N_3741);
or U8502 (N_8502,N_2118,N_1854);
nand U8503 (N_8503,N_3929,N_1699);
and U8504 (N_8504,N_3360,N_452);
or U8505 (N_8505,N_2415,N_4503);
nor U8506 (N_8506,N_1745,N_1968);
or U8507 (N_8507,N_1953,N_3987);
and U8508 (N_8508,N_2651,N_1528);
and U8509 (N_8509,N_4774,N_3158);
nor U8510 (N_8510,N_2721,N_126);
nor U8511 (N_8511,N_3136,N_1714);
and U8512 (N_8512,N_2840,N_3955);
nand U8513 (N_8513,N_4339,N_245);
nor U8514 (N_8514,N_307,N_107);
or U8515 (N_8515,N_1332,N_4894);
nor U8516 (N_8516,N_4077,N_2813);
or U8517 (N_8517,N_4236,N_4408);
nand U8518 (N_8518,N_231,N_4244);
nor U8519 (N_8519,N_1748,N_585);
and U8520 (N_8520,N_3096,N_1499);
nand U8521 (N_8521,N_1983,N_2623);
and U8522 (N_8522,N_2288,N_4082);
nor U8523 (N_8523,N_4417,N_2976);
nand U8524 (N_8524,N_339,N_1268);
nand U8525 (N_8525,N_578,N_2018);
and U8526 (N_8526,N_1446,N_4092);
or U8527 (N_8527,N_2415,N_3895);
and U8528 (N_8528,N_2117,N_2585);
or U8529 (N_8529,N_22,N_2976);
nand U8530 (N_8530,N_3179,N_687);
nand U8531 (N_8531,N_652,N_2195);
nand U8532 (N_8532,N_4510,N_3066);
and U8533 (N_8533,N_3964,N_2563);
and U8534 (N_8534,N_895,N_4187);
nand U8535 (N_8535,N_1042,N_263);
and U8536 (N_8536,N_2659,N_2922);
nand U8537 (N_8537,N_2971,N_1706);
nor U8538 (N_8538,N_230,N_18);
nand U8539 (N_8539,N_329,N_2493);
and U8540 (N_8540,N_3116,N_72);
nand U8541 (N_8541,N_4534,N_3861);
nand U8542 (N_8542,N_1763,N_1765);
and U8543 (N_8543,N_4228,N_4307);
nand U8544 (N_8544,N_4602,N_2652);
nor U8545 (N_8545,N_4694,N_4687);
nand U8546 (N_8546,N_4493,N_4083);
and U8547 (N_8547,N_1270,N_3357);
xnor U8548 (N_8548,N_3488,N_4360);
nor U8549 (N_8549,N_1744,N_4973);
nor U8550 (N_8550,N_2950,N_2377);
nand U8551 (N_8551,N_1229,N_380);
nor U8552 (N_8552,N_495,N_3289);
and U8553 (N_8553,N_1036,N_4531);
and U8554 (N_8554,N_48,N_3948);
nand U8555 (N_8555,N_2771,N_144);
nor U8556 (N_8556,N_3410,N_591);
nor U8557 (N_8557,N_3268,N_4374);
nand U8558 (N_8558,N_1300,N_2457);
nor U8559 (N_8559,N_1445,N_1443);
and U8560 (N_8560,N_1796,N_3594);
and U8561 (N_8561,N_848,N_1166);
nand U8562 (N_8562,N_2849,N_3248);
and U8563 (N_8563,N_4254,N_1994);
nand U8564 (N_8564,N_1277,N_3010);
nand U8565 (N_8565,N_892,N_247);
and U8566 (N_8566,N_1458,N_1401);
and U8567 (N_8567,N_2709,N_1845);
nand U8568 (N_8568,N_2990,N_3786);
and U8569 (N_8569,N_4464,N_1049);
or U8570 (N_8570,N_2548,N_1993);
nor U8571 (N_8571,N_2889,N_2435);
and U8572 (N_8572,N_2441,N_2358);
and U8573 (N_8573,N_2893,N_4451);
nor U8574 (N_8574,N_3699,N_4702);
or U8575 (N_8575,N_2995,N_1716);
nor U8576 (N_8576,N_4040,N_4487);
nand U8577 (N_8577,N_4614,N_2646);
xnor U8578 (N_8578,N_1723,N_623);
or U8579 (N_8579,N_3545,N_4848);
or U8580 (N_8580,N_4046,N_4395);
nand U8581 (N_8581,N_4573,N_189);
and U8582 (N_8582,N_294,N_2164);
nand U8583 (N_8583,N_1494,N_3378);
and U8584 (N_8584,N_4865,N_2560);
and U8585 (N_8585,N_1307,N_2100);
nor U8586 (N_8586,N_1418,N_939);
or U8587 (N_8587,N_932,N_3518);
nand U8588 (N_8588,N_2663,N_2759);
and U8589 (N_8589,N_4160,N_218);
and U8590 (N_8590,N_4151,N_3168);
or U8591 (N_8591,N_1285,N_3263);
nor U8592 (N_8592,N_4798,N_777);
and U8593 (N_8593,N_4952,N_4123);
nand U8594 (N_8594,N_74,N_3531);
and U8595 (N_8595,N_2376,N_504);
nand U8596 (N_8596,N_1402,N_3154);
and U8597 (N_8597,N_345,N_404);
or U8598 (N_8598,N_172,N_1704);
or U8599 (N_8599,N_3596,N_1991);
and U8600 (N_8600,N_4669,N_2010);
and U8601 (N_8601,N_3075,N_2366);
and U8602 (N_8602,N_1694,N_4085);
nand U8603 (N_8603,N_3490,N_4328);
or U8604 (N_8604,N_3187,N_1151);
and U8605 (N_8605,N_3367,N_3748);
and U8606 (N_8606,N_4158,N_1669);
nand U8607 (N_8607,N_3062,N_1150);
and U8608 (N_8608,N_3516,N_1703);
and U8609 (N_8609,N_3339,N_1404);
nor U8610 (N_8610,N_2635,N_4195);
or U8611 (N_8611,N_1659,N_4158);
xnor U8612 (N_8612,N_4389,N_1122);
nor U8613 (N_8613,N_666,N_2961);
nand U8614 (N_8614,N_3695,N_2821);
nor U8615 (N_8615,N_2626,N_2484);
or U8616 (N_8616,N_2621,N_3164);
and U8617 (N_8617,N_2522,N_949);
and U8618 (N_8618,N_1209,N_1184);
or U8619 (N_8619,N_1266,N_2601);
nand U8620 (N_8620,N_2583,N_2262);
or U8621 (N_8621,N_3092,N_973);
and U8622 (N_8622,N_3842,N_3337);
or U8623 (N_8623,N_3033,N_664);
nand U8624 (N_8624,N_715,N_4243);
nand U8625 (N_8625,N_3967,N_681);
nor U8626 (N_8626,N_2477,N_4088);
and U8627 (N_8627,N_3756,N_156);
nor U8628 (N_8628,N_1593,N_787);
and U8629 (N_8629,N_1151,N_593);
and U8630 (N_8630,N_1039,N_4594);
and U8631 (N_8631,N_2071,N_1736);
nor U8632 (N_8632,N_4253,N_2486);
or U8633 (N_8633,N_4658,N_3607);
or U8634 (N_8634,N_4574,N_788);
nand U8635 (N_8635,N_4601,N_466);
nor U8636 (N_8636,N_2810,N_663);
or U8637 (N_8637,N_4236,N_4343);
and U8638 (N_8638,N_1217,N_1520);
or U8639 (N_8639,N_2751,N_1083);
nor U8640 (N_8640,N_3812,N_66);
nand U8641 (N_8641,N_3961,N_2630);
and U8642 (N_8642,N_677,N_2564);
and U8643 (N_8643,N_549,N_1606);
or U8644 (N_8644,N_4893,N_1493);
nor U8645 (N_8645,N_1177,N_308);
nand U8646 (N_8646,N_487,N_3163);
nand U8647 (N_8647,N_1649,N_2932);
or U8648 (N_8648,N_3094,N_369);
and U8649 (N_8649,N_4901,N_3478);
nor U8650 (N_8650,N_1745,N_2184);
nor U8651 (N_8651,N_1005,N_48);
or U8652 (N_8652,N_3855,N_2929);
nor U8653 (N_8653,N_4707,N_4805);
nand U8654 (N_8654,N_2896,N_3964);
nand U8655 (N_8655,N_1016,N_1863);
or U8656 (N_8656,N_2461,N_4839);
nor U8657 (N_8657,N_762,N_2703);
or U8658 (N_8658,N_3326,N_3994);
nor U8659 (N_8659,N_1274,N_3653);
nor U8660 (N_8660,N_3006,N_661);
nand U8661 (N_8661,N_2057,N_1224);
or U8662 (N_8662,N_439,N_167);
nor U8663 (N_8663,N_3331,N_3832);
or U8664 (N_8664,N_3298,N_2856);
and U8665 (N_8665,N_4159,N_3032);
or U8666 (N_8666,N_1690,N_4356);
and U8667 (N_8667,N_1347,N_1222);
nor U8668 (N_8668,N_315,N_1840);
nor U8669 (N_8669,N_4440,N_2982);
or U8670 (N_8670,N_2530,N_1539);
or U8671 (N_8671,N_1070,N_2003);
nor U8672 (N_8672,N_4795,N_4014);
or U8673 (N_8673,N_36,N_1440);
and U8674 (N_8674,N_3681,N_3297);
nor U8675 (N_8675,N_1651,N_781);
nand U8676 (N_8676,N_4029,N_331);
and U8677 (N_8677,N_3521,N_1012);
nand U8678 (N_8678,N_4600,N_3726);
nor U8679 (N_8679,N_1741,N_3258);
nor U8680 (N_8680,N_1453,N_658);
and U8681 (N_8681,N_3217,N_4543);
or U8682 (N_8682,N_3920,N_2376);
or U8683 (N_8683,N_4089,N_2690);
or U8684 (N_8684,N_4763,N_2965);
nor U8685 (N_8685,N_4782,N_4950);
nor U8686 (N_8686,N_2017,N_2135);
nand U8687 (N_8687,N_4063,N_3494);
or U8688 (N_8688,N_2038,N_2314);
or U8689 (N_8689,N_4484,N_3025);
nand U8690 (N_8690,N_2025,N_747);
and U8691 (N_8691,N_2599,N_4948);
or U8692 (N_8692,N_4192,N_1519);
nand U8693 (N_8693,N_116,N_563);
nor U8694 (N_8694,N_1506,N_1656);
or U8695 (N_8695,N_2217,N_3878);
nand U8696 (N_8696,N_914,N_3732);
or U8697 (N_8697,N_942,N_3390);
nand U8698 (N_8698,N_684,N_3107);
nand U8699 (N_8699,N_2477,N_2315);
nor U8700 (N_8700,N_3706,N_4313);
or U8701 (N_8701,N_1280,N_3314);
nor U8702 (N_8702,N_4049,N_3168);
nor U8703 (N_8703,N_2702,N_486);
nor U8704 (N_8704,N_2938,N_3539);
nor U8705 (N_8705,N_1411,N_1333);
or U8706 (N_8706,N_4184,N_4322);
nor U8707 (N_8707,N_2572,N_2799);
nor U8708 (N_8708,N_4158,N_3483);
nor U8709 (N_8709,N_2878,N_1973);
and U8710 (N_8710,N_459,N_3832);
or U8711 (N_8711,N_4164,N_1067);
nand U8712 (N_8712,N_2099,N_4340);
nand U8713 (N_8713,N_415,N_3538);
and U8714 (N_8714,N_4837,N_3596);
or U8715 (N_8715,N_4928,N_3081);
and U8716 (N_8716,N_4483,N_245);
and U8717 (N_8717,N_1416,N_4527);
and U8718 (N_8718,N_4177,N_2892);
or U8719 (N_8719,N_150,N_2912);
or U8720 (N_8720,N_5,N_3517);
nor U8721 (N_8721,N_1559,N_113);
nand U8722 (N_8722,N_842,N_4707);
and U8723 (N_8723,N_2039,N_4446);
and U8724 (N_8724,N_4552,N_1820);
nor U8725 (N_8725,N_4226,N_1831);
or U8726 (N_8726,N_1357,N_141);
or U8727 (N_8727,N_4937,N_2803);
xnor U8728 (N_8728,N_450,N_2240);
xor U8729 (N_8729,N_267,N_4098);
nand U8730 (N_8730,N_3853,N_4204);
nand U8731 (N_8731,N_133,N_3942);
and U8732 (N_8732,N_576,N_1044);
nand U8733 (N_8733,N_4867,N_4848);
or U8734 (N_8734,N_76,N_1866);
nand U8735 (N_8735,N_4975,N_1587);
nand U8736 (N_8736,N_550,N_3331);
and U8737 (N_8737,N_1170,N_3300);
and U8738 (N_8738,N_4632,N_3262);
nand U8739 (N_8739,N_4772,N_4741);
or U8740 (N_8740,N_2779,N_1948);
nor U8741 (N_8741,N_1265,N_1117);
xnor U8742 (N_8742,N_3700,N_3453);
and U8743 (N_8743,N_1126,N_4720);
nand U8744 (N_8744,N_1960,N_4265);
nor U8745 (N_8745,N_3875,N_3739);
or U8746 (N_8746,N_1092,N_4724);
or U8747 (N_8747,N_3518,N_2914);
nor U8748 (N_8748,N_695,N_4835);
and U8749 (N_8749,N_686,N_440);
nand U8750 (N_8750,N_1939,N_1204);
and U8751 (N_8751,N_4097,N_208);
and U8752 (N_8752,N_2603,N_4330);
nand U8753 (N_8753,N_3949,N_4426);
or U8754 (N_8754,N_2486,N_3892);
or U8755 (N_8755,N_3443,N_2976);
or U8756 (N_8756,N_2884,N_1813);
nand U8757 (N_8757,N_985,N_811);
and U8758 (N_8758,N_305,N_3758);
nor U8759 (N_8759,N_4979,N_686);
or U8760 (N_8760,N_3383,N_1066);
or U8761 (N_8761,N_1547,N_2270);
nor U8762 (N_8762,N_151,N_4669);
nand U8763 (N_8763,N_3477,N_1299);
nor U8764 (N_8764,N_3031,N_43);
or U8765 (N_8765,N_2834,N_4838);
nor U8766 (N_8766,N_1316,N_994);
and U8767 (N_8767,N_844,N_57);
nor U8768 (N_8768,N_3207,N_3147);
nand U8769 (N_8769,N_242,N_3548);
or U8770 (N_8770,N_82,N_438);
nand U8771 (N_8771,N_333,N_1309);
and U8772 (N_8772,N_2937,N_2390);
nand U8773 (N_8773,N_1565,N_837);
and U8774 (N_8774,N_281,N_3382);
or U8775 (N_8775,N_566,N_2064);
and U8776 (N_8776,N_3961,N_4757);
nand U8777 (N_8777,N_2588,N_2064);
nand U8778 (N_8778,N_3183,N_2577);
nor U8779 (N_8779,N_2970,N_1172);
or U8780 (N_8780,N_1927,N_159);
and U8781 (N_8781,N_1255,N_3635);
nor U8782 (N_8782,N_3979,N_2022);
nand U8783 (N_8783,N_3310,N_4105);
and U8784 (N_8784,N_835,N_1508);
and U8785 (N_8785,N_3927,N_4001);
nand U8786 (N_8786,N_4877,N_4611);
nand U8787 (N_8787,N_3111,N_2379);
and U8788 (N_8788,N_2087,N_4275);
and U8789 (N_8789,N_2835,N_4016);
nand U8790 (N_8790,N_2205,N_403);
nand U8791 (N_8791,N_185,N_4742);
xor U8792 (N_8792,N_83,N_3490);
or U8793 (N_8793,N_684,N_786);
or U8794 (N_8794,N_985,N_1905);
and U8795 (N_8795,N_3402,N_4322);
and U8796 (N_8796,N_1839,N_704);
and U8797 (N_8797,N_2512,N_3316);
or U8798 (N_8798,N_2584,N_4566);
nand U8799 (N_8799,N_2608,N_4671);
or U8800 (N_8800,N_1019,N_3501);
and U8801 (N_8801,N_2213,N_4213);
or U8802 (N_8802,N_455,N_1838);
nand U8803 (N_8803,N_752,N_667);
nand U8804 (N_8804,N_3660,N_4586);
and U8805 (N_8805,N_1437,N_2401);
and U8806 (N_8806,N_4474,N_2435);
nand U8807 (N_8807,N_3793,N_193);
or U8808 (N_8808,N_4842,N_1458);
nand U8809 (N_8809,N_3867,N_4907);
and U8810 (N_8810,N_974,N_4694);
nor U8811 (N_8811,N_400,N_1139);
nor U8812 (N_8812,N_494,N_1369);
and U8813 (N_8813,N_4695,N_178);
nor U8814 (N_8814,N_4126,N_2132);
and U8815 (N_8815,N_1100,N_4222);
and U8816 (N_8816,N_4357,N_977);
nand U8817 (N_8817,N_4082,N_2397);
and U8818 (N_8818,N_1743,N_471);
nand U8819 (N_8819,N_175,N_3240);
or U8820 (N_8820,N_617,N_2899);
or U8821 (N_8821,N_3940,N_775);
or U8822 (N_8822,N_4409,N_1974);
and U8823 (N_8823,N_622,N_3944);
or U8824 (N_8824,N_3427,N_4000);
or U8825 (N_8825,N_4882,N_1277);
nand U8826 (N_8826,N_1913,N_1165);
nor U8827 (N_8827,N_47,N_4225);
and U8828 (N_8828,N_3707,N_3622);
or U8829 (N_8829,N_1634,N_233);
nor U8830 (N_8830,N_2687,N_894);
nand U8831 (N_8831,N_2774,N_4069);
or U8832 (N_8832,N_3166,N_3375);
nand U8833 (N_8833,N_2088,N_1177);
and U8834 (N_8834,N_4868,N_4899);
nor U8835 (N_8835,N_2632,N_1296);
and U8836 (N_8836,N_2316,N_2441);
and U8837 (N_8837,N_2796,N_4544);
nor U8838 (N_8838,N_2115,N_2263);
and U8839 (N_8839,N_3107,N_1766);
or U8840 (N_8840,N_4706,N_3138);
and U8841 (N_8841,N_68,N_3904);
nor U8842 (N_8842,N_4535,N_1852);
nor U8843 (N_8843,N_4691,N_4022);
nand U8844 (N_8844,N_356,N_827);
and U8845 (N_8845,N_4182,N_3550);
nor U8846 (N_8846,N_2493,N_1937);
or U8847 (N_8847,N_1464,N_1040);
nand U8848 (N_8848,N_1353,N_3462);
nand U8849 (N_8849,N_2992,N_4935);
nor U8850 (N_8850,N_862,N_4724);
or U8851 (N_8851,N_1615,N_2861);
and U8852 (N_8852,N_3285,N_3469);
or U8853 (N_8853,N_418,N_4272);
nor U8854 (N_8854,N_2310,N_3214);
nand U8855 (N_8855,N_3254,N_1608);
nand U8856 (N_8856,N_4270,N_3121);
or U8857 (N_8857,N_3876,N_3901);
nand U8858 (N_8858,N_3101,N_620);
or U8859 (N_8859,N_69,N_1767);
and U8860 (N_8860,N_959,N_1997);
and U8861 (N_8861,N_3901,N_614);
nor U8862 (N_8862,N_1826,N_1912);
nor U8863 (N_8863,N_2652,N_4096);
and U8864 (N_8864,N_3850,N_3349);
nor U8865 (N_8865,N_4396,N_456);
nand U8866 (N_8866,N_4204,N_1022);
nand U8867 (N_8867,N_4768,N_2539);
nor U8868 (N_8868,N_103,N_531);
nand U8869 (N_8869,N_622,N_3720);
and U8870 (N_8870,N_1309,N_4612);
and U8871 (N_8871,N_4611,N_3819);
or U8872 (N_8872,N_3190,N_3918);
or U8873 (N_8873,N_2456,N_2285);
nand U8874 (N_8874,N_4872,N_270);
or U8875 (N_8875,N_3023,N_473);
and U8876 (N_8876,N_324,N_2893);
nor U8877 (N_8877,N_2492,N_71);
and U8878 (N_8878,N_908,N_1789);
nor U8879 (N_8879,N_1851,N_3844);
nor U8880 (N_8880,N_327,N_3043);
nor U8881 (N_8881,N_812,N_3391);
or U8882 (N_8882,N_4194,N_190);
nand U8883 (N_8883,N_4363,N_511);
or U8884 (N_8884,N_1907,N_3882);
and U8885 (N_8885,N_4927,N_135);
or U8886 (N_8886,N_510,N_1885);
nand U8887 (N_8887,N_2432,N_2438);
nand U8888 (N_8888,N_1059,N_4137);
or U8889 (N_8889,N_2479,N_2960);
nand U8890 (N_8890,N_4235,N_672);
nand U8891 (N_8891,N_4415,N_605);
or U8892 (N_8892,N_1848,N_822);
or U8893 (N_8893,N_2947,N_4394);
and U8894 (N_8894,N_1117,N_4792);
and U8895 (N_8895,N_1029,N_135);
and U8896 (N_8896,N_1516,N_1971);
nor U8897 (N_8897,N_3978,N_292);
or U8898 (N_8898,N_1114,N_134);
and U8899 (N_8899,N_4085,N_3282);
and U8900 (N_8900,N_4398,N_704);
nand U8901 (N_8901,N_941,N_1199);
nand U8902 (N_8902,N_1447,N_3194);
nand U8903 (N_8903,N_4899,N_2070);
nor U8904 (N_8904,N_897,N_3626);
nor U8905 (N_8905,N_3141,N_2058);
and U8906 (N_8906,N_2241,N_3624);
or U8907 (N_8907,N_3971,N_3307);
nor U8908 (N_8908,N_4496,N_4133);
and U8909 (N_8909,N_2873,N_4552);
and U8910 (N_8910,N_3122,N_2803);
nor U8911 (N_8911,N_3445,N_520);
and U8912 (N_8912,N_953,N_4160);
and U8913 (N_8913,N_4616,N_32);
or U8914 (N_8914,N_118,N_3046);
or U8915 (N_8915,N_3404,N_4556);
nand U8916 (N_8916,N_2484,N_325);
nand U8917 (N_8917,N_4853,N_3701);
nor U8918 (N_8918,N_929,N_3728);
and U8919 (N_8919,N_1255,N_297);
nand U8920 (N_8920,N_2404,N_324);
nor U8921 (N_8921,N_3757,N_1132);
nor U8922 (N_8922,N_1394,N_4455);
nor U8923 (N_8923,N_185,N_418);
or U8924 (N_8924,N_3754,N_4403);
or U8925 (N_8925,N_4847,N_2710);
and U8926 (N_8926,N_1152,N_359);
or U8927 (N_8927,N_2254,N_504);
nor U8928 (N_8928,N_2025,N_3873);
or U8929 (N_8929,N_1181,N_2618);
or U8930 (N_8930,N_1258,N_4625);
or U8931 (N_8931,N_3153,N_3382);
and U8932 (N_8932,N_747,N_1727);
or U8933 (N_8933,N_4210,N_3886);
nor U8934 (N_8934,N_335,N_3694);
and U8935 (N_8935,N_4253,N_2521);
xnor U8936 (N_8936,N_2101,N_4533);
or U8937 (N_8937,N_4902,N_2628);
nor U8938 (N_8938,N_862,N_2060);
and U8939 (N_8939,N_1204,N_1151);
or U8940 (N_8940,N_85,N_3907);
nand U8941 (N_8941,N_428,N_1221);
and U8942 (N_8942,N_24,N_2843);
or U8943 (N_8943,N_334,N_1216);
or U8944 (N_8944,N_4165,N_1499);
and U8945 (N_8945,N_2829,N_3467);
nand U8946 (N_8946,N_253,N_2181);
nand U8947 (N_8947,N_876,N_4801);
or U8948 (N_8948,N_2071,N_3596);
nor U8949 (N_8949,N_96,N_179);
and U8950 (N_8950,N_1931,N_4313);
nor U8951 (N_8951,N_1809,N_3986);
nand U8952 (N_8952,N_1812,N_256);
and U8953 (N_8953,N_4022,N_1504);
nand U8954 (N_8954,N_2919,N_3539);
nand U8955 (N_8955,N_93,N_1046);
and U8956 (N_8956,N_1570,N_1344);
and U8957 (N_8957,N_4490,N_1257);
nor U8958 (N_8958,N_177,N_4225);
nor U8959 (N_8959,N_2283,N_1635);
nor U8960 (N_8960,N_1846,N_3467);
and U8961 (N_8961,N_535,N_2761);
and U8962 (N_8962,N_1183,N_3521);
nand U8963 (N_8963,N_2163,N_3087);
or U8964 (N_8964,N_4995,N_247);
nand U8965 (N_8965,N_25,N_4425);
and U8966 (N_8966,N_3256,N_4848);
nand U8967 (N_8967,N_2456,N_3465);
and U8968 (N_8968,N_3766,N_69);
and U8969 (N_8969,N_2909,N_2338);
or U8970 (N_8970,N_2977,N_4696);
or U8971 (N_8971,N_3891,N_4256);
and U8972 (N_8972,N_4444,N_2059);
nor U8973 (N_8973,N_2522,N_128);
or U8974 (N_8974,N_2040,N_3320);
or U8975 (N_8975,N_1862,N_2495);
nor U8976 (N_8976,N_622,N_961);
and U8977 (N_8977,N_2449,N_1820);
and U8978 (N_8978,N_2066,N_3711);
and U8979 (N_8979,N_4487,N_3748);
nand U8980 (N_8980,N_2320,N_4143);
and U8981 (N_8981,N_134,N_4239);
and U8982 (N_8982,N_1969,N_944);
nor U8983 (N_8983,N_4931,N_1392);
or U8984 (N_8984,N_1406,N_615);
nor U8985 (N_8985,N_4056,N_3618);
nand U8986 (N_8986,N_348,N_4474);
and U8987 (N_8987,N_42,N_3261);
and U8988 (N_8988,N_1078,N_1578);
nor U8989 (N_8989,N_2565,N_3237);
nor U8990 (N_8990,N_462,N_3166);
or U8991 (N_8991,N_2733,N_457);
nor U8992 (N_8992,N_190,N_995);
nand U8993 (N_8993,N_1902,N_4262);
and U8994 (N_8994,N_2972,N_3963);
nor U8995 (N_8995,N_4338,N_524);
and U8996 (N_8996,N_4127,N_299);
or U8997 (N_8997,N_4480,N_3327);
xor U8998 (N_8998,N_1755,N_3848);
nand U8999 (N_8999,N_2992,N_2864);
or U9000 (N_9000,N_1649,N_2983);
or U9001 (N_9001,N_1574,N_4262);
and U9002 (N_9002,N_1772,N_2136);
nand U9003 (N_9003,N_4434,N_1158);
nor U9004 (N_9004,N_4812,N_4288);
and U9005 (N_9005,N_2263,N_2023);
nand U9006 (N_9006,N_4366,N_586);
nand U9007 (N_9007,N_3280,N_1386);
and U9008 (N_9008,N_4764,N_292);
and U9009 (N_9009,N_4148,N_1812);
nor U9010 (N_9010,N_2796,N_2056);
xor U9011 (N_9011,N_3153,N_1840);
nor U9012 (N_9012,N_3295,N_3125);
or U9013 (N_9013,N_4338,N_1748);
or U9014 (N_9014,N_2891,N_117);
or U9015 (N_9015,N_4653,N_2485);
nand U9016 (N_9016,N_2848,N_3068);
and U9017 (N_9017,N_4952,N_2043);
and U9018 (N_9018,N_4844,N_4321);
and U9019 (N_9019,N_2841,N_3444);
nor U9020 (N_9020,N_3059,N_1415);
nor U9021 (N_9021,N_3461,N_2567);
nand U9022 (N_9022,N_1190,N_143);
nor U9023 (N_9023,N_3359,N_169);
nand U9024 (N_9024,N_1171,N_2019);
nor U9025 (N_9025,N_3283,N_2218);
and U9026 (N_9026,N_2516,N_4536);
or U9027 (N_9027,N_2480,N_2713);
nor U9028 (N_9028,N_2367,N_747);
or U9029 (N_9029,N_4101,N_4375);
or U9030 (N_9030,N_4407,N_2634);
nand U9031 (N_9031,N_3519,N_4553);
xnor U9032 (N_9032,N_2334,N_2608);
nand U9033 (N_9033,N_2397,N_3030);
nor U9034 (N_9034,N_1764,N_3656);
nor U9035 (N_9035,N_4970,N_4996);
nand U9036 (N_9036,N_712,N_4504);
or U9037 (N_9037,N_4451,N_4631);
nor U9038 (N_9038,N_4726,N_4076);
nand U9039 (N_9039,N_1600,N_974);
or U9040 (N_9040,N_660,N_1764);
nor U9041 (N_9041,N_3356,N_2261);
and U9042 (N_9042,N_1053,N_846);
nand U9043 (N_9043,N_2498,N_2384);
and U9044 (N_9044,N_3362,N_4688);
and U9045 (N_9045,N_1122,N_3764);
or U9046 (N_9046,N_2321,N_1156);
or U9047 (N_9047,N_3864,N_1835);
and U9048 (N_9048,N_2525,N_4679);
nor U9049 (N_9049,N_4867,N_2524);
and U9050 (N_9050,N_3993,N_2584);
and U9051 (N_9051,N_519,N_1450);
nor U9052 (N_9052,N_3768,N_4883);
or U9053 (N_9053,N_2986,N_4343);
and U9054 (N_9054,N_3279,N_3006);
nor U9055 (N_9055,N_41,N_3516);
and U9056 (N_9056,N_4733,N_4528);
and U9057 (N_9057,N_4635,N_2461);
or U9058 (N_9058,N_4640,N_3808);
nor U9059 (N_9059,N_3249,N_476);
or U9060 (N_9060,N_1689,N_465);
nand U9061 (N_9061,N_3687,N_3007);
nor U9062 (N_9062,N_496,N_3199);
nand U9063 (N_9063,N_3793,N_4180);
and U9064 (N_9064,N_3138,N_2974);
nor U9065 (N_9065,N_923,N_2636);
nor U9066 (N_9066,N_1834,N_1228);
and U9067 (N_9067,N_3408,N_1975);
nor U9068 (N_9068,N_3410,N_2444);
and U9069 (N_9069,N_4214,N_866);
nand U9070 (N_9070,N_3118,N_4698);
or U9071 (N_9071,N_1153,N_2984);
or U9072 (N_9072,N_2479,N_1941);
nand U9073 (N_9073,N_4585,N_1681);
and U9074 (N_9074,N_70,N_1190);
nor U9075 (N_9075,N_3524,N_3983);
and U9076 (N_9076,N_2305,N_2711);
nor U9077 (N_9077,N_468,N_702);
xnor U9078 (N_9078,N_2505,N_2287);
nand U9079 (N_9079,N_2267,N_4913);
and U9080 (N_9080,N_3982,N_4226);
nand U9081 (N_9081,N_1946,N_1952);
nor U9082 (N_9082,N_1856,N_3517);
and U9083 (N_9083,N_3350,N_967);
or U9084 (N_9084,N_3619,N_1477);
or U9085 (N_9085,N_2530,N_4490);
and U9086 (N_9086,N_118,N_1376);
xor U9087 (N_9087,N_2206,N_4709);
nand U9088 (N_9088,N_1072,N_1360);
and U9089 (N_9089,N_4667,N_595);
nor U9090 (N_9090,N_2610,N_1708);
nand U9091 (N_9091,N_4568,N_2886);
and U9092 (N_9092,N_3798,N_172);
nand U9093 (N_9093,N_1299,N_443);
nor U9094 (N_9094,N_763,N_4501);
nand U9095 (N_9095,N_3476,N_1614);
nor U9096 (N_9096,N_2856,N_2436);
or U9097 (N_9097,N_4519,N_3843);
nor U9098 (N_9098,N_2496,N_1345);
nand U9099 (N_9099,N_1016,N_2467);
nor U9100 (N_9100,N_2506,N_4174);
xnor U9101 (N_9101,N_3564,N_4390);
nor U9102 (N_9102,N_3601,N_4981);
or U9103 (N_9103,N_3795,N_2734);
nand U9104 (N_9104,N_40,N_3300);
nor U9105 (N_9105,N_915,N_4638);
or U9106 (N_9106,N_4768,N_3118);
and U9107 (N_9107,N_3252,N_1781);
or U9108 (N_9108,N_590,N_2604);
and U9109 (N_9109,N_1366,N_663);
nor U9110 (N_9110,N_4117,N_1168);
or U9111 (N_9111,N_4715,N_2763);
or U9112 (N_9112,N_4530,N_3852);
nand U9113 (N_9113,N_4223,N_4659);
nand U9114 (N_9114,N_2097,N_4457);
or U9115 (N_9115,N_2725,N_3333);
nor U9116 (N_9116,N_4053,N_1970);
nand U9117 (N_9117,N_4766,N_3047);
nor U9118 (N_9118,N_2615,N_3452);
and U9119 (N_9119,N_2114,N_4026);
or U9120 (N_9120,N_4898,N_1706);
xnor U9121 (N_9121,N_4392,N_2650);
nand U9122 (N_9122,N_3529,N_1471);
nand U9123 (N_9123,N_4290,N_4095);
nand U9124 (N_9124,N_1102,N_3541);
or U9125 (N_9125,N_4305,N_3307);
nand U9126 (N_9126,N_993,N_3192);
and U9127 (N_9127,N_3245,N_2820);
or U9128 (N_9128,N_4984,N_626);
and U9129 (N_9129,N_4203,N_1860);
nand U9130 (N_9130,N_1831,N_4679);
nor U9131 (N_9131,N_4908,N_923);
or U9132 (N_9132,N_4346,N_2259);
and U9133 (N_9133,N_2782,N_807);
nor U9134 (N_9134,N_2269,N_4410);
nor U9135 (N_9135,N_4811,N_3507);
xor U9136 (N_9136,N_85,N_2187);
and U9137 (N_9137,N_3203,N_670);
nor U9138 (N_9138,N_1679,N_3465);
and U9139 (N_9139,N_3387,N_4675);
and U9140 (N_9140,N_4414,N_2629);
and U9141 (N_9141,N_2258,N_3297);
or U9142 (N_9142,N_4718,N_660);
or U9143 (N_9143,N_1936,N_2976);
or U9144 (N_9144,N_4548,N_3213);
nand U9145 (N_9145,N_1081,N_4946);
or U9146 (N_9146,N_1818,N_3109);
nor U9147 (N_9147,N_4501,N_1650);
nor U9148 (N_9148,N_3763,N_2139);
nand U9149 (N_9149,N_3102,N_2801);
nand U9150 (N_9150,N_4825,N_4820);
or U9151 (N_9151,N_2843,N_226);
nor U9152 (N_9152,N_4166,N_4213);
and U9153 (N_9153,N_979,N_3292);
nor U9154 (N_9154,N_2246,N_2594);
and U9155 (N_9155,N_1936,N_4752);
nand U9156 (N_9156,N_3113,N_2743);
nor U9157 (N_9157,N_2732,N_4175);
and U9158 (N_9158,N_2589,N_1668);
nor U9159 (N_9159,N_4537,N_4375);
nand U9160 (N_9160,N_2031,N_951);
nor U9161 (N_9161,N_496,N_3628);
or U9162 (N_9162,N_1445,N_1057);
nand U9163 (N_9163,N_1206,N_697);
nor U9164 (N_9164,N_2322,N_4342);
or U9165 (N_9165,N_515,N_2922);
nor U9166 (N_9166,N_4037,N_1520);
or U9167 (N_9167,N_3078,N_4199);
or U9168 (N_9168,N_1535,N_243);
nor U9169 (N_9169,N_3670,N_1996);
nand U9170 (N_9170,N_1262,N_2437);
nand U9171 (N_9171,N_2606,N_3049);
and U9172 (N_9172,N_4032,N_1415);
or U9173 (N_9173,N_4897,N_3747);
and U9174 (N_9174,N_1091,N_360);
and U9175 (N_9175,N_4523,N_1580);
or U9176 (N_9176,N_1237,N_108);
nand U9177 (N_9177,N_1570,N_2844);
nor U9178 (N_9178,N_1342,N_393);
nor U9179 (N_9179,N_1046,N_3631);
nor U9180 (N_9180,N_2587,N_1512);
nand U9181 (N_9181,N_1004,N_3731);
or U9182 (N_9182,N_241,N_43);
nand U9183 (N_9183,N_2947,N_1594);
nand U9184 (N_9184,N_3426,N_2575);
and U9185 (N_9185,N_1800,N_3690);
nand U9186 (N_9186,N_4023,N_4694);
and U9187 (N_9187,N_3185,N_2201);
or U9188 (N_9188,N_3366,N_4305);
or U9189 (N_9189,N_575,N_1068);
and U9190 (N_9190,N_1884,N_547);
nand U9191 (N_9191,N_537,N_1057);
nand U9192 (N_9192,N_4706,N_4877);
and U9193 (N_9193,N_489,N_1455);
nor U9194 (N_9194,N_714,N_3130);
nor U9195 (N_9195,N_3313,N_4960);
and U9196 (N_9196,N_2659,N_1875);
nand U9197 (N_9197,N_1004,N_351);
or U9198 (N_9198,N_1985,N_1939);
and U9199 (N_9199,N_4811,N_3476);
or U9200 (N_9200,N_4881,N_3397);
or U9201 (N_9201,N_407,N_2057);
and U9202 (N_9202,N_143,N_3062);
nor U9203 (N_9203,N_4676,N_4692);
or U9204 (N_9204,N_4028,N_1158);
or U9205 (N_9205,N_241,N_4787);
nor U9206 (N_9206,N_3081,N_826);
and U9207 (N_9207,N_3396,N_1960);
nand U9208 (N_9208,N_4919,N_65);
and U9209 (N_9209,N_3794,N_2627);
or U9210 (N_9210,N_4138,N_3508);
nor U9211 (N_9211,N_3367,N_4677);
nand U9212 (N_9212,N_3483,N_2390);
nor U9213 (N_9213,N_3170,N_3561);
and U9214 (N_9214,N_2257,N_4094);
and U9215 (N_9215,N_293,N_2537);
or U9216 (N_9216,N_3899,N_900);
nor U9217 (N_9217,N_4997,N_2605);
nand U9218 (N_9218,N_4341,N_2584);
and U9219 (N_9219,N_1381,N_1841);
nand U9220 (N_9220,N_3035,N_3504);
nand U9221 (N_9221,N_4713,N_4516);
or U9222 (N_9222,N_3159,N_4975);
and U9223 (N_9223,N_899,N_3663);
nor U9224 (N_9224,N_504,N_4906);
nand U9225 (N_9225,N_1604,N_1406);
nor U9226 (N_9226,N_1965,N_1211);
nor U9227 (N_9227,N_1897,N_3619);
or U9228 (N_9228,N_4149,N_4306);
and U9229 (N_9229,N_2184,N_1394);
and U9230 (N_9230,N_141,N_4103);
and U9231 (N_9231,N_3313,N_4973);
nand U9232 (N_9232,N_2685,N_3490);
nand U9233 (N_9233,N_808,N_3684);
nand U9234 (N_9234,N_2086,N_4170);
or U9235 (N_9235,N_2225,N_1007);
or U9236 (N_9236,N_2376,N_2187);
or U9237 (N_9237,N_4612,N_1988);
or U9238 (N_9238,N_1528,N_3389);
nand U9239 (N_9239,N_1587,N_4279);
and U9240 (N_9240,N_1836,N_4311);
or U9241 (N_9241,N_2547,N_2619);
or U9242 (N_9242,N_3887,N_2133);
and U9243 (N_9243,N_1255,N_2183);
nand U9244 (N_9244,N_3720,N_4058);
nand U9245 (N_9245,N_2349,N_4125);
nor U9246 (N_9246,N_337,N_2839);
nand U9247 (N_9247,N_3952,N_2314);
nand U9248 (N_9248,N_376,N_3642);
and U9249 (N_9249,N_418,N_1631);
nand U9250 (N_9250,N_1518,N_24);
nand U9251 (N_9251,N_3327,N_198);
nand U9252 (N_9252,N_1760,N_4682);
nand U9253 (N_9253,N_3807,N_1926);
nor U9254 (N_9254,N_1319,N_1846);
and U9255 (N_9255,N_2877,N_3466);
or U9256 (N_9256,N_1619,N_4822);
and U9257 (N_9257,N_4507,N_42);
and U9258 (N_9258,N_3962,N_1934);
nand U9259 (N_9259,N_490,N_797);
nand U9260 (N_9260,N_2690,N_406);
nor U9261 (N_9261,N_353,N_3824);
nand U9262 (N_9262,N_1574,N_1619);
and U9263 (N_9263,N_3232,N_4840);
nor U9264 (N_9264,N_263,N_1975);
and U9265 (N_9265,N_1914,N_1107);
or U9266 (N_9266,N_1289,N_540);
nor U9267 (N_9267,N_2513,N_4025);
and U9268 (N_9268,N_3248,N_947);
nor U9269 (N_9269,N_3522,N_4858);
nor U9270 (N_9270,N_3814,N_1786);
nor U9271 (N_9271,N_149,N_3120);
or U9272 (N_9272,N_1393,N_3623);
nor U9273 (N_9273,N_1924,N_904);
nand U9274 (N_9274,N_4143,N_1788);
and U9275 (N_9275,N_3950,N_2404);
or U9276 (N_9276,N_2203,N_4803);
or U9277 (N_9277,N_359,N_2062);
and U9278 (N_9278,N_3809,N_3806);
nand U9279 (N_9279,N_3738,N_4815);
and U9280 (N_9280,N_3586,N_4689);
and U9281 (N_9281,N_2516,N_1966);
nand U9282 (N_9282,N_4394,N_3844);
and U9283 (N_9283,N_2393,N_1789);
or U9284 (N_9284,N_4864,N_4932);
and U9285 (N_9285,N_1056,N_3996);
or U9286 (N_9286,N_2124,N_1899);
and U9287 (N_9287,N_311,N_691);
or U9288 (N_9288,N_4440,N_34);
nand U9289 (N_9289,N_3409,N_4532);
nand U9290 (N_9290,N_2998,N_4716);
nor U9291 (N_9291,N_1744,N_4173);
or U9292 (N_9292,N_2994,N_3471);
or U9293 (N_9293,N_3417,N_2583);
or U9294 (N_9294,N_4466,N_748);
nor U9295 (N_9295,N_4856,N_4242);
nor U9296 (N_9296,N_3980,N_2529);
or U9297 (N_9297,N_4472,N_247);
nor U9298 (N_9298,N_50,N_1641);
or U9299 (N_9299,N_3439,N_3859);
nor U9300 (N_9300,N_1654,N_161);
nor U9301 (N_9301,N_1229,N_4100);
or U9302 (N_9302,N_4285,N_1440);
nor U9303 (N_9303,N_1448,N_2344);
nor U9304 (N_9304,N_974,N_528);
nand U9305 (N_9305,N_2512,N_2565);
or U9306 (N_9306,N_275,N_1259);
and U9307 (N_9307,N_4815,N_4300);
or U9308 (N_9308,N_524,N_1670);
and U9309 (N_9309,N_3193,N_4345);
nand U9310 (N_9310,N_2040,N_3267);
xnor U9311 (N_9311,N_1607,N_1168);
nand U9312 (N_9312,N_4321,N_1465);
nand U9313 (N_9313,N_706,N_2273);
and U9314 (N_9314,N_4465,N_3158);
and U9315 (N_9315,N_1014,N_767);
or U9316 (N_9316,N_4534,N_2360);
or U9317 (N_9317,N_2265,N_2221);
or U9318 (N_9318,N_3062,N_1941);
and U9319 (N_9319,N_4972,N_2084);
or U9320 (N_9320,N_3576,N_2230);
and U9321 (N_9321,N_4284,N_4427);
and U9322 (N_9322,N_3380,N_882);
nor U9323 (N_9323,N_3750,N_3337);
and U9324 (N_9324,N_2870,N_1953);
or U9325 (N_9325,N_2328,N_4833);
nor U9326 (N_9326,N_712,N_4317);
nand U9327 (N_9327,N_2389,N_3052);
nor U9328 (N_9328,N_4921,N_2372);
and U9329 (N_9329,N_2223,N_4563);
nor U9330 (N_9330,N_1105,N_1181);
nand U9331 (N_9331,N_827,N_4559);
and U9332 (N_9332,N_1014,N_3644);
nor U9333 (N_9333,N_4917,N_318);
nand U9334 (N_9334,N_1432,N_4288);
nor U9335 (N_9335,N_1723,N_1314);
and U9336 (N_9336,N_4830,N_1335);
and U9337 (N_9337,N_171,N_3978);
nand U9338 (N_9338,N_4418,N_2356);
and U9339 (N_9339,N_1005,N_4434);
and U9340 (N_9340,N_3930,N_2635);
nor U9341 (N_9341,N_3568,N_2552);
and U9342 (N_9342,N_3100,N_4218);
nor U9343 (N_9343,N_2678,N_132);
and U9344 (N_9344,N_2335,N_3112);
and U9345 (N_9345,N_644,N_2204);
or U9346 (N_9346,N_1363,N_3376);
and U9347 (N_9347,N_3065,N_2538);
and U9348 (N_9348,N_3573,N_1737);
or U9349 (N_9349,N_1650,N_3365);
and U9350 (N_9350,N_2397,N_4370);
nand U9351 (N_9351,N_271,N_3807);
or U9352 (N_9352,N_4774,N_2542);
nor U9353 (N_9353,N_3741,N_2505);
or U9354 (N_9354,N_653,N_2269);
or U9355 (N_9355,N_2447,N_2414);
or U9356 (N_9356,N_3549,N_125);
or U9357 (N_9357,N_1981,N_4434);
nand U9358 (N_9358,N_2647,N_4869);
nor U9359 (N_9359,N_3680,N_2995);
or U9360 (N_9360,N_4341,N_2506);
and U9361 (N_9361,N_614,N_3150);
and U9362 (N_9362,N_219,N_794);
nor U9363 (N_9363,N_2610,N_1624);
and U9364 (N_9364,N_1452,N_1364);
nor U9365 (N_9365,N_3510,N_3994);
or U9366 (N_9366,N_1748,N_1851);
or U9367 (N_9367,N_4922,N_1718);
nor U9368 (N_9368,N_3040,N_4350);
and U9369 (N_9369,N_1268,N_4835);
and U9370 (N_9370,N_3502,N_1121);
nand U9371 (N_9371,N_2986,N_431);
and U9372 (N_9372,N_1515,N_1645);
and U9373 (N_9373,N_1542,N_1037);
nand U9374 (N_9374,N_1127,N_1019);
or U9375 (N_9375,N_662,N_3438);
or U9376 (N_9376,N_27,N_559);
and U9377 (N_9377,N_1789,N_1180);
or U9378 (N_9378,N_2711,N_4944);
and U9379 (N_9379,N_901,N_1184);
or U9380 (N_9380,N_2343,N_1660);
nor U9381 (N_9381,N_3674,N_3839);
and U9382 (N_9382,N_2423,N_4909);
and U9383 (N_9383,N_404,N_1499);
nand U9384 (N_9384,N_1642,N_1353);
nand U9385 (N_9385,N_2989,N_843);
or U9386 (N_9386,N_444,N_3921);
and U9387 (N_9387,N_3760,N_3933);
nand U9388 (N_9388,N_4955,N_427);
nor U9389 (N_9389,N_1891,N_710);
nor U9390 (N_9390,N_132,N_1976);
nor U9391 (N_9391,N_2933,N_4861);
nand U9392 (N_9392,N_4761,N_1580);
and U9393 (N_9393,N_2335,N_4741);
or U9394 (N_9394,N_1033,N_3998);
nand U9395 (N_9395,N_663,N_3784);
or U9396 (N_9396,N_4624,N_1228);
and U9397 (N_9397,N_926,N_4710);
nor U9398 (N_9398,N_2683,N_1556);
or U9399 (N_9399,N_415,N_1951);
nor U9400 (N_9400,N_3905,N_3134);
or U9401 (N_9401,N_4335,N_4216);
or U9402 (N_9402,N_3824,N_2816);
and U9403 (N_9403,N_596,N_535);
nand U9404 (N_9404,N_2565,N_4716);
and U9405 (N_9405,N_4830,N_3630);
or U9406 (N_9406,N_599,N_3878);
and U9407 (N_9407,N_3513,N_1902);
or U9408 (N_9408,N_3813,N_2389);
xnor U9409 (N_9409,N_2215,N_1968);
nand U9410 (N_9410,N_3717,N_2418);
and U9411 (N_9411,N_3857,N_241);
and U9412 (N_9412,N_1539,N_3879);
nor U9413 (N_9413,N_4902,N_3804);
and U9414 (N_9414,N_1614,N_2724);
or U9415 (N_9415,N_4018,N_3337);
or U9416 (N_9416,N_138,N_3397);
and U9417 (N_9417,N_952,N_477);
nor U9418 (N_9418,N_4795,N_2623);
nand U9419 (N_9419,N_631,N_2567);
nand U9420 (N_9420,N_2185,N_3376);
or U9421 (N_9421,N_158,N_614);
or U9422 (N_9422,N_2727,N_122);
nor U9423 (N_9423,N_4723,N_3480);
and U9424 (N_9424,N_3038,N_117);
or U9425 (N_9425,N_2919,N_4797);
and U9426 (N_9426,N_3797,N_2966);
nor U9427 (N_9427,N_1639,N_4891);
nor U9428 (N_9428,N_3904,N_85);
or U9429 (N_9429,N_4999,N_988);
and U9430 (N_9430,N_4174,N_3646);
nor U9431 (N_9431,N_2512,N_1171);
nand U9432 (N_9432,N_4259,N_3563);
nor U9433 (N_9433,N_3194,N_287);
or U9434 (N_9434,N_3847,N_3580);
or U9435 (N_9435,N_1431,N_4777);
or U9436 (N_9436,N_1907,N_1077);
nand U9437 (N_9437,N_3230,N_652);
nand U9438 (N_9438,N_3828,N_1481);
and U9439 (N_9439,N_3863,N_2144);
nand U9440 (N_9440,N_4103,N_2162);
nor U9441 (N_9441,N_2976,N_88);
nor U9442 (N_9442,N_3448,N_3937);
nand U9443 (N_9443,N_4975,N_2061);
or U9444 (N_9444,N_333,N_2930);
nand U9445 (N_9445,N_2559,N_1190);
or U9446 (N_9446,N_4016,N_1534);
and U9447 (N_9447,N_87,N_2665);
nand U9448 (N_9448,N_813,N_3022);
or U9449 (N_9449,N_2662,N_3721);
or U9450 (N_9450,N_1024,N_684);
or U9451 (N_9451,N_4675,N_546);
or U9452 (N_9452,N_1235,N_1408);
or U9453 (N_9453,N_4706,N_837);
and U9454 (N_9454,N_394,N_3718);
or U9455 (N_9455,N_4957,N_2177);
nand U9456 (N_9456,N_3320,N_1992);
and U9457 (N_9457,N_4350,N_2727);
nor U9458 (N_9458,N_447,N_3624);
and U9459 (N_9459,N_2499,N_376);
and U9460 (N_9460,N_36,N_2600);
or U9461 (N_9461,N_784,N_2975);
nand U9462 (N_9462,N_3214,N_2593);
nand U9463 (N_9463,N_1254,N_2745);
or U9464 (N_9464,N_3953,N_1849);
nor U9465 (N_9465,N_1415,N_3);
or U9466 (N_9466,N_53,N_4281);
or U9467 (N_9467,N_291,N_1473);
nor U9468 (N_9468,N_3623,N_4538);
or U9469 (N_9469,N_3529,N_2196);
nand U9470 (N_9470,N_2142,N_4630);
nand U9471 (N_9471,N_1009,N_1080);
and U9472 (N_9472,N_1312,N_3453);
or U9473 (N_9473,N_685,N_378);
and U9474 (N_9474,N_439,N_1339);
or U9475 (N_9475,N_4233,N_3729);
nor U9476 (N_9476,N_973,N_2842);
nor U9477 (N_9477,N_2414,N_333);
nor U9478 (N_9478,N_4498,N_245);
nand U9479 (N_9479,N_754,N_2182);
or U9480 (N_9480,N_583,N_3994);
or U9481 (N_9481,N_2575,N_4724);
nand U9482 (N_9482,N_2214,N_3368);
or U9483 (N_9483,N_4973,N_1352);
and U9484 (N_9484,N_446,N_2988);
and U9485 (N_9485,N_352,N_1913);
nand U9486 (N_9486,N_1073,N_237);
nor U9487 (N_9487,N_1652,N_3781);
nor U9488 (N_9488,N_4694,N_1237);
and U9489 (N_9489,N_1215,N_3383);
and U9490 (N_9490,N_4302,N_0);
nor U9491 (N_9491,N_830,N_1015);
nand U9492 (N_9492,N_2616,N_3388);
and U9493 (N_9493,N_1709,N_4243);
nor U9494 (N_9494,N_2741,N_4113);
xor U9495 (N_9495,N_3433,N_3359);
or U9496 (N_9496,N_524,N_4108);
and U9497 (N_9497,N_976,N_2552);
nand U9498 (N_9498,N_3787,N_4029);
and U9499 (N_9499,N_230,N_2603);
nor U9500 (N_9500,N_1893,N_745);
and U9501 (N_9501,N_3305,N_4514);
or U9502 (N_9502,N_2223,N_446);
nand U9503 (N_9503,N_3180,N_776);
nor U9504 (N_9504,N_3741,N_1960);
nor U9505 (N_9505,N_3173,N_2119);
and U9506 (N_9506,N_438,N_4541);
nor U9507 (N_9507,N_2814,N_3307);
or U9508 (N_9508,N_1138,N_3685);
nor U9509 (N_9509,N_4845,N_4192);
and U9510 (N_9510,N_1874,N_2113);
nor U9511 (N_9511,N_3732,N_1331);
nor U9512 (N_9512,N_2617,N_2760);
nor U9513 (N_9513,N_2408,N_3207);
nor U9514 (N_9514,N_252,N_3497);
or U9515 (N_9515,N_1291,N_3681);
nor U9516 (N_9516,N_863,N_3585);
and U9517 (N_9517,N_2673,N_827);
nor U9518 (N_9518,N_2365,N_1544);
nor U9519 (N_9519,N_2191,N_1342);
nor U9520 (N_9520,N_4803,N_408);
and U9521 (N_9521,N_3971,N_4809);
or U9522 (N_9522,N_384,N_4378);
nand U9523 (N_9523,N_3416,N_4854);
nor U9524 (N_9524,N_796,N_498);
nand U9525 (N_9525,N_1671,N_4095);
or U9526 (N_9526,N_3073,N_2995);
and U9527 (N_9527,N_2158,N_4848);
and U9528 (N_9528,N_1840,N_4095);
and U9529 (N_9529,N_1308,N_4199);
nand U9530 (N_9530,N_882,N_103);
nor U9531 (N_9531,N_2413,N_4371);
nor U9532 (N_9532,N_1001,N_1171);
or U9533 (N_9533,N_1950,N_1065);
nand U9534 (N_9534,N_1144,N_3888);
or U9535 (N_9535,N_4740,N_4821);
or U9536 (N_9536,N_2774,N_4326);
or U9537 (N_9537,N_3653,N_3689);
nor U9538 (N_9538,N_1278,N_3349);
and U9539 (N_9539,N_252,N_4032);
and U9540 (N_9540,N_1289,N_2937);
nand U9541 (N_9541,N_3680,N_4187);
nand U9542 (N_9542,N_430,N_4733);
and U9543 (N_9543,N_776,N_2766);
nand U9544 (N_9544,N_3902,N_2373);
and U9545 (N_9545,N_2985,N_3554);
nand U9546 (N_9546,N_1063,N_1521);
and U9547 (N_9547,N_1344,N_2246);
nor U9548 (N_9548,N_4211,N_4825);
and U9549 (N_9549,N_3998,N_2321);
or U9550 (N_9550,N_1448,N_4591);
nand U9551 (N_9551,N_779,N_1786);
or U9552 (N_9552,N_4564,N_1101);
and U9553 (N_9553,N_4419,N_4);
and U9554 (N_9554,N_2963,N_213);
and U9555 (N_9555,N_661,N_178);
nand U9556 (N_9556,N_2964,N_2736);
nand U9557 (N_9557,N_2807,N_1094);
nand U9558 (N_9558,N_2231,N_1091);
or U9559 (N_9559,N_3667,N_3776);
nand U9560 (N_9560,N_3817,N_620);
and U9561 (N_9561,N_2527,N_719);
and U9562 (N_9562,N_1094,N_1750);
nor U9563 (N_9563,N_2642,N_1909);
nor U9564 (N_9564,N_2417,N_1579);
and U9565 (N_9565,N_2501,N_1834);
and U9566 (N_9566,N_580,N_3696);
nor U9567 (N_9567,N_1833,N_3104);
nor U9568 (N_9568,N_2344,N_1596);
and U9569 (N_9569,N_4961,N_3990);
nor U9570 (N_9570,N_1918,N_2070);
nor U9571 (N_9571,N_934,N_2012);
nor U9572 (N_9572,N_3787,N_3778);
and U9573 (N_9573,N_1697,N_838);
nor U9574 (N_9574,N_315,N_1395);
nand U9575 (N_9575,N_2626,N_348);
nand U9576 (N_9576,N_2616,N_3233);
nand U9577 (N_9577,N_1416,N_2108);
and U9578 (N_9578,N_3094,N_1692);
nand U9579 (N_9579,N_3138,N_3995);
nor U9580 (N_9580,N_158,N_1314);
or U9581 (N_9581,N_386,N_3507);
and U9582 (N_9582,N_3155,N_353);
and U9583 (N_9583,N_3106,N_564);
nand U9584 (N_9584,N_639,N_678);
nor U9585 (N_9585,N_2113,N_4271);
nor U9586 (N_9586,N_4319,N_1375);
nor U9587 (N_9587,N_1183,N_1703);
and U9588 (N_9588,N_3455,N_968);
and U9589 (N_9589,N_2563,N_3105);
and U9590 (N_9590,N_662,N_182);
xor U9591 (N_9591,N_2724,N_3915);
or U9592 (N_9592,N_3117,N_3064);
nand U9593 (N_9593,N_3749,N_3727);
xor U9594 (N_9594,N_4271,N_4135);
or U9595 (N_9595,N_236,N_1265);
and U9596 (N_9596,N_3620,N_717);
nand U9597 (N_9597,N_4497,N_1156);
nor U9598 (N_9598,N_1896,N_3137);
and U9599 (N_9599,N_359,N_3088);
nor U9600 (N_9600,N_1416,N_3732);
nor U9601 (N_9601,N_4333,N_166);
and U9602 (N_9602,N_4634,N_2465);
nand U9603 (N_9603,N_1636,N_4797);
or U9604 (N_9604,N_3237,N_4635);
xor U9605 (N_9605,N_1144,N_1222);
or U9606 (N_9606,N_2342,N_1174);
nand U9607 (N_9607,N_3441,N_4886);
and U9608 (N_9608,N_1689,N_927);
or U9609 (N_9609,N_1541,N_1755);
or U9610 (N_9610,N_4656,N_1748);
nand U9611 (N_9611,N_489,N_2668);
or U9612 (N_9612,N_4364,N_1632);
and U9613 (N_9613,N_1448,N_4038);
and U9614 (N_9614,N_4082,N_1319);
nor U9615 (N_9615,N_2563,N_3150);
nor U9616 (N_9616,N_1957,N_106);
nand U9617 (N_9617,N_460,N_1975);
and U9618 (N_9618,N_4182,N_4598);
and U9619 (N_9619,N_859,N_321);
nand U9620 (N_9620,N_2133,N_1890);
or U9621 (N_9621,N_910,N_2071);
and U9622 (N_9622,N_2641,N_3010);
nor U9623 (N_9623,N_3188,N_4256);
or U9624 (N_9624,N_3630,N_692);
or U9625 (N_9625,N_727,N_1523);
nand U9626 (N_9626,N_4339,N_1549);
nand U9627 (N_9627,N_682,N_3734);
and U9628 (N_9628,N_691,N_337);
nor U9629 (N_9629,N_1499,N_2318);
and U9630 (N_9630,N_1747,N_3303);
nor U9631 (N_9631,N_3124,N_3629);
or U9632 (N_9632,N_4946,N_4653);
and U9633 (N_9633,N_2980,N_4400);
nor U9634 (N_9634,N_1412,N_4621);
nand U9635 (N_9635,N_159,N_3604);
and U9636 (N_9636,N_1120,N_3644);
and U9637 (N_9637,N_3,N_941);
nor U9638 (N_9638,N_1189,N_1268);
or U9639 (N_9639,N_4760,N_4423);
and U9640 (N_9640,N_1733,N_363);
and U9641 (N_9641,N_3721,N_4497);
and U9642 (N_9642,N_1478,N_1318);
or U9643 (N_9643,N_964,N_848);
nand U9644 (N_9644,N_584,N_216);
or U9645 (N_9645,N_2190,N_4544);
nor U9646 (N_9646,N_4197,N_2274);
or U9647 (N_9647,N_4013,N_2311);
nor U9648 (N_9648,N_4157,N_2032);
and U9649 (N_9649,N_3433,N_1922);
nor U9650 (N_9650,N_4400,N_4354);
and U9651 (N_9651,N_272,N_3120);
or U9652 (N_9652,N_1222,N_1862);
nor U9653 (N_9653,N_3004,N_2272);
and U9654 (N_9654,N_3506,N_2475);
nand U9655 (N_9655,N_3787,N_2683);
and U9656 (N_9656,N_1005,N_2444);
and U9657 (N_9657,N_4054,N_339);
nor U9658 (N_9658,N_3460,N_3473);
nand U9659 (N_9659,N_3757,N_2660);
nor U9660 (N_9660,N_692,N_143);
and U9661 (N_9661,N_60,N_2630);
nor U9662 (N_9662,N_3634,N_315);
nand U9663 (N_9663,N_2903,N_3023);
nand U9664 (N_9664,N_4933,N_668);
nor U9665 (N_9665,N_2888,N_1361);
nor U9666 (N_9666,N_1852,N_1078);
and U9667 (N_9667,N_1248,N_2467);
nand U9668 (N_9668,N_3096,N_3442);
nand U9669 (N_9669,N_1064,N_3324);
and U9670 (N_9670,N_2787,N_259);
or U9671 (N_9671,N_1194,N_4363);
and U9672 (N_9672,N_3939,N_4004);
or U9673 (N_9673,N_3407,N_3364);
and U9674 (N_9674,N_1931,N_1038);
nand U9675 (N_9675,N_393,N_1606);
nor U9676 (N_9676,N_3430,N_875);
nand U9677 (N_9677,N_1569,N_966);
and U9678 (N_9678,N_3963,N_1680);
nor U9679 (N_9679,N_3846,N_3882);
nand U9680 (N_9680,N_2289,N_885);
or U9681 (N_9681,N_1488,N_2907);
nand U9682 (N_9682,N_3462,N_1470);
xnor U9683 (N_9683,N_3526,N_4358);
and U9684 (N_9684,N_383,N_1408);
and U9685 (N_9685,N_2376,N_2612);
or U9686 (N_9686,N_4491,N_2216);
nor U9687 (N_9687,N_3128,N_4410);
nand U9688 (N_9688,N_2937,N_4588);
and U9689 (N_9689,N_189,N_4863);
nor U9690 (N_9690,N_3407,N_4979);
and U9691 (N_9691,N_4948,N_1068);
and U9692 (N_9692,N_1139,N_1475);
and U9693 (N_9693,N_1006,N_238);
nor U9694 (N_9694,N_469,N_5);
nand U9695 (N_9695,N_527,N_4428);
nor U9696 (N_9696,N_1945,N_4203);
nand U9697 (N_9697,N_4148,N_2737);
nand U9698 (N_9698,N_3355,N_2680);
and U9699 (N_9699,N_774,N_2089);
and U9700 (N_9700,N_898,N_3881);
nor U9701 (N_9701,N_3088,N_2910);
or U9702 (N_9702,N_4647,N_3627);
or U9703 (N_9703,N_3538,N_2801);
nor U9704 (N_9704,N_4950,N_1287);
and U9705 (N_9705,N_1172,N_69);
nand U9706 (N_9706,N_2086,N_3449);
or U9707 (N_9707,N_4990,N_3564);
or U9708 (N_9708,N_2752,N_576);
nand U9709 (N_9709,N_3204,N_2434);
and U9710 (N_9710,N_117,N_1525);
nor U9711 (N_9711,N_4073,N_1634);
and U9712 (N_9712,N_1361,N_221);
nor U9713 (N_9713,N_633,N_1032);
and U9714 (N_9714,N_2982,N_3528);
nand U9715 (N_9715,N_530,N_345);
nand U9716 (N_9716,N_2736,N_4966);
or U9717 (N_9717,N_883,N_487);
nand U9718 (N_9718,N_4931,N_434);
and U9719 (N_9719,N_564,N_1457);
nand U9720 (N_9720,N_3843,N_1579);
nand U9721 (N_9721,N_2762,N_1530);
or U9722 (N_9722,N_2068,N_3950);
nand U9723 (N_9723,N_435,N_857);
and U9724 (N_9724,N_2363,N_1232);
and U9725 (N_9725,N_4116,N_1392);
nand U9726 (N_9726,N_4846,N_4343);
nor U9727 (N_9727,N_4168,N_1757);
or U9728 (N_9728,N_3944,N_3596);
nand U9729 (N_9729,N_3792,N_1325);
or U9730 (N_9730,N_4725,N_3097);
nor U9731 (N_9731,N_1161,N_4105);
or U9732 (N_9732,N_3374,N_2672);
and U9733 (N_9733,N_3505,N_3072);
nor U9734 (N_9734,N_1966,N_2547);
or U9735 (N_9735,N_3374,N_1373);
or U9736 (N_9736,N_2377,N_3335);
nor U9737 (N_9737,N_552,N_4359);
and U9738 (N_9738,N_196,N_176);
and U9739 (N_9739,N_4306,N_1118);
nor U9740 (N_9740,N_866,N_4765);
or U9741 (N_9741,N_926,N_3389);
nor U9742 (N_9742,N_2093,N_353);
and U9743 (N_9743,N_4284,N_4676);
and U9744 (N_9744,N_3231,N_2461);
or U9745 (N_9745,N_4748,N_2408);
xor U9746 (N_9746,N_2471,N_2694);
or U9747 (N_9747,N_1591,N_4212);
or U9748 (N_9748,N_2882,N_4017);
or U9749 (N_9749,N_3538,N_3190);
nor U9750 (N_9750,N_2227,N_517);
nand U9751 (N_9751,N_641,N_1620);
nor U9752 (N_9752,N_2682,N_1224);
or U9753 (N_9753,N_1310,N_92);
nor U9754 (N_9754,N_4358,N_4167);
and U9755 (N_9755,N_1612,N_1714);
nor U9756 (N_9756,N_4829,N_3729);
or U9757 (N_9757,N_2679,N_482);
and U9758 (N_9758,N_4724,N_1277);
or U9759 (N_9759,N_2972,N_1814);
nor U9760 (N_9760,N_1676,N_3276);
nand U9761 (N_9761,N_248,N_1561);
nor U9762 (N_9762,N_32,N_2193);
nand U9763 (N_9763,N_721,N_288);
and U9764 (N_9764,N_4690,N_818);
nor U9765 (N_9765,N_1424,N_332);
nand U9766 (N_9766,N_2168,N_3354);
or U9767 (N_9767,N_3253,N_2705);
or U9768 (N_9768,N_3242,N_1712);
nand U9769 (N_9769,N_104,N_1440);
nand U9770 (N_9770,N_90,N_1939);
or U9771 (N_9771,N_4704,N_4707);
nor U9772 (N_9772,N_3280,N_657);
nor U9773 (N_9773,N_2670,N_674);
and U9774 (N_9774,N_1674,N_2754);
nor U9775 (N_9775,N_4211,N_2506);
nand U9776 (N_9776,N_4989,N_4984);
nor U9777 (N_9777,N_2364,N_233);
or U9778 (N_9778,N_4549,N_691);
nor U9779 (N_9779,N_4875,N_499);
nand U9780 (N_9780,N_4140,N_729);
nor U9781 (N_9781,N_1669,N_29);
and U9782 (N_9782,N_666,N_4860);
and U9783 (N_9783,N_1553,N_3121);
nor U9784 (N_9784,N_3720,N_3715);
or U9785 (N_9785,N_1581,N_1783);
and U9786 (N_9786,N_2602,N_2886);
nand U9787 (N_9787,N_3119,N_473);
nand U9788 (N_9788,N_4335,N_691);
and U9789 (N_9789,N_2936,N_2041);
nor U9790 (N_9790,N_4119,N_2799);
nor U9791 (N_9791,N_4916,N_4971);
nand U9792 (N_9792,N_2669,N_2507);
and U9793 (N_9793,N_2572,N_1917);
or U9794 (N_9794,N_4451,N_1322);
nor U9795 (N_9795,N_2942,N_4096);
or U9796 (N_9796,N_3485,N_2305);
and U9797 (N_9797,N_1178,N_2386);
nand U9798 (N_9798,N_4240,N_4356);
nor U9799 (N_9799,N_40,N_3801);
nor U9800 (N_9800,N_988,N_4148);
nor U9801 (N_9801,N_4816,N_2118);
and U9802 (N_9802,N_3003,N_748);
nor U9803 (N_9803,N_1500,N_772);
and U9804 (N_9804,N_985,N_1330);
and U9805 (N_9805,N_4169,N_3700);
and U9806 (N_9806,N_1455,N_2585);
and U9807 (N_9807,N_56,N_4508);
nor U9808 (N_9808,N_4274,N_4451);
nand U9809 (N_9809,N_756,N_2747);
and U9810 (N_9810,N_2712,N_3111);
or U9811 (N_9811,N_4951,N_3105);
and U9812 (N_9812,N_1073,N_3001);
and U9813 (N_9813,N_4952,N_4437);
nor U9814 (N_9814,N_3391,N_692);
and U9815 (N_9815,N_1405,N_3005);
nor U9816 (N_9816,N_1039,N_4137);
and U9817 (N_9817,N_715,N_2680);
or U9818 (N_9818,N_3766,N_3931);
and U9819 (N_9819,N_4577,N_3572);
nor U9820 (N_9820,N_4702,N_463);
or U9821 (N_9821,N_4963,N_2145);
nor U9822 (N_9822,N_3683,N_3417);
nand U9823 (N_9823,N_14,N_2348);
nand U9824 (N_9824,N_611,N_1830);
nor U9825 (N_9825,N_2789,N_2575);
and U9826 (N_9826,N_530,N_2629);
and U9827 (N_9827,N_849,N_382);
nand U9828 (N_9828,N_4986,N_3631);
nor U9829 (N_9829,N_3235,N_3973);
nand U9830 (N_9830,N_3123,N_1909);
nand U9831 (N_9831,N_351,N_2337);
nor U9832 (N_9832,N_3689,N_1996);
or U9833 (N_9833,N_98,N_4839);
nor U9834 (N_9834,N_707,N_2805);
nand U9835 (N_9835,N_3318,N_4867);
nor U9836 (N_9836,N_1179,N_1919);
or U9837 (N_9837,N_4211,N_631);
or U9838 (N_9838,N_3199,N_4078);
or U9839 (N_9839,N_4004,N_171);
or U9840 (N_9840,N_4401,N_3671);
and U9841 (N_9841,N_1464,N_3697);
nor U9842 (N_9842,N_4181,N_2638);
and U9843 (N_9843,N_3912,N_0);
nand U9844 (N_9844,N_532,N_2461);
and U9845 (N_9845,N_1072,N_3189);
and U9846 (N_9846,N_3466,N_1924);
and U9847 (N_9847,N_2008,N_4896);
and U9848 (N_9848,N_4508,N_4337);
nand U9849 (N_9849,N_4985,N_984);
or U9850 (N_9850,N_3297,N_4341);
nand U9851 (N_9851,N_1375,N_3110);
nor U9852 (N_9852,N_3623,N_648);
and U9853 (N_9853,N_2823,N_1916);
and U9854 (N_9854,N_2797,N_2518);
nand U9855 (N_9855,N_4289,N_1657);
nor U9856 (N_9856,N_2854,N_2926);
nor U9857 (N_9857,N_3396,N_26);
nor U9858 (N_9858,N_1780,N_1138);
nand U9859 (N_9859,N_3427,N_2417);
and U9860 (N_9860,N_2270,N_2751);
nor U9861 (N_9861,N_3062,N_2645);
or U9862 (N_9862,N_4064,N_1850);
or U9863 (N_9863,N_3816,N_805);
nand U9864 (N_9864,N_1,N_924);
and U9865 (N_9865,N_1887,N_1675);
or U9866 (N_9866,N_200,N_2069);
nor U9867 (N_9867,N_3753,N_2860);
nor U9868 (N_9868,N_687,N_2171);
nor U9869 (N_9869,N_2701,N_3030);
and U9870 (N_9870,N_33,N_4752);
nand U9871 (N_9871,N_1276,N_454);
nor U9872 (N_9872,N_2389,N_1440);
nor U9873 (N_9873,N_2910,N_4522);
and U9874 (N_9874,N_162,N_3622);
and U9875 (N_9875,N_3887,N_3048);
nand U9876 (N_9876,N_3559,N_292);
nor U9877 (N_9877,N_4489,N_2325);
or U9878 (N_9878,N_2881,N_4414);
and U9879 (N_9879,N_1885,N_1995);
nand U9880 (N_9880,N_4379,N_1694);
and U9881 (N_9881,N_1916,N_3561);
nor U9882 (N_9882,N_2178,N_3533);
and U9883 (N_9883,N_137,N_740);
nor U9884 (N_9884,N_3357,N_2112);
and U9885 (N_9885,N_2454,N_3864);
nand U9886 (N_9886,N_4712,N_1547);
nand U9887 (N_9887,N_4220,N_3480);
nand U9888 (N_9888,N_3978,N_4866);
and U9889 (N_9889,N_2954,N_567);
nor U9890 (N_9890,N_544,N_60);
and U9891 (N_9891,N_1963,N_295);
or U9892 (N_9892,N_4586,N_3444);
nand U9893 (N_9893,N_3303,N_2989);
nand U9894 (N_9894,N_3313,N_2242);
and U9895 (N_9895,N_3782,N_1217);
or U9896 (N_9896,N_3284,N_2775);
nand U9897 (N_9897,N_517,N_1047);
and U9898 (N_9898,N_536,N_122);
nor U9899 (N_9899,N_1053,N_3249);
nand U9900 (N_9900,N_648,N_3294);
nor U9901 (N_9901,N_3146,N_808);
or U9902 (N_9902,N_3204,N_3977);
or U9903 (N_9903,N_1986,N_544);
or U9904 (N_9904,N_3247,N_91);
nor U9905 (N_9905,N_4084,N_873);
nand U9906 (N_9906,N_2063,N_2623);
nand U9907 (N_9907,N_4863,N_4855);
nand U9908 (N_9908,N_2095,N_1930);
nand U9909 (N_9909,N_544,N_1156);
nor U9910 (N_9910,N_3173,N_2278);
and U9911 (N_9911,N_3975,N_4853);
nor U9912 (N_9912,N_1164,N_2737);
and U9913 (N_9913,N_197,N_3861);
nand U9914 (N_9914,N_1787,N_461);
nand U9915 (N_9915,N_804,N_1397);
or U9916 (N_9916,N_3365,N_2666);
nor U9917 (N_9917,N_1137,N_965);
and U9918 (N_9918,N_2963,N_2035);
and U9919 (N_9919,N_239,N_4363);
nor U9920 (N_9920,N_219,N_1878);
nand U9921 (N_9921,N_658,N_4302);
and U9922 (N_9922,N_2874,N_4464);
and U9923 (N_9923,N_2661,N_958);
nor U9924 (N_9924,N_1542,N_3871);
nor U9925 (N_9925,N_113,N_1948);
xor U9926 (N_9926,N_4883,N_4366);
or U9927 (N_9927,N_4706,N_4790);
and U9928 (N_9928,N_2938,N_1024);
nand U9929 (N_9929,N_3925,N_3323);
or U9930 (N_9930,N_4965,N_217);
or U9931 (N_9931,N_49,N_3145);
or U9932 (N_9932,N_4627,N_1945);
or U9933 (N_9933,N_2688,N_2777);
or U9934 (N_9934,N_3546,N_1684);
or U9935 (N_9935,N_3309,N_1436);
and U9936 (N_9936,N_4084,N_4708);
and U9937 (N_9937,N_3867,N_1432);
nor U9938 (N_9938,N_4865,N_3908);
and U9939 (N_9939,N_2834,N_3299);
nand U9940 (N_9940,N_1267,N_3666);
nand U9941 (N_9941,N_3892,N_2986);
nand U9942 (N_9942,N_2086,N_1156);
or U9943 (N_9943,N_573,N_346);
or U9944 (N_9944,N_2517,N_4336);
and U9945 (N_9945,N_4424,N_1376);
nand U9946 (N_9946,N_4184,N_2251);
nor U9947 (N_9947,N_3138,N_1134);
or U9948 (N_9948,N_1816,N_2005);
or U9949 (N_9949,N_3909,N_4679);
and U9950 (N_9950,N_3169,N_3767);
nor U9951 (N_9951,N_3531,N_1897);
and U9952 (N_9952,N_2701,N_4463);
nand U9953 (N_9953,N_3033,N_2631);
or U9954 (N_9954,N_2549,N_1620);
and U9955 (N_9955,N_3270,N_4598);
or U9956 (N_9956,N_2008,N_4016);
nand U9957 (N_9957,N_1906,N_2954);
and U9958 (N_9958,N_3442,N_4228);
nor U9959 (N_9959,N_3633,N_3352);
and U9960 (N_9960,N_2402,N_3186);
and U9961 (N_9961,N_2778,N_4407);
or U9962 (N_9962,N_500,N_1321);
or U9963 (N_9963,N_3811,N_586);
or U9964 (N_9964,N_368,N_4739);
nand U9965 (N_9965,N_4872,N_1660);
xor U9966 (N_9966,N_125,N_4258);
nand U9967 (N_9967,N_4106,N_1369);
nor U9968 (N_9968,N_3105,N_924);
and U9969 (N_9969,N_2940,N_2659);
or U9970 (N_9970,N_2227,N_2502);
nor U9971 (N_9971,N_1228,N_3114);
and U9972 (N_9972,N_1231,N_4847);
nand U9973 (N_9973,N_4732,N_3068);
nand U9974 (N_9974,N_4699,N_4846);
or U9975 (N_9975,N_4210,N_721);
nand U9976 (N_9976,N_3438,N_3860);
or U9977 (N_9977,N_3248,N_510);
nand U9978 (N_9978,N_2936,N_3990);
or U9979 (N_9979,N_2536,N_99);
nor U9980 (N_9980,N_2700,N_1342);
and U9981 (N_9981,N_2086,N_3071);
nand U9982 (N_9982,N_39,N_792);
nor U9983 (N_9983,N_4011,N_2691);
nor U9984 (N_9984,N_3498,N_3710);
nand U9985 (N_9985,N_1785,N_1672);
and U9986 (N_9986,N_4670,N_261);
nand U9987 (N_9987,N_4091,N_1157);
nor U9988 (N_9988,N_4278,N_4681);
nand U9989 (N_9989,N_12,N_2637);
nor U9990 (N_9990,N_3762,N_2281);
or U9991 (N_9991,N_1338,N_2046);
nor U9992 (N_9992,N_2281,N_3117);
and U9993 (N_9993,N_3647,N_2111);
or U9994 (N_9994,N_3009,N_3381);
and U9995 (N_9995,N_4683,N_3011);
or U9996 (N_9996,N_3543,N_4988);
nand U9997 (N_9997,N_3976,N_1422);
nor U9998 (N_9998,N_262,N_1882);
or U9999 (N_9999,N_12,N_2859);
nand U10000 (N_10000,N_6023,N_9877);
or U10001 (N_10001,N_5833,N_6270);
and U10002 (N_10002,N_5568,N_9241);
nand U10003 (N_10003,N_6957,N_6018);
nor U10004 (N_10004,N_8569,N_7967);
nand U10005 (N_10005,N_8478,N_6642);
and U10006 (N_10006,N_8314,N_9891);
nor U10007 (N_10007,N_7752,N_5276);
or U10008 (N_10008,N_7651,N_8579);
and U10009 (N_10009,N_6946,N_7001);
or U10010 (N_10010,N_7061,N_6206);
and U10011 (N_10011,N_7251,N_9370);
or U10012 (N_10012,N_9402,N_6296);
and U10013 (N_10013,N_5404,N_6267);
nor U10014 (N_10014,N_6031,N_8455);
nand U10015 (N_10015,N_9478,N_9114);
or U10016 (N_10016,N_6523,N_5283);
nand U10017 (N_10017,N_6151,N_9300);
xnor U10018 (N_10018,N_9292,N_8610);
and U10019 (N_10019,N_6666,N_6036);
nand U10020 (N_10020,N_9349,N_7788);
nor U10021 (N_10021,N_9632,N_6974);
and U10022 (N_10022,N_9347,N_9919);
and U10023 (N_10023,N_5509,N_7910);
nand U10024 (N_10024,N_6803,N_9599);
or U10025 (N_10025,N_6375,N_9771);
and U10026 (N_10026,N_6188,N_5304);
or U10027 (N_10027,N_6086,N_7134);
and U10028 (N_10028,N_8309,N_9867);
nor U10029 (N_10029,N_8216,N_5146);
nand U10030 (N_10030,N_6937,N_8173);
and U10031 (N_10031,N_9480,N_9811);
or U10032 (N_10032,N_9000,N_6630);
and U10033 (N_10033,N_5908,N_5194);
nand U10034 (N_10034,N_5991,N_5686);
and U10035 (N_10035,N_5365,N_9812);
xnor U10036 (N_10036,N_9523,N_5047);
xnor U10037 (N_10037,N_6976,N_7580);
or U10038 (N_10038,N_7496,N_5101);
nor U10039 (N_10039,N_5263,N_9142);
and U10040 (N_10040,N_9094,N_5481);
or U10041 (N_10041,N_8007,N_6220);
or U10042 (N_10042,N_8636,N_5861);
or U10043 (N_10043,N_7575,N_6626);
nor U10044 (N_10044,N_7854,N_5403);
or U10045 (N_10045,N_6992,N_6410);
nor U10046 (N_10046,N_9073,N_5328);
or U10047 (N_10047,N_6875,N_7075);
nand U10048 (N_10048,N_6070,N_9514);
nor U10049 (N_10049,N_7582,N_8100);
nor U10050 (N_10050,N_9936,N_7637);
and U10051 (N_10051,N_5813,N_6495);
nand U10052 (N_10052,N_8312,N_8334);
nand U10053 (N_10053,N_8974,N_9497);
and U10054 (N_10054,N_9799,N_7319);
and U10055 (N_10055,N_6168,N_8036);
nand U10056 (N_10056,N_7674,N_5517);
and U10057 (N_10057,N_8500,N_8293);
nor U10058 (N_10058,N_5817,N_7190);
nand U10059 (N_10059,N_9009,N_7043);
and U10060 (N_10060,N_7783,N_6316);
or U10061 (N_10061,N_5102,N_6384);
or U10062 (N_10062,N_5784,N_6972);
nor U10063 (N_10063,N_8801,N_9285);
and U10064 (N_10064,N_8548,N_7911);
nand U10065 (N_10065,N_5225,N_5362);
nand U10066 (N_10066,N_6068,N_6228);
nand U10067 (N_10067,N_5027,N_9640);
nand U10068 (N_10068,N_7327,N_6598);
and U10069 (N_10069,N_7320,N_8797);
nand U10070 (N_10070,N_5448,N_9006);
or U10071 (N_10071,N_5918,N_5878);
and U10072 (N_10072,N_7488,N_5221);
or U10073 (N_10073,N_7232,N_5825);
nor U10074 (N_10074,N_7992,N_7712);
and U10075 (N_10075,N_7818,N_8744);
or U10076 (N_10076,N_8165,N_6386);
and U10077 (N_10077,N_7836,N_7521);
and U10078 (N_10078,N_6245,N_8715);
nor U10079 (N_10079,N_6475,N_5079);
or U10080 (N_10080,N_7690,N_8257);
nor U10081 (N_10081,N_6048,N_5342);
or U10082 (N_10082,N_5895,N_7466);
and U10083 (N_10083,N_5709,N_6981);
nor U10084 (N_10084,N_5153,N_7687);
or U10085 (N_10085,N_6576,N_6574);
or U10086 (N_10086,N_7194,N_6623);
or U10087 (N_10087,N_8783,N_7768);
nand U10088 (N_10088,N_7732,N_9984);
nand U10089 (N_10089,N_8174,N_5267);
nand U10090 (N_10090,N_9616,N_5692);
or U10091 (N_10091,N_5467,N_8458);
and U10092 (N_10092,N_5261,N_8897);
nor U10093 (N_10093,N_6804,N_9717);
and U10094 (N_10094,N_7328,N_5338);
and U10095 (N_10095,N_6873,N_5899);
or U10096 (N_10096,N_6312,N_5541);
and U10097 (N_10097,N_7868,N_7632);
and U10098 (N_10098,N_5869,N_9284);
or U10099 (N_10099,N_7760,N_8731);
and U10100 (N_10100,N_6140,N_5281);
nor U10101 (N_10101,N_6884,N_8289);
xnor U10102 (N_10102,N_5625,N_8241);
nor U10103 (N_10103,N_7014,N_7344);
nand U10104 (N_10104,N_8964,N_8973);
and U10105 (N_10105,N_7655,N_6369);
nor U10106 (N_10106,N_6066,N_5669);
or U10107 (N_10107,N_7299,N_9821);
or U10108 (N_10108,N_6802,N_7880);
nor U10109 (N_10109,N_7079,N_9422);
xor U10110 (N_10110,N_7937,N_7929);
and U10111 (N_10111,N_6178,N_9098);
nor U10112 (N_10112,N_6990,N_7173);
or U10113 (N_10113,N_7138,N_9360);
or U10114 (N_10114,N_6169,N_6497);
nand U10115 (N_10115,N_5030,N_8629);
or U10116 (N_10116,N_8613,N_9415);
and U10117 (N_10117,N_6822,N_5904);
nor U10118 (N_10118,N_7012,N_8196);
nand U10119 (N_10119,N_7119,N_8489);
nand U10120 (N_10120,N_7811,N_9917);
or U10121 (N_10121,N_6252,N_8518);
or U10122 (N_10122,N_5694,N_7996);
nand U10123 (N_10123,N_8941,N_9609);
and U10124 (N_10124,N_6989,N_5851);
or U10125 (N_10125,N_6439,N_9001);
or U10126 (N_10126,N_9206,N_5363);
or U10127 (N_10127,N_9535,N_5955);
nand U10128 (N_10128,N_5173,N_9395);
nand U10129 (N_10129,N_5288,N_9639);
nor U10130 (N_10130,N_9875,N_6665);
nand U10131 (N_10131,N_9448,N_9199);
nand U10132 (N_10132,N_8140,N_9100);
nor U10133 (N_10133,N_9011,N_7539);
nand U10134 (N_10134,N_5305,N_9755);
and U10135 (N_10135,N_6501,N_8741);
and U10136 (N_10136,N_8769,N_8528);
nand U10137 (N_10137,N_6028,N_5736);
and U10138 (N_10138,N_9081,N_7603);
or U10139 (N_10139,N_7882,N_6174);
nand U10140 (N_10140,N_8979,N_5648);
and U10141 (N_10141,N_5907,N_9179);
or U10142 (N_10142,N_5249,N_9087);
nor U10143 (N_10143,N_6340,N_6724);
or U10144 (N_10144,N_5280,N_9028);
and U10145 (N_10145,N_6812,N_6985);
and U10146 (N_10146,N_7865,N_6108);
nor U10147 (N_10147,N_9870,N_7004);
nand U10148 (N_10148,N_9683,N_5737);
or U10149 (N_10149,N_9680,N_9931);
nand U10150 (N_10150,N_8809,N_6322);
nand U10151 (N_10151,N_8496,N_7966);
and U10152 (N_10152,N_6117,N_5580);
and U10153 (N_10153,N_6717,N_5519);
and U10154 (N_10154,N_9981,N_7089);
nand U10155 (N_10155,N_7736,N_9730);
nor U10156 (N_10156,N_8480,N_7060);
nand U10157 (N_10157,N_9817,N_9298);
nand U10158 (N_10158,N_8089,N_6942);
or U10159 (N_10159,N_9871,N_7005);
xor U10160 (N_10160,N_9015,N_5191);
nor U10161 (N_10161,N_6686,N_7351);
nand U10162 (N_10162,N_8343,N_8142);
and U10163 (N_10163,N_5085,N_9439);
xor U10164 (N_10164,N_5087,N_6930);
or U10165 (N_10165,N_7955,N_6295);
nor U10166 (N_10166,N_8909,N_8333);
or U10167 (N_10167,N_6935,N_6622);
nand U10168 (N_10168,N_8191,N_5482);
or U10169 (N_10169,N_7963,N_8283);
nand U10170 (N_10170,N_6522,N_8713);
and U10171 (N_10171,N_6748,N_9033);
nor U10172 (N_10172,N_5126,N_8350);
and U10173 (N_10173,N_7162,N_5682);
or U10174 (N_10174,N_8073,N_8701);
or U10175 (N_10175,N_5368,N_9761);
or U10176 (N_10176,N_9092,N_9280);
or U10177 (N_10177,N_9058,N_7183);
nand U10178 (N_10178,N_9550,N_7893);
nor U10179 (N_10179,N_7777,N_8433);
or U10180 (N_10180,N_8252,N_7660);
nand U10181 (N_10181,N_7991,N_5593);
nor U10182 (N_10182,N_6399,N_7569);
or U10183 (N_10183,N_7873,N_7186);
nand U10184 (N_10184,N_5074,N_8234);
and U10185 (N_10185,N_9308,N_7830);
nand U10186 (N_10186,N_9432,N_5314);
nand U10187 (N_10187,N_9590,N_7791);
and U10188 (N_10188,N_9892,N_9608);
nor U10189 (N_10189,N_5166,N_6740);
nand U10190 (N_10190,N_9247,N_6703);
or U10191 (N_10191,N_7470,N_9797);
or U10192 (N_10192,N_7276,N_5549);
xnor U10193 (N_10193,N_9249,N_7944);
nand U10194 (N_10194,N_7504,N_7922);
and U10195 (N_10195,N_7512,N_7058);
or U10196 (N_10196,N_6283,N_8088);
or U10197 (N_10197,N_6530,N_6808);
nor U10198 (N_10198,N_5840,N_5800);
or U10199 (N_10199,N_8855,N_9014);
or U10200 (N_10200,N_9412,N_8201);
nor U10201 (N_10201,N_6547,N_7615);
and U10202 (N_10202,N_6357,N_8995);
nand U10203 (N_10203,N_6754,N_7832);
or U10204 (N_10204,N_6799,N_5697);
nor U10205 (N_10205,N_6398,N_6190);
or U10206 (N_10206,N_5954,N_5206);
nor U10207 (N_10207,N_9044,N_9474);
nor U10208 (N_10208,N_9966,N_6055);
nand U10209 (N_10209,N_6089,N_6741);
or U10210 (N_10210,N_5354,N_6466);
nand U10211 (N_10211,N_8661,N_8802);
and U10212 (N_10212,N_9752,N_5108);
and U10213 (N_10213,N_8609,N_7510);
or U10214 (N_10214,N_6215,N_8888);
nor U10215 (N_10215,N_6969,N_9907);
or U10216 (N_10216,N_5612,N_9372);
nor U10217 (N_10217,N_6033,N_7120);
nor U10218 (N_10218,N_9193,N_7477);
nand U10219 (N_10219,N_5139,N_7487);
nand U10220 (N_10220,N_8706,N_9473);
or U10221 (N_10221,N_7407,N_7041);
nor U10222 (N_10222,N_9604,N_5405);
nand U10223 (N_10223,N_8811,N_7750);
nand U10224 (N_10224,N_9065,N_9130);
and U10225 (N_10225,N_7146,N_9690);
and U10226 (N_10226,N_9406,N_9477);
and U10227 (N_10227,N_6424,N_7494);
or U10228 (N_10228,N_6241,N_8085);
nand U10229 (N_10229,N_9376,N_5491);
nand U10230 (N_10230,N_5243,N_5932);
or U10231 (N_10231,N_5708,N_9218);
nor U10232 (N_10232,N_8898,N_7142);
nand U10233 (N_10233,N_6577,N_9325);
nor U10234 (N_10234,N_8253,N_9460);
nand U10235 (N_10235,N_8491,N_9154);
and U10236 (N_10236,N_7782,N_8206);
xnor U10237 (N_10237,N_6402,N_7280);
nand U10238 (N_10238,N_7206,N_9196);
nand U10239 (N_10239,N_6155,N_7897);
and U10240 (N_10240,N_8880,N_8263);
nand U10241 (N_10241,N_6032,N_6918);
and U10242 (N_10242,N_8937,N_5691);
nand U10243 (N_10243,N_9289,N_5856);
nand U10244 (N_10244,N_5925,N_8294);
nor U10245 (N_10245,N_9855,N_5107);
nor U10246 (N_10246,N_5487,N_9768);
nor U10247 (N_10247,N_9270,N_7353);
or U10248 (N_10248,N_6680,N_7326);
nor U10249 (N_10249,N_6517,N_7890);
or U10250 (N_10250,N_7825,N_9296);
nand U10251 (N_10251,N_8127,N_6655);
nand U10252 (N_10252,N_8649,N_9784);
nor U10253 (N_10253,N_9568,N_6856);
and U10254 (N_10254,N_5723,N_7063);
or U10255 (N_10255,N_8817,N_9831);
or U10256 (N_10256,N_7331,N_8396);
nand U10257 (N_10257,N_7032,N_7971);
nor U10258 (N_10258,N_8700,N_7808);
nor U10259 (N_10259,N_5742,N_6756);
nand U10260 (N_10260,N_8389,N_6209);
or U10261 (N_10261,N_6051,N_5385);
or U10262 (N_10262,N_8120,N_9378);
and U10263 (N_10263,N_6759,N_9949);
and U10264 (N_10264,N_5988,N_9124);
nor U10265 (N_10265,N_9633,N_5607);
nor U10266 (N_10266,N_8187,N_7928);
or U10267 (N_10267,N_8482,N_7383);
nor U10268 (N_10268,N_9311,N_6940);
nor U10269 (N_10269,N_7303,N_9807);
nand U10270 (N_10270,N_6382,N_5661);
nor U10271 (N_10271,N_7531,N_5237);
and U10272 (N_10272,N_8235,N_7391);
nand U10273 (N_10273,N_7775,N_5485);
nor U10274 (N_10274,N_6778,N_7046);
nand U10275 (N_10275,N_7578,N_8074);
or U10276 (N_10276,N_7564,N_9565);
and U10277 (N_10277,N_9408,N_9042);
nand U10278 (N_10278,N_5406,N_8168);
xnor U10279 (N_10279,N_5984,N_9695);
or U10280 (N_10280,N_6641,N_5726);
or U10281 (N_10281,N_5091,N_8524);
nand U10282 (N_10282,N_9182,N_5934);
and U10283 (N_10283,N_7133,N_5431);
or U10284 (N_10284,N_6355,N_7434);
nor U10285 (N_10285,N_7608,N_8554);
nor U10286 (N_10286,N_5823,N_7015);
nor U10287 (N_10287,N_6869,N_6198);
or U10288 (N_10288,N_5914,N_8010);
nor U10289 (N_10289,N_8986,N_6512);
nor U10290 (N_10290,N_8767,N_9399);
or U10291 (N_10291,N_7695,N_7228);
or U10292 (N_10292,N_8822,N_5178);
nor U10293 (N_10293,N_8208,N_9783);
nor U10294 (N_10294,N_7287,N_5452);
and U10295 (N_10295,N_7392,N_5009);
nor U10296 (N_10296,N_6119,N_6005);
nor U10297 (N_10297,N_8938,N_6462);
and U10298 (N_10298,N_6762,N_6329);
nor U10299 (N_10299,N_6365,N_7964);
nor U10300 (N_10300,N_9923,N_8907);
nand U10301 (N_10301,N_5170,N_9209);
and U10302 (N_10302,N_9932,N_6154);
nor U10303 (N_10303,N_8096,N_9455);
nand U10304 (N_10304,N_6902,N_9970);
nor U10305 (N_10305,N_8793,N_7686);
nor U10306 (N_10306,N_9660,N_5804);
and U10307 (N_10307,N_7744,N_8572);
or U10308 (N_10308,N_8404,N_9269);
or U10309 (N_10309,N_8835,N_5443);
and U10310 (N_10310,N_6991,N_6385);
and U10311 (N_10311,N_6328,N_7681);
nor U10312 (N_10312,N_8550,N_5215);
or U10313 (N_10313,N_5436,N_9177);
nor U10314 (N_10314,N_7264,N_8968);
nor U10315 (N_10315,N_5688,N_6162);
nand U10316 (N_10316,N_5437,N_6818);
or U10317 (N_10317,N_8225,N_7553);
nand U10318 (N_10318,N_5290,N_8734);
and U10319 (N_10319,N_6960,N_5599);
nand U10320 (N_10320,N_9993,N_5507);
nor U10321 (N_10321,N_9885,N_9111);
and U10322 (N_10322,N_5883,N_9845);
or U10323 (N_10323,N_9818,N_6306);
nand U10324 (N_10324,N_5655,N_5829);
or U10325 (N_10325,N_9620,N_7505);
and U10326 (N_10326,N_8736,N_5421);
nand U10327 (N_10327,N_8094,N_6634);
nand U10328 (N_10328,N_7221,N_9089);
and U10329 (N_10329,N_5670,N_5802);
nand U10330 (N_10330,N_6900,N_9617);
nand U10331 (N_10331,N_9928,N_9531);
nor U10332 (N_10332,N_8538,N_6927);
and U10333 (N_10333,N_5967,N_5004);
and U10334 (N_10334,N_6753,N_9034);
nand U10335 (N_10335,N_7038,N_9418);
and U10336 (N_10336,N_7597,N_8141);
nand U10337 (N_10337,N_6079,N_8228);
and U10338 (N_10338,N_5204,N_5223);
nor U10339 (N_10339,N_6815,N_6107);
nor U10340 (N_10340,N_6760,N_5733);
and U10341 (N_10341,N_9409,N_6725);
and U10342 (N_10342,N_8400,N_8020);
or U10343 (N_10343,N_6370,N_8425);
or U10344 (N_10344,N_7499,N_6105);
and U10345 (N_10345,N_9461,N_5913);
nor U10346 (N_10346,N_8005,N_6862);
or U10347 (N_10347,N_8434,N_8521);
or U10348 (N_10348,N_6243,N_5378);
or U10349 (N_10349,N_6677,N_6944);
and U10350 (N_10350,N_8446,N_5930);
and U10351 (N_10351,N_9904,N_6941);
or U10352 (N_10352,N_8340,N_5372);
nand U10353 (N_10353,N_5537,N_8765);
or U10354 (N_10354,N_5623,N_7789);
nor U10355 (N_10355,N_8505,N_5344);
and U10356 (N_10356,N_7563,N_6579);
and U10357 (N_10357,N_6091,N_8657);
or U10358 (N_10358,N_5458,N_7551);
nor U10359 (N_10359,N_5573,N_9500);
nor U10360 (N_10360,N_6722,N_9290);
nor U10361 (N_10361,N_9693,N_6524);
nor U10362 (N_10362,N_8581,N_5209);
and U10363 (N_10363,N_9364,N_9563);
or U10364 (N_10364,N_9392,N_7692);
xor U10365 (N_10365,N_5945,N_9570);
xnor U10366 (N_10366,N_9521,N_9612);
and U10367 (N_10367,N_9989,N_7081);
nor U10368 (N_10368,N_7653,N_9753);
xor U10369 (N_10369,N_8121,N_7495);
xor U10370 (N_10370,N_8685,N_8213);
or U10371 (N_10371,N_8236,N_7869);
and U10372 (N_10372,N_6003,N_8601);
nor U10373 (N_10373,N_9317,N_9494);
and U10374 (N_10374,N_7355,N_7127);
nor U10375 (N_10375,N_9779,N_9594);
and U10376 (N_10376,N_9230,N_6310);
and U10377 (N_10377,N_8081,N_9839);
and U10378 (N_10378,N_6781,N_8692);
or U10379 (N_10379,N_6397,N_7364);
nand U10380 (N_10380,N_9012,N_5339);
or U10381 (N_10381,N_7570,N_8615);
or U10382 (N_10382,N_6840,N_9496);
or U10383 (N_10383,N_6225,N_6176);
and U10384 (N_10384,N_7057,N_8525);
nor U10385 (N_10385,N_7565,N_5167);
and U10386 (N_10386,N_7255,N_5712);
nor U10387 (N_10387,N_5316,N_7612);
and U10388 (N_10388,N_9048,N_5202);
nor U10389 (N_10389,N_9654,N_9067);
and U10390 (N_10390,N_5543,N_7034);
or U10391 (N_10391,N_8090,N_8896);
xnor U10392 (N_10392,N_5674,N_9687);
or U10393 (N_10393,N_5250,N_9518);
or U10394 (N_10394,N_6931,N_7150);
and U10395 (N_10395,N_7594,N_9980);
nand U10396 (N_10396,N_8212,N_9651);
nand U10397 (N_10397,N_7008,N_8607);
nor U10398 (N_10398,N_8456,N_8803);
or U10399 (N_10399,N_6094,N_9366);
xor U10400 (N_10400,N_6060,N_5787);
or U10401 (N_10401,N_8533,N_9635);
and U10402 (N_10402,N_6823,N_9527);
or U10403 (N_10403,N_9611,N_7288);
and U10404 (N_10404,N_9204,N_9056);
nor U10405 (N_10405,N_6463,N_9419);
nand U10406 (N_10406,N_8031,N_9624);
or U10407 (N_10407,N_7892,N_5024);
and U10408 (N_10408,N_9190,N_8998);
nor U10409 (N_10409,N_9004,N_9168);
or U10410 (N_10410,N_8232,N_7658);
or U10411 (N_10411,N_5123,N_8423);
or U10412 (N_10412,N_5425,N_5715);
and U10413 (N_10413,N_7593,N_8933);
or U10414 (N_10414,N_5763,N_5045);
and U10415 (N_10415,N_5680,N_7630);
nor U10416 (N_10416,N_5997,N_8368);
nand U10417 (N_10417,N_5631,N_6820);
and U10418 (N_10418,N_8985,N_9127);
nand U10419 (N_10419,N_8623,N_8418);
or U10420 (N_10420,N_9805,N_6257);
and U10421 (N_10421,N_8844,N_8291);
xor U10422 (N_10422,N_5253,N_6288);
or U10423 (N_10423,N_9742,N_5626);
nor U10424 (N_10424,N_5138,N_7780);
or U10425 (N_10425,N_6897,N_5843);
nor U10426 (N_10426,N_5810,N_8045);
nor U10427 (N_10427,N_8429,N_6115);
nand U10428 (N_10428,N_8409,N_9913);
and U10429 (N_10429,N_7755,N_9646);
and U10430 (N_10430,N_6083,N_6883);
nor U10431 (N_10431,N_8380,N_5968);
and U10432 (N_10432,N_9522,N_5315);
nor U10433 (N_10433,N_6745,N_7246);
nor U10434 (N_10434,N_5903,N_8112);
or U10435 (N_10435,N_8574,N_5970);
and U10436 (N_10436,N_6541,N_9454);
and U10437 (N_10437,N_8044,N_7624);
nor U10438 (N_10438,N_5216,N_6388);
and U10439 (N_10439,N_5873,N_8067);
nand U10440 (N_10440,N_6838,N_5113);
nor U10441 (N_10441,N_6562,N_5986);
or U10442 (N_10442,N_8954,N_7356);
or U10443 (N_10443,N_5322,N_6346);
nand U10444 (N_10444,N_8776,N_8475);
nor U10445 (N_10445,N_6307,N_5381);
or U10446 (N_10446,N_7231,N_8925);
and U10447 (N_10447,N_5001,N_6810);
and U10448 (N_10448,N_9947,N_8443);
nor U10449 (N_10449,N_8726,N_6583);
nand U10450 (N_10450,N_7380,N_7899);
and U10451 (N_10451,N_5335,N_9903);
nand U10452 (N_10452,N_5211,N_6956);
nand U10453 (N_10453,N_6984,N_6657);
or U10454 (N_10454,N_9211,N_7958);
or U10455 (N_10455,N_5190,N_6607);
or U10456 (N_10456,N_5373,N_9569);
nor U10457 (N_10457,N_5707,N_9827);
and U10458 (N_10458,N_5801,N_5564);
or U10459 (N_10459,N_5484,N_8481);
nor U10460 (N_10460,N_6996,N_5361);
and U10461 (N_10461,N_8021,N_6479);
or U10462 (N_10462,N_6337,N_8996);
nor U10463 (N_10463,N_8483,N_9720);
nand U10464 (N_10464,N_6082,N_5794);
nand U10465 (N_10465,N_8796,N_7396);
and U10466 (N_10466,N_7661,N_7985);
nor U10467 (N_10467,N_9800,N_8411);
and U10468 (N_10468,N_7511,N_6676);
and U10469 (N_10469,N_9748,N_9374);
and U10470 (N_10470,N_6166,N_8054);
nand U10471 (N_10471,N_7822,N_7562);
or U10472 (N_10472,N_7731,N_7175);
and U10473 (N_10473,N_5673,N_8867);
nor U10474 (N_10474,N_9954,N_7455);
nor U10475 (N_10475,N_6516,N_7095);
nand U10476 (N_10476,N_5889,N_8999);
nand U10477 (N_10477,N_9234,N_7091);
nor U10478 (N_10478,N_5795,N_8226);
nor U10479 (N_10479,N_8000,N_8808);
and U10480 (N_10480,N_7045,N_5195);
and U10481 (N_10481,N_9670,N_5524);
nor U10482 (N_10482,N_5128,N_5525);
or U10483 (N_10483,N_8714,N_7728);
and U10484 (N_10484,N_6567,N_6705);
nand U10485 (N_10485,N_6485,N_9759);
or U10486 (N_10486,N_6581,N_8420);
nand U10487 (N_10487,N_9967,N_9711);
or U10488 (N_10488,N_6792,N_5242);
and U10489 (N_10489,N_7121,N_8514);
nor U10490 (N_10490,N_8264,N_7529);
and U10491 (N_10491,N_5920,N_9872);
nand U10492 (N_10492,N_6711,N_6330);
and U10493 (N_10493,N_5656,N_6660);
nor U10494 (N_10494,N_9429,N_8588);
and U10495 (N_10495,N_8503,N_9769);
nor U10496 (N_10496,N_7476,N_6945);
nor U10497 (N_10497,N_5157,N_6120);
nand U10498 (N_10498,N_7387,N_6478);
or U10499 (N_10499,N_8686,N_9629);
nor U10500 (N_10500,N_6112,N_9754);
nand U10501 (N_10501,N_7253,N_7667);
xor U10502 (N_10502,N_6749,N_5793);
nor U10503 (N_10503,N_6208,N_8957);
nand U10504 (N_10504,N_7086,N_6560);
xor U10505 (N_10505,N_9834,N_7849);
or U10506 (N_10506,N_5016,N_5533);
nand U10507 (N_10507,N_9331,N_9836);
and U10508 (N_10508,N_8321,N_6319);
nor U10509 (N_10509,N_8494,N_9139);
nor U10510 (N_10510,N_5518,N_6716);
or U10511 (N_10511,N_7053,N_9975);
and U10512 (N_10512,N_7266,N_8600);
and U10513 (N_10513,N_5246,N_7573);
or U10514 (N_10514,N_7639,N_5463);
or U10515 (N_10515,N_6582,N_8024);
or U10516 (N_10516,N_8113,N_6039);
and U10517 (N_10517,N_8091,N_9210);
or U10518 (N_10518,N_9459,N_7109);
or U10519 (N_10519,N_9703,N_8377);
or U10520 (N_10520,N_9652,N_5069);
nand U10521 (N_10521,N_7341,N_9507);
nand U10522 (N_10522,N_9462,N_7177);
nor U10523 (N_10523,N_7337,N_5247);
and U10524 (N_10524,N_5578,N_9320);
nor U10525 (N_10525,N_7238,N_5606);
and U10526 (N_10526,N_9143,N_6729);
or U10527 (N_10527,N_8754,N_7277);
nor U10528 (N_10528,N_5460,N_6761);
and U10529 (N_10529,N_6798,N_9544);
and U10530 (N_10530,N_7815,N_9344);
and U10531 (N_10531,N_8328,N_6459);
nor U10532 (N_10532,N_7727,N_6496);
nand U10533 (N_10533,N_6709,N_5293);
or U10534 (N_10534,N_9697,N_7807);
nand U10535 (N_10535,N_6167,N_7968);
nand U10536 (N_10536,N_7098,N_5594);
and U10537 (N_10537,N_7203,N_6223);
or U10538 (N_10538,N_8002,N_5129);
or U10539 (N_10539,N_5395,N_9428);
and U10540 (N_10540,N_7691,N_5956);
nand U10541 (N_10541,N_5676,N_8852);
nand U10542 (N_10542,N_8819,N_8367);
nor U10543 (N_10543,N_9005,N_6194);
or U10544 (N_10544,N_8079,N_7472);
nand U10545 (N_10545,N_8510,N_9896);
nand U10546 (N_10546,N_6777,N_5364);
or U10547 (N_10547,N_5297,N_6564);
or U10548 (N_10548,N_9659,N_7805);
and U10549 (N_10549,N_8856,N_8272);
nand U10550 (N_10550,N_9804,N_8484);
or U10551 (N_10551,N_5398,N_6314);
or U10552 (N_10552,N_9281,N_8477);
and U10553 (N_10553,N_5587,N_9032);
or U10554 (N_10554,N_7066,N_9795);
xnor U10555 (N_10555,N_8781,N_6536);
and U10556 (N_10556,N_6229,N_8189);
nand U10557 (N_10557,N_6876,N_6266);
nor U10558 (N_10558,N_7093,N_8199);
or U10559 (N_10559,N_8637,N_9911);
nor U10560 (N_10560,N_7640,N_8705);
nand U10561 (N_10561,N_8317,N_7261);
nor U10562 (N_10562,N_6071,N_8237);
nand U10563 (N_10563,N_9943,N_7821);
and U10564 (N_10564,N_6246,N_5289);
or U10565 (N_10565,N_6250,N_8627);
nor U10566 (N_10566,N_7709,N_9901);
and U10567 (N_10567,N_5393,N_6401);
nand U10568 (N_10568,N_6011,N_7871);
and U10569 (N_10569,N_6587,N_5837);
nand U10570 (N_10570,N_6791,N_9369);
and U10571 (N_10571,N_7838,N_7983);
nand U10572 (N_10572,N_7743,N_8748);
or U10573 (N_10573,N_8442,N_5511);
and U10574 (N_10574,N_7201,N_8315);
or U10575 (N_10575,N_9156,N_7389);
nand U10576 (N_10576,N_7688,N_7544);
nor U10577 (N_10577,N_7406,N_5008);
nand U10578 (N_10578,N_5271,N_6787);
and U10579 (N_10579,N_8788,N_9365);
nand U10580 (N_10580,N_6837,N_6553);
and U10581 (N_10581,N_7101,N_8492);
nor U10582 (N_10582,N_6903,N_8919);
and U10583 (N_10583,N_6673,N_5468);
nor U10584 (N_10584,N_5589,N_5099);
nor U10585 (N_10585,N_8892,N_7258);
nor U10586 (N_10586,N_8375,N_6020);
or U10587 (N_10587,N_8826,N_9446);
nor U10588 (N_10588,N_9303,N_6796);
nor U10589 (N_10589,N_7701,N_9722);
nor U10590 (N_10590,N_5081,N_7614);
or U10591 (N_10591,N_7178,N_5332);
and U10592 (N_10592,N_8466,N_9996);
or U10593 (N_10593,N_7016,N_8812);
and U10594 (N_10594,N_9436,N_9942);
nand U10595 (N_10595,N_7433,N_6177);
nor U10596 (N_10596,N_7957,N_5958);
nor U10597 (N_10597,N_6612,N_8287);
or U10598 (N_10598,N_9760,N_7532);
nor U10599 (N_10599,N_8886,N_6784);
nand U10600 (N_10600,N_6616,N_7316);
or U10601 (N_10601,N_7459,N_9848);
and U10602 (N_10602,N_6647,N_5336);
and U10603 (N_10603,N_7309,N_7626);
nor U10604 (N_10604,N_9701,N_5514);
and U10605 (N_10605,N_9939,N_7618);
nand U10606 (N_10606,N_5959,N_5356);
nor U10607 (N_10607,N_8460,N_6009);
and U10608 (N_10608,N_7215,N_8388);
and U10609 (N_10609,N_8144,N_8318);
nor U10610 (N_10610,N_9623,N_8137);
or U10611 (N_10611,N_8238,N_8129);
nand U10612 (N_10612,N_5453,N_5893);
nor U10613 (N_10613,N_8260,N_6487);
nor U10614 (N_10614,N_5983,N_9010);
and U10615 (N_10615,N_6062,N_5026);
or U10616 (N_10616,N_7620,N_8628);
nand U10617 (N_10617,N_8761,N_5796);
and U10618 (N_10618,N_7621,N_6449);
nor U10619 (N_10619,N_7642,N_6262);
nand U10620 (N_10620,N_7414,N_5422);
nor U10621 (N_10621,N_9916,N_6299);
nand U10622 (N_10622,N_8504,N_7021);
and U10623 (N_10623,N_6438,N_9080);
or U10624 (N_10624,N_7410,N_9641);
nor U10625 (N_10625,N_9708,N_6444);
nand U10626 (N_10626,N_8772,N_8952);
nand U10627 (N_10627,N_5963,N_6110);
and U10628 (N_10628,N_8960,N_9564);
nor U10629 (N_10629,N_5960,N_9336);
and U10630 (N_10630,N_5056,N_9340);
or U10631 (N_10631,N_9467,N_7833);
and U10632 (N_10632,N_5132,N_5944);
nor U10633 (N_10633,N_8626,N_7935);
or U10634 (N_10634,N_7589,N_6016);
xnor U10635 (N_10635,N_9053,N_7155);
and U10636 (N_10636,N_9764,N_9472);
nand U10637 (N_10637,N_7244,N_8641);
nor U10638 (N_10638,N_8223,N_8565);
or U10639 (N_10639,N_9601,N_6008);
and U10640 (N_10640,N_5972,N_8766);
or U10641 (N_10641,N_8103,N_9707);
nand U10642 (N_10642,N_8192,N_8991);
and U10643 (N_10643,N_9229,N_7130);
nor U10644 (N_10644,N_5815,N_6603);
and U10645 (N_10645,N_7068,N_5042);
nand U10646 (N_10646,N_8487,N_5321);
and U10647 (N_10647,N_5111,N_6906);
and U10648 (N_10648,N_7954,N_7656);
and U10649 (N_10649,N_6650,N_9468);
and U10650 (N_10650,N_5179,N_8678);
or U10651 (N_10651,N_9791,N_6864);
nand U10652 (N_10652,N_5877,N_5124);
nor U10653 (N_10653,N_8281,N_5975);
and U10654 (N_10654,N_8681,N_8825);
or U10655 (N_10655,N_8947,N_9686);
and U10656 (N_10656,N_7125,N_8502);
nand U10657 (N_10657,N_9385,N_6293);
nand U10658 (N_10658,N_5619,N_7530);
nor U10659 (N_10659,N_8617,N_6922);
nor U10660 (N_10660,N_8977,N_6132);
or U10661 (N_10661,N_7105,N_8535);
and U10662 (N_10662,N_5554,N_9337);
and U10663 (N_10663,N_7623,N_6152);
and U10664 (N_10664,N_5105,N_8859);
and U10665 (N_10665,N_8945,N_8038);
and U10666 (N_10666,N_8961,N_7395);
and U10667 (N_10667,N_8256,N_6458);
and U10668 (N_10668,N_7605,N_7538);
nand U10669 (N_10669,N_7315,N_6004);
and U10670 (N_10670,N_6102,N_6075);
nor U10671 (N_10671,N_6965,N_7795);
nor U10672 (N_10672,N_5038,N_6706);
nand U10673 (N_10673,N_6320,N_6362);
or U10674 (N_10674,N_5394,N_8589);
or U10675 (N_10675,N_6372,N_8622);
or U10676 (N_10676,N_8575,N_7859);
nand U10677 (N_10677,N_6042,N_7219);
or U10678 (N_10678,N_5254,N_7307);
and U10679 (N_10679,N_7367,N_7934);
and U10680 (N_10680,N_6443,N_8558);
or U10681 (N_10681,N_9255,N_6125);
nor U10682 (N_10682,N_8479,N_7738);
and U10683 (N_10683,N_7054,N_9109);
or U10684 (N_10684,N_6889,N_7143);
and U10685 (N_10685,N_7463,N_8325);
nor U10686 (N_10686,N_9346,N_6271);
or U10687 (N_10687,N_5275,N_6515);
and U10688 (N_10688,N_5325,N_7349);
and U10689 (N_10689,N_8560,N_7814);
nand U10690 (N_10690,N_5531,N_7607);
nand U10691 (N_10691,N_5901,N_5755);
nand U10692 (N_10692,N_5808,N_8935);
and U10693 (N_10693,N_8393,N_5265);
nand U10694 (N_10694,N_5788,N_7598);
or U10695 (N_10695,N_6994,N_8905);
nand U10696 (N_10696,N_8331,N_7740);
and U10697 (N_10697,N_9968,N_7436);
nand U10698 (N_10698,N_9843,N_9756);
or U10699 (N_10699,N_6723,N_7776);
and U10700 (N_10700,N_7225,N_6498);
nand U10701 (N_10701,N_9673,N_9741);
nand U10702 (N_10702,N_5302,N_8583);
and U10703 (N_10703,N_9107,N_6636);
or U10704 (N_10704,N_6029,N_6109);
or U10705 (N_10705,N_5866,N_5186);
nand U10706 (N_10706,N_9200,N_9016);
and U10707 (N_10707,N_7450,N_5860);
and U10708 (N_10708,N_7431,N_5212);
or U10709 (N_10709,N_8540,N_8724);
or U10710 (N_10710,N_5743,N_6646);
or U10711 (N_10711,N_9902,N_6139);
xor U10712 (N_10712,N_6239,N_8753);
or U10713 (N_10713,N_5822,N_7198);
nand U10714 (N_10714,N_6216,N_6332);
nand U10715 (N_10715,N_5284,N_9426);
or U10716 (N_10716,N_7745,N_5327);
nand U10717 (N_10717,N_8777,N_7065);
and U10718 (N_10718,N_8774,N_6069);
nand U10719 (N_10719,N_5054,N_5703);
or U10720 (N_10720,N_5735,N_8449);
or U10721 (N_10721,N_6254,N_6453);
and U10722 (N_10722,N_9566,N_8914);
and U10723 (N_10723,N_8578,N_6834);
and U10724 (N_10724,N_8527,N_7154);
nor U10725 (N_10725,N_5188,N_5329);
nand U10726 (N_10726,N_6859,N_5521);
and U10727 (N_10727,N_5234,N_5862);
and U10728 (N_10728,N_9705,N_6899);
nand U10729 (N_10729,N_5657,N_5789);
nand U10730 (N_10730,N_6743,N_5664);
or U10731 (N_10731,N_7234,N_8182);
or U10732 (N_10732,N_6788,N_6057);
and U10733 (N_10733,N_6696,N_8546);
or U10734 (N_10734,N_6149,N_9861);
nand U10735 (N_10735,N_6012,N_7300);
nor U10736 (N_10736,N_5017,N_6970);
nor U10737 (N_10737,N_7716,N_6488);
nand U10738 (N_10738,N_7987,N_6667);
or U10739 (N_10739,N_7566,N_5390);
or U10740 (N_10740,N_7896,N_6908);
and U10741 (N_10741,N_8545,N_9508);
and U10742 (N_10742,N_7047,N_5110);
nand U10743 (N_10743,N_7696,N_5706);
nor U10744 (N_10744,N_7842,N_5546);
or U10745 (N_10745,N_7295,N_5434);
or U10746 (N_10746,N_6364,N_6024);
nor U10747 (N_10747,N_5240,N_9155);
and U10748 (N_10748,N_7223,N_6923);
and U10749 (N_10749,N_9171,N_7943);
and U10750 (N_10750,N_7972,N_8522);
nor U10751 (N_10751,N_6675,N_9960);
xor U10752 (N_10752,N_5671,N_9077);
or U10753 (N_10753,N_6275,N_8874);
and U10754 (N_10754,N_9489,N_7454);
nand U10755 (N_10755,N_6543,N_8230);
and U10756 (N_10756,N_8278,N_7774);
or U10757 (N_10757,N_5985,N_6211);
and U10758 (N_10758,N_6426,N_9043);
or U10759 (N_10759,N_6993,N_7916);
nor U10760 (N_10760,N_8344,N_5609);
and U10761 (N_10761,N_8051,N_5503);
nor U10762 (N_10762,N_5439,N_5219);
and U10763 (N_10763,N_6826,N_9195);
nor U10764 (N_10764,N_9676,N_5717);
or U10765 (N_10765,N_6833,N_9052);
or U10766 (N_10766,N_5020,N_6545);
nand U10767 (N_10767,N_6986,N_6187);
nand U10768 (N_10768,N_5888,N_7017);
nand U10769 (N_10769,N_7559,N_5312);
and U10770 (N_10770,N_9274,N_7111);
or U10771 (N_10771,N_6565,N_8669);
or U10772 (N_10772,N_5013,N_6074);
or U10773 (N_10773,N_8608,N_6327);
or U10774 (N_10774,N_6835,N_6932);
nor U10775 (N_10775,N_6437,N_8590);
nand U10776 (N_10776,N_6720,N_9275);
nor U10777 (N_10777,N_9039,N_9036);
nand U10778 (N_10778,N_6867,N_9329);
nand U10779 (N_10779,N_8787,N_7181);
nand U10780 (N_10780,N_8427,N_8923);
or U10781 (N_10781,N_6464,N_6195);
nor U10782 (N_10782,N_5785,N_8066);
nand U10783 (N_10783,N_5811,N_5605);
and U10784 (N_10784,N_6702,N_7191);
nand U10785 (N_10785,N_5198,N_7471);
nor U10786 (N_10786,N_5300,N_8004);
and U10787 (N_10787,N_5165,N_6237);
nand U10788 (N_10788,N_6095,N_9806);
nand U10789 (N_10789,N_7725,N_7770);
xor U10790 (N_10790,N_5072,N_9763);
and U10791 (N_10791,N_6046,N_7877);
nor U10792 (N_10792,N_6204,N_9537);
nand U10793 (N_10793,N_9951,N_8115);
nor U10794 (N_10794,N_6292,N_9045);
and U10795 (N_10795,N_9307,N_8901);
and U10796 (N_10796,N_9953,N_8338);
or U10797 (N_10797,N_6664,N_7020);
and U10798 (N_10798,N_9158,N_5571);
or U10799 (N_10799,N_7171,N_5003);
and U10800 (N_10800,N_9161,N_8490);
nand U10801 (N_10801,N_8987,N_9491);
and U10802 (N_10802,N_8301,N_5430);
and U10803 (N_10803,N_9776,N_8506);
and U10804 (N_10804,N_9972,N_8851);
and U10805 (N_10805,N_6035,N_5055);
or U10806 (N_10806,N_7489,N_8099);
nor U10807 (N_10807,N_9129,N_8980);
nor U10808 (N_10808,N_7677,N_8474);
nor U10809 (N_10809,N_6390,N_5351);
or U10810 (N_10810,N_6744,N_7816);
or U10811 (N_10811,N_7536,N_6713);
and U10812 (N_10812,N_6549,N_5995);
and U10813 (N_10813,N_9046,N_6409);
nand U10814 (N_10814,N_5266,N_7644);
nor U10815 (N_10815,N_7657,N_9207);
xor U10816 (N_10816,N_7210,N_8059);
nor U10817 (N_10817,N_6103,N_6662);
or U10818 (N_10818,N_8598,N_6831);
xnor U10819 (N_10819,N_5141,N_7915);
nand U10820 (N_10820,N_8139,N_9543);
nor U10821 (N_10821,N_5163,N_7698);
nand U10822 (N_10822,N_8353,N_5562);
and U10823 (N_10823,N_7137,N_6114);
and U10824 (N_10824,N_8737,N_8620);
nor U10825 (N_10825,N_8850,N_8335);
nand U10826 (N_10826,N_8976,N_5565);
nand U10827 (N_10827,N_5174,N_9528);
nor U10828 (N_10828,N_6958,N_9091);
and U10829 (N_10829,N_9287,N_5658);
and U10830 (N_10830,N_9488,N_8352);
or U10831 (N_10831,N_7469,N_8273);
or U10832 (N_10832,N_8512,N_5317);
nor U10833 (N_10833,N_9413,N_9267);
nor U10834 (N_10834,N_8942,N_8895);
and U10835 (N_10835,N_5311,N_7595);
nor U10836 (N_10836,N_7675,N_9746);
or U10837 (N_10837,N_7312,N_5700);
nand U10838 (N_10838,N_9481,N_6494);
nand U10839 (N_10839,N_6142,N_6030);
nor U10840 (N_10840,N_9485,N_6765);
xnor U10841 (N_10841,N_6303,N_6959);
nor U10842 (N_10842,N_9119,N_8062);
nand U10843 (N_10843,N_9820,N_6199);
nor U10844 (N_10844,N_5931,N_6511);
and U10845 (N_10845,N_7747,N_5906);
and U10846 (N_10846,N_7377,N_5196);
or U10847 (N_10847,N_5677,N_7317);
nand U10848 (N_10848,N_5058,N_6127);
and U10849 (N_10849,N_8943,N_9578);
nor U10850 (N_10850,N_9781,N_9495);
or U10851 (N_10851,N_5433,N_9808);
nand U10852 (N_10852,N_7817,N_7883);
and U10853 (N_10853,N_8320,N_6080);
nand U10854 (N_10854,N_5454,N_5644);
nor U10855 (N_10855,N_5545,N_8329);
nor U10856 (N_10856,N_9580,N_5665);
nor U10857 (N_10857,N_8014,N_8276);
nand U10858 (N_10858,N_5057,N_5049);
or U10859 (N_10859,N_5424,N_9121);
or U10860 (N_10860,N_8997,N_9060);
nand U10861 (N_10861,N_9160,N_6186);
nand U10862 (N_10862,N_9097,N_7974);
nor U10863 (N_10863,N_6698,N_8001);
nor U10864 (N_10864,N_6413,N_5078);
nand U10865 (N_10865,N_7085,N_9431);
or U10866 (N_10866,N_5953,N_8571);
and U10867 (N_10867,N_6145,N_7370);
or U10868 (N_10868,N_7853,N_6645);
and U10869 (N_10869,N_6391,N_5548);
and U10870 (N_10870,N_8111,N_7174);
or U10871 (N_10871,N_8310,N_7375);
nor U10872 (N_10872,N_5882,N_8846);
nor U10873 (N_10873,N_7528,N_6383);
nand U10874 (N_10874,N_5529,N_7705);
or U10875 (N_10875,N_7220,N_8936);
nor U10876 (N_10876,N_6769,N_9559);
nand U10877 (N_10877,N_5499,N_9167);
and U10878 (N_10878,N_6258,N_7668);
and U10879 (N_10879,N_8181,N_8780);
and U10880 (N_10880,N_8762,N_6521);
or U10881 (N_10881,N_9440,N_5150);
or U10882 (N_10882,N_9264,N_5905);
nand U10883 (N_10883,N_8648,N_5231);
or U10884 (N_10884,N_8614,N_6934);
nor U10885 (N_10885,N_5180,N_7819);
nand U10886 (N_10886,N_8379,N_9096);
and U10887 (N_10887,N_8163,N_7676);
nand U10888 (N_10888,N_9957,N_5438);
or U10889 (N_10889,N_5750,N_7903);
nor U10890 (N_10890,N_9330,N_5035);
xor U10891 (N_10891,N_6073,N_7664);
and U10892 (N_10892,N_9184,N_8647);
and U10893 (N_10893,N_8718,N_9288);
nor U10894 (N_10894,N_5292,N_9930);
and U10895 (N_10895,N_7646,N_9405);
or U10896 (N_10896,N_6894,N_9596);
and U10897 (N_10897,N_8247,N_5295);
nor U10898 (N_10898,N_7361,N_6321);
xnor U10899 (N_10899,N_8672,N_7110);
nor U10900 (N_10900,N_5282,N_8267);
nor U10901 (N_10901,N_7250,N_9961);
or U10902 (N_10902,N_5943,N_7581);
and U10903 (N_10903,N_6886,N_5268);
nor U10904 (N_10904,N_7306,N_9407);
or U10905 (N_10905,N_8721,N_7281);
nor U10906 (N_10906,N_9268,N_6751);
and U10907 (N_10907,N_8360,N_9021);
nand U10908 (N_10908,N_7988,N_6131);
nand U10909 (N_10909,N_6672,N_9888);
nor U10910 (N_10910,N_9955,N_8249);
or U10911 (N_10911,N_7723,N_8582);
or U10912 (N_10912,N_9476,N_5790);
nor U10913 (N_10913,N_6481,N_5993);
and U10914 (N_10914,N_9064,N_6841);
xor U10915 (N_10915,N_9236,N_6300);
and U10916 (N_10916,N_9194,N_8064);
or U10917 (N_10917,N_9883,N_9974);
and U10918 (N_10918,N_7199,N_6484);
or U10919 (N_10919,N_8770,N_8126);
and U10920 (N_10920,N_8606,N_7461);
and U10921 (N_10921,N_7336,N_7840);
nand U10922 (N_10922,N_8445,N_7586);
nand U10923 (N_10923,N_5029,N_6087);
nor U10924 (N_10924,N_8341,N_7724);
and U10925 (N_10925,N_7243,N_7652);
and U10926 (N_10926,N_5168,N_9120);
or U10927 (N_10927,N_6860,N_5824);
nor U10928 (N_10928,N_6376,N_8663);
and U10929 (N_10929,N_8029,N_7346);
and U10930 (N_10930,N_8082,N_6548);
and U10931 (N_10931,N_8205,N_6624);
nand U10932 (N_10932,N_9475,N_9963);
or U10933 (N_10933,N_5114,N_5061);
and U10934 (N_10934,N_6637,N_9253);
or U10935 (N_10935,N_8399,N_7102);
nand U10936 (N_10936,N_6797,N_9948);
nor U10937 (N_10937,N_6486,N_7135);
or U10938 (N_10938,N_6260,N_7984);
nand U10939 (N_10939,N_7035,N_7252);
and U10940 (N_10940,N_7112,N_7003);
nand U10941 (N_10941,N_8203,N_9973);
and U10942 (N_10942,N_5093,N_9093);
or U10943 (N_10943,N_9520,N_8308);
nand U10944 (N_10944,N_5513,N_5278);
or U10945 (N_10945,N_5879,N_5333);
and U10946 (N_10946,N_9842,N_7352);
or U10947 (N_10947,N_9780,N_8664);
nand U10948 (N_10948,N_8683,N_9698);
nor U10949 (N_10949,N_5241,N_5330);
nand U10950 (N_10950,N_9198,N_8022);
nor U10951 (N_10951,N_9886,N_7718);
and U10952 (N_10952,N_6263,N_8773);
nand U10953 (N_10953,N_9605,N_8439);
and U10954 (N_10954,N_8965,N_6473);
nor U10955 (N_10955,N_9299,N_8599);
and U10956 (N_10956,N_7685,N_8207);
nand U10957 (N_10957,N_9585,N_9263);
nand U10958 (N_10958,N_7749,N_7513);
nand U10959 (N_10959,N_8242,N_8469);
nor U10960 (N_10960,N_8269,N_9558);
nor U10961 (N_10961,N_8602,N_9790);
and U10962 (N_10962,N_7284,N_6483);
nand U10963 (N_10963,N_5727,N_6857);
nor U10964 (N_10964,N_7360,N_9835);
xnor U10965 (N_10965,N_7550,N_9862);
nor U10966 (N_10966,N_8424,N_9538);
and U10967 (N_10967,N_9483,N_9530);
or U10968 (N_10968,N_9050,N_5892);
and U10969 (N_10969,N_6829,N_9216);
and U10970 (N_10970,N_8034,N_9125);
nand U10971 (N_10971,N_7981,N_8757);
and U10972 (N_10972,N_6836,N_6007);
or U10973 (N_10973,N_5683,N_6627);
nor U10974 (N_10974,N_7611,N_9029);
nand U10975 (N_10975,N_5776,N_5650);
nand U10976 (N_10976,N_7260,N_8254);
nand U10977 (N_10977,N_9863,N_7412);
and U10978 (N_10978,N_5251,N_5569);
and U10979 (N_10979,N_5614,N_9546);
nand U10980 (N_10980,N_6136,N_9423);
nor U10981 (N_10981,N_7365,N_7070);
nand U10982 (N_10982,N_9825,N_6090);
and U10983 (N_10983,N_8832,N_5160);
nor U10984 (N_10984,N_8180,N_5258);
or U10985 (N_10985,N_8542,N_5505);
or U10986 (N_10986,N_9802,N_8464);
or U10987 (N_10987,N_7998,N_6064);
or U10988 (N_10988,N_5696,N_5855);
nand U10989 (N_10989,N_5033,N_7547);
nor U10990 (N_10990,N_6861,N_6084);
or U10991 (N_10991,N_9102,N_8292);
and U10992 (N_10992,N_7548,N_6592);
nor U10993 (N_10993,N_7864,N_7900);
nand U10994 (N_10994,N_8563,N_7385);
or U10995 (N_10995,N_5051,N_6381);
nor U10996 (N_10996,N_6507,N_7834);
nand U10997 (N_10997,N_5046,N_6593);
and U10998 (N_10998,N_5412,N_8485);
or U10999 (N_10999,N_8786,N_6455);
or U11000 (N_11000,N_5526,N_5257);
nor U11001 (N_11001,N_8557,N_9548);
nor U11002 (N_11002,N_9237,N_5501);
nand U11003 (N_11003,N_6128,N_9622);
nand U11004 (N_11004,N_5097,N_9293);
or U11005 (N_11005,N_9208,N_8507);
and U11006 (N_11006,N_7587,N_7693);
nand U11007 (N_11007,N_8049,N_9390);
and U11008 (N_11008,N_8624,N_5475);
nand U11009 (N_11009,N_8167,N_9095);
nand U11010 (N_11010,N_9541,N_9988);
or U11011 (N_11011,N_8202,N_9716);
nor U11012 (N_11012,N_8303,N_6249);
nor U11013 (N_11013,N_7371,N_9173);
or U11014 (N_11014,N_5536,N_8893);
or U11015 (N_11015,N_9254,N_8410);
nand U11016 (N_11016,N_5445,N_6021);
nor U11017 (N_11017,N_9310,N_5678);
or U11018 (N_11018,N_7720,N_9793);
nand U11019 (N_11019,N_5553,N_6041);
or U11020 (N_11020,N_9772,N_6874);
and U11021 (N_11021,N_5710,N_9529);
or U11022 (N_11022,N_9169,N_9059);
nand U11023 (N_11023,N_8468,N_9653);
nand U11024 (N_11024,N_7914,N_7523);
and U11025 (N_11025,N_9556,N_5949);
nor U11026 (N_11026,N_5598,N_5432);
nand U11027 (N_11027,N_8831,N_5370);
and U11028 (N_11028,N_5875,N_9625);
nor U11029 (N_11029,N_7024,N_9856);
and U11030 (N_11030,N_8463,N_6951);
or U11031 (N_11031,N_8076,N_9586);
nor U11032 (N_11032,N_7164,N_6811);
and U11033 (N_11033,N_8543,N_9647);
and U11034 (N_11034,N_7887,N_8633);
nand U11035 (N_11035,N_6904,N_5466);
or U11036 (N_11036,N_5495,N_9738);
nand U11037 (N_11037,N_7678,N_6737);
nand U11038 (N_11038,N_9815,N_5522);
nand U11039 (N_11039,N_7313,N_7751);
or U11040 (N_11040,N_9994,N_9959);
or U11041 (N_11041,N_9411,N_5640);
and U11042 (N_11042,N_9072,N_6482);
and U11043 (N_11043,N_9441,N_7088);
nand U11044 (N_11044,N_5291,N_7799);
or U11045 (N_11045,N_7719,N_8963);
and U11046 (N_11046,N_6159,N_8159);
nand U11047 (N_11047,N_6556,N_6658);
or U11048 (N_11048,N_6217,N_8611);
and U11049 (N_11049,N_8209,N_6878);
nand U11050 (N_11050,N_9847,N_8351);
nor U11051 (N_11051,N_5270,N_6843);
or U11052 (N_11052,N_5738,N_6920);
nor U11053 (N_11053,N_9022,N_9362);
and U11054 (N_11054,N_6747,N_9062);
or U11055 (N_11055,N_8019,N_5200);
or U11056 (N_11056,N_9250,N_8580);
or U11057 (N_11057,N_9700,N_9696);
or U11058 (N_11058,N_5377,N_8798);
nand U11059 (N_11059,N_7766,N_8092);
nor U11060 (N_11060,N_8397,N_7458);
and U11061 (N_11061,N_8346,N_9650);
nor U11062 (N_11062,N_5156,N_9146);
and U11063 (N_11063,N_9235,N_7823);
or U11064 (N_11064,N_9561,N_7148);
and U11065 (N_11065,N_8003,N_8666);
nand U11066 (N_11066,N_7742,N_8883);
or U11067 (N_11067,N_5756,N_8495);
and U11068 (N_11068,N_9516,N_5632);
nor U11069 (N_11069,N_8655,N_9343);
nand U11070 (N_11070,N_8680,N_6905);
or U11071 (N_11071,N_5624,N_7828);
nor U11072 (N_11072,N_8972,N_6691);
nor U11073 (N_11073,N_6851,N_9914);
or U11074 (N_11074,N_7082,N_6400);
and U11075 (N_11075,N_7176,N_8444);
xnor U11076 (N_11076,N_8011,N_6879);
nor U11077 (N_11077,N_6414,N_6251);
and U11078 (N_11078,N_7879,N_5183);
nor U11079 (N_11079,N_5350,N_7994);
nor U11080 (N_11080,N_5911,N_9243);
nor U11081 (N_11081,N_7340,N_8065);
nor U11082 (N_11082,N_7211,N_6663);
or U11083 (N_11083,N_6689,N_5048);
nand U11084 (N_11084,N_7729,N_5759);
nor U11085 (N_11085,N_5848,N_9575);
nand U11086 (N_11086,N_5535,N_9309);
or U11087 (N_11087,N_9074,N_8083);
or U11088 (N_11088,N_8017,N_5753);
or U11089 (N_11089,N_6882,N_6620);
nor U11090 (N_11090,N_8107,N_7478);
nand U11091 (N_11091,N_5144,N_7583);
or U11092 (N_11092,N_5301,N_6674);
nand U11093 (N_11093,N_8135,N_5112);
nor U11094 (N_11094,N_8259,N_9920);
nor U11095 (N_11095,N_5389,N_8966);
nor U11096 (N_11096,N_9918,N_6684);
nor U11097 (N_11097,N_7999,N_8654);
nand U11098 (N_11098,N_6916,N_5881);
nand U11099 (N_11099,N_5596,N_6456);
nor U11100 (N_11100,N_5239,N_6088);
nor U11101 (N_11101,N_6519,N_9471);
or U11102 (N_11102,N_5229,N_7113);
or U11103 (N_11103,N_9457,N_8023);
nor U11104 (N_11104,N_8032,N_9940);
nand U11105 (N_11105,N_8988,N_5608);
nand U11106 (N_11106,N_9458,N_9335);
nor U11107 (N_11107,N_5645,N_9279);
and U11108 (N_11108,N_7338,N_9965);
or U11109 (N_11109,N_7180,N_9261);
or U11110 (N_11110,N_6356,N_8027);
nand U11111 (N_11111,N_6508,N_6766);
nand U11112 (N_11112,N_5374,N_5838);
nand U11113 (N_11113,N_6682,N_8451);
nand U11114 (N_11114,N_6786,N_8488);
nor U11115 (N_11115,N_5349,N_9894);
or U11116 (N_11116,N_6561,N_8970);
and U11117 (N_11117,N_8366,N_8959);
nor U11118 (N_11118,N_9908,N_5136);
nor U11119 (N_11119,N_5620,N_9925);
nand U11120 (N_11120,N_8982,N_5397);
and U11121 (N_11121,N_6911,N_6953);
nand U11122 (N_11122,N_8217,N_5476);
nand U11123 (N_11123,N_9304,N_8183);
nand U11124 (N_11124,N_7379,N_6999);
and U11125 (N_11125,N_6282,N_9803);
and U11126 (N_11126,N_6265,N_7654);
nand U11127 (N_11127,N_5595,N_8369);
nand U11128 (N_11128,N_8372,N_8733);
or U11129 (N_11129,N_7452,N_5086);
nor U11130 (N_11130,N_6315,N_7975);
nand U11131 (N_11131,N_9868,N_8161);
and U11132 (N_11132,N_8638,N_8498);
nor U11133 (N_11133,N_9945,N_7305);
nor U11134 (N_11134,N_7274,N_7028);
nor U11135 (N_11135,N_8841,N_7713);
and U11136 (N_11136,N_5391,N_8807);
or U11137 (N_11137,N_7841,N_5769);
nand U11138 (N_11138,N_9239,N_8618);
nand U11139 (N_11139,N_7803,N_8833);
nand U11140 (N_11140,N_6236,N_6962);
nor U11141 (N_11141,N_8060,N_7025);
and U11142 (N_11142,N_5550,N_8447);
or U11143 (N_11143,N_7233,N_8114);
nor U11144 (N_11144,N_8740,N_6366);
and U11145 (N_11145,N_9401,N_5969);
or U11146 (N_11146,N_7771,N_6819);
nor U11147 (N_11147,N_8958,N_6415);
nor U11148 (N_11148,N_9934,N_7533);
or U11149 (N_11149,N_7293,N_6387);
or U11150 (N_11150,N_6943,N_5713);
nand U11151 (N_11151,N_5987,N_9400);
or U11152 (N_11152,N_6059,N_7860);
or U11153 (N_11153,N_6144,N_6774);
nand U11154 (N_11154,N_7628,N_7917);
nand U11155 (N_11155,N_5189,N_5310);
nand U11156 (N_11156,N_7217,N_8501);
nor U11157 (N_11157,N_9648,N_5826);
and U11158 (N_11158,N_9879,N_5287);
nor U11159 (N_11159,N_8037,N_5809);
nand U11160 (N_11160,N_6613,N_7535);
and U11161 (N_11161,N_7843,N_8436);
nor U11162 (N_11162,N_5902,N_6408);
and U11163 (N_11163,N_6568,N_5073);
nor U11164 (N_11164,N_7481,N_6858);
nand U11165 (N_11165,N_5642,N_7163);
xor U11166 (N_11166,N_8151,N_8381);
and U11167 (N_11167,N_5023,N_6054);
nand U11168 (N_11168,N_9899,N_8559);
xnor U11169 (N_11169,N_9628,N_7425);
or U11170 (N_11170,N_5917,N_5792);
or U11171 (N_11171,N_5900,N_8250);
and U11172 (N_11172,N_8994,N_8243);
nand U11173 (N_11173,N_5806,N_8910);
nand U11174 (N_11174,N_8789,N_6563);
or U11175 (N_11175,N_5457,N_8198);
and U11176 (N_11176,N_5754,N_6197);
nand U11177 (N_11177,N_9512,N_5854);
or U11178 (N_11178,N_8549,N_9221);
nand U11179 (N_11179,N_6367,N_5982);
nor U11180 (N_11180,N_6436,N_6085);
nand U11181 (N_11181,N_6554,N_9126);
and U11182 (N_11182,N_9860,N_7761);
nor U11183 (N_11183,N_8877,N_8908);
and U11184 (N_11184,N_7415,N_6948);
and U11185 (N_11185,N_8071,N_5131);
nor U11186 (N_11186,N_6975,N_6470);
nor U11187 (N_11187,N_8921,N_9099);
nor U11188 (N_11188,N_5557,N_5702);
and U11189 (N_11189,N_8211,N_5722);
and U11190 (N_11190,N_9944,N_7902);
nand U11191 (N_11191,N_7778,N_9987);
or U11192 (N_11192,N_8747,N_9822);
nand U11193 (N_11193,N_5411,N_8499);
nor U11194 (N_11194,N_5214,N_9393);
nor U11195 (N_11195,N_5919,N_7995);
nand U11196 (N_11196,N_8197,N_5158);
nor U11197 (N_11197,N_8928,N_9323);
or U11198 (N_11198,N_6343,N_6912);
nand U11199 (N_11199,N_8984,N_5641);
or U11200 (N_11200,N_6704,N_5603);
nand U11201 (N_11201,N_8266,N_6200);
and U11202 (N_11202,N_5068,N_7762);
nor U11203 (N_11203,N_5654,N_6358);
nor U11204 (N_11204,N_9787,N_9430);
and U11205 (N_11205,N_7462,N_9983);
nor U11206 (N_11206,N_6898,N_5880);
and U11207 (N_11207,N_6701,N_9258);
and U11208 (N_11208,N_5948,N_9592);
and U11209 (N_11209,N_5341,N_5865);
nor U11210 (N_11210,N_9164,N_9978);
nor U11211 (N_11211,N_5730,N_9851);
or U11212 (N_11212,N_7855,N_7265);
nor U11213 (N_11213,N_7094,N_6294);
nand U11214 (N_11214,N_7368,N_7298);
and U11215 (N_11215,N_6566,N_8188);
and U11216 (N_11216,N_7689,N_6750);
nand U11217 (N_11217,N_9595,N_8593);
and U11218 (N_11218,N_9338,N_8813);
nor U11219 (N_11219,N_6334,N_7188);
xnor U11220 (N_11220,N_6855,N_7421);
and U11221 (N_11221,N_5207,N_8497);
nand U11222 (N_11222,N_9398,N_8875);
and U11223 (N_11223,N_9487,N_6146);
nor U11224 (N_11224,N_6181,N_7579);
nor U11225 (N_11225,N_6963,N_9245);
and U11226 (N_11226,N_5273,N_5034);
or U11227 (N_11227,N_8324,N_7601);
nor U11228 (N_11228,N_6526,N_8072);
nor U11229 (N_11229,N_7270,N_5471);
nor U11230 (N_11230,N_8509,N_9657);
and U11231 (N_11231,N_9071,N_5923);
nor U11232 (N_11232,N_8670,N_5812);
and U11233 (N_11233,N_8166,N_5512);
nand U11234 (N_11234,N_5117,N_7939);
or U11235 (N_11235,N_9504,N_5819);
and U11236 (N_11236,N_5417,N_6342);
nor U11237 (N_11237,N_6785,N_9588);
nor U11238 (N_11238,N_5679,N_7087);
or U11239 (N_11239,N_7332,N_5090);
xor U11240 (N_11240,N_9606,N_8033);
nand U11241 (N_11241,N_9353,N_6350);
nand U11242 (N_11242,N_8847,N_7940);
or U11243 (N_11243,N_5575,N_9088);
and U11244 (N_11244,N_9115,N_5933);
nand U11245 (N_11245,N_7881,N_5597);
or U11246 (N_11246,N_8828,N_9248);
and U11247 (N_11247,N_5714,N_7889);
nand U11248 (N_11248,N_6242,N_6776);
nand U11249 (N_11249,N_8631,N_8716);
or U11250 (N_11250,N_8172,N_8026);
or U11251 (N_11251,N_7117,N_6967);
or U11252 (N_11252,N_5604,N_7990);
and U11253 (N_11253,N_7153,N_8775);
and U11254 (N_11254,N_7986,N_8164);
and U11255 (N_11255,N_5635,N_7806);
or U11256 (N_11256,N_5244,N_7218);
nand U11257 (N_11257,N_5627,N_5323);
nand U11258 (N_11258,N_6531,N_9149);
or U11259 (N_11259,N_9367,N_9416);
and U11260 (N_11260,N_5718,N_7949);
nand U11261 (N_11261,N_6185,N_6807);
or U11262 (N_11262,N_9991,N_9702);
and U11263 (N_11263,N_8251,N_9024);
and U11264 (N_11264,N_8704,N_5041);
nor U11265 (N_11265,N_8075,N_7721);
nand U11266 (N_11266,N_9832,N_5803);
nor U11267 (N_11267,N_8118,N_9453);
nor U11268 (N_11268,N_5782,N_5699);
nor U11269 (N_11269,N_7096,N_8702);
nand U11270 (N_11270,N_5367,N_9069);
nor U11271 (N_11271,N_6758,N_5874);
nand U11272 (N_11272,N_8280,N_7172);
or U11273 (N_11273,N_7697,N_7493);
nor U11274 (N_11274,N_7118,N_5711);
nor U11275 (N_11275,N_9727,N_7517);
and U11276 (N_11276,N_6557,N_6360);
nor U11277 (N_11277,N_9591,N_8300);
or U11278 (N_11278,N_9215,N_9971);
and U11279 (N_11279,N_9420,N_8639);
nand U11280 (N_11280,N_8842,N_9610);
nor U11281 (N_11281,N_5286,N_7157);
nor U11282 (N_11282,N_7224,N_6733);
nor U11283 (N_11283,N_6093,N_8763);
nand U11284 (N_11284,N_6363,N_9915);
nand U11285 (N_11285,N_5798,N_5964);
or U11286 (N_11286,N_6949,N_7160);
nand U11287 (N_11287,N_6844,N_8993);
or U11288 (N_11288,N_6351,N_5171);
nor U11289 (N_11289,N_6361,N_8453);
nor U11290 (N_11290,N_8042,N_7800);
or U11291 (N_11291,N_5408,N_5154);
or U11292 (N_11292,N_8332,N_8093);
nor U11293 (N_11293,N_6767,N_8122);
nand U11294 (N_11294,N_7097,N_7030);
nand U11295 (N_11295,N_8556,N_7479);
or U11296 (N_11296,N_5028,N_6440);
nor U11297 (N_11297,N_6964,N_6451);
nand U11298 (N_11298,N_5884,N_5387);
nor U11299 (N_11299,N_5410,N_9692);
and U11300 (N_11300,N_8371,N_6871);
nor U11301 (N_11301,N_5687,N_7271);
nor U11302 (N_11302,N_8750,N_6448);
nand U11303 (N_11303,N_5528,N_8863);
nand U11304 (N_11304,N_6734,N_8566);
nor U11305 (N_11305,N_9381,N_5621);
and U11306 (N_11306,N_6732,N_5701);
nand U11307 (N_11307,N_5493,N_9532);
nand U11308 (N_11308,N_7072,N_5731);
nor U11309 (N_11309,N_6058,N_6780);
or U11310 (N_11310,N_8899,N_7591);
nand U11311 (N_11311,N_5814,N_8147);
nand U11312 (N_11312,N_7888,N_7424);
nor U11313 (N_11313,N_9503,N_9777);
and U11314 (N_11314,N_9786,N_5106);
nand U11315 (N_11315,N_9644,N_6353);
nor U11316 (N_11316,N_9251,N_5544);
nand U11317 (N_11317,N_6779,N_5672);
nor U11318 (N_11318,N_5094,N_6393);
nor U11319 (N_11319,N_5210,N_6348);
and U11320 (N_11320,N_6076,N_9666);
or U11321 (N_11321,N_8110,N_7062);
and U11322 (N_11322,N_6573,N_8720);
nor U11323 (N_11323,N_8035,N_9185);
and U11324 (N_11324,N_7170,N_6183);
and U11325 (N_11325,N_5773,N_7717);
nor U11326 (N_11326,N_7073,N_7726);
nand U11327 (N_11327,N_5894,N_5721);
nand U11328 (N_11328,N_7577,N_6850);
and U11329 (N_11329,N_5259,N_7826);
nor U11330 (N_11330,N_6795,N_8738);
and U11331 (N_11331,N_7976,N_5849);
xor U11332 (N_11332,N_8676,N_8323);
or U11333 (N_11333,N_9846,N_5760);
nand U11334 (N_11334,N_6503,N_8526);
and U11335 (N_11335,N_9358,N_9933);
and U11336 (N_11336,N_9910,N_5556);
nand U11337 (N_11337,N_7700,N_7872);
or U11338 (N_11338,N_6492,N_7862);
and U11339 (N_11339,N_9540,N_9314);
nor U11340 (N_11340,N_5567,N_9715);
nor U11341 (N_11341,N_8915,N_7909);
xnor U11342 (N_11342,N_8290,N_9025);
nor U11343 (N_11343,N_8962,N_6100);
or U11344 (N_11344,N_7763,N_7002);
and U11345 (N_11345,N_7927,N_7204);
nand U11346 (N_11346,N_7543,N_6349);
nor U11347 (N_11347,N_5761,N_9688);
or U11348 (N_11348,N_7969,N_5313);
nor U11349 (N_11349,N_6138,N_7422);
or U11350 (N_11350,N_6163,N_9770);
and U11351 (N_11351,N_7417,N_9767);
and U11352 (N_11352,N_7453,N_9798);
and U11353 (N_11353,N_5382,N_8362);
nand U11354 (N_11354,N_6111,N_7945);
and U11355 (N_11355,N_6318,N_7567);
and U11356 (N_11356,N_6794,N_6499);
nor U11357 (N_11357,N_5610,N_8712);
and U11358 (N_11358,N_7519,N_6053);
nor U11359 (N_11359,N_7798,N_6143);
nor U11360 (N_11360,N_8547,N_6182);
nand U11361 (N_11361,N_9549,N_8370);
nor U11362 (N_11362,N_5386,N_6909);
and U11363 (N_11363,N_7506,N_9873);
and U11364 (N_11364,N_8586,N_5236);
nor U11365 (N_11365,N_5936,N_7374);
or U11366 (N_11366,N_7241,N_9946);
nand U11367 (N_11367,N_9348,N_7960);
nand U11368 (N_11368,N_5309,N_6668);
nand U11369 (N_11369,N_5928,N_6534);
nand U11370 (N_11370,N_6715,N_9394);
nand U11371 (N_11371,N_9869,N_8148);
and U11372 (N_11372,N_9377,N_5937);
or U11373 (N_11373,N_6038,N_6539);
nand U11374 (N_11374,N_9214,N_5492);
nor U11375 (N_11375,N_8068,N_7401);
nand U11376 (N_11376,N_8673,N_8727);
xnor U11377 (N_11377,N_5359,N_8426);
nand U11378 (N_11378,N_6687,N_5400);
nand U11379 (N_11379,N_7932,N_5577);
and U11380 (N_11380,N_9260,N_8337);
and U11381 (N_11381,N_9138,N_5886);
nor U11382 (N_11382,N_9794,N_5741);
nor U11383 (N_11383,N_9515,N_6392);
nand U11384 (N_11384,N_9859,N_7753);
and U11385 (N_11385,N_7439,N_6379);
or U11386 (N_11386,N_9140,N_9030);
nand U11387 (N_11387,N_9332,N_5637);
and U11388 (N_11388,N_7304,N_7936);
nand U11389 (N_11389,N_7213,N_5477);
or U11390 (N_11390,N_5724,N_9506);
and U11391 (N_11391,N_9630,N_5193);
nand U11392 (N_11392,N_5147,N_9524);
and U11393 (N_11393,N_6629,N_5065);
nand U11394 (N_11394,N_9313,N_5308);
nor U11395 (N_11395,N_9828,N_5402);
xor U11396 (N_11396,N_7354,N_5470);
nor U11397 (N_11397,N_8651,N_6301);
xor U11398 (N_11398,N_6210,N_8435);
nor U11399 (N_11399,N_7036,N_5177);
and U11400 (N_11400,N_6872,N_9881);
or U11401 (N_11401,N_6273,N_6892);
and U11402 (N_11402,N_7924,N_7764);
nor U11403 (N_11403,N_8815,N_6615);
nand U11404 (N_11404,N_5951,N_8239);
nand U11405 (N_11405,N_8894,N_5976);
and U11406 (N_11406,N_5145,N_6344);
nand U11407 (N_11407,N_7226,N_6335);
and U11408 (N_11408,N_7343,N_5561);
or U11409 (N_11409,N_6890,N_5508);
or U11410 (N_11410,N_8428,N_6901);
or U11411 (N_11411,N_6096,N_6736);
nand U11412 (N_11412,N_9240,N_9880);
and U11413 (N_11413,N_5002,N_9631);
nor U11414 (N_11414,N_9539,N_5371);
or U11415 (N_11415,N_6925,N_7145);
nor U11416 (N_11416,N_9165,N_6165);
nor U11417 (N_11417,N_6708,N_5419);
nand U11418 (N_11418,N_9810,N_5461);
nand U11419 (N_11419,N_6233,N_7007);
xnor U11420 (N_11420,N_7442,N_9762);
and U11421 (N_11421,N_5279,N_5080);
nor U11422 (N_11422,N_9427,N_9242);
or U11423 (N_11423,N_5182,N_6585);
and U11424 (N_11424,N_8361,N_6284);
nor U11425 (N_11425,N_9345,N_7613);
and U11426 (N_11426,N_9935,N_8171);
and U11427 (N_11427,N_5483,N_8268);
xnor U11428 (N_11428,N_9552,N_7084);
or U11429 (N_11429,N_9305,N_9757);
nand U11430 (N_11430,N_9765,N_7930);
nor U11431 (N_11431,N_5622,N_8667);
or U11432 (N_11432,N_6230,N_9057);
and U11433 (N_11433,N_5429,N_5887);
or U11434 (N_11434,N_9178,N_6160);
nor U11435 (N_11435,N_8876,N_8824);
nand U11436 (N_11436,N_6988,N_7633);
and U11437 (N_11437,N_6224,N_8311);
nor U11438 (N_11438,N_5994,N_6588);
nor U11439 (N_11439,N_9463,N_7554);
nor U11440 (N_11440,N_8591,N_7951);
nor U11441 (N_11441,N_8284,N_5076);
and U11442 (N_11442,N_6404,N_5264);
or U11443 (N_11443,N_6917,N_9719);
nor U11444 (N_11444,N_7071,N_5684);
nor U11445 (N_11445,N_7596,N_9113);
nor U11446 (N_11446,N_9890,N_7259);
nor U11447 (N_11447,N_9219,N_6998);
or U11448 (N_11448,N_5539,N_5455);
and U11449 (N_11449,N_9163,N_7216);
nand U11450 (N_11450,N_9642,N_5187);
nor U11451 (N_11451,N_8696,N_6323);
or U11452 (N_11452,N_6604,N_7342);
nor U11453 (N_11453,N_9223,N_5870);
or U11454 (N_11454,N_8412,N_7490);
nand U11455 (N_11455,N_9083,N_5052);
or U11456 (N_11456,N_8619,N_6433);
or U11457 (N_11457,N_9371,N_8722);
or U11458 (N_11458,N_7042,N_8108);
nand U11459 (N_11459,N_5414,N_5783);
nor U11460 (N_11460,N_9893,N_7973);
nand U11461 (N_11461,N_7980,N_8913);
or U11462 (N_11462,N_5941,N_6396);
nor U11463 (N_11463,N_8992,N_9517);
and U11464 (N_11464,N_8319,N_6685);
and U11465 (N_11465,N_6352,N_6052);
and U11466 (N_11466,N_7166,N_8592);
nor U11467 (N_11467,N_5500,N_8918);
nor U11468 (N_11468,N_5084,N_8246);
or U11469 (N_11469,N_9151,N_5118);
nand U11470 (N_11470,N_5277,N_7584);
or U11471 (N_11471,N_6019,N_6979);
or U11472 (N_11472,N_5070,N_5140);
and U11473 (N_11473,N_7706,N_8387);
and U11474 (N_11474,N_7080,N_7541);
nand U11475 (N_11475,N_8690,N_7480);
nand U11476 (N_11476,N_5355,N_9128);
nor U11477 (N_11477,N_8154,N_5590);
and U11478 (N_11478,N_6518,N_9858);
or U11479 (N_11479,N_5015,N_9225);
and U11480 (N_11480,N_8452,N_6281);
nor U11481 (N_11481,N_9112,N_9992);
or U11482 (N_11482,N_7104,N_9341);
nand U11483 (N_11483,N_9952,N_7023);
nor U11484 (N_11484,N_5857,N_9551);
nand U11485 (N_11485,N_9788,N_7961);
xnor U11486 (N_11486,N_6968,N_5100);
or U11487 (N_11487,N_7189,N_7754);
nand U11488 (N_11488,N_7139,N_6261);
nor U11489 (N_11489,N_5130,N_9675);
and U11490 (N_11490,N_9020,N_9665);
and U11491 (N_11491,N_6510,N_8134);
or U11492 (N_11492,N_7321,N_7345);
nand U11493 (N_11493,N_5527,N_6578);
and U11494 (N_11494,N_5867,N_7703);
nor U11495 (N_11495,N_6880,N_7599);
or U11496 (N_11496,N_9283,N_7029);
or U11497 (N_11497,N_5299,N_5479);
nand U11498 (N_11498,N_8612,N_5044);
and U11499 (N_11499,N_8210,N_7522);
and U11500 (N_11500,N_6467,N_6738);
nand U11501 (N_11501,N_6189,N_8967);
nor U11502 (N_11502,N_7106,N_9464);
nor U11503 (N_11503,N_9334,N_5092);
nand U11504 (N_11504,N_8513,N_8194);
or U11505 (N_11505,N_5653,N_6447);
or U11506 (N_11506,N_7381,N_9355);
nor U11507 (N_11507,N_8123,N_5871);
or U11508 (N_11508,N_9465,N_6212);
nand U11509 (N_11509,N_7447,N_9775);
nand U11510 (N_11510,N_5634,N_6538);
or U11511 (N_11511,N_7950,N_6631);
nor U11512 (N_11512,N_6121,N_6256);
or U11513 (N_11513,N_5135,N_9492);
nand U11514 (N_11514,N_6721,N_6147);
nor U11515 (N_11515,N_8743,N_5839);
nor U11516 (N_11516,N_6203,N_9662);
nand U11517 (N_11517,N_9636,N_7714);
and U11518 (N_11518,N_5462,N_7357);
or U11519 (N_11519,N_8771,N_9342);
and U11520 (N_11520,N_9553,N_9672);
xnor U11521 (N_11521,N_5885,N_6450);
nor U11522 (N_11522,N_5062,N_8912);
or U11523 (N_11523,N_6537,N_9511);
or U11524 (N_11524,N_9333,N_5816);
and U11525 (N_11525,N_8836,N_7684);
nand U11526 (N_11526,N_9486,N_5014);
nor U11527 (N_11527,N_8595,N_9536);
or U11528 (N_11528,N_7156,N_5162);
nor U11529 (N_11529,N_6092,N_6535);
nor U11530 (N_11530,N_7013,N_7359);
and U11531 (N_11531,N_5758,N_9964);
nand U11532 (N_11532,N_6423,N_5143);
nor U11533 (N_11533,N_9921,N_5863);
and U11534 (N_11534,N_7809,N_5739);
nand U11535 (N_11535,N_9854,N_8265);
or U11536 (N_11536,N_7149,N_7169);
or U11537 (N_11537,N_9047,N_6317);
nand U11538 (N_11538,N_5649,N_5752);
and U11539 (N_11539,N_6888,N_5762);
and U11540 (N_11540,N_9321,N_9510);
nand U11541 (N_11541,N_5748,N_7376);
nor U11542 (N_11542,N_6247,N_5064);
nand U11543 (N_11543,N_6045,N_8969);
and U11544 (N_11544,N_5152,N_9134);
nand U11545 (N_11545,N_5651,N_9384);
nand U11546 (N_11546,N_9613,N_7129);
nand U11547 (N_11547,N_5450,N_9437);
nor U11548 (N_11548,N_5472,N_5639);
nand U11549 (N_11549,N_9560,N_6814);
nor U11550 (N_11550,N_7205,N_8553);
xor U11551 (N_11551,N_7923,N_5992);
or U11552 (N_11552,N_8532,N_9682);
nand U11553 (N_11553,N_6710,N_6157);
and U11554 (N_11554,N_5618,N_8779);
nand U11555 (N_11555,N_7905,N_6514);
and U11556 (N_11556,N_8746,N_7609);
nand U11557 (N_11557,N_6842,N_8053);
nand U11558 (N_11558,N_8233,N_5704);
nor U11559 (N_11559,N_6572,N_9361);
nor U11560 (N_11560,N_8658,N_8849);
nand U11561 (N_11561,N_7161,N_6885);
nor U11562 (N_11562,N_9301,N_6040);
or U11563 (N_11563,N_9750,N_7941);
nor U11564 (N_11564,N_5576,N_7325);
nand U11565 (N_11565,N_8357,N_7334);
nor U11566 (N_11566,N_6727,N_9363);
nor U11567 (N_11567,N_5853,N_5077);
and U11568 (N_11568,N_8834,N_5095);
or U11569 (N_11569,N_8406,N_9737);
and U11570 (N_11570,N_9509,N_8462);
and U11571 (N_11571,N_9141,N_9286);
and U11572 (N_11572,N_5407,N_8316);
and U11573 (N_11573,N_7741,N_6416);
nand U11574 (N_11574,N_8376,N_8105);
or U11575 (N_11575,N_6635,N_8884);
and U11576 (N_11576,N_7861,N_9383);
or U11577 (N_11577,N_7643,N_5098);
nor U11578 (N_11578,N_7856,N_5765);
nor U11579 (N_11579,N_8916,N_6432);
or U11580 (N_11580,N_8820,N_6489);
nor U11581 (N_11581,N_5134,N_9212);
nor U11582 (N_11582,N_6865,N_8520);
or U11583 (N_11583,N_9226,N_6421);
nand U11584 (N_11584,N_9217,N_6752);
nand U11585 (N_11585,N_6692,N_9203);
nor U11586 (N_11586,N_9729,N_5306);
nor U11587 (N_11587,N_5778,N_7056);
nor U11588 (N_11588,N_7498,N_9233);
nand U11589 (N_11589,N_5272,N_7027);
and U11590 (N_11590,N_8800,N_9386);
or U11591 (N_11591,N_7600,N_7796);
and U11592 (N_11592,N_8390,N_8646);
nor U11593 (N_11593,N_9435,N_6509);
nor U11594 (N_11594,N_6304,N_5977);
or U11595 (N_11595,N_6098,N_7257);
or U11596 (N_11596,N_6044,N_8555);
nor U11597 (N_11597,N_6081,N_8756);
and U11598 (N_11598,N_7901,N_7508);
nand U11599 (N_11599,N_9291,N_5728);
and U11600 (N_11600,N_5847,N_8175);
or U11601 (N_11601,N_7486,N_5449);
or U11602 (N_11602,N_9995,N_6287);
and U11603 (N_11603,N_6887,N_7845);
or U11604 (N_11604,N_7048,N_7497);
or U11605 (N_11605,N_7645,N_7572);
nand U11606 (N_11606,N_9176,N_8006);
nor U11607 (N_11607,N_6828,N_8561);
nand U11608 (N_11608,N_6848,N_8837);
or U11609 (N_11609,N_8764,N_6928);
xnor U11610 (N_11610,N_8186,N_5668);
nand U11611 (N_11611,N_6527,N_7708);
nor U11612 (N_11612,N_9990,N_5256);
or U11613 (N_11613,N_6938,N_6150);
and U11614 (N_11614,N_5940,N_9008);
and U11615 (N_11615,N_5942,N_5747);
or U11616 (N_11616,N_6192,N_7942);
nand U11617 (N_11617,N_7947,N_8677);
nor U11618 (N_11618,N_7126,N_7009);
nand U11619 (N_11619,N_9017,N_7423);
nand U11620 (N_11620,N_8117,N_5037);
nor U11621 (N_11621,N_8568,N_7885);
or U11622 (N_11622,N_5532,N_6719);
or U11623 (N_11623,N_8156,N_6789);
and U11624 (N_11624,N_7179,N_5638);
and U11625 (N_11625,N_7663,N_8684);
nand U11626 (N_11626,N_7492,N_8050);
or U11627 (N_11627,N_8336,N_8792);
nand U11628 (N_11628,N_6718,N_8176);
and U11629 (N_11629,N_7031,N_8285);
or U11630 (N_11630,N_6643,N_8190);
and U11631 (N_11631,N_7147,N_6403);
and U11632 (N_11632,N_8838,N_6669);
nor U11633 (N_11633,N_9414,N_9272);
nand U11634 (N_11634,N_8200,N_7912);
nand U11635 (N_11635,N_6341,N_8106);
nand U11636 (N_11636,N_6825,N_5053);
nand U11637 (N_11637,N_9898,N_8759);
nand U11638 (N_11638,N_7978,N_6806);
nand U11639 (N_11639,N_5416,N_5000);
and U11640 (N_11640,N_7722,N_6771);
or U11641 (N_11641,N_8402,N_6278);
xor U11642 (N_11642,N_6707,N_5749);
nand U11643 (N_11643,N_6302,N_5274);
nand U11644 (N_11644,N_8348,N_8577);
nand U11645 (N_11645,N_5820,N_6153);
and U11646 (N_11646,N_5269,N_6500);
and U11647 (N_11647,N_5494,N_8299);
nor U11648 (N_11648,N_9745,N_9063);
nor U11649 (N_11649,N_9668,N_8133);
and U11650 (N_11650,N_9447,N_8215);
nand U11651 (N_11651,N_6374,N_7290);
and U11652 (N_11652,N_6731,N_7610);
nor U11653 (N_11653,N_7592,N_6693);
xor U11654 (N_11654,N_7673,N_5063);
or U11655 (N_11655,N_6373,N_9061);
or U11656 (N_11656,N_6156,N_6608);
or U11657 (N_11657,N_8244,N_8630);
nand U11658 (N_11658,N_9679,N_8749);
nand U11659 (N_11659,N_7482,N_6954);
nand U11660 (N_11660,N_7208,N_6763);
and U11661 (N_11661,N_8625,N_5586);
nand U11662 (N_11662,N_7474,N_6442);
or U11663 (N_11663,N_9681,N_7465);
or U11664 (N_11664,N_8138,N_8364);
nand U11665 (N_11665,N_8086,N_6595);
nor U11666 (N_11666,N_8124,N_7647);
or U11667 (N_11667,N_9876,N_6238);
nand U11668 (N_11668,N_7059,N_5021);
nand U11669 (N_11669,N_5767,N_6014);
and U11670 (N_11670,N_6002,N_7285);
nand U11671 (N_11671,N_6775,N_5841);
nor U11672 (N_11672,N_7542,N_9231);
and U11673 (N_11673,N_7292,N_6171);
nand U11674 (N_11674,N_8665,N_8848);
nor U11675 (N_11675,N_7426,N_5366);
or U11676 (N_11676,N_7197,N_7408);
and U11677 (N_11677,N_6219,N_9105);
nor U11678 (N_11678,N_7386,N_5478);
or U11679 (N_11679,N_8080,N_6196);
or U11680 (N_11680,N_7982,N_7568);
nor U11681 (N_11681,N_8871,N_6298);
and U11682 (N_11682,N_9927,N_6730);
nor U11683 (N_11683,N_7560,N_9583);
nand U11684 (N_11684,N_7184,N_9958);
and U11685 (N_11685,N_8515,N_8132);
nand U11686 (N_11686,N_9110,N_8768);
nand U11687 (N_11687,N_6394,N_5643);
nor U11688 (N_11688,N_7440,N_7116);
and U11689 (N_11689,N_5428,N_8473);
and U11690 (N_11690,N_8295,N_5989);
and U11691 (N_11691,N_9912,N_6971);
nor U11692 (N_11692,N_7503,N_7165);
nand U11693 (N_11693,N_8853,N_5939);
nor U11694 (N_11694,N_7526,N_7435);
nor U11695 (N_11695,N_9956,N_8603);
nor U11696 (N_11696,N_9002,N_9368);
nor U11697 (N_11697,N_8949,N_5298);
and U11698 (N_11698,N_5685,N_5104);
nand U11699 (N_11699,N_6939,N_8858);
xnor U11700 (N_11700,N_7867,N_8470);
and U11701 (N_11701,N_8048,N_9725);
nand U11702 (N_11702,N_8454,N_6594);
or U11703 (N_11703,N_9704,N_8924);
nand U11704 (N_11704,N_7151,N_7308);
nor U11705 (N_11705,N_7534,N_7847);
and U11706 (N_11706,N_8040,N_6446);
and U11707 (N_11707,N_5334,N_5127);
or U11708 (N_11708,N_8584,N_9614);
nand U11709 (N_11709,N_7362,N_5039);
xor U11710 (N_11710,N_8656,N_6529);
nor U11711 (N_11711,N_5558,N_5213);
or U11712 (N_11712,N_8472,N_6983);
and U11713 (N_11713,N_8229,N_6277);
or U11714 (N_11714,N_8097,N_9425);
or U11715 (N_11715,N_9049,N_9259);
and U11716 (N_11716,N_7283,N_6359);
and U11717 (N_11717,N_5636,N_6279);
nor U11718 (N_11718,N_6633,N_5459);
and U11719 (N_11719,N_7108,N_7852);
and U11720 (N_11720,N_5348,N_9318);
and U11721 (N_11721,N_9410,N_8861);
nand U11722 (N_11722,N_6982,N_9658);
nand U11723 (N_11723,N_6846,N_8359);
nor U11724 (N_11724,N_7441,N_7443);
and U11725 (N_11725,N_9906,N_7491);
nand U11726 (N_11726,N_7851,N_5978);
and U11727 (N_11727,N_9889,N_6533);
nand U11728 (N_11728,N_6135,N_6552);
and U11729 (N_11729,N_7757,N_5155);
and U11730 (N_11730,N_6559,N_6632);
nor U11731 (N_11731,N_9710,N_9849);
nor U11732 (N_11732,N_6712,N_9257);
nand U11733 (N_11733,N_9202,N_7576);
nor U11734 (N_11734,N_8327,N_9744);
or U11735 (N_11735,N_8419,N_7182);
or U11736 (N_11736,N_6977,N_5192);
nand U11737 (N_11737,N_6472,N_5025);
nand U11738 (N_11738,N_7240,N_5791);
nor U11739 (N_11739,N_5998,N_9778);
or U11740 (N_11740,N_8544,N_9424);
and U11741 (N_11741,N_8953,N_8179);
nor U11742 (N_11742,N_7734,N_8778);
or U11743 (N_11743,N_8422,N_5766);
nor U11744 (N_11744,N_9982,N_8286);
and U11745 (N_11745,N_9122,N_7590);
nand U11746 (N_11746,N_9359,N_6782);
nor U11747 (N_11747,N_9444,N_6193);
or U11748 (N_11748,N_7501,N_9108);
nand U11749 (N_11749,N_7765,N_9621);
or U11750 (N_11750,N_7680,N_7192);
nor U11751 (N_11751,N_6435,N_8095);
and U11752 (N_11752,N_9950,N_8162);
and U11753 (N_11753,N_9389,N_6493);
nor U11754 (N_11754,N_6202,N_7200);
nor U11755 (N_11755,N_5451,N_7730);
and U11756 (N_11756,N_5197,N_8830);
and U11757 (N_11757,N_9841,N_5442);
or U11758 (N_11758,N_8751,N_6852);
nand U11759 (N_11759,N_7272,N_7390);
or U11760 (N_11760,N_8519,N_9534);
xnor U11761 (N_11761,N_5659,N_7092);
and U11762 (N_11762,N_5115,N_7010);
nand U11763 (N_11763,N_6694,N_5836);
nor U11764 (N_11764,N_8864,N_6324);
nor U11765 (N_11765,N_6297,N_7527);
nor U11766 (N_11766,N_5159,N_5489);
nor U11767 (N_11767,N_6412,N_9969);
nor U11768 (N_11768,N_5441,N_8058);
nand U11769 (N_11769,N_5768,N_5262);
and U11770 (N_11770,N_6816,N_7659);
nor U11771 (N_11771,N_9747,N_8927);
or U11772 (N_11772,N_6173,N_9501);
nand U11773 (N_11773,N_9312,N_7473);
or U11774 (N_11774,N_7282,N_7388);
nor U11775 (N_11775,N_6280,N_9157);
nand U11776 (N_11776,N_9962,N_5646);
nand U11777 (N_11777,N_7874,N_9865);
or U11778 (N_11778,N_9013,N_7019);
nand U11779 (N_11779,N_8823,N_7339);
nand U11780 (N_11780,N_5384,N_5358);
or U11781 (N_11781,N_8302,N_7989);
nor U11782 (N_11782,N_9252,N_6805);
and U11783 (N_11783,N_9664,N_9864);
nor U11784 (N_11784,N_7515,N_5067);
nor U11785 (N_11785,N_6973,N_9685);
or U11786 (N_11786,N_7561,N_5974);
nand U11787 (N_11787,N_7616,N_5089);
and U11788 (N_11788,N_9175,N_8689);
nand U11789 (N_11789,N_9600,N_5006);
nor U11790 (N_11790,N_8552,N_7207);
nor U11791 (N_11791,N_8723,N_6377);
nand U11792 (N_11792,N_5208,N_6619);
or U11793 (N_11793,N_9315,N_6227);
nand U11794 (N_11794,N_5169,N_6017);
or U11795 (N_11795,N_7920,N_9826);
or U11796 (N_11796,N_8523,N_5852);
or U11797 (N_11797,N_9581,N_6452);
nand U11798 (N_11798,N_5502,N_7711);
and U11799 (N_11799,N_6609,N_7039);
or U11800 (N_11800,N_7428,N_8534);
nand U11801 (N_11801,N_5616,N_8691);
nand U11802 (N_11802,N_7756,N_7011);
nor U11803 (N_11803,N_6783,N_5777);
and U11804 (N_11804,N_6648,N_7636);
and U11805 (N_11805,N_5926,N_5582);
nor U11806 (N_11806,N_9075,N_8405);
nor U11807 (N_11807,N_6207,N_7347);
and U11808 (N_11808,N_8917,N_7631);
and U11809 (N_11809,N_6670,N_5199);
nand U11810 (N_11810,N_9180,N_9929);
nand U11811 (N_11811,N_9186,N_6997);
or U11812 (N_11812,N_9801,N_7931);
or U11813 (N_11813,N_7694,N_5523);
or U11814 (N_11814,N_6471,N_9375);
nand U11815 (N_11815,N_9197,N_8385);
or U11816 (N_11816,N_6354,N_6742);
nor U11817 (N_11817,N_7895,N_8981);
and U11818 (N_11818,N_5844,N_7979);
nand U11819 (N_11819,N_9271,N_5859);
and U11820 (N_11820,N_7262,N_5588);
and U11821 (N_11821,N_5392,N_7445);
and U11822 (N_11822,N_7699,N_8431);
nand U11823 (N_11823,N_7248,N_5318);
nand U11824 (N_11824,N_8881,N_6801);
nor U11825 (N_11825,N_9678,N_9643);
and U11826 (N_11826,N_6164,N_8018);
and U11827 (N_11827,N_5807,N_5891);
and U11828 (N_11828,N_7044,N_6248);
and U11829 (N_11829,N_7773,N_8275);
or U11830 (N_11830,N_8382,N_5633);
and U11831 (N_11831,N_6097,N_9796);
or U11832 (N_11832,N_7878,N_6309);
nor U11833 (N_11833,N_7956,N_9979);
xor U11834 (N_11834,N_9054,N_8616);
or U11835 (N_11835,N_8407,N_8975);
or U11836 (N_11836,N_5946,N_5456);
and U11837 (N_11837,N_6614,N_7187);
or U11838 (N_11838,N_9035,N_5504);
and U11839 (N_11839,N_5116,N_8573);
and U11840 (N_11840,N_8185,N_6043);
nor U11841 (N_11841,N_9598,N_9603);
or U11842 (N_11842,N_8926,N_8255);
nor U11843 (N_11843,N_8030,N_5303);
xor U11844 (N_11844,N_7574,N_8326);
and U11845 (N_11845,N_5161,N_6919);
and U11846 (N_11846,N_8948,N_9070);
or U11847 (N_11847,N_6118,N_6129);
and U11848 (N_11848,N_5496,N_8911);
or U11849 (N_11849,N_9766,N_5827);
or U11850 (N_11850,N_5232,N_7322);
nand U11851 (N_11851,N_7824,N_9442);
and U11852 (N_11852,N_7863,N_9699);
or U11853 (N_11853,N_9041,N_9986);
or U11854 (N_11854,N_5447,N_5233);
nand U11855 (N_11855,N_6625,N_5119);
nor U11856 (N_11856,N_8537,N_5516);
and U11857 (N_11857,N_8932,N_6980);
nor U11858 (N_11858,N_9256,N_8057);
or U11859 (N_11859,N_9132,N_8794);
nand U11860 (N_11860,N_8374,N_6290);
and U11861 (N_11861,N_8098,N_5530);
nor U11862 (N_11862,N_5835,N_8347);
or U11863 (N_11863,N_7546,N_8069);
or U11864 (N_11864,N_6926,N_7249);
and U11865 (N_11865,N_5540,N_9582);
nor U11866 (N_11866,N_6371,N_8077);
nand U11867 (N_11867,N_6726,N_5962);
and U11868 (N_11868,N_5498,N_7419);
nor U11869 (N_11869,N_5834,N_5845);
nor U11870 (N_11870,N_5469,N_8395);
nor U11871 (N_11871,N_6821,N_8635);
and U11872 (N_11872,N_8906,N_5698);
nand U11873 (N_11873,N_7430,N_6240);
nand U11874 (N_11874,N_8674,N_9572);
or U11875 (N_11875,N_7227,N_6434);
nand U11876 (N_11876,N_9905,N_7829);
and U11877 (N_11877,N_5551,N_9724);
and U11878 (N_11878,N_6457,N_5601);
and U11879 (N_11879,N_5950,N_8270);
and U11880 (N_11880,N_8799,N_7051);
or U11881 (N_11881,N_8872,N_7627);
nor U11882 (N_11882,N_7848,N_9382);
and U11883 (N_11883,N_9282,N_9162);
or U11884 (N_11884,N_9438,N_6845);
nand U11885 (N_11885,N_6491,N_7948);
nand U11886 (N_11886,N_7735,N_5238);
nor U11887 (N_11887,N_8865,N_6961);
or U11888 (N_11888,N_8313,N_8739);
nand U11889 (N_11889,N_9734,N_9824);
or U11890 (N_11890,N_5775,N_5555);
and U11891 (N_11891,N_8297,N_5331);
or U11892 (N_11892,N_8170,N_8009);
nor U11893 (N_11893,N_6050,N_6078);
nor U11894 (N_11894,N_7214,N_7672);
nand U11895 (N_11895,N_7394,N_9244);
nor U11896 (N_11896,N_6339,N_8585);
or U11897 (N_11897,N_6148,N_9449);
or U11898 (N_11898,N_5579,N_7870);
or U11899 (N_11899,N_6877,N_8013);
nor U11900 (N_11900,N_8752,N_6966);
and U11901 (N_11901,N_7168,N_6025);
nor U11902 (N_11902,N_9878,N_8814);
and U11903 (N_11903,N_9277,N_6770);
nand U11904 (N_11904,N_8711,N_7330);
nand U11905 (N_11905,N_8157,N_9404);
or U11906 (N_11906,N_6714,N_9153);
or U11907 (N_11907,N_9505,N_5176);
nor U11908 (N_11908,N_5979,N_7787);
and U11909 (N_11909,N_6285,N_9607);
or U11910 (N_11910,N_8944,N_8184);
nor U11911 (N_11911,N_7604,N_9192);
nor U11912 (N_11912,N_8274,N_7953);
and U11913 (N_11913,N_5326,N_6130);
xnor U11914 (N_11914,N_9792,N_7549);
and U11915 (N_11915,N_8845,N_6213);
xnor U11916 (N_11916,N_5380,N_5846);
nand U11917 (N_11917,N_6773,N_8437);
nor U11918 (N_11918,N_5340,N_9852);
or U11919 (N_11919,N_9227,N_9922);
nand U11920 (N_11920,N_8645,N_8708);
nand U11921 (N_11921,N_7335,N_7114);
and U11922 (N_11922,N_8682,N_8214);
and U11923 (N_11923,N_5383,N_5615);
nand U11924 (N_11924,N_9674,N_8695);
nand U11925 (N_11925,N_8047,N_8476);
or U11926 (N_11926,N_7275,N_5010);
or U11927 (N_11927,N_5497,N_7378);
or U11928 (N_11928,N_7507,N_8130);
or U11929 (N_11929,N_6768,N_8946);
and U11930 (N_11930,N_5602,N_9276);
nand U11931 (N_11931,N_9977,N_9999);
nor U11932 (N_11932,N_6870,N_7781);
or U11933 (N_11933,N_7078,N_7000);
nand U11934 (N_11934,N_6026,N_6460);
nor U11935 (N_11935,N_9602,N_7049);
nand U11936 (N_11936,N_7965,N_7710);
or U11937 (N_11937,N_6793,N_7558);
nor U11938 (N_11938,N_7074,N_9924);
nor U11939 (N_11939,N_7784,N_7235);
or U11940 (N_11940,N_9238,N_7635);
nor U11941 (N_11941,N_7907,N_8461);
xnor U11942 (N_11942,N_5652,N_8517);
or U11943 (N_11943,N_9627,N_8539);
nand U11944 (N_11944,N_7792,N_9137);
or U11945 (N_11945,N_7448,N_9078);
nand U11946 (N_11946,N_8570,N_9350);
and U11947 (N_11947,N_5751,N_5218);
nand U11948 (N_11948,N_5613,N_7918);
or U11949 (N_11949,N_5732,N_6525);
nand U11950 (N_11950,N_8632,N_5083);
or U11951 (N_11951,N_6218,N_6311);
nand U11952 (N_11952,N_5427,N_5486);
and U11953 (N_11953,N_7555,N_8955);
nand U11954 (N_11954,N_9222,N_7514);
nand U11955 (N_11955,N_9189,N_9838);
nor U11956 (N_11956,N_7456,N_9593);
nand U11957 (N_11957,N_8920,N_8873);
and U11958 (N_11958,N_7908,N_8150);
nand U11959 (N_11959,N_8417,N_6468);
nor U11960 (N_11960,N_6853,N_6231);
and U11961 (N_11961,N_9133,N_7793);
nor U11962 (N_11962,N_8594,N_8279);
nor U11963 (N_11963,N_9736,N_8432);
nor U11964 (N_11964,N_8516,N_7810);
nand U11965 (N_11965,N_5151,N_5357);
or U11966 (N_11966,N_8220,N_7212);
nor U11967 (N_11967,N_9554,N_6158);
nor U11968 (N_11968,N_9295,N_5396);
nand U11969 (N_11969,N_8675,N_8440);
and U11970 (N_11970,N_8195,N_6896);
and U11971 (N_11971,N_7136,N_9499);
nand U11972 (N_11972,N_9328,N_5729);
nor U11973 (N_11973,N_9220,N_8782);
or U11974 (N_11974,N_6063,N_8224);
nor U11975 (N_11975,N_9735,N_6839);
or U11976 (N_11976,N_7850,N_6000);
and U11977 (N_11977,N_5779,N_8227);
or U11978 (N_11978,N_5228,N_8862);
or U11979 (N_11979,N_9579,N_6868);
nor U11980 (N_11980,N_8450,N_7707);
nor U11981 (N_11981,N_7222,N_7846);
nor U11982 (N_11982,N_8193,N_8149);
nor U11983 (N_11983,N_8354,N_5032);
and U11984 (N_11984,N_9434,N_8804);
nand U11985 (N_11985,N_8791,N_7666);
nor U11986 (N_11986,N_9187,N_9166);
nor U11987 (N_11987,N_8869,N_5592);
and U11988 (N_11988,N_7242,N_5764);
nand U11989 (N_11989,N_9147,N_5662);
nor U11990 (N_11990,N_7446,N_8866);
and U11991 (N_11991,N_7263,N_9403);
nor U11992 (N_11992,N_7634,N_5375);
or U11993 (N_11993,N_9135,N_8795);
nor U11994 (N_11994,N_6072,N_6313);
nand U11995 (N_11995,N_8271,N_7876);
nor U11996 (N_11996,N_8401,N_7779);
nand U11997 (N_11997,N_5415,N_7269);
nand U11998 (N_11998,N_8531,N_8879);
or U11999 (N_11999,N_7100,N_8330);
nand U12000 (N_12000,N_5172,N_9519);
or U12001 (N_12001,N_6469,N_8342);
nor U12002 (N_12002,N_5566,N_7468);
and U12003 (N_12003,N_6172,N_6274);
nand U12004 (N_12004,N_9379,N_5719);
nor U12005 (N_12005,N_7906,N_7420);
and U12006 (N_12006,N_6617,N_5217);
and U12007 (N_12007,N_5075,N_9909);
nand U12008 (N_12008,N_9785,N_9031);
and U12009 (N_12009,N_6461,N_7518);
or U12010 (N_12010,N_8219,N_9084);
nand U12011 (N_12011,N_7429,N_5821);
nand U12012 (N_12012,N_6910,N_7348);
and U12013 (N_12013,N_7247,N_5120);
nand U12014 (N_12014,N_9076,N_5464);
nand U12015 (N_12015,N_7026,N_5506);
and U12016 (N_12016,N_9809,N_9116);
nand U12017 (N_12017,N_7785,N_8356);
nand U12018 (N_12018,N_5961,N_6606);
xor U12019 (N_12019,N_8158,N_5574);
nor U12020 (N_12020,N_9327,N_9573);
nor U12021 (N_12021,N_8169,N_6454);
nor U12022 (N_12022,N_6656,N_8288);
nor U12023 (N_12023,N_9262,N_5538);
nor U12024 (N_12024,N_8541,N_6222);
nand U12025 (N_12025,N_6611,N_9574);
nand U12026 (N_12026,N_6441,N_7052);
nor U12027 (N_12027,N_8306,N_5745);
nor U12028 (N_12028,N_9728,N_5864);
nor U12029 (N_12029,N_9213,N_9356);
or U12030 (N_12030,N_5830,N_5426);
nand U12031 (N_12031,N_5805,N_6690);
nand U12032 (N_12032,N_9294,N_9840);
or U12033 (N_12033,N_5780,N_6755);
and U12034 (N_12034,N_8441,N_5353);
nand U12035 (N_12035,N_7404,N_7050);
nand U12036 (N_12036,N_6584,N_6520);
or U12037 (N_12037,N_8136,N_9782);
and U12038 (N_12038,N_9445,N_7393);
or U12039 (N_12039,N_9326,N_6681);
and U12040 (N_12040,N_5103,N_5307);
nor U12041 (N_12041,N_6895,N_7302);
nor U12042 (N_12042,N_5542,N_9452);
nand U12043 (N_12043,N_5346,N_8070);
nand U12044 (N_12044,N_9829,N_9857);
and U12045 (N_12045,N_9351,N_7801);
or U12046 (N_12046,N_6506,N_7067);
and U12047 (N_12047,N_5220,N_9181);
and U12048 (N_12048,N_8063,N_7055);
nor U12049 (N_12049,N_5360,N_9387);
nor U12050 (N_12050,N_8486,N_7297);
or U12051 (N_12051,N_6253,N_6929);
and U12052 (N_12052,N_5480,N_6575);
and U12053 (N_12053,N_7358,N_6179);
nand U12054 (N_12054,N_6739,N_8349);
and U12055 (N_12055,N_9816,N_9205);
and U12056 (N_12056,N_6101,N_6597);
or U12057 (N_12057,N_5320,N_8028);
nand U12058 (N_12058,N_6122,N_7460);
or U12059 (N_12059,N_9671,N_6141);
nand U12060 (N_12060,N_7813,N_6817);
or U12061 (N_12061,N_6221,N_9850);
nor U12062 (N_12062,N_8597,N_6590);
and U12063 (N_12063,N_9450,N_7679);
nand U12064 (N_12064,N_5922,N_8511);
xnor U12065 (N_12065,N_5175,N_8012);
and U12066 (N_12066,N_7669,N_9068);
nor U12067 (N_12067,N_8177,N_5938);
or U12068 (N_12068,N_9637,N_5059);
nand U12069 (N_12069,N_5924,N_7159);
and U12070 (N_12070,N_8046,N_9615);
or U12071 (N_12071,N_8707,N_8643);
nand U12072 (N_12072,N_9555,N_6640);
and U12073 (N_12073,N_6699,N_9082);
nand U12074 (N_12074,N_8087,N_9689);
nand U12075 (N_12075,N_5423,N_6333);
nor U12076 (N_12076,N_7273,N_7416);
or U12077 (N_12077,N_6034,N_6830);
nor U12078 (N_12078,N_7946,N_7438);
or U12079 (N_12079,N_6001,N_6602);
or U12080 (N_12080,N_8790,N_6425);
nand U12081 (N_12081,N_8784,N_9677);
nand U12082 (N_12082,N_9278,N_7311);
or U12083 (N_12083,N_7239,N_9976);
or U12084 (N_12084,N_5996,N_5916);
and U12085 (N_12085,N_6955,N_7286);
or U12086 (N_12086,N_9814,N_7144);
and U12087 (N_12087,N_7209,N_8421);
nand U12088 (N_12088,N_7064,N_9837);
and U12089 (N_12089,N_9265,N_5440);
nand U12090 (N_12090,N_5040,N_9417);
or U12091 (N_12091,N_6201,N_9731);
or U12092 (N_12092,N_7898,N_8413);
and U12093 (N_12093,N_7786,N_7483);
xnor U12094 (N_12094,N_8940,N_9191);
nand U12095 (N_12095,N_6936,N_9397);
and U12096 (N_12096,N_7279,N_7037);
nor U12097 (N_12097,N_8891,N_5929);
nor U12098 (N_12098,N_7077,N_6893);
or U12099 (N_12099,N_7437,N_7400);
nand U12100 (N_12100,N_8408,N_8078);
and U12101 (N_12101,N_7373,N_8745);
nand U12102 (N_12102,N_7516,N_5137);
or U12103 (N_12103,N_9655,N_8296);
or U12104 (N_12104,N_9117,N_5227);
and U12105 (N_12105,N_9026,N_7683);
nor U12106 (N_12106,N_9433,N_9470);
nor U12107 (N_12107,N_8903,N_8688);
and U12108 (N_12108,N_7648,N_6134);
and U12109 (N_12109,N_7921,N_7256);
or U12110 (N_12110,N_8990,N_7237);
or U12111 (N_12111,N_5667,N_8015);
or U12112 (N_12112,N_6010,N_8178);
and U12113 (N_12113,N_8119,N_7278);
nand U12114 (N_12114,N_7467,N_8709);
or U12115 (N_12115,N_7875,N_5628);
nand U12116 (N_12116,N_8016,N_7769);
nand U12117 (N_12117,N_9732,N_5490);
nor U12118 (N_12118,N_6170,N_5832);
and U12119 (N_12119,N_7622,N_6368);
nor U12120 (N_12120,N_9897,N_7525);
and U12121 (N_12121,N_9136,N_6866);
and U12122 (N_12122,N_6264,N_7858);
nand U12123 (N_12123,N_8971,N_6420);
nor U12124 (N_12124,N_9170,N_7398);
nand U12125 (N_12125,N_9998,N_9456);
or U12126 (N_12126,N_6540,N_8660);
or U12127 (N_12127,N_6427,N_8277);
and U12128 (N_12128,N_7925,N_9723);
nor U12129 (N_12129,N_7977,N_6700);
and U12130 (N_12130,N_5420,N_6347);
nor U12131 (N_12131,N_5245,N_6015);
or U12132 (N_12132,N_6849,N_9201);
nor U12133 (N_12133,N_7585,N_6407);
nand U12134 (N_12134,N_6558,N_5121);
and U12135 (N_12135,N_5205,N_8131);
nand U12136 (N_12136,N_7333,N_7638);
and U12137 (N_12137,N_8061,N_7018);
and U12138 (N_12138,N_9306,N_6047);
nor U12139 (N_12139,N_7502,N_5831);
and U12140 (N_12140,N_9086,N_6600);
or U12141 (N_12141,N_6528,N_6137);
or U12142 (N_12142,N_6639,N_5858);
xor U12143 (N_12143,N_5947,N_5226);
and U12144 (N_12144,N_7746,N_5337);
nand U12145 (N_12145,N_5022,N_6126);
and U12146 (N_12146,N_7366,N_5474);
and U12147 (N_12147,N_8322,N_7891);
or U12148 (N_12148,N_5520,N_8536);
and U12149 (N_12149,N_7245,N_6735);
nor U12150 (N_12150,N_7267,N_9985);
or U12151 (N_12151,N_8102,N_7158);
or U12152 (N_12152,N_5515,N_6465);
or U12153 (N_12153,N_7140,N_7413);
nand U12154 (N_12154,N_8008,N_6419);
nor U12155 (N_12155,N_7794,N_7167);
nand U12156 (N_12156,N_8854,N_9174);
and U12157 (N_12157,N_7451,N_9844);
and U12158 (N_12158,N_6933,N_6924);
or U12159 (N_12159,N_7671,N_9937);
nor U12160 (N_12160,N_9051,N_5617);
or U12161 (N_12161,N_9526,N_5255);
nand U12162 (N_12162,N_7372,N_6987);
or U12163 (N_12163,N_8978,N_8530);
nor U12164 (N_12164,N_7195,N_6027);
nand U12165 (N_12165,N_9493,N_5181);
xnor U12166 (N_12166,N_8668,N_6544);
or U12167 (N_12167,N_7540,N_6474);
nand U12168 (N_12168,N_9103,N_5720);
nor U12169 (N_12169,N_8931,N_9451);
and U12170 (N_12170,N_9714,N_5036);
nand U12171 (N_12171,N_7537,N_7006);
nor U12172 (N_12172,N_7545,N_8567);
nand U12173 (N_12173,N_7403,N_5981);
or U12174 (N_12174,N_7132,N_5185);
nand U12175 (N_12175,N_9131,N_8143);
nand U12176 (N_12176,N_5559,N_8604);
or U12177 (N_12177,N_6695,N_5952);
nor U12178 (N_12178,N_6276,N_7500);
and U12179 (N_12179,N_8843,N_9339);
nor U12180 (N_12180,N_9525,N_6226);
nor U12181 (N_12181,N_5611,N_8465);
and U12182 (N_12182,N_9533,N_8956);
and U12183 (N_12183,N_6113,N_9066);
nor U12184 (N_12184,N_8508,N_8152);
nor U12185 (N_12185,N_5164,N_5018);
and U12186 (N_12186,N_6764,N_6336);
and U12187 (N_12187,N_8697,N_9023);
or U12188 (N_12188,N_9743,N_6116);
or U12189 (N_12189,N_7737,N_8231);
and U12190 (N_12190,N_6610,N_7839);
nand U12191 (N_12191,N_8378,N_9882);
nand U12192 (N_12192,N_7767,N_9758);
and U12193 (N_12193,N_5890,N_5842);
nand U12194 (N_12194,N_5965,N_9373);
nand U12195 (N_12195,N_5201,N_8742);
nand U12196 (N_12196,N_9466,N_8730);
nor U12197 (N_12197,N_7556,N_9684);
nand U12198 (N_12198,N_8339,N_6683);
and U12199 (N_12199,N_8052,N_9739);
or U12200 (N_12200,N_7301,N_8551);
and U12201 (N_12201,N_8839,N_6049);
nand U12202 (N_12202,N_6133,N_7837);
nand U12203 (N_12203,N_6235,N_7802);
and U12204 (N_12204,N_5695,N_8596);
nand U12205 (N_12205,N_5418,N_9656);
and U12206 (N_12206,N_8345,N_8109);
nor U12207 (N_12207,N_5203,N_8816);
nand U12208 (N_12208,N_6175,N_6728);
nand U12209 (N_12209,N_6652,N_5019);
nor U12210 (N_12210,N_9884,N_8383);
nand U12211 (N_12211,N_7324,N_6490);
nor U12212 (N_12212,N_6326,N_8902);
nor U12213 (N_12213,N_7122,N_7115);
and U12214 (N_12214,N_9853,N_9619);
and U12215 (N_12215,N_7524,N_8043);
nor U12216 (N_12216,N_6800,N_5572);
and U12217 (N_12217,N_6065,N_8398);
and U12218 (N_12218,N_5689,N_8448);
nor U12219 (N_12219,N_5740,N_6184);
nor U12220 (N_12220,N_5876,N_5584);
nor U12221 (N_12221,N_8989,N_9104);
or U12222 (N_12222,N_6950,N_6813);
and U12223 (N_12223,N_8889,N_6389);
nor U12224 (N_12224,N_6268,N_8605);
nor U12225 (N_12225,N_6325,N_9302);
and U12226 (N_12226,N_8694,N_8827);
nand U12227 (N_12227,N_8459,N_8365);
and U12228 (N_12228,N_8950,N_9443);
nand U12229 (N_12229,N_8621,N_6378);
nor U12230 (N_12230,N_8128,N_9712);
nand U12231 (N_12231,N_6555,N_8467);
and U12232 (N_12232,N_6380,N_8576);
and U12233 (N_12233,N_6601,N_6077);
nand U12234 (N_12234,N_9421,N_6289);
nor U12235 (N_12235,N_9997,N_7185);
or U12236 (N_12236,N_7606,N_7857);
nor U12237 (N_12237,N_6022,N_6331);
nand U12238 (N_12238,N_7402,N_9895);
or U12239 (N_12239,N_7397,N_6907);
and U12240 (N_12240,N_7193,N_6678);
nand U12241 (N_12241,N_6406,N_8282);
and U12242 (N_12242,N_8868,N_5388);
nand U12243 (N_12243,N_8416,N_8160);
or U12244 (N_12244,N_6395,N_9691);
or U12245 (N_12245,N_5369,N_7758);
nor U12246 (N_12246,N_9319,N_6291);
nand U12247 (N_12247,N_9040,N_8687);
and U12248 (N_12248,N_8145,N_9038);
nand U12249 (N_12249,N_6106,N_5082);
nor U12250 (N_12250,N_8729,N_6214);
nand U12251 (N_12251,N_7229,N_7625);
nand U12252 (N_12252,N_6599,N_5757);
and U12253 (N_12253,N_9152,N_7835);
and U12254 (N_12254,N_6591,N_7268);
or U12255 (N_12255,N_6161,N_5230);
or U12256 (N_12256,N_9547,N_6649);
or U12257 (N_12257,N_9718,N_6570);
nand U12258 (N_12258,N_5786,N_5818);
and U12259 (N_12259,N_9079,N_6232);
or U12260 (N_12260,N_9938,N_9773);
nor U12261 (N_12261,N_5149,N_7804);
nor U12262 (N_12262,N_5896,N_9567);
or U12263 (N_12263,N_9562,N_7733);
and U12264 (N_12264,N_7107,N_7411);
or U12265 (N_12265,N_7649,N_8101);
nor U12266 (N_12266,N_5957,N_5133);
nor U12267 (N_12267,N_8564,N_6476);
nor U12268 (N_12268,N_8146,N_7427);
and U12269 (N_12269,N_7033,N_5693);
nand U12270 (N_12270,N_5352,N_8699);
or U12271 (N_12271,N_6269,N_5927);
nor U12272 (N_12272,N_6445,N_8717);
nand U12273 (N_12273,N_9571,N_9584);
nor U12274 (N_12274,N_5446,N_5980);
nor U12275 (N_12275,N_7128,N_7831);
or U12276 (N_12276,N_6586,N_6338);
or U12277 (N_12277,N_7844,N_5647);
and U12278 (N_12278,N_7997,N_8363);
nand U12279 (N_12279,N_8386,N_5488);
nand U12280 (N_12280,N_8358,N_6542);
nor U12281 (N_12281,N_7457,N_9085);
or U12282 (N_12282,N_6505,N_8155);
nor U12283 (N_12283,N_7571,N_5868);
and U12284 (N_12284,N_5184,N_6659);
nor U12285 (N_12285,N_8829,N_8642);
nand U12286 (N_12286,N_6099,N_7866);
nor U12287 (N_12287,N_5005,N_5096);
nand U12288 (N_12288,N_7369,N_6809);
nor U12289 (N_12289,N_6417,N_8929);
or U12290 (N_12290,N_5222,N_9706);
and U12291 (N_12291,N_5413,N_9101);
nor U12292 (N_12292,N_9900,N_8725);
nand U12293 (N_12293,N_9018,N_9694);
and U12294 (N_12294,N_5122,N_7715);
or U12295 (N_12295,N_8818,N_7254);
or U12296 (N_12296,N_8951,N_6429);
nor U12297 (N_12297,N_7040,N_5031);
nor U12298 (N_12298,N_6477,N_5563);
or U12299 (N_12299,N_9733,N_7294);
nor U12300 (N_12300,N_5011,N_6502);
nor U12301 (N_12301,N_6978,N_5570);
nand U12302 (N_12302,N_8652,N_8261);
nor U12303 (N_12303,N_7926,N_5296);
nand U12304 (N_12304,N_8430,N_6589);
nor U12305 (N_12305,N_6272,N_7103);
and U12306 (N_12306,N_9123,N_5252);
nor U12307 (N_12307,N_8758,N_5746);
nand U12308 (N_12308,N_7552,N_5600);
nor U12309 (N_12309,N_8055,N_8805);
and U12310 (N_12310,N_7152,N_6305);
and U12311 (N_12311,N_9172,N_8039);
nand U12312 (N_12312,N_5444,N_7682);
nand U12313 (N_12313,N_6621,N_6921);
or U12314 (N_12314,N_8355,N_6824);
nand U12315 (N_12315,N_9273,N_6061);
nor U12316 (N_12316,N_6191,N_6551);
nor U12317 (N_12317,N_6947,N_5660);
and U12318 (N_12318,N_7484,N_8391);
nor U12319 (N_12319,N_8218,N_8394);
nor U12320 (N_12320,N_9638,N_9626);
or U12321 (N_12321,N_9159,N_5705);
and U12322 (N_12322,N_9830,N_5379);
nand U12323 (N_12323,N_7099,N_5912);
or U12324 (N_12324,N_6430,N_7617);
nor U12325 (N_12325,N_8934,N_9663);
nand U12326 (N_12326,N_5799,N_5473);
nand U12327 (N_12327,N_9813,N_9055);
and U12328 (N_12328,N_8882,N_5324);
nor U12329 (N_12329,N_7665,N_8305);
or U12330 (N_12330,N_6618,N_5060);
and U12331 (N_12331,N_7602,N_6697);
and U12332 (N_12332,N_6832,N_9721);
nor U12333 (N_12333,N_9037,N_8438);
nor U12334 (N_12334,N_5224,N_8041);
or U12335 (N_12335,N_8922,N_8653);
and U12336 (N_12336,N_7405,N_5409);
nor U12337 (N_12337,N_8728,N_9183);
nor U12338 (N_12338,N_8240,N_8153);
or U12339 (N_12339,N_7894,N_5774);
nand U12340 (N_12340,N_5552,N_7432);
or U12341 (N_12341,N_9774,N_7913);
nor U12342 (N_12342,N_9106,N_5294);
or U12343 (N_12343,N_5872,N_6651);
nor U12344 (N_12344,N_7797,N_8878);
nand U12345 (N_12345,N_9709,N_8659);
and U12346 (N_12346,N_5797,N_7123);
nor U12347 (N_12347,N_7884,N_8392);
nor U12348 (N_12348,N_5583,N_8640);
nor U12349 (N_12349,N_6644,N_7409);
or U12350 (N_12350,N_6638,N_5343);
or U12351 (N_12351,N_6234,N_7444);
nand U12352 (N_12352,N_8529,N_8939);
and U12353 (N_12353,N_7641,N_6881);
or U12354 (N_12354,N_6345,N_8904);
nor U12355 (N_12355,N_9228,N_9388);
or U12356 (N_12356,N_9396,N_5629);
or U12357 (N_12357,N_8821,N_6854);
nor U12358 (N_12358,N_8644,N_8104);
and U12359 (N_12359,N_9484,N_9542);
nor U12360 (N_12360,N_8634,N_8735);
nand U12361 (N_12361,N_5921,N_9577);
nor U12362 (N_12362,N_5772,N_7318);
nor U12363 (N_12363,N_9498,N_7310);
nor U12364 (N_12364,N_5966,N_7350);
nand U12365 (N_12365,N_9587,N_6123);
nand U12366 (N_12366,N_7418,N_8870);
nor U12367 (N_12367,N_7083,N_7329);
nor U12368 (N_12368,N_9479,N_6405);
or U12369 (N_12369,N_9246,N_6422);
nand U12370 (N_12370,N_6180,N_5675);
nor U12371 (N_12371,N_9713,N_5012);
nor U12372 (N_12372,N_5050,N_8785);
or U12373 (N_12373,N_6205,N_7772);
nand U12374 (N_12374,N_9823,N_8698);
nand U12375 (N_12375,N_7069,N_9297);
nor U12376 (N_12376,N_7827,N_8930);
nor U12377 (N_12377,N_9482,N_6013);
or U12378 (N_12378,N_7670,N_7131);
or U12379 (N_12379,N_9866,N_6952);
and U12380 (N_12380,N_8056,N_7485);
or U12381 (N_12381,N_9148,N_8860);
nand U12382 (N_12382,N_5910,N_5915);
nand U12383 (N_12383,N_6847,N_5681);
nor U12384 (N_12384,N_8116,N_8304);
and U12385 (N_12385,N_6653,N_5109);
nand U12386 (N_12386,N_9027,N_9391);
nor U12387 (N_12387,N_6628,N_7076);
xor U12388 (N_12388,N_9634,N_7933);
xor U12389 (N_12389,N_6418,N_8732);
nand U12390 (N_12390,N_7702,N_5690);
or U12391 (N_12391,N_7962,N_5043);
and U12392 (N_12392,N_8760,N_6661);
and U12393 (N_12393,N_6255,N_9232);
or U12394 (N_12394,N_6124,N_8084);
nand U12395 (N_12395,N_9352,N_9090);
nand U12396 (N_12396,N_8806,N_7363);
nor U12397 (N_12397,N_7629,N_6244);
nand U12398 (N_12398,N_5850,N_8887);
and U12399 (N_12399,N_9469,N_9354);
nor U12400 (N_12400,N_9726,N_7790);
nor U12401 (N_12401,N_9316,N_9941);
nor U12402 (N_12402,N_9150,N_9618);
nand U12403 (N_12403,N_8885,N_6580);
nand U12404 (N_12404,N_9589,N_7475);
and U12405 (N_12405,N_8373,N_6757);
and U12406 (N_12406,N_7399,N_5248);
and U12407 (N_12407,N_8662,N_6995);
or U12408 (N_12408,N_5071,N_9751);
nor U12409 (N_12409,N_6827,N_5771);
nor U12410 (N_12410,N_8025,N_6006);
nand U12411 (N_12411,N_6654,N_7520);
or U12412 (N_12412,N_5744,N_7202);
and U12413 (N_12413,N_6056,N_8221);
nand U12414 (N_12414,N_5973,N_8857);
or U12415 (N_12415,N_7650,N_7993);
nand U12416 (N_12416,N_9188,N_9576);
or U12417 (N_12417,N_8384,N_5560);
or U12418 (N_12418,N_8693,N_5897);
nor U12419 (N_12419,N_8890,N_7704);
nor U12420 (N_12420,N_5630,N_9003);
nand U12421 (N_12421,N_6746,N_6431);
and U12422 (N_12422,N_7509,N_6605);
or U12423 (N_12423,N_6504,N_6915);
nand U12424 (N_12424,N_9380,N_6679);
or U12425 (N_12425,N_7314,N_6480);
nand U12426 (N_12426,N_5399,N_7449);
nand U12427 (N_12427,N_8810,N_6428);
and U12428 (N_12428,N_7739,N_7090);
nand U12429 (N_12429,N_7748,N_7938);
nand U12430 (N_12430,N_8307,N_9357);
nand U12431 (N_12431,N_5347,N_6688);
nor U12432 (N_12432,N_6513,N_7323);
and U12433 (N_12433,N_9645,N_9502);
and U12434 (N_12434,N_5781,N_9118);
or U12435 (N_12435,N_8222,N_8493);
and U12436 (N_12436,N_7384,N_9597);
or U12437 (N_12437,N_9490,N_8840);
nor U12438 (N_12438,N_8204,N_6891);
nand U12439 (N_12439,N_8245,N_8983);
nor U12440 (N_12440,N_5345,N_8414);
and U12441 (N_12441,N_5435,N_5260);
and U12442 (N_12442,N_6259,N_5142);
nand U12443 (N_12443,N_9224,N_8703);
and U12444 (N_12444,N_6863,N_7296);
nand U12445 (N_12445,N_9740,N_6913);
nand U12446 (N_12446,N_7812,N_7124);
and U12447 (N_12447,N_9019,N_9819);
nand U12448 (N_12448,N_6286,N_9669);
or U12449 (N_12449,N_9144,N_6671);
and U12450 (N_12450,N_8900,N_6532);
nand U12451 (N_12451,N_8258,N_9513);
xnor U12452 (N_12452,N_8710,N_6790);
nand U12453 (N_12453,N_6569,N_8471);
and U12454 (N_12454,N_8679,N_9661);
nor U12455 (N_12455,N_7382,N_5401);
nand U12456 (N_12456,N_9749,N_5319);
nand U12457 (N_12457,N_8671,N_9145);
and U12458 (N_12458,N_5935,N_6571);
nor U12459 (N_12459,N_5971,N_5285);
or U12460 (N_12460,N_5666,N_7289);
and U12461 (N_12461,N_8562,N_5125);
nand U12462 (N_12462,N_5898,N_7886);
nor U12463 (N_12463,N_7820,N_8125);
and U12464 (N_12464,N_5534,N_7919);
nor U12465 (N_12465,N_8650,N_5088);
or U12466 (N_12466,N_5663,N_9667);
nand U12467 (N_12467,N_5066,N_9266);
nor U12468 (N_12468,N_6914,N_5585);
or U12469 (N_12469,N_7619,N_9887);
nand U12470 (N_12470,N_9649,N_6104);
nor U12471 (N_12471,N_5510,N_7291);
nor U12472 (N_12472,N_9833,N_6596);
and U12473 (N_12473,N_5581,N_5909);
nor U12474 (N_12474,N_5828,N_9874);
or U12475 (N_12475,N_7959,N_7141);
nand U12476 (N_12476,N_8298,N_7970);
or U12477 (N_12477,N_7557,N_5734);
and U12478 (N_12478,N_8248,N_5716);
nand U12479 (N_12479,N_5591,N_7952);
nand U12480 (N_12480,N_9324,N_5725);
and U12481 (N_12481,N_5465,N_5999);
or U12482 (N_12482,N_6037,N_8587);
xnor U12483 (N_12483,N_8415,N_7196);
nor U12484 (N_12484,N_8403,N_5547);
nand U12485 (N_12485,N_5990,N_9557);
nand U12486 (N_12486,N_6067,N_8262);
nand U12487 (N_12487,N_9545,N_6308);
or U12488 (N_12488,N_7236,N_8457);
nand U12489 (N_12489,N_7588,N_5770);
and U12490 (N_12490,N_7904,N_6546);
or U12491 (N_12491,N_5235,N_7662);
and U12492 (N_12492,N_5376,N_7230);
and U12493 (N_12493,N_9007,N_6550);
and U12494 (N_12494,N_9926,N_7759);
or U12495 (N_12495,N_5148,N_7022);
nor U12496 (N_12496,N_6772,N_5007);
nor U12497 (N_12497,N_7464,N_8755);
and U12498 (N_12498,N_6411,N_8719);
or U12499 (N_12499,N_9789,N_9322);
xnor U12500 (N_12500,N_5340,N_5673);
and U12501 (N_12501,N_6285,N_5813);
or U12502 (N_12502,N_5554,N_7396);
nand U12503 (N_12503,N_9369,N_6342);
and U12504 (N_12504,N_5078,N_9597);
nor U12505 (N_12505,N_7633,N_8346);
and U12506 (N_12506,N_7556,N_6126);
and U12507 (N_12507,N_5165,N_6327);
nand U12508 (N_12508,N_6695,N_6769);
or U12509 (N_12509,N_8312,N_9198);
and U12510 (N_12510,N_9701,N_8324);
nand U12511 (N_12511,N_6465,N_5211);
and U12512 (N_12512,N_8070,N_8190);
nor U12513 (N_12513,N_8900,N_6467);
and U12514 (N_12514,N_5757,N_9936);
and U12515 (N_12515,N_7129,N_6177);
nor U12516 (N_12516,N_8117,N_6954);
nand U12517 (N_12517,N_9000,N_5070);
and U12518 (N_12518,N_6879,N_7536);
or U12519 (N_12519,N_5096,N_6235);
nand U12520 (N_12520,N_6004,N_6644);
and U12521 (N_12521,N_6589,N_7470);
nand U12522 (N_12522,N_7717,N_6938);
nand U12523 (N_12523,N_7449,N_7163);
and U12524 (N_12524,N_8230,N_9689);
and U12525 (N_12525,N_7300,N_6670);
and U12526 (N_12526,N_6187,N_7936);
and U12527 (N_12527,N_9833,N_8651);
or U12528 (N_12528,N_8239,N_9273);
and U12529 (N_12529,N_9148,N_7482);
nor U12530 (N_12530,N_6964,N_9344);
and U12531 (N_12531,N_7994,N_6500);
or U12532 (N_12532,N_6181,N_5523);
or U12533 (N_12533,N_7671,N_5776);
or U12534 (N_12534,N_7659,N_7713);
and U12535 (N_12535,N_8109,N_9010);
and U12536 (N_12536,N_5613,N_6103);
or U12537 (N_12537,N_7898,N_9872);
or U12538 (N_12538,N_7288,N_9385);
or U12539 (N_12539,N_6937,N_8797);
nand U12540 (N_12540,N_5690,N_7170);
nor U12541 (N_12541,N_8705,N_5730);
and U12542 (N_12542,N_8178,N_6145);
or U12543 (N_12543,N_9813,N_9494);
nor U12544 (N_12544,N_8819,N_5679);
or U12545 (N_12545,N_9111,N_7838);
nand U12546 (N_12546,N_8064,N_8091);
nand U12547 (N_12547,N_5324,N_7933);
or U12548 (N_12548,N_7526,N_9587);
nand U12549 (N_12549,N_6902,N_5221);
and U12550 (N_12550,N_9222,N_6871);
or U12551 (N_12551,N_6203,N_7160);
nor U12552 (N_12552,N_7541,N_6557);
nor U12553 (N_12553,N_6803,N_6301);
nand U12554 (N_12554,N_7247,N_7401);
nor U12555 (N_12555,N_8032,N_8310);
nor U12556 (N_12556,N_6325,N_7923);
nand U12557 (N_12557,N_5957,N_5665);
and U12558 (N_12558,N_5933,N_7146);
nor U12559 (N_12559,N_7337,N_8214);
nand U12560 (N_12560,N_7391,N_5386);
or U12561 (N_12561,N_9759,N_6417);
nor U12562 (N_12562,N_9004,N_7295);
nand U12563 (N_12563,N_6321,N_9822);
nor U12564 (N_12564,N_5067,N_9694);
or U12565 (N_12565,N_6889,N_5603);
nand U12566 (N_12566,N_7085,N_7889);
nand U12567 (N_12567,N_9763,N_9728);
nand U12568 (N_12568,N_6168,N_5146);
and U12569 (N_12569,N_5485,N_8868);
or U12570 (N_12570,N_9981,N_9368);
nor U12571 (N_12571,N_9364,N_8019);
or U12572 (N_12572,N_5833,N_7850);
and U12573 (N_12573,N_8168,N_7153);
nor U12574 (N_12574,N_7771,N_7694);
nor U12575 (N_12575,N_8945,N_9506);
nand U12576 (N_12576,N_6443,N_6770);
and U12577 (N_12577,N_9382,N_9009);
and U12578 (N_12578,N_5526,N_7677);
and U12579 (N_12579,N_6886,N_9960);
nand U12580 (N_12580,N_6651,N_9252);
nor U12581 (N_12581,N_6296,N_7231);
nand U12582 (N_12582,N_9284,N_9566);
nand U12583 (N_12583,N_7697,N_6111);
or U12584 (N_12584,N_6162,N_9683);
and U12585 (N_12585,N_8531,N_6448);
or U12586 (N_12586,N_5928,N_9507);
and U12587 (N_12587,N_9881,N_9831);
nor U12588 (N_12588,N_8357,N_8252);
nand U12589 (N_12589,N_9968,N_8517);
nand U12590 (N_12590,N_8390,N_8491);
or U12591 (N_12591,N_9667,N_6837);
or U12592 (N_12592,N_9102,N_7277);
or U12593 (N_12593,N_8640,N_9350);
and U12594 (N_12594,N_6353,N_8673);
and U12595 (N_12595,N_7586,N_8174);
nor U12596 (N_12596,N_5566,N_7098);
nand U12597 (N_12597,N_7016,N_8056);
or U12598 (N_12598,N_6851,N_7551);
nor U12599 (N_12599,N_6333,N_5507);
or U12600 (N_12600,N_8593,N_8173);
nand U12601 (N_12601,N_9557,N_7670);
or U12602 (N_12602,N_9970,N_7449);
nor U12603 (N_12603,N_9850,N_6801);
or U12604 (N_12604,N_6529,N_5473);
nor U12605 (N_12605,N_7315,N_6404);
and U12606 (N_12606,N_6414,N_6462);
and U12607 (N_12607,N_5600,N_9758);
nor U12608 (N_12608,N_5185,N_7366);
or U12609 (N_12609,N_9056,N_8814);
nor U12610 (N_12610,N_9939,N_8612);
or U12611 (N_12611,N_6949,N_5743);
nand U12612 (N_12612,N_9916,N_7729);
nand U12613 (N_12613,N_9193,N_9262);
or U12614 (N_12614,N_7689,N_6811);
nand U12615 (N_12615,N_8920,N_8413);
nand U12616 (N_12616,N_9917,N_8203);
nor U12617 (N_12617,N_5409,N_9875);
and U12618 (N_12618,N_9822,N_8134);
or U12619 (N_12619,N_5278,N_5558);
or U12620 (N_12620,N_9921,N_8876);
and U12621 (N_12621,N_8378,N_7543);
nand U12622 (N_12622,N_7900,N_8354);
or U12623 (N_12623,N_6916,N_9451);
nor U12624 (N_12624,N_6742,N_6852);
nor U12625 (N_12625,N_8232,N_7466);
nand U12626 (N_12626,N_9503,N_5517);
or U12627 (N_12627,N_8273,N_6266);
or U12628 (N_12628,N_9866,N_7300);
or U12629 (N_12629,N_6190,N_6342);
nand U12630 (N_12630,N_9339,N_6423);
nor U12631 (N_12631,N_7359,N_8976);
nor U12632 (N_12632,N_5957,N_9541);
nand U12633 (N_12633,N_7090,N_5535);
and U12634 (N_12634,N_6287,N_5146);
nor U12635 (N_12635,N_8899,N_7935);
nor U12636 (N_12636,N_8647,N_6351);
xnor U12637 (N_12637,N_7119,N_7539);
and U12638 (N_12638,N_7806,N_5835);
nor U12639 (N_12639,N_8552,N_5694);
nor U12640 (N_12640,N_7030,N_6055);
nand U12641 (N_12641,N_8431,N_5268);
nand U12642 (N_12642,N_8385,N_7638);
or U12643 (N_12643,N_9475,N_6576);
and U12644 (N_12644,N_8536,N_5556);
and U12645 (N_12645,N_7153,N_8268);
nor U12646 (N_12646,N_9256,N_5487);
nand U12647 (N_12647,N_6649,N_5262);
nand U12648 (N_12648,N_7606,N_5454);
and U12649 (N_12649,N_9313,N_5237);
nor U12650 (N_12650,N_6986,N_6455);
nor U12651 (N_12651,N_7667,N_7184);
or U12652 (N_12652,N_7768,N_7332);
nand U12653 (N_12653,N_8393,N_5124);
nand U12654 (N_12654,N_9976,N_8607);
nor U12655 (N_12655,N_8694,N_7285);
and U12656 (N_12656,N_9271,N_8074);
nor U12657 (N_12657,N_7917,N_9384);
nor U12658 (N_12658,N_9554,N_8553);
nand U12659 (N_12659,N_6973,N_6199);
nor U12660 (N_12660,N_7848,N_5719);
or U12661 (N_12661,N_6351,N_7143);
or U12662 (N_12662,N_5827,N_7183);
nor U12663 (N_12663,N_8993,N_8984);
and U12664 (N_12664,N_8192,N_6628);
nand U12665 (N_12665,N_9099,N_6022);
nor U12666 (N_12666,N_8990,N_9926);
nand U12667 (N_12667,N_7962,N_8420);
nand U12668 (N_12668,N_5614,N_9254);
or U12669 (N_12669,N_9498,N_6981);
nand U12670 (N_12670,N_5852,N_9670);
and U12671 (N_12671,N_6474,N_9741);
and U12672 (N_12672,N_5479,N_6745);
or U12673 (N_12673,N_9812,N_9834);
or U12674 (N_12674,N_9415,N_9183);
and U12675 (N_12675,N_8121,N_6103);
and U12676 (N_12676,N_8692,N_6812);
nor U12677 (N_12677,N_6976,N_9085);
and U12678 (N_12678,N_7855,N_7417);
nor U12679 (N_12679,N_8942,N_9634);
nand U12680 (N_12680,N_9808,N_7787);
nand U12681 (N_12681,N_9560,N_8852);
nor U12682 (N_12682,N_9796,N_5371);
nand U12683 (N_12683,N_5842,N_5805);
nand U12684 (N_12684,N_8333,N_9963);
nand U12685 (N_12685,N_6627,N_6792);
nor U12686 (N_12686,N_5300,N_8597);
or U12687 (N_12687,N_6071,N_7752);
nor U12688 (N_12688,N_5999,N_7844);
nand U12689 (N_12689,N_9835,N_8022);
and U12690 (N_12690,N_6279,N_8727);
or U12691 (N_12691,N_7986,N_6751);
or U12692 (N_12692,N_7162,N_8669);
or U12693 (N_12693,N_6107,N_5643);
or U12694 (N_12694,N_5868,N_8625);
nor U12695 (N_12695,N_6052,N_7193);
or U12696 (N_12696,N_9780,N_6977);
or U12697 (N_12697,N_6578,N_5396);
nor U12698 (N_12698,N_8272,N_5595);
nand U12699 (N_12699,N_5711,N_6230);
nand U12700 (N_12700,N_9922,N_6091);
nor U12701 (N_12701,N_5200,N_5190);
nor U12702 (N_12702,N_9814,N_8535);
nor U12703 (N_12703,N_9781,N_5259);
nand U12704 (N_12704,N_5623,N_7622);
and U12705 (N_12705,N_8517,N_8717);
and U12706 (N_12706,N_6314,N_8078);
and U12707 (N_12707,N_8401,N_6119);
or U12708 (N_12708,N_9969,N_6488);
and U12709 (N_12709,N_6089,N_6784);
and U12710 (N_12710,N_6549,N_5688);
and U12711 (N_12711,N_9306,N_6145);
nor U12712 (N_12712,N_7403,N_7247);
nor U12713 (N_12713,N_5929,N_7870);
nor U12714 (N_12714,N_8677,N_5610);
nor U12715 (N_12715,N_9134,N_8040);
nand U12716 (N_12716,N_9660,N_8768);
and U12717 (N_12717,N_5336,N_9486);
or U12718 (N_12718,N_9269,N_7635);
and U12719 (N_12719,N_6198,N_5768);
and U12720 (N_12720,N_9001,N_5092);
nand U12721 (N_12721,N_7932,N_8264);
and U12722 (N_12722,N_9503,N_9511);
nand U12723 (N_12723,N_8345,N_8274);
and U12724 (N_12724,N_5897,N_8383);
or U12725 (N_12725,N_6377,N_9163);
nand U12726 (N_12726,N_8608,N_7834);
and U12727 (N_12727,N_7555,N_8470);
or U12728 (N_12728,N_7880,N_5691);
or U12729 (N_12729,N_5054,N_6059);
and U12730 (N_12730,N_9262,N_9342);
or U12731 (N_12731,N_8767,N_9299);
or U12732 (N_12732,N_9400,N_8648);
or U12733 (N_12733,N_8588,N_8555);
nand U12734 (N_12734,N_6964,N_8422);
nand U12735 (N_12735,N_8965,N_8834);
nor U12736 (N_12736,N_9399,N_9127);
nand U12737 (N_12737,N_8653,N_7974);
or U12738 (N_12738,N_6085,N_8462);
nand U12739 (N_12739,N_9819,N_7863);
and U12740 (N_12740,N_5956,N_5907);
and U12741 (N_12741,N_8884,N_5058);
nor U12742 (N_12742,N_8834,N_9219);
or U12743 (N_12743,N_9760,N_6715);
nor U12744 (N_12744,N_7653,N_9192);
or U12745 (N_12745,N_9930,N_6324);
nor U12746 (N_12746,N_5081,N_6872);
nand U12747 (N_12747,N_8603,N_8303);
nor U12748 (N_12748,N_9042,N_6513);
and U12749 (N_12749,N_8083,N_7085);
nor U12750 (N_12750,N_5947,N_9556);
nand U12751 (N_12751,N_8144,N_8729);
nand U12752 (N_12752,N_8328,N_9820);
or U12753 (N_12753,N_7867,N_9843);
nand U12754 (N_12754,N_8705,N_5319);
nor U12755 (N_12755,N_8886,N_7022);
and U12756 (N_12756,N_6899,N_6290);
nand U12757 (N_12757,N_5764,N_6479);
nand U12758 (N_12758,N_9660,N_7176);
nor U12759 (N_12759,N_5012,N_8965);
nand U12760 (N_12760,N_5712,N_5136);
nor U12761 (N_12761,N_7847,N_6168);
nand U12762 (N_12762,N_6408,N_9330);
nand U12763 (N_12763,N_6305,N_7915);
nand U12764 (N_12764,N_5532,N_6785);
and U12765 (N_12765,N_8605,N_9315);
and U12766 (N_12766,N_9523,N_6581);
nor U12767 (N_12767,N_6356,N_7207);
nand U12768 (N_12768,N_5858,N_8761);
nor U12769 (N_12769,N_9582,N_6764);
or U12770 (N_12770,N_9959,N_7164);
and U12771 (N_12771,N_8491,N_7619);
or U12772 (N_12772,N_9422,N_6473);
and U12773 (N_12773,N_7071,N_8119);
nand U12774 (N_12774,N_6895,N_8723);
nor U12775 (N_12775,N_8395,N_6845);
and U12776 (N_12776,N_5636,N_6894);
nand U12777 (N_12777,N_7649,N_9920);
nor U12778 (N_12778,N_6000,N_8675);
nand U12779 (N_12779,N_5482,N_8224);
nand U12780 (N_12780,N_7646,N_8718);
and U12781 (N_12781,N_8032,N_7351);
and U12782 (N_12782,N_6831,N_6817);
nand U12783 (N_12783,N_8343,N_6012);
or U12784 (N_12784,N_7329,N_9135);
or U12785 (N_12785,N_8991,N_8612);
or U12786 (N_12786,N_9510,N_9488);
nand U12787 (N_12787,N_5319,N_5822);
nand U12788 (N_12788,N_7930,N_7378);
and U12789 (N_12789,N_8201,N_5790);
nor U12790 (N_12790,N_8107,N_6781);
and U12791 (N_12791,N_6078,N_7859);
nand U12792 (N_12792,N_5410,N_8852);
nor U12793 (N_12793,N_5027,N_8715);
and U12794 (N_12794,N_7812,N_7521);
and U12795 (N_12795,N_6976,N_6736);
or U12796 (N_12796,N_7589,N_6574);
or U12797 (N_12797,N_5500,N_7017);
nand U12798 (N_12798,N_8396,N_9995);
nand U12799 (N_12799,N_8017,N_8432);
nor U12800 (N_12800,N_8176,N_9629);
nand U12801 (N_12801,N_5030,N_5763);
nand U12802 (N_12802,N_7476,N_6108);
nor U12803 (N_12803,N_8301,N_9198);
or U12804 (N_12804,N_6994,N_6223);
nand U12805 (N_12805,N_5973,N_6227);
and U12806 (N_12806,N_5612,N_9729);
nor U12807 (N_12807,N_9601,N_8028);
and U12808 (N_12808,N_7480,N_8379);
and U12809 (N_12809,N_7255,N_5026);
nor U12810 (N_12810,N_7781,N_6169);
or U12811 (N_12811,N_7127,N_5263);
or U12812 (N_12812,N_9835,N_8208);
nand U12813 (N_12813,N_8235,N_5481);
or U12814 (N_12814,N_5800,N_6245);
and U12815 (N_12815,N_5877,N_9766);
nor U12816 (N_12816,N_8316,N_5518);
nor U12817 (N_12817,N_5334,N_8216);
nor U12818 (N_12818,N_8931,N_8466);
nand U12819 (N_12819,N_9877,N_5599);
nand U12820 (N_12820,N_8035,N_7721);
and U12821 (N_12821,N_7142,N_7139);
and U12822 (N_12822,N_8919,N_9761);
nand U12823 (N_12823,N_7589,N_5000);
or U12824 (N_12824,N_5991,N_6692);
nor U12825 (N_12825,N_6685,N_7465);
or U12826 (N_12826,N_6931,N_7744);
and U12827 (N_12827,N_5895,N_9394);
and U12828 (N_12828,N_8854,N_7782);
and U12829 (N_12829,N_8470,N_5342);
nand U12830 (N_12830,N_8024,N_8098);
nor U12831 (N_12831,N_9062,N_8743);
nand U12832 (N_12832,N_8321,N_7765);
nand U12833 (N_12833,N_7687,N_5460);
nor U12834 (N_12834,N_9867,N_8344);
nand U12835 (N_12835,N_9733,N_8133);
or U12836 (N_12836,N_5615,N_8787);
nand U12837 (N_12837,N_7292,N_9474);
and U12838 (N_12838,N_6633,N_8631);
or U12839 (N_12839,N_6138,N_7574);
nor U12840 (N_12840,N_9368,N_8539);
nor U12841 (N_12841,N_8747,N_9121);
and U12842 (N_12842,N_7517,N_6241);
nand U12843 (N_12843,N_5318,N_9481);
and U12844 (N_12844,N_5231,N_8847);
nand U12845 (N_12845,N_7862,N_9584);
or U12846 (N_12846,N_6794,N_5685);
and U12847 (N_12847,N_5597,N_7432);
nand U12848 (N_12848,N_5236,N_6233);
and U12849 (N_12849,N_8841,N_7377);
and U12850 (N_12850,N_7643,N_6835);
and U12851 (N_12851,N_5058,N_7452);
and U12852 (N_12852,N_6795,N_8135);
and U12853 (N_12853,N_6575,N_5974);
and U12854 (N_12854,N_5736,N_5263);
nor U12855 (N_12855,N_9367,N_5008);
or U12856 (N_12856,N_5675,N_9185);
nand U12857 (N_12857,N_6985,N_9807);
nor U12858 (N_12858,N_7873,N_5507);
nand U12859 (N_12859,N_8677,N_9062);
nor U12860 (N_12860,N_7920,N_6112);
or U12861 (N_12861,N_7171,N_9959);
and U12862 (N_12862,N_6325,N_8480);
nand U12863 (N_12863,N_9463,N_8216);
or U12864 (N_12864,N_5726,N_6209);
or U12865 (N_12865,N_6025,N_9749);
or U12866 (N_12866,N_6446,N_6752);
nor U12867 (N_12867,N_7118,N_6404);
nand U12868 (N_12868,N_8730,N_9084);
and U12869 (N_12869,N_7218,N_7263);
or U12870 (N_12870,N_8000,N_7437);
xor U12871 (N_12871,N_9452,N_8892);
and U12872 (N_12872,N_6194,N_8871);
nor U12873 (N_12873,N_8810,N_5414);
xnor U12874 (N_12874,N_8154,N_6883);
nor U12875 (N_12875,N_8473,N_9998);
or U12876 (N_12876,N_5539,N_5010);
or U12877 (N_12877,N_8734,N_5986);
and U12878 (N_12878,N_7776,N_9258);
nand U12879 (N_12879,N_8726,N_7188);
or U12880 (N_12880,N_7255,N_6540);
and U12881 (N_12881,N_6142,N_6385);
and U12882 (N_12882,N_8095,N_9497);
xnor U12883 (N_12883,N_7312,N_8663);
or U12884 (N_12884,N_5944,N_6487);
or U12885 (N_12885,N_7229,N_7652);
nand U12886 (N_12886,N_7162,N_5230);
or U12887 (N_12887,N_6654,N_8969);
nand U12888 (N_12888,N_6744,N_5486);
or U12889 (N_12889,N_5231,N_5910);
or U12890 (N_12890,N_9584,N_8138);
or U12891 (N_12891,N_6462,N_5486);
or U12892 (N_12892,N_6344,N_7857);
and U12893 (N_12893,N_9996,N_7137);
nand U12894 (N_12894,N_8792,N_5692);
and U12895 (N_12895,N_7207,N_9802);
nand U12896 (N_12896,N_6803,N_7915);
and U12897 (N_12897,N_7223,N_8187);
nor U12898 (N_12898,N_9551,N_8211);
nor U12899 (N_12899,N_5296,N_5314);
or U12900 (N_12900,N_7571,N_5561);
nor U12901 (N_12901,N_8698,N_9625);
nor U12902 (N_12902,N_5470,N_7376);
nor U12903 (N_12903,N_8937,N_8816);
nor U12904 (N_12904,N_7410,N_5403);
and U12905 (N_12905,N_9741,N_8029);
and U12906 (N_12906,N_6442,N_5757);
nor U12907 (N_12907,N_5887,N_8579);
or U12908 (N_12908,N_5952,N_7895);
nand U12909 (N_12909,N_6662,N_5092);
or U12910 (N_12910,N_9142,N_9032);
or U12911 (N_12911,N_6623,N_9077);
nor U12912 (N_12912,N_6076,N_9046);
nand U12913 (N_12913,N_7309,N_5676);
or U12914 (N_12914,N_6193,N_5203);
nor U12915 (N_12915,N_6895,N_9246);
nand U12916 (N_12916,N_7378,N_8995);
and U12917 (N_12917,N_6433,N_5722);
and U12918 (N_12918,N_8806,N_8300);
and U12919 (N_12919,N_5055,N_9217);
nand U12920 (N_12920,N_6748,N_5201);
or U12921 (N_12921,N_9444,N_6916);
or U12922 (N_12922,N_7486,N_5039);
nor U12923 (N_12923,N_8488,N_9977);
nand U12924 (N_12924,N_7357,N_8960);
and U12925 (N_12925,N_7376,N_7962);
or U12926 (N_12926,N_5002,N_9872);
or U12927 (N_12927,N_8203,N_5810);
nor U12928 (N_12928,N_9185,N_8520);
nand U12929 (N_12929,N_5238,N_9857);
or U12930 (N_12930,N_9431,N_7507);
nor U12931 (N_12931,N_5771,N_7809);
nor U12932 (N_12932,N_8187,N_6366);
nor U12933 (N_12933,N_6139,N_5750);
nor U12934 (N_12934,N_6308,N_7501);
nor U12935 (N_12935,N_5587,N_9319);
and U12936 (N_12936,N_9756,N_5519);
nand U12937 (N_12937,N_5606,N_8187);
nand U12938 (N_12938,N_7674,N_6151);
and U12939 (N_12939,N_6845,N_8374);
and U12940 (N_12940,N_8821,N_9139);
or U12941 (N_12941,N_7361,N_5506);
nor U12942 (N_12942,N_6485,N_5525);
nor U12943 (N_12943,N_7463,N_8863);
or U12944 (N_12944,N_9887,N_8719);
and U12945 (N_12945,N_6104,N_6162);
nand U12946 (N_12946,N_6917,N_9658);
nor U12947 (N_12947,N_5400,N_9363);
or U12948 (N_12948,N_6889,N_8868);
nand U12949 (N_12949,N_6532,N_7720);
and U12950 (N_12950,N_6681,N_7763);
nor U12951 (N_12951,N_9056,N_6550);
nor U12952 (N_12952,N_5088,N_6936);
or U12953 (N_12953,N_8651,N_6434);
and U12954 (N_12954,N_6201,N_7390);
and U12955 (N_12955,N_5230,N_7633);
nand U12956 (N_12956,N_6320,N_5643);
and U12957 (N_12957,N_8459,N_8390);
and U12958 (N_12958,N_6270,N_9957);
xor U12959 (N_12959,N_7952,N_9610);
and U12960 (N_12960,N_7363,N_6367);
and U12961 (N_12961,N_6927,N_5742);
nor U12962 (N_12962,N_7041,N_5274);
and U12963 (N_12963,N_9478,N_9784);
nand U12964 (N_12964,N_6957,N_6333);
and U12965 (N_12965,N_8112,N_9890);
nor U12966 (N_12966,N_5471,N_7948);
nand U12967 (N_12967,N_9530,N_6206);
nor U12968 (N_12968,N_8145,N_8657);
or U12969 (N_12969,N_8631,N_8518);
nand U12970 (N_12970,N_7214,N_9559);
and U12971 (N_12971,N_6096,N_5214);
and U12972 (N_12972,N_7589,N_9703);
and U12973 (N_12973,N_8926,N_8558);
and U12974 (N_12974,N_7277,N_6555);
nand U12975 (N_12975,N_8277,N_8476);
nand U12976 (N_12976,N_5492,N_5627);
and U12977 (N_12977,N_5079,N_5900);
nand U12978 (N_12978,N_5457,N_6913);
or U12979 (N_12979,N_5559,N_5788);
nand U12980 (N_12980,N_9526,N_5734);
and U12981 (N_12981,N_8655,N_9742);
or U12982 (N_12982,N_5471,N_9334);
and U12983 (N_12983,N_7868,N_5239);
or U12984 (N_12984,N_9531,N_5360);
and U12985 (N_12985,N_7419,N_6023);
nor U12986 (N_12986,N_6790,N_9275);
and U12987 (N_12987,N_5296,N_7030);
nand U12988 (N_12988,N_7556,N_7966);
nor U12989 (N_12989,N_9328,N_5616);
nand U12990 (N_12990,N_6669,N_7726);
nor U12991 (N_12991,N_5535,N_5306);
nor U12992 (N_12992,N_8761,N_5296);
and U12993 (N_12993,N_5439,N_5277);
and U12994 (N_12994,N_6337,N_7501);
nand U12995 (N_12995,N_5727,N_5795);
nor U12996 (N_12996,N_6450,N_5931);
nand U12997 (N_12997,N_8152,N_7090);
xor U12998 (N_12998,N_9123,N_6845);
and U12999 (N_12999,N_6435,N_6128);
or U13000 (N_13000,N_8165,N_6272);
and U13001 (N_13001,N_6619,N_5125);
nand U13002 (N_13002,N_5728,N_6222);
nand U13003 (N_13003,N_7095,N_8338);
nand U13004 (N_13004,N_5464,N_8825);
nor U13005 (N_13005,N_7563,N_8782);
and U13006 (N_13006,N_7151,N_6566);
nor U13007 (N_13007,N_8153,N_7318);
and U13008 (N_13008,N_9926,N_5334);
and U13009 (N_13009,N_8085,N_8946);
or U13010 (N_13010,N_7011,N_5664);
nor U13011 (N_13011,N_7051,N_5165);
and U13012 (N_13012,N_8393,N_8278);
and U13013 (N_13013,N_9243,N_6413);
and U13014 (N_13014,N_6081,N_6593);
and U13015 (N_13015,N_8573,N_7474);
and U13016 (N_13016,N_6957,N_7536);
or U13017 (N_13017,N_5344,N_5321);
or U13018 (N_13018,N_5364,N_6061);
nand U13019 (N_13019,N_5567,N_8006);
or U13020 (N_13020,N_9891,N_5856);
xnor U13021 (N_13021,N_9660,N_6336);
nor U13022 (N_13022,N_5257,N_7294);
and U13023 (N_13023,N_9143,N_7416);
nand U13024 (N_13024,N_6613,N_9305);
nor U13025 (N_13025,N_8276,N_5504);
nand U13026 (N_13026,N_6980,N_6880);
or U13027 (N_13027,N_7921,N_8980);
and U13028 (N_13028,N_8886,N_5867);
or U13029 (N_13029,N_7610,N_7608);
or U13030 (N_13030,N_5192,N_9384);
nand U13031 (N_13031,N_8954,N_8515);
and U13032 (N_13032,N_8198,N_6712);
or U13033 (N_13033,N_8883,N_9037);
or U13034 (N_13034,N_6009,N_6264);
and U13035 (N_13035,N_5780,N_5705);
and U13036 (N_13036,N_9642,N_6273);
nor U13037 (N_13037,N_9233,N_6493);
nor U13038 (N_13038,N_6586,N_5400);
nor U13039 (N_13039,N_6449,N_9150);
or U13040 (N_13040,N_7998,N_6132);
nand U13041 (N_13041,N_9732,N_6999);
or U13042 (N_13042,N_5930,N_8120);
and U13043 (N_13043,N_9327,N_9969);
or U13044 (N_13044,N_6254,N_8180);
and U13045 (N_13045,N_9946,N_9399);
xor U13046 (N_13046,N_5398,N_6921);
nor U13047 (N_13047,N_9518,N_5349);
or U13048 (N_13048,N_8740,N_7594);
nand U13049 (N_13049,N_5453,N_7831);
or U13050 (N_13050,N_8258,N_7430);
or U13051 (N_13051,N_9998,N_6053);
or U13052 (N_13052,N_6693,N_8913);
nand U13053 (N_13053,N_7880,N_9308);
or U13054 (N_13054,N_6093,N_7198);
nor U13055 (N_13055,N_7119,N_5718);
nor U13056 (N_13056,N_6983,N_8086);
and U13057 (N_13057,N_9333,N_8727);
nand U13058 (N_13058,N_9912,N_6394);
and U13059 (N_13059,N_7404,N_8110);
or U13060 (N_13060,N_9191,N_6542);
nor U13061 (N_13061,N_5553,N_9687);
nor U13062 (N_13062,N_9416,N_6477);
and U13063 (N_13063,N_8648,N_8127);
nor U13064 (N_13064,N_8693,N_8193);
and U13065 (N_13065,N_6638,N_6433);
nand U13066 (N_13066,N_7893,N_7547);
and U13067 (N_13067,N_5579,N_5473);
or U13068 (N_13068,N_5058,N_8649);
and U13069 (N_13069,N_7912,N_9815);
nand U13070 (N_13070,N_6932,N_7035);
or U13071 (N_13071,N_8945,N_8273);
and U13072 (N_13072,N_8484,N_9943);
nor U13073 (N_13073,N_5447,N_5933);
or U13074 (N_13074,N_6314,N_5264);
nor U13075 (N_13075,N_6986,N_9203);
or U13076 (N_13076,N_5698,N_9334);
nand U13077 (N_13077,N_5944,N_8714);
and U13078 (N_13078,N_5049,N_7387);
and U13079 (N_13079,N_7659,N_7627);
nand U13080 (N_13080,N_7753,N_6410);
and U13081 (N_13081,N_8534,N_7281);
xor U13082 (N_13082,N_9641,N_5755);
nor U13083 (N_13083,N_8496,N_7974);
and U13084 (N_13084,N_5759,N_7622);
or U13085 (N_13085,N_7524,N_6946);
and U13086 (N_13086,N_7896,N_5898);
or U13087 (N_13087,N_7833,N_6897);
nor U13088 (N_13088,N_8565,N_6092);
and U13089 (N_13089,N_6129,N_7147);
nand U13090 (N_13090,N_9097,N_7316);
nor U13091 (N_13091,N_8792,N_8242);
or U13092 (N_13092,N_5533,N_9304);
or U13093 (N_13093,N_5218,N_5163);
or U13094 (N_13094,N_9670,N_9829);
and U13095 (N_13095,N_8714,N_9199);
nor U13096 (N_13096,N_7887,N_8904);
nand U13097 (N_13097,N_9710,N_6520);
and U13098 (N_13098,N_8955,N_6521);
and U13099 (N_13099,N_7624,N_6142);
or U13100 (N_13100,N_8845,N_8699);
and U13101 (N_13101,N_6735,N_7476);
nor U13102 (N_13102,N_6272,N_7284);
and U13103 (N_13103,N_7531,N_8643);
nor U13104 (N_13104,N_7728,N_9842);
or U13105 (N_13105,N_6729,N_5484);
and U13106 (N_13106,N_9725,N_8881);
or U13107 (N_13107,N_7205,N_9073);
and U13108 (N_13108,N_5717,N_6599);
and U13109 (N_13109,N_5638,N_5369);
nand U13110 (N_13110,N_8598,N_6389);
nor U13111 (N_13111,N_7908,N_8655);
or U13112 (N_13112,N_8954,N_6901);
nand U13113 (N_13113,N_5580,N_8282);
and U13114 (N_13114,N_7446,N_5983);
and U13115 (N_13115,N_9626,N_7041);
or U13116 (N_13116,N_8618,N_8363);
and U13117 (N_13117,N_6311,N_8717);
nor U13118 (N_13118,N_8126,N_8141);
or U13119 (N_13119,N_9992,N_8090);
nor U13120 (N_13120,N_5599,N_7470);
or U13121 (N_13121,N_8512,N_7668);
nor U13122 (N_13122,N_9161,N_7744);
or U13123 (N_13123,N_6313,N_8805);
and U13124 (N_13124,N_7425,N_7731);
or U13125 (N_13125,N_9606,N_6920);
and U13126 (N_13126,N_7530,N_9001);
or U13127 (N_13127,N_7685,N_5799);
or U13128 (N_13128,N_7417,N_6856);
nor U13129 (N_13129,N_5358,N_6419);
and U13130 (N_13130,N_5337,N_8671);
or U13131 (N_13131,N_6049,N_5076);
and U13132 (N_13132,N_6494,N_7588);
nor U13133 (N_13133,N_5836,N_6712);
nor U13134 (N_13134,N_5712,N_9448);
nor U13135 (N_13135,N_9059,N_5019);
or U13136 (N_13136,N_6671,N_9235);
or U13137 (N_13137,N_5678,N_6754);
or U13138 (N_13138,N_7120,N_9767);
nand U13139 (N_13139,N_8746,N_9476);
or U13140 (N_13140,N_9630,N_8729);
or U13141 (N_13141,N_8554,N_5714);
nand U13142 (N_13142,N_9111,N_8753);
nor U13143 (N_13143,N_7385,N_6403);
and U13144 (N_13144,N_5195,N_8666);
or U13145 (N_13145,N_8400,N_6272);
and U13146 (N_13146,N_5934,N_9153);
or U13147 (N_13147,N_7877,N_8950);
nand U13148 (N_13148,N_7855,N_9655);
or U13149 (N_13149,N_8305,N_7391);
and U13150 (N_13150,N_6026,N_7104);
or U13151 (N_13151,N_8436,N_5805);
and U13152 (N_13152,N_5153,N_7159);
and U13153 (N_13153,N_9611,N_8818);
nor U13154 (N_13154,N_8146,N_6616);
or U13155 (N_13155,N_7492,N_5234);
nor U13156 (N_13156,N_8901,N_8935);
or U13157 (N_13157,N_7147,N_5523);
or U13158 (N_13158,N_6983,N_9135);
and U13159 (N_13159,N_7443,N_6375);
and U13160 (N_13160,N_5326,N_5515);
nand U13161 (N_13161,N_6843,N_5862);
nand U13162 (N_13162,N_8035,N_5173);
and U13163 (N_13163,N_7157,N_6297);
xor U13164 (N_13164,N_5242,N_5099);
nor U13165 (N_13165,N_7600,N_8663);
nor U13166 (N_13166,N_5561,N_6405);
and U13167 (N_13167,N_7002,N_6849);
or U13168 (N_13168,N_6442,N_5119);
or U13169 (N_13169,N_9588,N_5456);
nand U13170 (N_13170,N_5082,N_5925);
nor U13171 (N_13171,N_5296,N_8453);
nand U13172 (N_13172,N_6858,N_8997);
nand U13173 (N_13173,N_8798,N_9312);
nor U13174 (N_13174,N_8281,N_8216);
nor U13175 (N_13175,N_8438,N_9729);
or U13176 (N_13176,N_8343,N_5091);
nand U13177 (N_13177,N_6266,N_8409);
or U13178 (N_13178,N_8531,N_6756);
or U13179 (N_13179,N_6879,N_7173);
or U13180 (N_13180,N_6783,N_7237);
and U13181 (N_13181,N_6098,N_7712);
or U13182 (N_13182,N_7787,N_8366);
nand U13183 (N_13183,N_8408,N_8320);
nand U13184 (N_13184,N_9084,N_6022);
nand U13185 (N_13185,N_9324,N_8035);
or U13186 (N_13186,N_5138,N_6414);
or U13187 (N_13187,N_8149,N_5590);
nor U13188 (N_13188,N_6428,N_7642);
nand U13189 (N_13189,N_7165,N_9250);
or U13190 (N_13190,N_6978,N_5755);
and U13191 (N_13191,N_9740,N_5879);
nor U13192 (N_13192,N_5917,N_8196);
and U13193 (N_13193,N_8107,N_6603);
nand U13194 (N_13194,N_9091,N_8382);
nand U13195 (N_13195,N_5843,N_8799);
and U13196 (N_13196,N_8463,N_8151);
or U13197 (N_13197,N_8536,N_5635);
and U13198 (N_13198,N_7773,N_7702);
and U13199 (N_13199,N_7022,N_8663);
nor U13200 (N_13200,N_5419,N_6859);
nand U13201 (N_13201,N_5833,N_5682);
or U13202 (N_13202,N_8243,N_9872);
or U13203 (N_13203,N_7451,N_8753);
nand U13204 (N_13204,N_8497,N_5126);
and U13205 (N_13205,N_7496,N_5047);
nor U13206 (N_13206,N_6451,N_5918);
nor U13207 (N_13207,N_5036,N_9140);
nand U13208 (N_13208,N_8316,N_7436);
or U13209 (N_13209,N_8446,N_6468);
and U13210 (N_13210,N_7845,N_9239);
or U13211 (N_13211,N_5207,N_7087);
or U13212 (N_13212,N_7257,N_8300);
nor U13213 (N_13213,N_5304,N_5285);
and U13214 (N_13214,N_8603,N_5391);
nand U13215 (N_13215,N_9674,N_5274);
and U13216 (N_13216,N_7476,N_6660);
and U13217 (N_13217,N_9654,N_9500);
and U13218 (N_13218,N_5034,N_6488);
nand U13219 (N_13219,N_6328,N_9435);
or U13220 (N_13220,N_5670,N_8837);
or U13221 (N_13221,N_7095,N_8343);
nand U13222 (N_13222,N_9751,N_8212);
nand U13223 (N_13223,N_9574,N_6838);
nor U13224 (N_13224,N_5230,N_5700);
nor U13225 (N_13225,N_9349,N_9843);
nor U13226 (N_13226,N_8908,N_7674);
and U13227 (N_13227,N_5174,N_6932);
nor U13228 (N_13228,N_7991,N_7056);
or U13229 (N_13229,N_8240,N_8938);
and U13230 (N_13230,N_7448,N_5130);
and U13231 (N_13231,N_6304,N_7726);
nor U13232 (N_13232,N_6942,N_7452);
nor U13233 (N_13233,N_5588,N_8936);
nor U13234 (N_13234,N_9167,N_7037);
and U13235 (N_13235,N_6150,N_8582);
nor U13236 (N_13236,N_9302,N_6086);
or U13237 (N_13237,N_6418,N_7085);
nor U13238 (N_13238,N_8365,N_7414);
nor U13239 (N_13239,N_7719,N_7096);
and U13240 (N_13240,N_9403,N_5307);
nand U13241 (N_13241,N_6365,N_5622);
nand U13242 (N_13242,N_6871,N_8717);
nor U13243 (N_13243,N_6719,N_8289);
xor U13244 (N_13244,N_8370,N_6134);
xor U13245 (N_13245,N_9568,N_7026);
nand U13246 (N_13246,N_8407,N_7815);
nand U13247 (N_13247,N_9259,N_7186);
nand U13248 (N_13248,N_5257,N_7388);
or U13249 (N_13249,N_9785,N_9161);
or U13250 (N_13250,N_9013,N_5249);
nand U13251 (N_13251,N_7344,N_6416);
nor U13252 (N_13252,N_5074,N_5313);
and U13253 (N_13253,N_8775,N_8026);
nor U13254 (N_13254,N_9738,N_7229);
xor U13255 (N_13255,N_7781,N_6728);
nor U13256 (N_13256,N_6440,N_5653);
nand U13257 (N_13257,N_8203,N_7793);
nor U13258 (N_13258,N_6900,N_5058);
nor U13259 (N_13259,N_5770,N_8839);
or U13260 (N_13260,N_8967,N_7863);
nand U13261 (N_13261,N_6876,N_8494);
nand U13262 (N_13262,N_9321,N_8277);
nand U13263 (N_13263,N_6349,N_8894);
nand U13264 (N_13264,N_5044,N_8360);
and U13265 (N_13265,N_6130,N_9613);
and U13266 (N_13266,N_9404,N_7823);
or U13267 (N_13267,N_9525,N_5412);
nand U13268 (N_13268,N_9061,N_5903);
or U13269 (N_13269,N_8396,N_5921);
nor U13270 (N_13270,N_8518,N_8796);
and U13271 (N_13271,N_6114,N_5865);
nor U13272 (N_13272,N_7371,N_9616);
and U13273 (N_13273,N_6719,N_6244);
nand U13274 (N_13274,N_8028,N_6196);
and U13275 (N_13275,N_8480,N_5519);
or U13276 (N_13276,N_9245,N_9578);
and U13277 (N_13277,N_8650,N_8078);
and U13278 (N_13278,N_6487,N_5474);
xor U13279 (N_13279,N_6568,N_9891);
nand U13280 (N_13280,N_8396,N_7139);
or U13281 (N_13281,N_5016,N_9970);
or U13282 (N_13282,N_6560,N_7906);
nor U13283 (N_13283,N_6552,N_9003);
and U13284 (N_13284,N_5206,N_8088);
nand U13285 (N_13285,N_8965,N_5573);
nand U13286 (N_13286,N_9198,N_9683);
or U13287 (N_13287,N_7423,N_7430);
and U13288 (N_13288,N_8570,N_7411);
and U13289 (N_13289,N_9162,N_5043);
nor U13290 (N_13290,N_8322,N_5102);
or U13291 (N_13291,N_8385,N_6917);
and U13292 (N_13292,N_5440,N_5127);
nand U13293 (N_13293,N_5010,N_8733);
nor U13294 (N_13294,N_8829,N_6977);
and U13295 (N_13295,N_8305,N_6503);
or U13296 (N_13296,N_6845,N_7544);
and U13297 (N_13297,N_9901,N_8761);
or U13298 (N_13298,N_9816,N_5018);
or U13299 (N_13299,N_8165,N_7069);
nand U13300 (N_13300,N_6183,N_8592);
nor U13301 (N_13301,N_9836,N_6584);
nand U13302 (N_13302,N_7998,N_5372);
nand U13303 (N_13303,N_9227,N_5046);
and U13304 (N_13304,N_8563,N_5125);
and U13305 (N_13305,N_7941,N_9873);
nand U13306 (N_13306,N_7573,N_6843);
and U13307 (N_13307,N_7102,N_5820);
nand U13308 (N_13308,N_7102,N_6713);
and U13309 (N_13309,N_7480,N_9058);
nand U13310 (N_13310,N_8544,N_9292);
nor U13311 (N_13311,N_9225,N_9434);
or U13312 (N_13312,N_9163,N_7962);
nand U13313 (N_13313,N_7448,N_9652);
and U13314 (N_13314,N_7663,N_9115);
or U13315 (N_13315,N_6833,N_8796);
or U13316 (N_13316,N_7745,N_8520);
nand U13317 (N_13317,N_6403,N_6810);
nand U13318 (N_13318,N_6056,N_6947);
or U13319 (N_13319,N_7385,N_6362);
or U13320 (N_13320,N_8616,N_9355);
and U13321 (N_13321,N_9041,N_9960);
and U13322 (N_13322,N_7712,N_8496);
and U13323 (N_13323,N_9265,N_7685);
nor U13324 (N_13324,N_8670,N_8250);
or U13325 (N_13325,N_5730,N_6700);
nor U13326 (N_13326,N_8315,N_6027);
nor U13327 (N_13327,N_6682,N_7016);
or U13328 (N_13328,N_9066,N_9859);
nor U13329 (N_13329,N_8905,N_6765);
nor U13330 (N_13330,N_6124,N_6426);
xor U13331 (N_13331,N_7001,N_7993);
and U13332 (N_13332,N_9777,N_8992);
or U13333 (N_13333,N_7080,N_9393);
nor U13334 (N_13334,N_5554,N_5885);
and U13335 (N_13335,N_5003,N_9181);
nor U13336 (N_13336,N_6380,N_5496);
or U13337 (N_13337,N_9313,N_6270);
nor U13338 (N_13338,N_6691,N_6897);
nor U13339 (N_13339,N_8092,N_5706);
or U13340 (N_13340,N_6631,N_5872);
nor U13341 (N_13341,N_9276,N_6384);
or U13342 (N_13342,N_8592,N_9419);
and U13343 (N_13343,N_9269,N_8078);
and U13344 (N_13344,N_8264,N_9748);
nor U13345 (N_13345,N_5407,N_6227);
or U13346 (N_13346,N_8602,N_6323);
xnor U13347 (N_13347,N_9800,N_7178);
nor U13348 (N_13348,N_5096,N_6838);
and U13349 (N_13349,N_7443,N_7604);
and U13350 (N_13350,N_8052,N_5680);
nand U13351 (N_13351,N_8107,N_7828);
nand U13352 (N_13352,N_7648,N_6987);
or U13353 (N_13353,N_6358,N_9136);
and U13354 (N_13354,N_8304,N_6683);
and U13355 (N_13355,N_8551,N_6965);
and U13356 (N_13356,N_5575,N_5178);
and U13357 (N_13357,N_9516,N_7448);
nand U13358 (N_13358,N_6719,N_7923);
nand U13359 (N_13359,N_7224,N_6020);
or U13360 (N_13360,N_9507,N_7020);
or U13361 (N_13361,N_7202,N_6123);
or U13362 (N_13362,N_8826,N_9147);
nand U13363 (N_13363,N_9394,N_5881);
nand U13364 (N_13364,N_7236,N_9503);
nand U13365 (N_13365,N_5340,N_7240);
or U13366 (N_13366,N_5392,N_6497);
or U13367 (N_13367,N_5187,N_5008);
nand U13368 (N_13368,N_7185,N_6695);
and U13369 (N_13369,N_8849,N_5886);
nor U13370 (N_13370,N_6003,N_6426);
nor U13371 (N_13371,N_7624,N_5851);
or U13372 (N_13372,N_8171,N_5744);
or U13373 (N_13373,N_9762,N_7136);
or U13374 (N_13374,N_7555,N_5988);
or U13375 (N_13375,N_9864,N_6922);
nor U13376 (N_13376,N_5144,N_7519);
nor U13377 (N_13377,N_7951,N_6349);
or U13378 (N_13378,N_5144,N_5162);
and U13379 (N_13379,N_7407,N_8342);
and U13380 (N_13380,N_9650,N_5546);
or U13381 (N_13381,N_7966,N_8504);
nor U13382 (N_13382,N_8786,N_9867);
nand U13383 (N_13383,N_9481,N_6650);
nor U13384 (N_13384,N_8238,N_9007);
and U13385 (N_13385,N_5803,N_7649);
nand U13386 (N_13386,N_8658,N_7603);
and U13387 (N_13387,N_5394,N_9283);
or U13388 (N_13388,N_5653,N_6949);
xor U13389 (N_13389,N_5247,N_6495);
nand U13390 (N_13390,N_8914,N_6748);
nand U13391 (N_13391,N_7826,N_8595);
nand U13392 (N_13392,N_7867,N_9295);
nor U13393 (N_13393,N_7685,N_5219);
nand U13394 (N_13394,N_9513,N_8665);
or U13395 (N_13395,N_7898,N_8396);
and U13396 (N_13396,N_5136,N_5026);
or U13397 (N_13397,N_5195,N_8612);
or U13398 (N_13398,N_9908,N_5202);
nand U13399 (N_13399,N_8451,N_8602);
and U13400 (N_13400,N_7454,N_9645);
nand U13401 (N_13401,N_8931,N_8221);
and U13402 (N_13402,N_7953,N_8489);
nand U13403 (N_13403,N_6969,N_9411);
and U13404 (N_13404,N_6283,N_7233);
nand U13405 (N_13405,N_7388,N_5748);
or U13406 (N_13406,N_5501,N_5684);
or U13407 (N_13407,N_8399,N_7079);
and U13408 (N_13408,N_6475,N_9030);
and U13409 (N_13409,N_6287,N_5785);
nor U13410 (N_13410,N_7117,N_9446);
or U13411 (N_13411,N_9288,N_9411);
nand U13412 (N_13412,N_7019,N_8016);
nand U13413 (N_13413,N_9263,N_6901);
and U13414 (N_13414,N_9572,N_6604);
nand U13415 (N_13415,N_6201,N_6159);
nor U13416 (N_13416,N_9421,N_8631);
xor U13417 (N_13417,N_6208,N_7086);
or U13418 (N_13418,N_8516,N_6816);
or U13419 (N_13419,N_9173,N_9146);
nand U13420 (N_13420,N_7010,N_5816);
nor U13421 (N_13421,N_9368,N_5920);
and U13422 (N_13422,N_7103,N_5365);
and U13423 (N_13423,N_8924,N_6923);
nor U13424 (N_13424,N_9960,N_8527);
and U13425 (N_13425,N_7855,N_6605);
nor U13426 (N_13426,N_6990,N_7161);
nor U13427 (N_13427,N_9995,N_7115);
nand U13428 (N_13428,N_9520,N_8990);
or U13429 (N_13429,N_6885,N_7539);
and U13430 (N_13430,N_8009,N_7791);
or U13431 (N_13431,N_8110,N_8621);
or U13432 (N_13432,N_6638,N_5983);
nand U13433 (N_13433,N_9076,N_6214);
nand U13434 (N_13434,N_9221,N_6377);
or U13435 (N_13435,N_5046,N_7442);
or U13436 (N_13436,N_8137,N_9914);
and U13437 (N_13437,N_5774,N_5273);
or U13438 (N_13438,N_5011,N_6766);
or U13439 (N_13439,N_5835,N_8059);
nor U13440 (N_13440,N_6019,N_8939);
or U13441 (N_13441,N_8342,N_5117);
xnor U13442 (N_13442,N_5629,N_6341);
or U13443 (N_13443,N_9840,N_6850);
nor U13444 (N_13444,N_7579,N_9460);
and U13445 (N_13445,N_5263,N_8861);
and U13446 (N_13446,N_9862,N_8256);
or U13447 (N_13447,N_7911,N_9355);
nand U13448 (N_13448,N_6944,N_6704);
and U13449 (N_13449,N_8137,N_9683);
or U13450 (N_13450,N_8392,N_7323);
nor U13451 (N_13451,N_5765,N_8902);
nor U13452 (N_13452,N_7008,N_6328);
nor U13453 (N_13453,N_8607,N_8525);
and U13454 (N_13454,N_6150,N_5325);
nor U13455 (N_13455,N_8173,N_5505);
or U13456 (N_13456,N_5129,N_6088);
nand U13457 (N_13457,N_9320,N_5916);
and U13458 (N_13458,N_9112,N_6441);
nand U13459 (N_13459,N_7274,N_6369);
and U13460 (N_13460,N_7452,N_7613);
nor U13461 (N_13461,N_6970,N_6342);
nor U13462 (N_13462,N_7221,N_7026);
and U13463 (N_13463,N_6252,N_8570);
and U13464 (N_13464,N_8992,N_9602);
nand U13465 (N_13465,N_6061,N_8257);
nor U13466 (N_13466,N_5582,N_9561);
and U13467 (N_13467,N_7893,N_9493);
or U13468 (N_13468,N_5387,N_6351);
nor U13469 (N_13469,N_6071,N_9386);
and U13470 (N_13470,N_7200,N_6888);
and U13471 (N_13471,N_7043,N_6606);
nand U13472 (N_13472,N_7716,N_9566);
and U13473 (N_13473,N_8840,N_6174);
nand U13474 (N_13474,N_9799,N_8699);
or U13475 (N_13475,N_7354,N_6828);
or U13476 (N_13476,N_7987,N_8525);
nand U13477 (N_13477,N_7330,N_9742);
and U13478 (N_13478,N_9395,N_6793);
nand U13479 (N_13479,N_6834,N_7707);
nand U13480 (N_13480,N_6489,N_8058);
nor U13481 (N_13481,N_5278,N_6843);
and U13482 (N_13482,N_7210,N_5222);
nor U13483 (N_13483,N_5365,N_6408);
nand U13484 (N_13484,N_6873,N_9581);
nand U13485 (N_13485,N_5456,N_7006);
nor U13486 (N_13486,N_6353,N_7883);
and U13487 (N_13487,N_5998,N_8813);
and U13488 (N_13488,N_6076,N_8722);
and U13489 (N_13489,N_9365,N_9055);
or U13490 (N_13490,N_6637,N_7419);
nand U13491 (N_13491,N_5817,N_8414);
nand U13492 (N_13492,N_5170,N_5923);
and U13493 (N_13493,N_7174,N_5215);
nand U13494 (N_13494,N_9208,N_7596);
nand U13495 (N_13495,N_7519,N_5048);
nand U13496 (N_13496,N_8104,N_8893);
nor U13497 (N_13497,N_5347,N_6928);
nor U13498 (N_13498,N_8149,N_7735);
nor U13499 (N_13499,N_6459,N_7483);
and U13500 (N_13500,N_9155,N_7255);
xnor U13501 (N_13501,N_9340,N_7868);
and U13502 (N_13502,N_5041,N_7600);
and U13503 (N_13503,N_7946,N_6940);
and U13504 (N_13504,N_8353,N_6029);
or U13505 (N_13505,N_8486,N_7788);
nand U13506 (N_13506,N_5045,N_6755);
nand U13507 (N_13507,N_8254,N_5624);
nor U13508 (N_13508,N_5958,N_7920);
nand U13509 (N_13509,N_8173,N_5448);
or U13510 (N_13510,N_9121,N_7468);
and U13511 (N_13511,N_5462,N_5817);
nand U13512 (N_13512,N_6428,N_5073);
nor U13513 (N_13513,N_5072,N_9019);
nand U13514 (N_13514,N_7391,N_8087);
nand U13515 (N_13515,N_5995,N_6325);
and U13516 (N_13516,N_5538,N_8458);
and U13517 (N_13517,N_8540,N_8490);
or U13518 (N_13518,N_9796,N_8105);
nor U13519 (N_13519,N_5915,N_9202);
and U13520 (N_13520,N_9704,N_8320);
nand U13521 (N_13521,N_8918,N_7201);
nor U13522 (N_13522,N_5033,N_6707);
or U13523 (N_13523,N_7747,N_9988);
nor U13524 (N_13524,N_9006,N_5557);
nor U13525 (N_13525,N_9322,N_9058);
xor U13526 (N_13526,N_6829,N_6277);
and U13527 (N_13527,N_9797,N_9096);
and U13528 (N_13528,N_5225,N_6891);
nor U13529 (N_13529,N_6880,N_9061);
and U13530 (N_13530,N_9824,N_5617);
nor U13531 (N_13531,N_5910,N_9149);
nor U13532 (N_13532,N_8545,N_5403);
or U13533 (N_13533,N_7406,N_8001);
nor U13534 (N_13534,N_9282,N_6012);
nand U13535 (N_13535,N_5626,N_5354);
nand U13536 (N_13536,N_8107,N_5955);
and U13537 (N_13537,N_9084,N_7165);
nand U13538 (N_13538,N_7842,N_9815);
nand U13539 (N_13539,N_6236,N_7297);
and U13540 (N_13540,N_6731,N_6854);
nand U13541 (N_13541,N_9001,N_9732);
or U13542 (N_13542,N_5319,N_8411);
or U13543 (N_13543,N_7034,N_5315);
or U13544 (N_13544,N_8575,N_6770);
or U13545 (N_13545,N_9492,N_8053);
and U13546 (N_13546,N_7760,N_5345);
nor U13547 (N_13547,N_5251,N_6986);
and U13548 (N_13548,N_9309,N_9653);
nor U13549 (N_13549,N_8819,N_6705);
or U13550 (N_13550,N_5199,N_5102);
nor U13551 (N_13551,N_5491,N_6831);
and U13552 (N_13552,N_6068,N_5225);
or U13553 (N_13553,N_7970,N_8564);
nand U13554 (N_13554,N_6179,N_6781);
or U13555 (N_13555,N_6385,N_7099);
nand U13556 (N_13556,N_8668,N_7076);
or U13557 (N_13557,N_6243,N_8735);
and U13558 (N_13558,N_9511,N_5499);
xnor U13559 (N_13559,N_8747,N_5120);
nand U13560 (N_13560,N_5500,N_8003);
nand U13561 (N_13561,N_5126,N_9348);
and U13562 (N_13562,N_9972,N_8922);
nor U13563 (N_13563,N_7786,N_8233);
nand U13564 (N_13564,N_7008,N_8719);
and U13565 (N_13565,N_5489,N_5872);
nand U13566 (N_13566,N_9783,N_9724);
xnor U13567 (N_13567,N_5272,N_9419);
and U13568 (N_13568,N_7382,N_5122);
and U13569 (N_13569,N_7821,N_8975);
nor U13570 (N_13570,N_6719,N_6092);
nor U13571 (N_13571,N_5236,N_8684);
nand U13572 (N_13572,N_8727,N_6649);
or U13573 (N_13573,N_9665,N_5091);
nor U13574 (N_13574,N_9779,N_8245);
nor U13575 (N_13575,N_8792,N_9413);
or U13576 (N_13576,N_7693,N_5278);
or U13577 (N_13577,N_5737,N_9102);
nor U13578 (N_13578,N_6387,N_6355);
nand U13579 (N_13579,N_6628,N_7357);
nor U13580 (N_13580,N_8653,N_7531);
nand U13581 (N_13581,N_8956,N_9332);
or U13582 (N_13582,N_5877,N_8731);
or U13583 (N_13583,N_8587,N_6553);
or U13584 (N_13584,N_9102,N_9455);
and U13585 (N_13585,N_9052,N_9562);
and U13586 (N_13586,N_5225,N_7066);
nand U13587 (N_13587,N_8532,N_9835);
nand U13588 (N_13588,N_7195,N_7181);
xnor U13589 (N_13589,N_8935,N_7160);
nor U13590 (N_13590,N_8396,N_7875);
nor U13591 (N_13591,N_5465,N_5130);
and U13592 (N_13592,N_5601,N_6238);
nand U13593 (N_13593,N_6753,N_9123);
nand U13594 (N_13594,N_8111,N_6314);
nor U13595 (N_13595,N_9668,N_9546);
nand U13596 (N_13596,N_7592,N_6162);
nand U13597 (N_13597,N_5699,N_6184);
nand U13598 (N_13598,N_7482,N_6714);
or U13599 (N_13599,N_5344,N_7916);
nand U13600 (N_13600,N_5096,N_7002);
xnor U13601 (N_13601,N_7034,N_5876);
and U13602 (N_13602,N_6109,N_5473);
nor U13603 (N_13603,N_5447,N_7752);
nand U13604 (N_13604,N_8396,N_6474);
and U13605 (N_13605,N_6195,N_6361);
or U13606 (N_13606,N_8624,N_9288);
nor U13607 (N_13607,N_5756,N_7931);
nor U13608 (N_13608,N_6826,N_7867);
nor U13609 (N_13609,N_5282,N_8578);
or U13610 (N_13610,N_8025,N_7082);
nand U13611 (N_13611,N_6493,N_7076);
or U13612 (N_13612,N_5131,N_9920);
nor U13613 (N_13613,N_6811,N_9003);
and U13614 (N_13614,N_7764,N_9857);
nor U13615 (N_13615,N_7067,N_5004);
nand U13616 (N_13616,N_5744,N_6052);
nand U13617 (N_13617,N_9596,N_9339);
nor U13618 (N_13618,N_9071,N_9579);
and U13619 (N_13619,N_5819,N_9739);
or U13620 (N_13620,N_6005,N_6776);
and U13621 (N_13621,N_6744,N_7212);
nor U13622 (N_13622,N_9924,N_7462);
nor U13623 (N_13623,N_7861,N_9635);
nor U13624 (N_13624,N_8153,N_9752);
nand U13625 (N_13625,N_6553,N_7083);
and U13626 (N_13626,N_6425,N_5920);
or U13627 (N_13627,N_9229,N_8774);
or U13628 (N_13628,N_7529,N_8342);
nand U13629 (N_13629,N_5175,N_9740);
and U13630 (N_13630,N_8907,N_7853);
nor U13631 (N_13631,N_5247,N_9901);
nand U13632 (N_13632,N_9316,N_5408);
and U13633 (N_13633,N_6597,N_6442);
nor U13634 (N_13634,N_5122,N_5979);
or U13635 (N_13635,N_9959,N_9686);
nand U13636 (N_13636,N_5745,N_8215);
nor U13637 (N_13637,N_7509,N_6090);
and U13638 (N_13638,N_5747,N_8685);
and U13639 (N_13639,N_9527,N_8586);
nor U13640 (N_13640,N_7173,N_5665);
nand U13641 (N_13641,N_7659,N_9449);
and U13642 (N_13642,N_8763,N_6354);
or U13643 (N_13643,N_5351,N_9376);
nor U13644 (N_13644,N_9179,N_6790);
and U13645 (N_13645,N_9277,N_8624);
and U13646 (N_13646,N_8726,N_9190);
nand U13647 (N_13647,N_8331,N_8484);
and U13648 (N_13648,N_8190,N_6052);
or U13649 (N_13649,N_9817,N_7544);
and U13650 (N_13650,N_9952,N_8170);
nor U13651 (N_13651,N_8455,N_5730);
and U13652 (N_13652,N_8644,N_6209);
nor U13653 (N_13653,N_8857,N_6178);
and U13654 (N_13654,N_5781,N_6766);
or U13655 (N_13655,N_8467,N_9359);
nand U13656 (N_13656,N_6498,N_8556);
nor U13657 (N_13657,N_9767,N_7103);
nand U13658 (N_13658,N_8578,N_8433);
nand U13659 (N_13659,N_5682,N_6008);
or U13660 (N_13660,N_7119,N_9248);
nor U13661 (N_13661,N_8655,N_5879);
or U13662 (N_13662,N_6210,N_9151);
nand U13663 (N_13663,N_5695,N_8132);
or U13664 (N_13664,N_5037,N_9610);
nand U13665 (N_13665,N_6342,N_6549);
nor U13666 (N_13666,N_6143,N_9495);
and U13667 (N_13667,N_8760,N_6135);
nor U13668 (N_13668,N_6260,N_5151);
nor U13669 (N_13669,N_9907,N_6999);
and U13670 (N_13670,N_7785,N_5940);
nor U13671 (N_13671,N_7820,N_6205);
nor U13672 (N_13672,N_7155,N_6406);
or U13673 (N_13673,N_8862,N_8718);
and U13674 (N_13674,N_7722,N_5676);
and U13675 (N_13675,N_5262,N_6096);
nor U13676 (N_13676,N_8421,N_7257);
or U13677 (N_13677,N_6148,N_7914);
nand U13678 (N_13678,N_6688,N_7798);
and U13679 (N_13679,N_5545,N_7148);
and U13680 (N_13680,N_5943,N_7740);
or U13681 (N_13681,N_6848,N_8347);
and U13682 (N_13682,N_5294,N_6441);
nor U13683 (N_13683,N_9933,N_7159);
xor U13684 (N_13684,N_8136,N_6536);
xor U13685 (N_13685,N_7736,N_5764);
or U13686 (N_13686,N_9051,N_8204);
or U13687 (N_13687,N_5806,N_6293);
and U13688 (N_13688,N_8434,N_5546);
and U13689 (N_13689,N_5489,N_6455);
nor U13690 (N_13690,N_9086,N_8096);
and U13691 (N_13691,N_5050,N_9294);
nand U13692 (N_13692,N_7652,N_9375);
and U13693 (N_13693,N_7102,N_7437);
xnor U13694 (N_13694,N_8787,N_7544);
nor U13695 (N_13695,N_7553,N_5310);
nand U13696 (N_13696,N_8478,N_8253);
or U13697 (N_13697,N_7531,N_7177);
nor U13698 (N_13698,N_6611,N_5076);
or U13699 (N_13699,N_9935,N_6163);
or U13700 (N_13700,N_9465,N_9168);
nand U13701 (N_13701,N_5004,N_8297);
nand U13702 (N_13702,N_6803,N_9522);
and U13703 (N_13703,N_5286,N_9782);
nand U13704 (N_13704,N_6574,N_9885);
nor U13705 (N_13705,N_8027,N_6214);
and U13706 (N_13706,N_5667,N_7054);
nand U13707 (N_13707,N_7711,N_8540);
or U13708 (N_13708,N_6759,N_6005);
nor U13709 (N_13709,N_9303,N_7303);
nand U13710 (N_13710,N_6768,N_6512);
nand U13711 (N_13711,N_6895,N_5418);
or U13712 (N_13712,N_7068,N_8784);
and U13713 (N_13713,N_9050,N_8526);
and U13714 (N_13714,N_6536,N_5794);
or U13715 (N_13715,N_9604,N_9138);
nand U13716 (N_13716,N_5729,N_7338);
nor U13717 (N_13717,N_9047,N_9704);
nor U13718 (N_13718,N_6170,N_7634);
nor U13719 (N_13719,N_8156,N_9106);
or U13720 (N_13720,N_5993,N_7963);
nor U13721 (N_13721,N_7617,N_8942);
or U13722 (N_13722,N_7512,N_6997);
or U13723 (N_13723,N_6033,N_5541);
and U13724 (N_13724,N_8113,N_6621);
or U13725 (N_13725,N_8928,N_8720);
or U13726 (N_13726,N_5831,N_9802);
nand U13727 (N_13727,N_6242,N_8978);
and U13728 (N_13728,N_9469,N_9619);
or U13729 (N_13729,N_9421,N_7444);
nand U13730 (N_13730,N_8898,N_7757);
and U13731 (N_13731,N_7078,N_6408);
nor U13732 (N_13732,N_8883,N_7602);
nand U13733 (N_13733,N_8258,N_9022);
nor U13734 (N_13734,N_8605,N_9707);
nand U13735 (N_13735,N_5901,N_9725);
nand U13736 (N_13736,N_6348,N_7499);
nand U13737 (N_13737,N_5989,N_8993);
nand U13738 (N_13738,N_6296,N_6100);
or U13739 (N_13739,N_8720,N_7628);
and U13740 (N_13740,N_5648,N_7192);
nand U13741 (N_13741,N_7549,N_5289);
and U13742 (N_13742,N_8175,N_9303);
nor U13743 (N_13743,N_9022,N_9303);
nand U13744 (N_13744,N_7443,N_9585);
nor U13745 (N_13745,N_7988,N_9579);
nor U13746 (N_13746,N_5435,N_7152);
and U13747 (N_13747,N_6416,N_8317);
or U13748 (N_13748,N_9930,N_8882);
nor U13749 (N_13749,N_8063,N_7026);
nand U13750 (N_13750,N_9514,N_7352);
nor U13751 (N_13751,N_9692,N_5821);
nor U13752 (N_13752,N_9853,N_6865);
nor U13753 (N_13753,N_9370,N_6562);
or U13754 (N_13754,N_8894,N_7525);
and U13755 (N_13755,N_6410,N_7894);
or U13756 (N_13756,N_8314,N_8691);
or U13757 (N_13757,N_5515,N_5544);
nor U13758 (N_13758,N_8299,N_8692);
nand U13759 (N_13759,N_7586,N_7241);
nor U13760 (N_13760,N_9441,N_5073);
and U13761 (N_13761,N_5661,N_7033);
nand U13762 (N_13762,N_7400,N_9506);
nor U13763 (N_13763,N_6274,N_7487);
or U13764 (N_13764,N_8830,N_7251);
or U13765 (N_13765,N_9113,N_6789);
or U13766 (N_13766,N_7365,N_9404);
nand U13767 (N_13767,N_9310,N_6836);
nand U13768 (N_13768,N_7931,N_5374);
nor U13769 (N_13769,N_6152,N_8545);
or U13770 (N_13770,N_6135,N_8297);
nor U13771 (N_13771,N_8462,N_5073);
nand U13772 (N_13772,N_6440,N_9335);
or U13773 (N_13773,N_8584,N_7576);
or U13774 (N_13774,N_7273,N_6793);
nor U13775 (N_13775,N_7588,N_5539);
xor U13776 (N_13776,N_5069,N_5487);
and U13777 (N_13777,N_7659,N_9763);
and U13778 (N_13778,N_8937,N_9549);
and U13779 (N_13779,N_8876,N_6121);
nand U13780 (N_13780,N_9563,N_9838);
nor U13781 (N_13781,N_6084,N_5384);
nor U13782 (N_13782,N_9093,N_7062);
nor U13783 (N_13783,N_7534,N_7716);
nor U13784 (N_13784,N_8301,N_8440);
and U13785 (N_13785,N_8482,N_5374);
or U13786 (N_13786,N_7918,N_8125);
nor U13787 (N_13787,N_7018,N_8669);
nor U13788 (N_13788,N_7962,N_7198);
nand U13789 (N_13789,N_6079,N_8792);
or U13790 (N_13790,N_9925,N_9610);
or U13791 (N_13791,N_5496,N_9286);
nand U13792 (N_13792,N_6474,N_9064);
and U13793 (N_13793,N_8995,N_5431);
or U13794 (N_13794,N_9894,N_7271);
nor U13795 (N_13795,N_8292,N_7162);
nor U13796 (N_13796,N_8927,N_8092);
or U13797 (N_13797,N_6187,N_8934);
or U13798 (N_13798,N_5626,N_8748);
and U13799 (N_13799,N_9840,N_8530);
or U13800 (N_13800,N_8326,N_6957);
nor U13801 (N_13801,N_9511,N_7317);
and U13802 (N_13802,N_9854,N_7654);
or U13803 (N_13803,N_9099,N_5493);
and U13804 (N_13804,N_6493,N_9720);
and U13805 (N_13805,N_5611,N_5762);
nand U13806 (N_13806,N_9400,N_6170);
nor U13807 (N_13807,N_8758,N_9441);
nor U13808 (N_13808,N_9601,N_9684);
nand U13809 (N_13809,N_8334,N_8130);
nand U13810 (N_13810,N_7250,N_8120);
xnor U13811 (N_13811,N_9306,N_5807);
or U13812 (N_13812,N_8541,N_9832);
nor U13813 (N_13813,N_5107,N_7194);
nor U13814 (N_13814,N_5249,N_8769);
nor U13815 (N_13815,N_7344,N_5659);
nand U13816 (N_13816,N_6617,N_5093);
and U13817 (N_13817,N_5303,N_6170);
and U13818 (N_13818,N_8837,N_6845);
and U13819 (N_13819,N_7583,N_5690);
and U13820 (N_13820,N_8372,N_8745);
nor U13821 (N_13821,N_9596,N_5015);
nor U13822 (N_13822,N_8789,N_7542);
nand U13823 (N_13823,N_8837,N_6775);
nand U13824 (N_13824,N_9715,N_8538);
or U13825 (N_13825,N_7730,N_6917);
nor U13826 (N_13826,N_6163,N_8008);
and U13827 (N_13827,N_6340,N_6556);
xnor U13828 (N_13828,N_9159,N_9021);
and U13829 (N_13829,N_6521,N_6277);
nand U13830 (N_13830,N_9482,N_8010);
nor U13831 (N_13831,N_9969,N_8899);
and U13832 (N_13832,N_7615,N_7695);
nand U13833 (N_13833,N_9573,N_5074);
nand U13834 (N_13834,N_8876,N_5529);
nor U13835 (N_13835,N_7458,N_5574);
or U13836 (N_13836,N_6673,N_7699);
nand U13837 (N_13837,N_7782,N_6886);
and U13838 (N_13838,N_5904,N_8848);
and U13839 (N_13839,N_8267,N_8093);
and U13840 (N_13840,N_8539,N_5047);
nor U13841 (N_13841,N_6561,N_9000);
and U13842 (N_13842,N_8837,N_7424);
and U13843 (N_13843,N_9319,N_5561);
nor U13844 (N_13844,N_7082,N_8683);
nor U13845 (N_13845,N_8924,N_7926);
and U13846 (N_13846,N_9830,N_5684);
and U13847 (N_13847,N_9514,N_6690);
nand U13848 (N_13848,N_9353,N_7778);
nand U13849 (N_13849,N_7140,N_6401);
and U13850 (N_13850,N_9031,N_8871);
and U13851 (N_13851,N_7284,N_5494);
or U13852 (N_13852,N_9732,N_9697);
or U13853 (N_13853,N_5652,N_8866);
or U13854 (N_13854,N_7911,N_5351);
nand U13855 (N_13855,N_6706,N_8375);
nor U13856 (N_13856,N_6025,N_5971);
or U13857 (N_13857,N_9632,N_9676);
nand U13858 (N_13858,N_8393,N_5007);
and U13859 (N_13859,N_5435,N_8567);
nand U13860 (N_13860,N_5217,N_5358);
or U13861 (N_13861,N_5501,N_9186);
nand U13862 (N_13862,N_8269,N_6669);
and U13863 (N_13863,N_7913,N_7520);
and U13864 (N_13864,N_5048,N_5894);
or U13865 (N_13865,N_9475,N_5801);
and U13866 (N_13866,N_8740,N_8953);
or U13867 (N_13867,N_7088,N_6307);
and U13868 (N_13868,N_7585,N_6632);
nand U13869 (N_13869,N_8567,N_6403);
nand U13870 (N_13870,N_7735,N_5330);
nor U13871 (N_13871,N_5286,N_9458);
nor U13872 (N_13872,N_9980,N_5167);
and U13873 (N_13873,N_8274,N_5966);
or U13874 (N_13874,N_6211,N_5511);
nand U13875 (N_13875,N_6254,N_6530);
and U13876 (N_13876,N_8797,N_9214);
or U13877 (N_13877,N_5048,N_9657);
or U13878 (N_13878,N_6430,N_8131);
nand U13879 (N_13879,N_9175,N_5198);
or U13880 (N_13880,N_8183,N_9228);
nand U13881 (N_13881,N_8239,N_8692);
or U13882 (N_13882,N_9913,N_5714);
and U13883 (N_13883,N_6603,N_8823);
or U13884 (N_13884,N_8882,N_6715);
and U13885 (N_13885,N_6587,N_9831);
nand U13886 (N_13886,N_7036,N_5671);
nor U13887 (N_13887,N_5419,N_8834);
or U13888 (N_13888,N_5898,N_8893);
nand U13889 (N_13889,N_8235,N_6099);
nand U13890 (N_13890,N_8934,N_6949);
xnor U13891 (N_13891,N_5515,N_6881);
nor U13892 (N_13892,N_7330,N_5882);
nand U13893 (N_13893,N_8067,N_6648);
nor U13894 (N_13894,N_7935,N_5651);
nand U13895 (N_13895,N_9782,N_5153);
nor U13896 (N_13896,N_9021,N_9313);
nand U13897 (N_13897,N_7788,N_5486);
or U13898 (N_13898,N_5412,N_8479);
nor U13899 (N_13899,N_5392,N_6029);
or U13900 (N_13900,N_7304,N_5860);
and U13901 (N_13901,N_8472,N_6909);
nor U13902 (N_13902,N_9203,N_6623);
and U13903 (N_13903,N_8314,N_9895);
and U13904 (N_13904,N_9739,N_7385);
or U13905 (N_13905,N_5175,N_5571);
nand U13906 (N_13906,N_9566,N_8567);
and U13907 (N_13907,N_6043,N_6759);
nor U13908 (N_13908,N_8098,N_7398);
and U13909 (N_13909,N_9954,N_9048);
nand U13910 (N_13910,N_8324,N_9824);
nand U13911 (N_13911,N_7264,N_8246);
nand U13912 (N_13912,N_8189,N_9902);
nor U13913 (N_13913,N_5139,N_8510);
and U13914 (N_13914,N_8792,N_7031);
nor U13915 (N_13915,N_9394,N_7642);
nor U13916 (N_13916,N_7033,N_7124);
nand U13917 (N_13917,N_7919,N_7293);
or U13918 (N_13918,N_5999,N_9982);
nor U13919 (N_13919,N_8608,N_8966);
nand U13920 (N_13920,N_7742,N_6469);
nand U13921 (N_13921,N_7589,N_9010);
nor U13922 (N_13922,N_9627,N_5240);
or U13923 (N_13923,N_8250,N_6816);
nor U13924 (N_13924,N_7486,N_8464);
nor U13925 (N_13925,N_5669,N_8660);
nor U13926 (N_13926,N_6487,N_7039);
nor U13927 (N_13927,N_6401,N_6030);
and U13928 (N_13928,N_7777,N_9687);
and U13929 (N_13929,N_8326,N_6494);
and U13930 (N_13930,N_7749,N_9832);
nand U13931 (N_13931,N_6980,N_8398);
nor U13932 (N_13932,N_5571,N_5598);
or U13933 (N_13933,N_7632,N_8437);
nor U13934 (N_13934,N_5003,N_9383);
nor U13935 (N_13935,N_6683,N_6501);
nor U13936 (N_13936,N_5166,N_6180);
nor U13937 (N_13937,N_8482,N_8209);
and U13938 (N_13938,N_6004,N_7011);
and U13939 (N_13939,N_5277,N_8510);
nand U13940 (N_13940,N_6999,N_8585);
nor U13941 (N_13941,N_9824,N_7877);
and U13942 (N_13942,N_9927,N_5200);
or U13943 (N_13943,N_8483,N_9035);
or U13944 (N_13944,N_9481,N_9624);
nand U13945 (N_13945,N_7069,N_6084);
nor U13946 (N_13946,N_8445,N_5664);
nand U13947 (N_13947,N_7145,N_6217);
nor U13948 (N_13948,N_5251,N_5821);
and U13949 (N_13949,N_5766,N_9747);
or U13950 (N_13950,N_5153,N_8348);
nor U13951 (N_13951,N_9344,N_6078);
nor U13952 (N_13952,N_6160,N_7365);
or U13953 (N_13953,N_5083,N_9568);
or U13954 (N_13954,N_5735,N_8247);
nand U13955 (N_13955,N_5406,N_7751);
nor U13956 (N_13956,N_7124,N_5455);
nor U13957 (N_13957,N_8655,N_6223);
or U13958 (N_13958,N_7820,N_5156);
nand U13959 (N_13959,N_9032,N_8901);
or U13960 (N_13960,N_6017,N_9135);
nor U13961 (N_13961,N_7615,N_5810);
nand U13962 (N_13962,N_7329,N_9156);
or U13963 (N_13963,N_6226,N_9800);
or U13964 (N_13964,N_5359,N_5001);
and U13965 (N_13965,N_7006,N_8127);
nor U13966 (N_13966,N_9858,N_5771);
nor U13967 (N_13967,N_5539,N_7671);
or U13968 (N_13968,N_9003,N_9045);
and U13969 (N_13969,N_5358,N_9125);
and U13970 (N_13970,N_9114,N_8547);
nand U13971 (N_13971,N_5440,N_7453);
nand U13972 (N_13972,N_5451,N_8206);
nand U13973 (N_13973,N_8692,N_8060);
nand U13974 (N_13974,N_5094,N_8186);
and U13975 (N_13975,N_6355,N_8102);
or U13976 (N_13976,N_8582,N_7977);
and U13977 (N_13977,N_8645,N_8091);
and U13978 (N_13978,N_9596,N_5107);
nor U13979 (N_13979,N_9620,N_9123);
or U13980 (N_13980,N_6335,N_6031);
nor U13981 (N_13981,N_8320,N_9115);
or U13982 (N_13982,N_7130,N_7012);
and U13983 (N_13983,N_8309,N_8014);
nand U13984 (N_13984,N_9926,N_7380);
and U13985 (N_13985,N_8065,N_9616);
nand U13986 (N_13986,N_9713,N_7913);
nand U13987 (N_13987,N_6638,N_5004);
nand U13988 (N_13988,N_8477,N_9632);
and U13989 (N_13989,N_7433,N_7804);
and U13990 (N_13990,N_5282,N_9976);
or U13991 (N_13991,N_8086,N_7680);
or U13992 (N_13992,N_7757,N_8831);
and U13993 (N_13993,N_8399,N_8414);
or U13994 (N_13994,N_6483,N_6963);
and U13995 (N_13995,N_8878,N_8595);
or U13996 (N_13996,N_9924,N_8983);
and U13997 (N_13997,N_8530,N_9899);
and U13998 (N_13998,N_8767,N_8332);
or U13999 (N_13999,N_5444,N_7942);
nor U14000 (N_14000,N_6563,N_6797);
and U14001 (N_14001,N_9744,N_7857);
nor U14002 (N_14002,N_6189,N_6108);
nand U14003 (N_14003,N_7791,N_6486);
nand U14004 (N_14004,N_9342,N_6435);
nand U14005 (N_14005,N_9974,N_5667);
and U14006 (N_14006,N_6486,N_8759);
and U14007 (N_14007,N_9717,N_6008);
nor U14008 (N_14008,N_9051,N_8497);
nor U14009 (N_14009,N_5422,N_6396);
or U14010 (N_14010,N_9652,N_5432);
and U14011 (N_14011,N_7807,N_7083);
and U14012 (N_14012,N_6544,N_6533);
or U14013 (N_14013,N_6129,N_7795);
nand U14014 (N_14014,N_8255,N_8235);
or U14015 (N_14015,N_7516,N_6418);
or U14016 (N_14016,N_6109,N_9276);
nand U14017 (N_14017,N_7440,N_9018);
and U14018 (N_14018,N_8872,N_7917);
nand U14019 (N_14019,N_5516,N_6037);
nor U14020 (N_14020,N_5516,N_8603);
and U14021 (N_14021,N_7346,N_9773);
nand U14022 (N_14022,N_5228,N_7243);
nand U14023 (N_14023,N_5508,N_8470);
and U14024 (N_14024,N_7805,N_7173);
and U14025 (N_14025,N_7100,N_8122);
or U14026 (N_14026,N_5442,N_9774);
and U14027 (N_14027,N_7051,N_9412);
nor U14028 (N_14028,N_7079,N_6609);
nand U14029 (N_14029,N_8556,N_5213);
nor U14030 (N_14030,N_9344,N_8065);
nor U14031 (N_14031,N_5753,N_5646);
nor U14032 (N_14032,N_5400,N_6330);
or U14033 (N_14033,N_5550,N_7437);
nand U14034 (N_14034,N_5142,N_5294);
nor U14035 (N_14035,N_8567,N_9074);
nand U14036 (N_14036,N_7474,N_7431);
or U14037 (N_14037,N_9667,N_8554);
and U14038 (N_14038,N_6755,N_9992);
nand U14039 (N_14039,N_7201,N_8585);
nor U14040 (N_14040,N_9702,N_8430);
nor U14041 (N_14041,N_8609,N_5258);
and U14042 (N_14042,N_9837,N_8474);
nand U14043 (N_14043,N_9149,N_7986);
nor U14044 (N_14044,N_6149,N_8246);
nor U14045 (N_14045,N_7218,N_7020);
or U14046 (N_14046,N_8229,N_9772);
and U14047 (N_14047,N_8650,N_5558);
nor U14048 (N_14048,N_5961,N_8908);
and U14049 (N_14049,N_9528,N_5734);
nor U14050 (N_14050,N_9073,N_9627);
and U14051 (N_14051,N_7460,N_6173);
or U14052 (N_14052,N_9855,N_6803);
and U14053 (N_14053,N_8124,N_6429);
nand U14054 (N_14054,N_9366,N_7527);
and U14055 (N_14055,N_8321,N_8932);
nand U14056 (N_14056,N_6909,N_8442);
nor U14057 (N_14057,N_6072,N_9610);
or U14058 (N_14058,N_7982,N_6001);
nand U14059 (N_14059,N_6753,N_9706);
nor U14060 (N_14060,N_8607,N_6742);
and U14061 (N_14061,N_5886,N_8399);
nor U14062 (N_14062,N_6806,N_6123);
or U14063 (N_14063,N_8870,N_9822);
nor U14064 (N_14064,N_9776,N_6214);
nand U14065 (N_14065,N_7122,N_6526);
nand U14066 (N_14066,N_9465,N_9756);
xor U14067 (N_14067,N_6922,N_5758);
nand U14068 (N_14068,N_8064,N_8219);
or U14069 (N_14069,N_7177,N_8649);
or U14070 (N_14070,N_5602,N_5215);
or U14071 (N_14071,N_6880,N_7056);
and U14072 (N_14072,N_7676,N_9257);
nand U14073 (N_14073,N_9464,N_9117);
or U14074 (N_14074,N_7260,N_8278);
nand U14075 (N_14075,N_7366,N_9288);
or U14076 (N_14076,N_6074,N_6819);
or U14077 (N_14077,N_9080,N_7400);
nor U14078 (N_14078,N_7668,N_7873);
or U14079 (N_14079,N_5773,N_9136);
nand U14080 (N_14080,N_9378,N_7319);
nand U14081 (N_14081,N_9075,N_5338);
or U14082 (N_14082,N_6055,N_5711);
nand U14083 (N_14083,N_8588,N_7047);
nor U14084 (N_14084,N_9271,N_6835);
or U14085 (N_14085,N_8290,N_9839);
nor U14086 (N_14086,N_5739,N_7596);
nand U14087 (N_14087,N_6963,N_6724);
or U14088 (N_14088,N_7450,N_9923);
nor U14089 (N_14089,N_9064,N_9435);
or U14090 (N_14090,N_7121,N_7912);
nor U14091 (N_14091,N_9690,N_7609);
nand U14092 (N_14092,N_9034,N_7935);
nand U14093 (N_14093,N_9538,N_6589);
and U14094 (N_14094,N_5765,N_7524);
or U14095 (N_14095,N_5395,N_5835);
or U14096 (N_14096,N_6169,N_9077);
nor U14097 (N_14097,N_9245,N_5738);
nor U14098 (N_14098,N_9298,N_5490);
and U14099 (N_14099,N_7328,N_9226);
nor U14100 (N_14100,N_6276,N_8232);
and U14101 (N_14101,N_9875,N_7585);
and U14102 (N_14102,N_8844,N_9416);
and U14103 (N_14103,N_7839,N_9345);
and U14104 (N_14104,N_5763,N_8970);
nand U14105 (N_14105,N_6785,N_6884);
or U14106 (N_14106,N_9091,N_9417);
and U14107 (N_14107,N_9095,N_8889);
and U14108 (N_14108,N_6983,N_9598);
and U14109 (N_14109,N_6180,N_9667);
nand U14110 (N_14110,N_5555,N_5814);
or U14111 (N_14111,N_9097,N_9249);
nor U14112 (N_14112,N_5718,N_5371);
nor U14113 (N_14113,N_5786,N_5314);
nor U14114 (N_14114,N_9474,N_9631);
nor U14115 (N_14115,N_9891,N_5918);
nor U14116 (N_14116,N_9710,N_7073);
or U14117 (N_14117,N_7381,N_6588);
nand U14118 (N_14118,N_9277,N_8453);
nand U14119 (N_14119,N_8584,N_5556);
nand U14120 (N_14120,N_8918,N_8278);
nor U14121 (N_14121,N_8366,N_9074);
nor U14122 (N_14122,N_5845,N_5873);
nor U14123 (N_14123,N_8528,N_8837);
or U14124 (N_14124,N_6888,N_5779);
and U14125 (N_14125,N_9550,N_6357);
or U14126 (N_14126,N_7988,N_6693);
nor U14127 (N_14127,N_9702,N_6410);
or U14128 (N_14128,N_8749,N_8200);
and U14129 (N_14129,N_6609,N_6268);
nor U14130 (N_14130,N_5759,N_5866);
nand U14131 (N_14131,N_9429,N_5965);
or U14132 (N_14132,N_7834,N_7485);
nor U14133 (N_14133,N_9587,N_8033);
or U14134 (N_14134,N_8945,N_6419);
nor U14135 (N_14135,N_9470,N_5069);
or U14136 (N_14136,N_6000,N_8435);
nor U14137 (N_14137,N_6020,N_9144);
and U14138 (N_14138,N_9706,N_9446);
or U14139 (N_14139,N_8757,N_5037);
nor U14140 (N_14140,N_7318,N_5200);
nor U14141 (N_14141,N_7470,N_9720);
and U14142 (N_14142,N_7854,N_8209);
xor U14143 (N_14143,N_8875,N_5329);
or U14144 (N_14144,N_5297,N_7077);
and U14145 (N_14145,N_9331,N_7781);
nor U14146 (N_14146,N_9579,N_8477);
nor U14147 (N_14147,N_6351,N_7974);
or U14148 (N_14148,N_5381,N_5504);
or U14149 (N_14149,N_7263,N_7280);
nor U14150 (N_14150,N_6063,N_6500);
nand U14151 (N_14151,N_9128,N_8006);
nor U14152 (N_14152,N_6979,N_5399);
and U14153 (N_14153,N_7886,N_8169);
nand U14154 (N_14154,N_6557,N_7309);
nand U14155 (N_14155,N_6232,N_7863);
nor U14156 (N_14156,N_6695,N_9381);
and U14157 (N_14157,N_6150,N_5179);
nor U14158 (N_14158,N_6619,N_8965);
xor U14159 (N_14159,N_6349,N_8662);
nor U14160 (N_14160,N_8905,N_8099);
nor U14161 (N_14161,N_9686,N_7914);
and U14162 (N_14162,N_6505,N_8068);
nand U14163 (N_14163,N_7873,N_8655);
and U14164 (N_14164,N_7961,N_6671);
nor U14165 (N_14165,N_7089,N_7804);
or U14166 (N_14166,N_5726,N_9732);
or U14167 (N_14167,N_6208,N_6275);
nor U14168 (N_14168,N_7013,N_7840);
or U14169 (N_14169,N_8563,N_6266);
or U14170 (N_14170,N_5109,N_5501);
nor U14171 (N_14171,N_5386,N_7842);
nand U14172 (N_14172,N_7335,N_8498);
and U14173 (N_14173,N_6276,N_6264);
nand U14174 (N_14174,N_9898,N_6790);
nand U14175 (N_14175,N_5292,N_8676);
or U14176 (N_14176,N_5258,N_7877);
and U14177 (N_14177,N_6649,N_9247);
and U14178 (N_14178,N_5252,N_5227);
nor U14179 (N_14179,N_6586,N_5287);
and U14180 (N_14180,N_7695,N_5728);
and U14181 (N_14181,N_9716,N_7447);
and U14182 (N_14182,N_6700,N_6871);
nor U14183 (N_14183,N_9949,N_5319);
and U14184 (N_14184,N_9842,N_8108);
nor U14185 (N_14185,N_6429,N_6414);
or U14186 (N_14186,N_8796,N_6684);
and U14187 (N_14187,N_7617,N_8753);
or U14188 (N_14188,N_7915,N_6661);
nor U14189 (N_14189,N_6708,N_7557);
nand U14190 (N_14190,N_5144,N_6001);
nor U14191 (N_14191,N_7948,N_8896);
nor U14192 (N_14192,N_6307,N_6015);
and U14193 (N_14193,N_7565,N_8772);
nor U14194 (N_14194,N_6669,N_9180);
xnor U14195 (N_14195,N_9348,N_7717);
and U14196 (N_14196,N_6941,N_8598);
nor U14197 (N_14197,N_5896,N_8457);
nor U14198 (N_14198,N_5460,N_5248);
nor U14199 (N_14199,N_5500,N_7452);
nand U14200 (N_14200,N_7153,N_8081);
nand U14201 (N_14201,N_7270,N_6367);
nor U14202 (N_14202,N_9871,N_9124);
nand U14203 (N_14203,N_9303,N_5190);
nand U14204 (N_14204,N_7908,N_6813);
nor U14205 (N_14205,N_9595,N_9563);
and U14206 (N_14206,N_7165,N_7918);
and U14207 (N_14207,N_6259,N_7393);
and U14208 (N_14208,N_9686,N_6674);
and U14209 (N_14209,N_5662,N_9461);
and U14210 (N_14210,N_5800,N_7117);
nand U14211 (N_14211,N_9132,N_5939);
nor U14212 (N_14212,N_7125,N_5710);
nor U14213 (N_14213,N_5833,N_8195);
nor U14214 (N_14214,N_7589,N_7533);
or U14215 (N_14215,N_8077,N_7680);
nor U14216 (N_14216,N_8761,N_9387);
and U14217 (N_14217,N_9567,N_5172);
nor U14218 (N_14218,N_9661,N_6663);
nand U14219 (N_14219,N_8155,N_8990);
and U14220 (N_14220,N_6968,N_9416);
nor U14221 (N_14221,N_5002,N_5286);
or U14222 (N_14222,N_6294,N_6199);
or U14223 (N_14223,N_8388,N_7536);
and U14224 (N_14224,N_7107,N_8897);
nand U14225 (N_14225,N_8305,N_7309);
nor U14226 (N_14226,N_9718,N_7608);
nand U14227 (N_14227,N_6288,N_5545);
nor U14228 (N_14228,N_9794,N_5443);
nor U14229 (N_14229,N_8537,N_8899);
nor U14230 (N_14230,N_5189,N_9545);
nor U14231 (N_14231,N_8059,N_7696);
nand U14232 (N_14232,N_8320,N_7605);
nor U14233 (N_14233,N_5306,N_8876);
and U14234 (N_14234,N_7264,N_5038);
and U14235 (N_14235,N_9980,N_7566);
nand U14236 (N_14236,N_6388,N_8905);
nand U14237 (N_14237,N_6825,N_6957);
nor U14238 (N_14238,N_9668,N_7584);
or U14239 (N_14239,N_5346,N_6434);
nor U14240 (N_14240,N_5828,N_6553);
or U14241 (N_14241,N_9652,N_7162);
and U14242 (N_14242,N_5974,N_6411);
and U14243 (N_14243,N_8088,N_9802);
nand U14244 (N_14244,N_5910,N_9698);
and U14245 (N_14245,N_7738,N_6196);
nand U14246 (N_14246,N_7214,N_7501);
and U14247 (N_14247,N_5374,N_8924);
and U14248 (N_14248,N_6951,N_6369);
nor U14249 (N_14249,N_5962,N_8896);
nand U14250 (N_14250,N_7384,N_9555);
or U14251 (N_14251,N_9726,N_9252);
nand U14252 (N_14252,N_8630,N_8081);
or U14253 (N_14253,N_8132,N_8639);
nor U14254 (N_14254,N_5026,N_8212);
nor U14255 (N_14255,N_8336,N_7164);
or U14256 (N_14256,N_7599,N_6473);
nor U14257 (N_14257,N_9134,N_9593);
and U14258 (N_14258,N_8992,N_8873);
nand U14259 (N_14259,N_7722,N_6533);
and U14260 (N_14260,N_5592,N_6432);
nand U14261 (N_14261,N_5034,N_8261);
nand U14262 (N_14262,N_9542,N_7190);
nor U14263 (N_14263,N_8550,N_7898);
nand U14264 (N_14264,N_6286,N_7941);
nor U14265 (N_14265,N_7129,N_7076);
nand U14266 (N_14266,N_9785,N_7620);
or U14267 (N_14267,N_7278,N_5121);
nor U14268 (N_14268,N_6698,N_8139);
nand U14269 (N_14269,N_9731,N_9664);
and U14270 (N_14270,N_5046,N_8153);
and U14271 (N_14271,N_7938,N_7387);
nor U14272 (N_14272,N_5801,N_6792);
and U14273 (N_14273,N_6555,N_5196);
nor U14274 (N_14274,N_8056,N_8951);
nor U14275 (N_14275,N_6188,N_9293);
and U14276 (N_14276,N_5868,N_8383);
and U14277 (N_14277,N_8656,N_9536);
or U14278 (N_14278,N_5349,N_6702);
nor U14279 (N_14279,N_9955,N_6542);
nor U14280 (N_14280,N_6143,N_8361);
nor U14281 (N_14281,N_9994,N_6232);
nand U14282 (N_14282,N_9780,N_5709);
or U14283 (N_14283,N_5263,N_7368);
nor U14284 (N_14284,N_8098,N_9671);
nand U14285 (N_14285,N_6820,N_7055);
and U14286 (N_14286,N_9997,N_6879);
nand U14287 (N_14287,N_7798,N_9016);
nor U14288 (N_14288,N_6844,N_8167);
nor U14289 (N_14289,N_5671,N_8573);
nor U14290 (N_14290,N_6625,N_7419);
nor U14291 (N_14291,N_8782,N_8579);
and U14292 (N_14292,N_9162,N_9645);
nor U14293 (N_14293,N_6013,N_8822);
or U14294 (N_14294,N_7383,N_9793);
and U14295 (N_14295,N_8879,N_5485);
and U14296 (N_14296,N_7658,N_8657);
nand U14297 (N_14297,N_8462,N_8206);
nand U14298 (N_14298,N_9895,N_8006);
nand U14299 (N_14299,N_6592,N_9913);
or U14300 (N_14300,N_7229,N_9602);
nand U14301 (N_14301,N_7706,N_8479);
and U14302 (N_14302,N_9301,N_7213);
nand U14303 (N_14303,N_5490,N_6544);
nand U14304 (N_14304,N_7734,N_9850);
nor U14305 (N_14305,N_6195,N_5987);
nor U14306 (N_14306,N_8771,N_7004);
or U14307 (N_14307,N_9681,N_8230);
and U14308 (N_14308,N_9126,N_9788);
nand U14309 (N_14309,N_8798,N_8504);
xnor U14310 (N_14310,N_9743,N_8514);
nand U14311 (N_14311,N_5632,N_5631);
and U14312 (N_14312,N_9720,N_8909);
nand U14313 (N_14313,N_8849,N_8152);
and U14314 (N_14314,N_5512,N_7248);
nand U14315 (N_14315,N_5216,N_6391);
nor U14316 (N_14316,N_9344,N_8820);
or U14317 (N_14317,N_7838,N_8794);
or U14318 (N_14318,N_7566,N_7372);
or U14319 (N_14319,N_5815,N_6573);
nand U14320 (N_14320,N_5245,N_8829);
and U14321 (N_14321,N_9934,N_9944);
nand U14322 (N_14322,N_7534,N_5711);
or U14323 (N_14323,N_9150,N_7244);
or U14324 (N_14324,N_7026,N_5292);
nor U14325 (N_14325,N_9893,N_8744);
nor U14326 (N_14326,N_8982,N_5454);
nand U14327 (N_14327,N_5707,N_7022);
and U14328 (N_14328,N_7791,N_5685);
and U14329 (N_14329,N_5438,N_6831);
nand U14330 (N_14330,N_7928,N_6917);
and U14331 (N_14331,N_9801,N_7266);
nor U14332 (N_14332,N_5519,N_5826);
nand U14333 (N_14333,N_6047,N_7825);
nor U14334 (N_14334,N_7555,N_9059);
or U14335 (N_14335,N_6062,N_7275);
nor U14336 (N_14336,N_9678,N_7783);
xnor U14337 (N_14337,N_5392,N_8587);
and U14338 (N_14338,N_9606,N_9445);
nor U14339 (N_14339,N_9796,N_8388);
or U14340 (N_14340,N_9136,N_6538);
or U14341 (N_14341,N_6372,N_5828);
and U14342 (N_14342,N_5974,N_9053);
nor U14343 (N_14343,N_7690,N_6202);
nor U14344 (N_14344,N_8890,N_9433);
or U14345 (N_14345,N_8383,N_6488);
nor U14346 (N_14346,N_7050,N_5028);
nand U14347 (N_14347,N_9089,N_6384);
nand U14348 (N_14348,N_5546,N_6924);
or U14349 (N_14349,N_5598,N_9215);
or U14350 (N_14350,N_6704,N_7889);
or U14351 (N_14351,N_8422,N_6965);
and U14352 (N_14352,N_9409,N_8351);
nor U14353 (N_14353,N_6770,N_6748);
or U14354 (N_14354,N_5967,N_9732);
nand U14355 (N_14355,N_5391,N_5257);
nor U14356 (N_14356,N_8144,N_7899);
nor U14357 (N_14357,N_8748,N_6000);
and U14358 (N_14358,N_5835,N_7543);
nor U14359 (N_14359,N_6981,N_6698);
nand U14360 (N_14360,N_7151,N_6105);
and U14361 (N_14361,N_6262,N_5880);
and U14362 (N_14362,N_7583,N_8071);
or U14363 (N_14363,N_5546,N_8185);
nor U14364 (N_14364,N_8523,N_7332);
nand U14365 (N_14365,N_6934,N_9634);
nand U14366 (N_14366,N_9198,N_9614);
and U14367 (N_14367,N_5405,N_5374);
nor U14368 (N_14368,N_5283,N_7111);
and U14369 (N_14369,N_9564,N_8933);
and U14370 (N_14370,N_7454,N_6258);
or U14371 (N_14371,N_9674,N_7977);
nor U14372 (N_14372,N_8014,N_7496);
nor U14373 (N_14373,N_5672,N_5919);
and U14374 (N_14374,N_9014,N_7589);
or U14375 (N_14375,N_6615,N_7959);
nor U14376 (N_14376,N_8708,N_5815);
and U14377 (N_14377,N_8781,N_7242);
or U14378 (N_14378,N_9105,N_8056);
nor U14379 (N_14379,N_8881,N_6862);
and U14380 (N_14380,N_5773,N_9292);
nand U14381 (N_14381,N_7723,N_9710);
or U14382 (N_14382,N_5743,N_9372);
nand U14383 (N_14383,N_7566,N_9912);
nand U14384 (N_14384,N_7693,N_8944);
nand U14385 (N_14385,N_8711,N_7190);
and U14386 (N_14386,N_8444,N_7668);
and U14387 (N_14387,N_7707,N_7388);
and U14388 (N_14388,N_8396,N_9375);
nor U14389 (N_14389,N_6312,N_7165);
nand U14390 (N_14390,N_9345,N_7540);
or U14391 (N_14391,N_5050,N_7858);
nand U14392 (N_14392,N_6613,N_5277);
or U14393 (N_14393,N_7246,N_6790);
or U14394 (N_14394,N_6118,N_9416);
and U14395 (N_14395,N_8341,N_8573);
and U14396 (N_14396,N_6642,N_7758);
nor U14397 (N_14397,N_5713,N_5302);
nor U14398 (N_14398,N_8291,N_8796);
nand U14399 (N_14399,N_9628,N_6726);
nor U14400 (N_14400,N_8666,N_8761);
or U14401 (N_14401,N_7074,N_9810);
and U14402 (N_14402,N_6903,N_9735);
or U14403 (N_14403,N_8883,N_9272);
nor U14404 (N_14404,N_8244,N_9284);
or U14405 (N_14405,N_9623,N_5682);
nand U14406 (N_14406,N_6173,N_5604);
nand U14407 (N_14407,N_5501,N_7167);
nor U14408 (N_14408,N_7015,N_5935);
and U14409 (N_14409,N_6672,N_7164);
and U14410 (N_14410,N_6652,N_6761);
or U14411 (N_14411,N_6793,N_5549);
and U14412 (N_14412,N_9582,N_7010);
nand U14413 (N_14413,N_8051,N_7258);
or U14414 (N_14414,N_7913,N_5850);
or U14415 (N_14415,N_5095,N_7572);
nand U14416 (N_14416,N_9011,N_9572);
nand U14417 (N_14417,N_6484,N_6926);
nand U14418 (N_14418,N_7582,N_6904);
nand U14419 (N_14419,N_8320,N_6394);
nand U14420 (N_14420,N_5846,N_9710);
and U14421 (N_14421,N_8716,N_8605);
or U14422 (N_14422,N_8239,N_9036);
nand U14423 (N_14423,N_8884,N_7468);
or U14424 (N_14424,N_8468,N_8182);
and U14425 (N_14425,N_6809,N_5901);
nor U14426 (N_14426,N_9538,N_5783);
or U14427 (N_14427,N_8716,N_6812);
or U14428 (N_14428,N_8035,N_6406);
and U14429 (N_14429,N_7650,N_5011);
or U14430 (N_14430,N_6931,N_5583);
nor U14431 (N_14431,N_6515,N_8740);
and U14432 (N_14432,N_8047,N_5072);
nor U14433 (N_14433,N_7716,N_5609);
and U14434 (N_14434,N_7394,N_6764);
and U14435 (N_14435,N_5438,N_8538);
nand U14436 (N_14436,N_7817,N_6398);
or U14437 (N_14437,N_7987,N_6195);
nand U14438 (N_14438,N_9620,N_7597);
nand U14439 (N_14439,N_9475,N_6716);
and U14440 (N_14440,N_8246,N_8202);
or U14441 (N_14441,N_5265,N_6811);
or U14442 (N_14442,N_8492,N_8968);
nor U14443 (N_14443,N_6476,N_8043);
nor U14444 (N_14444,N_7077,N_7830);
and U14445 (N_14445,N_5497,N_8121);
nor U14446 (N_14446,N_9559,N_6051);
nand U14447 (N_14447,N_6778,N_7959);
nor U14448 (N_14448,N_9917,N_9317);
nor U14449 (N_14449,N_9148,N_5463);
nand U14450 (N_14450,N_8689,N_8645);
nand U14451 (N_14451,N_6623,N_8118);
nand U14452 (N_14452,N_9142,N_7455);
and U14453 (N_14453,N_6850,N_6306);
or U14454 (N_14454,N_5225,N_8535);
nor U14455 (N_14455,N_6477,N_5145);
nor U14456 (N_14456,N_8951,N_9597);
or U14457 (N_14457,N_5091,N_8421);
nand U14458 (N_14458,N_6532,N_9574);
and U14459 (N_14459,N_9989,N_8896);
or U14460 (N_14460,N_8861,N_5812);
or U14461 (N_14461,N_8030,N_5687);
or U14462 (N_14462,N_7631,N_7624);
nor U14463 (N_14463,N_9755,N_6833);
or U14464 (N_14464,N_6971,N_6961);
nor U14465 (N_14465,N_8553,N_8494);
and U14466 (N_14466,N_8674,N_6631);
nor U14467 (N_14467,N_8357,N_8427);
nor U14468 (N_14468,N_5693,N_7397);
nand U14469 (N_14469,N_6593,N_8651);
nand U14470 (N_14470,N_5058,N_8320);
nor U14471 (N_14471,N_9485,N_8923);
nand U14472 (N_14472,N_8089,N_8638);
nand U14473 (N_14473,N_8066,N_6596);
and U14474 (N_14474,N_7497,N_9634);
nor U14475 (N_14475,N_6094,N_8935);
and U14476 (N_14476,N_9528,N_8364);
nand U14477 (N_14477,N_8689,N_7796);
nand U14478 (N_14478,N_9483,N_9128);
or U14479 (N_14479,N_6993,N_5864);
nand U14480 (N_14480,N_6433,N_8594);
or U14481 (N_14481,N_5820,N_5112);
or U14482 (N_14482,N_9067,N_9426);
nor U14483 (N_14483,N_7254,N_9131);
or U14484 (N_14484,N_5328,N_7615);
or U14485 (N_14485,N_5354,N_6931);
or U14486 (N_14486,N_7673,N_8396);
or U14487 (N_14487,N_5407,N_6978);
or U14488 (N_14488,N_7531,N_6397);
and U14489 (N_14489,N_9906,N_6634);
or U14490 (N_14490,N_6292,N_6801);
and U14491 (N_14491,N_8548,N_6153);
nand U14492 (N_14492,N_9254,N_7064);
and U14493 (N_14493,N_6904,N_9942);
or U14494 (N_14494,N_7088,N_6819);
nor U14495 (N_14495,N_8192,N_9318);
and U14496 (N_14496,N_6826,N_6360);
and U14497 (N_14497,N_9226,N_6424);
or U14498 (N_14498,N_7830,N_8096);
nor U14499 (N_14499,N_5129,N_9698);
nor U14500 (N_14500,N_6197,N_9335);
nor U14501 (N_14501,N_8580,N_9807);
or U14502 (N_14502,N_5770,N_9580);
and U14503 (N_14503,N_6255,N_8176);
and U14504 (N_14504,N_5117,N_6928);
and U14505 (N_14505,N_5286,N_8665);
and U14506 (N_14506,N_6623,N_6855);
and U14507 (N_14507,N_5608,N_6958);
nor U14508 (N_14508,N_5258,N_6325);
or U14509 (N_14509,N_5797,N_8581);
nand U14510 (N_14510,N_9914,N_6839);
and U14511 (N_14511,N_6157,N_7964);
nand U14512 (N_14512,N_9990,N_5949);
and U14513 (N_14513,N_8046,N_8359);
nor U14514 (N_14514,N_7674,N_8223);
nor U14515 (N_14515,N_7004,N_9051);
or U14516 (N_14516,N_7916,N_8910);
and U14517 (N_14517,N_9083,N_8483);
and U14518 (N_14518,N_8077,N_7079);
nor U14519 (N_14519,N_5465,N_6189);
nor U14520 (N_14520,N_6346,N_7146);
or U14521 (N_14521,N_8141,N_5941);
nor U14522 (N_14522,N_6771,N_9532);
or U14523 (N_14523,N_6376,N_8166);
nor U14524 (N_14524,N_9277,N_6652);
nor U14525 (N_14525,N_9647,N_6849);
nor U14526 (N_14526,N_5825,N_6122);
and U14527 (N_14527,N_8356,N_8156);
nor U14528 (N_14528,N_8711,N_5925);
and U14529 (N_14529,N_8896,N_9143);
nand U14530 (N_14530,N_8617,N_9291);
or U14531 (N_14531,N_7975,N_6491);
or U14532 (N_14532,N_8253,N_9880);
nand U14533 (N_14533,N_9635,N_7298);
or U14534 (N_14534,N_7604,N_9342);
nand U14535 (N_14535,N_6435,N_6463);
and U14536 (N_14536,N_6388,N_5489);
nor U14537 (N_14537,N_9431,N_7809);
xnor U14538 (N_14538,N_7371,N_7981);
or U14539 (N_14539,N_8325,N_7684);
nand U14540 (N_14540,N_6720,N_5812);
and U14541 (N_14541,N_9897,N_7308);
and U14542 (N_14542,N_8632,N_8025);
nand U14543 (N_14543,N_8376,N_7175);
and U14544 (N_14544,N_6116,N_7642);
or U14545 (N_14545,N_8019,N_9085);
nor U14546 (N_14546,N_8182,N_5513);
or U14547 (N_14547,N_7997,N_7920);
nand U14548 (N_14548,N_7652,N_5400);
and U14549 (N_14549,N_9796,N_9358);
nor U14550 (N_14550,N_8502,N_8235);
or U14551 (N_14551,N_8582,N_8010);
or U14552 (N_14552,N_7785,N_9998);
or U14553 (N_14553,N_6703,N_5192);
nand U14554 (N_14554,N_5579,N_5950);
nor U14555 (N_14555,N_9663,N_8987);
and U14556 (N_14556,N_8021,N_8232);
nand U14557 (N_14557,N_6048,N_6874);
or U14558 (N_14558,N_8414,N_5500);
or U14559 (N_14559,N_8897,N_6729);
nand U14560 (N_14560,N_8037,N_8948);
and U14561 (N_14561,N_9867,N_7770);
nor U14562 (N_14562,N_9736,N_8426);
nand U14563 (N_14563,N_8359,N_5610);
nand U14564 (N_14564,N_6668,N_7111);
nand U14565 (N_14565,N_6587,N_6426);
and U14566 (N_14566,N_7199,N_8157);
or U14567 (N_14567,N_6977,N_6007);
and U14568 (N_14568,N_7188,N_6034);
nor U14569 (N_14569,N_9620,N_8179);
and U14570 (N_14570,N_8950,N_8376);
or U14571 (N_14571,N_8594,N_6789);
nand U14572 (N_14572,N_9242,N_7346);
nand U14573 (N_14573,N_8118,N_7999);
nor U14574 (N_14574,N_6896,N_7839);
nor U14575 (N_14575,N_7013,N_8491);
and U14576 (N_14576,N_7458,N_8915);
or U14577 (N_14577,N_5681,N_8240);
nor U14578 (N_14578,N_7910,N_6976);
and U14579 (N_14579,N_5306,N_7763);
nand U14580 (N_14580,N_7486,N_8216);
or U14581 (N_14581,N_5495,N_7577);
and U14582 (N_14582,N_7532,N_5569);
nor U14583 (N_14583,N_7151,N_9065);
and U14584 (N_14584,N_7159,N_7222);
or U14585 (N_14585,N_9108,N_6176);
or U14586 (N_14586,N_7660,N_7261);
and U14587 (N_14587,N_6778,N_8713);
and U14588 (N_14588,N_7040,N_9497);
xnor U14589 (N_14589,N_7909,N_5852);
nand U14590 (N_14590,N_6919,N_5393);
nor U14591 (N_14591,N_8509,N_7226);
nand U14592 (N_14592,N_8080,N_8307);
nand U14593 (N_14593,N_5679,N_8247);
nor U14594 (N_14594,N_6136,N_6190);
nand U14595 (N_14595,N_9644,N_7348);
and U14596 (N_14596,N_7017,N_9539);
nand U14597 (N_14597,N_8638,N_9906);
and U14598 (N_14598,N_7107,N_8371);
or U14599 (N_14599,N_9556,N_6594);
or U14600 (N_14600,N_8646,N_6626);
nor U14601 (N_14601,N_5822,N_9341);
nor U14602 (N_14602,N_6921,N_9065);
nand U14603 (N_14603,N_6270,N_7144);
nor U14604 (N_14604,N_7924,N_9822);
or U14605 (N_14605,N_8964,N_6195);
and U14606 (N_14606,N_7405,N_6448);
nand U14607 (N_14607,N_6131,N_9874);
nor U14608 (N_14608,N_7224,N_8937);
and U14609 (N_14609,N_6056,N_8354);
nor U14610 (N_14610,N_6250,N_7803);
or U14611 (N_14611,N_6448,N_9008);
nand U14612 (N_14612,N_6587,N_8661);
or U14613 (N_14613,N_9516,N_7437);
nor U14614 (N_14614,N_5190,N_5673);
or U14615 (N_14615,N_6083,N_6646);
nor U14616 (N_14616,N_6462,N_7582);
nor U14617 (N_14617,N_6816,N_6680);
nand U14618 (N_14618,N_5604,N_6495);
nor U14619 (N_14619,N_5987,N_9273);
nand U14620 (N_14620,N_8229,N_6691);
nor U14621 (N_14621,N_9064,N_8298);
and U14622 (N_14622,N_9374,N_9676);
and U14623 (N_14623,N_8725,N_8076);
or U14624 (N_14624,N_7755,N_6185);
or U14625 (N_14625,N_6455,N_7653);
and U14626 (N_14626,N_9850,N_7878);
and U14627 (N_14627,N_8979,N_6393);
nand U14628 (N_14628,N_7342,N_9911);
or U14629 (N_14629,N_7257,N_8030);
or U14630 (N_14630,N_5281,N_5724);
nor U14631 (N_14631,N_5801,N_6256);
and U14632 (N_14632,N_5250,N_8259);
or U14633 (N_14633,N_8009,N_6112);
and U14634 (N_14634,N_8339,N_5754);
nor U14635 (N_14635,N_8099,N_8709);
and U14636 (N_14636,N_9413,N_9744);
and U14637 (N_14637,N_9873,N_6621);
nand U14638 (N_14638,N_6027,N_6123);
and U14639 (N_14639,N_6110,N_7996);
xnor U14640 (N_14640,N_8758,N_7401);
and U14641 (N_14641,N_9628,N_5589);
or U14642 (N_14642,N_5931,N_5337);
nand U14643 (N_14643,N_5695,N_5260);
nand U14644 (N_14644,N_9646,N_7906);
or U14645 (N_14645,N_9082,N_5627);
or U14646 (N_14646,N_9159,N_6196);
and U14647 (N_14647,N_8989,N_9834);
and U14648 (N_14648,N_9119,N_6320);
nand U14649 (N_14649,N_8369,N_5309);
and U14650 (N_14650,N_7032,N_8546);
nor U14651 (N_14651,N_6216,N_7486);
or U14652 (N_14652,N_5455,N_8593);
and U14653 (N_14653,N_8050,N_8342);
xnor U14654 (N_14654,N_9686,N_6673);
nor U14655 (N_14655,N_7339,N_5790);
or U14656 (N_14656,N_5095,N_6875);
or U14657 (N_14657,N_5006,N_6976);
nand U14658 (N_14658,N_5900,N_9576);
nand U14659 (N_14659,N_9984,N_7648);
nand U14660 (N_14660,N_5127,N_9001);
nor U14661 (N_14661,N_6260,N_7108);
and U14662 (N_14662,N_6623,N_6471);
or U14663 (N_14663,N_7818,N_9695);
and U14664 (N_14664,N_8633,N_9681);
nor U14665 (N_14665,N_6971,N_5539);
nor U14666 (N_14666,N_7832,N_8131);
or U14667 (N_14667,N_5871,N_7150);
or U14668 (N_14668,N_5068,N_6001);
or U14669 (N_14669,N_5553,N_8233);
and U14670 (N_14670,N_6430,N_9952);
nor U14671 (N_14671,N_5893,N_8586);
and U14672 (N_14672,N_9813,N_7177);
and U14673 (N_14673,N_9403,N_6133);
nand U14674 (N_14674,N_5980,N_8344);
nor U14675 (N_14675,N_7030,N_6065);
or U14676 (N_14676,N_5895,N_7062);
nand U14677 (N_14677,N_7333,N_5426);
and U14678 (N_14678,N_9046,N_9170);
nor U14679 (N_14679,N_7139,N_6693);
nand U14680 (N_14680,N_8625,N_9865);
nand U14681 (N_14681,N_5777,N_5660);
and U14682 (N_14682,N_8369,N_8291);
and U14683 (N_14683,N_7147,N_5138);
and U14684 (N_14684,N_7695,N_7160);
or U14685 (N_14685,N_5356,N_5158);
and U14686 (N_14686,N_7532,N_5207);
or U14687 (N_14687,N_9684,N_7654);
nand U14688 (N_14688,N_6116,N_7063);
and U14689 (N_14689,N_5429,N_8556);
nor U14690 (N_14690,N_9576,N_9894);
nand U14691 (N_14691,N_8056,N_8611);
nand U14692 (N_14692,N_5957,N_7438);
nand U14693 (N_14693,N_7812,N_8750);
and U14694 (N_14694,N_8279,N_5540);
and U14695 (N_14695,N_8826,N_5381);
or U14696 (N_14696,N_8289,N_7253);
and U14697 (N_14697,N_5416,N_9882);
nand U14698 (N_14698,N_6776,N_7843);
or U14699 (N_14699,N_9179,N_9520);
nor U14700 (N_14700,N_5085,N_7582);
and U14701 (N_14701,N_7554,N_5076);
or U14702 (N_14702,N_5229,N_7506);
nor U14703 (N_14703,N_9134,N_7047);
or U14704 (N_14704,N_9201,N_7273);
nand U14705 (N_14705,N_7907,N_9097);
and U14706 (N_14706,N_6724,N_9975);
or U14707 (N_14707,N_9164,N_9517);
nand U14708 (N_14708,N_8541,N_5423);
or U14709 (N_14709,N_8130,N_5177);
and U14710 (N_14710,N_5828,N_9744);
nor U14711 (N_14711,N_7256,N_8688);
and U14712 (N_14712,N_5090,N_6636);
or U14713 (N_14713,N_8333,N_8123);
or U14714 (N_14714,N_9305,N_9724);
nor U14715 (N_14715,N_7233,N_7719);
nand U14716 (N_14716,N_7950,N_6724);
nand U14717 (N_14717,N_8078,N_8387);
or U14718 (N_14718,N_8216,N_6316);
nor U14719 (N_14719,N_7580,N_7052);
and U14720 (N_14720,N_8812,N_5813);
or U14721 (N_14721,N_6525,N_9303);
and U14722 (N_14722,N_8346,N_5353);
nand U14723 (N_14723,N_9776,N_5007);
and U14724 (N_14724,N_7591,N_7571);
nand U14725 (N_14725,N_5297,N_7730);
or U14726 (N_14726,N_9076,N_7223);
nand U14727 (N_14727,N_8953,N_6863);
and U14728 (N_14728,N_8011,N_5433);
nand U14729 (N_14729,N_7561,N_9788);
nor U14730 (N_14730,N_8559,N_9355);
nand U14731 (N_14731,N_6990,N_7250);
nand U14732 (N_14732,N_8633,N_9784);
xor U14733 (N_14733,N_9772,N_5598);
or U14734 (N_14734,N_5763,N_5946);
and U14735 (N_14735,N_5095,N_5077);
nand U14736 (N_14736,N_6909,N_5350);
nor U14737 (N_14737,N_8028,N_5162);
nor U14738 (N_14738,N_5216,N_5093);
and U14739 (N_14739,N_9963,N_9259);
nand U14740 (N_14740,N_5488,N_9963);
or U14741 (N_14741,N_9076,N_7661);
or U14742 (N_14742,N_5909,N_7936);
nand U14743 (N_14743,N_6186,N_9201);
nor U14744 (N_14744,N_5813,N_6560);
nor U14745 (N_14745,N_5426,N_5808);
or U14746 (N_14746,N_8879,N_7283);
and U14747 (N_14747,N_8830,N_7750);
nand U14748 (N_14748,N_7448,N_7371);
nand U14749 (N_14749,N_7355,N_7762);
nor U14750 (N_14750,N_8952,N_6442);
nor U14751 (N_14751,N_9693,N_9172);
nor U14752 (N_14752,N_7442,N_6249);
or U14753 (N_14753,N_6354,N_9165);
nor U14754 (N_14754,N_7590,N_6036);
nor U14755 (N_14755,N_8780,N_9863);
nor U14756 (N_14756,N_9082,N_6586);
xor U14757 (N_14757,N_8068,N_5691);
nor U14758 (N_14758,N_6476,N_6495);
or U14759 (N_14759,N_6400,N_5427);
nand U14760 (N_14760,N_6274,N_8118);
or U14761 (N_14761,N_7216,N_6380);
or U14762 (N_14762,N_9348,N_6686);
nand U14763 (N_14763,N_6141,N_9311);
or U14764 (N_14764,N_6666,N_5222);
and U14765 (N_14765,N_7275,N_7774);
nor U14766 (N_14766,N_9148,N_5423);
and U14767 (N_14767,N_7015,N_6289);
nor U14768 (N_14768,N_8757,N_6811);
nand U14769 (N_14769,N_8263,N_9650);
and U14770 (N_14770,N_9327,N_7942);
and U14771 (N_14771,N_8435,N_8976);
or U14772 (N_14772,N_7798,N_8169);
or U14773 (N_14773,N_7672,N_6423);
nor U14774 (N_14774,N_9754,N_6361);
and U14775 (N_14775,N_6697,N_5287);
nand U14776 (N_14776,N_7521,N_9672);
nor U14777 (N_14777,N_6632,N_8044);
and U14778 (N_14778,N_5652,N_8951);
nor U14779 (N_14779,N_6684,N_5721);
nand U14780 (N_14780,N_8230,N_5078);
and U14781 (N_14781,N_7102,N_7140);
nor U14782 (N_14782,N_5152,N_8955);
nand U14783 (N_14783,N_9946,N_9392);
and U14784 (N_14784,N_6506,N_8800);
nand U14785 (N_14785,N_5293,N_9075);
nor U14786 (N_14786,N_9648,N_6163);
nor U14787 (N_14787,N_5421,N_8901);
and U14788 (N_14788,N_8401,N_5219);
nand U14789 (N_14789,N_6109,N_6490);
nor U14790 (N_14790,N_5924,N_8608);
nor U14791 (N_14791,N_7477,N_5283);
and U14792 (N_14792,N_5319,N_5307);
nand U14793 (N_14793,N_9528,N_8812);
nor U14794 (N_14794,N_6148,N_8621);
or U14795 (N_14795,N_7038,N_8421);
or U14796 (N_14796,N_8308,N_8368);
nor U14797 (N_14797,N_9451,N_7412);
and U14798 (N_14798,N_8773,N_9147);
nand U14799 (N_14799,N_8531,N_8038);
or U14800 (N_14800,N_6952,N_5344);
nand U14801 (N_14801,N_9487,N_9405);
nand U14802 (N_14802,N_9332,N_7362);
or U14803 (N_14803,N_6175,N_9942);
or U14804 (N_14804,N_9988,N_6918);
nor U14805 (N_14805,N_5516,N_9415);
nor U14806 (N_14806,N_8624,N_9685);
or U14807 (N_14807,N_7278,N_5834);
and U14808 (N_14808,N_5496,N_7477);
nor U14809 (N_14809,N_5432,N_8761);
or U14810 (N_14810,N_6725,N_5150);
or U14811 (N_14811,N_5414,N_8175);
nand U14812 (N_14812,N_9730,N_6863);
nand U14813 (N_14813,N_8095,N_7032);
or U14814 (N_14814,N_6680,N_6725);
nand U14815 (N_14815,N_8888,N_9566);
or U14816 (N_14816,N_9415,N_5540);
and U14817 (N_14817,N_6715,N_5366);
and U14818 (N_14818,N_7927,N_5927);
nor U14819 (N_14819,N_8964,N_6935);
nand U14820 (N_14820,N_7032,N_5790);
or U14821 (N_14821,N_7555,N_9280);
nand U14822 (N_14822,N_8811,N_9462);
nor U14823 (N_14823,N_8350,N_5652);
nor U14824 (N_14824,N_9169,N_9323);
and U14825 (N_14825,N_8568,N_8420);
and U14826 (N_14826,N_7043,N_8087);
nor U14827 (N_14827,N_8881,N_7852);
nand U14828 (N_14828,N_7799,N_9669);
and U14829 (N_14829,N_9632,N_6613);
nor U14830 (N_14830,N_9360,N_9819);
nand U14831 (N_14831,N_7417,N_9909);
nor U14832 (N_14832,N_7105,N_6124);
nand U14833 (N_14833,N_9066,N_6091);
or U14834 (N_14834,N_8262,N_7721);
and U14835 (N_14835,N_5727,N_7100);
or U14836 (N_14836,N_7730,N_6190);
nand U14837 (N_14837,N_5129,N_7001);
nand U14838 (N_14838,N_9322,N_8934);
nor U14839 (N_14839,N_8313,N_9417);
nand U14840 (N_14840,N_7418,N_7238);
nor U14841 (N_14841,N_9915,N_5649);
and U14842 (N_14842,N_5479,N_5066);
and U14843 (N_14843,N_6709,N_5116);
or U14844 (N_14844,N_9445,N_8926);
nor U14845 (N_14845,N_9887,N_6251);
and U14846 (N_14846,N_9346,N_8972);
nor U14847 (N_14847,N_8102,N_9088);
and U14848 (N_14848,N_8630,N_9988);
or U14849 (N_14849,N_7414,N_7422);
nand U14850 (N_14850,N_6263,N_6574);
nand U14851 (N_14851,N_7887,N_9664);
nor U14852 (N_14852,N_9779,N_8747);
and U14853 (N_14853,N_8267,N_7605);
or U14854 (N_14854,N_5148,N_6648);
nand U14855 (N_14855,N_7866,N_6051);
or U14856 (N_14856,N_5198,N_9653);
nand U14857 (N_14857,N_9239,N_6217);
nand U14858 (N_14858,N_7701,N_9706);
nand U14859 (N_14859,N_8428,N_7111);
or U14860 (N_14860,N_6367,N_9631);
nor U14861 (N_14861,N_6452,N_9392);
nor U14862 (N_14862,N_8876,N_7967);
nand U14863 (N_14863,N_8464,N_7730);
or U14864 (N_14864,N_9122,N_8654);
or U14865 (N_14865,N_6544,N_8360);
and U14866 (N_14866,N_5915,N_9839);
nor U14867 (N_14867,N_6905,N_8368);
nand U14868 (N_14868,N_6182,N_6869);
or U14869 (N_14869,N_6140,N_5959);
and U14870 (N_14870,N_9465,N_5124);
nor U14871 (N_14871,N_5274,N_9827);
and U14872 (N_14872,N_8511,N_7071);
nor U14873 (N_14873,N_7598,N_7009);
nand U14874 (N_14874,N_9899,N_5303);
nand U14875 (N_14875,N_9946,N_7044);
or U14876 (N_14876,N_9099,N_5831);
nand U14877 (N_14877,N_8833,N_7478);
or U14878 (N_14878,N_5841,N_6399);
nor U14879 (N_14879,N_8203,N_9575);
or U14880 (N_14880,N_6790,N_6611);
nand U14881 (N_14881,N_6219,N_9707);
or U14882 (N_14882,N_9459,N_9340);
nand U14883 (N_14883,N_7145,N_8291);
and U14884 (N_14884,N_8886,N_5317);
and U14885 (N_14885,N_9298,N_5600);
nand U14886 (N_14886,N_6805,N_7468);
and U14887 (N_14887,N_8662,N_5317);
and U14888 (N_14888,N_8182,N_9702);
nand U14889 (N_14889,N_5623,N_5008);
or U14890 (N_14890,N_9901,N_9444);
or U14891 (N_14891,N_6086,N_9135);
or U14892 (N_14892,N_8068,N_7789);
nor U14893 (N_14893,N_8106,N_9650);
or U14894 (N_14894,N_8392,N_7660);
or U14895 (N_14895,N_7246,N_9427);
nand U14896 (N_14896,N_9670,N_8465);
and U14897 (N_14897,N_7381,N_9643);
or U14898 (N_14898,N_8560,N_9053);
and U14899 (N_14899,N_5488,N_9686);
and U14900 (N_14900,N_8946,N_5198);
and U14901 (N_14901,N_9565,N_9761);
nor U14902 (N_14902,N_9783,N_5777);
nor U14903 (N_14903,N_9321,N_9619);
or U14904 (N_14904,N_9283,N_6541);
and U14905 (N_14905,N_5344,N_8855);
nand U14906 (N_14906,N_9401,N_6154);
and U14907 (N_14907,N_9387,N_5632);
nor U14908 (N_14908,N_6882,N_5544);
or U14909 (N_14909,N_8125,N_6196);
or U14910 (N_14910,N_7976,N_8647);
and U14911 (N_14911,N_5731,N_6547);
and U14912 (N_14912,N_7955,N_5571);
and U14913 (N_14913,N_9860,N_9268);
nor U14914 (N_14914,N_6739,N_7691);
nor U14915 (N_14915,N_7879,N_5009);
and U14916 (N_14916,N_7031,N_6961);
nand U14917 (N_14917,N_7075,N_6517);
nand U14918 (N_14918,N_6832,N_5792);
nand U14919 (N_14919,N_7386,N_6889);
or U14920 (N_14920,N_6194,N_7766);
nor U14921 (N_14921,N_8076,N_7757);
nor U14922 (N_14922,N_5749,N_9261);
or U14923 (N_14923,N_8393,N_8920);
and U14924 (N_14924,N_6582,N_6469);
nand U14925 (N_14925,N_9024,N_9026);
and U14926 (N_14926,N_6362,N_9076);
nor U14927 (N_14927,N_6124,N_6340);
and U14928 (N_14928,N_6230,N_6910);
or U14929 (N_14929,N_8164,N_8324);
or U14930 (N_14930,N_6150,N_6156);
and U14931 (N_14931,N_7307,N_6846);
nor U14932 (N_14932,N_8214,N_8690);
nand U14933 (N_14933,N_5342,N_9333);
nand U14934 (N_14934,N_9681,N_8250);
nand U14935 (N_14935,N_7673,N_5105);
nand U14936 (N_14936,N_6801,N_5952);
and U14937 (N_14937,N_6087,N_6635);
and U14938 (N_14938,N_8053,N_7845);
nor U14939 (N_14939,N_6544,N_7029);
and U14940 (N_14940,N_6583,N_6539);
or U14941 (N_14941,N_7129,N_6626);
and U14942 (N_14942,N_5367,N_9728);
or U14943 (N_14943,N_7334,N_7505);
and U14944 (N_14944,N_8914,N_7628);
nand U14945 (N_14945,N_6450,N_8326);
nor U14946 (N_14946,N_9302,N_6046);
or U14947 (N_14947,N_8045,N_5220);
nor U14948 (N_14948,N_6460,N_7627);
or U14949 (N_14949,N_8542,N_6862);
and U14950 (N_14950,N_8070,N_6137);
or U14951 (N_14951,N_7020,N_8645);
or U14952 (N_14952,N_8198,N_7668);
or U14953 (N_14953,N_5027,N_5714);
or U14954 (N_14954,N_5651,N_8865);
or U14955 (N_14955,N_6624,N_6645);
or U14956 (N_14956,N_7221,N_9502);
or U14957 (N_14957,N_5765,N_5571);
nor U14958 (N_14958,N_8591,N_8843);
or U14959 (N_14959,N_8622,N_9329);
or U14960 (N_14960,N_7713,N_8546);
and U14961 (N_14961,N_8052,N_8218);
nor U14962 (N_14962,N_6830,N_6806);
nand U14963 (N_14963,N_8750,N_7620);
or U14964 (N_14964,N_5348,N_8093);
and U14965 (N_14965,N_7574,N_8420);
xor U14966 (N_14966,N_8629,N_7646);
nand U14967 (N_14967,N_7087,N_5852);
and U14968 (N_14968,N_7647,N_9051);
nand U14969 (N_14969,N_7330,N_7181);
or U14970 (N_14970,N_9048,N_5355);
or U14971 (N_14971,N_5837,N_9021);
or U14972 (N_14972,N_7776,N_6799);
nor U14973 (N_14973,N_5839,N_6239);
nor U14974 (N_14974,N_9440,N_5694);
or U14975 (N_14975,N_9726,N_9570);
nor U14976 (N_14976,N_6456,N_8979);
nor U14977 (N_14977,N_9538,N_9748);
or U14978 (N_14978,N_8025,N_7688);
and U14979 (N_14979,N_6443,N_5188);
or U14980 (N_14980,N_5161,N_5886);
nand U14981 (N_14981,N_7267,N_8204);
or U14982 (N_14982,N_5469,N_7784);
or U14983 (N_14983,N_8405,N_6392);
nand U14984 (N_14984,N_6824,N_6264);
nand U14985 (N_14985,N_9491,N_7653);
and U14986 (N_14986,N_6240,N_8611);
nor U14987 (N_14987,N_8869,N_5336);
nand U14988 (N_14988,N_8592,N_6207);
nand U14989 (N_14989,N_6625,N_8417);
and U14990 (N_14990,N_7457,N_5274);
or U14991 (N_14991,N_8582,N_5527);
nand U14992 (N_14992,N_8236,N_5247);
nand U14993 (N_14993,N_6312,N_9096);
nor U14994 (N_14994,N_7204,N_7302);
or U14995 (N_14995,N_5538,N_5850);
nand U14996 (N_14996,N_9998,N_8244);
nor U14997 (N_14997,N_8126,N_6113);
nor U14998 (N_14998,N_7630,N_7928);
or U14999 (N_14999,N_9182,N_6148);
nand U15000 (N_15000,N_11656,N_12189);
nand U15001 (N_15001,N_11730,N_13237);
or U15002 (N_15002,N_10625,N_10354);
nor U15003 (N_15003,N_11584,N_12955);
and U15004 (N_15004,N_14293,N_10996);
or U15005 (N_15005,N_10328,N_13456);
and U15006 (N_15006,N_10304,N_10926);
and U15007 (N_15007,N_11694,N_10373);
or U15008 (N_15008,N_14738,N_14660);
nor U15009 (N_15009,N_13881,N_13426);
and U15010 (N_15010,N_13789,N_13411);
nand U15011 (N_15011,N_10013,N_11477);
nor U15012 (N_15012,N_14836,N_13035);
or U15013 (N_15013,N_12765,N_14379);
and U15014 (N_15014,N_10028,N_10042);
nand U15015 (N_15015,N_12799,N_13433);
and U15016 (N_15016,N_12656,N_14462);
or U15017 (N_15017,N_10342,N_14346);
nand U15018 (N_15018,N_13571,N_14850);
nor U15019 (N_15019,N_13765,N_11524);
nor U15020 (N_15020,N_12824,N_10064);
and U15021 (N_15021,N_12355,N_13444);
nor U15022 (N_15022,N_13914,N_10363);
nand U15023 (N_15023,N_14819,N_13125);
nand U15024 (N_15024,N_11707,N_13905);
or U15025 (N_15025,N_10571,N_10254);
nand U15026 (N_15026,N_13590,N_12285);
nand U15027 (N_15027,N_12769,N_11251);
nor U15028 (N_15028,N_12051,N_10447);
nor U15029 (N_15029,N_12046,N_10375);
and U15030 (N_15030,N_11666,N_11916);
nand U15031 (N_15031,N_11057,N_11008);
or U15032 (N_15032,N_12359,N_12144);
nand U15033 (N_15033,N_10728,N_10557);
or U15034 (N_15034,N_12622,N_11897);
xnor U15035 (N_15035,N_14874,N_10259);
or U15036 (N_15036,N_14244,N_13672);
and U15037 (N_15037,N_11580,N_10843);
nor U15038 (N_15038,N_11602,N_13155);
nor U15039 (N_15039,N_10652,N_10924);
and U15040 (N_15040,N_13229,N_12097);
and U15041 (N_15041,N_14133,N_12443);
nor U15042 (N_15042,N_14938,N_11404);
or U15043 (N_15043,N_10885,N_10852);
nor U15044 (N_15044,N_13458,N_11724);
nand U15045 (N_15045,N_13561,N_12791);
nand U15046 (N_15046,N_11984,N_10025);
nand U15047 (N_15047,N_11550,N_12773);
nor U15048 (N_15048,N_10473,N_11114);
and U15049 (N_15049,N_12534,N_14191);
xnor U15050 (N_15050,N_10786,N_11779);
nor U15051 (N_15051,N_10287,N_12269);
or U15052 (N_15052,N_14114,N_12209);
nand U15053 (N_15053,N_12047,N_12204);
and U15054 (N_15054,N_14980,N_11051);
nand U15055 (N_15055,N_12558,N_12075);
nand U15056 (N_15056,N_10832,N_11179);
and U15057 (N_15057,N_11879,N_10070);
nor U15058 (N_15058,N_13546,N_14473);
nor U15059 (N_15059,N_14446,N_11520);
nand U15060 (N_15060,N_12758,N_14219);
and U15061 (N_15061,N_10682,N_10718);
or U15062 (N_15062,N_14677,N_11096);
nand U15063 (N_15063,N_10892,N_10331);
nand U15064 (N_15064,N_11327,N_11507);
and U15065 (N_15065,N_13328,N_12587);
nor U15066 (N_15066,N_13532,N_14782);
nand U15067 (N_15067,N_14882,N_10585);
nand U15068 (N_15068,N_12108,N_14106);
nor U15069 (N_15069,N_10821,N_13732);
and U15070 (N_15070,N_13017,N_13714);
and U15071 (N_15071,N_13564,N_12977);
nor U15072 (N_15072,N_13357,N_13497);
nand U15073 (N_15073,N_10871,N_14008);
nor U15074 (N_15074,N_14924,N_12673);
and U15075 (N_15075,N_10362,N_13390);
and U15076 (N_15076,N_13077,N_14931);
and U15077 (N_15077,N_14117,N_10664);
nand U15078 (N_15078,N_11934,N_10290);
nand U15079 (N_15079,N_14139,N_11444);
nand U15080 (N_15080,N_14072,N_12412);
nand U15081 (N_15081,N_13431,N_11660);
or U15082 (N_15082,N_12055,N_10462);
nor U15083 (N_15083,N_13309,N_13159);
nor U15084 (N_15084,N_13998,N_10492);
nor U15085 (N_15085,N_12542,N_10207);
and U15086 (N_15086,N_14774,N_12211);
nor U15087 (N_15087,N_13629,N_12239);
and U15088 (N_15088,N_13931,N_13953);
and U15089 (N_15089,N_10189,N_12107);
nor U15090 (N_15090,N_13582,N_12631);
nand U15091 (N_15091,N_14189,N_11826);
and U15092 (N_15092,N_10041,N_10299);
nor U15093 (N_15093,N_10910,N_10612);
and U15094 (N_15094,N_13701,N_11955);
or U15095 (N_15095,N_13259,N_12248);
and U15096 (N_15096,N_11437,N_14044);
or U15097 (N_15097,N_12668,N_13432);
nand U15098 (N_15098,N_14640,N_11433);
and U15099 (N_15099,N_11554,N_10534);
nand U15100 (N_15100,N_11812,N_13508);
or U15101 (N_15101,N_11213,N_12585);
nand U15102 (N_15102,N_14406,N_14916);
or U15103 (N_15103,N_10734,N_11195);
nor U15104 (N_15104,N_11918,N_11650);
nor U15105 (N_15105,N_11962,N_12577);
nor U15106 (N_15106,N_14136,N_11242);
nor U15107 (N_15107,N_10601,N_10976);
nand U15108 (N_15108,N_14923,N_12284);
or U15109 (N_15109,N_11162,N_10093);
or U15110 (N_15110,N_11224,N_10168);
nor U15111 (N_15111,N_11170,N_11058);
nand U15112 (N_15112,N_14689,N_13037);
and U15113 (N_15113,N_11727,N_10729);
xnor U15114 (N_15114,N_13145,N_13785);
and U15115 (N_15115,N_14225,N_14342);
and U15116 (N_15116,N_12245,N_10719);
nand U15117 (N_15117,N_14616,N_10243);
nand U15118 (N_15118,N_14273,N_10449);
and U15119 (N_15119,N_14697,N_11490);
nor U15120 (N_15120,N_11546,N_14703);
nand U15121 (N_15121,N_11463,N_13646);
nor U15122 (N_15122,N_14325,N_13831);
and U15123 (N_15123,N_12254,N_13245);
or U15124 (N_15124,N_13522,N_14538);
and U15125 (N_15125,N_12212,N_11377);
or U15126 (N_15126,N_13032,N_13971);
or U15127 (N_15127,N_10182,N_10387);
and U15128 (N_15128,N_13066,N_10886);
xor U15129 (N_15129,N_14474,N_10800);
or U15130 (N_15130,N_13673,N_13584);
or U15131 (N_15131,N_14706,N_10115);
or U15132 (N_15132,N_11809,N_10895);
and U15133 (N_15133,N_12948,N_14213);
or U15134 (N_15134,N_10381,N_10395);
and U15135 (N_15135,N_14339,N_12009);
and U15136 (N_15136,N_12167,N_14130);
nor U15137 (N_15137,N_12506,N_10574);
or U15138 (N_15138,N_14297,N_10099);
xor U15139 (N_15139,N_12807,N_13733);
nand U15140 (N_15140,N_11810,N_11345);
nand U15141 (N_15141,N_12295,N_11940);
nor U15142 (N_15142,N_11359,N_14651);
or U15143 (N_15143,N_13056,N_10079);
nand U15144 (N_15144,N_13791,N_10412);
or U15145 (N_15145,N_11119,N_11022);
nor U15146 (N_15146,N_11418,N_14852);
or U15147 (N_15147,N_12195,N_10106);
nand U15148 (N_15148,N_12404,N_12405);
and U15149 (N_15149,N_13302,N_14613);
and U15150 (N_15150,N_14120,N_10069);
nand U15151 (N_15151,N_13844,N_11850);
or U15152 (N_15152,N_13788,N_14915);
and U15153 (N_15153,N_12532,N_12117);
or U15154 (N_15154,N_11115,N_10994);
or U15155 (N_15155,N_13742,N_13902);
nand U15156 (N_15156,N_13345,N_10993);
and U15157 (N_15157,N_10162,N_12710);
nor U15158 (N_15158,N_14202,N_11732);
or U15159 (N_15159,N_14499,N_13285);
nand U15160 (N_15160,N_13641,N_13869);
and U15161 (N_15161,N_10450,N_11612);
nand U15162 (N_15162,N_11113,N_14003);
or U15163 (N_15163,N_10742,N_10642);
and U15164 (N_15164,N_11691,N_11018);
nand U15165 (N_15165,N_13917,N_10284);
and U15166 (N_15166,N_10679,N_11384);
nand U15167 (N_15167,N_13516,N_14144);
nand U15168 (N_15168,N_11878,N_13787);
or U15169 (N_15169,N_11438,N_12216);
or U15170 (N_15170,N_12401,N_11871);
and U15171 (N_15171,N_13738,N_14283);
nand U15172 (N_15172,N_11798,N_11748);
or U15173 (N_15173,N_12899,N_10442);
and U15174 (N_15174,N_11336,N_12645);
and U15175 (N_15175,N_10399,N_12784);
and U15176 (N_15176,N_10978,N_14833);
nand U15177 (N_15177,N_11606,N_12669);
and U15178 (N_15178,N_10890,N_13545);
and U15179 (N_15179,N_14374,N_14679);
nor U15180 (N_15180,N_13635,N_12941);
and U15181 (N_15181,N_10195,N_10723);
nand U15182 (N_15182,N_10086,N_11079);
nor U15183 (N_15183,N_11501,N_12989);
or U15184 (N_15184,N_13081,N_13779);
and U15185 (N_15185,N_12725,N_13230);
nor U15186 (N_15186,N_12099,N_12711);
or U15187 (N_15187,N_12741,N_12023);
nor U15188 (N_15188,N_14211,N_12070);
nor U15189 (N_15189,N_10253,N_10605);
nand U15190 (N_15190,N_12696,N_13075);
nand U15191 (N_15191,N_11328,N_10181);
xor U15192 (N_15192,N_10623,N_14624);
nor U15193 (N_15193,N_11664,N_10215);
and U15194 (N_15194,N_13303,N_11919);
and U15195 (N_15195,N_11196,N_10797);
or U15196 (N_15196,N_10756,N_14414);
nor U15197 (N_15197,N_11159,N_14308);
or U15198 (N_15198,N_13956,N_13731);
nand U15199 (N_15199,N_13558,N_10113);
nand U15200 (N_15200,N_12984,N_11853);
nand U15201 (N_15201,N_10445,N_11150);
nor U15202 (N_15202,N_12054,N_10527);
nor U15203 (N_15203,N_14444,N_14470);
nand U15204 (N_15204,N_10698,N_12927);
nor U15205 (N_15205,N_12887,N_12383);
nor U15206 (N_15206,N_13148,N_11800);
or U15207 (N_15207,N_11639,N_11402);
and U15208 (N_15208,N_12796,N_10572);
and U15209 (N_15209,N_14585,N_12249);
nand U15210 (N_15210,N_10731,N_12351);
nor U15211 (N_15211,N_12516,N_14386);
nand U15212 (N_15212,N_10114,N_14298);
and U15213 (N_15213,N_14806,N_14242);
or U15214 (N_15214,N_13932,N_11725);
nand U15215 (N_15215,N_10245,N_11396);
nor U15216 (N_15216,N_10884,N_14844);
and U15217 (N_15217,N_11737,N_14927);
and U15218 (N_15218,N_12064,N_14764);
and U15219 (N_15219,N_13815,N_10372);
nor U15220 (N_15220,N_13832,N_12588);
or U15221 (N_15221,N_13270,N_13154);
and U15222 (N_15222,N_14741,N_12568);
or U15223 (N_15223,N_11997,N_11849);
or U15224 (N_15224,N_14231,N_13140);
nor U15225 (N_15225,N_10177,N_14049);
nor U15226 (N_15226,N_12974,N_13517);
nor U15227 (N_15227,N_10861,N_10704);
nor U15228 (N_15228,N_13419,N_12283);
nor U15229 (N_15229,N_12403,N_10736);
nor U15230 (N_15230,N_14509,N_14593);
and U15231 (N_15231,N_13397,N_12502);
and U15232 (N_15232,N_12485,N_12119);
nor U15233 (N_15233,N_13033,N_14055);
nand U15234 (N_15234,N_14476,N_13316);
and U15235 (N_15235,N_11803,N_13760);
nor U15236 (N_15236,N_14389,N_10520);
or U15237 (N_15237,N_13863,N_12338);
and U15238 (N_15238,N_12730,N_11065);
or U15239 (N_15239,N_12426,N_14318);
and U15240 (N_15240,N_10564,N_13857);
and U15241 (N_15241,N_13298,N_13467);
and U15242 (N_15242,N_12081,N_12832);
and U15243 (N_15243,N_11434,N_13795);
nor U15244 (N_15244,N_10616,N_13067);
nand U15245 (N_15245,N_10913,N_11852);
nor U15246 (N_15246,N_12361,N_13833);
nor U15247 (N_15247,N_14766,N_13801);
nor U15248 (N_15248,N_13818,N_11883);
or U15249 (N_15249,N_13836,N_11263);
nand U15250 (N_15250,N_12994,N_12931);
nor U15251 (N_15251,N_10754,N_11376);
nor U15252 (N_15252,N_13220,N_12803);
nand U15253 (N_15253,N_12679,N_11840);
and U15254 (N_15254,N_11152,N_10098);
and U15255 (N_15255,N_13978,N_13211);
and U15256 (N_15256,N_12146,N_10006);
nor U15257 (N_15257,N_12919,N_13721);
nor U15258 (N_15258,N_14917,N_13550);
nor U15259 (N_15259,N_10319,N_10095);
nor U15260 (N_15260,N_10888,N_14983);
and U15261 (N_15261,N_13860,N_13492);
nor U15262 (N_15262,N_12510,N_11275);
or U15263 (N_15263,N_12190,N_11975);
or U15264 (N_15264,N_13805,N_14456);
and U15265 (N_15265,N_11998,N_14925);
nor U15266 (N_15266,N_14175,N_10847);
and U15267 (N_15267,N_12021,N_12397);
nor U15268 (N_15268,N_10353,N_11721);
and U15269 (N_15269,N_12855,N_11312);
nand U15270 (N_15270,N_11027,N_12004);
or U15271 (N_15271,N_14570,N_10056);
nand U15272 (N_15272,N_11020,N_14512);
nor U15273 (N_15273,N_13612,N_10104);
and U15274 (N_15274,N_14370,N_14837);
nor U15275 (N_15275,N_10638,N_13999);
nor U15276 (N_15276,N_14718,N_11190);
or U15277 (N_15277,N_13218,N_10084);
nand U15278 (N_15278,N_10474,N_10906);
or U15279 (N_15279,N_14188,N_14641);
or U15280 (N_15280,N_10173,N_11227);
or U15281 (N_15281,N_13617,N_14327);
nand U15282 (N_15282,N_13124,N_11217);
or U15283 (N_15283,N_10646,N_12032);
or U15284 (N_15284,N_10551,N_11856);
and U15285 (N_15285,N_10080,N_14279);
or U15286 (N_15286,N_10203,N_11534);
and U15287 (N_15287,N_14477,N_10456);
nor U15288 (N_15288,N_12777,N_11106);
nor U15289 (N_15289,N_13942,N_14036);
nand U15290 (N_15290,N_11149,N_11999);
nor U15291 (N_15291,N_12252,N_14042);
and U15292 (N_15292,N_10929,N_13628);
and U15293 (N_15293,N_12851,N_10295);
nor U15294 (N_15294,N_11705,N_12810);
nor U15295 (N_15295,N_11910,N_10012);
and U15296 (N_15296,N_12837,N_10665);
and U15297 (N_15297,N_13587,N_14469);
nand U15298 (N_15298,N_14942,N_10337);
nand U15299 (N_15299,N_10784,N_12050);
or U15300 (N_15300,N_10066,N_11514);
or U15301 (N_15301,N_12115,N_14866);
and U15302 (N_15302,N_13768,N_12828);
nor U15303 (N_15303,N_13880,N_14184);
and U15304 (N_15304,N_14162,N_12056);
and U15305 (N_15305,N_10981,N_14407);
or U15306 (N_15306,N_11802,N_13735);
and U15307 (N_15307,N_12491,N_10773);
and U15308 (N_15308,N_11073,N_10726);
nand U15309 (N_15309,N_13115,N_10586);
nand U15310 (N_15310,N_13105,N_14333);
nand U15311 (N_15311,N_11936,N_11432);
or U15312 (N_15312,N_11188,N_12482);
and U15313 (N_15313,N_12650,N_11382);
or U15314 (N_15314,N_13227,N_10887);
or U15315 (N_15315,N_13350,N_11258);
and U15316 (N_15316,N_13726,N_14261);
and U15317 (N_15317,N_10127,N_13078);
or U15318 (N_15318,N_12610,N_10516);
or U15319 (N_15319,N_14131,N_13622);
or U15320 (N_15320,N_14760,N_13424);
nand U15321 (N_15321,N_11768,N_12893);
nor U15322 (N_15322,N_12736,N_12935);
or U15323 (N_15323,N_12808,N_12366);
nand U15324 (N_15324,N_10713,N_12451);
and U15325 (N_15325,N_14877,N_10628);
nand U15326 (N_15326,N_10277,N_14128);
nand U15327 (N_15327,N_13773,N_10406);
or U15328 (N_15328,N_11101,N_14142);
nor U15329 (N_15329,N_12231,N_12185);
and U15330 (N_15330,N_12597,N_14002);
or U15331 (N_15331,N_12966,N_13690);
nor U15332 (N_15332,N_11193,N_14071);
or U15333 (N_15333,N_13042,N_12895);
nor U15334 (N_15334,N_10034,N_11753);
nor U15335 (N_15335,N_11718,N_11220);
nand U15336 (N_15336,N_11349,N_14217);
and U15337 (N_15337,N_12821,N_10251);
nand U15338 (N_15338,N_10468,N_12771);
xor U15339 (N_15339,N_13798,N_14296);
nor U15340 (N_15340,N_11371,N_12907);
nand U15341 (N_15341,N_14412,N_10389);
or U15342 (N_15342,N_13594,N_14839);
or U15343 (N_15343,N_11482,N_14830);
nand U15344 (N_15344,N_14945,N_11372);
and U15345 (N_15345,N_10178,N_11052);
nand U15346 (N_15346,N_10928,N_10766);
or U15347 (N_15347,N_11898,N_11129);
nand U15348 (N_15348,N_13537,N_13184);
and U15349 (N_15349,N_10831,N_10689);
or U15350 (N_15350,N_12681,N_13347);
nand U15351 (N_15351,N_14629,N_13473);
nor U15352 (N_15352,N_13406,N_13210);
nor U15353 (N_15353,N_14549,N_14522);
nand U15354 (N_15354,N_10804,N_12546);
or U15355 (N_15355,N_11357,N_11938);
nand U15356 (N_15356,N_10889,N_11623);
nor U15357 (N_15357,N_12719,N_13987);
and U15358 (N_15358,N_13087,N_12398);
and U15359 (N_15359,N_14434,N_11497);
and U15360 (N_15360,N_10092,N_11502);
nand U15361 (N_15361,N_13378,N_14439);
nand U15362 (N_15362,N_11568,N_12200);
nand U15363 (N_15363,N_12950,N_13712);
nor U15364 (N_15364,N_13711,N_13653);
and U15365 (N_15365,N_12233,N_11704);
nand U15366 (N_15366,N_11487,N_12220);
nand U15367 (N_15367,N_10699,N_12724);
or U15368 (N_15368,N_10645,N_12991);
and U15369 (N_15369,N_11561,N_12813);
and U15370 (N_15370,N_10673,N_13856);
nor U15371 (N_15371,N_12559,N_13514);
and U15372 (N_15372,N_14362,N_13970);
nor U15373 (N_15373,N_14978,N_14194);
or U15374 (N_15374,N_14930,N_13146);
nor U15375 (N_15375,N_10859,N_12634);
nor U15376 (N_15376,N_14387,N_12467);
nor U15377 (N_15377,N_10404,N_13648);
or U15378 (N_15378,N_11875,N_13169);
and U15379 (N_15379,N_14530,N_10058);
or U15380 (N_15380,N_11836,N_11624);
and U15381 (N_15381,N_13552,N_13752);
or U15382 (N_15382,N_11176,N_13219);
or U15383 (N_15383,N_12944,N_11331);
and U15384 (N_15384,N_12170,N_11401);
or U15385 (N_15385,N_10772,N_14702);
or U15386 (N_15386,N_14801,N_11743);
nor U15387 (N_15387,N_10512,N_14572);
or U15388 (N_15388,N_10082,N_13083);
nand U15389 (N_15389,N_10522,N_10150);
nor U15390 (N_15390,N_10008,N_14529);
xor U15391 (N_15391,N_13827,N_11711);
nor U15392 (N_15392,N_10932,N_12531);
nor U15393 (N_15393,N_13638,N_12509);
and U15394 (N_15394,N_14986,N_12225);
nor U15395 (N_15395,N_10562,N_10968);
and U15396 (N_15396,N_10838,N_12296);
and U15397 (N_15397,N_14310,N_13474);
nor U15398 (N_15398,N_14501,N_11831);
or U15399 (N_15399,N_14223,N_11925);
or U15400 (N_15400,N_13415,N_10970);
nand U15401 (N_15401,N_10307,N_12374);
nand U15402 (N_15402,N_12477,N_11285);
or U15403 (N_15403,N_13939,N_10286);
nor U15404 (N_15404,N_11722,N_14332);
nor U15405 (N_15405,N_13767,N_13040);
or U15406 (N_15406,N_12794,N_12762);
nand U15407 (N_15407,N_11557,N_10757);
nand U15408 (N_15408,N_14912,N_13174);
nand U15409 (N_15409,N_13570,N_11063);
nor U15410 (N_15410,N_10204,N_13092);
or U15411 (N_15411,N_13504,N_10191);
and U15412 (N_15412,N_14622,N_14547);
nor U15413 (N_15413,N_13873,N_13841);
nand U15414 (N_15414,N_14770,N_14396);
or U15415 (N_15415,N_14436,N_13329);
nand U15416 (N_15416,N_14426,N_12949);
or U15417 (N_15417,N_10853,N_13023);
or U15418 (N_15418,N_10244,N_12702);
and U15419 (N_15419,N_12697,N_13919);
nor U15420 (N_15420,N_10015,N_10707);
nor U15421 (N_15421,N_12447,N_10427);
and U15422 (N_15422,N_12793,N_11523);
nand U15423 (N_15423,N_10903,N_12078);
xor U15424 (N_15424,N_10803,N_13104);
and U15425 (N_15425,N_14534,N_13911);
nor U15426 (N_15426,N_13206,N_11784);
or U15427 (N_15427,N_12104,N_14047);
or U15428 (N_15428,N_13591,N_12377);
and U15429 (N_15429,N_11511,N_13363);
nor U15430 (N_15430,N_14209,N_14252);
nand U15431 (N_15431,N_14233,N_13756);
nor U15432 (N_15432,N_14807,N_14102);
and U15433 (N_15433,N_12957,N_13876);
and U15434 (N_15434,N_12446,N_10550);
nand U15435 (N_15435,N_14575,N_14926);
and U15436 (N_15436,N_13213,N_14857);
and U15437 (N_15437,N_13465,N_12300);
nor U15438 (N_15438,N_12782,N_10019);
nand U15439 (N_15439,N_11549,N_14574);
nand U15440 (N_15440,N_10769,N_14793);
and U15441 (N_15441,N_12779,N_14580);
nor U15442 (N_15442,N_13671,N_11254);
nand U15443 (N_15443,N_10700,N_11178);
and U15444 (N_15444,N_13694,N_11140);
and U15445 (N_15445,N_10722,N_10298);
and U15446 (N_15446,N_10635,N_11665);
nand U15447 (N_15447,N_14847,N_13740);
or U15448 (N_15448,N_14894,N_13233);
and U15449 (N_15449,N_13668,N_14638);
and U15450 (N_15450,N_12569,N_10305);
or U15451 (N_15451,N_11047,N_11413);
and U15452 (N_15452,N_12852,N_12207);
nor U15453 (N_15453,N_10129,N_13607);
nor U15454 (N_15454,N_14784,N_12859);
and U15455 (N_15455,N_13758,N_11130);
and U15456 (N_15456,N_12294,N_13743);
or U15457 (N_15457,N_11683,N_13557);
nor U15458 (N_15458,N_11629,N_13024);
or U15459 (N_15459,N_10324,N_11653);
nor U15460 (N_15460,N_11844,N_13374);
nor U15461 (N_15461,N_13292,N_14902);
nor U15462 (N_15462,N_14554,N_10949);
or U15463 (N_15463,N_12507,N_10814);
and U15464 (N_15464,N_11741,N_11636);
nor U15465 (N_15465,N_14745,N_12689);
and U15466 (N_15466,N_14306,N_11239);
nor U15467 (N_15467,N_10827,N_10882);
nor U15468 (N_15468,N_12661,N_14809);
or U15469 (N_15469,N_13534,N_12879);
nand U15470 (N_15470,N_12838,N_10010);
or U15471 (N_15471,N_14132,N_13348);
or U15472 (N_15472,N_10555,N_12834);
nand U15473 (N_15473,N_14300,N_12947);
nor U15474 (N_15474,N_12210,N_12116);
and U15475 (N_15475,N_12923,N_11111);
and U15476 (N_15476,N_10280,N_11295);
or U15477 (N_15477,N_12926,N_10566);
nor U15478 (N_15478,N_10631,N_10320);
nor U15479 (N_15479,N_13021,N_10402);
and U15480 (N_15480,N_11086,N_11300);
and U15481 (N_15481,N_11191,N_12809);
nor U15482 (N_15482,N_14557,N_12778);
and U15483 (N_15483,N_13886,N_14253);
and U15484 (N_15484,N_11137,N_12048);
and U15485 (N_15485,N_13392,N_13071);
or U15486 (N_15486,N_12692,N_14259);
and U15487 (N_15487,N_11590,N_14832);
and U15488 (N_15488,N_10538,N_11670);
and U15489 (N_15489,N_11344,N_13187);
nor U15490 (N_15490,N_10500,N_13012);
nor U15491 (N_15491,N_14686,N_11105);
or U15492 (N_15492,N_13490,N_11778);
or U15493 (N_15493,N_12040,N_11642);
and U15494 (N_15494,N_14970,N_10274);
nand U15495 (N_15495,N_12968,N_11728);
or U15496 (N_15496,N_14670,N_14060);
or U15497 (N_15497,N_13178,N_10687);
or U15498 (N_15498,N_12652,N_13807);
or U15499 (N_15499,N_12647,N_14249);
and U15500 (N_15500,N_12399,N_12664);
or U15501 (N_15501,N_11977,N_11001);
nor U15502 (N_15502,N_10107,N_12636);
or U15503 (N_15503,N_10164,N_12174);
nor U15504 (N_15504,N_12277,N_10143);
nand U15505 (N_15505,N_14422,N_11333);
or U15506 (N_15506,N_14783,N_13643);
nand U15507 (N_15507,N_13749,N_12083);
or U15508 (N_15508,N_13908,N_10458);
nor U15509 (N_15509,N_10065,N_11895);
and U15510 (N_15510,N_10959,N_10246);
nand U15511 (N_15511,N_12928,N_12089);
and U15512 (N_15512,N_11060,N_10709);
nand U15513 (N_15513,N_14180,N_12264);
nor U15514 (N_15514,N_14787,N_14424);
and U15515 (N_15515,N_11143,N_11405);
and U15516 (N_15516,N_10917,N_11318);
nand U15517 (N_15517,N_11608,N_10193);
or U15518 (N_15518,N_11603,N_11392);
or U15519 (N_15519,N_11112,N_11877);
or U15520 (N_15520,N_12801,N_10539);
or U15521 (N_15521,N_13858,N_12537);
nand U15522 (N_15522,N_12240,N_11745);
nand U15523 (N_15523,N_13099,N_13022);
nor U15524 (N_15524,N_10325,N_12726);
nand U15525 (N_15525,N_12184,N_14376);
nand U15526 (N_15526,N_13152,N_13242);
or U15527 (N_15527,N_14255,N_11099);
and U15528 (N_15528,N_11174,N_10333);
and U15529 (N_15529,N_10488,N_10209);
nor U15530 (N_15530,N_11041,N_10424);
nand U15531 (N_15531,N_10643,N_10948);
and U15532 (N_15532,N_13295,N_14357);
or U15533 (N_15533,N_11369,N_13739);
nand U15534 (N_15534,N_13461,N_11596);
nor U15535 (N_15535,N_10142,N_12118);
nor U15536 (N_15536,N_13102,N_14519);
and U15537 (N_15537,N_14910,N_14602);
or U15538 (N_15538,N_12543,N_12437);
or U15539 (N_15539,N_10229,N_13884);
nor U15540 (N_15540,N_13372,N_10275);
nand U15541 (N_15541,N_11573,N_13006);
and U15542 (N_15542,N_13770,N_10636);
and U15543 (N_15543,N_11702,N_11367);
and U15544 (N_15544,N_12253,N_12131);
or U15545 (N_15545,N_11839,N_10338);
nand U15546 (N_15546,N_12459,N_14435);
and U15547 (N_15547,N_13766,N_12978);
nand U15548 (N_15548,N_14543,N_14150);
nor U15549 (N_15549,N_12554,N_14587);
and U15550 (N_15550,N_10820,N_11576);
nand U15551 (N_15551,N_13747,N_11915);
nor U15552 (N_15552,N_11921,N_13980);
nor U15553 (N_15553,N_11564,N_13626);
and U15554 (N_15554,N_13388,N_10523);
nor U15555 (N_15555,N_12958,N_12783);
nand U15556 (N_15556,N_11067,N_12385);
nand U15557 (N_15557,N_13179,N_13535);
nor U15558 (N_15558,N_11183,N_12255);
or U15559 (N_15559,N_11627,N_14315);
and U15560 (N_15560,N_14448,N_11474);
and U15561 (N_15561,N_12266,N_12498);
nand U15562 (N_15562,N_10345,N_11657);
nor U15563 (N_15563,N_12316,N_14179);
and U15564 (N_15564,N_10388,N_11565);
or U15565 (N_15565,N_14463,N_12604);
nand U15566 (N_15566,N_13068,N_14533);
nand U15567 (N_15567,N_12229,N_13647);
and U15568 (N_15568,N_14550,N_10235);
or U15569 (N_15569,N_10116,N_12909);
nand U15570 (N_15570,N_14692,N_13501);
nor U15571 (N_15571,N_13396,N_10124);
nor U15572 (N_15572,N_14385,N_12572);
nand U15573 (N_15573,N_11460,N_12053);
and U15574 (N_15574,N_11085,N_13427);
or U15575 (N_15575,N_10659,N_10167);
and U15576 (N_15576,N_10282,N_14069);
or U15577 (N_15577,N_14540,N_14663);
nor U15578 (N_15578,N_14311,N_10556);
or U15579 (N_15579,N_12221,N_10750);
or U15580 (N_15580,N_12637,N_12698);
and U15581 (N_15581,N_11846,N_11771);
nand U15582 (N_15582,N_14779,N_10690);
and U15583 (N_15583,N_11185,N_10130);
nand U15584 (N_15584,N_10405,N_13903);
nand U15585 (N_15585,N_13586,N_11816);
or U15586 (N_15586,N_11054,N_14568);
and U15587 (N_15587,N_14730,N_10187);
or U15588 (N_15588,N_13536,N_10444);
and U15589 (N_15589,N_12001,N_10619);
or U15590 (N_15590,N_10180,N_14729);
and U15591 (N_15591,N_14941,N_10666);
nand U15592 (N_15592,N_13581,N_10608);
xnor U15593 (N_15593,N_13569,N_14590);
nor U15594 (N_15594,N_12512,N_14099);
and U15595 (N_15595,N_12905,N_10945);
or U15596 (N_15596,N_13069,N_13777);
nand U15597 (N_15597,N_11954,N_14317);
and U15598 (N_15598,N_12561,N_13150);
and U15599 (N_15599,N_10453,N_14654);
and U15600 (N_15600,N_12257,N_12387);
or U15601 (N_15601,N_14603,N_14747);
nand U15602 (N_15602,N_14596,N_10536);
and U15603 (N_15603,N_11594,N_13127);
nand U15604 (N_15604,N_11062,N_12671);
nor U15605 (N_15605,N_14367,N_11411);
or U15606 (N_15606,N_14892,N_10367);
and U15607 (N_15607,N_13769,N_10807);
or U15608 (N_15608,N_14571,N_11973);
and U15609 (N_15609,N_10826,N_12100);
and U15610 (N_15610,N_12894,N_14058);
or U15611 (N_15611,N_13598,N_10860);
or U15612 (N_15612,N_14662,N_13757);
and U15613 (N_15613,N_11232,N_11484);
nor U15614 (N_15614,N_12161,N_10669);
or U15615 (N_15615,N_13008,N_10873);
nand U15616 (N_15616,N_14478,N_13291);
nor U15617 (N_15617,N_12324,N_10966);
or U15618 (N_15618,N_10946,N_11770);
nor U15619 (N_15619,N_11772,N_11374);
and U15620 (N_15620,N_13825,N_13226);
nand U15621 (N_15621,N_14371,N_11076);
and U15622 (N_15622,N_13470,N_13192);
nor U15623 (N_15623,N_13551,N_12609);
nor U15624 (N_15624,N_12840,N_14085);
or U15625 (N_15625,N_13682,N_13385);
and U15626 (N_15626,N_10285,N_10368);
nor U15627 (N_15627,N_11951,N_11033);
and U15628 (N_15628,N_14467,N_11701);
nor U15629 (N_15629,N_10428,N_13859);
or U15630 (N_15630,N_12270,N_14174);
or U15631 (N_15631,N_12780,N_11031);
nor U15632 (N_15632,N_14763,N_11266);
nand U15633 (N_15633,N_13719,N_14022);
and U15634 (N_15634,N_14581,N_10262);
and U15635 (N_15635,N_12074,N_11466);
and U15636 (N_15636,N_13039,N_13639);
nand U15637 (N_15637,N_11091,N_10017);
nor U15638 (N_15638,N_13923,N_12731);
nand U15639 (N_15639,N_11994,N_14086);
or U15640 (N_15640,N_13110,N_13351);
nand U15641 (N_15641,N_10489,N_10049);
nand U15642 (N_15642,N_13894,N_11760);
or U15643 (N_15643,N_14377,N_14932);
nand U15644 (N_15644,N_13964,N_14987);
and U15645 (N_15645,N_13799,N_10618);
and U15646 (N_15646,N_11519,N_11407);
and U15647 (N_15647,N_13936,N_13602);
and U15648 (N_15648,N_12917,N_10501);
nor U15649 (N_15649,N_10222,N_14145);
or U15650 (N_15650,N_13051,N_13614);
nor U15651 (N_15651,N_13867,N_11698);
or U15652 (N_15652,N_12427,N_10448);
nand U15653 (N_15653,N_11648,N_11610);
nor U15654 (N_15654,N_14421,N_10485);
nor U15655 (N_15655,N_10747,N_14964);
nand U15656 (N_15656,N_11212,N_11505);
nor U15657 (N_15657,N_14073,N_10225);
nand U15658 (N_15658,N_13986,N_11643);
and U15659 (N_15659,N_11833,N_13592);
or U15660 (N_15660,N_10477,N_12583);
or U15661 (N_15661,N_14417,N_13754);
or U15662 (N_15662,N_10934,N_14247);
nand U15663 (N_15663,N_12036,N_14754);
or U15664 (N_15664,N_13052,N_13486);
and U15665 (N_15665,N_13118,N_11780);
and U15666 (N_15666,N_12910,N_14751);
nor U15667 (N_15667,N_12193,N_14454);
nor U15668 (N_15668,N_14307,N_10971);
or U15669 (N_15669,N_13208,N_13910);
nor U15670 (N_15670,N_10386,N_10937);
and U15671 (N_15671,N_10196,N_11307);
or U15672 (N_15672,N_14944,N_11671);
xnor U15673 (N_15673,N_12902,N_10779);
nor U15674 (N_15674,N_13959,N_14748);
and U15675 (N_15675,N_12723,N_11465);
nand U15676 (N_15676,N_11738,N_12886);
and U15677 (N_15677,N_11399,N_10809);
or U15678 (N_15678,N_10002,N_14445);
nor U15679 (N_15679,N_13111,N_14739);
nor U15680 (N_15680,N_12343,N_12878);
and U15681 (N_15681,N_14301,N_11024);
and U15682 (N_15682,N_13173,N_10125);
nand U15683 (N_15683,N_13829,N_10241);
nor U15684 (N_15684,N_10661,N_13354);
nand U15685 (N_15685,N_13877,N_10261);
or U15686 (N_15686,N_14843,N_13823);
or U15687 (N_15687,N_11245,N_14858);
nor U15688 (N_15688,N_12219,N_12395);
nor U15689 (N_15689,N_14324,N_14186);
and U15690 (N_15690,N_14100,N_12013);
nand U15691 (N_15691,N_10877,N_14045);
or U15692 (N_15692,N_10438,N_11851);
nor U15693 (N_15693,N_12648,N_13846);
nor U15694 (N_15694,N_10451,N_11214);
or U15695 (N_15695,N_10611,N_10001);
nand U15696 (N_15696,N_11423,N_11966);
nor U15697 (N_15697,N_11457,N_11427);
nor U15698 (N_15698,N_12557,N_12429);
or U15699 (N_15699,N_13518,N_13197);
or U15700 (N_15700,N_11635,N_11735);
or U15701 (N_15701,N_13225,N_11456);
or U15702 (N_15702,N_10597,N_13929);
nor U15703 (N_15703,N_10911,N_10061);
and U15704 (N_15704,N_13700,N_14080);
nor U15705 (N_15705,N_11284,N_10716);
or U15706 (N_15706,N_12178,N_11082);
or U15707 (N_15707,N_10393,N_11990);
nor U15708 (N_15708,N_12675,N_12900);
and U15709 (N_15709,N_10863,N_11416);
or U15710 (N_15710,N_14220,N_11620);
nor U15711 (N_15711,N_11663,N_11075);
nand U15712 (N_15712,N_10224,N_14200);
and U15713 (N_15713,N_10007,N_14955);
nor U15714 (N_15714,N_14583,N_13308);
nor U15715 (N_15715,N_14159,N_10219);
nand U15716 (N_15716,N_13004,N_13321);
or U15717 (N_15717,N_14630,N_12712);
and U15718 (N_15718,N_14735,N_13138);
nor U15719 (N_15719,N_11237,N_11522);
xnor U15720 (N_15720,N_11177,N_11552);
nand U15721 (N_15721,N_14569,N_10024);
and U15722 (N_15722,N_14487,N_13510);
and U15723 (N_15723,N_11583,N_10226);
nand U15724 (N_15724,N_14780,N_10793);
nor U15725 (N_15725,N_13993,N_13519);
nor U15726 (N_15726,N_11361,N_10732);
and U15727 (N_15727,N_12739,N_14816);
nand U15728 (N_15728,N_12027,N_10783);
nand U15729 (N_15729,N_13542,N_11788);
nand U15730 (N_15730,N_13853,N_14701);
nand U15731 (N_15731,N_11755,N_12582);
and U15732 (N_15732,N_10158,N_12329);
nor U15733 (N_15733,N_12518,N_11845);
nand U15734 (N_15734,N_14316,N_14715);
and U15735 (N_15735,N_11393,N_11389);
and U15736 (N_15736,N_14664,N_13147);
nand U15737 (N_15737,N_11793,N_13356);
and U15738 (N_15738,N_12595,N_14411);
nand U15739 (N_15739,N_14129,N_10118);
or U15740 (N_15740,N_12314,N_13002);
nand U15741 (N_15741,N_14352,N_13728);
and U15742 (N_15742,N_14378,N_12686);
or U15743 (N_15743,N_12876,N_12987);
and U15744 (N_15744,N_13265,N_10965);
xnor U15745 (N_15745,N_11498,N_13073);
nor U15746 (N_15746,N_10810,N_11941);
or U15747 (N_15747,N_12079,N_10408);
nor U15748 (N_15748,N_10385,N_11893);
and U15749 (N_15749,N_13402,N_14280);
nor U15750 (N_15750,N_12932,N_12352);
nand U15751 (N_15751,N_11834,N_13975);
and U15752 (N_15752,N_13257,N_12344);
or U15753 (N_15753,N_14323,N_10192);
and U15754 (N_15754,N_10712,N_10339);
and U15755 (N_15755,N_10613,N_11297);
nor U15756 (N_15756,N_14795,N_13421);
nand U15757 (N_15757,N_12431,N_12608);
and U15758 (N_15758,N_10370,N_12845);
nand U15759 (N_15759,N_12961,N_10604);
nand U15760 (N_15760,N_13272,N_12842);
nor U15761 (N_15761,N_12218,N_12382);
and U15762 (N_15762,N_10174,N_11323);
or U15763 (N_15763,N_13549,N_10579);
or U15764 (N_15764,N_10227,N_13191);
nor U15765 (N_15765,N_14940,N_12735);
nand U15766 (N_15766,N_13478,N_11283);
nor U15767 (N_15767,N_10134,N_10437);
or U15768 (N_15768,N_13588,N_11094);
and U15769 (N_15769,N_13692,N_14012);
or U15770 (N_15770,N_12244,N_10755);
and U15771 (N_15771,N_10144,N_14732);
or U15772 (N_15772,N_13717,N_11061);
nand U15773 (N_15773,N_10925,N_14799);
or U15774 (N_15774,N_10815,N_10606);
and U15775 (N_15775,N_10413,N_12754);
nor U15776 (N_15776,N_14646,N_11981);
and U15777 (N_15777,N_13450,N_12060);
and U15778 (N_15778,N_14699,N_10759);
and U15779 (N_15779,N_14391,N_14450);
or U15780 (N_15780,N_14048,N_14402);
or U15781 (N_15781,N_12963,N_13307);
and U15782 (N_15782,N_11461,N_12135);
and U15783 (N_15783,N_13512,N_12157);
nor U15784 (N_15784,N_12908,N_12822);
or U15785 (N_15785,N_13744,N_12494);
or U15786 (N_15786,N_14197,N_13207);
or U15787 (N_15787,N_14500,N_11873);
or U15788 (N_15788,N_13352,N_10421);
and U15789 (N_15789,N_12873,N_13834);
or U15790 (N_15790,N_11277,N_13640);
xnor U15791 (N_15791,N_13389,N_14578);
nor U15792 (N_15792,N_12705,N_12490);
or U15793 (N_15793,N_14636,N_12775);
nor U15794 (N_15794,N_13418,N_14895);
or U15795 (N_15795,N_12708,N_14871);
and U15796 (N_15796,N_10390,N_14722);
nand U15797 (N_15797,N_11542,N_10875);
and U15798 (N_15798,N_13967,N_13142);
nand U15799 (N_15799,N_13812,N_14274);
and U15800 (N_15800,N_14666,N_12340);
or U15801 (N_15801,N_12576,N_13391);
nor U15802 (N_15802,N_12843,N_11709);
nand U15803 (N_15803,N_12030,N_10674);
nand U15804 (N_15804,N_14257,N_11726);
and U15805 (N_15805,N_11272,N_14285);
xnor U15806 (N_15806,N_12483,N_11644);
nand U15807 (N_15807,N_13090,N_10239);
and U15808 (N_15808,N_14264,N_11708);
and U15809 (N_15809,N_13930,N_14721);
or U15810 (N_15810,N_13000,N_11509);
or U15811 (N_15811,N_11920,N_13809);
and U15812 (N_15812,N_12520,N_10845);
or U15813 (N_15813,N_13940,N_10464);
and U15814 (N_15814,N_11452,N_10009);
and U15815 (N_15815,N_14291,N_14430);
or U15816 (N_15816,N_13655,N_14913);
or U15817 (N_15817,N_11578,N_14693);
and U15818 (N_15818,N_12599,N_11510);
nor U15819 (N_15819,N_12005,N_13416);
or U15820 (N_15820,N_13074,N_12544);
nand U15821 (N_15821,N_10647,N_12953);
nor U15822 (N_15822,N_11862,N_13380);
nand U15823 (N_15823,N_13362,N_12278);
nor U15824 (N_15824,N_12700,N_13882);
nand U15825 (N_15825,N_12368,N_10584);
or U15826 (N_15826,N_12448,N_12499);
nor U15827 (N_15827,N_14864,N_11619);
nor U15828 (N_15828,N_13585,N_12372);
or U15829 (N_15829,N_12370,N_11861);
and U15830 (N_15830,N_13997,N_12620);
nor U15831 (N_15831,N_13493,N_13865);
nor U15832 (N_15832,N_10655,N_14172);
nor U15833 (N_15833,N_11448,N_11483);
or U15834 (N_15834,N_11209,N_11992);
nand U15835 (N_15835,N_11689,N_14453);
nand U15836 (N_15836,N_14127,N_14988);
nor U15837 (N_15837,N_11540,N_13737);
and U15838 (N_15838,N_14861,N_10982);
nand U15839 (N_15839,N_10837,N_12386);
nand U15840 (N_15840,N_13005,N_10990);
nand U15841 (N_15841,N_11805,N_10470);
or U15842 (N_15842,N_12390,N_13304);
nor U15843 (N_15843,N_14643,N_14959);
nand U15844 (N_15844,N_10288,N_10380);
and U15845 (N_15845,N_13423,N_12102);
and U15846 (N_15846,N_11256,N_14804);
nor U15847 (N_15847,N_14064,N_14789);
and U15848 (N_15848,N_13079,N_13521);
and U15849 (N_15849,N_13377,N_10033);
and U15850 (N_15850,N_12112,N_12922);
nand U15851 (N_15851,N_13709,N_11334);
nor U15852 (N_15852,N_11006,N_11591);
or U15853 (N_15853,N_13144,N_12400);
nor U15854 (N_15854,N_10048,N_11016);
or U15855 (N_15855,N_14828,N_14755);
nand U15856 (N_15856,N_12006,N_14420);
nor U15857 (N_15857,N_14979,N_11166);
and U15858 (N_15858,N_14289,N_12163);
or U15859 (N_15859,N_14239,N_13193);
or U15860 (N_15860,N_12098,N_14438);
or U15861 (N_15861,N_12181,N_12706);
or U15862 (N_15862,N_14812,N_11104);
nand U15863 (N_15863,N_12912,N_11806);
or U15864 (N_15864,N_10364,N_14967);
nor U15865 (N_15865,N_14447,N_11582);
nor U15866 (N_15866,N_11706,N_10715);
or U15867 (N_15867,N_14826,N_13201);
nor U15868 (N_15868,N_14455,N_13893);
and U15869 (N_15869,N_11678,N_10541);
nand U15870 (N_15870,N_12303,N_11373);
nand U15871 (N_15871,N_13489,N_11604);
nand U15872 (N_15872,N_13574,N_10980);
nand U15873 (N_15873,N_12728,N_10311);
and U15874 (N_15874,N_12541,N_11503);
nand U15875 (N_15875,N_12495,N_11661);
nand U15876 (N_15876,N_14005,N_12898);
nand U15877 (N_15877,N_13091,N_11518);
nor U15878 (N_15878,N_12356,N_12789);
and U15879 (N_15879,N_14946,N_14528);
or U15880 (N_15880,N_12464,N_13553);
or U15881 (N_15881,N_13333,N_13874);
nand U15882 (N_15882,N_13875,N_12707);
nor U15883 (N_15883,N_14258,N_14750);
nor U15884 (N_15884,N_14566,N_10194);
or U15885 (N_15885,N_13398,N_11792);
nor U15886 (N_15886,N_11202,N_11731);
nand U15887 (N_15887,N_12194,N_11471);
nor U15888 (N_15888,N_12301,N_14535);
or U15889 (N_15889,N_10973,N_10670);
nand U15890 (N_15890,N_14025,N_11733);
and U15891 (N_15891,N_13122,N_10540);
and U15892 (N_15892,N_12619,N_14562);
nor U15893 (N_15893,N_12293,N_10938);
or U15894 (N_15894,N_13417,N_14845);
nand U15895 (N_15895,N_10575,N_11662);
nor U15896 (N_15896,N_12085,N_10315);
and U15897 (N_15897,N_11077,N_13185);
nor U15898 (N_15898,N_14711,N_10183);
nand U15899 (N_15899,N_12197,N_10480);
nand U15900 (N_15900,N_14918,N_13063);
nand U15901 (N_15901,N_10133,N_13963);
nor U15902 (N_15902,N_12147,N_10697);
nor U15903 (N_15903,N_14384,N_11435);
or U15904 (N_15904,N_14495,N_11495);
nor U15905 (N_15905,N_11136,N_13160);
nand U15906 (N_15906,N_10498,N_13228);
and U15907 (N_15907,N_13725,N_14177);
nor U15908 (N_15908,N_14337,N_10179);
nor U15909 (N_15909,N_14449,N_10554);
and U15910 (N_15910,N_13382,N_13072);
nor U15911 (N_15911,N_12094,N_11588);
nand U15912 (N_15912,N_11181,N_13706);
nor U15913 (N_15913,N_12547,N_13180);
or U15914 (N_15914,N_11625,N_10721);
nand U15915 (N_15915,N_10858,N_11515);
or U15916 (N_15916,N_13681,N_12035);
nor U15917 (N_15917,N_11221,N_13868);
and U15918 (N_15918,N_11231,N_11400);
nand U15919 (N_15919,N_10260,N_10459);
nor U15920 (N_15920,N_10073,N_13727);
xnor U15921 (N_15921,N_14262,N_12755);
or U15922 (N_15922,N_14304,N_14645);
and U15923 (N_15923,N_13786,N_14458);
nand U15924 (N_15924,N_13311,N_14680);
and U15925 (N_15925,N_13541,N_13481);
or U15926 (N_15926,N_13495,N_14542);
or U15927 (N_15927,N_12402,N_14124);
and U15928 (N_15928,N_13053,N_10985);
nand U15929 (N_15929,N_14633,N_12918);
nor U15930 (N_15930,N_10880,N_13907);
and U15931 (N_15931,N_12884,N_14632);
and U15932 (N_15932,N_14981,N_10933);
nor U15933 (N_15933,N_12575,N_10202);
or U15934 (N_15934,N_13195,N_14786);
or U15935 (N_15935,N_12198,N_14373);
nor U15936 (N_15936,N_12761,N_14433);
nor U15937 (N_15937,N_12176,N_11713);
and U15938 (N_15938,N_10300,N_12150);
nand U15939 (N_15939,N_10184,N_13477);
and U15940 (N_15940,N_13630,N_12424);
or U15941 (N_15941,N_14695,N_11783);
nand U15942 (N_15942,N_13775,N_10278);
nor U15943 (N_15943,N_12924,N_10467);
nand U15944 (N_15944,N_14010,N_13520);
or U15945 (N_15945,N_12757,N_13778);
nand U15946 (N_15946,N_11004,N_10781);
nor U15947 (N_15947,N_11090,N_14284);
and U15948 (N_15948,N_12214,N_11303);
nor U15949 (N_15949,N_14404,N_14138);
and U15950 (N_15950,N_14742,N_11913);
or U15951 (N_15951,N_11468,N_14427);
nor U15952 (N_15952,N_13973,N_12921);
and U15953 (N_15953,N_11028,N_12049);
or U15954 (N_15954,N_13290,N_11964);
nand U15955 (N_15955,N_12388,N_11097);
nor U15956 (N_15956,N_11180,N_13360);
nand U15957 (N_15957,N_10535,N_10657);
or U15958 (N_15958,N_12750,N_10366);
and U15959 (N_15959,N_11649,N_12470);
or U15960 (N_15960,N_11010,N_13263);
and U15961 (N_15961,N_10738,N_12581);
nor U15962 (N_15962,N_13158,N_10172);
or U15963 (N_15963,N_10237,N_14712);
nor U15964 (N_15964,N_11881,N_13826);
or U15965 (N_15965,N_14416,N_10443);
or U15966 (N_15966,N_13010,N_10767);
nand U15967 (N_15967,N_13468,N_12945);
and U15968 (N_15968,N_11184,N_14260);
or U15969 (N_15969,N_12863,N_14153);
or U15970 (N_15970,N_14250,N_11622);
and U15971 (N_15971,N_11598,N_14440);
or U15972 (N_15972,N_13163,N_10147);
nor U15973 (N_15973,N_11479,N_13204);
or U15974 (N_15974,N_13790,N_12442);
and U15975 (N_15975,N_10198,N_13358);
or U15976 (N_15976,N_12882,N_12763);
or U15977 (N_15977,N_14195,N_13500);
nor U15978 (N_15978,N_12419,N_10974);
and U15979 (N_15979,N_10400,N_13476);
nor U15980 (N_15980,N_12109,N_11886);
nand U15981 (N_15981,N_12187,N_13306);
nor U15982 (N_15982,N_13436,N_14952);
nand U15983 (N_15983,N_10035,N_11824);
nand U15984 (N_15984,N_12320,N_13429);
or U15985 (N_15985,N_14312,N_11695);
and U15986 (N_15986,N_11988,N_10951);
nor U15987 (N_15987,N_10620,N_12916);
nor U15988 (N_15988,N_11421,N_10258);
nor U15989 (N_15989,N_14011,N_10904);
or U15990 (N_15990,N_13043,N_11128);
or U15991 (N_15991,N_11198,N_10919);
and U15992 (N_15992,N_10330,N_14517);
nand U15993 (N_15993,N_10161,N_12025);
or U15994 (N_15994,N_12261,N_10703);
or U15995 (N_15995,N_12202,N_10940);
and U15996 (N_15996,N_12939,N_12633);
and U15997 (N_15997,N_13296,N_11789);
or U15998 (N_15998,N_14119,N_11949);
or U15999 (N_15999,N_13892,N_11252);
and U16000 (N_16000,N_10455,N_14224);
nand U16001 (N_16001,N_13540,N_12524);
nand U16002 (N_16002,N_13475,N_12827);
and U16003 (N_16003,N_12029,N_14769);
nand U16004 (N_16004,N_13484,N_13422);
nand U16005 (N_16005,N_10587,N_11756);
nand U16006 (N_16006,N_11676,N_12841);
nor U16007 (N_16007,N_10250,N_12805);
or U16008 (N_16008,N_10296,N_11259);
or U16009 (N_16009,N_12445,N_10374);
or U16010 (N_16010,N_13414,N_11310);
nor U16011 (N_16011,N_13029,N_13176);
and U16012 (N_16012,N_10004,N_11486);
nand U16013 (N_16013,N_10292,N_13962);
or U16014 (N_16014,N_10216,N_10740);
and U16015 (N_16015,N_10775,N_10120);
xnor U16016 (N_16016,N_13948,N_13912);
and U16017 (N_16017,N_12139,N_13531);
or U16018 (N_16018,N_10491,N_11775);
nand U16019 (N_16019,N_11761,N_12096);
nand U16020 (N_16020,N_10508,N_12137);
and U16021 (N_16021,N_10420,N_14218);
nand U16022 (N_16022,N_11684,N_12786);
nand U16023 (N_16023,N_12693,N_14813);
and U16024 (N_16024,N_12438,N_10346);
nor U16025 (N_16025,N_14479,N_14901);
and U16026 (N_16026,N_13273,N_10927);
nand U16027 (N_16027,N_10119,N_10930);
and U16028 (N_16028,N_12996,N_11462);
and U16029 (N_16029,N_11240,N_12549);
and U16030 (N_16030,N_11517,N_10855);
nor U16031 (N_16031,N_11821,N_12653);
and U16032 (N_16032,N_14846,N_10394);
nand U16033 (N_16033,N_10276,N_14425);
or U16034 (N_16034,N_10502,N_12556);
nand U16035 (N_16035,N_10270,N_14393);
nor U16036 (N_16036,N_14505,N_10695);
and U16037 (N_16037,N_12205,N_10774);
nand U16038 (N_16038,N_11338,N_13633);
or U16039 (N_16039,N_10506,N_13697);
and U16040 (N_16040,N_14146,N_14198);
or U16041 (N_16041,N_14607,N_13960);
or U16042 (N_16042,N_14170,N_14842);
nor U16043 (N_16043,N_10044,N_14382);
nor U16044 (N_16044,N_11876,N_11356);
nor U16045 (N_16045,N_14811,N_12331);
nor U16046 (N_16046,N_12322,N_12363);
and U16047 (N_16047,N_14221,N_14056);
and U16048 (N_16048,N_14634,N_12747);
or U16049 (N_16049,N_13036,N_10289);
nand U16050 (N_16050,N_10899,N_12247);
nand U16051 (N_16051,N_13281,N_11847);
or U16052 (N_16052,N_11135,N_14466);
nor U16053 (N_16053,N_14392,N_11358);
and U16054 (N_16054,N_14889,N_10864);
nand U16055 (N_16055,N_11354,N_14791);
or U16056 (N_16056,N_11289,N_11243);
nand U16057 (N_16057,N_12230,N_12621);
and U16058 (N_16058,N_12660,N_12038);
nand U16059 (N_16059,N_11420,N_11971);
xor U16060 (N_16060,N_12717,N_12975);
nand U16061 (N_16061,N_14428,N_12971);
xor U16062 (N_16062,N_11903,N_14321);
nor U16063 (N_16063,N_12142,N_14269);
nand U16064 (N_16064,N_11383,N_13554);
and U16065 (N_16065,N_13149,N_10291);
nor U16066 (N_16066,N_12920,N_12829);
nand U16067 (N_16067,N_13261,N_10504);
nor U16068 (N_16068,N_13248,N_14091);
nand U16069 (N_16069,N_11163,N_11957);
nand U16070 (N_16070,N_12555,N_10081);
nand U16071 (N_16071,N_13969,N_13691);
nand U16072 (N_16072,N_13820,N_12328);
nor U16073 (N_16073,N_11924,N_12392);
and U16074 (N_16074,N_13762,N_10801);
and U16075 (N_16075,N_10908,N_12486);
nand U16076 (N_16076,N_12274,N_14511);
and U16077 (N_16077,N_12422,N_14388);
nor U16078 (N_16078,N_11021,N_13080);
or U16079 (N_16079,N_13751,N_13763);
nand U16080 (N_16080,N_13299,N_11907);
or U16081 (N_16081,N_11342,N_13089);
and U16082 (N_16082,N_12348,N_13983);
and U16083 (N_16083,N_14594,N_10031);
or U16084 (N_16084,N_11032,N_11817);
nor U16085 (N_16085,N_11403,N_12330);
nor U16086 (N_16086,N_13575,N_14203);
or U16087 (N_16087,N_10415,N_14489);
nand U16088 (N_16088,N_11906,N_11044);
or U16089 (N_16089,N_10694,N_11424);
nand U16090 (N_16090,N_10155,N_14672);
xnor U16091 (N_16091,N_14898,N_11370);
nor U16092 (N_16092,N_10943,N_13399);
or U16093 (N_16093,N_13047,N_12063);
nor U16094 (N_16094,N_12373,N_14954);
and U16095 (N_16095,N_14887,N_10921);
or U16096 (N_16096,N_14230,N_13196);
and U16097 (N_16097,N_13677,N_11690);
nor U16098 (N_16098,N_11659,N_11088);
nor U16099 (N_16099,N_10914,N_14481);
or U16100 (N_16100,N_12980,N_12563);
and U16101 (N_16101,N_13657,N_12481);
or U16102 (N_16102,N_14508,N_12073);
nor U16103 (N_16103,N_14237,N_11250);
nor U16104 (N_16104,N_11560,N_14778);
nand U16105 (N_16105,N_13990,N_13025);
and U16106 (N_16106,N_13580,N_11720);
or U16107 (N_16107,N_11688,N_13020);
or U16108 (N_16108,N_12849,N_13485);
nor U16109 (N_16109,N_12848,N_13157);
nor U16110 (N_16110,N_13610,N_10795);
or U16111 (N_16111,N_10796,N_14116);
and U16112 (N_16112,N_14725,N_13278);
nand U16113 (N_16113,N_11562,N_12839);
nand U16114 (N_16114,N_14911,N_12466);
nand U16115 (N_16115,N_10446,N_12105);
xnor U16116 (N_16116,N_12463,N_10866);
or U16117 (N_16117,N_12456,N_11262);
nor U16118 (N_16118,N_10240,N_13027);
nand U16119 (N_16119,N_12797,N_10798);
and U16120 (N_16120,N_14818,N_10590);
or U16121 (N_16121,N_14103,N_12280);
nand U16122 (N_16122,N_14728,N_14827);
or U16123 (N_16123,N_11896,N_14176);
nor U16124 (N_16124,N_14169,N_12820);
and U16125 (N_16125,N_13645,N_13215);
nor U16126 (N_16126,N_14437,N_13724);
nand U16127 (N_16127,N_14620,N_13267);
nor U16128 (N_16128,N_12488,N_12072);
nand U16129 (N_16129,N_13530,N_11443);
nand U16130 (N_16130,N_11394,N_10548);
and U16131 (N_16131,N_10764,N_12458);
and U16132 (N_16132,N_13277,N_14849);
nand U16133 (N_16133,N_13403,N_13560);
or U16134 (N_16134,N_11829,N_13817);
nor U16135 (N_16135,N_13946,N_10874);
nor U16136 (N_16136,N_10533,N_14740);
and U16137 (N_16137,N_12265,N_12493);
nor U16138 (N_16138,N_13764,N_11007);
nor U16139 (N_16139,N_12925,N_13386);
and U16140 (N_16140,N_14363,N_14349);
xnor U16141 (N_16141,N_12242,N_14158);
nor U16142 (N_16142,N_13370,N_14870);
or U16143 (N_16143,N_11440,N_13720);
nor U16144 (N_16144,N_11172,N_11107);
nor U16145 (N_16145,N_12678,N_10829);
nor U16146 (N_16146,N_10872,N_14611);
nand U16147 (N_16147,N_10221,N_10672);
nor U16148 (N_16148,N_10060,N_11011);
nand U16149 (N_16149,N_12129,N_14521);
and U16150 (N_16150,N_11124,N_12024);
and U16151 (N_16151,N_14656,N_10211);
nand U16152 (N_16152,N_12312,N_10857);
or U16153 (N_16153,N_11808,N_11759);
nor U16154 (N_16154,N_13181,N_13096);
nor U16155 (N_16155,N_13596,N_13529);
and U16156 (N_16156,N_11734,N_10808);
nand U16157 (N_16157,N_12680,N_12003);
nor U16158 (N_16158,N_14815,N_13202);
and U16159 (N_16159,N_12565,N_13933);
nor U16160 (N_16160,N_12788,N_11908);
nand U16161 (N_16161,N_13685,N_14295);
or U16162 (N_16162,N_13784,N_14070);
and U16163 (N_16163,N_13636,N_13446);
nor U16164 (N_16164,N_11811,N_13018);
and U16165 (N_16165,N_14334,N_12956);
nand U16166 (N_16166,N_10515,N_10668);
nor U16167 (N_16167,N_14733,N_11566);
nor U16168 (N_16168,N_13106,N_10436);
or U16169 (N_16169,N_11631,N_12566);
or U16170 (N_16170,N_13611,N_10813);
nand U16171 (N_16171,N_14256,N_13664);
or U16172 (N_16172,N_11264,N_10947);
or U16173 (N_16173,N_11319,N_11723);
nand U16174 (N_16174,N_13434,N_10281);
nor U16175 (N_16175,N_13313,N_14909);
or U16176 (N_16176,N_12018,N_10332);
nor U16177 (N_16177,N_11446,N_12562);
nor U16178 (N_16178,N_10062,N_11947);
and U16179 (N_16179,N_10952,N_12578);
nor U16180 (N_16180,N_10637,N_12580);
and U16181 (N_16181,N_11611,N_12687);
nor U16182 (N_16182,N_14514,N_14336);
nand U16183 (N_16183,N_13523,N_10111);
or U16184 (N_16184,N_12360,N_10883);
nor U16185 (N_16185,N_14805,N_14271);
nor U16186 (N_16186,N_12243,N_11799);
or U16187 (N_16187,N_10089,N_13100);
nand U16188 (N_16188,N_13927,N_14859);
or U16189 (N_16189,N_13260,N_11587);
or U16190 (N_16190,N_12790,N_11304);
nor U16191 (N_16191,N_13330,N_11638);
nand U16192 (N_16192,N_13048,N_14820);
nand U16193 (N_16193,N_14338,N_13659);
nand U16194 (N_16194,N_12616,N_14151);
nand U16195 (N_16195,N_14043,N_12764);
and U16196 (N_16196,N_10741,N_13117);
nor U16197 (N_16197,N_13046,N_14920);
nor U16198 (N_16198,N_13780,N_12173);
and U16199 (N_16199,N_12232,N_14181);
nor U16200 (N_16200,N_12856,N_10272);
or U16201 (N_16201,N_11454,N_13824);
nand U16202 (N_16202,N_11864,N_10909);
nand U16203 (N_16203,N_11362,N_10457);
and U16204 (N_16204,N_11492,N_14084);
nor U16205 (N_16205,N_12826,N_10897);
nor U16206 (N_16206,N_12836,N_14375);
and U16207 (N_16207,N_13600,N_13713);
nor U16208 (N_16208,N_11686,N_11249);
nor U16209 (N_16209,N_13442,N_11822);
nor U16210 (N_16210,N_12529,N_12452);
or U16211 (N_16211,N_14984,N_13821);
and U16212 (N_16212,N_13539,N_11571);
nand U16213 (N_16213,N_11848,N_11045);
nor U16214 (N_16214,N_12305,N_10343);
nor U16215 (N_16215,N_10955,N_11049);
or U16216 (N_16216,N_10936,N_13462);
nand U16217 (N_16217,N_10361,N_14113);
nand U16218 (N_16218,N_13044,N_13955);
nand U16219 (N_16219,N_12259,N_12365);
nor U16220 (N_16220,N_11081,N_10653);
nor U16221 (N_16221,N_11513,N_12045);
nand U16222 (N_16222,N_14518,N_14737);
and U16223 (N_16223,N_10493,N_11569);
nand U16224 (N_16224,N_11538,N_10984);
and U16225 (N_16225,N_14515,N_12999);
or U16226 (N_16226,N_11013,N_10432);
or U16227 (N_16227,N_11675,N_13252);
or U16228 (N_16228,N_11870,N_12515);
or U16229 (N_16229,N_14890,N_14394);
and U16230 (N_16230,N_13693,N_12237);
nor U16231 (N_16231,N_13007,N_11282);
or U16232 (N_16232,N_10360,N_12376);
or U16233 (N_16233,N_11009,N_10357);
nand U16234 (N_16234,N_13041,N_11473);
nor U16235 (N_16235,N_10771,N_14504);
nor U16236 (N_16236,N_14147,N_10140);
or U16237 (N_16237,N_10561,N_11147);
or U16238 (N_16238,N_14908,N_14053);
or U16239 (N_16239,N_10486,N_10530);
nand U16240 (N_16240,N_10977,N_12134);
nand U16241 (N_16241,N_10744,N_10075);
or U16242 (N_16242,N_13941,N_13730);
or U16243 (N_16243,N_13094,N_11346);
and U16244 (N_16244,N_13164,N_13904);
and U16245 (N_16245,N_11029,N_14497);
nor U16246 (N_16246,N_12774,N_10159);
or U16247 (N_16247,N_14734,N_13782);
nand U16248 (N_16248,N_10341,N_13814);
nor U16249 (N_16249,N_14598,N_10479);
xor U16250 (N_16250,N_11667,N_11982);
or U16251 (N_16251,N_13344,N_11253);
nor U16252 (N_16252,N_14507,N_14246);
nor U16253 (N_16253,N_14781,N_10020);
nor U16254 (N_16254,N_14282,N_10054);
and U16255 (N_16255,N_13221,N_12127);
nor U16256 (N_16256,N_12088,N_10879);
and U16257 (N_16257,N_11293,N_12492);
nor U16258 (N_16258,N_10768,N_13654);
or U16259 (N_16259,N_10067,N_11858);
and U16260 (N_16260,N_12629,N_12744);
nor U16261 (N_16261,N_11255,N_12896);
and U16262 (N_16262,N_12627,N_12440);
nand U16263 (N_16263,N_10175,N_13451);
and U16264 (N_16264,N_12990,N_14951);
or U16265 (N_16265,N_13597,N_11109);
and U16266 (N_16266,N_13899,N_12830);
nor U16267 (N_16267,N_13491,N_12649);
nor U16268 (N_16268,N_13842,N_13435);
nor U16269 (N_16269,N_14558,N_13961);
nand U16270 (N_16270,N_14212,N_10799);
and U16271 (N_16271,N_11015,N_10185);
and U16272 (N_16272,N_13852,N_14001);
nor U16273 (N_16273,N_12101,N_12804);
and U16274 (N_16274,N_13384,N_10760);
and U16275 (N_16275,N_10149,N_10137);
or U16276 (N_16276,N_12449,N_11548);
nand U16277 (N_16277,N_14838,N_14031);
nand U16278 (N_16278,N_11218,N_10745);
nor U16279 (N_16279,N_12165,N_10365);
nor U16280 (N_16280,N_11506,N_12002);
and U16281 (N_16281,N_13583,N_10156);
nor U16282 (N_16282,N_14694,N_14004);
nor U16283 (N_16283,N_13251,N_10708);
nor U16284 (N_16284,N_11952,N_11156);
and U16285 (N_16285,N_10570,N_11763);
nand U16286 (N_16286,N_11750,N_11794);
or U16287 (N_16287,N_10939,N_10988);
nor U16288 (N_16288,N_12286,N_12913);
nor U16289 (N_16289,N_13601,N_10518);
nor U16290 (N_16290,N_12976,N_12267);
or U16291 (N_16291,N_11679,N_12858);
nand U16292 (N_16292,N_11120,N_12371);
nand U16293 (N_16293,N_12833,N_14893);
nor U16294 (N_16294,N_12889,N_11070);
and U16295 (N_16295,N_11134,N_11944);
nor U16296 (N_16296,N_12508,N_12484);
nor U16297 (N_16297,N_10152,N_12141);
or U16298 (N_16298,N_12965,N_13198);
xor U16299 (N_16299,N_14943,N_10264);
and U16300 (N_16300,N_12954,N_10894);
or U16301 (N_16301,N_13748,N_12866);
nand U16302 (N_16302,N_12903,N_14101);
or U16303 (N_16303,N_14210,N_11017);
or U16304 (N_16304,N_12358,N_12823);
nor U16305 (N_16305,N_12743,N_11978);
and U16306 (N_16306,N_11819,N_13627);
or U16307 (N_16307,N_14776,N_14982);
or U16308 (N_16308,N_12156,N_12263);
xor U16309 (N_16309,N_14358,N_13239);
nand U16310 (N_16310,N_10407,N_10739);
and U16311 (N_16311,N_10811,N_10589);
or U16312 (N_16312,N_12022,N_14243);
and U16313 (N_16313,N_10735,N_14834);
nor U16314 (N_16314,N_11740,N_12222);
or U16315 (N_16315,N_11138,N_10979);
and U16316 (N_16316,N_14746,N_12334);
nor U16317 (N_16317,N_10350,N_13667);
and U16318 (N_16318,N_13686,N_12258);
nand U16319 (N_16319,N_10454,N_11368);
nand U16320 (N_16320,N_12897,N_14126);
and U16321 (N_16321,N_10998,N_14415);
or U16322 (N_16322,N_10944,N_13835);
or U16323 (N_16323,N_10231,N_12684);
nor U16324 (N_16324,N_11431,N_10171);
or U16325 (N_16325,N_12880,N_12430);
nand U16326 (N_16326,N_10496,N_13151);
and U16327 (N_16327,N_14888,N_14600);
nor U16328 (N_16328,N_13565,N_13699);
and U16329 (N_16329,N_11989,N_14896);
nand U16330 (N_16330,N_12103,N_13199);
nand U16331 (N_16331,N_11710,N_11902);
or U16332 (N_16332,N_13593,N_14553);
and U16333 (N_16333,N_14502,N_12420);
nor U16334 (N_16334,N_14266,N_13085);
or U16335 (N_16335,N_14094,N_10391);
and U16336 (N_16336,N_14937,N_12182);
and U16337 (N_16337,N_12406,N_14078);
and U16338 (N_16338,N_12028,N_10792);
nor U16339 (N_16339,N_14496,N_12423);
nor U16340 (N_16340,N_12069,N_12623);
nand U16341 (N_16341,N_13676,N_13368);
and U16342 (N_16342,N_13573,N_10138);
and U16343 (N_16343,N_12536,N_11270);
nor U16344 (N_16344,N_14134,N_11929);
and U16345 (N_16345,N_14122,N_13957);
nor U16346 (N_16346,N_13342,N_10654);
nor U16347 (N_16347,N_14057,N_11074);
and U16348 (N_16348,N_14671,N_10109);
nor U16349 (N_16349,N_11025,N_14688);
nand U16350 (N_16350,N_13412,N_10578);
or U16351 (N_16351,N_14187,N_14510);
nor U16352 (N_16352,N_11194,N_14989);
nand U16353 (N_16353,N_13013,N_10969);
and U16354 (N_16354,N_10249,N_10598);
nor U16355 (N_16355,N_14822,N_12476);
nand U16356 (N_16356,N_11332,N_14853);
nor U16357 (N_16357,N_12279,N_11765);
nor U16358 (N_16358,N_13506,N_12617);
and U16359 (N_16359,N_14548,N_12519);
nor U16360 (N_16360,N_14149,N_14567);
or U16361 (N_16361,N_13816,N_11036);
or U16362 (N_16362,N_14228,N_14235);
nor U16363 (N_16363,N_14977,N_12806);
nor U16364 (N_16364,N_12946,N_14639);
and U16365 (N_16365,N_14140,N_13808);
xnor U16366 (N_16366,N_12008,N_10308);
nand U16367 (N_16367,N_11528,N_12302);
and U16368 (N_16368,N_10507,N_12172);
or U16369 (N_16369,N_10762,N_13243);
nor U16370 (N_16370,N_12818,N_11880);
nor U16371 (N_16371,N_13335,N_10422);
nor U16372 (N_16372,N_10050,N_10717);
and U16373 (N_16373,N_11341,N_10151);
nand U16374 (N_16374,N_13683,N_14028);
nor U16375 (N_16375,N_12505,N_10835);
nor U16376 (N_16376,N_10384,N_12753);
nand U16377 (N_16377,N_11558,N_13139);
and U16378 (N_16378,N_14030,N_11494);
nor U16379 (N_16379,N_13171,N_14545);
or U16380 (N_16380,N_12228,N_14975);
or U16381 (N_16381,N_12465,N_10052);
or U16382 (N_16382,N_12760,N_12670);
and U16383 (N_16383,N_11682,N_13678);
nand U16384 (N_16384,N_11640,N_12857);
xnor U16385 (N_16385,N_11330,N_10021);
xor U16386 (N_16386,N_11901,N_13935);
nor U16387 (N_16387,N_13533,N_14344);
and U16388 (N_16388,N_10379,N_11537);
nor U16389 (N_16389,N_14609,N_14773);
and U16390 (N_16390,N_11791,N_11169);
nand U16391 (N_16391,N_14589,N_13200);
and U16392 (N_16392,N_11586,N_12450);
nand U16393 (N_16393,N_12655,N_14366);
nand U16394 (N_16394,N_13703,N_14359);
and U16395 (N_16395,N_13968,N_10891);
nand U16396 (N_16396,N_13966,N_10117);
nand U16397 (N_16397,N_14840,N_14865);
and U16398 (N_16398,N_11030,N_13241);
or U16399 (N_16399,N_12408,N_11570);
nor U16400 (N_16400,N_12310,N_12007);
nand U16401 (N_16401,N_11378,N_11488);
nor U16402 (N_16402,N_14027,N_14418);
and U16403 (N_16403,N_11942,N_12986);
nor U16404 (N_16404,N_14040,N_10484);
xor U16405 (N_16405,N_12960,N_11589);
nor U16406 (N_16406,N_14875,N_13830);
or U16407 (N_16407,N_12067,N_13112);
nand U16408 (N_16408,N_12906,N_11419);
or U16409 (N_16409,N_12315,N_14661);
nand U16410 (N_16410,N_12428,N_13375);
nand U16411 (N_16411,N_13297,N_13850);
nand U16412 (N_16412,N_11417,N_10529);
or U16413 (N_16413,N_13794,N_13280);
or U16414 (N_16414,N_10603,N_13460);
and U16415 (N_16415,N_11380,N_10465);
nor U16416 (N_16416,N_13235,N_12227);
or U16417 (N_16417,N_12814,N_14560);
and U16418 (N_16418,N_11677,N_12685);
nor U16419 (N_16419,N_14109,N_14105);
nand U16420 (N_16420,N_11716,N_12904);
nand U16421 (N_16421,N_12188,N_14088);
or U16422 (N_16422,N_13466,N_13205);
nor U16423 (N_16423,N_10102,N_13445);
and U16424 (N_16424,N_10720,N_10753);
nand U16425 (N_16425,N_12973,N_14125);
or U16426 (N_16426,N_11658,N_11531);
or U16427 (N_16427,N_10865,N_12734);
nand U16428 (N_16428,N_14682,N_11958);
and U16429 (N_16429,N_13819,N_13723);
and U16430 (N_16430,N_14491,N_13322);
nand U16431 (N_16431,N_12291,N_14305);
or U16432 (N_16432,N_13503,N_11715);
or U16433 (N_16433,N_11547,N_12164);
nand U16434 (N_16434,N_10960,N_11397);
or U16435 (N_16435,N_12122,N_12017);
nor U16436 (N_16436,N_12171,N_14192);
and U16437 (N_16437,N_14704,N_13177);
nand U16438 (N_16438,N_14226,N_13264);
nor U16439 (N_16439,N_12625,N_10997);
nor U16440 (N_16440,N_11807,N_11472);
nor U16441 (N_16441,N_13578,N_11776);
and U16442 (N_16442,N_11337,N_11203);
or U16443 (N_16443,N_11205,N_14708);
nor U16444 (N_16444,N_10003,N_11974);
or U16445 (N_16445,N_13182,N_11260);
or U16446 (N_16446,N_14193,N_14856);
nor U16447 (N_16447,N_12703,N_10096);
nand U16448 (N_16448,N_11100,N_14299);
or U16449 (N_16449,N_12337,N_13502);
nor U16450 (N_16450,N_14356,N_10051);
or U16451 (N_16451,N_11773,N_14019);
nand U16452 (N_16452,N_12339,N_10435);
or U16453 (N_16453,N_11301,N_12816);
and U16454 (N_16454,N_14724,N_11410);
or U16455 (N_16455,N_13891,N_14597);
and U16456 (N_16456,N_13972,N_13093);
nor U16457 (N_16457,N_14855,N_12480);
nor U16458 (N_16458,N_12624,N_10238);
nor U16459 (N_16459,N_13359,N_12323);
nand U16460 (N_16460,N_11296,N_11968);
or U16461 (N_16461,N_13704,N_11820);
nand U16462 (N_16462,N_11699,N_12530);
nand U16463 (N_16463,N_14976,N_12126);
nand U16464 (N_16464,N_10513,N_11703);
and U16465 (N_16465,N_13232,N_10497);
nor U16466 (N_16466,N_13663,N_10090);
or U16467 (N_16467,N_14083,N_10956);
or U16468 (N_16468,N_14051,N_11388);
nor U16469 (N_16469,N_10263,N_12436);
or U16470 (N_16470,N_10256,N_12168);
and U16471 (N_16471,N_14013,N_14561);
nor U16472 (N_16472,N_11628,N_11455);
and U16473 (N_16473,N_11867,N_12441);
and U16474 (N_16474,N_11267,N_12911);
or U16475 (N_16475,N_13800,N_14674);
nand U16476 (N_16476,N_10881,N_14276);
and U16477 (N_16477,N_13448,N_14251);
nand U16478 (N_16478,N_11056,N_12738);
nand U16479 (N_16479,N_11144,N_10577);
or U16480 (N_16480,N_11003,N_11888);
nand U16481 (N_16481,N_10356,N_14577);
nor U16482 (N_16482,N_11412,N_10675);
or U16483 (N_16483,N_14023,N_14152);
and U16484 (N_16484,N_10691,N_14196);
and U16485 (N_16485,N_11108,N_12854);
nand U16486 (N_16486,N_14957,N_12704);
or U16487 (N_16487,N_11986,N_11316);
or U16488 (N_16488,N_11887,N_10558);
or U16489 (N_16489,N_11948,N_10429);
nand U16490 (N_16490,N_12781,N_14621);
or U16491 (N_16491,N_14792,N_13190);
nand U16492 (N_16492,N_12756,N_13837);
nor U16493 (N_16493,N_10822,N_14537);
nand U16494 (N_16494,N_12460,N_13318);
or U16495 (N_16495,N_10824,N_14050);
nor U16496 (N_16496,N_10018,N_11911);
nor U16497 (N_16497,N_12545,N_11972);
nor U16498 (N_16498,N_11089,N_13548);
and U16499 (N_16499,N_11428,N_12864);
nor U16500 (N_16500,N_13889,N_11116);
nor U16501 (N_16501,N_11796,N_11496);
and U16502 (N_16502,N_10472,N_14971);
and U16503 (N_16503,N_14135,N_10053);
or U16504 (N_16504,N_10248,N_13275);
nor U16505 (N_16505,N_11685,N_14277);
or U16506 (N_16506,N_10526,N_14263);
and U16507 (N_16507,N_12933,N_11956);
and U16508 (N_16508,N_12694,N_14360);
nor U16509 (N_16509,N_14527,N_13952);
and U16510 (N_16510,N_13538,N_11192);
and U16511 (N_16511,N_14684,N_14314);
and U16512 (N_16512,N_11182,N_12297);
nor U16513 (N_16513,N_12654,N_11599);
nor U16514 (N_16514,N_13310,N_12059);
or U16515 (N_16515,N_11269,N_11395);
nand U16516 (N_16516,N_11855,N_13979);
nor U16517 (N_16517,N_11607,N_12307);
nor U16518 (N_16518,N_10392,N_14390);
or U16519 (N_16519,N_12967,N_13097);
and U16520 (N_16520,N_11026,N_12125);
nand U16521 (N_16521,N_11917,N_10139);
or U16522 (N_16522,N_12872,N_11050);
and U16523 (N_16523,N_11930,N_13253);
nand U16524 (N_16524,N_13843,N_10146);
nand U16525 (N_16525,N_11616,N_13387);
or U16526 (N_16526,N_13604,N_10902);
nor U16527 (N_16527,N_12057,N_14956);
or U16528 (N_16528,N_13577,N_13924);
and U16529 (N_16529,N_11257,N_13828);
or U16530 (N_16530,N_14076,N_12275);
or U16531 (N_16531,N_12169,N_11068);
and U16532 (N_16532,N_14431,N_10854);
nand U16533 (N_16533,N_12523,N_13175);
nor U16534 (N_16534,N_10322,N_11553);
nor U16535 (N_16535,N_13938,N_13471);
or U16536 (N_16536,N_14717,N_12870);
and U16537 (N_16537,N_11167,N_10743);
nor U16538 (N_16538,N_10433,N_12357);
or U16539 (N_16539,N_10752,N_14115);
nor U16540 (N_16540,N_10790,N_13249);
nor U16541 (N_16541,N_10410,N_10671);
or U16542 (N_16542,N_14354,N_12584);
and U16543 (N_16543,N_12533,N_13606);
nor U16544 (N_16544,N_14710,N_13361);
nand U16545 (N_16545,N_10532,N_11967);
nor U16546 (N_16546,N_11645,N_13811);
nand U16547 (N_16547,N_10416,N_11476);
nand U16548 (N_16548,N_13119,N_10293);
nand U16549 (N_16549,N_13928,N_11894);
nand U16550 (N_16550,N_11837,N_12574);
or U16551 (N_16551,N_11891,N_11442);
nor U16552 (N_16552,N_11545,N_10950);
nand U16553 (N_16553,N_12110,N_13279);
nor U16554 (N_16554,N_10469,N_14405);
or U16555 (N_16555,N_14166,N_12276);
or U16556 (N_16556,N_11801,N_12672);
nor U16557 (N_16557,N_13088,N_13796);
nand U16558 (N_16558,N_13750,N_11874);
nand U16559 (N_16559,N_10876,N_10475);
nand U16560 (N_16560,N_13082,N_12496);
or U16561 (N_16561,N_13016,N_11071);
or U16562 (N_16562,N_13223,N_12663);
nand U16563 (N_16563,N_13231,N_11206);
nor U16564 (N_16564,N_13095,N_14905);
nand U16565 (N_16565,N_10046,N_11945);
or U16566 (N_16566,N_14605,N_10503);
and U16567 (N_16567,N_13098,N_14685);
and U16568 (N_16568,N_13153,N_14353);
nand U16569 (N_16569,N_10931,N_12742);
and U16570 (N_16570,N_11577,N_10758);
nand U16571 (N_16571,N_12058,N_11781);
nand U16572 (N_16572,N_14555,N_10802);
nand U16573 (N_16573,N_11315,N_10916);
nor U16574 (N_16574,N_12881,N_11621);
nand U16575 (N_16575,N_13001,N_13839);
nand U16576 (N_16576,N_10805,N_12883);
nor U16577 (N_16577,N_11600,N_14199);
or U16578 (N_16578,N_12586,N_13576);
or U16579 (N_16579,N_10651,N_12011);
nor U16580 (N_16580,N_10045,N_10565);
and U16581 (N_16581,N_14460,N_14216);
nor U16582 (N_16582,N_12819,N_13026);
nor U16583 (N_16583,N_11023,N_11317);
nor U16584 (N_16584,N_12415,N_11365);
nand U16585 (N_16585,N_10582,N_10514);
and U16586 (N_16586,N_10121,N_10396);
or U16587 (N_16587,N_13463,N_11430);
nor U16588 (N_16588,N_13337,N_14006);
nand U16589 (N_16589,N_13440,N_14997);
and U16590 (N_16590,N_12642,N_11863);
and U16591 (N_16591,N_11204,N_12571);
and U16592 (N_16592,N_12598,N_14468);
or U16593 (N_16593,N_11098,N_12607);
nand U16594 (N_16594,N_14328,N_14891);
nor U16595 (N_16595,N_14880,N_13855);
nand U16596 (N_16596,N_11302,N_14020);
or U16597 (N_16597,N_11693,N_13890);
or U16598 (N_16598,N_14403,N_11912);
or U16599 (N_16599,N_10166,N_11572);
or U16600 (N_16600,N_14757,N_11146);
nor U16601 (N_16601,N_12658,N_13364);
or U16602 (N_16602,N_12439,N_11932);
nand U16603 (N_16603,N_10409,N_11597);
nor U16604 (N_16604,N_11757,N_11391);
nor U16605 (N_16605,N_11749,N_10957);
or U16606 (N_16606,N_10153,N_12601);
and U16607 (N_16607,N_14329,N_14112);
or U16608 (N_16608,N_10267,N_14532);
nor U16609 (N_16609,N_12487,N_10901);
nand U16610 (N_16610,N_13130,N_11637);
and U16611 (N_16611,N_11335,N_14104);
nor U16612 (N_16612,N_12983,N_14873);
and U16613 (N_16613,N_14524,N_10954);
nand U16614 (N_16614,N_11823,N_11288);
and U16615 (N_16615,N_11069,N_11767);
or U16616 (N_16616,N_11500,N_13702);
or U16617 (N_16617,N_14236,N_11882);
and U16618 (N_16618,N_11199,N_11700);
nand U16619 (N_16619,N_14934,N_10629);
and U16620 (N_16620,N_13945,N_12475);
or U16621 (N_16621,N_11229,N_10083);
and U16622 (N_16622,N_14171,N_10316);
or U16623 (N_16623,N_11408,N_10678);
or U16624 (N_16624,N_13054,N_13925);
nand U16625 (N_16625,N_10856,N_12319);
nand U16626 (N_16626,N_13312,N_11087);
nor U16627 (N_16627,N_11236,N_11585);
and U16628 (N_16628,N_12525,N_13488);
and U16629 (N_16629,N_10312,N_13338);
or U16630 (N_16630,N_13861,N_14998);
nand U16631 (N_16631,N_13848,N_10685);
nor U16632 (N_16632,N_11211,N_14275);
nor U16633 (N_16633,N_10425,N_11521);
and U16634 (N_16634,N_10011,N_10806);
nand U16635 (N_16635,N_11298,N_14879);
and U16636 (N_16636,N_12548,N_11053);
and U16637 (N_16637,N_10825,N_10791);
or U16638 (N_16638,N_11535,N_12995);
nor U16639 (N_16639,N_14401,N_11790);
nor U16640 (N_16640,N_13810,N_11499);
and U16641 (N_16641,N_13030,N_11996);
nor U16642 (N_16642,N_10145,N_14313);
nand U16643 (N_16643,N_11828,N_14201);
or U16644 (N_16644,N_10841,N_12982);
nor U16645 (N_16645,N_13064,N_12721);
nor U16646 (N_16646,N_12288,N_14029);
nor U16647 (N_16647,N_14465,N_14744);
and U16648 (N_16648,N_14716,N_13616);
nand U16649 (N_16649,N_13128,N_10188);
nor U16650 (N_16650,N_13483,N_12602);
or U16651 (N_16651,N_11593,N_13776);
nand U16652 (N_16652,N_12662,N_11226);
nor U16653 (N_16653,N_13896,N_13634);
or U16654 (N_16654,N_14756,N_12354);
nand U16655 (N_16655,N_14904,N_10271);
or U16656 (N_16656,N_12026,N_14749);
or U16657 (N_16657,N_10528,N_10964);
nor U16658 (N_16658,N_10836,N_14690);
nor U16659 (N_16659,N_13715,N_10846);
or U16660 (N_16660,N_12092,N_10549);
nand U16661 (N_16661,N_14992,N_12152);
nand U16662 (N_16662,N_14141,N_13511);
nor U16663 (N_16663,N_10094,N_14383);
nor U16664 (N_16664,N_14498,N_10614);
nand U16665 (N_16665,N_10649,N_13217);
or U16666 (N_16666,N_13705,N_13194);
or U16667 (N_16667,N_14525,N_11379);
and U16668 (N_16668,N_12128,N_12615);
nor U16669 (N_16669,N_11991,N_13527);
or U16670 (N_16670,N_10103,N_12196);
and U16671 (N_16671,N_12273,N_13061);
nor U16672 (N_16672,N_12407,N_11084);
nor U16673 (N_16673,N_11409,N_10915);
and U16674 (N_16674,N_12644,N_12042);
nand U16675 (N_16675,N_13528,N_14655);
and U16676 (N_16676,N_12336,N_14867);
or U16677 (N_16677,N_14014,N_12677);
nand U16678 (N_16678,N_14731,N_14848);
nor U16679 (N_16679,N_12538,N_11533);
and U16680 (N_16680,N_14287,N_13383);
nand U16681 (N_16681,N_12349,N_11634);
nor U16682 (N_16682,N_12815,N_10128);
nand U16683 (N_16683,N_13034,N_14648);
and U16684 (N_16684,N_13049,N_11436);
and U16685 (N_16685,N_11605,N_13336);
and U16686 (N_16686,N_11038,N_13393);
or U16687 (N_16687,N_13323,N_12517);
nor U16688 (N_16688,N_13661,N_14614);
and U16689 (N_16689,N_13135,N_14167);
and U16690 (N_16690,N_10898,N_12130);
nor U16691 (N_16691,N_10190,N_14759);
nor U16692 (N_16692,N_12433,N_10344);
nor U16693 (N_16693,N_11613,N_13214);
nand U16694 (N_16694,N_14046,N_10461);
or U16695 (N_16695,N_14168,N_12086);
and U16696 (N_16696,N_13680,N_10987);
nor U16697 (N_16697,N_12111,N_14669);
and U16698 (N_16698,N_13469,N_14066);
nor U16699 (N_16699,N_13137,N_13745);
or U16700 (N_16700,N_14206,N_11102);
nand U16701 (N_16701,N_14488,N_10063);
nor U16702 (N_16702,N_14626,N_11804);
nor U16703 (N_16703,N_11131,N_12062);
nand U16704 (N_16704,N_13624,N_10693);
and U16705 (N_16705,N_14691,N_14016);
or U16706 (N_16706,N_11072,N_13507);
and U16707 (N_16707,N_12759,N_14972);
nand U16708 (N_16708,N_10452,N_13555);
nor U16709 (N_16709,N_10573,N_12367);
nor U16710 (N_16710,N_14808,N_12120);
and U16711 (N_16711,N_12590,N_10397);
and U16712 (N_16712,N_13870,N_14876);
nor U16713 (N_16713,N_14111,N_11223);
and U16714 (N_16714,N_11238,N_11343);
nor U16715 (N_16715,N_14062,N_11674);
or U16716 (N_16716,N_10487,N_10851);
nor U16717 (N_16717,N_13183,N_11993);
nor U16718 (N_16718,N_11207,N_12043);
nor U16719 (N_16719,N_13057,N_12016);
and U16720 (N_16720,N_11390,N_14922);
nand U16721 (N_16721,N_13060,N_12489);
nor U16722 (N_16722,N_14208,N_13305);
or U16723 (N_16723,N_14794,N_11005);
nand U16724 (N_16724,N_10029,N_11601);
and U16725 (N_16725,N_12457,N_11292);
nor U16726 (N_16726,N_13965,N_14635);
or U16727 (N_16727,N_12121,N_10923);
nor U16728 (N_16728,N_12682,N_12158);
and U16729 (N_16729,N_10896,N_13381);
or U16730 (N_16730,N_12350,N_14884);
nor U16731 (N_16731,N_10816,N_11366);
nand U16732 (N_16732,N_10658,N_13803);
nand U16733 (N_16733,N_10205,N_10505);
nor U16734 (N_16734,N_12860,N_10317);
or U16735 (N_16735,N_13162,N_14472);
and U16736 (N_16736,N_13696,N_14485);
and U16737 (N_16737,N_14154,N_11976);
nand U16738 (N_16738,N_14623,N_11019);
nand U16739 (N_16739,N_11387,N_14355);
or U16740 (N_16740,N_14024,N_12000);
nand U16741 (N_16741,N_13332,N_14657);
or U16742 (N_16742,N_10186,N_10686);
nor U16743 (N_16743,N_10519,N_12226);
nand U16744 (N_16744,N_13559,N_10351);
nand U16745 (N_16745,N_10542,N_11225);
or U16746 (N_16746,N_10633,N_10868);
nand U16747 (N_16747,N_11340,N_10047);
nor U16748 (N_16748,N_13543,N_10730);
or U16749 (N_16749,N_13404,N_13428);
nor U16750 (N_16750,N_11508,N_12885);
nor U16751 (N_16751,N_13695,N_13755);
nor U16752 (N_16752,N_14281,N_13400);
or U16753 (N_16753,N_13437,N_10214);
nand U16754 (N_16754,N_13120,N_14294);
nor U16755 (N_16755,N_10430,N_11652);
nand U16756 (N_16756,N_11078,N_10592);
or U16757 (N_16757,N_13343,N_10265);
nand U16758 (N_16758,N_12143,N_14347);
nor U16759 (N_16759,N_13736,N_11815);
or U16760 (N_16760,N_11946,N_14451);
and U16761 (N_16761,N_12770,N_11626);
or U16762 (N_16762,N_13058,N_11123);
nor U16763 (N_16763,N_10201,N_11914);
nand U16764 (N_16764,N_10085,N_13430);
nand U16765 (N_16765,N_10431,N_14272);
or U16766 (N_16766,N_12262,N_13605);
and U16767 (N_16767,N_13407,N_14990);
and U16768 (N_16768,N_10627,N_13716);
nor U16769 (N_16769,N_10016,N_11165);
and U16770 (N_16770,N_14546,N_11980);
or U16771 (N_16771,N_11040,N_10714);
or U16772 (N_16772,N_13888,N_13637);
or U16773 (N_16773,N_10108,N_13133);
or U16774 (N_16774,N_12037,N_14161);
or U16775 (N_16775,N_12019,N_13976);
or U16776 (N_16776,N_11000,N_11937);
and U16777 (N_16777,N_13339,N_12540);
nand U16778 (N_16778,N_10850,N_12915);
or U16779 (N_16779,N_12504,N_14714);
and U16780 (N_16780,N_10848,N_14400);
nor U16781 (N_16781,N_10812,N_11467);
or U16782 (N_16782,N_13849,N_13906);
nand U16783 (N_16783,N_10537,N_10576);
nor U16784 (N_16784,N_11842,N_12140);
and U16785 (N_16785,N_13293,N_10076);
nor U16786 (N_16786,N_14017,N_10681);
nor U16787 (N_16787,N_14950,N_13123);
or U16788 (N_16788,N_10834,N_10110);
or U16789 (N_16789,N_10233,N_10607);
or U16790 (N_16790,N_12714,N_10912);
xor U16791 (N_16791,N_14090,N_11491);
nor U16792 (N_16792,N_11064,N_14907);
or U16793 (N_16793,N_14947,N_13269);
and U16794 (N_16794,N_13995,N_14092);
and U16795 (N_16795,N_11818,N_12579);
nor U16796 (N_16796,N_11439,N_14810);
nand U16797 (N_16797,N_10663,N_14595);
nand U16798 (N_16798,N_12970,N_11832);
and U16799 (N_16799,N_14423,N_11859);
and U16800 (N_16800,N_11208,N_11526);
nand U16801 (N_16801,N_14958,N_11364);
nor U16802 (N_16802,N_12375,N_14486);
nand U16803 (N_16803,N_11164,N_11892);
and U16804 (N_16804,N_13922,N_10398);
or U16805 (N_16805,N_12318,N_14991);
nor U16806 (N_16806,N_10963,N_14817);
nor U16807 (N_16807,N_10840,N_13621);
or U16808 (N_16808,N_13050,N_13454);
nand U16809 (N_16809,N_10495,N_10610);
and U16810 (N_16810,N_14309,N_14248);
and U16811 (N_16811,N_11244,N_12347);
or U16812 (N_16812,N_13515,N_13441);
or U16813 (N_16813,N_10358,N_11905);
and U16814 (N_16814,N_10460,N_11762);
and U16815 (N_16815,N_12527,N_11532);
nand U16816 (N_16816,N_14183,N_13689);
nor U16817 (N_16817,N_13168,N_14351);
nand U16818 (N_16818,N_10032,N_10383);
nand U16819 (N_16819,N_11543,N_10335);
or U16820 (N_16820,N_14961,N_12972);
nand U16821 (N_16821,N_11278,N_10907);
nor U16822 (N_16822,N_12136,N_14288);
nand U16823 (N_16823,N_10005,N_14160);
and U16824 (N_16824,N_14667,N_13015);
nor U16825 (N_16825,N_12455,N_10228);
and U16826 (N_16826,N_11869,N_13289);
and U16827 (N_16827,N_13974,N_13951);
nand U16828 (N_16828,N_11066,N_11037);
and U16829 (N_16829,N_13662,N_13642);
and U16830 (N_16830,N_12251,N_14531);
and U16831 (N_16831,N_10641,N_13141);
nand U16832 (N_16832,N_11219,N_14556);
nand U16833 (N_16833,N_10441,N_10521);
nand U16834 (N_16834,N_13367,N_13107);
nor U16835 (N_16835,N_11216,N_11426);
nor U16836 (N_16836,N_10220,N_12199);
or U16837 (N_16837,N_10525,N_13544);
and U16838 (N_16838,N_14118,N_13921);
nand U16839 (N_16839,N_11398,N_14929);
nor U16840 (N_16840,N_14536,N_12934);
nand U16841 (N_16841,N_13526,N_10662);
and U16842 (N_16842,N_13452,N_10266);
and U16843 (N_16843,N_12638,N_12394);
nand U16844 (N_16844,N_13186,N_12114);
or U16845 (N_16845,N_11825,N_14380);
and U16846 (N_16846,N_12600,N_11782);
nand U16847 (N_16847,N_13619,N_12564);
nor U16848 (N_16848,N_12867,N_12192);
or U16849 (N_16849,N_10706,N_13003);
or U16850 (N_16850,N_10230,N_14936);
or U16851 (N_16851,N_10546,N_12015);
or U16852 (N_16852,N_12175,N_12521);
nand U16853 (N_16853,N_14185,N_13632);
nand U16854 (N_16854,N_12936,N_10749);
nor U16855 (N_16855,N_13879,N_11747);
or U16856 (N_16856,N_10559,N_14240);
and U16857 (N_16857,N_11581,N_11995);
nand U16858 (N_16858,N_13494,N_12317);
nand U16859 (N_16859,N_13992,N_14108);
and U16860 (N_16860,N_14164,N_11668);
nor U16861 (N_16861,N_13011,N_13482);
nor U16862 (N_16862,N_10327,N_12132);
or U16863 (N_16863,N_12020,N_13480);
and U16864 (N_16864,N_10517,N_12071);
nand U16865 (N_16865,N_14665,N_14948);
and U16866 (N_16866,N_13792,N_14081);
or U16867 (N_16867,N_11889,N_12177);
and U16868 (N_16868,N_11276,N_11928);
nor U16869 (N_16869,N_14966,N_11979);
nor U16870 (N_16870,N_12528,N_12659);
nor U16871 (N_16871,N_11681,N_12084);
and U16872 (N_16872,N_11672,N_10382);
nand U16873 (N_16873,N_12560,N_12959);
nor U16874 (N_16874,N_13729,N_10748);
and U16875 (N_16875,N_14054,N_12342);
and U16876 (N_16876,N_14032,N_12208);
and U16877 (N_16877,N_11729,N_11305);
nand U16878 (N_16878,N_11347,N_11838);
or U16879 (N_16879,N_13405,N_10326);
or U16880 (N_16880,N_10499,N_11758);
or U16881 (N_16881,N_14523,N_14687);
and U16882 (N_16882,N_14335,N_10232);
or U16883 (N_16883,N_12106,N_13772);
nand U16884 (N_16884,N_10580,N_12186);
or U16885 (N_16885,N_12869,N_12552);
nand U16886 (N_16886,N_12454,N_12626);
nand U16887 (N_16887,N_14752,N_10059);
nand U16888 (N_16888,N_12888,N_12473);
nand U16889 (N_16889,N_12497,N_10761);
nand U16890 (N_16890,N_14678,N_11133);
or U16891 (N_16891,N_13797,N_11464);
and U16892 (N_16892,N_13761,N_10310);
and U16893 (N_16893,N_11363,N_11201);
and U16894 (N_16894,N_14601,N_14644);
or U16895 (N_16895,N_10828,N_11127);
and U16896 (N_16896,N_14588,N_12666);
nand U16897 (N_16897,N_14331,N_11161);
nor U16898 (N_16898,N_10359,N_11034);
nand U16899 (N_16899,N_13203,N_13132);
nor U16900 (N_16900,N_14506,N_10588);
xor U16901 (N_16901,N_11595,N_13258);
or U16902 (N_16902,N_14604,N_11118);
nor U16903 (N_16903,N_14503,N_14245);
nand U16904 (N_16904,N_13613,N_10242);
and U16905 (N_16905,N_12846,N_13567);
nand U16906 (N_16906,N_12160,N_12113);
or U16907 (N_16907,N_10869,N_12952);
nor U16908 (N_16908,N_12844,N_11451);
nor U16909 (N_16909,N_12513,N_12290);
or U16910 (N_16910,N_13547,N_14241);
nand U16911 (N_16911,N_10101,N_10683);
xor U16912 (N_16912,N_12981,N_12868);
and U16913 (N_16913,N_12432,N_14222);
or U16914 (N_16914,N_13595,N_11592);
nand U16915 (N_16915,N_13373,N_13101);
or U16916 (N_16916,N_14322,N_11449);
nor U16917 (N_16917,N_14107,N_11866);
or U16918 (N_16918,N_14723,N_12306);
or U16919 (N_16919,N_13167,N_13589);
and U16920 (N_16920,N_14227,N_11386);
nor U16921 (N_16921,N_13753,N_11814);
nor U16922 (N_16922,N_14302,N_12930);
nand U16923 (N_16923,N_14606,N_10989);
or U16924 (N_16924,N_12612,N_11872);
and U16925 (N_16925,N_10563,N_14872);
nand U16926 (N_16926,N_10782,N_10776);
xor U16927 (N_16927,N_11935,N_13947);
and U16928 (N_16928,N_14059,N_12462);
nor U16929 (N_16929,N_13341,N_10531);
nor U16930 (N_16930,N_13247,N_12474);
or U16931 (N_16931,N_13172,N_10819);
or U16932 (N_16932,N_12871,N_12068);
nor U16933 (N_16933,N_10763,N_11093);
nor U16934 (N_16934,N_10862,N_14903);
nor U16935 (N_16935,N_12162,N_13376);
nor U16936 (N_16936,N_12817,N_13369);
or U16937 (N_16937,N_13045,N_14034);
nor U16938 (N_16938,N_13287,N_13126);
nor U16939 (N_16939,N_14869,N_13887);
nor U16940 (N_16940,N_11551,N_11355);
and U16941 (N_16941,N_13883,N_14775);
nand U16942 (N_16942,N_12962,N_13898);
and U16943 (N_16943,N_10334,N_11286);
or U16944 (N_16944,N_11719,N_14061);
or U16945 (N_16945,N_12800,N_10789);
nor U16946 (N_16946,N_10154,N_11480);
or U16947 (N_16947,N_10867,N_14234);
nand U16948 (N_16948,N_11615,N_10839);
and U16949 (N_16949,N_14707,N_14350);
and U16950 (N_16950,N_13918,N_10055);
nor U16951 (N_16951,N_14267,N_11274);
or U16952 (N_16952,N_13684,N_13114);
and U16953 (N_16953,N_12346,N_12335);
nand U16954 (N_16954,N_14767,N_12381);
or U16955 (N_16955,N_14484,N_11567);
or U16956 (N_16956,N_12041,N_13862);
nand U16957 (N_16957,N_13781,N_11655);
or U16958 (N_16958,N_13625,N_10918);
nor U16959 (N_16959,N_14564,N_10440);
or U16960 (N_16960,N_14615,N_11429);
nand U16961 (N_16961,N_10778,N_13479);
nand U16962 (N_16962,N_13353,N_14565);
nand U16963 (N_16963,N_13806,N_14835);
nand U16964 (N_16964,N_12732,N_14039);
nand U16965 (N_16965,N_10000,N_14698);
or U16966 (N_16966,N_14483,N_10727);
nand U16967 (N_16967,N_13447,N_12378);
or U16968 (N_16968,N_10626,N_11563);
or U16969 (N_16969,N_14077,N_14994);
nor U16970 (N_16970,N_12891,N_13934);
nand U16971 (N_16971,N_13599,N_10294);
and U16972 (N_16972,N_12124,N_13845);
or U16973 (N_16973,N_11556,N_12592);
and U16974 (N_16974,N_12091,N_13579);
and U16975 (N_16975,N_13209,N_14814);
nor U16976 (N_16976,N_12729,N_12413);
nor U16977 (N_16977,N_14618,N_12299);
and U16978 (N_16978,N_10077,N_13188);
and U16979 (N_16979,N_13950,N_13566);
or U16980 (N_16980,N_10900,N_10223);
or U16981 (N_16981,N_14409,N_12630);
nand U16982 (N_16982,N_10206,N_13319);
or U16983 (N_16983,N_13076,N_12901);
or U16984 (N_16984,N_13954,N_14254);
nor U16985 (N_16985,N_14928,N_13062);
nor U16986 (N_16986,N_14178,N_10197);
and U16987 (N_16987,N_14962,N_12605);
or U16988 (N_16988,N_11375,N_12461);
or U16989 (N_16989,N_13425,N_11900);
nand U16990 (N_16990,N_12416,N_14579);
xor U16991 (N_16991,N_11261,N_14343);
nand U16992 (N_16992,N_14413,N_13065);
or U16993 (N_16993,N_11151,N_10026);
and U16994 (N_16994,N_13346,N_12281);
and U16995 (N_16995,N_12940,N_14883);
nand U16996 (N_16996,N_10640,N_14494);
nor U16997 (N_16997,N_14074,N_14627);
or U16998 (N_16998,N_14683,N_10132);
nor U16999 (N_16999,N_14591,N_11890);
or U17000 (N_17000,N_13652,N_14969);
or U17001 (N_17001,N_14480,N_13878);
and U17002 (N_17002,N_11353,N_13926);
and U17003 (N_17003,N_10302,N_10323);
and U17004 (N_17004,N_14617,N_10349);
or U17005 (N_17005,N_12699,N_10552);
nor U17006 (N_17006,N_14182,N_12014);
nor U17007 (N_17007,N_12469,N_14459);
or U17008 (N_17008,N_14326,N_10676);
and U17009 (N_17009,N_14429,N_11459);
and U17010 (N_17010,N_11308,N_14065);
and U17011 (N_17011,N_11265,N_10014);
or U17012 (N_17012,N_14586,N_10995);
or U17013 (N_17013,N_13669,N_12223);
nand U17014 (N_17014,N_10126,N_11854);
nor U17015 (N_17015,N_10953,N_12526);
or U17016 (N_17016,N_13371,N_14551);
and U17017 (N_17017,N_10463,N_13365);
and U17018 (N_17018,N_14156,N_14862);
or U17019 (N_17019,N_12992,N_12674);
or U17020 (N_17020,N_13288,N_11035);
or U17021 (N_17021,N_14768,N_13649);
nor U17022 (N_17022,N_12326,N_12611);
and U17023 (N_17023,N_14121,N_14796);
and U17024 (N_17024,N_12594,N_13913);
nor U17025 (N_17025,N_11048,N_10208);
or U17026 (N_17026,N_12133,N_13325);
and U17027 (N_17027,N_14758,N_13840);
nor U17028 (N_17028,N_12034,N_14829);
nor U17029 (N_17029,N_13958,N_13901);
and U17030 (N_17030,N_11646,N_13262);
nand U17031 (N_17031,N_10701,N_12304);
nor U17032 (N_17032,N_10941,N_12052);
or U17033 (N_17033,N_10160,N_12665);
or U17034 (N_17034,N_11478,N_11158);
or U17035 (N_17035,N_11014,N_14526);
and U17036 (N_17036,N_14038,N_14798);
nand U17037 (N_17037,N_10321,N_13734);
nor U17038 (N_17038,N_13301,N_14996);
nor U17039 (N_17039,N_11360,N_13920);
nand U17040 (N_17040,N_10639,N_14788);
nor U17041 (N_17041,N_11215,N_10163);
or U17042 (N_17042,N_10920,N_11339);
and U17043 (N_17043,N_10905,N_11083);
nand U17044 (N_17044,N_13937,N_10567);
nand U17045 (N_17045,N_12183,N_13804);
xnor U17046 (N_17046,N_13895,N_11961);
nand U17047 (N_17047,N_11654,N_10725);
nand U17048 (N_17048,N_11769,N_14516);
or U17049 (N_17049,N_13284,N_10483);
nand U17050 (N_17050,N_13395,N_12993);
and U17051 (N_17051,N_10986,N_11157);
nand U17052 (N_17052,N_13222,N_10684);
nor U17053 (N_17053,N_14771,N_11291);
nor U17054 (N_17054,N_11055,N_12409);
or U17055 (N_17055,N_12641,N_14096);
nand U17056 (N_17056,N_14610,N_14700);
nand U17057 (N_17057,N_10780,N_13977);
or U17058 (N_17058,N_12748,N_13134);
nor U17059 (N_17059,N_14442,N_10596);
or U17060 (N_17060,N_13340,N_13771);
nand U17061 (N_17061,N_13505,N_12550);
and U17062 (N_17062,N_14963,N_11039);
and U17063 (N_17063,N_14399,N_10991);
or U17064 (N_17064,N_11235,N_13216);
nor U17065 (N_17065,N_13009,N_11117);
nand U17066 (N_17066,N_11618,N_13513);
or U17067 (N_17067,N_11080,N_12206);
and U17068 (N_17068,N_14148,N_11970);
and U17069 (N_17069,N_10591,N_11306);
or U17070 (N_17070,N_12688,N_11712);
nand U17071 (N_17071,N_14933,N_14270);
nor U17072 (N_17072,N_11279,N_12292);
and U17073 (N_17073,N_12718,N_14067);
nand U17074 (N_17074,N_13331,N_13019);
or U17075 (N_17075,N_11673,N_13847);
nand U17076 (N_17076,N_14831,N_10688);
or U17077 (N_17077,N_10524,N_13698);
nand U17078 (N_17078,N_12180,N_11574);
nor U17079 (N_17079,N_11110,N_10329);
nor U17080 (N_17080,N_14290,N_14649);
nand U17081 (N_17081,N_12155,N_10434);
nand U17082 (N_17082,N_11450,N_12256);
and U17083 (N_17083,N_11228,N_14544);
or U17084 (N_17084,N_12166,N_12123);
or U17085 (N_17085,N_10038,N_14513);
nor U17086 (N_17086,N_11145,N_11609);
or U17087 (N_17087,N_12061,N_13286);
nand U17088 (N_17088,N_14676,N_11329);
or U17089 (N_17089,N_14584,N_14659);
or U17090 (N_17090,N_12260,N_10377);
nand U17091 (N_17091,N_14668,N_10794);
or U17092 (N_17092,N_13718,N_10710);
and U17093 (N_17093,N_13236,N_10692);
or U17094 (N_17094,N_14985,N_10958);
nand U17095 (N_17095,N_10595,N_11777);
and U17096 (N_17096,N_10482,N_12369);
and U17097 (N_17097,N_12776,N_13086);
or U17098 (N_17098,N_13525,N_10141);
nand U17099 (N_17099,N_11795,N_13449);
nand U17100 (N_17100,N_11280,N_11960);
nand U17101 (N_17101,N_10787,N_12511);
nand U17102 (N_17102,N_12012,N_10490);
nor U17103 (N_17103,N_11579,N_13562);
or U17104 (N_17104,N_11647,N_12514);
nand U17105 (N_17105,N_12591,N_11385);
nor U17106 (N_17106,N_10724,N_11324);
nor U17107 (N_17107,N_12802,N_11233);
nor U17108 (N_17108,N_11953,N_10352);
nand U17109 (N_17109,N_12831,N_11059);
and U17110 (N_17110,N_10074,N_10972);
nor U17111 (N_17111,N_12282,N_14900);
or U17112 (N_17112,N_14939,N_10511);
nor U17113 (N_17113,N_10268,N_12596);
nand U17114 (N_17114,N_12414,N_13900);
nand U17115 (N_17115,N_10303,N_12865);
nor U17116 (N_17116,N_12676,N_10347);
nor U17117 (N_17117,N_12241,N_12640);
nor U17118 (N_17118,N_10609,N_13563);
nand U17119 (N_17119,N_12417,N_13254);
nand U17120 (N_17120,N_12268,N_14232);
nor U17121 (N_17121,N_10426,N_14087);
nor U17122 (N_17122,N_10680,N_11736);
and U17123 (N_17123,N_12434,N_12215);
or U17124 (N_17124,N_12080,N_14089);
nand U17125 (N_17125,N_12768,N_14173);
or U17126 (N_17126,N_12695,N_13409);
nor U17127 (N_17127,N_14709,N_13650);
or U17128 (N_17128,N_11348,N_10942);
nor U17129 (N_17129,N_12746,N_10040);
or U17130 (N_17130,N_11969,N_10068);
or U17131 (N_17131,N_13618,N_10348);
or U17132 (N_17132,N_10702,N_13121);
and U17133 (N_17133,N_11126,N_14110);
and U17134 (N_17134,N_13741,N_12690);
or U17135 (N_17135,N_13413,N_12246);
or U17136 (N_17136,N_13300,N_12988);
or U17137 (N_17137,N_10785,N_10961);
and U17138 (N_17138,N_10593,N_11155);
nand U17139 (N_17139,N_12151,N_14675);
and U17140 (N_17140,N_10279,N_10419);
or U17141 (N_17141,N_12835,N_10355);
nand U17142 (N_17142,N_14265,N_11234);
nor U17143 (N_17143,N_10078,N_13989);
or U17144 (N_17144,N_13283,N_14082);
nor U17145 (N_17145,N_14753,N_12691);
or U17146 (N_17146,N_10696,N_14471);
nor U17147 (N_17147,N_14207,N_14559);
or U17148 (N_17148,N_13439,N_13038);
nor U17149 (N_17149,N_13059,N_10023);
and U17150 (N_17150,N_10471,N_11241);
or U17151 (N_17151,N_11141,N_11268);
nor U17152 (N_17152,N_11186,N_11987);
or U17153 (N_17153,N_11633,N_12635);
and U17154 (N_17154,N_12985,N_12798);
and U17155 (N_17155,N_11281,N_11132);
and U17156 (N_17156,N_12308,N_10022);
or U17157 (N_17157,N_12792,N_11939);
or U17158 (N_17158,N_14215,N_11680);
or U17159 (N_17159,N_11697,N_13568);
nand U17160 (N_17160,N_10213,N_13620);
or U17161 (N_17161,N_10088,N_11904);
and U17162 (N_17162,N_14841,N_11797);
nand U17163 (N_17163,N_11441,N_10983);
nor U17164 (N_17164,N_10599,N_13320);
or U17165 (N_17165,N_12287,N_13326);
nor U17166 (N_17166,N_14492,N_10547);
nand U17167 (N_17167,N_10935,N_10112);
and U17168 (N_17168,N_12478,N_13774);
and U17169 (N_17169,N_13498,N_10371);
and U17170 (N_17170,N_13666,N_11950);
nor U17171 (N_17171,N_13129,N_13496);
nor U17172 (N_17172,N_10544,N_13984);
nor U17173 (N_17173,N_13317,N_13410);
and U17174 (N_17174,N_12643,N_11922);
and U17175 (N_17175,N_12639,N_12785);
and U17176 (N_17176,N_14960,N_10439);
nor U17177 (N_17177,N_12535,N_11959);
nand U17178 (N_17178,N_11885,N_11415);
nand U17179 (N_17179,N_12418,N_10560);
nand U17180 (N_17180,N_13722,N_10478);
nand U17181 (N_17181,N_13234,N_13014);
and U17182 (N_17182,N_10036,N_14035);
or U17183 (N_17183,N_12472,N_12861);
nor U17184 (N_17184,N_12745,N_11175);
and U17185 (N_17185,N_12603,N_14395);
and U17186 (N_17186,N_14935,N_13710);
nand U17187 (N_17187,N_12364,N_10615);
nor U17188 (N_17188,N_12010,N_14348);
nor U17189 (N_17189,N_10071,N_10176);
nor U17190 (N_17190,N_14968,N_14999);
nand U17191 (N_17191,N_14520,N_12825);
and U17192 (N_17192,N_14919,N_10823);
or U17193 (N_17193,N_11290,N_13499);
nor U17194 (N_17194,N_11860,N_14443);
nand U17195 (N_17195,N_13556,N_13472);
nor U17196 (N_17196,N_10581,N_14736);
nor U17197 (N_17197,N_11985,N_12411);
or U17198 (N_17198,N_14823,N_11764);
nand U17199 (N_17199,N_14009,N_11943);
and U17200 (N_17200,N_12235,N_12298);
nand U17201 (N_17201,N_11311,N_13324);
and U17202 (N_17202,N_12795,N_11168);
or U17203 (N_17203,N_10602,N_12646);
xnor U17204 (N_17204,N_10476,N_12553);
nor U17205 (N_17205,N_14341,N_14319);
nor U17206 (N_17206,N_11485,N_11187);
or U17207 (N_17207,N_14652,N_10770);
nor U17208 (N_17208,N_11868,N_14854);
and U17209 (N_17209,N_10136,N_11103);
xnor U17210 (N_17210,N_10369,N_14320);
nand U17211 (N_17211,N_14163,N_14539);
nand U17212 (N_17212,N_11717,N_14095);
nand U17213 (N_17213,N_14432,N_11933);
and U17214 (N_17214,N_10833,N_13189);
and U17215 (N_17215,N_10236,N_13623);
or U17216 (N_17216,N_12522,N_13644);
or U17217 (N_17217,N_11617,N_12853);
or U17218 (N_17218,N_10039,N_13420);
nand U17219 (N_17219,N_14974,N_14921);
and U17220 (N_17220,N_13688,N_14190);
nand U17221 (N_17221,N_11469,N_14229);
nand U17222 (N_17222,N_10494,N_14137);
or U17223 (N_17223,N_13108,N_12787);
nand U17224 (N_17224,N_11447,N_10634);
and U17225 (N_17225,N_12766,N_10423);
and U17226 (N_17226,N_14441,N_13487);
and U17227 (N_17227,N_12149,N_14340);
and U17228 (N_17228,N_10711,N_14599);
and U17229 (N_17229,N_11153,N_14785);
nor U17230 (N_17230,N_12937,N_14552);
and U17231 (N_17231,N_10650,N_13651);
or U17232 (N_17232,N_14461,N_11122);
nor U17233 (N_17233,N_12044,N_13864);
nand U17234 (N_17234,N_14015,N_11425);
nor U17235 (N_17235,N_13897,N_10992);
or U17236 (N_17236,N_10510,N_11632);
and U17237 (N_17237,N_13355,N_14079);
and U17238 (N_17238,N_13143,N_14863);
or U17239 (N_17239,N_11714,N_13802);
nand U17240 (N_17240,N_12667,N_10148);
or U17241 (N_17241,N_14143,N_13459);
nand U17242 (N_17242,N_13255,N_12570);
or U17243 (N_17243,N_13871,N_10309);
or U17244 (N_17244,N_10922,N_10660);
or U17245 (N_17245,N_12213,N_14214);
or U17246 (N_17246,N_13793,N_12031);
nor U17247 (N_17247,N_12333,N_11739);
and U17248 (N_17248,N_13294,N_11744);
xor U17249 (N_17249,N_13165,N_11171);
nor U17250 (N_17250,N_11884,N_14278);
nor U17251 (N_17251,N_11002,N_11899);
or U17252 (N_17252,N_10414,N_13070);
nand U17253 (N_17253,N_12628,N_13524);
nor U17254 (N_17254,N_12309,N_13854);
or U17255 (N_17255,N_12812,N_13851);
nor U17256 (N_17256,N_10746,N_12767);
and U17257 (N_17257,N_10313,N_11481);
nand U17258 (N_17258,N_11641,N_11222);
or U17259 (N_17259,N_13982,N_12191);
nand U17260 (N_17260,N_13915,N_12862);
or U17261 (N_17261,N_14292,N_12722);
nand U17262 (N_17262,N_11046,N_12551);
nand U17263 (N_17263,N_14797,N_12410);
nor U17264 (N_17264,N_14068,N_11154);
xor U17265 (N_17265,N_13885,N_12964);
and U17266 (N_17266,N_12391,N_14765);
nor U17267 (N_17267,N_10297,N_12087);
and U17268 (N_17268,N_14761,N_10218);
and U17269 (N_17269,N_14238,N_12951);
and U17270 (N_17270,N_10418,N_12224);
or U17271 (N_17271,N_10975,N_13988);
or U17272 (N_17272,N_13572,N_11931);
or U17273 (N_17273,N_11043,N_10849);
and U17274 (N_17274,N_11095,N_12969);
or U17275 (N_17275,N_13687,N_12093);
and U17276 (N_17276,N_13349,N_13981);
nand U17277 (N_17277,N_12153,N_12444);
nand U17278 (N_17278,N_12589,N_13055);
nor U17279 (N_17279,N_12234,N_14410);
or U17280 (N_17280,N_13240,N_11909);
or U17281 (N_17281,N_11766,N_14330);
nor U17282 (N_17282,N_14800,N_12272);
nand U17283 (N_17283,N_12632,N_14906);
nor U17284 (N_17284,N_10257,N_11012);
nand U17285 (N_17285,N_11830,N_10817);
xnor U17286 (N_17286,N_14653,N_12201);
or U17287 (N_17287,N_10210,N_13943);
and U17288 (N_17288,N_10027,N_10967);
nor U17289 (N_17289,N_11042,N_13315);
and U17290 (N_17290,N_12039,N_10543);
nor U17291 (N_17291,N_12618,N_13271);
or U17292 (N_17292,N_14642,N_10401);
or U17293 (N_17293,N_11350,N_14041);
nor U17294 (N_17294,N_14625,N_11841);
nand U17295 (N_17295,N_12683,N_13996);
nor U17296 (N_17296,N_12752,N_14973);
nand U17297 (N_17297,N_11687,N_12657);
and U17298 (N_17298,N_14949,N_11525);
nand U17299 (N_17299,N_14720,N_13314);
or U17300 (N_17300,N_13675,N_12353);
or U17301 (N_17301,N_13674,N_12145);
or U17302 (N_17302,N_12138,N_10999);
nand U17303 (N_17303,N_11406,N_14303);
nand U17304 (N_17304,N_10594,N_14965);
nand U17305 (N_17305,N_13136,N_12749);
or U17306 (N_17306,N_11445,N_13166);
nor U17307 (N_17307,N_12500,N_11923);
and U17308 (N_17308,N_10072,N_10481);
or U17309 (N_17309,N_12850,N_10273);
nor U17310 (N_17310,N_10568,N_13031);
nor U17311 (N_17311,N_10777,N_14681);
nand U17312 (N_17312,N_11669,N_13916);
and U17313 (N_17313,N_10200,N_12311);
nand U17314 (N_17314,N_12421,N_10091);
and U17315 (N_17315,N_13985,N_11754);
nand U17316 (N_17316,N_12325,N_10378);
and U17317 (N_17317,N_11555,N_13453);
nand U17318 (N_17318,N_14592,N_10135);
nand U17319 (N_17319,N_13759,N_14993);
nor U17320 (N_17320,N_12573,N_13707);
or U17321 (N_17321,N_12942,N_12877);
nor U17322 (N_17322,N_14885,N_10630);
or U17323 (N_17323,N_13084,N_11536);
nor U17324 (N_17324,N_10252,N_11414);
and U17325 (N_17325,N_13156,N_12938);
nand U17326 (N_17326,N_13746,N_12203);
nor U17327 (N_17327,N_11325,N_10037);
or U17328 (N_17328,N_11470,N_13266);
or U17329 (N_17329,N_14372,N_12095);
and U17330 (N_17330,N_12979,N_14790);
or U17331 (N_17331,N_10170,N_11248);
nor U17332 (N_17332,N_13670,N_10466);
and U17333 (N_17333,N_11230,N_14719);
nor U17334 (N_17334,N_12435,N_10234);
nand U17335 (N_17335,N_14361,N_10617);
and U17336 (N_17336,N_12271,N_12914);
nand U17337 (N_17337,N_13509,N_11530);
or U17338 (N_17338,N_13708,N_14608);
nand U17339 (N_17339,N_12345,N_11504);
nor U17340 (N_17340,N_11857,N_12929);
or U17341 (N_17341,N_14821,N_12892);
or U17342 (N_17342,N_14021,N_10376);
nand U17343 (N_17343,N_13658,N_13028);
and U17344 (N_17344,N_14052,N_14165);
and U17345 (N_17345,N_10842,N_12501);
nand U17346 (N_17346,N_11247,N_14878);
or U17347 (N_17347,N_12503,N_10199);
nand U17348 (N_17348,N_12614,N_10123);
or U17349 (N_17349,N_14037,N_11200);
nand U17350 (N_17350,N_10624,N_12179);
or U17351 (N_17351,N_13994,N_12425);
nand U17352 (N_17352,N_13282,N_14286);
nor U17353 (N_17353,N_12606,N_11125);
and U17354 (N_17354,N_12998,N_14825);
or U17355 (N_17355,N_10097,N_12362);
nor U17356 (N_17356,N_14886,N_11752);
and U17357 (N_17357,N_10403,N_14762);
nor U17358 (N_17358,N_12077,N_12066);
nand U17359 (N_17359,N_14612,N_14803);
and U17360 (N_17360,N_11926,N_10878);
nor U17361 (N_17361,N_11835,N_10336);
and U17362 (N_17362,N_14772,N_11197);
or U17363 (N_17363,N_10621,N_13212);
nor U17364 (N_17364,N_12593,N_12396);
and U17365 (N_17365,N_12737,N_10733);
or U17366 (N_17366,N_12943,N_14097);
nand U17367 (N_17367,N_10644,N_11351);
nand U17368 (N_17368,N_14365,N_10165);
and U17369 (N_17369,N_10553,N_14899);
nand U17370 (N_17370,N_10283,N_13838);
or U17371 (N_17371,N_13109,N_13256);
nand U17372 (N_17372,N_14018,N_14650);
nand U17373 (N_17373,N_14475,N_13366);
and U17374 (N_17374,N_10043,N_14576);
nor U17375 (N_17375,N_11287,N_10105);
and U17376 (N_17376,N_12393,N_12327);
nand U17377 (N_17377,N_11786,N_14368);
and U17378 (N_17378,N_14582,N_12740);
or U17379 (N_17379,N_11320,N_13866);
or U17380 (N_17380,N_12713,N_14619);
nand U17381 (N_17381,N_14860,N_12709);
nand U17382 (N_17382,N_13909,N_12772);
or U17383 (N_17383,N_13224,N_11575);
nor U17384 (N_17384,N_13443,N_13401);
nor U17385 (N_17385,N_13464,N_10411);
and U17386 (N_17386,N_12468,N_11121);
and U17387 (N_17387,N_10157,N_13250);
and U17388 (N_17388,N_12321,N_10100);
nor U17389 (N_17389,N_12154,N_10306);
or U17390 (N_17390,N_13379,N_12341);
nand U17391 (N_17391,N_14696,N_12289);
nand U17392 (N_17392,N_12453,N_10818);
nand U17393 (N_17393,N_11422,N_11246);
or U17394 (N_17394,N_14063,N_12236);
and U17395 (N_17395,N_12733,N_11746);
nand U17396 (N_17396,N_10247,N_10830);
and U17397 (N_17397,N_12380,N_11527);
nor U17398 (N_17398,N_14157,N_12720);
nor U17399 (N_17399,N_11189,N_11458);
nor U17400 (N_17400,N_14093,N_14658);
and U17401 (N_17401,N_14397,N_11314);
or U17402 (N_17402,N_13103,N_13238);
and U17403 (N_17403,N_13631,N_12890);
nor U17404 (N_17404,N_14705,N_11696);
nand U17405 (N_17405,N_12379,N_14647);
and U17406 (N_17406,N_10788,N_13991);
nand U17407 (N_17407,N_14713,N_10583);
and U17408 (N_17408,N_11352,N_11843);
or U17409 (N_17409,N_14573,N_12567);
or U17410 (N_17410,N_11313,N_13603);
and U17411 (N_17411,N_14381,N_11092);
nand U17412 (N_17412,N_13394,N_13656);
nor U17413 (N_17413,N_11827,N_10751);
nand U17414 (N_17414,N_12217,N_11148);
nand U17415 (N_17415,N_14743,N_10648);
nand U17416 (N_17416,N_11541,N_10705);
and U17417 (N_17417,N_10667,N_10656);
nand U17418 (N_17418,N_12751,N_11751);
nor U17419 (N_17419,N_13608,N_10870);
nor U17420 (N_17420,N_14452,N_10737);
nand U17421 (N_17421,N_14563,N_13244);
or U17422 (N_17422,N_11322,N_14026);
nor U17423 (N_17423,N_12875,N_11787);
or U17424 (N_17424,N_14123,N_13660);
nor U17425 (N_17425,N_10545,N_10122);
and U17426 (N_17426,N_12076,N_14995);
or U17427 (N_17427,N_14637,N_13131);
nor U17428 (N_17428,N_10340,N_12471);
nand U17429 (N_17429,N_14000,N_10169);
and U17430 (N_17430,N_12384,N_10844);
nor U17431 (N_17431,N_14914,N_14631);
nand U17432 (N_17432,N_10318,N_11381);
nand U17433 (N_17433,N_14204,N_10269);
nor U17434 (N_17434,N_11142,N_11630);
nor U17435 (N_17435,N_12389,N_11299);
or U17436 (N_17436,N_11983,N_11965);
nor U17437 (N_17437,N_14205,N_11516);
nor U17438 (N_17438,N_10087,N_14881);
nor U17439 (N_17439,N_14726,N_11271);
nor U17440 (N_17440,N_11294,N_11614);
nand U17441 (N_17441,N_13170,N_14457);
and U17442 (N_17442,N_14268,N_14953);
and U17443 (N_17443,N_12651,N_12332);
nor U17444 (N_17444,N_11493,N_14419);
nand U17445 (N_17445,N_11529,N_12701);
and U17446 (N_17446,N_13609,N_10677);
or U17447 (N_17447,N_10600,N_14628);
or U17448 (N_17448,N_12874,N_14464);
nor U17449 (N_17449,N_13116,N_11321);
or U17450 (N_17450,N_14490,N_10622);
or U17451 (N_17451,N_14033,N_11559);
nand U17452 (N_17452,N_12613,N_14345);
nand U17453 (N_17453,N_11160,N_13813);
nand U17454 (N_17454,N_13268,N_13276);
or U17455 (N_17455,N_14075,N_11273);
and U17456 (N_17456,N_14802,N_13822);
or U17457 (N_17457,N_13679,N_11651);
or U17458 (N_17458,N_14155,N_10569);
nor U17459 (N_17459,N_11512,N_10893);
nand U17460 (N_17460,N_12065,N_12033);
nor U17461 (N_17461,N_14482,N_14851);
or U17462 (N_17462,N_12997,N_14541);
or U17463 (N_17463,N_13457,N_12727);
and U17464 (N_17464,N_14824,N_11173);
or U17465 (N_17465,N_11139,N_12716);
nand U17466 (N_17466,N_13246,N_14398);
nand U17467 (N_17467,N_13327,N_13455);
and U17468 (N_17468,N_10212,N_14673);
nand U17469 (N_17469,N_10765,N_11326);
and U17470 (N_17470,N_10301,N_13438);
nor U17471 (N_17471,N_14897,N_11742);
nand U17472 (N_17472,N_10632,N_14369);
xor U17473 (N_17473,N_14493,N_12250);
and U17474 (N_17474,N_12313,N_11692);
nand U17475 (N_17475,N_14868,N_13872);
and U17476 (N_17476,N_10131,N_13615);
or U17477 (N_17477,N_11489,N_11774);
or U17478 (N_17478,N_10314,N_13665);
and U17479 (N_17479,N_13334,N_11865);
nand U17480 (N_17480,N_11785,N_14007);
or U17481 (N_17481,N_12539,N_11813);
or U17482 (N_17482,N_13949,N_14098);
nor U17483 (N_17483,N_11309,N_10509);
and U17484 (N_17484,N_12159,N_13944);
and U17485 (N_17485,N_10030,N_12238);
nor U17486 (N_17486,N_12847,N_11475);
nand U17487 (N_17487,N_12148,N_11539);
or U17488 (N_17488,N_13113,N_10417);
nand U17489 (N_17489,N_11544,N_12082);
or U17490 (N_17490,N_14727,N_12090);
or U17491 (N_17491,N_12715,N_10217);
or U17492 (N_17492,N_12811,N_13274);
and U17493 (N_17493,N_11453,N_11927);
nand U17494 (N_17494,N_14777,N_14364);
or U17495 (N_17495,N_13161,N_10255);
nand U17496 (N_17496,N_11210,N_14408);
or U17497 (N_17497,N_13408,N_12479);
and U17498 (N_17498,N_13783,N_11963);
nand U17499 (N_17499,N_10962,N_10057);
nand U17500 (N_17500,N_12009,N_11544);
or U17501 (N_17501,N_14800,N_13754);
nor U17502 (N_17502,N_14897,N_10950);
nor U17503 (N_17503,N_14075,N_12754);
nand U17504 (N_17504,N_10602,N_13842);
nor U17505 (N_17505,N_10142,N_10309);
nand U17506 (N_17506,N_11732,N_10633);
nand U17507 (N_17507,N_11568,N_10261);
nor U17508 (N_17508,N_12925,N_13202);
or U17509 (N_17509,N_12562,N_10187);
and U17510 (N_17510,N_14116,N_14084);
nor U17511 (N_17511,N_10733,N_11105);
and U17512 (N_17512,N_13713,N_10744);
nand U17513 (N_17513,N_12279,N_13267);
or U17514 (N_17514,N_13438,N_13674);
or U17515 (N_17515,N_10708,N_12052);
or U17516 (N_17516,N_14227,N_10128);
and U17517 (N_17517,N_13208,N_12318);
and U17518 (N_17518,N_12468,N_11363);
and U17519 (N_17519,N_12993,N_14612);
and U17520 (N_17520,N_13369,N_14534);
nand U17521 (N_17521,N_12112,N_11520);
or U17522 (N_17522,N_13466,N_12994);
nor U17523 (N_17523,N_10150,N_10726);
nand U17524 (N_17524,N_14363,N_11595);
nor U17525 (N_17525,N_12391,N_13807);
nor U17526 (N_17526,N_11655,N_11331);
nor U17527 (N_17527,N_13800,N_10909);
nor U17528 (N_17528,N_14115,N_14973);
nand U17529 (N_17529,N_14894,N_14191);
nand U17530 (N_17530,N_14262,N_14945);
nor U17531 (N_17531,N_11571,N_12750);
nor U17532 (N_17532,N_10304,N_11436);
nor U17533 (N_17533,N_10630,N_10683);
nor U17534 (N_17534,N_12745,N_11704);
or U17535 (N_17535,N_10219,N_13317);
nor U17536 (N_17536,N_12775,N_12645);
nor U17537 (N_17537,N_14923,N_11399);
nor U17538 (N_17538,N_13641,N_11564);
or U17539 (N_17539,N_12564,N_14335);
nand U17540 (N_17540,N_10637,N_11985);
and U17541 (N_17541,N_13415,N_11452);
nand U17542 (N_17542,N_11533,N_12962);
nand U17543 (N_17543,N_10618,N_14724);
and U17544 (N_17544,N_13372,N_14809);
or U17545 (N_17545,N_12652,N_11254);
nand U17546 (N_17546,N_11879,N_14659);
or U17547 (N_17547,N_12125,N_14792);
nor U17548 (N_17548,N_13305,N_12465);
and U17549 (N_17549,N_12632,N_13543);
nor U17550 (N_17550,N_10237,N_10303);
or U17551 (N_17551,N_10797,N_12870);
and U17552 (N_17552,N_10389,N_11073);
or U17553 (N_17553,N_10403,N_10516);
and U17554 (N_17554,N_13468,N_11297);
and U17555 (N_17555,N_11341,N_11065);
nor U17556 (N_17556,N_12087,N_13614);
nand U17557 (N_17557,N_13952,N_10692);
nand U17558 (N_17558,N_12529,N_10821);
nor U17559 (N_17559,N_12539,N_14322);
and U17560 (N_17560,N_14842,N_14123);
and U17561 (N_17561,N_14169,N_12954);
or U17562 (N_17562,N_12617,N_13453);
or U17563 (N_17563,N_14411,N_10083);
nor U17564 (N_17564,N_10454,N_13400);
nor U17565 (N_17565,N_11807,N_12849);
nor U17566 (N_17566,N_11328,N_11217);
or U17567 (N_17567,N_14310,N_10857);
nor U17568 (N_17568,N_14879,N_14559);
or U17569 (N_17569,N_13890,N_13512);
or U17570 (N_17570,N_14279,N_11781);
nand U17571 (N_17571,N_10653,N_12078);
and U17572 (N_17572,N_12871,N_12136);
nor U17573 (N_17573,N_12516,N_11269);
or U17574 (N_17574,N_10326,N_12244);
and U17575 (N_17575,N_13750,N_13019);
and U17576 (N_17576,N_10025,N_12140);
and U17577 (N_17577,N_14203,N_10114);
or U17578 (N_17578,N_11513,N_14712);
nor U17579 (N_17579,N_12198,N_13153);
or U17580 (N_17580,N_11999,N_14013);
and U17581 (N_17581,N_10881,N_13861);
and U17582 (N_17582,N_13279,N_13415);
and U17583 (N_17583,N_10075,N_13113);
nand U17584 (N_17584,N_14464,N_12601);
or U17585 (N_17585,N_11822,N_12657);
nor U17586 (N_17586,N_11489,N_14710);
nor U17587 (N_17587,N_13471,N_13793);
nor U17588 (N_17588,N_12639,N_11098);
or U17589 (N_17589,N_14672,N_10973);
nor U17590 (N_17590,N_12749,N_14352);
nand U17591 (N_17591,N_11200,N_14297);
nor U17592 (N_17592,N_10558,N_11004);
nand U17593 (N_17593,N_13143,N_14960);
xnor U17594 (N_17594,N_13872,N_12439);
nand U17595 (N_17595,N_10776,N_14203);
and U17596 (N_17596,N_12584,N_10882);
or U17597 (N_17597,N_13722,N_14063);
and U17598 (N_17598,N_13053,N_11926);
nand U17599 (N_17599,N_14022,N_14528);
and U17600 (N_17600,N_14578,N_12566);
nor U17601 (N_17601,N_12085,N_11337);
nand U17602 (N_17602,N_13257,N_13116);
or U17603 (N_17603,N_12168,N_10342);
and U17604 (N_17604,N_14724,N_12479);
or U17605 (N_17605,N_10821,N_12568);
nor U17606 (N_17606,N_11356,N_13807);
nand U17607 (N_17607,N_13249,N_11929);
and U17608 (N_17608,N_13534,N_14120);
nor U17609 (N_17609,N_13940,N_11796);
or U17610 (N_17610,N_11663,N_12882);
or U17611 (N_17611,N_13383,N_12355);
or U17612 (N_17612,N_10897,N_10574);
nand U17613 (N_17613,N_12101,N_13886);
nor U17614 (N_17614,N_10071,N_12982);
nor U17615 (N_17615,N_14766,N_13602);
and U17616 (N_17616,N_11073,N_10009);
xnor U17617 (N_17617,N_12423,N_13042);
or U17618 (N_17618,N_12464,N_13644);
and U17619 (N_17619,N_14593,N_10293);
nand U17620 (N_17620,N_12946,N_13496);
or U17621 (N_17621,N_10309,N_14453);
nor U17622 (N_17622,N_14207,N_11489);
or U17623 (N_17623,N_14686,N_11868);
and U17624 (N_17624,N_14863,N_10165);
nand U17625 (N_17625,N_13899,N_11378);
and U17626 (N_17626,N_11294,N_10124);
and U17627 (N_17627,N_14321,N_12349);
nor U17628 (N_17628,N_12785,N_14673);
and U17629 (N_17629,N_14286,N_13023);
nor U17630 (N_17630,N_11323,N_10075);
and U17631 (N_17631,N_10515,N_10355);
and U17632 (N_17632,N_12163,N_11957);
nand U17633 (N_17633,N_11970,N_12412);
nor U17634 (N_17634,N_14718,N_10692);
and U17635 (N_17635,N_14163,N_11328);
and U17636 (N_17636,N_12663,N_10549);
nand U17637 (N_17637,N_11309,N_10500);
and U17638 (N_17638,N_14910,N_12786);
nand U17639 (N_17639,N_13910,N_10799);
and U17640 (N_17640,N_13741,N_13823);
or U17641 (N_17641,N_13378,N_13878);
nand U17642 (N_17642,N_13720,N_10419);
nor U17643 (N_17643,N_11493,N_10001);
and U17644 (N_17644,N_10865,N_12790);
or U17645 (N_17645,N_11310,N_10646);
and U17646 (N_17646,N_11262,N_12945);
nand U17647 (N_17647,N_13872,N_14559);
or U17648 (N_17648,N_11469,N_10920);
xor U17649 (N_17649,N_11996,N_11022);
nand U17650 (N_17650,N_13150,N_12957);
nor U17651 (N_17651,N_12875,N_11087);
or U17652 (N_17652,N_14420,N_14473);
and U17653 (N_17653,N_13619,N_10838);
and U17654 (N_17654,N_13369,N_14287);
nor U17655 (N_17655,N_13415,N_12617);
and U17656 (N_17656,N_10668,N_11890);
nand U17657 (N_17657,N_13661,N_10780);
and U17658 (N_17658,N_14083,N_11274);
nand U17659 (N_17659,N_14961,N_13732);
nor U17660 (N_17660,N_10653,N_13314);
or U17661 (N_17661,N_12257,N_10563);
xnor U17662 (N_17662,N_12784,N_11120);
and U17663 (N_17663,N_12456,N_14432);
nand U17664 (N_17664,N_12143,N_14358);
or U17665 (N_17665,N_13451,N_10303);
nor U17666 (N_17666,N_11193,N_12489);
or U17667 (N_17667,N_10597,N_10425);
and U17668 (N_17668,N_10052,N_12688);
nor U17669 (N_17669,N_10102,N_13049);
nor U17670 (N_17670,N_11429,N_13324);
nor U17671 (N_17671,N_13106,N_10652);
nor U17672 (N_17672,N_10310,N_12249);
nor U17673 (N_17673,N_13066,N_14737);
or U17674 (N_17674,N_14481,N_14291);
or U17675 (N_17675,N_14403,N_10153);
and U17676 (N_17676,N_12560,N_11304);
and U17677 (N_17677,N_10682,N_13066);
nor U17678 (N_17678,N_13434,N_11815);
and U17679 (N_17679,N_13002,N_14841);
or U17680 (N_17680,N_10120,N_13312);
xor U17681 (N_17681,N_13673,N_11388);
and U17682 (N_17682,N_14857,N_12896);
nor U17683 (N_17683,N_11155,N_13585);
nor U17684 (N_17684,N_12546,N_10055);
nand U17685 (N_17685,N_10181,N_12055);
or U17686 (N_17686,N_11260,N_12587);
or U17687 (N_17687,N_14295,N_14559);
or U17688 (N_17688,N_12833,N_13847);
or U17689 (N_17689,N_10828,N_12366);
or U17690 (N_17690,N_12713,N_10295);
nor U17691 (N_17691,N_14804,N_12763);
nand U17692 (N_17692,N_13586,N_14390);
nand U17693 (N_17693,N_11118,N_12864);
nand U17694 (N_17694,N_13077,N_12548);
or U17695 (N_17695,N_12780,N_12774);
nor U17696 (N_17696,N_10153,N_14651);
and U17697 (N_17697,N_14150,N_14061);
and U17698 (N_17698,N_11516,N_11080);
and U17699 (N_17699,N_12484,N_10495);
or U17700 (N_17700,N_13135,N_10565);
or U17701 (N_17701,N_14341,N_14099);
and U17702 (N_17702,N_13589,N_13151);
or U17703 (N_17703,N_11582,N_11064);
nand U17704 (N_17704,N_12181,N_11346);
nand U17705 (N_17705,N_12791,N_10864);
nor U17706 (N_17706,N_11899,N_12207);
and U17707 (N_17707,N_10420,N_12017);
nand U17708 (N_17708,N_13717,N_12329);
nor U17709 (N_17709,N_11179,N_11580);
nand U17710 (N_17710,N_10960,N_11115);
nand U17711 (N_17711,N_11508,N_14658);
nor U17712 (N_17712,N_11725,N_11487);
nor U17713 (N_17713,N_12521,N_12461);
and U17714 (N_17714,N_13104,N_11585);
nor U17715 (N_17715,N_13106,N_12515);
nor U17716 (N_17716,N_10677,N_14594);
or U17717 (N_17717,N_11172,N_12661);
or U17718 (N_17718,N_10450,N_11371);
and U17719 (N_17719,N_11392,N_11062);
nand U17720 (N_17720,N_14240,N_14411);
or U17721 (N_17721,N_10452,N_14273);
nand U17722 (N_17722,N_14773,N_14734);
and U17723 (N_17723,N_14543,N_12311);
and U17724 (N_17724,N_12803,N_10589);
or U17725 (N_17725,N_14152,N_12633);
and U17726 (N_17726,N_13322,N_14183);
and U17727 (N_17727,N_14357,N_12766);
and U17728 (N_17728,N_10915,N_14010);
nor U17729 (N_17729,N_12915,N_11505);
or U17730 (N_17730,N_14665,N_10035);
or U17731 (N_17731,N_11626,N_11954);
and U17732 (N_17732,N_10845,N_14113);
and U17733 (N_17733,N_11595,N_12801);
and U17734 (N_17734,N_10424,N_13725);
nand U17735 (N_17735,N_10066,N_14595);
nand U17736 (N_17736,N_12828,N_14036);
nand U17737 (N_17737,N_11524,N_10409);
nor U17738 (N_17738,N_11369,N_14546);
or U17739 (N_17739,N_10857,N_13453);
nand U17740 (N_17740,N_11268,N_11799);
nor U17741 (N_17741,N_13915,N_13107);
nand U17742 (N_17742,N_10970,N_10158);
nor U17743 (N_17743,N_10728,N_11415);
or U17744 (N_17744,N_14512,N_11282);
or U17745 (N_17745,N_13780,N_14178);
nand U17746 (N_17746,N_14794,N_12216);
and U17747 (N_17747,N_10091,N_10394);
and U17748 (N_17748,N_11690,N_12242);
nor U17749 (N_17749,N_10736,N_10705);
nor U17750 (N_17750,N_13533,N_13707);
nor U17751 (N_17751,N_10877,N_14965);
and U17752 (N_17752,N_10715,N_10481);
and U17753 (N_17753,N_14191,N_10985);
or U17754 (N_17754,N_14494,N_11163);
and U17755 (N_17755,N_13235,N_10289);
nand U17756 (N_17756,N_14557,N_12975);
nand U17757 (N_17757,N_10984,N_14691);
and U17758 (N_17758,N_11073,N_11564);
nand U17759 (N_17759,N_13745,N_11421);
or U17760 (N_17760,N_13298,N_13242);
or U17761 (N_17761,N_14685,N_13759);
or U17762 (N_17762,N_12970,N_11690);
nor U17763 (N_17763,N_11420,N_12704);
and U17764 (N_17764,N_13788,N_11318);
nor U17765 (N_17765,N_10789,N_13337);
nor U17766 (N_17766,N_10177,N_12129);
nand U17767 (N_17767,N_11327,N_12885);
nor U17768 (N_17768,N_13842,N_14130);
or U17769 (N_17769,N_12259,N_12789);
and U17770 (N_17770,N_14670,N_10614);
nor U17771 (N_17771,N_11310,N_13927);
or U17772 (N_17772,N_12904,N_12440);
nand U17773 (N_17773,N_14845,N_11023);
nand U17774 (N_17774,N_10597,N_13153);
or U17775 (N_17775,N_11178,N_13049);
nor U17776 (N_17776,N_12022,N_14915);
nor U17777 (N_17777,N_10759,N_13975);
nor U17778 (N_17778,N_11162,N_11183);
and U17779 (N_17779,N_10743,N_14857);
nand U17780 (N_17780,N_11953,N_13052);
nor U17781 (N_17781,N_12695,N_14752);
and U17782 (N_17782,N_13333,N_11506);
and U17783 (N_17783,N_11706,N_13405);
and U17784 (N_17784,N_12620,N_13136);
nor U17785 (N_17785,N_12830,N_11108);
and U17786 (N_17786,N_11403,N_13369);
nor U17787 (N_17787,N_10225,N_13913);
or U17788 (N_17788,N_14770,N_12746);
nand U17789 (N_17789,N_12901,N_14907);
nand U17790 (N_17790,N_12946,N_13217);
and U17791 (N_17791,N_10810,N_13912);
nor U17792 (N_17792,N_13432,N_10519);
nand U17793 (N_17793,N_11112,N_13694);
nand U17794 (N_17794,N_11818,N_11358);
nor U17795 (N_17795,N_14897,N_14914);
nand U17796 (N_17796,N_10562,N_11358);
and U17797 (N_17797,N_12318,N_13126);
and U17798 (N_17798,N_13728,N_11559);
nor U17799 (N_17799,N_14349,N_11032);
nand U17800 (N_17800,N_13218,N_12384);
nor U17801 (N_17801,N_13349,N_12294);
nor U17802 (N_17802,N_14452,N_14865);
nor U17803 (N_17803,N_13478,N_14695);
or U17804 (N_17804,N_11241,N_13366);
nor U17805 (N_17805,N_12010,N_12966);
or U17806 (N_17806,N_10746,N_11880);
nor U17807 (N_17807,N_12870,N_12971);
and U17808 (N_17808,N_10454,N_10149);
and U17809 (N_17809,N_10164,N_13002);
nand U17810 (N_17810,N_11388,N_11902);
and U17811 (N_17811,N_12921,N_13638);
nor U17812 (N_17812,N_12738,N_11058);
and U17813 (N_17813,N_13664,N_13534);
nand U17814 (N_17814,N_12936,N_11356);
or U17815 (N_17815,N_10052,N_10589);
nand U17816 (N_17816,N_12112,N_13063);
and U17817 (N_17817,N_12699,N_10208);
and U17818 (N_17818,N_13468,N_10971);
or U17819 (N_17819,N_13047,N_12382);
or U17820 (N_17820,N_11719,N_13427);
nand U17821 (N_17821,N_13305,N_14477);
nor U17822 (N_17822,N_12030,N_13589);
or U17823 (N_17823,N_13554,N_13458);
nor U17824 (N_17824,N_12068,N_12062);
nor U17825 (N_17825,N_10822,N_13628);
nor U17826 (N_17826,N_13769,N_14322);
nand U17827 (N_17827,N_14500,N_14303);
nor U17828 (N_17828,N_14010,N_10802);
or U17829 (N_17829,N_10598,N_14039);
nand U17830 (N_17830,N_13169,N_13849);
and U17831 (N_17831,N_12524,N_14601);
and U17832 (N_17832,N_14535,N_12814);
nor U17833 (N_17833,N_11284,N_11148);
nor U17834 (N_17834,N_10136,N_10582);
nand U17835 (N_17835,N_14797,N_11862);
nor U17836 (N_17836,N_12465,N_12997);
and U17837 (N_17837,N_11795,N_13219);
nor U17838 (N_17838,N_11790,N_13347);
nand U17839 (N_17839,N_11303,N_12431);
and U17840 (N_17840,N_13302,N_12080);
nor U17841 (N_17841,N_11369,N_12355);
and U17842 (N_17842,N_14181,N_14793);
nor U17843 (N_17843,N_14848,N_14267);
nor U17844 (N_17844,N_13115,N_14689);
or U17845 (N_17845,N_14296,N_11391);
nor U17846 (N_17846,N_14983,N_12811);
and U17847 (N_17847,N_14027,N_11033);
or U17848 (N_17848,N_12496,N_13389);
nand U17849 (N_17849,N_13129,N_14607);
and U17850 (N_17850,N_11605,N_14730);
nand U17851 (N_17851,N_11997,N_14948);
nand U17852 (N_17852,N_12997,N_14507);
and U17853 (N_17853,N_12262,N_12677);
or U17854 (N_17854,N_10903,N_12450);
and U17855 (N_17855,N_14181,N_10707);
nor U17856 (N_17856,N_11642,N_12477);
or U17857 (N_17857,N_13687,N_11142);
nand U17858 (N_17858,N_12662,N_10490);
or U17859 (N_17859,N_11023,N_12401);
nor U17860 (N_17860,N_14160,N_11055);
or U17861 (N_17861,N_12448,N_10400);
nor U17862 (N_17862,N_12087,N_10942);
or U17863 (N_17863,N_12560,N_11669);
or U17864 (N_17864,N_11684,N_13453);
and U17865 (N_17865,N_13260,N_12749);
or U17866 (N_17866,N_12032,N_12030);
or U17867 (N_17867,N_14018,N_12206);
nand U17868 (N_17868,N_14393,N_14734);
and U17869 (N_17869,N_14235,N_13595);
and U17870 (N_17870,N_10301,N_11338);
or U17871 (N_17871,N_14383,N_14135);
nor U17872 (N_17872,N_10737,N_14309);
and U17873 (N_17873,N_12757,N_11671);
nand U17874 (N_17874,N_11980,N_12319);
and U17875 (N_17875,N_10491,N_13668);
nor U17876 (N_17876,N_14971,N_12615);
or U17877 (N_17877,N_12471,N_13338);
and U17878 (N_17878,N_14218,N_13795);
or U17879 (N_17879,N_12655,N_11693);
or U17880 (N_17880,N_14344,N_11496);
or U17881 (N_17881,N_11889,N_14207);
or U17882 (N_17882,N_14835,N_14052);
nor U17883 (N_17883,N_11265,N_11083);
nor U17884 (N_17884,N_14823,N_14607);
nand U17885 (N_17885,N_13739,N_14883);
nor U17886 (N_17886,N_11141,N_13613);
and U17887 (N_17887,N_12891,N_14771);
or U17888 (N_17888,N_14938,N_11634);
xor U17889 (N_17889,N_13822,N_11704);
or U17890 (N_17890,N_12065,N_13759);
nand U17891 (N_17891,N_11486,N_14395);
or U17892 (N_17892,N_13125,N_13604);
or U17893 (N_17893,N_10295,N_14673);
nor U17894 (N_17894,N_10728,N_10082);
nor U17895 (N_17895,N_11838,N_11739);
or U17896 (N_17896,N_14557,N_14980);
nor U17897 (N_17897,N_10743,N_12599);
nand U17898 (N_17898,N_14478,N_11031);
and U17899 (N_17899,N_10070,N_11638);
or U17900 (N_17900,N_12554,N_11167);
nor U17901 (N_17901,N_12389,N_14916);
and U17902 (N_17902,N_13460,N_11627);
nand U17903 (N_17903,N_11233,N_14383);
and U17904 (N_17904,N_10830,N_10494);
and U17905 (N_17905,N_14021,N_14915);
nand U17906 (N_17906,N_13293,N_12661);
and U17907 (N_17907,N_10613,N_11092);
nand U17908 (N_17908,N_13154,N_13296);
or U17909 (N_17909,N_14857,N_14898);
or U17910 (N_17910,N_13994,N_14021);
or U17911 (N_17911,N_14573,N_10091);
or U17912 (N_17912,N_12195,N_13282);
and U17913 (N_17913,N_14622,N_14952);
nor U17914 (N_17914,N_11138,N_13404);
or U17915 (N_17915,N_11881,N_13022);
nor U17916 (N_17916,N_11053,N_12787);
or U17917 (N_17917,N_14156,N_11895);
and U17918 (N_17918,N_12799,N_10334);
nand U17919 (N_17919,N_11233,N_13957);
and U17920 (N_17920,N_10902,N_11349);
nand U17921 (N_17921,N_11507,N_14785);
nand U17922 (N_17922,N_12720,N_14261);
nand U17923 (N_17923,N_12991,N_13607);
and U17924 (N_17924,N_12024,N_13339);
or U17925 (N_17925,N_14696,N_12898);
and U17926 (N_17926,N_11157,N_13464);
nand U17927 (N_17927,N_13671,N_11391);
nand U17928 (N_17928,N_12452,N_11787);
nand U17929 (N_17929,N_12024,N_10412);
or U17930 (N_17930,N_12042,N_12991);
nand U17931 (N_17931,N_11115,N_13192);
and U17932 (N_17932,N_11922,N_13640);
nand U17933 (N_17933,N_10046,N_11233);
and U17934 (N_17934,N_13481,N_13938);
nor U17935 (N_17935,N_11577,N_14770);
or U17936 (N_17936,N_12258,N_13015);
nand U17937 (N_17937,N_12746,N_10877);
xnor U17938 (N_17938,N_11183,N_14450);
and U17939 (N_17939,N_12118,N_13105);
and U17940 (N_17940,N_11921,N_11889);
nand U17941 (N_17941,N_13829,N_13240);
nor U17942 (N_17942,N_14083,N_12885);
and U17943 (N_17943,N_12259,N_10587);
and U17944 (N_17944,N_14577,N_12776);
and U17945 (N_17945,N_14782,N_12711);
nor U17946 (N_17946,N_14687,N_11606);
nor U17947 (N_17947,N_12956,N_13876);
nor U17948 (N_17948,N_14230,N_14375);
nor U17949 (N_17949,N_14610,N_14912);
nor U17950 (N_17950,N_13377,N_14479);
nor U17951 (N_17951,N_10127,N_13491);
or U17952 (N_17952,N_11792,N_10324);
or U17953 (N_17953,N_12277,N_10137);
and U17954 (N_17954,N_10431,N_13982);
nor U17955 (N_17955,N_12997,N_11883);
and U17956 (N_17956,N_13116,N_10194);
or U17957 (N_17957,N_11114,N_12845);
nor U17958 (N_17958,N_12781,N_11958);
or U17959 (N_17959,N_11299,N_10842);
or U17960 (N_17960,N_13537,N_14626);
and U17961 (N_17961,N_10903,N_14124);
nand U17962 (N_17962,N_12587,N_14433);
or U17963 (N_17963,N_10777,N_10534);
nand U17964 (N_17964,N_10379,N_11089);
and U17965 (N_17965,N_11755,N_10166);
nand U17966 (N_17966,N_13992,N_14200);
or U17967 (N_17967,N_10339,N_12865);
and U17968 (N_17968,N_13623,N_10223);
and U17969 (N_17969,N_11756,N_13691);
nand U17970 (N_17970,N_11190,N_14248);
or U17971 (N_17971,N_13457,N_11491);
nor U17972 (N_17972,N_10889,N_11628);
or U17973 (N_17973,N_10645,N_12379);
nor U17974 (N_17974,N_13694,N_12151);
xor U17975 (N_17975,N_12272,N_14807);
nand U17976 (N_17976,N_13565,N_12939);
or U17977 (N_17977,N_14032,N_12966);
nor U17978 (N_17978,N_10672,N_12017);
nor U17979 (N_17979,N_11484,N_13766);
nor U17980 (N_17980,N_12640,N_12016);
xor U17981 (N_17981,N_10576,N_14371);
nand U17982 (N_17982,N_11878,N_11479);
or U17983 (N_17983,N_11540,N_12969);
and U17984 (N_17984,N_11782,N_12697);
and U17985 (N_17985,N_10758,N_12037);
xnor U17986 (N_17986,N_12895,N_12775);
nand U17987 (N_17987,N_11213,N_12602);
nor U17988 (N_17988,N_12760,N_13964);
and U17989 (N_17989,N_13178,N_14792);
or U17990 (N_17990,N_13838,N_11222);
nor U17991 (N_17991,N_10864,N_13298);
or U17992 (N_17992,N_12842,N_14020);
or U17993 (N_17993,N_11077,N_10567);
nor U17994 (N_17994,N_10178,N_13728);
or U17995 (N_17995,N_13252,N_10026);
and U17996 (N_17996,N_13692,N_11357);
or U17997 (N_17997,N_10897,N_11081);
or U17998 (N_17998,N_11698,N_13659);
nand U17999 (N_17999,N_13787,N_13050);
and U18000 (N_18000,N_11115,N_14738);
or U18001 (N_18001,N_12919,N_11616);
nor U18002 (N_18002,N_11257,N_14729);
nor U18003 (N_18003,N_12300,N_13447);
nand U18004 (N_18004,N_13124,N_12683);
nand U18005 (N_18005,N_11616,N_10192);
nand U18006 (N_18006,N_11291,N_11633);
and U18007 (N_18007,N_10343,N_12103);
nor U18008 (N_18008,N_12217,N_10903);
and U18009 (N_18009,N_14005,N_12684);
or U18010 (N_18010,N_13776,N_11218);
nor U18011 (N_18011,N_11484,N_12058);
or U18012 (N_18012,N_11984,N_12169);
and U18013 (N_18013,N_11658,N_13306);
nand U18014 (N_18014,N_11702,N_14330);
nor U18015 (N_18015,N_12427,N_13363);
nand U18016 (N_18016,N_14381,N_12356);
or U18017 (N_18017,N_13085,N_13621);
and U18018 (N_18018,N_13882,N_14587);
nand U18019 (N_18019,N_14152,N_10253);
or U18020 (N_18020,N_12852,N_11621);
nor U18021 (N_18021,N_12757,N_10194);
nand U18022 (N_18022,N_13658,N_10688);
nand U18023 (N_18023,N_11050,N_10082);
xnor U18024 (N_18024,N_12848,N_14971);
or U18025 (N_18025,N_11608,N_13685);
and U18026 (N_18026,N_13025,N_13923);
nand U18027 (N_18027,N_13819,N_12965);
and U18028 (N_18028,N_13166,N_10420);
or U18029 (N_18029,N_11523,N_12226);
nor U18030 (N_18030,N_12347,N_10694);
or U18031 (N_18031,N_11591,N_12935);
nand U18032 (N_18032,N_12844,N_10348);
nand U18033 (N_18033,N_14286,N_14268);
nor U18034 (N_18034,N_10013,N_12921);
or U18035 (N_18035,N_14762,N_10526);
or U18036 (N_18036,N_10694,N_14533);
nor U18037 (N_18037,N_14025,N_12452);
nand U18038 (N_18038,N_10354,N_10002);
nand U18039 (N_18039,N_14134,N_11985);
nand U18040 (N_18040,N_13402,N_14540);
and U18041 (N_18041,N_10907,N_10671);
and U18042 (N_18042,N_10259,N_11573);
nand U18043 (N_18043,N_13265,N_13147);
and U18044 (N_18044,N_12611,N_11306);
nor U18045 (N_18045,N_11290,N_13125);
nand U18046 (N_18046,N_10684,N_14154);
nor U18047 (N_18047,N_10342,N_10621);
or U18048 (N_18048,N_12149,N_13924);
nand U18049 (N_18049,N_10711,N_14206);
nand U18050 (N_18050,N_11454,N_10805);
or U18051 (N_18051,N_10470,N_10322);
nor U18052 (N_18052,N_14273,N_12815);
nand U18053 (N_18053,N_11110,N_12459);
nor U18054 (N_18054,N_10798,N_10147);
nor U18055 (N_18055,N_13339,N_11434);
nor U18056 (N_18056,N_10768,N_14794);
nor U18057 (N_18057,N_12191,N_14027);
nand U18058 (N_18058,N_10964,N_12485);
or U18059 (N_18059,N_11938,N_12619);
or U18060 (N_18060,N_12805,N_10914);
nor U18061 (N_18061,N_14827,N_10653);
or U18062 (N_18062,N_14949,N_13883);
or U18063 (N_18063,N_12230,N_10707);
or U18064 (N_18064,N_14152,N_13587);
nand U18065 (N_18065,N_10928,N_12295);
nor U18066 (N_18066,N_10473,N_10368);
nand U18067 (N_18067,N_12565,N_13496);
or U18068 (N_18068,N_11870,N_10848);
nor U18069 (N_18069,N_12818,N_12618);
or U18070 (N_18070,N_12195,N_12986);
nor U18071 (N_18071,N_12828,N_11397);
xnor U18072 (N_18072,N_10791,N_11940);
and U18073 (N_18073,N_10225,N_14940);
or U18074 (N_18074,N_11824,N_14143);
nor U18075 (N_18075,N_10065,N_14961);
or U18076 (N_18076,N_12548,N_14794);
nand U18077 (N_18077,N_11176,N_13475);
and U18078 (N_18078,N_12686,N_12860);
and U18079 (N_18079,N_10731,N_11953);
and U18080 (N_18080,N_10667,N_12000);
or U18081 (N_18081,N_10773,N_13432);
or U18082 (N_18082,N_13178,N_14832);
or U18083 (N_18083,N_14629,N_13713);
or U18084 (N_18084,N_13142,N_10825);
nor U18085 (N_18085,N_13269,N_12818);
and U18086 (N_18086,N_14896,N_13624);
or U18087 (N_18087,N_12903,N_13969);
and U18088 (N_18088,N_11968,N_12438);
and U18089 (N_18089,N_12229,N_11521);
nand U18090 (N_18090,N_11075,N_13057);
and U18091 (N_18091,N_12755,N_11665);
nor U18092 (N_18092,N_10251,N_14253);
nand U18093 (N_18093,N_12708,N_11590);
or U18094 (N_18094,N_11936,N_14260);
nor U18095 (N_18095,N_11291,N_11007);
nand U18096 (N_18096,N_11473,N_14219);
or U18097 (N_18097,N_10112,N_11436);
nand U18098 (N_18098,N_14148,N_13716);
or U18099 (N_18099,N_10936,N_11217);
nand U18100 (N_18100,N_10059,N_11977);
and U18101 (N_18101,N_10815,N_14443);
and U18102 (N_18102,N_11160,N_14005);
and U18103 (N_18103,N_12644,N_14547);
nand U18104 (N_18104,N_11025,N_14781);
nand U18105 (N_18105,N_11127,N_13910);
nand U18106 (N_18106,N_13816,N_12797);
or U18107 (N_18107,N_12952,N_10387);
nor U18108 (N_18108,N_12656,N_14117);
and U18109 (N_18109,N_10907,N_13402);
nor U18110 (N_18110,N_12522,N_11175);
nor U18111 (N_18111,N_12365,N_13159);
xnor U18112 (N_18112,N_14836,N_13505);
or U18113 (N_18113,N_10826,N_12826);
or U18114 (N_18114,N_10785,N_12680);
nand U18115 (N_18115,N_11596,N_11007);
and U18116 (N_18116,N_14472,N_13425);
nand U18117 (N_18117,N_11841,N_14944);
or U18118 (N_18118,N_14625,N_13811);
or U18119 (N_18119,N_10624,N_12967);
nor U18120 (N_18120,N_14439,N_10712);
or U18121 (N_18121,N_12278,N_14385);
and U18122 (N_18122,N_10485,N_10616);
nor U18123 (N_18123,N_10166,N_14694);
and U18124 (N_18124,N_13661,N_12518);
nor U18125 (N_18125,N_11277,N_13278);
or U18126 (N_18126,N_11728,N_10989);
nand U18127 (N_18127,N_13248,N_12966);
nand U18128 (N_18128,N_10487,N_11223);
nor U18129 (N_18129,N_11847,N_10965);
or U18130 (N_18130,N_14584,N_13877);
nor U18131 (N_18131,N_13127,N_12989);
nor U18132 (N_18132,N_11136,N_12857);
nand U18133 (N_18133,N_13757,N_10603);
and U18134 (N_18134,N_12475,N_14043);
or U18135 (N_18135,N_13395,N_12141);
nor U18136 (N_18136,N_13050,N_12575);
and U18137 (N_18137,N_11904,N_14368);
and U18138 (N_18138,N_14001,N_14941);
or U18139 (N_18139,N_13700,N_12391);
nor U18140 (N_18140,N_12229,N_13548);
nand U18141 (N_18141,N_14033,N_13227);
nor U18142 (N_18142,N_10013,N_10211);
nand U18143 (N_18143,N_13914,N_14980);
or U18144 (N_18144,N_11313,N_11340);
nor U18145 (N_18145,N_10751,N_14547);
and U18146 (N_18146,N_10271,N_12954);
or U18147 (N_18147,N_13546,N_12938);
or U18148 (N_18148,N_10237,N_12946);
and U18149 (N_18149,N_13246,N_10875);
or U18150 (N_18150,N_14330,N_14934);
and U18151 (N_18151,N_12930,N_14258);
nor U18152 (N_18152,N_10742,N_13727);
nor U18153 (N_18153,N_10925,N_11108);
or U18154 (N_18154,N_10515,N_11679);
nor U18155 (N_18155,N_14288,N_13488);
and U18156 (N_18156,N_13332,N_10072);
nor U18157 (N_18157,N_11304,N_14838);
and U18158 (N_18158,N_11893,N_13473);
nand U18159 (N_18159,N_13766,N_12846);
and U18160 (N_18160,N_13909,N_10534);
and U18161 (N_18161,N_11593,N_12776);
or U18162 (N_18162,N_13276,N_12080);
and U18163 (N_18163,N_13933,N_10154);
nand U18164 (N_18164,N_11954,N_10358);
and U18165 (N_18165,N_11680,N_11947);
nor U18166 (N_18166,N_11438,N_12925);
nor U18167 (N_18167,N_10471,N_10632);
nand U18168 (N_18168,N_11171,N_12242);
nand U18169 (N_18169,N_13009,N_11812);
and U18170 (N_18170,N_11532,N_11958);
and U18171 (N_18171,N_12387,N_11587);
or U18172 (N_18172,N_13750,N_14167);
or U18173 (N_18173,N_11877,N_13931);
or U18174 (N_18174,N_13805,N_10079);
nor U18175 (N_18175,N_14600,N_12793);
nand U18176 (N_18176,N_14367,N_12343);
or U18177 (N_18177,N_10077,N_11263);
and U18178 (N_18178,N_11295,N_14391);
nor U18179 (N_18179,N_12325,N_10144);
nor U18180 (N_18180,N_14750,N_12526);
nand U18181 (N_18181,N_12771,N_11701);
nand U18182 (N_18182,N_10576,N_13612);
nor U18183 (N_18183,N_12032,N_12099);
nor U18184 (N_18184,N_10474,N_10896);
and U18185 (N_18185,N_11505,N_12634);
nand U18186 (N_18186,N_10278,N_14113);
nand U18187 (N_18187,N_13892,N_12897);
or U18188 (N_18188,N_11547,N_14952);
and U18189 (N_18189,N_14178,N_14556);
or U18190 (N_18190,N_11836,N_12988);
or U18191 (N_18191,N_12214,N_14283);
nand U18192 (N_18192,N_10496,N_10728);
and U18193 (N_18193,N_10655,N_13013);
and U18194 (N_18194,N_13143,N_13795);
and U18195 (N_18195,N_11613,N_11642);
nor U18196 (N_18196,N_13817,N_10723);
nor U18197 (N_18197,N_14150,N_11693);
nor U18198 (N_18198,N_12585,N_11582);
and U18199 (N_18199,N_12622,N_12640);
or U18200 (N_18200,N_12538,N_13799);
nor U18201 (N_18201,N_12000,N_12616);
nand U18202 (N_18202,N_14703,N_11272);
and U18203 (N_18203,N_10519,N_11166);
nand U18204 (N_18204,N_10374,N_13018);
nor U18205 (N_18205,N_12557,N_10324);
or U18206 (N_18206,N_14125,N_14262);
nor U18207 (N_18207,N_13218,N_12783);
and U18208 (N_18208,N_13969,N_14856);
or U18209 (N_18209,N_11976,N_11561);
nor U18210 (N_18210,N_10607,N_14141);
and U18211 (N_18211,N_10496,N_10046);
nand U18212 (N_18212,N_14972,N_11470);
and U18213 (N_18213,N_10828,N_11376);
nor U18214 (N_18214,N_13934,N_14517);
and U18215 (N_18215,N_12193,N_11149);
nand U18216 (N_18216,N_13367,N_12044);
or U18217 (N_18217,N_10260,N_11403);
nor U18218 (N_18218,N_12965,N_11953);
or U18219 (N_18219,N_13795,N_13256);
nor U18220 (N_18220,N_14863,N_12811);
nand U18221 (N_18221,N_13412,N_12969);
nand U18222 (N_18222,N_12674,N_12587);
or U18223 (N_18223,N_10238,N_12441);
nor U18224 (N_18224,N_11748,N_11393);
and U18225 (N_18225,N_14947,N_13687);
and U18226 (N_18226,N_13584,N_13416);
or U18227 (N_18227,N_12599,N_13905);
nor U18228 (N_18228,N_14559,N_14952);
or U18229 (N_18229,N_13755,N_10289);
nand U18230 (N_18230,N_10658,N_13828);
or U18231 (N_18231,N_13131,N_11627);
xor U18232 (N_18232,N_14272,N_13063);
nand U18233 (N_18233,N_12005,N_10580);
nor U18234 (N_18234,N_13173,N_14558);
or U18235 (N_18235,N_12168,N_11032);
or U18236 (N_18236,N_13526,N_13908);
or U18237 (N_18237,N_10577,N_11755);
and U18238 (N_18238,N_14607,N_12177);
and U18239 (N_18239,N_13783,N_12791);
and U18240 (N_18240,N_14631,N_11764);
nor U18241 (N_18241,N_10869,N_14582);
nand U18242 (N_18242,N_14767,N_12764);
nand U18243 (N_18243,N_11853,N_11002);
or U18244 (N_18244,N_10089,N_10224);
and U18245 (N_18245,N_14459,N_10249);
or U18246 (N_18246,N_10251,N_10334);
or U18247 (N_18247,N_13769,N_11469);
and U18248 (N_18248,N_12636,N_12598);
nand U18249 (N_18249,N_10134,N_13452);
and U18250 (N_18250,N_11640,N_12889);
and U18251 (N_18251,N_14561,N_11163);
or U18252 (N_18252,N_11206,N_12957);
nand U18253 (N_18253,N_12760,N_14187);
nor U18254 (N_18254,N_11513,N_13410);
or U18255 (N_18255,N_12053,N_13234);
nand U18256 (N_18256,N_12324,N_12320);
and U18257 (N_18257,N_13610,N_14394);
nor U18258 (N_18258,N_11266,N_12094);
or U18259 (N_18259,N_14032,N_11128);
and U18260 (N_18260,N_14826,N_13722);
nand U18261 (N_18261,N_12864,N_12985);
nand U18262 (N_18262,N_12315,N_11809);
or U18263 (N_18263,N_14971,N_14349);
or U18264 (N_18264,N_13257,N_14752);
and U18265 (N_18265,N_12604,N_14080);
and U18266 (N_18266,N_14807,N_10451);
or U18267 (N_18267,N_14078,N_12985);
or U18268 (N_18268,N_12412,N_14118);
or U18269 (N_18269,N_14649,N_13162);
nand U18270 (N_18270,N_13199,N_12266);
or U18271 (N_18271,N_11233,N_14043);
nand U18272 (N_18272,N_11353,N_11518);
nor U18273 (N_18273,N_11913,N_12253);
and U18274 (N_18274,N_10926,N_10524);
nand U18275 (N_18275,N_13945,N_13015);
and U18276 (N_18276,N_12070,N_14228);
and U18277 (N_18277,N_13360,N_13042);
nand U18278 (N_18278,N_13985,N_10713);
nand U18279 (N_18279,N_14164,N_13622);
and U18280 (N_18280,N_10241,N_11545);
or U18281 (N_18281,N_13261,N_11416);
nor U18282 (N_18282,N_14290,N_10623);
nand U18283 (N_18283,N_13451,N_10098);
and U18284 (N_18284,N_14407,N_13730);
nand U18285 (N_18285,N_11441,N_14683);
nand U18286 (N_18286,N_10500,N_11787);
nor U18287 (N_18287,N_13914,N_12937);
xnor U18288 (N_18288,N_12758,N_13337);
or U18289 (N_18289,N_12504,N_10166);
or U18290 (N_18290,N_11422,N_11910);
nor U18291 (N_18291,N_12603,N_14132);
nor U18292 (N_18292,N_12851,N_11474);
nand U18293 (N_18293,N_10335,N_14920);
or U18294 (N_18294,N_10313,N_13640);
and U18295 (N_18295,N_13337,N_11388);
and U18296 (N_18296,N_10645,N_12610);
and U18297 (N_18297,N_11249,N_14885);
nand U18298 (N_18298,N_14358,N_11264);
nor U18299 (N_18299,N_10767,N_12674);
nor U18300 (N_18300,N_12808,N_14706);
or U18301 (N_18301,N_10835,N_10905);
or U18302 (N_18302,N_14930,N_11079);
or U18303 (N_18303,N_11577,N_13050);
or U18304 (N_18304,N_10075,N_14370);
nand U18305 (N_18305,N_10108,N_10266);
and U18306 (N_18306,N_12098,N_14263);
or U18307 (N_18307,N_11133,N_13492);
and U18308 (N_18308,N_13621,N_12334);
and U18309 (N_18309,N_10610,N_10985);
nor U18310 (N_18310,N_13375,N_11822);
and U18311 (N_18311,N_10705,N_13950);
nand U18312 (N_18312,N_12306,N_11062);
and U18313 (N_18313,N_13635,N_10990);
nand U18314 (N_18314,N_10143,N_12981);
and U18315 (N_18315,N_14764,N_14839);
or U18316 (N_18316,N_11254,N_11810);
and U18317 (N_18317,N_11068,N_13880);
nand U18318 (N_18318,N_10421,N_11165);
or U18319 (N_18319,N_11900,N_10661);
nor U18320 (N_18320,N_12011,N_14756);
nand U18321 (N_18321,N_11240,N_11401);
or U18322 (N_18322,N_13275,N_14289);
nor U18323 (N_18323,N_13403,N_10094);
or U18324 (N_18324,N_12907,N_13933);
or U18325 (N_18325,N_13168,N_12617);
or U18326 (N_18326,N_14585,N_10583);
or U18327 (N_18327,N_13971,N_12061);
and U18328 (N_18328,N_12839,N_11480);
and U18329 (N_18329,N_13074,N_11022);
or U18330 (N_18330,N_12703,N_13228);
nand U18331 (N_18331,N_11291,N_12781);
nor U18332 (N_18332,N_10440,N_14696);
nor U18333 (N_18333,N_10638,N_12741);
nor U18334 (N_18334,N_11805,N_10503);
or U18335 (N_18335,N_10106,N_12553);
and U18336 (N_18336,N_10296,N_11580);
or U18337 (N_18337,N_14189,N_11261);
or U18338 (N_18338,N_12395,N_13791);
nand U18339 (N_18339,N_10824,N_12444);
and U18340 (N_18340,N_14721,N_10872);
nor U18341 (N_18341,N_10312,N_12916);
or U18342 (N_18342,N_11045,N_11638);
or U18343 (N_18343,N_14064,N_13625);
or U18344 (N_18344,N_13904,N_12403);
and U18345 (N_18345,N_11943,N_14070);
nand U18346 (N_18346,N_13160,N_10201);
nor U18347 (N_18347,N_14247,N_10628);
nand U18348 (N_18348,N_12872,N_10850);
and U18349 (N_18349,N_11556,N_14368);
nand U18350 (N_18350,N_14180,N_11728);
and U18351 (N_18351,N_13934,N_12642);
nor U18352 (N_18352,N_12500,N_14967);
or U18353 (N_18353,N_11348,N_10312);
nor U18354 (N_18354,N_11575,N_12755);
nand U18355 (N_18355,N_14981,N_12046);
and U18356 (N_18356,N_10288,N_13992);
nand U18357 (N_18357,N_12669,N_14690);
nand U18358 (N_18358,N_11544,N_13042);
nor U18359 (N_18359,N_13812,N_13197);
or U18360 (N_18360,N_10913,N_11060);
nand U18361 (N_18361,N_10558,N_12816);
nor U18362 (N_18362,N_12796,N_12350);
or U18363 (N_18363,N_14044,N_14960);
nor U18364 (N_18364,N_10186,N_12850);
nand U18365 (N_18365,N_11064,N_10187);
nand U18366 (N_18366,N_10007,N_14708);
or U18367 (N_18367,N_13980,N_13644);
nor U18368 (N_18368,N_14292,N_14824);
nand U18369 (N_18369,N_11240,N_13554);
and U18370 (N_18370,N_12621,N_11469);
xnor U18371 (N_18371,N_13350,N_12689);
or U18372 (N_18372,N_13288,N_12805);
nor U18373 (N_18373,N_14153,N_12000);
and U18374 (N_18374,N_13576,N_11202);
nand U18375 (N_18375,N_10200,N_12236);
or U18376 (N_18376,N_13128,N_13324);
nand U18377 (N_18377,N_11660,N_14826);
or U18378 (N_18378,N_13558,N_12446);
and U18379 (N_18379,N_13198,N_12927);
and U18380 (N_18380,N_14424,N_10092);
or U18381 (N_18381,N_10168,N_14875);
and U18382 (N_18382,N_12235,N_12008);
nand U18383 (N_18383,N_14791,N_11777);
nand U18384 (N_18384,N_14117,N_14312);
nor U18385 (N_18385,N_12389,N_12099);
or U18386 (N_18386,N_13712,N_13689);
nand U18387 (N_18387,N_14929,N_11496);
nand U18388 (N_18388,N_10227,N_10312);
or U18389 (N_18389,N_12699,N_10632);
and U18390 (N_18390,N_12018,N_12399);
nand U18391 (N_18391,N_13879,N_14684);
or U18392 (N_18392,N_11563,N_14362);
nand U18393 (N_18393,N_13459,N_13895);
and U18394 (N_18394,N_11171,N_10383);
nand U18395 (N_18395,N_13235,N_10374);
nor U18396 (N_18396,N_12123,N_14560);
and U18397 (N_18397,N_11130,N_14517);
nand U18398 (N_18398,N_12285,N_14319);
nand U18399 (N_18399,N_10055,N_12355);
nor U18400 (N_18400,N_13355,N_10769);
and U18401 (N_18401,N_12942,N_11305);
nor U18402 (N_18402,N_13289,N_12550);
and U18403 (N_18403,N_14302,N_13210);
and U18404 (N_18404,N_13554,N_12305);
nor U18405 (N_18405,N_14861,N_12521);
nand U18406 (N_18406,N_14206,N_12169);
nand U18407 (N_18407,N_11108,N_11364);
xnor U18408 (N_18408,N_11478,N_13149);
and U18409 (N_18409,N_11846,N_11721);
or U18410 (N_18410,N_11039,N_12727);
nand U18411 (N_18411,N_14635,N_14873);
nor U18412 (N_18412,N_13305,N_10503);
nor U18413 (N_18413,N_13542,N_11304);
or U18414 (N_18414,N_14918,N_12535);
and U18415 (N_18415,N_13101,N_11350);
nand U18416 (N_18416,N_11808,N_13771);
nand U18417 (N_18417,N_14391,N_11519);
nor U18418 (N_18418,N_12514,N_11288);
nand U18419 (N_18419,N_12573,N_10683);
nor U18420 (N_18420,N_11671,N_10168);
nor U18421 (N_18421,N_12619,N_14730);
and U18422 (N_18422,N_10276,N_10324);
nand U18423 (N_18423,N_10851,N_13577);
nand U18424 (N_18424,N_13243,N_10165);
and U18425 (N_18425,N_13874,N_11306);
nand U18426 (N_18426,N_14189,N_11386);
nor U18427 (N_18427,N_12393,N_10957);
nand U18428 (N_18428,N_12174,N_14170);
or U18429 (N_18429,N_11662,N_10020);
and U18430 (N_18430,N_13536,N_13656);
and U18431 (N_18431,N_14025,N_13589);
nor U18432 (N_18432,N_10267,N_14969);
or U18433 (N_18433,N_10210,N_10766);
and U18434 (N_18434,N_13895,N_11007);
or U18435 (N_18435,N_14309,N_13448);
nand U18436 (N_18436,N_10495,N_11760);
nor U18437 (N_18437,N_13139,N_12526);
nor U18438 (N_18438,N_14325,N_13068);
nor U18439 (N_18439,N_11476,N_13952);
nand U18440 (N_18440,N_11823,N_14766);
or U18441 (N_18441,N_10890,N_12186);
and U18442 (N_18442,N_11134,N_14686);
nor U18443 (N_18443,N_10980,N_13506);
nand U18444 (N_18444,N_13124,N_11398);
and U18445 (N_18445,N_14541,N_10717);
and U18446 (N_18446,N_13210,N_13341);
or U18447 (N_18447,N_14066,N_13879);
or U18448 (N_18448,N_11236,N_13016);
or U18449 (N_18449,N_14750,N_10051);
or U18450 (N_18450,N_12993,N_12483);
nor U18451 (N_18451,N_13954,N_11196);
nor U18452 (N_18452,N_10132,N_12273);
nand U18453 (N_18453,N_12977,N_12309);
and U18454 (N_18454,N_11063,N_14301);
and U18455 (N_18455,N_13460,N_13892);
or U18456 (N_18456,N_12065,N_14846);
nor U18457 (N_18457,N_10907,N_10285);
or U18458 (N_18458,N_10685,N_12077);
or U18459 (N_18459,N_12254,N_10479);
or U18460 (N_18460,N_13308,N_11957);
or U18461 (N_18461,N_14334,N_10588);
and U18462 (N_18462,N_12654,N_13339);
nand U18463 (N_18463,N_10121,N_13384);
and U18464 (N_18464,N_11323,N_12085);
and U18465 (N_18465,N_13853,N_13437);
nor U18466 (N_18466,N_10797,N_13196);
nand U18467 (N_18467,N_12031,N_12036);
nand U18468 (N_18468,N_14421,N_12165);
or U18469 (N_18469,N_14640,N_13063);
nand U18470 (N_18470,N_14095,N_13297);
nand U18471 (N_18471,N_12881,N_12859);
nand U18472 (N_18472,N_10473,N_14488);
nor U18473 (N_18473,N_11221,N_13884);
and U18474 (N_18474,N_14065,N_12244);
or U18475 (N_18475,N_14675,N_13608);
nand U18476 (N_18476,N_11362,N_13240);
and U18477 (N_18477,N_12926,N_13134);
or U18478 (N_18478,N_13951,N_11354);
nand U18479 (N_18479,N_14285,N_11708);
or U18480 (N_18480,N_13177,N_11006);
or U18481 (N_18481,N_14111,N_12641);
and U18482 (N_18482,N_10623,N_10577);
or U18483 (N_18483,N_12659,N_11516);
nand U18484 (N_18484,N_12198,N_12836);
or U18485 (N_18485,N_11052,N_10448);
and U18486 (N_18486,N_11939,N_12614);
nor U18487 (N_18487,N_13797,N_12662);
or U18488 (N_18488,N_13560,N_10763);
nor U18489 (N_18489,N_12571,N_11670);
and U18490 (N_18490,N_12070,N_10012);
nand U18491 (N_18491,N_11954,N_12556);
nand U18492 (N_18492,N_14206,N_12373);
or U18493 (N_18493,N_10115,N_10095);
nand U18494 (N_18494,N_14354,N_13472);
nor U18495 (N_18495,N_12700,N_13591);
and U18496 (N_18496,N_12815,N_12504);
or U18497 (N_18497,N_13517,N_13625);
nand U18498 (N_18498,N_13613,N_11799);
or U18499 (N_18499,N_14214,N_12588);
or U18500 (N_18500,N_12726,N_12166);
nor U18501 (N_18501,N_14132,N_11551);
xor U18502 (N_18502,N_13777,N_14513);
nand U18503 (N_18503,N_10090,N_14345);
nand U18504 (N_18504,N_13426,N_13824);
and U18505 (N_18505,N_10442,N_12750);
nand U18506 (N_18506,N_14029,N_10966);
or U18507 (N_18507,N_14692,N_10071);
or U18508 (N_18508,N_12479,N_14950);
and U18509 (N_18509,N_10568,N_12217);
nand U18510 (N_18510,N_11567,N_14228);
nor U18511 (N_18511,N_12294,N_10759);
or U18512 (N_18512,N_12402,N_12145);
and U18513 (N_18513,N_10411,N_13906);
nand U18514 (N_18514,N_14903,N_10335);
or U18515 (N_18515,N_11299,N_11269);
nand U18516 (N_18516,N_12860,N_12643);
nand U18517 (N_18517,N_12997,N_11546);
nand U18518 (N_18518,N_13836,N_13208);
nor U18519 (N_18519,N_14481,N_11795);
nor U18520 (N_18520,N_12894,N_13455);
nor U18521 (N_18521,N_10751,N_12746);
nand U18522 (N_18522,N_11489,N_14620);
nor U18523 (N_18523,N_14904,N_11198);
and U18524 (N_18524,N_13066,N_11137);
and U18525 (N_18525,N_13618,N_14135);
and U18526 (N_18526,N_12348,N_11102);
and U18527 (N_18527,N_13800,N_10093);
or U18528 (N_18528,N_12322,N_14903);
or U18529 (N_18529,N_12200,N_10504);
nand U18530 (N_18530,N_14637,N_13183);
and U18531 (N_18531,N_14737,N_14105);
and U18532 (N_18532,N_14881,N_12954);
and U18533 (N_18533,N_10322,N_11729);
nand U18534 (N_18534,N_12827,N_14985);
or U18535 (N_18535,N_10462,N_11715);
nand U18536 (N_18536,N_11208,N_10773);
nor U18537 (N_18537,N_14774,N_11516);
and U18538 (N_18538,N_10738,N_10377);
nand U18539 (N_18539,N_14199,N_14866);
and U18540 (N_18540,N_12276,N_14967);
and U18541 (N_18541,N_13174,N_11123);
nor U18542 (N_18542,N_10467,N_10717);
and U18543 (N_18543,N_10380,N_13100);
nand U18544 (N_18544,N_10509,N_12238);
or U18545 (N_18545,N_13646,N_11531);
or U18546 (N_18546,N_12639,N_10693);
nor U18547 (N_18547,N_13053,N_11822);
nand U18548 (N_18548,N_11445,N_14988);
or U18549 (N_18549,N_12606,N_10725);
and U18550 (N_18550,N_10916,N_11864);
and U18551 (N_18551,N_14575,N_12441);
nor U18552 (N_18552,N_12130,N_10441);
or U18553 (N_18553,N_13271,N_13676);
or U18554 (N_18554,N_10175,N_11323);
and U18555 (N_18555,N_12776,N_13398);
nor U18556 (N_18556,N_13277,N_14047);
or U18557 (N_18557,N_14338,N_11154);
or U18558 (N_18558,N_10978,N_13250);
or U18559 (N_18559,N_10620,N_10525);
or U18560 (N_18560,N_11432,N_10143);
and U18561 (N_18561,N_14582,N_13469);
and U18562 (N_18562,N_14087,N_12295);
and U18563 (N_18563,N_13108,N_14278);
nand U18564 (N_18564,N_13431,N_14748);
or U18565 (N_18565,N_14456,N_14542);
nand U18566 (N_18566,N_14094,N_12518);
or U18567 (N_18567,N_14950,N_12470);
nor U18568 (N_18568,N_11138,N_14476);
nand U18569 (N_18569,N_11366,N_10672);
and U18570 (N_18570,N_10938,N_14512);
nor U18571 (N_18571,N_12452,N_11655);
or U18572 (N_18572,N_14033,N_11508);
and U18573 (N_18573,N_11308,N_11324);
nor U18574 (N_18574,N_13052,N_12084);
and U18575 (N_18575,N_13344,N_14270);
and U18576 (N_18576,N_12511,N_14496);
and U18577 (N_18577,N_10948,N_10923);
nand U18578 (N_18578,N_14411,N_12296);
nand U18579 (N_18579,N_10512,N_10758);
nor U18580 (N_18580,N_13480,N_14111);
and U18581 (N_18581,N_13663,N_11811);
nor U18582 (N_18582,N_12072,N_13384);
nor U18583 (N_18583,N_13322,N_13855);
nor U18584 (N_18584,N_14028,N_12801);
nand U18585 (N_18585,N_12598,N_11793);
nor U18586 (N_18586,N_14925,N_12574);
and U18587 (N_18587,N_11796,N_14922);
nand U18588 (N_18588,N_12677,N_11382);
and U18589 (N_18589,N_13747,N_11992);
or U18590 (N_18590,N_14115,N_10338);
nor U18591 (N_18591,N_10263,N_13685);
or U18592 (N_18592,N_14740,N_13483);
and U18593 (N_18593,N_14575,N_11624);
nand U18594 (N_18594,N_13466,N_10009);
or U18595 (N_18595,N_13281,N_10251);
or U18596 (N_18596,N_11739,N_14322);
or U18597 (N_18597,N_14042,N_10622);
or U18598 (N_18598,N_12534,N_12608);
nand U18599 (N_18599,N_13486,N_13367);
nand U18600 (N_18600,N_14192,N_10286);
nand U18601 (N_18601,N_12996,N_12571);
nand U18602 (N_18602,N_10602,N_14294);
nor U18603 (N_18603,N_10671,N_14026);
and U18604 (N_18604,N_13915,N_11335);
nor U18605 (N_18605,N_11981,N_10460);
and U18606 (N_18606,N_13484,N_13258);
or U18607 (N_18607,N_13695,N_14056);
or U18608 (N_18608,N_13997,N_11862);
and U18609 (N_18609,N_11234,N_12256);
nor U18610 (N_18610,N_12969,N_13054);
and U18611 (N_18611,N_12119,N_14506);
or U18612 (N_18612,N_11063,N_12051);
nand U18613 (N_18613,N_11966,N_11283);
nand U18614 (N_18614,N_11517,N_12089);
and U18615 (N_18615,N_12003,N_12455);
nand U18616 (N_18616,N_14377,N_11961);
nand U18617 (N_18617,N_14058,N_14024);
nor U18618 (N_18618,N_10506,N_10842);
nand U18619 (N_18619,N_12020,N_12633);
or U18620 (N_18620,N_12716,N_13403);
or U18621 (N_18621,N_14802,N_13831);
nor U18622 (N_18622,N_13833,N_14439);
nor U18623 (N_18623,N_10991,N_12056);
or U18624 (N_18624,N_11565,N_12246);
nor U18625 (N_18625,N_11071,N_12283);
nand U18626 (N_18626,N_14676,N_14069);
nand U18627 (N_18627,N_14394,N_10690);
or U18628 (N_18628,N_12450,N_10079);
and U18629 (N_18629,N_13478,N_13008);
or U18630 (N_18630,N_11127,N_10539);
nand U18631 (N_18631,N_10250,N_14597);
or U18632 (N_18632,N_12352,N_10725);
nor U18633 (N_18633,N_12111,N_10241);
nor U18634 (N_18634,N_13186,N_13807);
nor U18635 (N_18635,N_12000,N_12166);
and U18636 (N_18636,N_10362,N_14469);
nor U18637 (N_18637,N_14672,N_10962);
and U18638 (N_18638,N_11378,N_12314);
or U18639 (N_18639,N_11772,N_12292);
nand U18640 (N_18640,N_14957,N_10818);
nor U18641 (N_18641,N_13534,N_13211);
and U18642 (N_18642,N_13477,N_12261);
and U18643 (N_18643,N_10162,N_12320);
or U18644 (N_18644,N_12186,N_13332);
nand U18645 (N_18645,N_10172,N_11930);
and U18646 (N_18646,N_12476,N_12383);
or U18647 (N_18647,N_10534,N_14209);
and U18648 (N_18648,N_12412,N_12622);
nand U18649 (N_18649,N_11856,N_11732);
nand U18650 (N_18650,N_10069,N_11981);
nor U18651 (N_18651,N_13858,N_14225);
or U18652 (N_18652,N_12719,N_11141);
nor U18653 (N_18653,N_14036,N_14526);
or U18654 (N_18654,N_10536,N_13417);
nand U18655 (N_18655,N_10177,N_13099);
nor U18656 (N_18656,N_14083,N_13755);
and U18657 (N_18657,N_14768,N_11659);
or U18658 (N_18658,N_13890,N_14787);
and U18659 (N_18659,N_13836,N_11461);
nor U18660 (N_18660,N_14299,N_11515);
or U18661 (N_18661,N_12650,N_10006);
or U18662 (N_18662,N_10791,N_10684);
nor U18663 (N_18663,N_10974,N_10957);
nor U18664 (N_18664,N_13022,N_13387);
and U18665 (N_18665,N_13193,N_11799);
nand U18666 (N_18666,N_10465,N_10419);
nand U18667 (N_18667,N_14619,N_14864);
nand U18668 (N_18668,N_12749,N_10222);
or U18669 (N_18669,N_14197,N_13873);
or U18670 (N_18670,N_14647,N_12886);
and U18671 (N_18671,N_13156,N_14317);
nor U18672 (N_18672,N_13220,N_10469);
and U18673 (N_18673,N_10281,N_10490);
or U18674 (N_18674,N_10117,N_13052);
nor U18675 (N_18675,N_11425,N_11313);
or U18676 (N_18676,N_13901,N_14352);
nand U18677 (N_18677,N_11568,N_13253);
nand U18678 (N_18678,N_10552,N_13341);
nor U18679 (N_18679,N_12791,N_12589);
nand U18680 (N_18680,N_14935,N_14617);
or U18681 (N_18681,N_10426,N_13888);
or U18682 (N_18682,N_14627,N_12002);
nor U18683 (N_18683,N_13918,N_14311);
nor U18684 (N_18684,N_10223,N_13180);
nand U18685 (N_18685,N_14548,N_14879);
nor U18686 (N_18686,N_10847,N_13390);
and U18687 (N_18687,N_12863,N_13162);
and U18688 (N_18688,N_13699,N_11489);
or U18689 (N_18689,N_10029,N_12314);
nand U18690 (N_18690,N_13029,N_11951);
nor U18691 (N_18691,N_10300,N_11880);
and U18692 (N_18692,N_13630,N_11682);
nor U18693 (N_18693,N_10789,N_14052);
and U18694 (N_18694,N_12819,N_12553);
nor U18695 (N_18695,N_14765,N_10249);
nand U18696 (N_18696,N_12094,N_13435);
nor U18697 (N_18697,N_13433,N_14527);
or U18698 (N_18698,N_12190,N_10701);
or U18699 (N_18699,N_12209,N_14531);
and U18700 (N_18700,N_14329,N_13257);
and U18701 (N_18701,N_13110,N_12698);
and U18702 (N_18702,N_14176,N_12236);
nand U18703 (N_18703,N_10074,N_13792);
nand U18704 (N_18704,N_12328,N_10827);
and U18705 (N_18705,N_11556,N_14735);
or U18706 (N_18706,N_14912,N_12263);
nand U18707 (N_18707,N_11042,N_11271);
nand U18708 (N_18708,N_13537,N_10272);
nor U18709 (N_18709,N_13460,N_13293);
nor U18710 (N_18710,N_14709,N_13102);
xnor U18711 (N_18711,N_11078,N_14771);
nand U18712 (N_18712,N_14930,N_12133);
or U18713 (N_18713,N_11243,N_12763);
nand U18714 (N_18714,N_11012,N_14121);
nand U18715 (N_18715,N_13345,N_10411);
or U18716 (N_18716,N_13633,N_14112);
or U18717 (N_18717,N_12897,N_14618);
nand U18718 (N_18718,N_11124,N_14463);
and U18719 (N_18719,N_11593,N_14640);
and U18720 (N_18720,N_13167,N_12050);
or U18721 (N_18721,N_14833,N_11933);
or U18722 (N_18722,N_13429,N_13466);
nand U18723 (N_18723,N_14736,N_14976);
and U18724 (N_18724,N_11786,N_14958);
and U18725 (N_18725,N_11098,N_11799);
and U18726 (N_18726,N_14418,N_10011);
or U18727 (N_18727,N_13428,N_13000);
or U18728 (N_18728,N_11739,N_11732);
nand U18729 (N_18729,N_12224,N_13764);
or U18730 (N_18730,N_11486,N_13072);
or U18731 (N_18731,N_14140,N_14565);
nand U18732 (N_18732,N_14211,N_14023);
nand U18733 (N_18733,N_14356,N_14279);
nor U18734 (N_18734,N_11367,N_13098);
nor U18735 (N_18735,N_11130,N_13260);
nand U18736 (N_18736,N_11349,N_11052);
or U18737 (N_18737,N_10392,N_12087);
or U18738 (N_18738,N_14170,N_11778);
and U18739 (N_18739,N_11355,N_10631);
or U18740 (N_18740,N_12664,N_11511);
and U18741 (N_18741,N_10749,N_13057);
nand U18742 (N_18742,N_14075,N_11999);
or U18743 (N_18743,N_11912,N_11975);
or U18744 (N_18744,N_12951,N_13879);
nor U18745 (N_18745,N_12745,N_10491);
nor U18746 (N_18746,N_14100,N_13588);
nand U18747 (N_18747,N_14282,N_10141);
nor U18748 (N_18748,N_13247,N_13813);
nor U18749 (N_18749,N_10538,N_12808);
or U18750 (N_18750,N_13890,N_14478);
and U18751 (N_18751,N_11535,N_14660);
nor U18752 (N_18752,N_13171,N_10315);
nand U18753 (N_18753,N_13353,N_12303);
and U18754 (N_18754,N_13850,N_10003);
nor U18755 (N_18755,N_12296,N_10798);
nand U18756 (N_18756,N_14429,N_11824);
nor U18757 (N_18757,N_14149,N_14854);
nand U18758 (N_18758,N_12544,N_11621);
or U18759 (N_18759,N_11589,N_10215);
or U18760 (N_18760,N_12199,N_14333);
or U18761 (N_18761,N_14340,N_13623);
or U18762 (N_18762,N_13812,N_12519);
nand U18763 (N_18763,N_14125,N_11172);
or U18764 (N_18764,N_11630,N_10691);
nor U18765 (N_18765,N_10939,N_13510);
nand U18766 (N_18766,N_12251,N_11697);
or U18767 (N_18767,N_12530,N_11368);
and U18768 (N_18768,N_14428,N_13330);
nor U18769 (N_18769,N_11995,N_12895);
nor U18770 (N_18770,N_13408,N_12924);
and U18771 (N_18771,N_14595,N_12660);
nand U18772 (N_18772,N_11381,N_13587);
nor U18773 (N_18773,N_12938,N_14435);
nand U18774 (N_18774,N_12107,N_11584);
and U18775 (N_18775,N_11715,N_11228);
and U18776 (N_18776,N_11986,N_10256);
nand U18777 (N_18777,N_13214,N_11459);
or U18778 (N_18778,N_11627,N_11658);
or U18779 (N_18779,N_14336,N_10974);
or U18780 (N_18780,N_14322,N_13857);
nand U18781 (N_18781,N_14015,N_12177);
nand U18782 (N_18782,N_14940,N_13608);
nor U18783 (N_18783,N_12038,N_10347);
nand U18784 (N_18784,N_13168,N_13073);
and U18785 (N_18785,N_12666,N_12874);
and U18786 (N_18786,N_13242,N_10389);
xnor U18787 (N_18787,N_13570,N_13402);
and U18788 (N_18788,N_13734,N_10563);
or U18789 (N_18789,N_13757,N_14702);
and U18790 (N_18790,N_13770,N_14148);
nand U18791 (N_18791,N_10506,N_12243);
nor U18792 (N_18792,N_10266,N_13625);
nand U18793 (N_18793,N_12386,N_13269);
nor U18794 (N_18794,N_11240,N_13706);
nor U18795 (N_18795,N_13272,N_11754);
nor U18796 (N_18796,N_13254,N_12422);
or U18797 (N_18797,N_14857,N_10360);
and U18798 (N_18798,N_10601,N_12267);
and U18799 (N_18799,N_11627,N_13378);
nor U18800 (N_18800,N_13975,N_11125);
nand U18801 (N_18801,N_13160,N_10170);
nor U18802 (N_18802,N_13040,N_14444);
and U18803 (N_18803,N_13093,N_11151);
nand U18804 (N_18804,N_10089,N_12829);
or U18805 (N_18805,N_11229,N_12117);
nor U18806 (N_18806,N_13856,N_13806);
nor U18807 (N_18807,N_11157,N_10758);
or U18808 (N_18808,N_14302,N_11793);
and U18809 (N_18809,N_10344,N_14317);
nand U18810 (N_18810,N_12929,N_14513);
nor U18811 (N_18811,N_10773,N_12357);
or U18812 (N_18812,N_14336,N_11495);
or U18813 (N_18813,N_13025,N_11807);
nor U18814 (N_18814,N_14503,N_14230);
xnor U18815 (N_18815,N_14762,N_13986);
or U18816 (N_18816,N_13038,N_10308);
or U18817 (N_18817,N_10441,N_10155);
nor U18818 (N_18818,N_10585,N_11201);
nand U18819 (N_18819,N_12181,N_14573);
and U18820 (N_18820,N_13301,N_13531);
nand U18821 (N_18821,N_14247,N_10175);
and U18822 (N_18822,N_11117,N_14790);
nand U18823 (N_18823,N_11485,N_10539);
or U18824 (N_18824,N_13108,N_14031);
or U18825 (N_18825,N_13249,N_13362);
and U18826 (N_18826,N_11371,N_14837);
nand U18827 (N_18827,N_13189,N_13977);
nor U18828 (N_18828,N_12578,N_11918);
or U18829 (N_18829,N_14073,N_13221);
or U18830 (N_18830,N_13620,N_10605);
nand U18831 (N_18831,N_13144,N_11240);
nor U18832 (N_18832,N_13699,N_11675);
and U18833 (N_18833,N_11552,N_14751);
nand U18834 (N_18834,N_12781,N_12542);
and U18835 (N_18835,N_10117,N_13393);
nand U18836 (N_18836,N_14564,N_13839);
or U18837 (N_18837,N_11970,N_14944);
or U18838 (N_18838,N_11615,N_12337);
nand U18839 (N_18839,N_12549,N_10940);
and U18840 (N_18840,N_10585,N_14884);
and U18841 (N_18841,N_10297,N_13503);
nand U18842 (N_18842,N_13689,N_13652);
or U18843 (N_18843,N_11221,N_14474);
or U18844 (N_18844,N_13708,N_11161);
nor U18845 (N_18845,N_14081,N_11528);
nand U18846 (N_18846,N_12256,N_12748);
nor U18847 (N_18847,N_14084,N_10536);
nand U18848 (N_18848,N_10407,N_12026);
nand U18849 (N_18849,N_12952,N_12525);
or U18850 (N_18850,N_14908,N_12953);
or U18851 (N_18851,N_14356,N_13953);
nand U18852 (N_18852,N_11090,N_10350);
or U18853 (N_18853,N_13177,N_14932);
and U18854 (N_18854,N_13698,N_13043);
or U18855 (N_18855,N_10655,N_13317);
and U18856 (N_18856,N_11080,N_12681);
nor U18857 (N_18857,N_10100,N_11582);
nor U18858 (N_18858,N_12661,N_10667);
and U18859 (N_18859,N_10358,N_13358);
nand U18860 (N_18860,N_12590,N_14210);
or U18861 (N_18861,N_12463,N_14115);
or U18862 (N_18862,N_13262,N_13644);
or U18863 (N_18863,N_12762,N_14901);
nand U18864 (N_18864,N_13567,N_13878);
or U18865 (N_18865,N_14344,N_12728);
nand U18866 (N_18866,N_11823,N_10119);
or U18867 (N_18867,N_13605,N_13563);
or U18868 (N_18868,N_13233,N_10729);
or U18869 (N_18869,N_14924,N_12880);
or U18870 (N_18870,N_10991,N_14358);
nor U18871 (N_18871,N_10092,N_11752);
nor U18872 (N_18872,N_10088,N_10470);
or U18873 (N_18873,N_12687,N_10508);
nor U18874 (N_18874,N_14796,N_13179);
nand U18875 (N_18875,N_11731,N_12033);
nand U18876 (N_18876,N_13247,N_14423);
nor U18877 (N_18877,N_13000,N_10496);
and U18878 (N_18878,N_13324,N_12326);
and U18879 (N_18879,N_14640,N_10606);
nand U18880 (N_18880,N_14154,N_12594);
nor U18881 (N_18881,N_10403,N_12692);
or U18882 (N_18882,N_13222,N_12242);
and U18883 (N_18883,N_11166,N_10343);
or U18884 (N_18884,N_10463,N_13943);
nor U18885 (N_18885,N_12101,N_14348);
nand U18886 (N_18886,N_10121,N_13520);
and U18887 (N_18887,N_10173,N_11194);
or U18888 (N_18888,N_14707,N_12707);
nor U18889 (N_18889,N_13962,N_11891);
xnor U18890 (N_18890,N_13033,N_11884);
or U18891 (N_18891,N_14305,N_10418);
nor U18892 (N_18892,N_12779,N_11547);
nor U18893 (N_18893,N_11894,N_12623);
nand U18894 (N_18894,N_10860,N_12928);
and U18895 (N_18895,N_12389,N_14025);
nand U18896 (N_18896,N_13525,N_13860);
or U18897 (N_18897,N_14782,N_13144);
or U18898 (N_18898,N_13501,N_11503);
and U18899 (N_18899,N_14278,N_12067);
or U18900 (N_18900,N_13260,N_10723);
or U18901 (N_18901,N_14745,N_13582);
nor U18902 (N_18902,N_14330,N_14896);
and U18903 (N_18903,N_12963,N_13381);
xor U18904 (N_18904,N_10025,N_14344);
and U18905 (N_18905,N_12024,N_10531);
or U18906 (N_18906,N_12929,N_12662);
and U18907 (N_18907,N_14882,N_11817);
or U18908 (N_18908,N_14993,N_10407);
nor U18909 (N_18909,N_11663,N_14211);
nor U18910 (N_18910,N_11226,N_12349);
nand U18911 (N_18911,N_14407,N_11571);
nand U18912 (N_18912,N_14499,N_14179);
or U18913 (N_18913,N_11900,N_12161);
or U18914 (N_18914,N_11603,N_10918);
nor U18915 (N_18915,N_14766,N_14444);
nand U18916 (N_18916,N_14474,N_10417);
nand U18917 (N_18917,N_13181,N_12663);
nor U18918 (N_18918,N_11602,N_14929);
nand U18919 (N_18919,N_13977,N_10636);
or U18920 (N_18920,N_10158,N_13293);
and U18921 (N_18921,N_14485,N_14355);
nand U18922 (N_18922,N_12879,N_11167);
nor U18923 (N_18923,N_12299,N_11427);
and U18924 (N_18924,N_10420,N_12980);
or U18925 (N_18925,N_10487,N_14145);
nand U18926 (N_18926,N_10734,N_10391);
nor U18927 (N_18927,N_11171,N_12768);
or U18928 (N_18928,N_11996,N_10754);
nand U18929 (N_18929,N_11026,N_12118);
nor U18930 (N_18930,N_12689,N_10415);
nor U18931 (N_18931,N_12640,N_14040);
and U18932 (N_18932,N_10123,N_12318);
or U18933 (N_18933,N_12216,N_10777);
or U18934 (N_18934,N_11082,N_14381);
nor U18935 (N_18935,N_12763,N_12145);
and U18936 (N_18936,N_14992,N_14955);
nand U18937 (N_18937,N_13623,N_11246);
nor U18938 (N_18938,N_11424,N_13489);
and U18939 (N_18939,N_10958,N_13858);
and U18940 (N_18940,N_14016,N_12253);
nor U18941 (N_18941,N_12451,N_13306);
and U18942 (N_18942,N_13970,N_10975);
nand U18943 (N_18943,N_14972,N_10508);
and U18944 (N_18944,N_13256,N_13985);
nand U18945 (N_18945,N_10879,N_14790);
or U18946 (N_18946,N_11341,N_10387);
nand U18947 (N_18947,N_10118,N_11150);
and U18948 (N_18948,N_13076,N_10460);
or U18949 (N_18949,N_11079,N_14826);
nand U18950 (N_18950,N_14025,N_14421);
or U18951 (N_18951,N_14827,N_13860);
nor U18952 (N_18952,N_11704,N_12166);
or U18953 (N_18953,N_12085,N_10766);
and U18954 (N_18954,N_13272,N_13626);
nor U18955 (N_18955,N_12260,N_10696);
and U18956 (N_18956,N_11188,N_14811);
nor U18957 (N_18957,N_12898,N_13739);
and U18958 (N_18958,N_14907,N_12230);
nand U18959 (N_18959,N_13126,N_12633);
nand U18960 (N_18960,N_12711,N_10864);
or U18961 (N_18961,N_12193,N_14183);
nand U18962 (N_18962,N_10140,N_12045);
and U18963 (N_18963,N_11352,N_10982);
or U18964 (N_18964,N_12995,N_11891);
and U18965 (N_18965,N_12901,N_12218);
or U18966 (N_18966,N_10782,N_12746);
or U18967 (N_18967,N_11782,N_14551);
nor U18968 (N_18968,N_14125,N_10246);
nand U18969 (N_18969,N_11711,N_14780);
nand U18970 (N_18970,N_14982,N_10616);
nand U18971 (N_18971,N_10853,N_10002);
and U18972 (N_18972,N_12646,N_12036);
and U18973 (N_18973,N_13563,N_12262);
or U18974 (N_18974,N_12155,N_10364);
nand U18975 (N_18975,N_14040,N_11723);
nor U18976 (N_18976,N_10038,N_14501);
nand U18977 (N_18977,N_14441,N_13090);
nand U18978 (N_18978,N_10271,N_11090);
nor U18979 (N_18979,N_14570,N_10032);
and U18980 (N_18980,N_13054,N_12375);
nand U18981 (N_18981,N_11865,N_13857);
or U18982 (N_18982,N_14158,N_11119);
nand U18983 (N_18983,N_14088,N_13050);
nor U18984 (N_18984,N_14123,N_10609);
and U18985 (N_18985,N_10536,N_11493);
nor U18986 (N_18986,N_10328,N_14454);
or U18987 (N_18987,N_13766,N_12853);
and U18988 (N_18988,N_12752,N_13146);
nor U18989 (N_18989,N_12330,N_14437);
and U18990 (N_18990,N_13294,N_14421);
or U18991 (N_18991,N_14956,N_14996);
nor U18992 (N_18992,N_11908,N_11089);
nor U18993 (N_18993,N_11988,N_13834);
or U18994 (N_18994,N_14032,N_11568);
or U18995 (N_18995,N_11929,N_13700);
and U18996 (N_18996,N_10273,N_11886);
or U18997 (N_18997,N_10361,N_12181);
xor U18998 (N_18998,N_10430,N_13850);
or U18999 (N_18999,N_14449,N_10452);
nor U19000 (N_19000,N_14801,N_13623);
or U19001 (N_19001,N_14591,N_11195);
or U19002 (N_19002,N_12997,N_10311);
nand U19003 (N_19003,N_14451,N_12057);
and U19004 (N_19004,N_13701,N_14724);
nand U19005 (N_19005,N_14644,N_10506);
nor U19006 (N_19006,N_10975,N_14014);
and U19007 (N_19007,N_10402,N_13024);
xnor U19008 (N_19008,N_14832,N_11819);
or U19009 (N_19009,N_12326,N_12609);
or U19010 (N_19010,N_13546,N_12303);
or U19011 (N_19011,N_10200,N_11867);
nor U19012 (N_19012,N_12658,N_11051);
nand U19013 (N_19013,N_12019,N_11590);
and U19014 (N_19014,N_14451,N_11765);
nor U19015 (N_19015,N_14458,N_14733);
and U19016 (N_19016,N_14112,N_10780);
nor U19017 (N_19017,N_10609,N_13760);
or U19018 (N_19018,N_11780,N_14796);
nor U19019 (N_19019,N_11732,N_12525);
and U19020 (N_19020,N_14217,N_14110);
nor U19021 (N_19021,N_13782,N_11789);
or U19022 (N_19022,N_13987,N_13829);
nand U19023 (N_19023,N_13845,N_13586);
nand U19024 (N_19024,N_10907,N_13960);
or U19025 (N_19025,N_11121,N_12141);
and U19026 (N_19026,N_14642,N_12592);
nand U19027 (N_19027,N_13695,N_11362);
and U19028 (N_19028,N_10699,N_10945);
nand U19029 (N_19029,N_13479,N_11515);
nand U19030 (N_19030,N_13811,N_12960);
or U19031 (N_19031,N_12880,N_11441);
nand U19032 (N_19032,N_14582,N_10794);
and U19033 (N_19033,N_13293,N_11378);
or U19034 (N_19034,N_12873,N_13989);
nor U19035 (N_19035,N_14345,N_14967);
and U19036 (N_19036,N_14892,N_12663);
and U19037 (N_19037,N_10466,N_12051);
nor U19038 (N_19038,N_13162,N_10782);
and U19039 (N_19039,N_10585,N_14466);
nand U19040 (N_19040,N_11246,N_14735);
nor U19041 (N_19041,N_10735,N_11008);
or U19042 (N_19042,N_14351,N_10139);
or U19043 (N_19043,N_13035,N_11183);
nor U19044 (N_19044,N_12091,N_11942);
nor U19045 (N_19045,N_12465,N_11175);
nand U19046 (N_19046,N_10720,N_11104);
or U19047 (N_19047,N_13896,N_10877);
nor U19048 (N_19048,N_13932,N_14922);
nand U19049 (N_19049,N_14381,N_13490);
nand U19050 (N_19050,N_12106,N_10596);
nor U19051 (N_19051,N_13477,N_13463);
or U19052 (N_19052,N_11220,N_14399);
and U19053 (N_19053,N_13576,N_13308);
or U19054 (N_19054,N_11792,N_13529);
and U19055 (N_19055,N_11335,N_14676);
nand U19056 (N_19056,N_13256,N_14343);
nor U19057 (N_19057,N_13259,N_13482);
nor U19058 (N_19058,N_11033,N_12720);
nor U19059 (N_19059,N_11646,N_14678);
and U19060 (N_19060,N_10608,N_14886);
nor U19061 (N_19061,N_14670,N_12684);
or U19062 (N_19062,N_11222,N_12737);
and U19063 (N_19063,N_14193,N_13155);
and U19064 (N_19064,N_11767,N_10522);
and U19065 (N_19065,N_13951,N_11136);
nand U19066 (N_19066,N_11828,N_14407);
or U19067 (N_19067,N_10759,N_10127);
and U19068 (N_19068,N_10196,N_14636);
or U19069 (N_19069,N_14253,N_14931);
nand U19070 (N_19070,N_12934,N_14416);
and U19071 (N_19071,N_10824,N_14562);
or U19072 (N_19072,N_12778,N_12884);
nand U19073 (N_19073,N_12682,N_13248);
or U19074 (N_19074,N_10123,N_10860);
nor U19075 (N_19075,N_12205,N_12565);
and U19076 (N_19076,N_12906,N_12805);
nand U19077 (N_19077,N_14750,N_14649);
nor U19078 (N_19078,N_12623,N_11505);
and U19079 (N_19079,N_14366,N_12826);
and U19080 (N_19080,N_11209,N_12484);
nand U19081 (N_19081,N_12063,N_10496);
nor U19082 (N_19082,N_11004,N_11225);
nand U19083 (N_19083,N_14999,N_14936);
nand U19084 (N_19084,N_11111,N_12663);
nor U19085 (N_19085,N_13592,N_10714);
or U19086 (N_19086,N_14713,N_13069);
or U19087 (N_19087,N_12860,N_12653);
nor U19088 (N_19088,N_14690,N_11029);
nand U19089 (N_19089,N_11279,N_14685);
and U19090 (N_19090,N_13578,N_10583);
nand U19091 (N_19091,N_14668,N_10385);
or U19092 (N_19092,N_12165,N_13645);
nand U19093 (N_19093,N_10060,N_13551);
or U19094 (N_19094,N_10591,N_11619);
nor U19095 (N_19095,N_14605,N_12979);
and U19096 (N_19096,N_11655,N_14951);
or U19097 (N_19097,N_13507,N_13176);
nor U19098 (N_19098,N_12858,N_11728);
nor U19099 (N_19099,N_14948,N_13428);
or U19100 (N_19100,N_14792,N_14859);
nand U19101 (N_19101,N_14172,N_13125);
nor U19102 (N_19102,N_13284,N_13168);
xnor U19103 (N_19103,N_12710,N_12222);
or U19104 (N_19104,N_11753,N_13784);
nor U19105 (N_19105,N_14246,N_14256);
and U19106 (N_19106,N_11547,N_12985);
and U19107 (N_19107,N_13742,N_14128);
and U19108 (N_19108,N_12270,N_10748);
or U19109 (N_19109,N_10999,N_13542);
nor U19110 (N_19110,N_12450,N_12999);
nor U19111 (N_19111,N_10838,N_10105);
and U19112 (N_19112,N_13785,N_14875);
nand U19113 (N_19113,N_12098,N_13871);
or U19114 (N_19114,N_13076,N_14327);
and U19115 (N_19115,N_13802,N_13009);
nand U19116 (N_19116,N_14492,N_10448);
nand U19117 (N_19117,N_12617,N_12471);
and U19118 (N_19118,N_12678,N_10369);
and U19119 (N_19119,N_13287,N_13164);
nand U19120 (N_19120,N_13239,N_10469);
and U19121 (N_19121,N_10932,N_10584);
nand U19122 (N_19122,N_11016,N_13460);
nor U19123 (N_19123,N_10109,N_13334);
nand U19124 (N_19124,N_10051,N_10717);
nand U19125 (N_19125,N_10311,N_12877);
or U19126 (N_19126,N_11775,N_10012);
nand U19127 (N_19127,N_14057,N_13601);
and U19128 (N_19128,N_11652,N_10106);
and U19129 (N_19129,N_10709,N_11427);
nor U19130 (N_19130,N_14167,N_14735);
or U19131 (N_19131,N_10620,N_13690);
nor U19132 (N_19132,N_11980,N_14150);
and U19133 (N_19133,N_13157,N_11867);
or U19134 (N_19134,N_14729,N_11125);
nor U19135 (N_19135,N_14126,N_11601);
nand U19136 (N_19136,N_14668,N_13288);
nor U19137 (N_19137,N_13706,N_12404);
nand U19138 (N_19138,N_11414,N_10529);
nand U19139 (N_19139,N_13267,N_12362);
and U19140 (N_19140,N_13254,N_13136);
nor U19141 (N_19141,N_11332,N_11602);
or U19142 (N_19142,N_13973,N_13361);
nor U19143 (N_19143,N_13908,N_12254);
and U19144 (N_19144,N_10017,N_12953);
nand U19145 (N_19145,N_13504,N_12184);
or U19146 (N_19146,N_12677,N_14301);
or U19147 (N_19147,N_14005,N_10717);
nor U19148 (N_19148,N_10283,N_12698);
or U19149 (N_19149,N_11409,N_10681);
and U19150 (N_19150,N_12245,N_13988);
or U19151 (N_19151,N_11697,N_13700);
or U19152 (N_19152,N_10841,N_14769);
nand U19153 (N_19153,N_10670,N_11467);
nand U19154 (N_19154,N_10696,N_13827);
and U19155 (N_19155,N_13065,N_14620);
nand U19156 (N_19156,N_10241,N_10539);
nand U19157 (N_19157,N_11042,N_13222);
or U19158 (N_19158,N_11625,N_11459);
nor U19159 (N_19159,N_12910,N_14517);
nor U19160 (N_19160,N_10124,N_14608);
or U19161 (N_19161,N_10838,N_11814);
nor U19162 (N_19162,N_11797,N_12587);
nor U19163 (N_19163,N_14741,N_10731);
nor U19164 (N_19164,N_13881,N_10966);
nor U19165 (N_19165,N_13322,N_14353);
and U19166 (N_19166,N_13618,N_12745);
nand U19167 (N_19167,N_12874,N_13167);
nand U19168 (N_19168,N_14035,N_10642);
nor U19169 (N_19169,N_10215,N_11703);
and U19170 (N_19170,N_14073,N_12364);
or U19171 (N_19171,N_11040,N_11097);
and U19172 (N_19172,N_10906,N_12063);
nor U19173 (N_19173,N_11403,N_13051);
or U19174 (N_19174,N_14424,N_14718);
and U19175 (N_19175,N_14072,N_14275);
or U19176 (N_19176,N_11834,N_14716);
and U19177 (N_19177,N_11917,N_14986);
or U19178 (N_19178,N_11351,N_12220);
nand U19179 (N_19179,N_14339,N_14441);
and U19180 (N_19180,N_14060,N_11913);
nand U19181 (N_19181,N_13090,N_12528);
nand U19182 (N_19182,N_14379,N_12146);
or U19183 (N_19183,N_14150,N_12664);
and U19184 (N_19184,N_14549,N_14945);
and U19185 (N_19185,N_13288,N_14453);
and U19186 (N_19186,N_10480,N_12665);
and U19187 (N_19187,N_14720,N_14971);
nor U19188 (N_19188,N_11436,N_12721);
or U19189 (N_19189,N_12100,N_10564);
or U19190 (N_19190,N_12095,N_11894);
and U19191 (N_19191,N_10111,N_10208);
or U19192 (N_19192,N_12982,N_12611);
xnor U19193 (N_19193,N_10392,N_10908);
nand U19194 (N_19194,N_14959,N_13671);
nand U19195 (N_19195,N_12357,N_14746);
nand U19196 (N_19196,N_13795,N_14301);
nor U19197 (N_19197,N_13604,N_14246);
or U19198 (N_19198,N_10417,N_11687);
nand U19199 (N_19199,N_11655,N_14317);
nor U19200 (N_19200,N_12515,N_13687);
nor U19201 (N_19201,N_11272,N_14124);
nand U19202 (N_19202,N_11084,N_12048);
nor U19203 (N_19203,N_10336,N_14653);
nor U19204 (N_19204,N_12970,N_11353);
or U19205 (N_19205,N_12683,N_12573);
nand U19206 (N_19206,N_10434,N_14202);
nor U19207 (N_19207,N_12988,N_10482);
or U19208 (N_19208,N_14671,N_10041);
nor U19209 (N_19209,N_13131,N_14646);
nor U19210 (N_19210,N_10407,N_13455);
or U19211 (N_19211,N_12025,N_11449);
and U19212 (N_19212,N_13755,N_11761);
nand U19213 (N_19213,N_13811,N_12258);
and U19214 (N_19214,N_11562,N_12876);
nand U19215 (N_19215,N_11098,N_10188);
and U19216 (N_19216,N_11226,N_11360);
nor U19217 (N_19217,N_14958,N_12775);
nor U19218 (N_19218,N_13080,N_12193);
or U19219 (N_19219,N_10558,N_10637);
and U19220 (N_19220,N_10192,N_13922);
or U19221 (N_19221,N_13357,N_10371);
or U19222 (N_19222,N_14029,N_10496);
and U19223 (N_19223,N_12442,N_12540);
nand U19224 (N_19224,N_10697,N_13818);
or U19225 (N_19225,N_10387,N_11320);
nor U19226 (N_19226,N_10544,N_14801);
nor U19227 (N_19227,N_12973,N_11467);
nor U19228 (N_19228,N_14941,N_12806);
or U19229 (N_19229,N_10485,N_10834);
nand U19230 (N_19230,N_11188,N_10365);
or U19231 (N_19231,N_13607,N_11956);
nand U19232 (N_19232,N_13463,N_13693);
nand U19233 (N_19233,N_13758,N_11128);
or U19234 (N_19234,N_14497,N_14030);
and U19235 (N_19235,N_12632,N_14281);
nor U19236 (N_19236,N_11672,N_11234);
nand U19237 (N_19237,N_14045,N_12795);
or U19238 (N_19238,N_11633,N_11855);
or U19239 (N_19239,N_13942,N_13680);
or U19240 (N_19240,N_13914,N_12417);
and U19241 (N_19241,N_14444,N_14581);
nor U19242 (N_19242,N_10562,N_14614);
or U19243 (N_19243,N_11727,N_14380);
nand U19244 (N_19244,N_12581,N_10245);
nand U19245 (N_19245,N_11395,N_11090);
and U19246 (N_19246,N_13483,N_10222);
nand U19247 (N_19247,N_12088,N_10310);
nand U19248 (N_19248,N_12511,N_10522);
nand U19249 (N_19249,N_12578,N_13591);
nand U19250 (N_19250,N_14363,N_11888);
or U19251 (N_19251,N_13375,N_13078);
or U19252 (N_19252,N_11953,N_12972);
nor U19253 (N_19253,N_14673,N_14335);
or U19254 (N_19254,N_14192,N_12096);
nor U19255 (N_19255,N_10311,N_13903);
nand U19256 (N_19256,N_13575,N_13496);
and U19257 (N_19257,N_13255,N_12864);
nand U19258 (N_19258,N_11160,N_13614);
nand U19259 (N_19259,N_11660,N_12718);
and U19260 (N_19260,N_14722,N_14270);
or U19261 (N_19261,N_12357,N_12838);
and U19262 (N_19262,N_13867,N_12123);
nor U19263 (N_19263,N_13843,N_13343);
and U19264 (N_19264,N_13754,N_11811);
nor U19265 (N_19265,N_14508,N_11911);
nand U19266 (N_19266,N_10674,N_14039);
nor U19267 (N_19267,N_11750,N_13836);
nor U19268 (N_19268,N_14756,N_13279);
nand U19269 (N_19269,N_12531,N_11427);
or U19270 (N_19270,N_13789,N_14585);
nand U19271 (N_19271,N_12917,N_14280);
nand U19272 (N_19272,N_13541,N_14145);
and U19273 (N_19273,N_12521,N_10387);
or U19274 (N_19274,N_11390,N_11059);
nor U19275 (N_19275,N_14589,N_10727);
nor U19276 (N_19276,N_10888,N_12410);
and U19277 (N_19277,N_10892,N_10092);
or U19278 (N_19278,N_11471,N_10617);
nor U19279 (N_19279,N_11454,N_13032);
nor U19280 (N_19280,N_12826,N_10139);
nand U19281 (N_19281,N_10327,N_10363);
or U19282 (N_19282,N_11281,N_13949);
nand U19283 (N_19283,N_13428,N_13762);
and U19284 (N_19284,N_10274,N_12478);
nor U19285 (N_19285,N_13967,N_14802);
nor U19286 (N_19286,N_12894,N_13411);
or U19287 (N_19287,N_11491,N_12761);
nand U19288 (N_19288,N_13902,N_12650);
or U19289 (N_19289,N_13603,N_11356);
or U19290 (N_19290,N_13464,N_13069);
and U19291 (N_19291,N_13498,N_12336);
or U19292 (N_19292,N_11746,N_14221);
or U19293 (N_19293,N_10154,N_10710);
xor U19294 (N_19294,N_11495,N_11602);
nor U19295 (N_19295,N_14055,N_13533);
and U19296 (N_19296,N_12735,N_11125);
or U19297 (N_19297,N_14696,N_14049);
nand U19298 (N_19298,N_13163,N_14620);
nand U19299 (N_19299,N_13043,N_10088);
and U19300 (N_19300,N_12308,N_10952);
nor U19301 (N_19301,N_13634,N_10926);
nor U19302 (N_19302,N_12204,N_10689);
nor U19303 (N_19303,N_10735,N_14162);
and U19304 (N_19304,N_11590,N_13474);
and U19305 (N_19305,N_11039,N_12980);
and U19306 (N_19306,N_13078,N_10531);
nor U19307 (N_19307,N_10333,N_14098);
nor U19308 (N_19308,N_14709,N_14193);
nand U19309 (N_19309,N_10571,N_14516);
nor U19310 (N_19310,N_12001,N_11128);
and U19311 (N_19311,N_13480,N_10878);
nor U19312 (N_19312,N_11064,N_11252);
nand U19313 (N_19313,N_13349,N_12559);
or U19314 (N_19314,N_12179,N_12739);
nor U19315 (N_19315,N_14963,N_14326);
or U19316 (N_19316,N_11135,N_10637);
and U19317 (N_19317,N_12211,N_13790);
nand U19318 (N_19318,N_11092,N_12117);
or U19319 (N_19319,N_11484,N_13477);
nand U19320 (N_19320,N_11714,N_12984);
and U19321 (N_19321,N_13055,N_12466);
nor U19322 (N_19322,N_14614,N_11628);
nand U19323 (N_19323,N_10104,N_13422);
and U19324 (N_19324,N_10284,N_14217);
or U19325 (N_19325,N_11084,N_10736);
nand U19326 (N_19326,N_11097,N_14622);
and U19327 (N_19327,N_13420,N_10871);
or U19328 (N_19328,N_12633,N_12453);
nor U19329 (N_19329,N_14651,N_13963);
and U19330 (N_19330,N_12461,N_10608);
nor U19331 (N_19331,N_11940,N_12076);
nand U19332 (N_19332,N_11480,N_12305);
or U19333 (N_19333,N_11415,N_10689);
and U19334 (N_19334,N_12619,N_11787);
or U19335 (N_19335,N_12250,N_12984);
or U19336 (N_19336,N_11416,N_13254);
nand U19337 (N_19337,N_14936,N_14818);
and U19338 (N_19338,N_12785,N_11301);
nor U19339 (N_19339,N_13526,N_10751);
or U19340 (N_19340,N_10130,N_12971);
or U19341 (N_19341,N_11605,N_11360);
and U19342 (N_19342,N_11352,N_11323);
nor U19343 (N_19343,N_10230,N_12744);
nor U19344 (N_19344,N_12546,N_12432);
or U19345 (N_19345,N_12787,N_11663);
nand U19346 (N_19346,N_10538,N_10937);
or U19347 (N_19347,N_14507,N_12280);
or U19348 (N_19348,N_14050,N_14645);
and U19349 (N_19349,N_12356,N_13446);
nor U19350 (N_19350,N_12012,N_12606);
or U19351 (N_19351,N_12414,N_12726);
nand U19352 (N_19352,N_14756,N_14332);
nand U19353 (N_19353,N_10353,N_12207);
nor U19354 (N_19354,N_10183,N_12709);
or U19355 (N_19355,N_10742,N_11214);
and U19356 (N_19356,N_12042,N_10218);
nor U19357 (N_19357,N_14319,N_12368);
or U19358 (N_19358,N_14260,N_13234);
nand U19359 (N_19359,N_14734,N_12690);
nand U19360 (N_19360,N_14898,N_14749);
nand U19361 (N_19361,N_14641,N_14436);
nand U19362 (N_19362,N_11913,N_10646);
or U19363 (N_19363,N_14051,N_13215);
nand U19364 (N_19364,N_14251,N_11017);
and U19365 (N_19365,N_13967,N_10985);
or U19366 (N_19366,N_10110,N_12563);
or U19367 (N_19367,N_14998,N_14959);
or U19368 (N_19368,N_10151,N_10399);
nor U19369 (N_19369,N_11926,N_12222);
nand U19370 (N_19370,N_14080,N_10750);
or U19371 (N_19371,N_10215,N_10770);
or U19372 (N_19372,N_13428,N_11856);
nand U19373 (N_19373,N_13838,N_14585);
nand U19374 (N_19374,N_12683,N_10354);
or U19375 (N_19375,N_14151,N_11604);
and U19376 (N_19376,N_11702,N_13351);
nor U19377 (N_19377,N_13608,N_14886);
and U19378 (N_19378,N_13927,N_12886);
nor U19379 (N_19379,N_14843,N_10255);
and U19380 (N_19380,N_10212,N_13184);
nand U19381 (N_19381,N_12140,N_10714);
nand U19382 (N_19382,N_11775,N_14244);
nor U19383 (N_19383,N_11746,N_11104);
or U19384 (N_19384,N_10615,N_10273);
nor U19385 (N_19385,N_11915,N_11396);
nand U19386 (N_19386,N_12753,N_11329);
or U19387 (N_19387,N_13065,N_14580);
nor U19388 (N_19388,N_10059,N_14477);
nor U19389 (N_19389,N_13902,N_13230);
nor U19390 (N_19390,N_10030,N_13930);
or U19391 (N_19391,N_11345,N_14218);
nand U19392 (N_19392,N_11896,N_12518);
or U19393 (N_19393,N_12430,N_11452);
or U19394 (N_19394,N_10766,N_10733);
nor U19395 (N_19395,N_14821,N_13684);
and U19396 (N_19396,N_12590,N_12050);
nand U19397 (N_19397,N_10403,N_10338);
nand U19398 (N_19398,N_14055,N_14863);
and U19399 (N_19399,N_14809,N_14693);
nor U19400 (N_19400,N_10318,N_10071);
and U19401 (N_19401,N_11703,N_10102);
nor U19402 (N_19402,N_13270,N_10759);
or U19403 (N_19403,N_12555,N_11402);
nor U19404 (N_19404,N_14705,N_14866);
and U19405 (N_19405,N_14109,N_14338);
nor U19406 (N_19406,N_13333,N_13357);
nand U19407 (N_19407,N_13254,N_10180);
nand U19408 (N_19408,N_11258,N_12602);
and U19409 (N_19409,N_13152,N_11886);
nand U19410 (N_19410,N_14036,N_14867);
and U19411 (N_19411,N_13180,N_13617);
and U19412 (N_19412,N_13758,N_13794);
and U19413 (N_19413,N_13131,N_12174);
nor U19414 (N_19414,N_11734,N_11874);
or U19415 (N_19415,N_14142,N_13895);
or U19416 (N_19416,N_13300,N_12009);
nor U19417 (N_19417,N_11516,N_11181);
or U19418 (N_19418,N_14977,N_10209);
and U19419 (N_19419,N_14325,N_13617);
nor U19420 (N_19420,N_12364,N_14958);
or U19421 (N_19421,N_10299,N_11195);
xor U19422 (N_19422,N_13107,N_13939);
or U19423 (N_19423,N_13398,N_13409);
or U19424 (N_19424,N_11885,N_11425);
nand U19425 (N_19425,N_11137,N_11196);
and U19426 (N_19426,N_13736,N_14219);
nand U19427 (N_19427,N_11013,N_13958);
nand U19428 (N_19428,N_12548,N_10431);
nand U19429 (N_19429,N_14597,N_13764);
or U19430 (N_19430,N_11793,N_12603);
and U19431 (N_19431,N_11183,N_13825);
nor U19432 (N_19432,N_11481,N_14435);
and U19433 (N_19433,N_13104,N_10393);
and U19434 (N_19434,N_11876,N_10494);
or U19435 (N_19435,N_11737,N_14671);
and U19436 (N_19436,N_11661,N_12255);
nand U19437 (N_19437,N_12582,N_10521);
nand U19438 (N_19438,N_10152,N_13260);
nor U19439 (N_19439,N_11200,N_13625);
nand U19440 (N_19440,N_10431,N_11786);
nand U19441 (N_19441,N_12019,N_11879);
and U19442 (N_19442,N_10127,N_10045);
or U19443 (N_19443,N_14091,N_10260);
or U19444 (N_19444,N_10171,N_14133);
or U19445 (N_19445,N_12477,N_14090);
nand U19446 (N_19446,N_13527,N_10802);
and U19447 (N_19447,N_14752,N_13180);
nor U19448 (N_19448,N_13707,N_13747);
nor U19449 (N_19449,N_13210,N_13289);
nor U19450 (N_19450,N_13650,N_14211);
or U19451 (N_19451,N_14371,N_13531);
xnor U19452 (N_19452,N_11431,N_10230);
and U19453 (N_19453,N_11894,N_13482);
and U19454 (N_19454,N_11639,N_12565);
nand U19455 (N_19455,N_10117,N_10214);
and U19456 (N_19456,N_14778,N_13394);
and U19457 (N_19457,N_10005,N_13080);
nor U19458 (N_19458,N_12396,N_10701);
nor U19459 (N_19459,N_10373,N_14230);
nand U19460 (N_19460,N_14044,N_14962);
nor U19461 (N_19461,N_14032,N_11279);
nor U19462 (N_19462,N_14406,N_13908);
and U19463 (N_19463,N_14112,N_13915);
nand U19464 (N_19464,N_11159,N_12954);
and U19465 (N_19465,N_12632,N_14203);
and U19466 (N_19466,N_13044,N_10928);
nand U19467 (N_19467,N_14953,N_12611);
and U19468 (N_19468,N_10549,N_10205);
or U19469 (N_19469,N_14460,N_10110);
or U19470 (N_19470,N_10980,N_11235);
nand U19471 (N_19471,N_11466,N_14464);
and U19472 (N_19472,N_10863,N_12015);
nand U19473 (N_19473,N_14951,N_12963);
nand U19474 (N_19474,N_12356,N_10948);
nand U19475 (N_19475,N_11490,N_10230);
nor U19476 (N_19476,N_12226,N_13079);
or U19477 (N_19477,N_12017,N_11597);
nor U19478 (N_19478,N_11409,N_11093);
nand U19479 (N_19479,N_14703,N_11251);
or U19480 (N_19480,N_13705,N_11698);
and U19481 (N_19481,N_14910,N_12767);
nand U19482 (N_19482,N_14078,N_14922);
nand U19483 (N_19483,N_13261,N_11770);
nand U19484 (N_19484,N_11901,N_13306);
or U19485 (N_19485,N_13732,N_10478);
or U19486 (N_19486,N_12180,N_14230);
nand U19487 (N_19487,N_13374,N_12786);
nor U19488 (N_19488,N_11465,N_10640);
nand U19489 (N_19489,N_14708,N_14500);
or U19490 (N_19490,N_11138,N_14817);
or U19491 (N_19491,N_11143,N_10346);
nor U19492 (N_19492,N_12501,N_10655);
nor U19493 (N_19493,N_10905,N_11354);
nand U19494 (N_19494,N_11160,N_12452);
nor U19495 (N_19495,N_13082,N_14269);
xor U19496 (N_19496,N_14041,N_12273);
and U19497 (N_19497,N_14980,N_11850);
or U19498 (N_19498,N_13280,N_14336);
nor U19499 (N_19499,N_14507,N_11852);
nor U19500 (N_19500,N_13034,N_10106);
nor U19501 (N_19501,N_14806,N_10396);
nor U19502 (N_19502,N_13237,N_11026);
nand U19503 (N_19503,N_12110,N_11703);
nor U19504 (N_19504,N_14412,N_14698);
nor U19505 (N_19505,N_10723,N_10026);
xor U19506 (N_19506,N_10847,N_10792);
nor U19507 (N_19507,N_13519,N_10771);
nor U19508 (N_19508,N_13742,N_12690);
and U19509 (N_19509,N_12314,N_14361);
or U19510 (N_19510,N_11759,N_10915);
nor U19511 (N_19511,N_13534,N_11145);
nand U19512 (N_19512,N_11365,N_12170);
nor U19513 (N_19513,N_10346,N_12998);
nor U19514 (N_19514,N_11350,N_13640);
nor U19515 (N_19515,N_13388,N_13977);
and U19516 (N_19516,N_13550,N_12892);
nor U19517 (N_19517,N_14287,N_12874);
nor U19518 (N_19518,N_12760,N_11817);
or U19519 (N_19519,N_12131,N_12125);
xnor U19520 (N_19520,N_14280,N_12536);
nand U19521 (N_19521,N_13488,N_10014);
nor U19522 (N_19522,N_14422,N_10327);
and U19523 (N_19523,N_14510,N_11183);
and U19524 (N_19524,N_12382,N_13897);
and U19525 (N_19525,N_14725,N_10631);
and U19526 (N_19526,N_13477,N_11690);
and U19527 (N_19527,N_13550,N_12581);
nor U19528 (N_19528,N_10066,N_12019);
nand U19529 (N_19529,N_11034,N_10322);
nor U19530 (N_19530,N_12160,N_14363);
nand U19531 (N_19531,N_13210,N_10443);
nand U19532 (N_19532,N_11457,N_11586);
nand U19533 (N_19533,N_14041,N_12616);
or U19534 (N_19534,N_10841,N_10370);
and U19535 (N_19535,N_14733,N_10226);
or U19536 (N_19536,N_13742,N_11996);
or U19537 (N_19537,N_10599,N_11449);
nand U19538 (N_19538,N_11167,N_14417);
and U19539 (N_19539,N_14699,N_12576);
and U19540 (N_19540,N_13898,N_13581);
nand U19541 (N_19541,N_14250,N_10445);
nand U19542 (N_19542,N_12016,N_13060);
nand U19543 (N_19543,N_13377,N_14331);
nand U19544 (N_19544,N_10450,N_10679);
and U19545 (N_19545,N_12234,N_10061);
nor U19546 (N_19546,N_12194,N_14387);
or U19547 (N_19547,N_12284,N_14269);
nand U19548 (N_19548,N_13392,N_10811);
and U19549 (N_19549,N_10600,N_14946);
nand U19550 (N_19550,N_11197,N_13862);
nor U19551 (N_19551,N_14297,N_11289);
nand U19552 (N_19552,N_10008,N_14361);
and U19553 (N_19553,N_13148,N_14740);
or U19554 (N_19554,N_12831,N_13939);
and U19555 (N_19555,N_14613,N_11369);
and U19556 (N_19556,N_10503,N_11859);
and U19557 (N_19557,N_14895,N_14698);
nor U19558 (N_19558,N_14727,N_12628);
nor U19559 (N_19559,N_13622,N_12130);
and U19560 (N_19560,N_12784,N_11867);
nor U19561 (N_19561,N_12623,N_10512);
or U19562 (N_19562,N_12523,N_13239);
xnor U19563 (N_19563,N_11698,N_10270);
and U19564 (N_19564,N_13851,N_14543);
and U19565 (N_19565,N_11300,N_11000);
and U19566 (N_19566,N_12879,N_11349);
or U19567 (N_19567,N_13760,N_14670);
or U19568 (N_19568,N_12942,N_11365);
or U19569 (N_19569,N_14618,N_12336);
or U19570 (N_19570,N_13506,N_13417);
nor U19571 (N_19571,N_14845,N_11754);
or U19572 (N_19572,N_11624,N_12473);
xor U19573 (N_19573,N_11956,N_12339);
or U19574 (N_19574,N_12941,N_11151);
nand U19575 (N_19575,N_12034,N_13186);
nor U19576 (N_19576,N_14833,N_14528);
nor U19577 (N_19577,N_10305,N_13045);
nor U19578 (N_19578,N_11401,N_12492);
and U19579 (N_19579,N_12469,N_13663);
or U19580 (N_19580,N_12162,N_14575);
or U19581 (N_19581,N_11477,N_10322);
nand U19582 (N_19582,N_14652,N_10103);
nor U19583 (N_19583,N_13154,N_11212);
and U19584 (N_19584,N_11801,N_12840);
nor U19585 (N_19585,N_13773,N_12327);
or U19586 (N_19586,N_10385,N_10509);
nand U19587 (N_19587,N_11237,N_10009);
nor U19588 (N_19588,N_12601,N_14394);
and U19589 (N_19589,N_10469,N_10142);
nand U19590 (N_19590,N_11400,N_10231);
nand U19591 (N_19591,N_12576,N_13967);
nand U19592 (N_19592,N_10736,N_10047);
or U19593 (N_19593,N_10516,N_10624);
nor U19594 (N_19594,N_12020,N_12179);
or U19595 (N_19595,N_12236,N_10139);
nand U19596 (N_19596,N_14809,N_11726);
nor U19597 (N_19597,N_13586,N_13304);
or U19598 (N_19598,N_14953,N_11297);
xnor U19599 (N_19599,N_10822,N_13553);
or U19600 (N_19600,N_10670,N_14692);
and U19601 (N_19601,N_11784,N_10332);
and U19602 (N_19602,N_10409,N_11617);
and U19603 (N_19603,N_14111,N_11598);
nor U19604 (N_19604,N_12702,N_10221);
nor U19605 (N_19605,N_11804,N_12376);
and U19606 (N_19606,N_10156,N_14548);
nand U19607 (N_19607,N_12851,N_14191);
nor U19608 (N_19608,N_13588,N_14804);
or U19609 (N_19609,N_13279,N_12696);
nand U19610 (N_19610,N_11683,N_14590);
and U19611 (N_19611,N_12580,N_13272);
or U19612 (N_19612,N_14015,N_12713);
nand U19613 (N_19613,N_10758,N_11000);
or U19614 (N_19614,N_10314,N_11643);
or U19615 (N_19615,N_10466,N_12057);
or U19616 (N_19616,N_11012,N_13890);
nor U19617 (N_19617,N_14830,N_12413);
nor U19618 (N_19618,N_10261,N_12491);
and U19619 (N_19619,N_12321,N_13992);
or U19620 (N_19620,N_11004,N_10377);
or U19621 (N_19621,N_12818,N_10998);
nor U19622 (N_19622,N_14316,N_14720);
nand U19623 (N_19623,N_11429,N_11202);
nand U19624 (N_19624,N_14030,N_10914);
or U19625 (N_19625,N_10483,N_11787);
or U19626 (N_19626,N_10311,N_11960);
nand U19627 (N_19627,N_10261,N_12610);
nor U19628 (N_19628,N_11190,N_10086);
and U19629 (N_19629,N_12258,N_12609);
and U19630 (N_19630,N_13637,N_11883);
nor U19631 (N_19631,N_14787,N_12179);
and U19632 (N_19632,N_14820,N_11390);
or U19633 (N_19633,N_11908,N_11820);
nor U19634 (N_19634,N_13248,N_11111);
or U19635 (N_19635,N_14810,N_11448);
or U19636 (N_19636,N_11667,N_11977);
or U19637 (N_19637,N_10102,N_14016);
or U19638 (N_19638,N_11440,N_13331);
and U19639 (N_19639,N_12933,N_12505);
nand U19640 (N_19640,N_14084,N_13444);
nand U19641 (N_19641,N_13424,N_12363);
nor U19642 (N_19642,N_12811,N_14855);
nor U19643 (N_19643,N_11264,N_13590);
nor U19644 (N_19644,N_13322,N_14369);
nor U19645 (N_19645,N_10620,N_13437);
nor U19646 (N_19646,N_10496,N_13943);
or U19647 (N_19647,N_10930,N_13752);
nor U19648 (N_19648,N_12354,N_14747);
or U19649 (N_19649,N_12626,N_13169);
nor U19650 (N_19650,N_11538,N_14153);
and U19651 (N_19651,N_14553,N_11317);
and U19652 (N_19652,N_10218,N_12814);
nor U19653 (N_19653,N_14822,N_12247);
or U19654 (N_19654,N_12951,N_11520);
or U19655 (N_19655,N_13775,N_13517);
nor U19656 (N_19656,N_11210,N_11127);
nand U19657 (N_19657,N_13731,N_13689);
nor U19658 (N_19658,N_14280,N_13461);
nand U19659 (N_19659,N_12095,N_14395);
and U19660 (N_19660,N_14142,N_12716);
nand U19661 (N_19661,N_13756,N_14417);
nand U19662 (N_19662,N_14357,N_10403);
nor U19663 (N_19663,N_12094,N_13000);
nand U19664 (N_19664,N_14632,N_14939);
nor U19665 (N_19665,N_11676,N_14551);
and U19666 (N_19666,N_11104,N_13516);
nand U19667 (N_19667,N_10732,N_12370);
nand U19668 (N_19668,N_11532,N_13034);
nor U19669 (N_19669,N_11378,N_13582);
and U19670 (N_19670,N_13409,N_12689);
nor U19671 (N_19671,N_10674,N_13734);
or U19672 (N_19672,N_12634,N_10997);
or U19673 (N_19673,N_13191,N_13278);
nand U19674 (N_19674,N_10185,N_10616);
and U19675 (N_19675,N_10724,N_11595);
or U19676 (N_19676,N_14935,N_13473);
xnor U19677 (N_19677,N_11736,N_10598);
or U19678 (N_19678,N_10733,N_13373);
nand U19679 (N_19679,N_11864,N_11907);
or U19680 (N_19680,N_10035,N_10550);
and U19681 (N_19681,N_10504,N_10831);
nor U19682 (N_19682,N_10622,N_11895);
and U19683 (N_19683,N_10025,N_13301);
and U19684 (N_19684,N_14090,N_12174);
nor U19685 (N_19685,N_11233,N_10261);
nor U19686 (N_19686,N_10012,N_10027);
and U19687 (N_19687,N_11900,N_14905);
and U19688 (N_19688,N_12395,N_14010);
nand U19689 (N_19689,N_13463,N_12640);
nor U19690 (N_19690,N_14681,N_10241);
nor U19691 (N_19691,N_10007,N_14204);
nor U19692 (N_19692,N_14541,N_11023);
nand U19693 (N_19693,N_10643,N_12847);
nor U19694 (N_19694,N_12957,N_13459);
xnor U19695 (N_19695,N_14888,N_11663);
nor U19696 (N_19696,N_12544,N_10883);
and U19697 (N_19697,N_12785,N_14224);
nand U19698 (N_19698,N_11986,N_12899);
nor U19699 (N_19699,N_10097,N_10304);
nand U19700 (N_19700,N_12836,N_11023);
or U19701 (N_19701,N_11189,N_10461);
and U19702 (N_19702,N_11772,N_10001);
and U19703 (N_19703,N_12583,N_13710);
nand U19704 (N_19704,N_14209,N_10704);
and U19705 (N_19705,N_10200,N_10313);
nand U19706 (N_19706,N_11533,N_11218);
and U19707 (N_19707,N_10503,N_11974);
nor U19708 (N_19708,N_11138,N_11196);
or U19709 (N_19709,N_14362,N_10209);
nand U19710 (N_19710,N_14099,N_10554);
or U19711 (N_19711,N_14763,N_11265);
nand U19712 (N_19712,N_11046,N_12729);
nand U19713 (N_19713,N_12778,N_14142);
or U19714 (N_19714,N_14339,N_13957);
nor U19715 (N_19715,N_11225,N_11449);
and U19716 (N_19716,N_11795,N_14581);
nor U19717 (N_19717,N_10518,N_13989);
nand U19718 (N_19718,N_10438,N_12475);
nand U19719 (N_19719,N_10293,N_10387);
and U19720 (N_19720,N_14655,N_14873);
or U19721 (N_19721,N_13085,N_13630);
and U19722 (N_19722,N_12015,N_14964);
nand U19723 (N_19723,N_13679,N_13294);
nor U19724 (N_19724,N_11443,N_11358);
and U19725 (N_19725,N_13463,N_13564);
or U19726 (N_19726,N_11850,N_11279);
or U19727 (N_19727,N_11106,N_11441);
and U19728 (N_19728,N_14754,N_13170);
or U19729 (N_19729,N_11307,N_11401);
xnor U19730 (N_19730,N_12001,N_14668);
or U19731 (N_19731,N_13874,N_12662);
or U19732 (N_19732,N_12175,N_13262);
nand U19733 (N_19733,N_11722,N_13014);
nor U19734 (N_19734,N_14806,N_13209);
or U19735 (N_19735,N_12401,N_12313);
and U19736 (N_19736,N_10996,N_13138);
and U19737 (N_19737,N_13437,N_10346);
and U19738 (N_19738,N_10367,N_10750);
nand U19739 (N_19739,N_11215,N_10050);
or U19740 (N_19740,N_10741,N_14877);
nand U19741 (N_19741,N_12763,N_13930);
and U19742 (N_19742,N_13512,N_14184);
and U19743 (N_19743,N_10775,N_11417);
nand U19744 (N_19744,N_12419,N_14893);
or U19745 (N_19745,N_10180,N_14011);
and U19746 (N_19746,N_14426,N_12732);
nor U19747 (N_19747,N_12509,N_12598);
or U19748 (N_19748,N_14087,N_13179);
and U19749 (N_19749,N_12873,N_10768);
or U19750 (N_19750,N_11695,N_12842);
nand U19751 (N_19751,N_12222,N_11112);
xor U19752 (N_19752,N_14697,N_11276);
and U19753 (N_19753,N_11256,N_13447);
nand U19754 (N_19754,N_13655,N_14705);
nor U19755 (N_19755,N_14743,N_13075);
or U19756 (N_19756,N_13760,N_10063);
or U19757 (N_19757,N_10133,N_13553);
nor U19758 (N_19758,N_11894,N_13434);
or U19759 (N_19759,N_12144,N_10101);
and U19760 (N_19760,N_13540,N_11856);
nand U19761 (N_19761,N_11242,N_14031);
or U19762 (N_19762,N_13415,N_12272);
and U19763 (N_19763,N_10943,N_10416);
nand U19764 (N_19764,N_12633,N_11321);
nor U19765 (N_19765,N_12607,N_12088);
or U19766 (N_19766,N_12564,N_11205);
and U19767 (N_19767,N_13238,N_13293);
nand U19768 (N_19768,N_14735,N_10052);
nor U19769 (N_19769,N_10992,N_12567);
nor U19770 (N_19770,N_12139,N_12742);
nand U19771 (N_19771,N_12740,N_12257);
nand U19772 (N_19772,N_11648,N_13391);
or U19773 (N_19773,N_10564,N_11275);
nor U19774 (N_19774,N_10887,N_13726);
or U19775 (N_19775,N_12241,N_10704);
or U19776 (N_19776,N_10919,N_10081);
nor U19777 (N_19777,N_11333,N_12683);
and U19778 (N_19778,N_14865,N_10447);
and U19779 (N_19779,N_14081,N_10286);
nand U19780 (N_19780,N_10184,N_12757);
nand U19781 (N_19781,N_13017,N_13138);
or U19782 (N_19782,N_12021,N_13757);
or U19783 (N_19783,N_12672,N_13890);
nand U19784 (N_19784,N_14826,N_13645);
and U19785 (N_19785,N_12606,N_13741);
nand U19786 (N_19786,N_11587,N_12197);
nand U19787 (N_19787,N_13517,N_13075);
nand U19788 (N_19788,N_12647,N_11326);
nor U19789 (N_19789,N_14408,N_11132);
nor U19790 (N_19790,N_10925,N_11750);
nor U19791 (N_19791,N_13357,N_10587);
nor U19792 (N_19792,N_13494,N_13576);
nand U19793 (N_19793,N_13968,N_10781);
and U19794 (N_19794,N_12235,N_13261);
nor U19795 (N_19795,N_11016,N_14037);
nor U19796 (N_19796,N_10963,N_13170);
or U19797 (N_19797,N_11356,N_12796);
and U19798 (N_19798,N_12750,N_10922);
and U19799 (N_19799,N_13658,N_12523);
or U19800 (N_19800,N_12216,N_11327);
and U19801 (N_19801,N_10484,N_12253);
and U19802 (N_19802,N_13394,N_12863);
or U19803 (N_19803,N_10023,N_12442);
nand U19804 (N_19804,N_14341,N_13380);
nand U19805 (N_19805,N_14068,N_13858);
or U19806 (N_19806,N_13236,N_12561);
nor U19807 (N_19807,N_13085,N_13721);
nand U19808 (N_19808,N_11208,N_10682);
and U19809 (N_19809,N_12113,N_11967);
and U19810 (N_19810,N_14752,N_14854);
or U19811 (N_19811,N_11406,N_14638);
nand U19812 (N_19812,N_11606,N_12665);
nor U19813 (N_19813,N_10509,N_12029);
and U19814 (N_19814,N_13376,N_13509);
nand U19815 (N_19815,N_14903,N_12771);
nand U19816 (N_19816,N_12721,N_11075);
nand U19817 (N_19817,N_12217,N_12955);
nand U19818 (N_19818,N_10883,N_13065);
nor U19819 (N_19819,N_11407,N_13778);
nor U19820 (N_19820,N_14434,N_14793);
nand U19821 (N_19821,N_10860,N_14890);
nand U19822 (N_19822,N_11617,N_12589);
nand U19823 (N_19823,N_14801,N_13453);
or U19824 (N_19824,N_14834,N_14294);
nand U19825 (N_19825,N_10340,N_10707);
and U19826 (N_19826,N_12031,N_12467);
or U19827 (N_19827,N_10874,N_14136);
and U19828 (N_19828,N_11087,N_14405);
or U19829 (N_19829,N_13709,N_10317);
nor U19830 (N_19830,N_14356,N_10595);
nor U19831 (N_19831,N_14490,N_11528);
and U19832 (N_19832,N_12239,N_10749);
nor U19833 (N_19833,N_14946,N_13248);
and U19834 (N_19834,N_12041,N_13982);
or U19835 (N_19835,N_10570,N_13408);
and U19836 (N_19836,N_13423,N_13818);
nand U19837 (N_19837,N_10034,N_14308);
or U19838 (N_19838,N_11399,N_11345);
xnor U19839 (N_19839,N_13875,N_14546);
nand U19840 (N_19840,N_12096,N_10100);
nor U19841 (N_19841,N_12117,N_13292);
nand U19842 (N_19842,N_13164,N_14151);
or U19843 (N_19843,N_11512,N_10086);
nand U19844 (N_19844,N_11853,N_14127);
and U19845 (N_19845,N_10721,N_11062);
and U19846 (N_19846,N_13879,N_14115);
and U19847 (N_19847,N_10827,N_11163);
nor U19848 (N_19848,N_13387,N_10632);
nor U19849 (N_19849,N_11426,N_12572);
and U19850 (N_19850,N_13428,N_14944);
or U19851 (N_19851,N_12857,N_10423);
or U19852 (N_19852,N_11816,N_11170);
nor U19853 (N_19853,N_11788,N_14943);
or U19854 (N_19854,N_10282,N_14016);
nand U19855 (N_19855,N_11069,N_11551);
nor U19856 (N_19856,N_14701,N_11324);
or U19857 (N_19857,N_10391,N_12097);
and U19858 (N_19858,N_13314,N_10485);
nor U19859 (N_19859,N_14651,N_12966);
nand U19860 (N_19860,N_14362,N_11357);
nor U19861 (N_19861,N_11758,N_13083);
nor U19862 (N_19862,N_14420,N_11041);
nand U19863 (N_19863,N_12156,N_10004);
nor U19864 (N_19864,N_13811,N_10011);
and U19865 (N_19865,N_14983,N_10942);
xnor U19866 (N_19866,N_14868,N_12075);
nor U19867 (N_19867,N_13660,N_11741);
or U19868 (N_19868,N_11992,N_13833);
nand U19869 (N_19869,N_12275,N_12811);
or U19870 (N_19870,N_13135,N_12411);
nor U19871 (N_19871,N_10299,N_13941);
or U19872 (N_19872,N_11060,N_12616);
nand U19873 (N_19873,N_14461,N_12782);
or U19874 (N_19874,N_10345,N_10876);
nor U19875 (N_19875,N_13756,N_12090);
or U19876 (N_19876,N_13725,N_13764);
nand U19877 (N_19877,N_12752,N_13085);
and U19878 (N_19878,N_11982,N_13558);
and U19879 (N_19879,N_11548,N_12538);
and U19880 (N_19880,N_10524,N_14798);
or U19881 (N_19881,N_12208,N_13342);
and U19882 (N_19882,N_12206,N_10374);
and U19883 (N_19883,N_14432,N_11833);
nor U19884 (N_19884,N_11488,N_13860);
nand U19885 (N_19885,N_10059,N_12229);
or U19886 (N_19886,N_12588,N_13354);
and U19887 (N_19887,N_13891,N_14100);
and U19888 (N_19888,N_11547,N_12465);
nor U19889 (N_19889,N_10326,N_14916);
nand U19890 (N_19890,N_14218,N_12853);
nand U19891 (N_19891,N_11761,N_12236);
nand U19892 (N_19892,N_11850,N_12090);
xnor U19893 (N_19893,N_14420,N_14648);
or U19894 (N_19894,N_14838,N_12754);
nand U19895 (N_19895,N_11701,N_10283);
nand U19896 (N_19896,N_13946,N_14473);
or U19897 (N_19897,N_12569,N_13841);
nor U19898 (N_19898,N_10591,N_11818);
or U19899 (N_19899,N_13810,N_12296);
nor U19900 (N_19900,N_13938,N_10126);
nor U19901 (N_19901,N_11425,N_11838);
nand U19902 (N_19902,N_11660,N_13182);
nor U19903 (N_19903,N_14414,N_13989);
and U19904 (N_19904,N_11742,N_10576);
nand U19905 (N_19905,N_13053,N_10495);
or U19906 (N_19906,N_10988,N_14971);
or U19907 (N_19907,N_12582,N_13876);
nor U19908 (N_19908,N_13200,N_12739);
nand U19909 (N_19909,N_14034,N_11410);
nor U19910 (N_19910,N_10935,N_14054);
or U19911 (N_19911,N_13350,N_14381);
nor U19912 (N_19912,N_13733,N_14214);
or U19913 (N_19913,N_14258,N_11242);
nor U19914 (N_19914,N_11896,N_11485);
nor U19915 (N_19915,N_13307,N_11413);
nor U19916 (N_19916,N_10255,N_11662);
nand U19917 (N_19917,N_11813,N_11784);
and U19918 (N_19918,N_14664,N_14070);
nor U19919 (N_19919,N_12680,N_13062);
nand U19920 (N_19920,N_10366,N_13534);
nand U19921 (N_19921,N_12955,N_10644);
nor U19922 (N_19922,N_10215,N_14994);
or U19923 (N_19923,N_14247,N_13522);
nor U19924 (N_19924,N_14115,N_10619);
nor U19925 (N_19925,N_14633,N_13161);
or U19926 (N_19926,N_14324,N_10524);
nand U19927 (N_19927,N_11907,N_13840);
nor U19928 (N_19928,N_10148,N_11187);
and U19929 (N_19929,N_13978,N_10494);
and U19930 (N_19930,N_14618,N_12761);
nor U19931 (N_19931,N_11996,N_11456);
nor U19932 (N_19932,N_10035,N_11678);
or U19933 (N_19933,N_14016,N_12266);
or U19934 (N_19934,N_10792,N_12376);
and U19935 (N_19935,N_10578,N_12220);
and U19936 (N_19936,N_10799,N_13873);
nand U19937 (N_19937,N_12086,N_13452);
nor U19938 (N_19938,N_12789,N_12108);
or U19939 (N_19939,N_12819,N_10585);
or U19940 (N_19940,N_14288,N_10313);
or U19941 (N_19941,N_11329,N_14356);
nand U19942 (N_19942,N_11927,N_13803);
nor U19943 (N_19943,N_13019,N_12695);
nor U19944 (N_19944,N_12188,N_11337);
or U19945 (N_19945,N_14691,N_11093);
nor U19946 (N_19946,N_10653,N_13528);
nand U19947 (N_19947,N_10185,N_13820);
or U19948 (N_19948,N_13698,N_14950);
and U19949 (N_19949,N_14260,N_14881);
nand U19950 (N_19950,N_14348,N_12159);
nor U19951 (N_19951,N_14771,N_12985);
nor U19952 (N_19952,N_11431,N_10498);
and U19953 (N_19953,N_12576,N_10575);
and U19954 (N_19954,N_12198,N_12741);
or U19955 (N_19955,N_12906,N_13806);
nand U19956 (N_19956,N_14291,N_14836);
nand U19957 (N_19957,N_14730,N_10581);
nor U19958 (N_19958,N_13880,N_10548);
nand U19959 (N_19959,N_12167,N_13965);
nor U19960 (N_19960,N_11916,N_12142);
and U19961 (N_19961,N_13243,N_14826);
nand U19962 (N_19962,N_13719,N_14586);
and U19963 (N_19963,N_10584,N_13478);
and U19964 (N_19964,N_11585,N_11605);
nor U19965 (N_19965,N_11073,N_12316);
nand U19966 (N_19966,N_10446,N_11176);
or U19967 (N_19967,N_12259,N_12114);
nor U19968 (N_19968,N_13083,N_12028);
or U19969 (N_19969,N_10517,N_13831);
or U19970 (N_19970,N_14632,N_13409);
nand U19971 (N_19971,N_12998,N_12991);
or U19972 (N_19972,N_10649,N_11299);
nor U19973 (N_19973,N_14553,N_13749);
nand U19974 (N_19974,N_14317,N_14224);
and U19975 (N_19975,N_11646,N_10234);
or U19976 (N_19976,N_10067,N_14166);
or U19977 (N_19977,N_13222,N_10172);
or U19978 (N_19978,N_14415,N_12254);
and U19979 (N_19979,N_13904,N_10394);
nor U19980 (N_19980,N_12385,N_11002);
nand U19981 (N_19981,N_12489,N_10716);
nor U19982 (N_19982,N_12377,N_10981);
or U19983 (N_19983,N_12183,N_11954);
nand U19984 (N_19984,N_12295,N_11840);
nand U19985 (N_19985,N_13773,N_11042);
or U19986 (N_19986,N_13880,N_10958);
or U19987 (N_19987,N_13629,N_11368);
and U19988 (N_19988,N_14438,N_14578);
nor U19989 (N_19989,N_12397,N_14800);
nor U19990 (N_19990,N_11534,N_13734);
or U19991 (N_19991,N_11956,N_12333);
or U19992 (N_19992,N_14657,N_11139);
and U19993 (N_19993,N_12233,N_11315);
nand U19994 (N_19994,N_10557,N_14549);
or U19995 (N_19995,N_12388,N_14584);
nand U19996 (N_19996,N_10926,N_10202);
xnor U19997 (N_19997,N_13848,N_10884);
and U19998 (N_19998,N_13667,N_11135);
nand U19999 (N_19999,N_13193,N_10490);
nor UO_0 (O_0,N_18577,N_15944);
nor UO_1 (O_1,N_18004,N_18758);
or UO_2 (O_2,N_18088,N_17802);
nand UO_3 (O_3,N_19986,N_18309);
nor UO_4 (O_4,N_16543,N_18036);
or UO_5 (O_5,N_15644,N_15545);
nor UO_6 (O_6,N_19019,N_18259);
or UO_7 (O_7,N_16532,N_15012);
nand UO_8 (O_8,N_15098,N_15950);
nand UO_9 (O_9,N_15170,N_16736);
nand UO_10 (O_10,N_15404,N_18189);
nor UO_11 (O_11,N_17613,N_15078);
or UO_12 (O_12,N_19065,N_19604);
and UO_13 (O_13,N_17856,N_17783);
or UO_14 (O_14,N_19896,N_15532);
and UO_15 (O_15,N_15051,N_19420);
and UO_16 (O_16,N_17209,N_18879);
nor UO_17 (O_17,N_19423,N_17732);
nand UO_18 (O_18,N_18103,N_19723);
and UO_19 (O_19,N_19006,N_17649);
nand UO_20 (O_20,N_19419,N_19522);
nor UO_21 (O_21,N_16089,N_17887);
and UO_22 (O_22,N_15216,N_17340);
and UO_23 (O_23,N_19035,N_17761);
or UO_24 (O_24,N_18342,N_18028);
nor UO_25 (O_25,N_17187,N_15708);
or UO_26 (O_26,N_16769,N_18391);
and UO_27 (O_27,N_18407,N_17450);
and UO_28 (O_28,N_18565,N_18414);
nand UO_29 (O_29,N_19753,N_16560);
and UO_30 (O_30,N_17113,N_16962);
nor UO_31 (O_31,N_15229,N_15022);
nand UO_32 (O_32,N_17075,N_17134);
or UO_33 (O_33,N_17698,N_15328);
and UO_34 (O_34,N_18473,N_15983);
and UO_35 (O_35,N_17301,N_15332);
nor UO_36 (O_36,N_17695,N_16339);
or UO_37 (O_37,N_15611,N_17911);
and UO_38 (O_38,N_17499,N_16287);
and UO_39 (O_39,N_16763,N_19718);
nor UO_40 (O_40,N_18294,N_19754);
nor UO_41 (O_41,N_18078,N_19495);
and UO_42 (O_42,N_18285,N_18753);
nand UO_43 (O_43,N_19483,N_17399);
or UO_44 (O_44,N_16268,N_18889);
or UO_45 (O_45,N_18510,N_16284);
nand UO_46 (O_46,N_17051,N_15812);
nand UO_47 (O_47,N_15824,N_16124);
or UO_48 (O_48,N_18919,N_17728);
nand UO_49 (O_49,N_18578,N_19952);
and UO_50 (O_50,N_15972,N_19379);
nand UO_51 (O_51,N_15114,N_16487);
nand UO_52 (O_52,N_15093,N_15493);
nor UO_53 (O_53,N_18549,N_18821);
or UO_54 (O_54,N_19913,N_19563);
or UO_55 (O_55,N_16976,N_16886);
or UO_56 (O_56,N_17666,N_19623);
or UO_57 (O_57,N_17950,N_18156);
nand UO_58 (O_58,N_15206,N_16889);
or UO_59 (O_59,N_16171,N_17417);
and UO_60 (O_60,N_16282,N_17391);
nor UO_61 (O_61,N_15584,N_17617);
nor UO_62 (O_62,N_16159,N_19333);
and UO_63 (O_63,N_16020,N_19611);
nand UO_64 (O_64,N_19036,N_19650);
or UO_65 (O_65,N_18283,N_16387);
and UO_66 (O_66,N_17740,N_16685);
and UO_67 (O_67,N_19371,N_19814);
nand UO_68 (O_68,N_19429,N_19910);
and UO_69 (O_69,N_16117,N_16190);
and UO_70 (O_70,N_17658,N_18470);
and UO_71 (O_71,N_16181,N_18823);
nand UO_72 (O_72,N_16194,N_17982);
and UO_73 (O_73,N_17276,N_19820);
nor UO_74 (O_74,N_16998,N_19552);
nor UO_75 (O_75,N_19266,N_19220);
and UO_76 (O_76,N_17112,N_19962);
nand UO_77 (O_77,N_15041,N_15962);
nor UO_78 (O_78,N_17337,N_18187);
nand UO_79 (O_79,N_19147,N_18454);
nand UO_80 (O_80,N_16196,N_17049);
or UO_81 (O_81,N_15279,N_18999);
nand UO_82 (O_82,N_18747,N_18094);
and UO_83 (O_83,N_18692,N_19564);
nand UO_84 (O_84,N_18574,N_19346);
or UO_85 (O_85,N_18878,N_15221);
and UO_86 (O_86,N_19424,N_16508);
nand UO_87 (O_87,N_18296,N_15113);
nand UO_88 (O_88,N_17852,N_19710);
or UO_89 (O_89,N_17779,N_15571);
or UO_90 (O_90,N_15029,N_17387);
or UO_91 (O_91,N_15747,N_18116);
and UO_92 (O_92,N_18093,N_15265);
nand UO_93 (O_93,N_15560,N_18442);
nor UO_94 (O_94,N_18964,N_16659);
nand UO_95 (O_95,N_15361,N_16728);
nand UO_96 (O_96,N_17412,N_18907);
and UO_97 (O_97,N_19457,N_16254);
nor UO_98 (O_98,N_15499,N_18828);
or UO_99 (O_99,N_15855,N_18430);
nor UO_100 (O_100,N_18066,N_17124);
and UO_101 (O_101,N_18491,N_16338);
or UO_102 (O_102,N_18948,N_19943);
and UO_103 (O_103,N_19201,N_17586);
or UO_104 (O_104,N_18979,N_16442);
nor UO_105 (O_105,N_18820,N_18906);
nand UO_106 (O_106,N_16208,N_17904);
nor UO_107 (O_107,N_17273,N_16071);
nor UO_108 (O_108,N_19629,N_17826);
nand UO_109 (O_109,N_16365,N_19100);
and UO_110 (O_110,N_15432,N_15788);
and UO_111 (O_111,N_18554,N_19123);
or UO_112 (O_112,N_18630,N_18838);
and UO_113 (O_113,N_17096,N_19174);
and UO_114 (O_114,N_18928,N_17549);
or UO_115 (O_115,N_15874,N_15862);
nor UO_116 (O_116,N_17961,N_19772);
and UO_117 (O_117,N_19211,N_15414);
nor UO_118 (O_118,N_19187,N_17180);
and UO_119 (O_119,N_17667,N_18800);
and UO_120 (O_120,N_18083,N_15700);
or UO_121 (O_121,N_19183,N_19776);
and UO_122 (O_122,N_19177,N_17889);
and UO_123 (O_123,N_15075,N_18397);
or UO_124 (O_124,N_15223,N_19080);
and UO_125 (O_125,N_16872,N_16090);
and UO_126 (O_126,N_19242,N_15460);
and UO_127 (O_127,N_19778,N_18737);
or UO_128 (O_128,N_18529,N_18263);
and UO_129 (O_129,N_18084,N_16575);
or UO_130 (O_130,N_18045,N_19515);
or UO_131 (O_131,N_18846,N_19658);
nor UO_132 (O_132,N_18598,N_19181);
nand UO_133 (O_133,N_16537,N_16372);
nor UO_134 (O_134,N_19317,N_18129);
nor UO_135 (O_135,N_16906,N_16966);
nor UO_136 (O_136,N_17197,N_15924);
nand UO_137 (O_137,N_16642,N_19341);
nor UO_138 (O_138,N_19111,N_18572);
and UO_139 (O_139,N_18749,N_15082);
nand UO_140 (O_140,N_16264,N_19672);
nand UO_141 (O_141,N_15524,N_18362);
nor UO_142 (O_142,N_16926,N_17108);
or UO_143 (O_143,N_18789,N_17932);
nor UO_144 (O_144,N_17820,N_19037);
nor UO_145 (O_145,N_16014,N_15539);
or UO_146 (O_146,N_18575,N_17179);
nor UO_147 (O_147,N_16959,N_18541);
and UO_148 (O_148,N_16648,N_18787);
or UO_149 (O_149,N_19781,N_18883);
and UO_150 (O_150,N_15503,N_17804);
and UO_151 (O_151,N_15110,N_18620);
nand UO_152 (O_152,N_15322,N_17263);
nand UO_153 (O_153,N_16592,N_17748);
and UO_154 (O_154,N_15932,N_15392);
and UO_155 (O_155,N_18134,N_15405);
nor UO_156 (O_156,N_15912,N_16542);
nand UO_157 (O_157,N_18849,N_15429);
nand UO_158 (O_158,N_15522,N_17336);
nand UO_159 (O_159,N_18278,N_15242);
or UO_160 (O_160,N_16199,N_17511);
or UO_161 (O_161,N_18122,N_19408);
or UO_162 (O_162,N_16871,N_17342);
and UO_163 (O_163,N_19439,N_17780);
nor UO_164 (O_164,N_17490,N_15165);
or UO_165 (O_165,N_15709,N_19709);
or UO_166 (O_166,N_19933,N_15016);
nand UO_167 (O_167,N_19360,N_18546);
and UO_168 (O_168,N_18322,N_16121);
and UO_169 (O_169,N_16384,N_15890);
nand UO_170 (O_170,N_17442,N_16974);
nor UO_171 (O_171,N_17668,N_16803);
nand UO_172 (O_172,N_15379,N_15713);
nand UO_173 (O_173,N_15336,N_15500);
and UO_174 (O_174,N_19873,N_19173);
and UO_175 (O_175,N_18911,N_18232);
or UO_176 (O_176,N_17097,N_18276);
nand UO_177 (O_177,N_17758,N_16333);
nor UO_178 (O_178,N_15739,N_17947);
and UO_179 (O_179,N_18933,N_19344);
nand UO_180 (O_180,N_15084,N_16513);
and UO_181 (O_181,N_16309,N_16658);
nand UO_182 (O_182,N_19142,N_19272);
or UO_183 (O_183,N_19740,N_17217);
or UO_184 (O_184,N_16001,N_16169);
nand UO_185 (O_185,N_16224,N_16305);
nor UO_186 (O_186,N_17120,N_16297);
nand UO_187 (O_187,N_17058,N_19205);
or UO_188 (O_188,N_18857,N_19406);
or UO_189 (O_189,N_17080,N_16928);
or UO_190 (O_190,N_18042,N_17327);
and UO_191 (O_191,N_17561,N_16478);
nand UO_192 (O_192,N_18059,N_19306);
and UO_193 (O_193,N_18010,N_19127);
nor UO_194 (O_194,N_16447,N_15344);
and UO_195 (O_195,N_15507,N_17492);
and UO_196 (O_196,N_16055,N_17772);
nor UO_197 (O_197,N_17365,N_19176);
and UO_198 (O_198,N_16337,N_18405);
nor UO_199 (O_199,N_19885,N_15620);
nand UO_200 (O_200,N_18568,N_16600);
xor UO_201 (O_201,N_16450,N_18102);
nor UO_202 (O_202,N_16942,N_17648);
nor UO_203 (O_203,N_18241,N_16646);
nor UO_204 (O_204,N_18333,N_15062);
nor UO_205 (O_205,N_17101,N_19322);
xnor UO_206 (O_206,N_17584,N_19471);
and UO_207 (O_207,N_19315,N_18623);
or UO_208 (O_208,N_16587,N_15005);
and UO_209 (O_209,N_17150,N_16416);
and UO_210 (O_210,N_18786,N_15849);
nand UO_211 (O_211,N_15761,N_18996);
or UO_212 (O_212,N_17782,N_15948);
nor UO_213 (O_213,N_18387,N_16901);
nor UO_214 (O_214,N_19761,N_16366);
nor UO_215 (O_215,N_18480,N_16556);
nand UO_216 (O_216,N_17017,N_15616);
nand UO_217 (O_217,N_18131,N_18663);
and UO_218 (O_218,N_17743,N_17121);
and UO_219 (O_219,N_16348,N_17725);
nor UO_220 (O_220,N_18633,N_17752);
nand UO_221 (O_221,N_18525,N_17324);
or UO_222 (O_222,N_18386,N_16484);
nor UO_223 (O_223,N_18647,N_17624);
or UO_224 (O_224,N_18538,N_17266);
nand UO_225 (O_225,N_16098,N_18897);
or UO_226 (O_226,N_15196,N_15888);
nand UO_227 (O_227,N_18658,N_18221);
nor UO_228 (O_228,N_16645,N_16637);
nand UO_229 (O_229,N_16903,N_15796);
nor UO_230 (O_230,N_18389,N_16713);
and UO_231 (O_231,N_15696,N_18269);
nor UO_232 (O_232,N_16409,N_17127);
nor UO_233 (O_233,N_19641,N_17690);
xor UO_234 (O_234,N_16475,N_17000);
or UO_235 (O_235,N_16156,N_16899);
nand UO_236 (O_236,N_15273,N_16306);
nor UO_237 (O_237,N_18429,N_16065);
nor UO_238 (O_238,N_18238,N_17956);
or UO_239 (O_239,N_16651,N_17929);
and UO_240 (O_240,N_19869,N_19179);
and UO_241 (O_241,N_19250,N_16390);
nor UO_242 (O_242,N_19367,N_15635);
and UO_243 (O_243,N_17600,N_18893);
or UO_244 (O_244,N_18351,N_18356);
nand UO_245 (O_245,N_17840,N_19531);
nor UO_246 (O_246,N_18245,N_17583);
nor UO_247 (O_247,N_18484,N_16617);
or UO_248 (O_248,N_17456,N_18959);
nor UO_249 (O_249,N_19535,N_15204);
nand UO_250 (O_250,N_18884,N_15154);
or UO_251 (O_251,N_18409,N_15529);
nand UO_252 (O_252,N_18475,N_15418);
nor UO_253 (O_253,N_15348,N_17445);
and UO_254 (O_254,N_18839,N_19235);
nand UO_255 (O_255,N_15986,N_18812);
nor UO_256 (O_256,N_18360,N_19874);
and UO_257 (O_257,N_15810,N_19064);
and UO_258 (O_258,N_16405,N_17713);
and UO_259 (O_259,N_18783,N_18446);
nand UO_260 (O_260,N_16813,N_16673);
nand UO_261 (O_261,N_17859,N_15249);
nand UO_262 (O_262,N_17107,N_17654);
nand UO_263 (O_263,N_15658,N_17102);
nor UO_264 (O_264,N_18697,N_16107);
nand UO_265 (O_265,N_16495,N_17827);
or UO_266 (O_266,N_19878,N_19972);
or UO_267 (O_267,N_17634,N_18069);
nor UO_268 (O_268,N_19503,N_19270);
and UO_269 (O_269,N_19796,N_16539);
nor UO_270 (O_270,N_15570,N_15054);
nor UO_271 (O_271,N_17003,N_16005);
nor UO_272 (O_272,N_19588,N_16512);
and UO_273 (O_273,N_15157,N_16332);
and UO_274 (O_274,N_18383,N_17449);
nor UO_275 (O_275,N_16606,N_17906);
nor UO_276 (O_276,N_18530,N_19391);
nor UO_277 (O_277,N_18335,N_15859);
nor UO_278 (O_278,N_16815,N_15281);
or UO_279 (O_279,N_17063,N_15046);
or UO_280 (O_280,N_18885,N_16310);
nor UO_281 (O_281,N_17152,N_17937);
nor UO_282 (O_282,N_15125,N_17454);
and UO_283 (O_283,N_16170,N_18166);
and UO_284 (O_284,N_19131,N_18348);
or UO_285 (O_285,N_18349,N_18234);
nand UO_286 (O_286,N_18868,N_18141);
xor UO_287 (O_287,N_18662,N_16747);
nand UO_288 (O_288,N_18656,N_15673);
nand UO_289 (O_289,N_15509,N_19296);
and UO_290 (O_290,N_15171,N_18972);
or UO_291 (O_291,N_19219,N_15003);
and UO_292 (O_292,N_19448,N_19128);
nand UO_293 (O_293,N_18251,N_15166);
and UO_294 (O_294,N_16672,N_16158);
nor UO_295 (O_295,N_18524,N_15870);
and UO_296 (O_296,N_18412,N_18910);
nand UO_297 (O_297,N_17371,N_17665);
or UO_298 (O_298,N_19414,N_16355);
nand UO_299 (O_299,N_17248,N_15438);
or UO_300 (O_300,N_18695,N_19530);
or UO_301 (O_301,N_15080,N_19729);
nand UO_302 (O_302,N_16230,N_17216);
nor UO_303 (O_303,N_19657,N_19829);
nor UO_304 (O_304,N_15423,N_19840);
or UO_305 (O_305,N_16795,N_19038);
nand UO_306 (O_306,N_16127,N_18855);
nor UO_307 (O_307,N_17588,N_18952);
nand UO_308 (O_308,N_15536,N_18895);
nand UO_309 (O_309,N_19576,N_16443);
and UO_310 (O_310,N_18768,N_15366);
or UO_311 (O_311,N_17105,N_17086);
or UO_312 (O_312,N_15095,N_17558);
and UO_313 (O_313,N_19892,N_16589);
nand UO_314 (O_314,N_18138,N_16981);
and UO_315 (O_315,N_17957,N_19899);
or UO_316 (O_316,N_18628,N_19160);
nor UO_317 (O_317,N_16425,N_19090);
or UO_318 (O_318,N_17858,N_16419);
nand UO_319 (O_319,N_16357,N_16370);
or UO_320 (O_320,N_16270,N_17033);
or UO_321 (O_321,N_19711,N_17547);
and UO_322 (O_322,N_19567,N_19022);
nand UO_323 (O_323,N_16200,N_18767);
nand UO_324 (O_324,N_15711,N_19186);
and UO_325 (O_325,N_16367,N_16327);
nand UO_326 (O_326,N_15934,N_16953);
nand UO_327 (O_327,N_19669,N_17531);
or UO_328 (O_328,N_19852,N_19903);
nor UO_329 (O_329,N_17182,N_18898);
or UO_330 (O_330,N_19033,N_19700);
nor UO_331 (O_331,N_15868,N_18012);
and UO_332 (O_332,N_17200,N_17045);
or UO_333 (O_333,N_17855,N_16923);
nand UO_334 (O_334,N_17343,N_16979);
nand UO_335 (O_335,N_18621,N_19553);
or UO_336 (O_336,N_17990,N_18239);
nor UO_337 (O_337,N_18642,N_15559);
and UO_338 (O_338,N_16920,N_19598);
and UO_339 (O_339,N_17059,N_15145);
nor UO_340 (O_340,N_18992,N_19927);
nor UO_341 (O_341,N_18261,N_17238);
nand UO_342 (O_342,N_17622,N_19880);
and UO_343 (O_343,N_17874,N_17031);
or UO_344 (O_344,N_15454,N_15317);
or UO_345 (O_345,N_16079,N_19476);
nand UO_346 (O_346,N_17981,N_15502);
or UO_347 (O_347,N_17186,N_19170);
nand UO_348 (O_348,N_18727,N_19214);
nand UO_349 (O_349,N_15383,N_16661);
or UO_350 (O_350,N_15059,N_17447);
nor UO_351 (O_351,N_18773,N_15879);
and UO_352 (O_352,N_19436,N_17978);
and UO_353 (O_353,N_18536,N_16892);
nor UO_354 (O_354,N_15137,N_15428);
nor UO_355 (O_355,N_15629,N_16640);
nor UO_356 (O_356,N_17015,N_15451);
or UO_357 (O_357,N_16571,N_16324);
or UO_358 (O_358,N_19861,N_19671);
nand UO_359 (O_359,N_18504,N_15515);
nand UO_360 (O_360,N_19664,N_15079);
nand UO_361 (O_361,N_17892,N_17679);
and UO_362 (O_362,N_18458,N_16040);
or UO_363 (O_363,N_16582,N_17395);
nand UO_364 (O_364,N_18483,N_17202);
nand UO_365 (O_365,N_15477,N_19758);
and UO_366 (O_366,N_15642,N_19256);
nor UO_367 (O_367,N_17287,N_15627);
or UO_368 (O_368,N_15806,N_19286);
nand UO_369 (O_369,N_17935,N_18128);
or UO_370 (O_370,N_16438,N_19921);
nor UO_371 (O_371,N_19615,N_16485);
or UO_372 (O_372,N_18160,N_19410);
nor UO_373 (O_373,N_19676,N_16061);
or UO_374 (O_374,N_16376,N_19180);
and UO_375 (O_375,N_15027,N_15226);
nand UO_376 (O_376,N_19898,N_19893);
nand UO_377 (O_377,N_15094,N_18751);
or UO_378 (O_378,N_17686,N_19118);
nand UO_379 (O_379,N_18746,N_16328);
nor UO_380 (O_380,N_19248,N_17192);
or UO_381 (O_381,N_18619,N_15025);
and UO_382 (O_382,N_18210,N_18946);
nand UO_383 (O_383,N_19807,N_19724);
and UO_384 (O_384,N_15774,N_15891);
or UO_385 (O_385,N_16466,N_16745);
nand UO_386 (O_386,N_15353,N_19164);
nor UO_387 (O_387,N_16233,N_15970);
nor UO_388 (O_388,N_15973,N_18961);
or UO_389 (O_389,N_15933,N_17267);
and UO_390 (O_390,N_15795,N_18939);
nor UO_391 (O_391,N_16657,N_19162);
and UO_392 (O_392,N_15942,N_18958);
or UO_393 (O_393,N_18831,N_17446);
nor UO_394 (O_394,N_16641,N_16549);
nand UO_395 (O_395,N_16832,N_16567);
nand UO_396 (O_396,N_15207,N_19975);
and UO_397 (O_397,N_18610,N_15304);
nor UO_398 (O_398,N_18091,N_19244);
xor UO_399 (O_399,N_15666,N_15367);
and UO_400 (O_400,N_15519,N_16380);
and UO_401 (O_401,N_16799,N_17065);
or UO_402 (O_402,N_19839,N_15960);
or UO_403 (O_403,N_17060,N_19113);
and UO_404 (O_404,N_16807,N_16797);
or UO_405 (O_405,N_17355,N_16498);
nor UO_406 (O_406,N_15060,N_17463);
or UO_407 (O_407,N_19786,N_17281);
or UO_408 (O_408,N_18905,N_17744);
nand UO_409 (O_409,N_18203,N_15832);
and UO_410 (O_410,N_16474,N_15087);
or UO_411 (O_411,N_16113,N_17602);
nand UO_412 (O_412,N_19846,N_18861);
or UO_413 (O_413,N_16688,N_18158);
nand UO_414 (O_414,N_18039,N_17711);
nand UO_415 (O_415,N_17401,N_19905);
and UO_416 (O_416,N_16619,N_19649);
or UO_417 (O_417,N_17350,N_19459);
and UO_418 (O_418,N_17146,N_16655);
nand UO_419 (O_419,N_15587,N_16302);
nand UO_420 (O_420,N_17345,N_19045);
or UO_421 (O_421,N_17056,N_19145);
or UO_422 (O_422,N_15877,N_17380);
nor UO_423 (O_423,N_15038,N_16440);
or UO_424 (O_424,N_16334,N_15531);
or UO_425 (O_425,N_18167,N_16031);
and UO_426 (O_426,N_19210,N_15319);
nand UO_427 (O_427,N_16149,N_15566);
nor UO_428 (O_428,N_16004,N_19493);
nand UO_429 (O_429,N_18709,N_15132);
and UO_430 (O_430,N_16585,N_16929);
or UO_431 (O_431,N_17148,N_17372);
nand UO_432 (O_432,N_16064,N_19215);
nor UO_433 (O_433,N_19432,N_15471);
or UO_434 (O_434,N_15638,N_16530);
and UO_435 (O_435,N_15254,N_17661);
or UO_436 (O_436,N_15364,N_16449);
or UO_437 (O_437,N_16205,N_18627);
nor UO_438 (O_438,N_17509,N_17841);
nand UO_439 (O_439,N_18151,N_16433);
nand UO_440 (O_440,N_18657,N_18526);
nand UO_441 (O_441,N_15525,N_16679);
or UO_442 (O_442,N_15469,N_16683);
or UO_443 (O_443,N_15142,N_19224);
and UO_444 (O_444,N_15401,N_17198);
nand UO_445 (O_445,N_15321,N_17409);
nor UO_446 (O_446,N_15825,N_15993);
nor UO_447 (O_447,N_18481,N_15966);
and UO_448 (O_448,N_18731,N_19120);
or UO_449 (O_449,N_15742,N_19620);
or UO_450 (O_450,N_16228,N_17540);
xor UO_451 (O_451,N_17696,N_16588);
nand UO_452 (O_452,N_19354,N_15841);
nand UO_453 (O_453,N_15189,N_18306);
or UO_454 (O_454,N_16767,N_18206);
nor UO_455 (O_455,N_18708,N_15569);
or UO_456 (O_456,N_17895,N_16185);
nor UO_457 (O_457,N_15362,N_16082);
and UO_458 (O_458,N_17270,N_15352);
nand UO_459 (O_459,N_18415,N_19098);
and UO_460 (O_460,N_19345,N_15535);
and UO_461 (O_461,N_15826,N_17898);
and UO_462 (O_462,N_17411,N_17153);
or UO_463 (O_463,N_15955,N_17335);
nor UO_464 (O_464,N_19619,N_18495);
nand UO_465 (O_465,N_19453,N_15453);
nand UO_466 (O_466,N_17007,N_19271);
nand UO_467 (O_467,N_17918,N_19373);
and UO_468 (O_468,N_15886,N_16457);
and UO_469 (O_469,N_17778,N_18410);
and UO_470 (O_470,N_15577,N_15836);
or UO_471 (O_471,N_17203,N_19381);
nand UO_472 (O_472,N_19343,N_15914);
or UO_473 (O_473,N_19216,N_19894);
nand UO_474 (O_474,N_19759,N_18226);
nand UO_475 (O_475,N_16276,N_16599);
and UO_476 (O_476,N_15015,N_17268);
or UO_477 (O_477,N_19188,N_17422);
and UO_478 (O_478,N_18909,N_19714);
nor UO_479 (O_479,N_19475,N_15691);
or UO_480 (O_480,N_17448,N_16103);
or UO_481 (O_481,N_18970,N_15882);
nand UO_482 (O_482,N_16362,N_15119);
nor UO_483 (O_483,N_19883,N_19512);
and UO_484 (O_484,N_17520,N_17754);
nand UO_485 (O_485,N_18579,N_19252);
nand UO_486 (O_486,N_18850,N_18328);
nand UO_487 (O_487,N_15552,N_16676);
nand UO_488 (O_488,N_19764,N_15275);
nand UO_489 (O_489,N_16748,N_17388);
and UO_490 (O_490,N_15308,N_15476);
and UO_491 (O_491,N_19716,N_17765);
nand UO_492 (O_492,N_17819,N_16033);
and UO_493 (O_493,N_17694,N_18608);
or UO_494 (O_494,N_19397,N_16142);
nand UO_495 (O_495,N_16080,N_15656);
or UO_496 (O_496,N_16373,N_18368);
or UO_497 (O_497,N_19196,N_16534);
nand UO_498 (O_498,N_18449,N_18808);
nor UO_499 (O_499,N_17604,N_15619);
or UO_500 (O_500,N_16781,N_15447);
nor UO_501 (O_501,N_16710,N_19284);
nand UO_502 (O_502,N_15719,N_15623);
or UO_503 (O_503,N_16184,N_15402);
nor UO_504 (O_504,N_15875,N_17538);
or UO_505 (O_505,N_17229,N_15801);
nand UO_506 (O_506,N_19940,N_15071);
or UO_507 (O_507,N_18683,N_16323);
xor UO_508 (O_508,N_16250,N_17710);
nor UO_509 (O_509,N_15478,N_15178);
and UO_510 (O_510,N_16482,N_17405);
or UO_511 (O_511,N_16441,N_18308);
xnor UO_512 (O_512,N_15574,N_18533);
nand UO_513 (O_513,N_15480,N_16467);
nand UO_514 (O_514,N_19957,N_19402);
nand UO_515 (O_515,N_15981,N_15406);
or UO_516 (O_516,N_15586,N_16347);
or UO_517 (O_517,N_19290,N_18456);
nand UO_518 (O_518,N_16193,N_19227);
nor UO_519 (O_519,N_17389,N_15491);
and UO_520 (O_520,N_16675,N_19585);
nor UO_521 (O_521,N_17702,N_16201);
or UO_522 (O_522,N_17004,N_16432);
nor UO_523 (O_523,N_15091,N_15576);
nand UO_524 (O_524,N_18341,N_19101);
or UO_525 (O_525,N_16206,N_17322);
nand UO_526 (O_526,N_18997,N_18372);
and UO_527 (O_527,N_16211,N_15228);
nand UO_528 (O_528,N_16609,N_15508);
or UO_529 (O_529,N_15318,N_19960);
and UO_530 (O_530,N_18327,N_17062);
or UO_531 (O_531,N_18025,N_16209);
and UO_532 (O_532,N_16147,N_15904);
or UO_533 (O_533,N_15064,N_19150);
and UO_534 (O_534,N_18521,N_16690);
nor UO_535 (O_535,N_16011,N_17067);
nand UO_536 (O_536,N_15013,N_19509);
and UO_537 (O_537,N_16921,N_19279);
or UO_538 (O_538,N_16361,N_18264);
nand UO_539 (O_539,N_19813,N_15816);
nor UO_540 (O_540,N_15732,N_18790);
or UO_541 (O_541,N_15595,N_16346);
nand UO_542 (O_542,N_17441,N_15813);
nand UO_543 (O_543,N_17505,N_19914);
nor UO_544 (O_544,N_18371,N_17341);
nand UO_545 (O_545,N_19437,N_17620);
and UO_546 (O_546,N_18392,N_18431);
and UO_547 (O_547,N_15293,N_18803);
nand UO_548 (O_548,N_18394,N_15847);
nand UO_549 (O_549,N_17542,N_17529);
or UO_550 (O_550,N_18586,N_18459);
and UO_551 (O_551,N_19646,N_15112);
or UO_552 (O_552,N_15705,N_19027);
or UO_553 (O_553,N_17770,N_19977);
nor UO_554 (O_554,N_16021,N_15072);
or UO_555 (O_555,N_17873,N_19207);
and UO_556 (O_556,N_16895,N_19991);
nand UO_557 (O_557,N_15880,N_18848);
nand UO_558 (O_558,N_19025,N_18321);
or UO_559 (O_559,N_16612,N_19338);
nor UO_560 (O_560,N_17800,N_18570);
and UO_561 (O_561,N_18988,N_16825);
and UO_562 (O_562,N_19541,N_15939);
nand UO_563 (O_563,N_16751,N_15906);
and UO_564 (O_564,N_16766,N_18581);
nand UO_565 (O_565,N_18289,N_19403);
and UO_566 (O_566,N_17199,N_16702);
nand UO_567 (O_567,N_15272,N_17236);
or UO_568 (O_568,N_19044,N_17771);
and UO_569 (O_569,N_16291,N_17607);
and UO_570 (O_570,N_17418,N_16489);
nand UO_571 (O_571,N_16322,N_19855);
nand UO_572 (O_572,N_18195,N_17709);
and UO_573 (O_573,N_17587,N_17862);
or UO_574 (O_574,N_15007,N_16106);
nor UO_575 (O_575,N_15534,N_19158);
nor UO_576 (O_576,N_18917,N_18140);
nor UO_577 (O_577,N_19501,N_16595);
or UO_578 (O_578,N_19607,N_16697);
or UO_579 (O_579,N_16120,N_17635);
or UO_580 (O_580,N_16488,N_15244);
or UO_581 (O_581,N_17924,N_17810);
or UO_582 (O_582,N_18990,N_17513);
or UO_583 (O_583,N_16550,N_18105);
or UO_584 (O_584,N_16491,N_15606);
xor UO_585 (O_585,N_16653,N_17041);
nand UO_586 (O_586,N_18743,N_18987);
nand UO_587 (O_587,N_15585,N_17550);
nand UO_588 (O_588,N_16918,N_16051);
nor UO_589 (O_589,N_18488,N_15150);
nor UO_590 (O_590,N_16706,N_16598);
and UO_591 (O_591,N_16738,N_15057);
nand UO_592 (O_592,N_18466,N_18024);
or UO_593 (O_593,N_15878,N_17557);
nand UO_594 (O_594,N_15643,N_15397);
nor UO_595 (O_595,N_19032,N_17662);
or UO_596 (O_596,N_15685,N_16884);
or UO_597 (O_597,N_18750,N_19715);
or UO_598 (O_598,N_17460,N_15030);
or UO_599 (O_599,N_15484,N_18563);
nand UO_600 (O_600,N_19871,N_17682);
nand UO_601 (O_601,N_16418,N_17023);
nor UO_602 (O_602,N_19217,N_15530);
or UO_603 (O_603,N_19931,N_17193);
nand UO_604 (O_604,N_19015,N_16701);
or UO_605 (O_605,N_18912,N_15702);
nand UO_606 (O_606,N_19490,N_18200);
or UO_607 (O_607,N_19386,N_15608);
nand UO_608 (O_608,N_18676,N_16189);
or UO_609 (O_609,N_18260,N_15769);
nand UO_610 (O_610,N_19732,N_16620);
or UO_611 (O_611,N_19735,N_15692);
nand UO_612 (O_612,N_18778,N_16897);
nand UO_613 (O_613,N_16796,N_16544);
nand UO_614 (O_614,N_17585,N_16671);
nor UO_615 (O_615,N_16364,N_17647);
or UO_616 (O_616,N_15548,N_18926);
nor UO_617 (O_617,N_16172,N_18614);
nor UO_618 (O_618,N_17878,N_15996);
and UO_619 (O_619,N_19788,N_16108);
and UO_620 (O_620,N_17219,N_15804);
nand UO_621 (O_621,N_16198,N_17443);
nor UO_622 (O_622,N_19946,N_17618);
and UO_623 (O_623,N_15725,N_16336);
nor UO_624 (O_624,N_16504,N_18871);
or UO_625 (O_625,N_18824,N_19949);
nor UO_626 (O_626,N_16952,N_16192);
nand UO_627 (O_627,N_16025,N_16614);
nand UO_628 (O_628,N_19602,N_19152);
nand UO_629 (O_629,N_18179,N_15665);
nor UO_630 (O_630,N_19730,N_17357);
nor UO_631 (O_631,N_18337,N_18908);
and UO_632 (O_632,N_15128,N_19085);
or UO_633 (O_633,N_17722,N_15090);
or UO_634 (O_634,N_16951,N_15122);
nor UO_635 (O_635,N_15938,N_16077);
nor UO_636 (O_636,N_16410,N_16036);
and UO_637 (O_637,N_16932,N_18227);
nand UO_638 (O_638,N_15325,N_16798);
nand UO_639 (O_639,N_16581,N_19845);
nor UO_640 (O_640,N_19292,N_16817);
nor UO_641 (O_641,N_19347,N_16398);
nand UO_642 (O_642,N_16015,N_19575);
nor UO_643 (O_643,N_16887,N_17118);
nand UO_644 (O_644,N_15802,N_15674);
and UO_645 (O_645,N_18983,N_15437);
and UO_646 (O_646,N_16772,N_19692);
or UO_647 (O_647,N_18482,N_19133);
nor UO_648 (O_648,N_17328,N_19046);
nand UO_649 (O_649,N_18589,N_17569);
and UO_650 (O_650,N_15235,N_16426);
nand UO_651 (O_651,N_16345,N_16656);
nor UO_652 (O_652,N_19388,N_19529);
nor UO_653 (O_653,N_17057,N_16866);
and UO_654 (O_654,N_16680,N_16350);
nor UO_655 (O_655,N_15833,N_19295);
nand UO_656 (O_656,N_16829,N_17201);
or UO_657 (O_657,N_18213,N_15389);
nand UO_658 (O_658,N_15413,N_18977);
or UO_659 (O_659,N_19278,N_19119);
and UO_660 (O_660,N_16665,N_16486);
and UO_661 (O_661,N_18262,N_17608);
nand UO_662 (O_662,N_15305,N_17481);
and UO_663 (O_663,N_17700,N_17566);
or UO_664 (O_664,N_15045,N_15134);
and UO_665 (O_665,N_17949,N_16050);
and UO_666 (O_666,N_15393,N_19148);
or UO_667 (O_667,N_19968,N_16842);
and UO_668 (O_668,N_16203,N_15593);
nor UO_669 (O_669,N_19003,N_15468);
or UO_670 (O_670,N_19502,N_19433);
or UO_671 (O_671,N_16636,N_15929);
nand UO_672 (O_672,N_18573,N_18096);
nand UO_673 (O_673,N_17246,N_19745);
nor UO_674 (O_674,N_17329,N_16148);
nor UO_675 (O_675,N_15276,N_17533);
and UO_676 (O_676,N_19798,N_17465);
nand UO_677 (O_677,N_15654,N_16983);
and UO_678 (O_678,N_16757,N_19321);
nand UO_679 (O_679,N_16937,N_16547);
or UO_680 (O_680,N_16756,N_17130);
nor UO_681 (O_681,N_15065,N_17736);
or UO_682 (O_682,N_17699,N_15430);
and UO_683 (O_683,N_17299,N_15417);
nor UO_684 (O_684,N_18188,N_15667);
and UO_685 (O_685,N_16873,N_15217);
nor UO_686 (O_686,N_16439,N_18085);
and UO_687 (O_687,N_19990,N_18223);
and UO_688 (O_688,N_18235,N_15035);
or UO_689 (O_689,N_18191,N_17678);
nand UO_690 (O_690,N_17907,N_15307);
nor UO_691 (O_691,N_17166,N_17601);
nand UO_692 (O_692,N_15215,N_19765);
nand UO_693 (O_693,N_18081,N_19261);
nand UO_694 (O_694,N_17261,N_19538);
nand UO_695 (O_695,N_17142,N_17999);
nor UO_696 (O_696,N_17504,N_19835);
nor UO_697 (O_697,N_18476,N_15779);
nor UO_698 (O_698,N_16940,N_18154);
nor UO_699 (O_699,N_18301,N_16404);
and UO_700 (O_700,N_18165,N_16326);
or UO_701 (O_701,N_19327,N_17379);
nand UO_702 (O_702,N_16851,N_16273);
nand UO_703 (O_703,N_15959,N_16427);
or UO_704 (O_704,N_16822,N_18361);
and UO_705 (O_705,N_15734,N_15850);
nor UO_706 (O_706,N_18492,N_16818);
xor UO_707 (O_707,N_16984,N_16758);
and UO_708 (O_708,N_19245,N_15817);
nand UO_709 (O_709,N_16994,N_17727);
and UO_710 (O_710,N_17178,N_17785);
nand UO_711 (O_711,N_19443,N_18418);
or UO_712 (O_712,N_17038,N_15033);
or UO_713 (O_713,N_18303,N_15175);
nor UO_714 (O_714,N_19956,N_18949);
nand UO_715 (O_715,N_17094,N_15211);
and UO_716 (O_716,N_16008,N_18845);
and UO_717 (O_717,N_17882,N_19609);
nor UO_718 (O_718,N_15693,N_16891);
nand UO_719 (O_719,N_15495,N_17131);
nor UO_720 (O_720,N_19633,N_16607);
and UO_721 (O_721,N_15865,N_16591);
nand UO_722 (O_722,N_19578,N_17279);
nor UO_723 (O_723,N_17141,N_15575);
and UO_724 (O_724,N_15230,N_19577);
nand UO_725 (O_725,N_16408,N_19225);
or UO_726 (O_726,N_19587,N_19137);
nor UO_727 (O_727,N_15537,N_17953);
nand UO_728 (O_728,N_18528,N_18090);
nand UO_729 (O_729,N_19837,N_18268);
nor UO_730 (O_730,N_17589,N_15391);
or UO_731 (O_731,N_15210,N_17310);
or UO_732 (O_732,N_15147,N_17792);
nand UO_733 (O_733,N_18969,N_19738);
and UO_734 (O_734,N_16808,N_19140);
or UO_735 (O_735,N_16517,N_17917);
nor UO_736 (O_736,N_19365,N_15956);
or UO_737 (O_737,N_16075,N_17663);
and UO_738 (O_738,N_19395,N_16002);
nor UO_739 (O_739,N_15913,N_17087);
and UO_740 (O_740,N_18719,N_15042);
nor UO_741 (O_741,N_15731,N_16593);
and UO_742 (O_742,N_16719,N_16067);
nor UO_743 (O_743,N_18689,N_15444);
and UO_744 (O_744,N_18745,N_16259);
nor UO_745 (O_745,N_16933,N_16225);
or UO_746 (O_746,N_18043,N_18265);
or UO_747 (O_747,N_15101,N_18257);
and UO_748 (O_748,N_15594,N_17407);
or UO_749 (O_749,N_15756,N_15829);
and UO_750 (O_750,N_17471,N_15023);
and UO_751 (O_751,N_15937,N_18671);
or UO_752 (O_752,N_17296,N_16633);
nand UO_753 (O_753,N_18702,N_15243);
nor UO_754 (O_754,N_16342,N_16826);
and UO_755 (O_755,N_15919,N_17410);
and UO_756 (O_756,N_19193,N_17029);
and UO_757 (O_757,N_19223,N_16022);
or UO_758 (O_758,N_19048,N_19309);
or UO_759 (O_759,N_15604,N_19519);
or UO_760 (O_760,N_17637,N_19487);
nor UO_761 (O_761,N_15680,N_16820);
nor UO_762 (O_762,N_16074,N_15940);
nor UO_763 (O_763,N_19654,N_19750);
or UO_764 (O_764,N_15155,N_17375);
or UO_765 (O_765,N_19887,N_17352);
or UO_766 (O_766,N_17891,N_18101);
nand UO_767 (O_767,N_18068,N_17879);
or UO_768 (O_768,N_15320,N_17222);
and UO_769 (O_769,N_19107,N_16191);
or UO_770 (O_770,N_19191,N_15289);
and UO_771 (O_771,N_19656,N_16922);
or UO_772 (O_772,N_16644,N_17543);
and UO_773 (O_773,N_17052,N_17019);
and UO_774 (O_774,N_18903,N_15306);
nand UO_775 (O_775,N_15528,N_18740);
nand UO_776 (O_776,N_18854,N_16980);
or UO_777 (O_777,N_19886,N_16666);
and UO_778 (O_778,N_16411,N_19438);
nand UO_779 (O_779,N_18772,N_18307);
and UO_780 (O_780,N_15152,N_15634);
nand UO_781 (O_781,N_19954,N_16616);
or UO_782 (O_782,N_19265,N_19590);
or UO_783 (O_783,N_16515,N_17811);
xor UO_784 (O_784,N_19178,N_17987);
and UO_785 (O_785,N_16565,N_17995);
or UO_786 (O_786,N_19428,N_15753);
nor UO_787 (O_787,N_17707,N_18074);
nor UO_788 (O_788,N_17484,N_19533);
or UO_789 (O_789,N_15180,N_15350);
nand UO_790 (O_790,N_16212,N_15590);
and UO_791 (O_791,N_16470,N_15077);
and UO_792 (O_792,N_18461,N_19685);
nand UO_793 (O_793,N_17283,N_17208);
and UO_794 (O_794,N_18117,N_18804);
and UO_795 (O_795,N_17383,N_15994);
nor UO_796 (O_796,N_19694,N_15612);
nand UO_797 (O_797,N_16845,N_17636);
nand UO_798 (O_798,N_16317,N_18971);
and UO_799 (O_799,N_15511,N_19659);
nor UO_800 (O_800,N_18557,N_18457);
or UO_801 (O_801,N_16741,N_16856);
nand UO_802 (O_802,N_19249,N_18777);
and UO_803 (O_803,N_19783,N_17482);
nor UO_804 (O_804,N_17733,N_18672);
nor UO_805 (O_805,N_18793,N_19630);
or UO_806 (O_806,N_16464,N_19690);
or UO_807 (O_807,N_19200,N_17085);
nand UO_808 (O_808,N_15185,N_16258);
nand UO_809 (O_809,N_19746,N_19362);
nor UO_810 (O_810,N_16237,N_16625);
nor UO_811 (O_811,N_17292,N_19866);
nand UO_812 (O_812,N_18780,N_17374);
nor UO_813 (O_813,N_17363,N_16091);
nand UO_814 (O_814,N_18425,N_19255);
nor UO_815 (O_815,N_16062,N_17794);
xor UO_816 (O_816,N_16776,N_18182);
or UO_817 (O_817,N_18030,N_17272);
and UO_818 (O_818,N_18532,N_18542);
or UO_819 (O_819,N_19847,N_16931);
nor UO_820 (O_820,N_18655,N_16782);
nor UO_821 (O_821,N_16558,N_17010);
or UO_822 (O_822,N_19213,N_17514);
or UO_823 (O_823,N_16275,N_15607);
nand UO_824 (O_824,N_17020,N_17701);
nand UO_825 (O_825,N_18782,N_15969);
nor UO_826 (O_826,N_16678,N_19078);
or UO_827 (O_827,N_16583,N_16660);
xor UO_828 (O_828,N_15416,N_15592);
and UO_829 (O_829,N_15127,N_19404);
or UO_830 (O_830,N_18252,N_18467);
nor UO_831 (O_831,N_18401,N_19665);
nor UO_832 (O_832,N_17582,N_17390);
nand UO_833 (O_833,N_17524,N_16481);
nand UO_834 (O_834,N_16574,N_17125);
nor UO_835 (O_835,N_15011,N_18560);
and UO_836 (O_836,N_18624,N_16604);
or UO_837 (O_837,N_18762,N_16436);
nor UO_838 (O_838,N_17224,N_16572);
nand UO_839 (O_839,N_17068,N_19028);
or UO_840 (O_840,N_17119,N_15840);
nand UO_841 (O_841,N_18847,N_17851);
nand UO_842 (O_842,N_17486,N_19728);
nand UO_843 (O_843,N_19780,N_15737);
and UO_844 (O_844,N_15807,N_18046);
or UO_845 (O_845,N_17872,N_19281);
or UO_846 (O_846,N_16078,N_18133);
nor UO_847 (O_847,N_15808,N_16311);
or UO_848 (O_848,N_19784,N_16533);
and UO_849 (O_849,N_15008,N_18286);
nand UO_850 (O_850,N_19841,N_19639);
or UO_851 (O_851,N_15446,N_17726);
and UO_852 (O_852,N_18650,N_15809);
or UO_853 (O_853,N_17815,N_15542);
or UO_854 (O_854,N_16840,N_17084);
nand UO_855 (O_855,N_19713,N_15772);
and UO_856 (O_856,N_17609,N_15897);
and UO_857 (O_857,N_17347,N_19924);
or UO_858 (O_858,N_15312,N_15497);
nand UO_859 (O_859,N_18588,N_18423);
nor UO_860 (O_860,N_17436,N_16610);
and UO_861 (O_861,N_16833,N_19026);
nor UO_862 (O_862,N_19074,N_15735);
nor UO_863 (O_863,N_19267,N_18686);
and UO_864 (O_864,N_15070,N_19226);
nand UO_865 (O_865,N_17865,N_15412);
nand UO_866 (O_866,N_17077,N_19087);
and UO_867 (O_867,N_16765,N_17559);
or UO_868 (O_868,N_19581,N_16308);
or UO_869 (O_869,N_15031,N_16522);
and UO_870 (O_870,N_19431,N_15259);
nand UO_871 (O_871,N_16375,N_19524);
or UO_872 (O_872,N_17210,N_19951);
nor UO_873 (O_873,N_15848,N_17572);
nand UO_874 (O_874,N_19877,N_16269);
nor UO_875 (O_875,N_19826,N_17474);
nand UO_876 (O_876,N_15789,N_18302);
and UO_877 (O_877,N_18497,N_17451);
xnor UO_878 (O_878,N_19703,N_19425);
and UO_879 (O_879,N_18056,N_15034);
nor UO_880 (O_880,N_16087,N_15017);
and UO_881 (O_881,N_17759,N_19491);
nor UO_882 (O_882,N_17156,N_15050);
or UO_883 (O_883,N_19310,N_15936);
nor UO_884 (O_884,N_18146,N_19416);
nand UO_885 (O_885,N_17556,N_19599);
nand UO_886 (O_886,N_19282,N_19539);
nor UO_887 (O_887,N_18474,N_15470);
and UO_888 (O_888,N_15896,N_15436);
or UO_889 (O_889,N_17438,N_15990);
nor UO_890 (O_890,N_18559,N_19029);
and UO_891 (O_891,N_18724,N_16729);
nor UO_892 (O_892,N_15728,N_15464);
nor UO_893 (O_893,N_15853,N_16179);
nor UO_894 (O_894,N_18955,N_17043);
and UO_895 (O_895,N_15978,N_17691);
and UO_896 (O_896,N_18517,N_17606);
or UO_897 (O_897,N_16292,N_15382);
or UO_898 (O_898,N_17307,N_16972);
nand UO_899 (O_899,N_17139,N_15723);
or UO_900 (O_900,N_18806,N_16267);
or UO_901 (O_901,N_18819,N_19548);
nor UO_902 (O_902,N_18514,N_16229);
or UO_903 (O_903,N_19095,N_19299);
and UO_904 (O_904,N_18272,N_17250);
and UO_905 (O_905,N_18796,N_17459);
nor UO_906 (O_906,N_15295,N_17610);
xor UO_907 (O_907,N_19906,N_17980);
nor UO_908 (O_908,N_19208,N_17983);
nor UO_909 (O_909,N_17669,N_19355);
nor UO_910 (O_910,N_18704,N_16234);
nand UO_911 (O_911,N_19904,N_18369);
or UO_912 (O_912,N_16875,N_16982);
or UO_913 (O_913,N_18050,N_19280);
nand UO_914 (O_914,N_17814,N_17218);
nor UO_915 (O_915,N_17674,N_15284);
nor UO_916 (O_916,N_16854,N_16711);
nor UO_917 (O_917,N_15267,N_15927);
nand UO_918 (O_918,N_17922,N_15283);
or UO_919 (O_919,N_17971,N_18797);
nor UO_920 (O_920,N_17378,N_16186);
nand UO_921 (O_921,N_15296,N_18716);
and UO_922 (O_922,N_19971,N_15191);
or UO_923 (O_923,N_15752,N_16253);
nand UO_924 (O_924,N_17364,N_15252);
and UO_925 (O_925,N_18852,N_15467);
nor UO_926 (O_926,N_18211,N_15058);
nand UO_927 (O_927,N_19151,N_18938);
nor UO_928 (O_928,N_17517,N_18665);
nand UO_929 (O_929,N_18587,N_19236);
nor UO_930 (O_930,N_16421,N_16037);
and UO_931 (O_931,N_18114,N_15411);
nand UO_932 (O_932,N_16392,N_15327);
nor UO_933 (O_933,N_16118,N_16682);
and UO_934 (O_934,N_16301,N_16114);
and UO_935 (O_935,N_15533,N_15561);
and UO_936 (O_936,N_18011,N_18520);
nand UO_937 (O_937,N_18537,N_18345);
and UO_938 (O_938,N_15231,N_18003);
or UO_939 (O_939,N_18755,N_16784);
and UO_940 (O_940,N_18366,N_18607);
nand UO_941 (O_941,N_18965,N_19129);
or UO_942 (O_942,N_17697,N_17416);
and UO_943 (O_943,N_15907,N_15456);
or UO_944 (O_944,N_18157,N_16216);
nor UO_945 (O_945,N_18612,N_18645);
and UO_946 (O_946,N_18827,N_18127);
or UO_947 (O_947,N_17920,N_19721);
nor UO_948 (O_948,N_16725,N_15985);
and UO_949 (O_949,N_19568,N_18694);
or UO_950 (O_950,N_19138,N_19190);
nor UO_951 (O_951,N_19768,N_16777);
and UO_952 (O_952,N_19169,N_17265);
nand UO_953 (O_953,N_18567,N_16786);
nand UO_954 (O_954,N_15203,N_15618);
and UO_955 (O_955,N_16139,N_17493);
nand UO_956 (O_956,N_16835,N_15842);
and UO_957 (O_957,N_19771,N_15766);
nand UO_958 (O_958,N_19736,N_17249);
or UO_959 (O_959,N_17116,N_18637);
or UO_960 (O_960,N_15963,N_16060);
nor UO_961 (O_961,N_19209,N_15682);
nand UO_962 (O_962,N_19542,N_15375);
nand UO_963 (O_963,N_16843,N_18636);
nand UO_964 (O_964,N_16667,N_17432);
nor UO_965 (O_965,N_16576,N_16936);
or UO_966 (O_966,N_19104,N_16987);
nor UO_967 (O_967,N_17991,N_16638);
or UO_968 (O_968,N_18125,N_18669);
nand UO_969 (O_969,N_18019,N_17469);
nor UO_970 (O_970,N_18222,N_17595);
or UO_971 (O_971,N_17188,N_16602);
nor UO_972 (O_972,N_18896,N_18698);
xor UO_973 (O_973,N_15099,N_17143);
nand UO_974 (O_974,N_18305,N_15750);
and UO_975 (O_975,N_17477,N_18998);
and UO_976 (O_976,N_19779,N_16502);
or UO_977 (O_977,N_17546,N_18053);
and UO_978 (O_978,N_17928,N_19110);
nand UO_979 (O_979,N_19258,N_19999);
or UO_980 (O_980,N_19451,N_16570);
and UO_981 (O_981,N_17313,N_16883);
and UO_982 (O_982,N_18060,N_15895);
and UO_983 (O_983,N_18679,N_17824);
or UO_984 (O_984,N_17829,N_15856);
and UO_985 (O_985,N_19613,N_17818);
nor UO_986 (O_986,N_19484,N_19259);
nand UO_987 (O_987,N_17821,N_17464);
nand UO_988 (O_988,N_15946,N_15311);
nand UO_989 (O_989,N_18681,N_16045);
or UO_990 (O_990,N_19558,N_17429);
nor UO_991 (O_991,N_17958,N_17262);
or UO_992 (O_992,N_19304,N_17403);
nor UO_993 (O_993,N_16954,N_19018);
and UO_994 (O_994,N_15439,N_17093);
and UO_995 (O_995,N_16461,N_17870);
nor UO_996 (O_996,N_17944,N_15765);
nor UO_997 (O_997,N_19600,N_19836);
nand UO_998 (O_998,N_18705,N_15102);
and UO_999 (O_999,N_19762,N_17822);
nor UO_1000 (O_1000,N_15814,N_19550);
xnor UO_1001 (O_1001,N_16885,N_17361);
or UO_1002 (O_1002,N_19544,N_19467);
nor UO_1003 (O_1003,N_16030,N_18355);
and UO_1004 (O_1004,N_19314,N_19859);
nand UO_1005 (O_1005,N_15019,N_15582);
nor UO_1006 (O_1006,N_18130,N_19017);
nand UO_1007 (O_1007,N_15967,N_15931);
nor UO_1008 (O_1008,N_15073,N_16775);
and UO_1009 (O_1009,N_19966,N_17402);
or UO_1010 (O_1010,N_19378,N_16076);
and UO_1011 (O_1011,N_15236,N_18534);
and UO_1012 (O_1012,N_15360,N_16423);
or UO_1013 (O_1013,N_16122,N_17321);
nor UO_1014 (O_1014,N_15381,N_19114);
and UO_1015 (O_1015,N_19393,N_17022);
xnor UO_1016 (O_1016,N_15126,N_19202);
nor UO_1017 (O_1017,N_19051,N_19061);
nor UO_1018 (O_1018,N_18000,N_19130);
and UO_1019 (O_1019,N_17367,N_18108);
nand UO_1020 (O_1020,N_17413,N_19460);
or UO_1021 (O_1021,N_19532,N_16371);
nor UO_1022 (O_1022,N_19755,N_16358);
nand UO_1023 (O_1023,N_18438,N_15194);
nand UO_1024 (O_1024,N_16459,N_19413);
nor UO_1025 (O_1025,N_16262,N_16430);
nor UO_1026 (O_1026,N_17320,N_19442);
nand UO_1027 (O_1027,N_19323,N_19042);
and UO_1028 (O_1028,N_18564,N_18815);
and UO_1029 (O_1029,N_18121,N_15746);
nand UO_1030 (O_1030,N_19039,N_15266);
and UO_1031 (O_1031,N_17472,N_19640);
or UO_1032 (O_1032,N_15300,N_16904);
or UO_1033 (O_1033,N_18795,N_19447);
nor UO_1034 (O_1034,N_17868,N_19739);
nor UO_1035 (O_1035,N_16551,N_16806);
or UO_1036 (O_1036,N_16072,N_16707);
or UO_1037 (O_1037,N_17571,N_18247);
nand UO_1038 (O_1038,N_16814,N_16819);
nor UO_1039 (O_1039,N_15159,N_19523);
nor UO_1040 (O_1040,N_18923,N_16472);
or UO_1041 (O_1041,N_16621,N_16227);
nand UO_1042 (O_1042,N_19864,N_15457);
nand UO_1043 (O_1043,N_15257,N_18175);
and UO_1044 (O_1044,N_18214,N_19232);
nor UO_1045 (O_1045,N_15338,N_16810);
nor UO_1046 (O_1046,N_15893,N_18112);
xor UO_1047 (O_1047,N_16764,N_15255);
xor UO_1048 (O_1048,N_18810,N_15710);
nor UO_1049 (O_1049,N_16377,N_18177);
nor UO_1050 (O_1050,N_18098,N_17181);
nand UO_1051 (O_1051,N_18957,N_19559);
nand UO_1052 (O_1052,N_17293,N_17718);
and UO_1053 (O_1053,N_15562,N_17805);
nand UO_1054 (O_1054,N_15151,N_19197);
and UO_1055 (O_1055,N_16670,N_19815);
nand UO_1056 (O_1056,N_17256,N_18164);
nand UO_1057 (O_1057,N_17431,N_18984);
nand UO_1058 (O_1058,N_15957,N_15626);
nor UO_1059 (O_1059,N_19810,N_19923);
or UO_1060 (O_1060,N_17857,N_18034);
nor UO_1061 (O_1061,N_15589,N_17468);
or UO_1062 (O_1062,N_15701,N_18763);
or UO_1063 (O_1063,N_15871,N_19117);
nor UO_1064 (O_1064,N_15274,N_16278);
nor UO_1065 (O_1065,N_15501,N_19149);
or UO_1066 (O_1066,N_16010,N_15744);
xnor UO_1067 (O_1067,N_17104,N_15771);
nand UO_1068 (O_1068,N_19474,N_16400);
and UO_1069 (O_1069,N_15964,N_19336);
and UO_1070 (O_1070,N_17223,N_17790);
and UO_1071 (O_1071,N_16454,N_15258);
or UO_1072 (O_1072,N_17630,N_18013);
or UO_1073 (O_1073,N_16934,N_17175);
nand UO_1074 (O_1074,N_16100,N_17848);
nor UO_1075 (O_1075,N_18215,N_15683);
nor UO_1076 (O_1076,N_15176,N_19823);
and UO_1077 (O_1077,N_16579,N_18144);
nor UO_1078 (O_1078,N_18674,N_15679);
and UO_1079 (O_1079,N_15496,N_15741);
and UO_1080 (O_1080,N_18712,N_15250);
nor UO_1081 (O_1081,N_16285,N_16514);
or UO_1082 (O_1082,N_16219,N_18020);
or UO_1083 (O_1083,N_18402,N_17526);
or UO_1084 (O_1084,N_18248,N_16496);
and UO_1085 (O_1085,N_18100,N_18334);
and UO_1086 (O_1086,N_19867,N_15791);
and UO_1087 (O_1087,N_18142,N_16834);
or UO_1088 (O_1088,N_19978,N_17715);
nor UO_1089 (O_1089,N_18314,N_16088);
and UO_1090 (O_1090,N_16153,N_19806);
and UO_1091 (O_1091,N_15650,N_16038);
nand UO_1092 (O_1092,N_19011,N_18664);
nor UO_1093 (O_1093,N_18818,N_15998);
nand UO_1094 (O_1094,N_16989,N_18732);
nor UO_1095 (O_1095,N_17479,N_19144);
nand UO_1096 (O_1096,N_17834,N_17470);
nor UO_1097 (O_1097,N_17677,N_17359);
or UO_1098 (O_1098,N_16395,N_15908);
nor UO_1099 (O_1099,N_17315,N_15780);
and UO_1100 (O_1100,N_17082,N_18813);
and UO_1101 (O_1101,N_17680,N_19072);
xor UO_1102 (O_1102,N_16608,N_19274);
nand UO_1103 (O_1103,N_15063,N_15793);
and UO_1104 (O_1104,N_15565,N_18801);
or UO_1105 (O_1105,N_18448,N_16700);
nand UO_1106 (O_1106,N_16908,N_19891);
and UO_1107 (O_1107,N_15186,N_16717);
nand UO_1108 (O_1108,N_18876,N_15153);
and UO_1109 (O_1109,N_18914,N_18077);
and UO_1110 (O_1110,N_16343,N_19626);
nand UO_1111 (O_1111,N_15000,N_18670);
nand UO_1112 (O_1112,N_19888,N_18330);
nor UO_1113 (O_1113,N_16601,N_18052);
nor UO_1114 (O_1114,N_15610,N_17838);
nor UO_1115 (O_1115,N_18590,N_15422);
or UO_1116 (O_1116,N_18651,N_16452);
nand UO_1117 (O_1117,N_17955,N_16130);
nor UO_1118 (O_1118,N_17286,N_15541);
and UO_1119 (O_1119,N_17440,N_15462);
xnor UO_1120 (O_1120,N_17073,N_18502);
and UO_1121 (O_1121,N_18877,N_18325);
or UO_1122 (O_1122,N_19536,N_17480);
nor UO_1123 (O_1123,N_17362,N_17762);
nor UO_1124 (O_1124,N_16964,N_17106);
and UO_1125 (O_1125,N_15026,N_19518);
or UO_1126 (O_1126,N_19239,N_15486);
or UO_1127 (O_1127,N_19291,N_16924);
or UO_1128 (O_1128,N_18079,N_16893);
or UO_1129 (O_1129,N_18202,N_18503);
nor UO_1130 (O_1130,N_19234,N_19947);
or UO_1131 (O_1131,N_18453,N_15489);
nand UO_1132 (O_1132,N_19494,N_15523);
or UO_1133 (O_1133,N_15291,N_17685);
or UO_1134 (O_1134,N_19752,N_16941);
nand UO_1135 (O_1135,N_15184,N_19288);
nand UO_1136 (O_1136,N_16580,N_17032);
nand UO_1137 (O_1137,N_19696,N_16277);
or UO_1138 (O_1138,N_16730,N_16948);
or UO_1139 (O_1139,N_15578,N_15167);
or UO_1140 (O_1140,N_19634,N_16180);
and UO_1141 (O_1141,N_16223,N_16303);
or UO_1142 (O_1142,N_16852,N_18553);
and UO_1143 (O_1143,N_18816,N_15652);
nor UO_1144 (O_1144,N_17775,N_17306);
and UO_1145 (O_1145,N_18288,N_15066);
nor UO_1146 (O_1146,N_18212,N_15085);
and UO_1147 (O_1147,N_15052,N_15603);
nor UO_1148 (O_1148,N_16465,N_17693);
and UO_1149 (O_1149,N_18180,N_17228);
nand UO_1150 (O_1150,N_16662,N_16684);
and UO_1151 (O_1151,N_16509,N_16749);
nand UO_1152 (O_1152,N_17864,N_18548);
nand UO_1153 (O_1153,N_17423,N_15369);
and UO_1154 (O_1154,N_19369,N_18582);
nor UO_1155 (O_1155,N_18205,N_16821);
and UO_1156 (O_1156,N_17831,N_19384);
nand UO_1157 (O_1157,N_19631,N_17338);
nor UO_1158 (O_1158,N_18953,N_16687);
and UO_1159 (O_1159,N_17137,N_19198);
nor UO_1160 (O_1160,N_18540,N_15310);
or UO_1161 (O_1161,N_19936,N_16188);
nor UO_1162 (O_1162,N_18378,N_15513);
or UO_1163 (O_1163,N_16220,N_17867);
nand UO_1164 (O_1164,N_15730,N_16562);
nand UO_1165 (O_1165,N_17719,N_18092);
nor UO_1166 (O_1166,N_19666,N_18174);
nand UO_1167 (O_1167,N_18439,N_18324);
nor UO_1168 (O_1168,N_16909,N_17817);
and UO_1169 (O_1169,N_16536,N_15120);
nor UO_1170 (O_1170,N_18172,N_15776);
nand UO_1171 (O_1171,N_15941,N_16946);
and UO_1172 (O_1172,N_15409,N_19998);
nand UO_1173 (O_1173,N_17717,N_15921);
nand UO_1174 (O_1174,N_15601,N_16026);
nor UO_1175 (O_1175,N_18791,N_15588);
or UO_1176 (O_1176,N_15628,N_18975);
and UO_1177 (O_1177,N_16634,N_16000);
nor UO_1178 (O_1178,N_18710,N_16791);
or UO_1179 (O_1179,N_16573,N_15997);
or UO_1180 (O_1180,N_15688,N_19096);
nor UO_1181 (O_1181,N_15294,N_15260);
nor UO_1182 (O_1182,N_15609,N_16905);
nor UO_1183 (O_1183,N_15140,N_16256);
nand UO_1184 (O_1184,N_18316,N_15787);
and UO_1185 (O_1185,N_19773,N_17832);
or UO_1186 (O_1186,N_19742,N_16788);
xnor UO_1187 (O_1187,N_18859,N_16349);
and UO_1188 (O_1188,N_18945,N_19167);
and UO_1189 (O_1189,N_16281,N_19636);
and UO_1190 (O_1190,N_19141,N_15212);
nor UO_1191 (O_1191,N_16627,N_17220);
or UO_1192 (O_1192,N_19115,N_15129);
or UO_1193 (O_1193,N_17245,N_18437);
or UO_1194 (O_1194,N_18754,N_16312);
or UO_1195 (O_1195,N_19099,N_17425);
nor UO_1196 (O_1196,N_16009,N_19907);
nor UO_1197 (O_1197,N_17288,N_17491);
and UO_1198 (O_1198,N_18864,N_16265);
or UO_1199 (O_1199,N_18382,N_18315);
nand UO_1200 (O_1200,N_19967,N_17334);
or UO_1201 (O_1201,N_17896,N_17973);
or UO_1202 (O_1202,N_18765,N_16925);
and UO_1203 (O_1203,N_17264,N_17021);
nor UO_1204 (O_1204,N_16094,N_16146);
nand UO_1205 (O_1205,N_17519,N_18569);
nor UO_1206 (O_1206,N_19543,N_17899);
nand UO_1207 (O_1207,N_18363,N_19070);
and UO_1208 (O_1208,N_16694,N_18054);
or UO_1209 (O_1209,N_19108,N_16787);
nand UO_1210 (O_1210,N_16041,N_17157);
nand UO_1211 (O_1211,N_18137,N_16207);
or UO_1212 (O_1212,N_15657,N_19890);
and UO_1213 (O_1213,N_15190,N_15156);
and UO_1214 (O_1214,N_17214,N_16458);
or UO_1215 (O_1215,N_18870,N_19005);
or UO_1216 (O_1216,N_18644,N_19596);
nor UO_1217 (O_1217,N_16943,N_16737);
and UO_1218 (O_1218,N_18539,N_18061);
nand UO_1219 (O_1219,N_15004,N_15442);
nand UO_1220 (O_1220,N_18275,N_17730);
nand UO_1221 (O_1221,N_15797,N_17376);
or UO_1222 (O_1222,N_16493,N_16363);
or UO_1223 (O_1223,N_15333,N_18500);
or UO_1224 (O_1224,N_18411,N_17289);
and UO_1225 (O_1225,N_17506,N_18380);
nand UO_1226 (O_1226,N_16176,N_18989);
nor UO_1227 (O_1227,N_18270,N_18109);
and UO_1228 (O_1228,N_15916,N_15790);
or UO_1229 (O_1229,N_17839,N_17184);
nand UO_1230 (O_1230,N_19320,N_19168);
or UO_1231 (O_1231,N_16731,N_15475);
nor UO_1232 (O_1232,N_16525,N_18748);
nor UO_1233 (O_1233,N_15386,N_19302);
or UO_1234 (O_1234,N_16378,N_19517);
nand UO_1235 (O_1235,N_17962,N_18479);
nor UO_1236 (O_1236,N_17194,N_15123);
nor UO_1237 (O_1237,N_15118,N_18781);
nand UO_1238 (O_1238,N_16266,N_18064);
nand UO_1239 (O_1239,N_17404,N_19000);
nand UO_1240 (O_1240,N_15754,N_19312);
nand UO_1241 (O_1241,N_17008,N_18622);
or UO_1242 (O_1242,N_15323,N_18722);
nor UO_1243 (O_1243,N_17303,N_17185);
and UO_1244 (O_1244,N_15474,N_17331);
nor UO_1245 (O_1245,N_16151,N_19655);
and UO_1246 (O_1246,N_18915,N_19283);
nor UO_1247 (O_1247,N_17452,N_16161);
xnor UO_1248 (O_1248,N_18943,N_19276);
nor UO_1249 (O_1249,N_17496,N_18890);
and UO_1250 (O_1250,N_19625,N_18343);
and UO_1251 (O_1251,N_15861,N_17952);
nand UO_1252 (O_1252,N_15555,N_18377);
and UO_1253 (O_1253,N_18424,N_17527);
or UO_1254 (O_1254,N_16839,N_18617);
nand UO_1255 (O_1255,N_17593,N_19353);
and UO_1256 (O_1256,N_18240,N_16727);
and UO_1257 (O_1257,N_16780,N_19297);
or UO_1258 (O_1258,N_18229,N_17466);
or UO_1259 (O_1259,N_16353,N_18435);
nand UO_1260 (O_1260,N_19031,N_15130);
nand UO_1261 (O_1261,N_16293,N_18150);
or UO_1262 (O_1262,N_16420,N_18400);
nor UO_1263 (O_1263,N_18832,N_18720);
nand UO_1264 (O_1264,N_15699,N_19192);
and UO_1265 (O_1265,N_19155,N_16134);
xnor UO_1266 (O_1266,N_17535,N_17430);
nand UO_1267 (O_1267,N_15415,N_15143);
or UO_1268 (O_1268,N_17117,N_15342);
and UO_1269 (O_1269,N_15357,N_15831);
xnor UO_1270 (O_1270,N_18690,N_15396);
nand UO_1271 (O_1271,N_16446,N_19010);
nand UO_1272 (O_1272,N_18318,N_17930);
or UO_1273 (O_1273,N_19427,N_16524);
or UO_1274 (O_1274,N_18444,N_19789);
and UO_1275 (O_1275,N_16912,N_16445);
nor UO_1276 (O_1276,N_16878,N_18374);
nand UO_1277 (O_1277,N_18406,N_15920);
nor UO_1278 (O_1278,N_17590,N_18111);
nor UO_1279 (O_1279,N_17426,N_18065);
and UO_1280 (O_1280,N_17753,N_17392);
nor UO_1281 (O_1281,N_19357,N_15864);
nor UO_1282 (O_1282,N_16613,N_17325);
and UO_1283 (O_1283,N_17078,N_17683);
nor UO_1284 (O_1284,N_17284,N_17619);
nor UO_1285 (O_1285,N_19525,N_19580);
and UO_1286 (O_1286,N_19941,N_17398);
and UO_1287 (O_1287,N_18331,N_18027);
nor UO_1288 (O_1288,N_15851,N_15828);
nand UO_1289 (O_1289,N_19818,N_18320);
nand UO_1290 (O_1290,N_15835,N_15285);
nand UO_1291 (O_1291,N_18929,N_16044);
or UO_1292 (O_1292,N_18840,N_15762);
and UO_1293 (O_1293,N_16760,N_15922);
nand UO_1294 (O_1294,N_16453,N_19112);
and UO_1295 (O_1295,N_15722,N_15887);
nand UO_1296 (O_1296,N_19434,N_15505);
or UO_1297 (O_1297,N_18317,N_15647);
nand UO_1298 (O_1298,N_16315,N_19135);
or UO_1299 (O_1299,N_16068,N_15910);
nand UO_1300 (O_1300,N_19106,N_18641);
and UO_1301 (O_1301,N_18701,N_16401);
nand UO_1302 (O_1302,N_15512,N_15928);
and UO_1303 (O_1303,N_18604,N_15521);
or UO_1304 (O_1304,N_16511,N_16382);
or UO_1305 (O_1305,N_19527,N_19569);
or UO_1306 (O_1306,N_15358,N_19919);
nor UO_1307 (O_1307,N_16528,N_19787);
nor UO_1308 (O_1308,N_15636,N_19726);
and UO_1309 (O_1309,N_19462,N_15043);
nor UO_1310 (O_1310,N_17035,N_18413);
nand UO_1311 (O_1311,N_17312,N_18163);
and UO_1312 (O_1312,N_18344,N_18049);
or UO_1313 (O_1313,N_15169,N_15314);
nor UO_1314 (O_1314,N_15076,N_18044);
or UO_1315 (O_1315,N_15615,N_19863);
nor UO_1316 (O_1316,N_16162,N_17897);
or UO_1317 (O_1317,N_15777,N_18836);
nand UO_1318 (O_1318,N_17936,N_18599);
or UO_1319 (O_1319,N_16016,N_18312);
and UO_1320 (O_1320,N_16590,N_16635);
nand UO_1321 (O_1321,N_16913,N_16816);
and UO_1322 (O_1322,N_18654,N_19705);
or UO_1323 (O_1323,N_15949,N_18340);
nor UO_1324 (O_1324,N_17326,N_19848);
and UO_1325 (O_1325,N_19237,N_17729);
nand UO_1326 (O_1326,N_17749,N_15270);
nand UO_1327 (O_1327,N_19350,N_17420);
nand UO_1328 (O_1328,N_15408,N_19583);
nor UO_1329 (O_1329,N_19677,N_17394);
nand UO_1330 (O_1330,N_16520,N_17798);
or UO_1331 (O_1331,N_16286,N_19809);
or UO_1332 (O_1332,N_16759,N_16894);
and UO_1333 (O_1333,N_15443,N_17969);
nor UO_1334 (O_1334,N_16957,N_15690);
and UO_1335 (O_1335,N_17439,N_17776);
and UO_1336 (O_1336,N_15668,N_16732);
or UO_1337 (O_1337,N_16911,N_19632);
nor UO_1338 (O_1338,N_17577,N_16858);
nand UO_1339 (O_1339,N_18089,N_16864);
nand UO_1340 (O_1340,N_16099,N_18858);
xnor UO_1341 (O_1341,N_16251,N_15845);
or UO_1342 (O_1342,N_15740,N_18236);
nor UO_1343 (O_1343,N_15219,N_16135);
or UO_1344 (O_1344,N_18660,N_15827);
or UO_1345 (O_1345,N_16374,N_17090);
nor UO_1346 (O_1346,N_17145,N_18779);
and UO_1347 (O_1347,N_17894,N_19822);
nand UO_1348 (O_1348,N_16692,N_15543);
nand UO_1349 (O_1349,N_19528,N_16774);
nand UO_1350 (O_1350,N_15995,N_19230);
and UO_1351 (O_1351,N_16304,N_18373);
and UO_1352 (O_1352,N_15309,N_16396);
nor UO_1353 (O_1353,N_16428,N_17036);
and UO_1354 (O_1354,N_19069,N_17984);
and UO_1355 (O_1355,N_15434,N_18792);
nor UO_1356 (O_1356,N_17760,N_19126);
nor UO_1357 (O_1357,N_18652,N_17247);
nand UO_1358 (O_1358,N_19492,N_15103);
or UO_1359 (O_1359,N_17578,N_17333);
nand UO_1360 (O_1360,N_19500,N_19418);
or UO_1361 (O_1361,N_18436,N_16991);
nand UO_1362 (O_1362,N_15748,N_16049);
nor UO_1363 (O_1363,N_17960,N_15487);
nor UO_1364 (O_1364,N_17515,N_15247);
nand UO_1365 (O_1365,N_19767,N_15786);
and UO_1366 (O_1366,N_19821,N_16649);
or UO_1367 (O_1367,N_16217,N_16753);
nand UO_1368 (O_1368,N_17475,N_15639);
and UO_1369 (O_1369,N_19794,N_16863);
and UO_1370 (O_1370,N_19748,N_19614);
nand UO_1371 (O_1371,N_15820,N_16622);
nor UO_1372 (O_1372,N_18609,N_19592);
nand UO_1373 (O_1373,N_17110,N_19047);
or UO_1374 (O_1374,N_15718,N_16559);
and UO_1375 (O_1375,N_19610,N_19727);
and UO_1376 (O_1376,N_17731,N_19161);
and UO_1377 (O_1377,N_19706,N_16039);
or UO_1378 (O_1378,N_15445,N_18421);
and UO_1379 (O_1379,N_18843,N_17939);
or UO_1380 (O_1380,N_17234,N_17227);
or UO_1381 (O_1381,N_15518,N_18230);
or UO_1382 (O_1382,N_17836,N_16800);
nand UO_1383 (O_1383,N_17173,N_19328);
nor UO_1384 (O_1384,N_17244,N_19488);
and UO_1385 (O_1385,N_17594,N_18550);
and UO_1386 (O_1386,N_16876,N_16095);
nor UO_1387 (O_1387,N_18493,N_15760);
and UO_1388 (O_1388,N_19348,N_18192);
or UO_1389 (O_1389,N_19791,N_18733);
nor UO_1390 (O_1390,N_15316,N_19545);
nor UO_1391 (O_1391,N_17755,N_15370);
and UO_1392 (O_1392,N_19097,N_15455);
nand UO_1393 (O_1393,N_17970,N_19686);
nor UO_1394 (O_1394,N_15473,N_18974);
or UO_1395 (O_1395,N_17614,N_18888);
or UO_1396 (O_1396,N_18584,N_19964);
or UO_1397 (O_1397,N_19638,N_17485);
and UO_1398 (O_1398,N_17386,N_17539);
and UO_1399 (O_1399,N_18626,N_17495);
and UO_1400 (O_1400,N_16143,N_17434);
nand UO_1401 (O_1401,N_16540,N_15869);
and UO_1402 (O_1402,N_15498,N_16722);
or UO_1403 (O_1403,N_15006,N_15377);
nor UO_1404 (O_1404,N_16950,N_18518);
and UO_1405 (O_1405,N_16874,N_18347);
nand UO_1406 (O_1406,N_18936,N_15745);
xnor UO_1407 (O_1407,N_15514,N_18699);
or UO_1408 (O_1408,N_15706,N_17252);
or UO_1409 (O_1409,N_19858,N_17847);
and UO_1410 (O_1410,N_19697,N_16988);
nor UO_1411 (O_1411,N_18017,N_18029);
or UO_1412 (O_1412,N_18616,N_19253);
or UO_1413 (O_1413,N_18246,N_18485);
nor UO_1414 (O_1414,N_18785,N_19862);
and UO_1415 (O_1415,N_17996,N_19770);
nand UO_1416 (O_1416,N_17828,N_15372);
nor UO_1417 (O_1417,N_16383,N_17494);
nand UO_1418 (O_1418,N_16804,N_16054);
nand UO_1419 (O_1419,N_15024,N_17652);
nor UO_1420 (O_1420,N_17453,N_19699);
or UO_1421 (O_1421,N_16985,N_15202);
or UO_1422 (O_1422,N_16735,N_15334);
and UO_1423 (O_1423,N_16561,N_15901);
or UO_1424 (O_1424,N_17034,N_18659);
nor UO_1425 (O_1425,N_18545,N_18390);
nand UO_1426 (O_1426,N_15131,N_17737);
nand UO_1427 (O_1427,N_19264,N_16444);
and UO_1428 (O_1428,N_17168,N_19884);
or UO_1429 (O_1429,N_15863,N_17189);
nand UO_1430 (O_1430,N_16801,N_17741);
nand UO_1431 (O_1431,N_17912,N_16145);
and UO_1432 (O_1432,N_17763,N_17579);
nor UO_1433 (O_1433,N_17660,N_19950);
nand UO_1434 (O_1434,N_15703,N_19572);
nand UO_1435 (O_1435,N_16668,N_18512);
or UO_1436 (O_1436,N_18721,N_19058);
nand UO_1437 (O_1437,N_16150,N_19842);
nor UO_1438 (O_1438,N_16516,N_17356);
or UO_1439 (O_1439,N_15068,N_18016);
or UO_1440 (O_1440,N_19812,N_18561);
nand UO_1441 (O_1441,N_17915,N_19582);
nand UO_1442 (O_1442,N_19693,N_18682);
or UO_1443 (O_1443,N_16173,N_16320);
nand UO_1444 (O_1444,N_15238,N_15331);
or UO_1445 (O_1445,N_17860,N_18197);
nor UO_1446 (O_1446,N_18080,N_15209);
and UO_1447 (O_1447,N_18523,N_19549);
and UO_1448 (O_1448,N_15074,N_19828);
nor UO_1449 (O_1449,N_15822,N_17866);
nand UO_1450 (O_1450,N_19231,N_18170);
or UO_1451 (O_1451,N_15540,N_17914);
or UO_1452 (O_1452,N_16669,N_18841);
or UO_1453 (O_1453,N_19335,N_17825);
and UO_1454 (O_1454,N_16546,N_17002);
and UO_1455 (O_1455,N_17959,N_15163);
nand UO_1456 (O_1456,N_16247,N_17909);
nand UO_1457 (O_1457,N_17881,N_15188);
and UO_1458 (O_1458,N_19725,N_18190);
nor UO_1459 (O_1459,N_16456,N_18807);
or UO_1460 (O_1460,N_18169,N_16154);
or UO_1461 (O_1461,N_17965,N_19463);
nor UO_1462 (O_1462,N_17926,N_19872);
nor UO_1463 (O_1463,N_15290,N_15197);
and UO_1464 (O_1464,N_19645,N_17162);
or UO_1465 (O_1465,N_19660,N_19329);
and UO_1466 (O_1466,N_19269,N_17183);
or UO_1467 (O_1467,N_15233,N_19628);
nand UO_1468 (O_1468,N_19799,N_18973);
and UO_1469 (O_1469,N_15792,N_19673);
and UO_1470 (O_1470,N_19831,N_15775);
and UO_1471 (O_1471,N_18145,N_17756);
nand UO_1472 (O_1472,N_17672,N_16652);
or UO_1473 (O_1473,N_18761,N_17369);
or UO_1474 (O_1474,N_16415,N_17171);
or UO_1475 (O_1475,N_18798,N_17621);
or UO_1476 (O_1476,N_15622,N_17724);
and UO_1477 (O_1477,N_15926,N_19797);
and UO_1478 (O_1478,N_17129,N_18715);
nor UO_1479 (O_1479,N_17323,N_18963);
and UO_1480 (O_1480,N_16043,N_18058);
nand UO_1481 (O_1481,N_19199,N_17573);
or UO_1482 (O_1482,N_19132,N_19364);
and UO_1483 (O_1483,N_19651,N_18207);
or UO_1484 (O_1484,N_16584,N_17808);
nor UO_1485 (O_1485,N_15909,N_19593);
or UO_1486 (O_1486,N_16960,N_16750);
nor UO_1487 (O_1487,N_19562,N_16059);
nor UO_1488 (O_1488,N_17242,N_19701);
nor UO_1489 (O_1489,N_19415,N_18899);
and UO_1490 (O_1490,N_18072,N_19040);
or UO_1491 (O_1491,N_17580,N_17670);
or UO_1492 (O_1492,N_18126,N_15784);
nand UO_1493 (O_1493,N_17807,N_18873);
and UO_1494 (O_1494,N_15551,N_19608);
or UO_1495 (O_1495,N_17295,N_15538);
or UO_1496 (O_1496,N_19668,N_15782);
nor UO_1497 (O_1497,N_15567,N_15083);
or UO_1498 (O_1498,N_17989,N_15553);
nor UO_1499 (O_1499,N_16526,N_18580);
nand UO_1500 (O_1500,N_17597,N_19358);
nor UO_1501 (O_1501,N_17837,N_18298);
nand UO_1502 (O_1502,N_19330,N_16298);
or UO_1503 (O_1503,N_17006,N_17934);
nand UO_1504 (O_1504,N_18759,N_17455);
and UO_1505 (O_1505,N_19257,N_16414);
or UO_1506 (O_1506,N_16012,N_18194);
nand UO_1507 (O_1507,N_17437,N_17974);
nand UO_1508 (O_1508,N_15288,N_18143);
or UO_1509 (O_1509,N_18930,N_19351);
nand UO_1510 (O_1510,N_19154,N_15410);
nor UO_1511 (O_1511,N_18118,N_17099);
nor UO_1512 (O_1512,N_15527,N_16178);
or UO_1513 (O_1513,N_16479,N_15351);
nand UO_1514 (O_1514,N_17976,N_17603);
nor UO_1515 (O_1515,N_18496,N_17853);
nand UO_1516 (O_1516,N_16992,N_18615);
nor UO_1517 (O_1517,N_15199,N_19684);
nand UO_1518 (O_1518,N_15139,N_17028);
and UO_1519 (O_1519,N_19480,N_19704);
or UO_1520 (O_1520,N_17788,N_16714);
and UO_1521 (O_1521,N_19401,N_15234);
nor UO_1522 (O_1522,N_17046,N_15398);
or UO_1523 (O_1523,N_18277,N_17042);
or UO_1524 (O_1524,N_18026,N_19520);
or UO_1525 (O_1525,N_17014,N_15096);
and UO_1526 (O_1526,N_19653,N_19319);
and UO_1527 (O_1527,N_17133,N_19251);
and UO_1528 (O_1528,N_15426,N_15637);
and UO_1529 (O_1529,N_17071,N_18040);
nor UO_1530 (O_1530,N_18703,N_17319);
nor UO_1531 (O_1531,N_18460,N_16210);
or UO_1532 (O_1532,N_15208,N_19300);
and UO_1533 (O_1533,N_16919,N_18594);
nor UO_1534 (O_1534,N_19763,N_16771);
or UO_1535 (O_1535,N_16402,N_17257);
nor UO_1536 (O_1536,N_16898,N_15876);
or UO_1537 (O_1537,N_19382,N_15440);
or UO_1538 (O_1538,N_17147,N_15253);
or UO_1539 (O_1539,N_16197,N_17633);
xnor UO_1540 (O_1540,N_15449,N_15490);
or UO_1541 (O_1541,N_19849,N_15645);
or UO_1542 (O_1542,N_19067,N_18469);
and UO_1543 (O_1543,N_16101,N_17237);
or UO_1544 (O_1544,N_15675,N_15935);
nand UO_1545 (O_1545,N_15661,N_17626);
or UO_1546 (O_1546,N_15105,N_19441);
and UO_1547 (O_1547,N_18723,N_16794);
or UO_1548 (O_1548,N_19313,N_19383);
nand UO_1549 (O_1549,N_15363,N_17919);
nor UO_1550 (O_1550,N_19331,N_16024);
nor UO_1551 (O_1551,N_17746,N_19785);
or UO_1552 (O_1552,N_17774,N_17575);
nor UO_1553 (O_1553,N_16978,N_16880);
or UO_1554 (O_1554,N_17373,N_19175);
nor UO_1555 (O_1555,N_19189,N_15492);
and UO_1556 (O_1556,N_17349,N_15329);
and UO_1557 (O_1557,N_16603,N_16137);
nand UO_1558 (O_1558,N_18292,N_18736);
nand UO_1559 (O_1559,N_16182,N_16056);
or UO_1560 (O_1560,N_19825,N_17172);
and UO_1561 (O_1561,N_18505,N_18370);
nor UO_1562 (O_1562,N_19937,N_15282);
nor UO_1563 (O_1563,N_19203,N_15991);
nor UO_1564 (O_1564,N_15671,N_17553);
and UO_1565 (O_1565,N_19565,N_18835);
and UO_1566 (O_1566,N_16831,N_15407);
nor UO_1567 (O_1567,N_16469,N_16949);
nand UO_1568 (O_1568,N_17801,N_16492);
nand UO_1569 (O_1569,N_16915,N_16429);
nor UO_1570 (O_1570,N_17835,N_19055);
and UO_1571 (O_1571,N_15450,N_16723);
nand UO_1572 (O_1572,N_16063,N_17813);
nand UO_1573 (O_1573,N_15526,N_18856);
or UO_1574 (O_1574,N_19667,N_19766);
nor UO_1575 (O_1575,N_17714,N_17923);
and UO_1576 (O_1576,N_18522,N_15695);
nor UO_1577 (O_1577,N_17123,N_16890);
or UO_1578 (O_1578,N_15857,N_16477);
nand UO_1579 (O_1579,N_16110,N_15354);
nand UO_1580 (O_1580,N_17476,N_17773);
and UO_1581 (O_1581,N_19221,N_17190);
nor UO_1582 (O_1582,N_16965,N_17945);
nor UO_1583 (O_1583,N_17545,N_15961);
or UO_1584 (O_1584,N_15770,N_19454);
or UO_1585 (O_1585,N_18070,N_18937);
or UO_1586 (O_1586,N_16762,N_16018);
nand UO_1587 (O_1587,N_16471,N_16999);
or UO_1588 (O_1588,N_15716,N_18892);
and UO_1589 (O_1589,N_16870,N_15504);
and UO_1590 (O_1590,N_16518,N_18597);
nand UO_1591 (O_1591,N_18339,N_18244);
nor UO_1592 (O_1592,N_19308,N_19163);
nand UO_1593 (O_1593,N_15546,N_16437);
nand UO_1594 (O_1594,N_18095,N_18123);
or UO_1595 (O_1595,N_15481,N_16240);
or UO_1596 (O_1596,N_15399,N_15297);
nor UO_1597 (O_1597,N_19233,N_18139);
or UO_1598 (O_1598,N_18281,N_17536);
nor UO_1599 (O_1599,N_19377,N_16837);
nor UO_1600 (O_1600,N_17642,N_19332);
or UO_1601 (O_1601,N_16081,N_19561);
nand UO_1602 (O_1602,N_16235,N_15805);
nand UO_1603 (O_1603,N_15917,N_19897);
nand UO_1604 (O_1604,N_19469,N_19409);
nor UO_1605 (O_1605,N_19622,N_15689);
nand UO_1606 (O_1606,N_18440,N_17457);
nor UO_1607 (O_1607,N_16568,N_18527);
and UO_1608 (O_1608,N_16335,N_16360);
and UO_1609 (O_1609,N_16003,N_19247);
and UO_1610 (O_1610,N_16131,N_19733);
and UO_1611 (O_1611,N_15303,N_18427);
nand UO_1612 (O_1612,N_16097,N_19963);
nor UO_1613 (O_1613,N_19741,N_17791);
nand UO_1614 (O_1614,N_19513,N_17883);
and UO_1615 (O_1615,N_19458,N_18711);
and UO_1616 (O_1616,N_17599,N_18067);
and UO_1617 (O_1617,N_18501,N_19497);
and UO_1618 (O_1618,N_16354,N_18395);
nor UO_1619 (O_1619,N_17348,N_18178);
and UO_1620 (O_1620,N_15100,N_19411);
nand UO_1621 (O_1621,N_15174,N_18811);
and UO_1622 (O_1622,N_15466,N_17297);
or UO_1623 (O_1623,N_16531,N_17135);
nor UO_1624 (O_1624,N_17908,N_19063);
and UO_1625 (O_1625,N_17570,N_17159);
or UO_1626 (O_1626,N_19056,N_16824);
nor UO_1627 (O_1627,N_18432,N_16746);
nor UO_1628 (O_1628,N_17061,N_18593);
and UO_1629 (O_1629,N_15028,N_15374);
and UO_1630 (O_1630,N_15069,N_17523);
nor UO_1631 (O_1631,N_16677,N_18199);
and UO_1632 (O_1632,N_15141,N_17745);
and UO_1633 (O_1633,N_17793,N_18055);
or UO_1634 (O_1634,N_18666,N_16035);
or UO_1635 (O_1635,N_18552,N_19792);
or UO_1636 (O_1636,N_15482,N_17512);
nand UO_1637 (O_1637,N_15149,N_18097);
and UO_1638 (O_1638,N_19206,N_19618);
and UO_1639 (O_1639,N_16623,N_15193);
and UO_1640 (O_1640,N_18865,N_17396);
or UO_1641 (O_1641,N_16865,N_17013);
and UO_1642 (O_1642,N_16506,N_17195);
nand UO_1643 (O_1643,N_16990,N_18976);
nor UO_1644 (O_1644,N_16830,N_15915);
and UO_1645 (O_1645,N_17072,N_16861);
nand UO_1646 (O_1646,N_18931,N_16279);
and UO_1647 (O_1647,N_17231,N_17498);
and UO_1648 (O_1648,N_19675,N_18287);
or UO_1649 (O_1649,N_17639,N_16116);
nand UO_1650 (O_1650,N_18420,N_16330);
and UO_1651 (O_1651,N_15261,N_16639);
or UO_1652 (O_1652,N_16836,N_15394);
nand UO_1653 (O_1653,N_15621,N_15930);
or UO_1654 (O_1654,N_15378,N_19521);
nand UO_1655 (O_1655,N_19925,N_17803);
or UO_1656 (O_1656,N_19979,N_17503);
nor UO_1657 (O_1657,N_19551,N_15262);
xnor UO_1658 (O_1658,N_17100,N_17098);
nand UO_1659 (O_1659,N_18770,N_15162);
and UO_1660 (O_1660,N_17069,N_15550);
or UO_1661 (O_1661,N_17207,N_18216);
and UO_1662 (O_1662,N_17992,N_18249);
or UO_1663 (O_1663,N_18124,N_15371);
and UO_1664 (O_1664,N_19262,N_15182);
nand UO_1665 (O_1665,N_18002,N_17628);
nand UO_1666 (O_1666,N_18729,N_18384);
or UO_1667 (O_1667,N_19734,N_19339);
or UO_1668 (O_1668,N_16846,N_17169);
nor UO_1669 (O_1669,N_19430,N_16093);
nand UO_1670 (O_1670,N_19540,N_15684);
and UO_1671 (O_1671,N_16497,N_17294);
nor UO_1672 (O_1672,N_15039,N_15195);
and UO_1673 (O_1673,N_17001,N_19712);
nor UO_1674 (O_1674,N_15660,N_15630);
nand UO_1675 (O_1675,N_19663,N_19606);
or UO_1676 (O_1676,N_15648,N_17053);
nand UO_1677 (O_1677,N_19637,N_18585);
and UO_1678 (O_1678,N_18332,N_18555);
nor UO_1679 (O_1679,N_15146,N_17875);
nand UO_1680 (O_1680,N_16252,N_16963);
nand UO_1681 (O_1681,N_16969,N_16451);
nor UO_1682 (O_1682,N_17592,N_15107);
nand UO_1683 (O_1683,N_19555,N_19997);
and UO_1684 (O_1684,N_16510,N_16017);
or UO_1685 (O_1685,N_16900,N_16654);
xor UO_1686 (O_1686,N_18225,N_19844);
and UO_1687 (O_1687,N_18106,N_19387);
nand UO_1688 (O_1688,N_17954,N_19081);
and UO_1689 (O_1689,N_15510,N_15951);
nor UO_1690 (O_1690,N_15452,N_17854);
nor UO_1691 (O_1691,N_15698,N_19926);
nand UO_1692 (O_1692,N_19832,N_19624);
or UO_1693 (O_1693,N_19464,N_17768);
nand UO_1694 (O_1694,N_16195,N_16715);
and UO_1695 (O_1695,N_15965,N_18640);
or UO_1696 (O_1696,N_19970,N_16626);
nor UO_1697 (O_1697,N_16221,N_15021);
or UO_1698 (O_1698,N_19374,N_15714);
nor UO_1699 (O_1699,N_16236,N_18940);
and UO_1700 (O_1700,N_15579,N_18379);
nor UO_1701 (O_1701,N_15465,N_18021);
nor UO_1702 (O_1702,N_15427,N_18894);
or UO_1703 (O_1703,N_19229,N_16693);
nor UO_1704 (O_1704,N_19591,N_16555);
and UO_1705 (O_1705,N_17986,N_16802);
nand UO_1706 (O_1706,N_19294,N_17534);
or UO_1707 (O_1707,N_18120,N_19955);
and UO_1708 (O_1708,N_19456,N_15121);
nor UO_1709 (O_1709,N_15097,N_15721);
and UO_1710 (O_1710,N_18822,N_15677);
or UO_1711 (O_1711,N_19661,N_15664);
nand UO_1712 (O_1712,N_15263,N_18738);
and UO_1713 (O_1713,N_16166,N_19089);
and UO_1714 (O_1714,N_16703,N_18051);
nand UO_1715 (O_1715,N_15181,N_18757);
nand UO_1716 (O_1716,N_18487,N_16877);
or UO_1717 (O_1717,N_18506,N_18183);
nand UO_1718 (O_1718,N_18001,N_15712);
and UO_1719 (O_1719,N_17913,N_15335);
nor UO_1720 (O_1720,N_17144,N_15269);
nand UO_1721 (O_1721,N_15715,N_15704);
nand UO_1722 (O_1722,N_19399,N_17681);
and UO_1723 (O_1723,N_19751,N_19902);
and UO_1724 (O_1724,N_17548,N_17330);
or UO_1725 (O_1725,N_15547,N_18243);
nand UO_1726 (O_1726,N_17076,N_17951);
or UO_1727 (O_1727,N_18942,N_18771);
nor UO_1728 (O_1728,N_15384,N_15349);
nand UO_1729 (O_1729,N_19860,N_17419);
nor UO_1730 (O_1730,N_15727,N_15958);
nand UO_1731 (O_1731,N_19498,N_18282);
and UO_1732 (O_1732,N_19838,N_18326);
nor UO_1733 (O_1733,N_19635,N_15681);
xor UO_1734 (O_1734,N_18441,N_15458);
nand UO_1735 (O_1735,N_17884,N_19811);
nor UO_1736 (O_1736,N_19156,N_16724);
xnor UO_1737 (O_1737,N_16566,N_19289);
nand UO_1738 (O_1738,N_15558,N_18148);
or UO_1739 (O_1739,N_16862,N_18119);
nor UO_1740 (O_1740,N_15198,N_18224);
nand UO_1741 (O_1741,N_18507,N_19719);
nor UO_1742 (O_1742,N_19325,N_19385);
nor UO_1743 (O_1743,N_15898,N_16529);
and UO_1744 (O_1744,N_15757,N_17757);
nand UO_1745 (O_1745,N_17400,N_18693);
nor UO_1746 (O_1746,N_15330,N_15854);
nor UO_1747 (O_1747,N_15755,N_18927);
xnor UO_1748 (O_1748,N_18643,N_17581);
nand UO_1749 (O_1749,N_17738,N_18714);
nand UO_1750 (O_1750,N_19066,N_19969);
nor UO_1751 (O_1751,N_18023,N_19125);
or UO_1752 (O_1752,N_15952,N_19254);
nand UO_1753 (O_1753,N_17612,N_19139);
xor UO_1754 (O_1754,N_16222,N_18752);
nand UO_1755 (O_1755,N_15763,N_15846);
and UO_1756 (O_1756,N_17111,N_15980);
and UO_1757 (O_1757,N_19340,N_19356);
nor UO_1758 (O_1758,N_15036,N_18625);
and UO_1759 (O_1759,N_19146,N_19153);
and UO_1760 (O_1760,N_15048,N_18336);
nor UO_1761 (O_1761,N_15053,N_18784);
and UO_1762 (O_1762,N_18110,N_15738);
or UO_1763 (O_1763,N_18220,N_19644);
and UO_1764 (O_1764,N_17039,N_18204);
nand UO_1765 (O_1765,N_15148,N_18874);
and UO_1766 (O_1766,N_16888,N_19091);
or UO_1767 (O_1767,N_16263,N_16752);
nor UO_1768 (O_1768,N_18329,N_18993);
nor UO_1769 (O_1769,N_18962,N_15014);
nand UO_1770 (O_1770,N_18404,N_18494);
nor UO_1771 (O_1771,N_16102,N_19805);
nor UO_1772 (O_1772,N_16734,N_17298);
and UO_1773 (O_1773,N_17488,N_19983);
nor UO_1774 (O_1774,N_18147,N_19584);
and UO_1775 (O_1775,N_18218,N_15368);
and UO_1776 (O_1776,N_18035,N_18985);
and UO_1777 (O_1777,N_19407,N_19942);
or UO_1778 (O_1778,N_18551,N_16869);
nand UO_1779 (O_1779,N_15056,N_16385);
or UO_1780 (O_1780,N_15568,N_17921);
nor UO_1781 (O_1781,N_17054,N_17863);
and UO_1782 (O_1782,N_15687,N_19077);
or UO_1783 (O_1783,N_18728,N_15894);
nor UO_1784 (O_1784,N_18104,N_18136);
nor UO_1785 (O_1785,N_19426,N_17507);
and UO_1786 (O_1786,N_15343,N_19928);
nor UO_1787 (O_1787,N_16272,N_17066);
nand UO_1788 (O_1788,N_16848,N_18280);
or UO_1789 (O_1789,N_19930,N_17525);
and UO_1790 (O_1790,N_18233,N_19246);
nor UO_1791 (O_1791,N_16790,N_19688);
nor UO_1792 (O_1792,N_15625,N_18600);
or UO_1793 (O_1793,N_15424,N_18075);
nor UO_1794 (O_1794,N_17766,N_15089);
nand UO_1795 (O_1795,N_19901,N_18531);
and UO_1796 (O_1796,N_19366,N_16138);
nor UO_1797 (O_1797,N_19359,N_19363);
and UO_1798 (O_1798,N_15720,N_15819);
or UO_1799 (O_1799,N_19024,N_19477);
or UO_1800 (O_1800,N_17943,N_19993);
or UO_1801 (O_1801,N_17302,N_17174);
nor UO_1802 (O_1802,N_15425,N_16902);
nand UO_1803 (O_1803,N_17427,N_19911);
nand UO_1804 (O_1804,N_15271,N_19507);
nor UO_1805 (O_1805,N_15655,N_17366);
nor UO_1806 (O_1806,N_18515,N_18766);
and UO_1807 (O_1807,N_15885,N_15002);
and UO_1808 (O_1808,N_19749,N_15461);
nand UO_1809 (O_1809,N_15954,N_19586);
nand UO_1810 (O_1810,N_16144,N_18606);
nand UO_1811 (O_1811,N_16006,N_18602);
or UO_1812 (O_1812,N_17846,N_18826);
nor UO_1813 (O_1813,N_19589,N_16455);
and UO_1814 (O_1814,N_16046,N_17518);
nor UO_1815 (O_1815,N_15902,N_18450);
nor UO_1816 (O_1816,N_18718,N_16773);
nor UO_1817 (O_1817,N_16109,N_17720);
and UO_1818 (O_1818,N_16823,N_15999);
and UO_1819 (O_1819,N_19380,N_15355);
nor UO_1820 (O_1820,N_16615,N_19774);
or UO_1821 (O_1821,N_19243,N_16379);
and UO_1822 (O_1822,N_15900,N_19060);
nor UO_1823 (O_1823,N_16084,N_18434);
and UO_1824 (O_1824,N_15843,N_16352);
nand UO_1825 (O_1825,N_16535,N_19238);
nor UO_1826 (O_1826,N_15979,N_18162);
and UO_1827 (O_1827,N_16554,N_15707);
or UO_1828 (O_1828,N_16047,N_16793);
nand UO_1829 (O_1829,N_16541,N_17938);
nand UO_1830 (O_1830,N_16359,N_16828);
or UO_1831 (O_1831,N_15783,N_19008);
and UO_1832 (O_1832,N_15614,N_18193);
or UO_1833 (O_1833,N_18601,N_19417);
nor UO_1834 (O_1834,N_16288,N_19681);
or UO_1835 (O_1835,N_16961,N_18451);
or UO_1836 (O_1836,N_16388,N_18591);
and UO_1837 (O_1837,N_16500,N_15213);
nand UO_1838 (O_1838,N_15136,N_17251);
nand UO_1839 (O_1839,N_17946,N_17081);
and UO_1840 (O_1840,N_16473,N_19449);
nand UO_1841 (O_1841,N_16628,N_19920);
or UO_1842 (O_1842,N_16460,N_19324);
nand UO_1843 (O_1843,N_19041,N_19305);
nand UO_1844 (O_1844,N_15161,N_17122);
nand UO_1845 (O_1845,N_19547,N_19777);
and UO_1846 (O_1846,N_17305,N_19012);
nor UO_1847 (O_1847,N_17074,N_19307);
nand UO_1848 (O_1848,N_17353,N_18613);
nand UO_1849 (O_1849,N_18966,N_19895);
nor UO_1850 (O_1850,N_18880,N_19184);
nand UO_1851 (O_1851,N_19298,N_18886);
nand UO_1852 (O_1852,N_16841,N_18403);
or UO_1853 (O_1853,N_15278,N_16248);
nand UO_1854 (O_1854,N_15420,N_15403);
or UO_1855 (O_1855,N_15726,N_19143);
nor UO_1856 (O_1856,N_17360,N_18171);
nor UO_1857 (O_1857,N_15597,N_15984);
or UO_1858 (O_1858,N_18295,N_19994);
or UO_1859 (O_1859,N_16553,N_16742);
nor UO_1860 (O_1860,N_15923,N_19717);
nor UO_1861 (O_1861,N_18149,N_16721);
and UO_1862 (O_1862,N_16674,N_17703);
and UO_1863 (O_1863,N_19136,N_18516);
and UO_1864 (O_1864,N_17734,N_19030);
nor UO_1865 (O_1865,N_16681,N_17861);
nor UO_1866 (O_1866,N_18271,N_19285);
or UO_1867 (O_1867,N_16708,N_17467);
xnor UO_1868 (O_1868,N_16695,N_18794);
and UO_1869 (O_1869,N_19194,N_15116);
or UO_1870 (O_1870,N_18760,N_17510);
or UO_1871 (O_1871,N_17346,N_19013);
nand UO_1872 (O_1872,N_16691,N_19398);
and UO_1873 (O_1873,N_17641,N_18596);
or UO_1874 (O_1874,N_16271,N_18231);
nor UO_1875 (O_1875,N_18678,N_19103);
nand UO_1876 (O_1876,N_17705,N_19973);
or UO_1877 (O_1877,N_17011,N_16412);
nand UO_1878 (O_1878,N_19082,N_19976);
or UO_1879 (O_1879,N_18471,N_16104);
and UO_1880 (O_1880,N_17016,N_19687);
nor UO_1881 (O_1881,N_16029,N_16916);
nor UO_1882 (O_1882,N_17688,N_17565);
nor UO_1883 (O_1883,N_17787,N_18725);
or UO_1884 (O_1884,N_19817,N_16689);
and UO_1885 (O_1885,N_16838,N_15838);
or UO_1886 (O_1886,N_15485,N_18155);
or UO_1887 (O_1887,N_18556,N_16716);
or UO_1888 (O_1888,N_16709,N_17568);
nand UO_1889 (O_1889,N_17280,N_19682);
nand UO_1890 (O_1890,N_15225,N_19489);
nor UO_1891 (O_1891,N_15773,N_16650);
nand UO_1892 (O_1892,N_19486,N_18358);
nor UO_1893 (O_1893,N_17502,N_17876);
nor UO_1894 (O_1894,N_19680,N_17344);
nand UO_1895 (O_1895,N_18385,N_15117);
and UO_1896 (O_1896,N_15326,N_16165);
and UO_1897 (O_1897,N_18860,N_17968);
and UO_1898 (O_1898,N_16505,N_18950);
nor UO_1899 (O_1899,N_18359,N_19958);
or UO_1900 (O_1900,N_16896,N_18508);
and UO_1901 (O_1901,N_17692,N_18994);
xor UO_1902 (O_1902,N_19695,N_16855);
or UO_1903 (O_1903,N_15758,N_17903);
and UO_1904 (O_1904,N_16296,N_19800);
or UO_1905 (O_1905,N_16519,N_16261);
nor UO_1906 (O_1906,N_19982,N_19316);
nor UO_1907 (O_1907,N_19938,N_17521);
nand UO_1908 (O_1908,N_18920,N_15844);
nor UO_1909 (O_1909,N_19376,N_15600);
or UO_1910 (O_1910,N_16136,N_16468);
nand UO_1911 (O_1911,N_15839,N_17114);
or UO_1912 (O_1912,N_15245,N_16105);
or UO_1913 (O_1913,N_18741,N_16368);
nand UO_1914 (O_1914,N_16859,N_19301);
nand UO_1915 (O_1915,N_15943,N_17869);
nand UO_1916 (O_1916,N_17657,N_15280);
nor UO_1917 (O_1917,N_17241,N_16391);
nor UO_1918 (O_1918,N_16739,N_19775);
and UO_1919 (O_1919,N_16499,N_18242);
xnor UO_1920 (O_1920,N_18047,N_16712);
nor UO_1921 (O_1921,N_19793,N_18916);
nand UO_1922 (O_1922,N_19989,N_18219);
nand UO_1923 (O_1923,N_19801,N_18463);
nor UO_1924 (O_1924,N_17138,N_19674);
and UO_1925 (O_1925,N_16664,N_17871);
and UO_1926 (O_1926,N_18511,N_17025);
and UO_1927 (O_1927,N_16907,N_16958);
or UO_1928 (O_1928,N_18986,N_16119);
xor UO_1929 (O_1929,N_16917,N_16624);
or UO_1930 (O_1930,N_17964,N_17742);
and UO_1931 (O_1931,N_16501,N_19122);
nand UO_1932 (O_1932,N_16740,N_17933);
and UO_1933 (O_1933,N_17902,N_19918);
nor UO_1934 (O_1934,N_15086,N_18031);
nand UO_1935 (O_1935,N_15724,N_19001);
nor UO_1936 (O_1936,N_16698,N_19833);
and UO_1937 (O_1937,N_16331,N_18605);
nor UO_1938 (O_1938,N_19273,N_16431);
nand UO_1939 (O_1939,N_18408,N_16630);
and UO_1940 (O_1940,N_19988,N_17977);
nor UO_1941 (O_1941,N_16019,N_17567);
and UO_1942 (O_1942,N_16231,N_15672);
and UO_1943 (O_1943,N_15248,N_18266);
nor UO_1944 (O_1944,N_15866,N_18805);
xor UO_1945 (O_1945,N_18968,N_15669);
nand UO_1946 (O_1946,N_18869,N_15463);
and UO_1947 (O_1947,N_16993,N_16521);
nor UO_1948 (O_1948,N_17126,N_17850);
and UO_1949 (O_1949,N_19482,N_16947);
nand UO_1950 (O_1950,N_16494,N_17316);
or UO_1951 (O_1951,N_18279,N_19579);
nor UO_1952 (O_1952,N_16995,N_15892);
and UO_1953 (O_1953,N_16218,N_19195);
and UO_1954 (O_1954,N_18073,N_16257);
nor UO_1955 (O_1955,N_15044,N_17985);
nor UO_1956 (O_1956,N_19546,N_18900);
nor UO_1957 (O_1957,N_18680,N_18393);
or UO_1958 (O_1958,N_16643,N_15778);
nor UO_1959 (O_1959,N_18198,N_17274);
nand UO_1960 (O_1960,N_16155,N_16058);
nand UO_1961 (O_1961,N_19505,N_17886);
or UO_1962 (O_1962,N_17408,N_15858);
or UO_1963 (O_1963,N_16696,N_15651);
nand UO_1964 (O_1964,N_19337,N_16939);
or UO_1965 (O_1965,N_15599,N_18472);
nor UO_1966 (O_1966,N_19932,N_17931);
or UO_1967 (O_1967,N_17645,N_15632);
or UO_1968 (O_1968,N_16586,N_17109);
and UO_1969 (O_1969,N_19134,N_15988);
and UO_1970 (O_1970,N_15337,N_17018);
and UO_1971 (O_1971,N_16811,N_18925);
xor UO_1972 (O_1972,N_17781,N_19679);
and UO_1973 (O_1973,N_16879,N_19959);
and UO_1974 (O_1974,N_17115,N_15520);
and UO_1975 (O_1975,N_16329,N_18982);
nor UO_1976 (O_1976,N_15020,N_15729);
or UO_1977 (O_1977,N_17421,N_18954);
or UO_1978 (O_1978,N_18675,N_19444);
nor UO_1979 (O_1979,N_18634,N_19370);
nor UO_1980 (O_1980,N_15889,N_17089);
and UO_1981 (O_1981,N_15365,N_18082);
nor UO_1982 (O_1982,N_17975,N_19485);
nor UO_1983 (O_1983,N_18595,N_19043);
nand UO_1984 (O_1984,N_18375,N_15506);
or UO_1985 (O_1985,N_17799,N_17215);
and UO_1986 (O_1986,N_15104,N_16605);
nand UO_1987 (O_1987,N_17483,N_17176);
or UO_1988 (O_1988,N_15220,N_15483);
nand UO_1989 (O_1989,N_15239,N_16164);
nor UO_1990 (O_1990,N_17478,N_19303);
nand UO_1991 (O_1991,N_17812,N_17151);
and UO_1992 (O_1992,N_18428,N_18041);
nand UO_1993 (O_1993,N_15799,N_16413);
or UO_1994 (O_1994,N_15324,N_17998);
nand UO_1995 (O_1995,N_19537,N_17308);
or UO_1996 (O_1996,N_18862,N_16476);
and UO_1997 (O_1997,N_17554,N_17155);
nor UO_1998 (O_1998,N_16563,N_15811);
or UO_1999 (O_1999,N_15494,N_17988);
or UO_2000 (O_2000,N_18775,N_15292);
nand UO_2001 (O_2001,N_17721,N_17967);
xnor UO_2002 (O_2002,N_15388,N_16792);
or UO_2003 (O_2003,N_15187,N_15572);
and UO_2004 (O_2004,N_15815,N_16369);
nor UO_2005 (O_2005,N_19222,N_18995);
nand UO_2006 (O_2006,N_17910,N_16720);
and UO_2007 (O_2007,N_15649,N_16705);
or UO_2008 (O_2008,N_17656,N_19708);
or UO_2009 (O_2009,N_18006,N_19616);
xnor UO_2010 (O_2010,N_17751,N_19934);
or UO_2011 (O_2011,N_19803,N_17687);
or UO_2012 (O_2012,N_16548,N_18875);
and UO_2013 (O_2013,N_17880,N_18381);
nand UO_2014 (O_2014,N_18519,N_16152);
and UO_2015 (O_2015,N_18799,N_15133);
or UO_2016 (O_2016,N_18646,N_19731);
nand UO_2017 (O_2017,N_19908,N_15192);
and UO_2018 (O_2018,N_16132,N_16483);
nand UO_2019 (O_2019,N_15953,N_15214);
nor UO_2020 (O_2020,N_17591,N_19496);
or UO_2021 (O_2021,N_15158,N_18365);
and UO_2022 (O_2022,N_18455,N_17627);
or UO_2023 (O_2023,N_17927,N_15109);
and UO_2024 (O_2024,N_19652,N_15067);
and UO_2025 (O_2025,N_17314,N_18464);
nor UO_2026 (O_2026,N_18902,N_17196);
and UO_2027 (O_2027,N_19445,N_19185);
and UO_2028 (O_2028,N_15346,N_16955);
nor UO_2029 (O_2029,N_19076,N_16289);
nor UO_2030 (O_2030,N_17901,N_17444);
and UO_2031 (O_2031,N_16686,N_16868);
nor UO_2032 (O_2032,N_16351,N_16125);
or UO_2033 (O_2033,N_15286,N_18173);
or UO_2034 (O_2034,N_19075,N_18153);
nand UO_2035 (O_2035,N_15172,N_19698);
and UO_2036 (O_2036,N_18941,N_16070);
and UO_2037 (O_2037,N_16238,N_15177);
xnor UO_2038 (O_2038,N_17277,N_16394);
nand UO_2039 (O_2039,N_16552,N_18913);
nand UO_2040 (O_2040,N_17797,N_15767);
nor UO_2041 (O_2041,N_18947,N_15264);
nand UO_2042 (O_2042,N_17433,N_15345);
nand UO_2043 (O_2043,N_17243,N_15061);
and UO_2044 (O_2044,N_17629,N_15837);
nor UO_2045 (O_2045,N_19995,N_15018);
and UO_2046 (O_2046,N_19478,N_15516);
nand UO_2047 (O_2047,N_16255,N_17497);
or UO_2048 (O_2048,N_17979,N_18918);
nor UO_2049 (O_2049,N_17528,N_15088);
and UO_2050 (O_2050,N_16596,N_18181);
nor UO_2051 (O_2051,N_16183,N_17128);
or UO_2052 (O_2052,N_18653,N_16028);
nor UO_2053 (O_2053,N_15268,N_15138);
nand UO_2054 (O_2054,N_17596,N_15823);
and UO_2055 (O_2055,N_17644,N_18416);
and UO_2056 (O_2056,N_19557,N_15421);
or UO_2057 (O_2057,N_18744,N_18274);
nand UO_2058 (O_2058,N_17269,N_17625);
or UO_2059 (O_2059,N_17332,N_16927);
nand UO_2060 (O_2060,N_18684,N_18833);
nor UO_2061 (O_2061,N_18981,N_18978);
nor UO_2062 (O_2062,N_17796,N_17300);
or UO_2063 (O_2063,N_16141,N_19648);
and UO_2064 (O_2064,N_15653,N_17948);
nor UO_2065 (O_2065,N_17598,N_15431);
and UO_2066 (O_2066,N_16809,N_16663);
nor UO_2067 (O_2067,N_15563,N_16967);
and UO_2068 (O_2068,N_19165,N_18255);
nor UO_2069 (O_2069,N_19466,N_19275);
nand UO_2070 (O_2070,N_17564,N_17230);
and UO_2071 (O_2071,N_17381,N_19009);
or UO_2072 (O_2072,N_18649,N_16260);
or UO_2073 (O_2073,N_17544,N_19744);
nor UO_2074 (O_2074,N_19707,N_16944);
and UO_2075 (O_2075,N_16202,N_17877);
or UO_2076 (O_2076,N_17009,N_19263);
nor UO_2077 (O_2077,N_19405,N_17640);
nor UO_2078 (O_2078,N_18135,N_17638);
nor UO_2079 (O_2079,N_17291,N_18618);
or UO_2080 (O_2080,N_18814,N_15678);
xor UO_2081 (O_2081,N_16406,N_15975);
or UO_2082 (O_2082,N_18688,N_16594);
or UO_2083 (O_2083,N_15662,N_19062);
nor UO_2084 (O_2084,N_15591,N_19086);
nand UO_2085 (O_2085,N_17676,N_15976);
nor UO_2086 (O_2086,N_16086,N_17235);
nand UO_2087 (O_2087,N_15301,N_17940);
and UO_2088 (O_2088,N_17226,N_17309);
nor UO_2089 (O_2089,N_18008,N_19935);
nand UO_2090 (O_2090,N_19400,N_18267);
and UO_2091 (O_2091,N_16249,N_15676);
nand UO_2092 (O_2092,N_19014,N_19882);
and UO_2093 (O_2093,N_19057,N_19455);
nor UO_2094 (O_2094,N_19352,N_15010);
nand UO_2095 (O_2095,N_17149,N_16314);
nand UO_2096 (O_2096,N_15047,N_18168);
nor UO_2097 (O_2097,N_18924,N_15232);
and UO_2098 (O_2098,N_17563,N_19116);
and UO_2099 (O_2099,N_16213,N_16569);
and UO_2100 (O_2100,N_19757,N_17317);
and UO_2101 (O_2101,N_17070,N_17655);
nor UO_2102 (O_2102,N_16073,N_17205);
nand UO_2103 (O_2103,N_17551,N_15124);
nor UO_2104 (O_2104,N_16938,N_19974);
nor UO_2105 (O_2105,N_15764,N_17204);
nand UO_2106 (O_2106,N_19079,N_18176);
nor UO_2107 (O_2107,N_19594,N_17140);
or UO_2108 (O_2108,N_19670,N_18842);
nor UO_2109 (O_2109,N_15554,N_19782);
or UO_2110 (O_2110,N_17795,N_16294);
or UO_2111 (O_2111,N_18087,N_17370);
and UO_2112 (O_2112,N_15144,N_17351);
or UO_2113 (O_2113,N_18707,N_17963);
or UO_2114 (O_2114,N_15800,N_19916);
xor UO_2115 (O_2115,N_16316,N_16631);
or UO_2116 (O_2116,N_19088,N_16733);
and UO_2117 (O_2117,N_15359,N_19605);
xor UO_2118 (O_2118,N_17508,N_16718);
nor UO_2119 (O_2119,N_17489,N_19945);
or UO_2120 (O_2120,N_19981,N_18113);
nand UO_2121 (O_2121,N_16325,N_15733);
nand UO_2122 (O_2122,N_19879,N_19944);
or UO_2123 (O_2123,N_18706,N_19662);
nand UO_2124 (O_2124,N_18544,N_16034);
nor UO_2125 (O_2125,N_18788,N_17532);
or UO_2126 (O_2126,N_18290,N_16827);
and UO_2127 (O_2127,N_17221,N_15968);
or UO_2128 (O_2128,N_15246,N_16448);
nand UO_2129 (O_2129,N_16069,N_15395);
and UO_2130 (O_2130,N_15179,N_16242);
nand UO_2131 (O_2131,N_19595,N_18015);
and UO_2132 (O_2132,N_15785,N_15390);
nand UO_2133 (O_2133,N_18756,N_15299);
nor UO_2134 (O_2134,N_15873,N_18944);
xnor UO_2135 (O_2135,N_18254,N_16434);
nand UO_2136 (O_2136,N_17651,N_17424);
or UO_2137 (O_2137,N_19465,N_18443);
nand UO_2138 (O_2138,N_19311,N_16042);
nand UO_2139 (O_2139,N_17684,N_18185);
nor UO_2140 (O_2140,N_18201,N_16381);
nor UO_2141 (O_2141,N_16997,N_18921);
and UO_2142 (O_2142,N_18465,N_15222);
and UO_2143 (O_2143,N_17397,N_18776);
or UO_2144 (O_2144,N_17161,N_16140);
or UO_2145 (O_2145,N_19769,N_19996);
and UO_2146 (O_2146,N_17167,N_19850);
and UO_2147 (O_2147,N_16860,N_19526);
nor UO_2148 (O_2148,N_19159,N_16545);
nand UO_2149 (O_2149,N_19683,N_16066);
nand UO_2150 (O_2150,N_16507,N_17769);
and UO_2151 (O_2151,N_17318,N_18057);
and UO_2152 (O_2152,N_18872,N_19023);
nand UO_2153 (O_2153,N_16280,N_19603);
and UO_2154 (O_2154,N_17377,N_18513);
xnor UO_2155 (O_2155,N_15341,N_19900);
nand UO_2156 (O_2156,N_19881,N_18152);
and UO_2157 (O_2157,N_17664,N_19470);
and UO_2158 (O_2158,N_18661,N_19182);
or UO_2159 (O_2159,N_15830,N_19461);
xor UO_2160 (O_2160,N_18639,N_18115);
nor UO_2161 (O_2161,N_17473,N_17212);
nand UO_2162 (O_2162,N_18764,N_19597);
or UO_2163 (O_2163,N_16910,N_19368);
or UO_2164 (O_2164,N_19021,N_16849);
and UO_2165 (O_2165,N_16783,N_18284);
nand UO_2166 (O_2166,N_19511,N_15556);
nand UO_2167 (O_2167,N_17290,N_18477);
and UO_2168 (O_2168,N_19743,N_17562);
nand UO_2169 (O_2169,N_17673,N_17177);
or UO_2170 (O_2170,N_16480,N_15743);
nand UO_2171 (O_2171,N_19171,N_19737);
nand UO_2172 (O_2172,N_17232,N_18062);
and UO_2173 (O_2173,N_19720,N_17103);
or UO_2174 (O_2174,N_18071,N_17789);
nand UO_2175 (O_2175,N_19870,N_18901);
nand UO_2176 (O_2176,N_17905,N_15834);
and UO_2177 (O_2177,N_17706,N_19790);
nor UO_2178 (O_2178,N_16083,N_18882);
and UO_2179 (O_2179,N_17994,N_19504);
nand UO_2180 (O_2180,N_18904,N_17739);
nor UO_2181 (O_2181,N_15218,N_16112);
nor UO_2182 (O_2182,N_17833,N_18991);
or UO_2183 (O_2183,N_15717,N_16290);
nand UO_2184 (O_2184,N_18237,N_16564);
or UO_2185 (O_2185,N_16970,N_17631);
nand UO_2186 (O_2186,N_17675,N_19912);
and UO_2187 (O_2187,N_18350,N_18558);
or UO_2188 (O_2188,N_19985,N_18486);
nor UO_2189 (O_2189,N_15549,N_18346);
or UO_2190 (O_2190,N_16397,N_18834);
or UO_2191 (O_2191,N_15315,N_15227);
nor UO_2192 (O_2192,N_18499,N_16128);
nor UO_2193 (O_2193,N_16761,N_19612);
nand UO_2194 (O_2194,N_18611,N_19102);
nand UO_2195 (O_2195,N_19499,N_19939);
or UO_2196 (O_2196,N_16882,N_19240);
or UO_2197 (O_2197,N_18313,N_15032);
or UO_2198 (O_2198,N_16274,N_15617);
nand UO_2199 (O_2199,N_18713,N_18844);
and UO_2200 (O_2200,N_17650,N_19566);
and UO_2201 (O_2201,N_19260,N_17282);
or UO_2202 (O_2202,N_17165,N_15613);
nor UO_2203 (O_2203,N_19506,N_16935);
nor UO_2204 (O_2204,N_17040,N_16111);
nor UO_2205 (O_2205,N_17030,N_18399);
nand UO_2206 (O_2206,N_15387,N_16168);
or UO_2207 (O_2207,N_16968,N_16053);
nand UO_2208 (O_2208,N_18293,N_16389);
or UO_2209 (O_2209,N_17260,N_18388);
and UO_2210 (O_2210,N_19446,N_18576);
nor UO_2211 (O_2211,N_18509,N_15251);
or UO_2212 (O_2212,N_18830,N_15633);
nand UO_2213 (O_2213,N_19218,N_18417);
or UO_2214 (O_2214,N_19396,N_19479);
nand UO_2215 (O_2215,N_15646,N_18426);
and UO_2216 (O_2216,N_17239,N_16027);
or UO_2217 (O_2217,N_17384,N_19212);
or UO_2218 (O_2218,N_19702,N_18592);
nand UO_2219 (O_2219,N_17842,N_19909);
nor UO_2220 (O_2220,N_19084,N_17211);
nor UO_2221 (O_2221,N_18132,N_19450);
and UO_2222 (O_2222,N_15640,N_17646);
or UO_2223 (O_2223,N_16881,N_16704);
and UO_2224 (O_2224,N_18635,N_18817);
or UO_2225 (O_2225,N_17064,N_15224);
nand UO_2226 (O_2226,N_18396,N_16578);
or UO_2227 (O_2227,N_17154,N_18629);
nand UO_2228 (O_2228,N_17890,N_16341);
or UO_2229 (O_2229,N_18304,N_18956);
or UO_2230 (O_2230,N_19050,N_18228);
nor UO_2231 (O_2231,N_16313,N_19268);
nor UO_2232 (O_2232,N_15899,N_18809);
or UO_2233 (O_2233,N_19804,N_15340);
nor UO_2234 (O_2234,N_16503,N_17233);
or UO_2235 (O_2235,N_18951,N_18867);
nand UO_2236 (O_2236,N_16245,N_15373);
nand UO_2237 (O_2237,N_15287,N_16755);
or UO_2238 (O_2238,N_17830,N_18677);
and UO_2239 (O_2239,N_16435,N_18825);
nand UO_2240 (O_2240,N_17462,N_19105);
nor UO_2241 (O_2241,N_19929,N_18734);
or UO_2242 (O_2242,N_17806,N_19318);
nand UO_2243 (O_2243,N_19049,N_16177);
nor UO_2244 (O_2244,N_15903,N_16618);
and UO_2245 (O_2245,N_19390,N_19854);
or UO_2246 (O_2246,N_19834,N_16867);
and UO_2247 (O_2247,N_18922,N_18323);
or UO_2248 (O_2248,N_18038,N_16319);
or UO_2249 (O_2249,N_19349,N_17712);
or UO_2250 (O_2250,N_18291,N_19965);
or UO_2251 (O_2251,N_16812,N_16167);
or UO_2252 (O_2252,N_15686,N_18376);
or UO_2253 (O_2253,N_15631,N_19068);
nand UO_2254 (O_2254,N_15663,N_18967);
nor UO_2255 (O_2255,N_18037,N_17048);
and UO_2256 (O_2256,N_19856,N_17092);
or UO_2257 (O_2257,N_15302,N_15200);
nand UO_2258 (O_2258,N_15376,N_17259);
nand UO_2259 (O_2259,N_18354,N_18419);
nand UO_2260 (O_2260,N_17163,N_15581);
nor UO_2261 (O_2261,N_15040,N_17026);
nand UO_2262 (O_2262,N_16986,N_15605);
nand UO_2263 (O_2263,N_18367,N_16340);
and UO_2264 (O_2264,N_18566,N_19293);
nand UO_2265 (O_2265,N_16996,N_17671);
or UO_2266 (O_2266,N_16971,N_15821);
nor UO_2267 (O_2267,N_15488,N_17643);
nand UO_2268 (O_2268,N_16092,N_17027);
and UO_2269 (O_2269,N_17777,N_18462);
nor UO_2270 (O_2270,N_19816,N_19922);
nor UO_2271 (O_2271,N_15298,N_18107);
or UO_2272 (O_2272,N_17164,N_15759);
and UO_2273 (O_2273,N_18853,N_19992);
nor UO_2274 (O_2274,N_18863,N_18258);
and UO_2275 (O_2275,N_17809,N_15872);
nand UO_2276 (O_2276,N_19054,N_19287);
nor UO_2277 (O_2277,N_19166,N_15135);
and UO_2278 (O_2278,N_16945,N_18717);
and UO_2279 (O_2279,N_16023,N_18742);
or UO_2280 (O_2280,N_17414,N_16085);
and UO_2281 (O_2281,N_18735,N_18352);
nand UO_2282 (O_2282,N_18099,N_17415);
or UO_2283 (O_2283,N_18250,N_15641);
nor UO_2284 (O_2284,N_17764,N_17500);
nand UO_2285 (O_2285,N_19412,N_19034);
and UO_2286 (O_2286,N_17158,N_17132);
nor UO_2287 (O_2287,N_18452,N_16244);
and UO_2288 (O_2288,N_18687,N_18007);
and UO_2289 (O_2289,N_17160,N_17393);
and UO_2290 (O_2290,N_15081,N_19889);
and UO_2291 (O_2291,N_18685,N_19016);
and UO_2292 (O_2292,N_17659,N_17254);
nand UO_2293 (O_2293,N_19204,N_16770);
and UO_2294 (O_2294,N_15201,N_15624);
or UO_2295 (O_2295,N_15768,N_17574);
nor UO_2296 (O_2296,N_19830,N_19083);
or UO_2297 (O_2297,N_16215,N_15472);
nor UO_2298 (O_2298,N_19843,N_19627);
and UO_2299 (O_2299,N_18338,N_18273);
or UO_2300 (O_2300,N_17522,N_19795);
and UO_2301 (O_2301,N_19508,N_15971);
nand UO_2302 (O_2302,N_17708,N_17368);
nand UO_2303 (O_2303,N_18730,N_16914);
nand UO_2304 (O_2304,N_19342,N_17170);
and UO_2305 (O_2305,N_16538,N_16300);
and UO_2306 (O_2306,N_15803,N_19059);
nor UO_2307 (O_2307,N_17516,N_19394);
and UO_2308 (O_2308,N_15479,N_15598);
or UO_2309 (O_2309,N_17689,N_17849);
and UO_2310 (O_2310,N_18186,N_16743);
nand UO_2311 (O_2311,N_15049,N_18445);
and UO_2312 (O_2312,N_16175,N_19481);
nand UO_2313 (O_2313,N_15884,N_18208);
nand UO_2314 (O_2314,N_16157,N_16123);
nor UO_2315 (O_2315,N_16399,N_15945);
nor UO_2316 (O_2316,N_16356,N_19865);
nor UO_2317 (O_2317,N_15852,N_16126);
or UO_2318 (O_2318,N_15339,N_16463);
or UO_2319 (O_2319,N_19157,N_16930);
nand UO_2320 (O_2320,N_18196,N_16973);
nand UO_2321 (O_2321,N_16129,N_17047);
and UO_2322 (O_2322,N_17055,N_19915);
and UO_2323 (O_2323,N_16417,N_19802);
nor UO_2324 (O_2324,N_15736,N_17253);
nand UO_2325 (O_2325,N_19002,N_17024);
nand UO_2326 (O_2326,N_15580,N_16214);
nor UO_2327 (O_2327,N_19643,N_17044);
nor UO_2328 (O_2328,N_18769,N_17091);
nand UO_2329 (O_2329,N_17358,N_17406);
nand UO_2330 (O_2330,N_18299,N_16611);
or UO_2331 (O_2331,N_16013,N_15055);
nor UO_2332 (O_2332,N_18562,N_16744);
and UO_2333 (O_2333,N_15183,N_18700);
nand UO_2334 (O_2334,N_16490,N_16321);
or UO_2335 (O_2335,N_15867,N_17767);
or UO_2336 (O_2336,N_17844,N_19510);
nor UO_2337 (O_2337,N_16778,N_18086);
nor UO_2338 (O_2338,N_18802,N_16779);
and UO_2339 (O_2339,N_15749,N_19722);
nand UO_2340 (O_2340,N_15433,N_17972);
and UO_2341 (O_2341,N_17716,N_16239);
nor UO_2342 (O_2342,N_17942,N_18297);
nand UO_2343 (O_2343,N_15385,N_19853);
nor UO_2344 (O_2344,N_16163,N_17653);
or UO_2345 (O_2345,N_18217,N_18256);
nor UO_2346 (O_2346,N_17255,N_17191);
and UO_2347 (O_2347,N_18048,N_19808);
nor UO_2348 (O_2348,N_16246,N_17916);
or UO_2349 (O_2349,N_19109,N_17083);
nor UO_2350 (O_2350,N_19334,N_17458);
nand UO_2351 (O_2351,N_16232,N_19574);
or UO_2352 (O_2352,N_19953,N_18851);
or UO_2353 (O_2353,N_18468,N_17615);
nor UO_2354 (O_2354,N_17278,N_17845);
and UO_2355 (O_2355,N_15602,N_18009);
nand UO_2356 (O_2356,N_17240,N_18005);
nor UO_2357 (O_2357,N_15987,N_15313);
and UO_2358 (O_2358,N_19819,N_16295);
nor UO_2359 (O_2359,N_19948,N_15659);
or UO_2360 (O_2360,N_17735,N_18478);
nand UO_2361 (O_2361,N_19827,N_15911);
nor UO_2362 (O_2362,N_17616,N_18960);
and UO_2363 (O_2363,N_17632,N_16057);
nor UO_2364 (O_2364,N_16523,N_19472);
nand UO_2365 (O_2365,N_19421,N_17560);
nand UO_2366 (O_2366,N_15583,N_15694);
nor UO_2367 (O_2367,N_18696,N_15419);
nor UO_2368 (O_2368,N_17893,N_19875);
nor UO_2369 (O_2369,N_15751,N_17823);
and UO_2370 (O_2370,N_16007,N_18490);
and UO_2371 (O_2371,N_19375,N_16847);
nand UO_2372 (O_2372,N_16785,N_17339);
nor UO_2373 (O_2373,N_17382,N_15441);
and UO_2374 (O_2374,N_18357,N_18887);
nor UO_2375 (O_2375,N_18032,N_15544);
nand UO_2376 (O_2376,N_16577,N_19617);
nor UO_2377 (O_2377,N_15164,N_16422);
and UO_2378 (O_2378,N_15115,N_15596);
nor UO_2379 (O_2379,N_17213,N_19747);
nand UO_2380 (O_2380,N_17611,N_17530);
nor UO_2381 (O_2381,N_18891,N_18076);
nor UO_2382 (O_2382,N_18583,N_16243);
or UO_2383 (O_2383,N_17723,N_19052);
nor UO_2384 (O_2384,N_18353,N_18543);
nand UO_2385 (O_2385,N_16975,N_15160);
and UO_2386 (O_2386,N_17537,N_19094);
or UO_2387 (O_2387,N_15380,N_16048);
nor UO_2388 (O_2388,N_17311,N_15989);
nor UO_2389 (O_2389,N_18547,N_19980);
nand UO_2390 (O_2390,N_19516,N_19917);
nor UO_2391 (O_2391,N_19422,N_19868);
nand UO_2392 (O_2392,N_16299,N_15009);
nor UO_2393 (O_2393,N_17095,N_19571);
and UO_2394 (O_2394,N_17900,N_18739);
and UO_2395 (O_2395,N_18632,N_19228);
and UO_2396 (O_2396,N_16393,N_18638);
xor UO_2397 (O_2397,N_18311,N_19372);
and UO_2398 (O_2398,N_17050,N_17037);
and UO_2399 (O_2399,N_19473,N_15173);
nor UO_2400 (O_2400,N_17816,N_17225);
or UO_2401 (O_2401,N_15517,N_17941);
or UO_2402 (O_2402,N_16768,N_16789);
nor UO_2403 (O_2403,N_16032,N_18184);
nand UO_2404 (O_2404,N_19601,N_15670);
nand UO_2405 (O_2405,N_16527,N_18932);
or UO_2406 (O_2406,N_18014,N_17888);
nor UO_2407 (O_2407,N_18535,N_17275);
nand UO_2408 (O_2408,N_19689,N_18829);
nand UO_2409 (O_2409,N_19004,N_15092);
nand UO_2410 (O_2410,N_17784,N_16850);
nor UO_2411 (O_2411,N_17271,N_19570);
or UO_2412 (O_2412,N_15977,N_17285);
nand UO_2413 (O_2413,N_18631,N_19556);
nand UO_2414 (O_2414,N_18364,N_17206);
nor UO_2415 (O_2415,N_18161,N_15992);
xor UO_2416 (O_2416,N_15918,N_18489);
and UO_2417 (O_2417,N_19389,N_16307);
nand UO_2418 (O_2418,N_19647,N_19452);
and UO_2419 (O_2419,N_18866,N_16241);
nor UO_2420 (O_2420,N_17925,N_18726);
or UO_2421 (O_2421,N_17605,N_15883);
or UO_2422 (O_2422,N_18691,N_18253);
and UO_2423 (O_2423,N_19277,N_16283);
or UO_2424 (O_2424,N_16096,N_15557);
and UO_2425 (O_2425,N_18667,N_18673);
nor UO_2426 (O_2426,N_17704,N_17079);
or UO_2427 (O_2427,N_17993,N_19987);
nand UO_2428 (O_2428,N_17555,N_19440);
nor UO_2429 (O_2429,N_18603,N_19241);
nor UO_2430 (O_2430,N_17136,N_19824);
or UO_2431 (O_2431,N_15237,N_16403);
or UO_2432 (O_2432,N_15564,N_19172);
or UO_2433 (O_2433,N_18648,N_18300);
and UO_2434 (O_2434,N_17005,N_19984);
nor UO_2435 (O_2435,N_17552,N_19851);
nand UO_2436 (O_2436,N_15111,N_18774);
and UO_2437 (O_2437,N_19007,N_15240);
or UO_2438 (O_2438,N_18935,N_19020);
and UO_2439 (O_2439,N_19691,N_17786);
nand UO_2440 (O_2440,N_15205,N_18433);
and UO_2441 (O_2441,N_18881,N_17997);
nor UO_2442 (O_2442,N_18033,N_19621);
nand UO_2443 (O_2443,N_19121,N_16318);
and UO_2444 (O_2444,N_15881,N_19554);
nor UO_2445 (O_2445,N_15459,N_15818);
or UO_2446 (O_2446,N_17385,N_19534);
xor UO_2447 (O_2447,N_16160,N_18159);
and UO_2448 (O_2448,N_16699,N_16647);
or UO_2449 (O_2449,N_15400,N_17428);
and UO_2450 (O_2450,N_18209,N_17623);
or UO_2451 (O_2451,N_17304,N_19468);
nor UO_2452 (O_2452,N_15347,N_16115);
nand UO_2453 (O_2453,N_19573,N_19560);
xnor UO_2454 (O_2454,N_15106,N_18063);
nor UO_2455 (O_2455,N_18447,N_16407);
and UO_2456 (O_2456,N_15947,N_15982);
or UO_2457 (O_2457,N_19642,N_17501);
nor UO_2458 (O_2458,N_16424,N_16853);
and UO_2459 (O_2459,N_15256,N_17088);
or UO_2460 (O_2460,N_15241,N_19514);
nand UO_2461 (O_2461,N_19073,N_15573);
nand UO_2462 (O_2462,N_17747,N_16344);
nor UO_2463 (O_2463,N_16844,N_16386);
and UO_2464 (O_2464,N_17487,N_16857);
nor UO_2465 (O_2465,N_16226,N_17885);
and UO_2466 (O_2466,N_18668,N_17354);
and UO_2467 (O_2467,N_16133,N_16597);
and UO_2468 (O_2468,N_17012,N_15356);
nor UO_2469 (O_2469,N_18571,N_16204);
nor UO_2470 (O_2470,N_19678,N_19124);
nor UO_2471 (O_2471,N_19071,N_17843);
nor UO_2472 (O_2472,N_19093,N_18980);
nor UO_2473 (O_2473,N_16956,N_19756);
nor UO_2474 (O_2474,N_15168,N_15860);
and UO_2475 (O_2475,N_19435,N_16726);
nand UO_2476 (O_2476,N_18310,N_16632);
and UO_2477 (O_2477,N_18319,N_15794);
and UO_2478 (O_2478,N_19392,N_15108);
or UO_2479 (O_2479,N_15781,N_17435);
and UO_2480 (O_2480,N_19961,N_15697);
nor UO_2481 (O_2481,N_16462,N_19876);
nor UO_2482 (O_2482,N_19760,N_18018);
nor UO_2483 (O_2483,N_16187,N_15001);
and UO_2484 (O_2484,N_15798,N_15277);
and UO_2485 (O_2485,N_17461,N_15448);
nor UO_2486 (O_2486,N_18498,N_16754);
nand UO_2487 (O_2487,N_15435,N_15905);
nand UO_2488 (O_2488,N_16052,N_17966);
or UO_2489 (O_2489,N_17750,N_19053);
and UO_2490 (O_2490,N_15925,N_17258);
nor UO_2491 (O_2491,N_16977,N_16557);
and UO_2492 (O_2492,N_16805,N_16629);
and UO_2493 (O_2493,N_18934,N_17576);
and UO_2494 (O_2494,N_19857,N_19361);
nand UO_2495 (O_2495,N_15974,N_19092);
nor UO_2496 (O_2496,N_15037,N_17541);
or UO_2497 (O_2497,N_18398,N_18022);
and UO_2498 (O_2498,N_18422,N_16174);
or UO_2499 (O_2499,N_18837,N_19326);
endmodule