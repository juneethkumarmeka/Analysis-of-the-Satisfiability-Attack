module basic_2000_20000_2500_5_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_383,In_129);
nor U1 (N_1,In_1839,In_1731);
and U2 (N_2,In_1151,In_1272);
xor U3 (N_3,In_1665,In_1998);
nor U4 (N_4,In_970,In_1369);
and U5 (N_5,In_1754,In_286);
nor U6 (N_6,In_1389,In_713);
nor U7 (N_7,In_1489,In_333);
and U8 (N_8,In_620,In_1917);
nor U9 (N_9,In_1908,In_1596);
xnor U10 (N_10,In_362,In_1959);
or U11 (N_11,In_322,In_56);
or U12 (N_12,In_1221,In_1643);
nand U13 (N_13,In_1978,In_1104);
nor U14 (N_14,In_1184,In_196);
nand U15 (N_15,In_572,In_267);
and U16 (N_16,In_1758,In_1520);
nand U17 (N_17,In_25,In_991);
nor U18 (N_18,In_1505,In_1124);
xnor U19 (N_19,In_101,In_1916);
or U20 (N_20,In_59,In_928);
nor U21 (N_21,In_1242,In_776);
and U22 (N_22,In_31,In_901);
and U23 (N_23,In_526,In_847);
nand U24 (N_24,In_1987,In_1085);
nor U25 (N_25,In_1941,In_468);
xor U26 (N_26,In_1663,In_752);
and U27 (N_27,In_1670,In_161);
and U28 (N_28,In_1289,In_1140);
or U29 (N_29,In_792,In_1641);
xor U30 (N_30,In_12,In_95);
or U31 (N_31,In_354,In_222);
and U32 (N_32,In_555,In_865);
nor U33 (N_33,In_771,In_108);
nor U34 (N_34,In_1247,In_1580);
or U35 (N_35,In_379,In_520);
and U36 (N_36,In_1239,In_1254);
xor U37 (N_37,In_884,In_820);
and U38 (N_38,In_937,In_149);
nor U39 (N_39,In_1760,In_471);
xnor U40 (N_40,In_413,In_660);
nand U41 (N_41,In_1411,In_621);
and U42 (N_42,In_1900,In_260);
nor U43 (N_43,In_1069,In_1743);
xor U44 (N_44,In_1874,In_1409);
nor U45 (N_45,In_715,In_378);
nand U46 (N_46,In_1963,In_995);
nand U47 (N_47,In_919,In_144);
or U48 (N_48,In_274,In_93);
and U49 (N_49,In_1677,In_978);
nand U50 (N_50,In_627,In_192);
nand U51 (N_51,In_1716,In_1092);
nor U52 (N_52,In_1983,In_864);
xor U53 (N_53,In_1189,In_1444);
and U54 (N_54,In_32,In_1410);
and U55 (N_55,In_183,In_603);
and U56 (N_56,In_525,In_1887);
and U57 (N_57,In_1138,In_916);
and U58 (N_58,In_1326,In_1644);
nand U59 (N_59,In_1044,In_1307);
xor U60 (N_60,In_833,In_1684);
nand U61 (N_61,In_134,In_1014);
or U62 (N_62,In_1428,In_723);
and U63 (N_63,In_102,In_1989);
and U64 (N_64,In_508,In_567);
and U65 (N_65,In_597,In_1858);
or U66 (N_66,In_1047,In_1820);
and U67 (N_67,In_1485,In_881);
nand U68 (N_68,In_546,In_45);
nand U69 (N_69,In_1176,In_373);
or U70 (N_70,In_721,In_871);
and U71 (N_71,In_1400,In_287);
nand U72 (N_72,In_807,In_163);
nand U73 (N_73,In_513,In_242);
or U74 (N_74,In_1359,In_122);
nor U75 (N_75,In_1056,In_1732);
and U76 (N_76,In_1283,In_50);
xnor U77 (N_77,In_1600,In_1609);
nor U78 (N_78,In_1769,In_1315);
or U79 (N_79,In_812,In_1507);
nor U80 (N_80,In_414,In_1220);
nor U81 (N_81,In_841,In_1374);
nor U82 (N_82,In_29,In_213);
nand U83 (N_83,In_1686,In_1840);
and U84 (N_84,In_206,In_593);
and U85 (N_85,In_832,In_1667);
and U86 (N_86,In_74,In_1346);
nand U87 (N_87,In_113,In_1035);
or U88 (N_88,In_1564,In_1844);
nor U89 (N_89,In_810,In_693);
or U90 (N_90,In_550,In_214);
nor U91 (N_91,In_1961,In_1569);
nand U92 (N_92,In_39,In_175);
nand U93 (N_93,In_846,In_1304);
and U94 (N_94,In_498,In_439);
and U95 (N_95,In_70,In_283);
and U96 (N_96,In_840,In_1251);
or U97 (N_97,In_1404,In_856);
nand U98 (N_98,In_690,In_749);
and U99 (N_99,In_1435,In_1477);
or U100 (N_100,In_275,In_862);
nand U101 (N_101,In_756,In_446);
or U102 (N_102,In_1182,In_1061);
nand U103 (N_103,In_1353,In_1636);
or U104 (N_104,In_1943,In_731);
xnor U105 (N_105,In_651,In_1067);
nor U106 (N_106,In_172,In_412);
and U107 (N_107,In_582,In_328);
or U108 (N_108,In_392,In_1432);
and U109 (N_109,In_1300,In_123);
xor U110 (N_110,In_658,In_868);
nand U111 (N_111,In_1867,In_366);
nor U112 (N_112,In_141,In_878);
nand U113 (N_113,In_1417,In_1468);
or U114 (N_114,In_1088,In_1697);
and U115 (N_115,In_139,In_1985);
nor U116 (N_116,In_5,In_542);
and U117 (N_117,In_1537,In_1872);
nor U118 (N_118,In_1386,In_1962);
nor U119 (N_119,In_674,In_1431);
nor U120 (N_120,In_630,In_635);
and U121 (N_121,In_823,In_1334);
nand U122 (N_122,In_1121,In_1788);
nor U123 (N_123,In_592,In_1871);
or U124 (N_124,In_1311,In_836);
xor U125 (N_125,In_1995,In_1271);
or U126 (N_126,In_1367,In_228);
nor U127 (N_127,In_949,In_1804);
nand U128 (N_128,In_1826,In_1179);
xnor U129 (N_129,In_1079,In_1378);
nand U130 (N_130,In_939,In_685);
nand U131 (N_131,In_1063,In_1745);
and U132 (N_132,In_1647,In_1341);
nor U133 (N_133,In_1183,In_882);
and U134 (N_134,In_631,In_510);
or U135 (N_135,In_1778,In_57);
xnor U136 (N_136,In_1125,In_1098);
nand U137 (N_137,In_1497,In_107);
nand U138 (N_138,In_662,In_1650);
and U139 (N_139,In_464,In_1122);
nand U140 (N_140,In_1504,In_505);
and U141 (N_141,In_376,In_473);
and U142 (N_142,In_162,In_855);
and U143 (N_143,In_1610,In_1907);
or U144 (N_144,In_1118,In_585);
nand U145 (N_145,In_1591,In_1691);
xor U146 (N_146,In_115,In_705);
nand U147 (N_147,In_1335,In_1688);
nor U148 (N_148,In_1449,In_1893);
or U149 (N_149,In_607,In_1819);
nor U150 (N_150,In_1398,In_1479);
and U151 (N_151,In_231,In_825);
and U152 (N_152,In_536,In_358);
nor U153 (N_153,In_1055,In_600);
xor U154 (N_154,In_1534,In_169);
xnor U155 (N_155,In_350,In_1704);
and U156 (N_156,In_1744,In_641);
or U157 (N_157,In_1236,In_187);
or U158 (N_158,In_1679,In_1040);
and U159 (N_159,In_73,In_639);
or U160 (N_160,In_1921,In_707);
and U161 (N_161,In_1034,In_415);
or U162 (N_162,In_1484,In_1838);
and U163 (N_163,In_1136,In_979);
xnor U164 (N_164,In_1896,In_352);
or U165 (N_165,In_1719,In_209);
or U166 (N_166,In_992,In_461);
nor U167 (N_167,In_33,In_459);
nor U168 (N_168,In_360,In_1499);
nand U169 (N_169,In_1037,In_179);
nand U170 (N_170,In_7,In_1408);
or U171 (N_171,In_176,In_409);
nand U172 (N_172,In_1224,In_581);
nand U173 (N_173,In_529,In_433);
or U174 (N_174,In_1891,In_1022);
xnor U175 (N_175,In_1482,In_858);
or U176 (N_176,In_706,In_809);
or U177 (N_177,In_469,In_610);
and U178 (N_178,In_1146,In_1747);
nand U179 (N_179,In_457,In_1116);
nor U180 (N_180,In_906,In_338);
and U181 (N_181,In_1646,In_1909);
or U182 (N_182,In_61,In_1781);
nand U183 (N_183,In_734,In_1493);
or U184 (N_184,In_454,In_128);
or U185 (N_185,In_241,In_445);
or U186 (N_186,In_1013,In_349);
nor U187 (N_187,In_393,In_925);
and U188 (N_188,In_1205,In_769);
nand U189 (N_189,In_1093,In_186);
nand U190 (N_190,In_1991,In_540);
xor U191 (N_191,In_324,In_745);
nand U192 (N_192,In_357,In_1293);
and U193 (N_193,In_710,In_1199);
nand U194 (N_194,In_897,In_915);
nor U195 (N_195,In_975,In_152);
nand U196 (N_196,In_1828,In_1049);
xnor U197 (N_197,In_1020,In_1120);
or U198 (N_198,In_1860,In_815);
nor U199 (N_199,In_813,In_1005);
nor U200 (N_200,In_1194,In_1469);
and U201 (N_201,In_740,In_427);
and U202 (N_202,In_528,In_1883);
and U203 (N_203,In_1773,In_1946);
and U204 (N_204,In_1405,In_575);
or U205 (N_205,In_938,In_1654);
xor U206 (N_206,In_14,In_558);
nor U207 (N_207,In_1944,In_1217);
or U208 (N_208,In_1514,In_625);
xor U209 (N_209,In_1529,In_647);
and U210 (N_210,In_435,In_1280);
and U211 (N_211,In_561,In_1656);
and U212 (N_212,In_480,In_1738);
and U213 (N_213,In_310,In_748);
xor U214 (N_214,In_950,In_185);
and U215 (N_215,In_1866,In_1388);
nor U216 (N_216,In_634,In_1969);
and U217 (N_217,In_83,In_1624);
nor U218 (N_218,In_1458,In_1281);
or U219 (N_219,In_564,In_46);
and U220 (N_220,In_402,In_1175);
nand U221 (N_221,In_1561,In_1267);
or U222 (N_222,In_1793,In_391);
or U223 (N_223,In_262,In_910);
xnor U224 (N_224,In_1051,In_1734);
xor U225 (N_225,In_1545,In_1824);
nand U226 (N_226,In_772,In_606);
nor U227 (N_227,In_791,In_1581);
nand U228 (N_228,In_802,In_1859);
nor U229 (N_229,In_808,In_1814);
nor U230 (N_230,In_1786,In_1972);
nor U231 (N_231,In_1160,In_84);
nand U232 (N_232,In_1099,In_372);
and U233 (N_233,In_726,In_1421);
nand U234 (N_234,In_720,In_37);
or U235 (N_235,In_211,In_1533);
nand U236 (N_236,In_1238,In_766);
or U237 (N_237,In_1815,In_13);
and U238 (N_238,In_676,In_1546);
nand U239 (N_239,In_237,In_504);
nand U240 (N_240,In_418,In_1555);
and U241 (N_241,In_460,In_28);
and U242 (N_242,In_238,In_335);
or U243 (N_243,In_254,In_250);
and U244 (N_244,In_859,In_1938);
or U245 (N_245,In_556,In_885);
nor U246 (N_246,In_1174,In_1787);
nor U247 (N_247,In_1064,In_1023);
nand U248 (N_248,In_1225,In_448);
xnor U249 (N_249,In_340,In_1631);
xnor U250 (N_250,In_1953,In_518);
xor U251 (N_251,In_1358,In_235);
and U252 (N_252,In_1578,In_1523);
nor U253 (N_253,In_424,In_797);
nand U254 (N_254,In_680,In_1592);
and U255 (N_255,In_1095,In_611);
nor U256 (N_256,In_120,In_282);
nor U257 (N_257,In_400,In_1375);
or U258 (N_258,In_1920,In_1904);
xnor U259 (N_259,In_1930,In_534);
and U260 (N_260,In_533,In_71);
nand U261 (N_261,In_1133,In_1735);
nor U262 (N_262,In_401,In_436);
and U263 (N_263,In_531,In_778);
nor U264 (N_264,In_1748,In_1019);
or U265 (N_265,In_1892,In_1733);
or U266 (N_266,In_1567,In_997);
xnor U267 (N_267,In_232,In_1384);
and U268 (N_268,In_784,In_1572);
nor U269 (N_269,In_1889,In_612);
or U270 (N_270,In_568,In_694);
nand U271 (N_271,In_1925,In_1750);
nand U272 (N_272,In_1777,In_466);
nand U273 (N_273,In_828,In_353);
and U274 (N_274,In_423,In_375);
nor U275 (N_275,In_87,In_1390);
nor U276 (N_276,In_741,In_1041);
or U277 (N_277,In_487,In_921);
nor U278 (N_278,In_1956,In_1807);
and U279 (N_279,In_1509,In_408);
nand U280 (N_280,In_1577,In_381);
xor U281 (N_281,In_1779,In_574);
nor U282 (N_282,In_276,In_1864);
or U283 (N_283,In_596,In_775);
and U284 (N_284,In_1594,In_1086);
and U285 (N_285,In_180,In_1492);
nand U286 (N_286,In_1424,In_1651);
xnor U287 (N_287,In_347,In_1336);
nor U288 (N_288,In_1999,In_1616);
nand U289 (N_289,In_946,In_936);
and U290 (N_290,In_472,In_1898);
and U291 (N_291,In_1439,In_1597);
nand U292 (N_292,In_1462,In_119);
and U293 (N_293,In_655,In_875);
nand U294 (N_294,In_1377,In_1002);
nand U295 (N_295,In_764,In_1323);
or U296 (N_296,In_21,In_1396);
nand U297 (N_297,In_800,In_1290);
or U298 (N_298,In_1268,In_768);
nor U299 (N_299,In_1234,In_233);
and U300 (N_300,In_58,In_1699);
or U301 (N_301,In_30,In_10);
and U302 (N_302,In_1994,In_757);
and U303 (N_303,In_1081,In_532);
and U304 (N_304,In_1027,In_168);
and U305 (N_305,In_500,In_1463);
and U306 (N_306,In_1689,In_1541);
or U307 (N_307,In_1822,In_1169);
and U308 (N_308,In_1071,In_1172);
xor U309 (N_309,In_202,In_1123);
and U310 (N_310,In_1440,In_1046);
and U311 (N_311,In_331,In_566);
and U312 (N_312,In_626,In_1940);
or U313 (N_313,In_314,In_1834);
or U314 (N_314,In_1980,In_1601);
or U315 (N_315,In_1903,In_1693);
and U316 (N_316,In_40,In_1584);
nor U317 (N_317,In_109,In_577);
nor U318 (N_318,In_1633,In_1583);
and U319 (N_319,In_1001,In_1302);
or U320 (N_320,In_763,In_1059);
nor U321 (N_321,In_1416,In_245);
or U322 (N_322,In_1134,In_96);
nand U323 (N_323,In_1441,In_1589);
xor U324 (N_324,In_893,In_648);
nand U325 (N_325,In_1451,In_319);
nor U326 (N_326,In_1399,In_348);
xor U327 (N_327,In_22,In_1329);
xor U328 (N_328,In_765,In_675);
and U329 (N_329,In_266,In_259);
nand U330 (N_330,In_1923,In_1842);
nor U331 (N_331,In_587,In_482);
nor U332 (N_332,In_200,In_1318);
nand U333 (N_333,In_735,In_996);
nand U334 (N_334,In_1167,In_867);
or U335 (N_335,In_382,In_1881);
or U336 (N_336,In_1918,In_1762);
or U337 (N_337,In_441,In_1582);
and U338 (N_338,In_956,In_537);
nor U339 (N_339,In_1127,In_1250);
xnor U340 (N_340,In_204,In_1371);
or U341 (N_341,In_1950,In_304);
nand U342 (N_342,In_1705,In_485);
xor U343 (N_343,In_1683,In_456);
nand U344 (N_344,In_886,In_1515);
nor U345 (N_345,In_229,In_1391);
and U346 (N_346,In_329,In_1948);
xor U347 (N_347,In_1203,In_790);
nand U348 (N_348,In_920,In_663);
xor U349 (N_349,In_609,In_1548);
and U350 (N_350,In_1158,In_133);
nor U351 (N_351,In_1796,In_1422);
nand U352 (N_352,In_594,In_1926);
nor U353 (N_353,In_296,In_940);
or U354 (N_354,In_1540,In_1658);
nand U355 (N_355,In_394,In_1986);
or U356 (N_356,In_747,In_1967);
and U357 (N_357,In_1278,In_221);
nand U358 (N_358,In_1437,In_554);
nor U359 (N_359,In_852,In_223);
and U360 (N_360,In_984,In_805);
nor U361 (N_361,In_293,In_279);
and U362 (N_362,In_150,In_1736);
and U363 (N_363,In_285,In_780);
or U364 (N_364,In_417,In_1206);
and U365 (N_365,In_346,In_1749);
and U366 (N_366,In_614,In_1246);
or U367 (N_367,In_494,In_686);
and U368 (N_368,In_742,In_1464);
or U369 (N_369,In_1869,In_272);
or U370 (N_370,In_1818,In_1782);
and U371 (N_371,In_1894,In_1718);
nand U372 (N_372,In_794,In_151);
nor U373 (N_373,In_584,In_746);
nor U374 (N_374,In_848,In_1078);
nand U375 (N_375,In_1722,In_1080);
and U376 (N_376,In_1165,In_1803);
xnor U377 (N_377,In_1666,In_1007);
xor U378 (N_378,In_361,In_1108);
nor U379 (N_379,In_945,In_704);
and U380 (N_380,In_935,In_1958);
nand U381 (N_381,In_1102,In_1614);
or U382 (N_382,In_499,In_1370);
or U383 (N_383,In_944,In_1201);
or U384 (N_384,In_1681,In_1106);
nand U385 (N_385,In_1368,In_672);
nand U386 (N_386,In_19,In_1695);
or U387 (N_387,In_908,In_1456);
nor U388 (N_388,In_1992,In_1296);
and U389 (N_389,In_1621,In_1087);
and U390 (N_390,In_269,In_579);
nand U391 (N_391,In_873,In_1314);
nand U392 (N_392,In_1342,In_1645);
or U393 (N_393,In_1915,In_243);
nor U394 (N_394,In_263,In_1284);
nand U395 (N_395,In_1954,In_955);
nand U396 (N_396,In_1157,In_1951);
or U397 (N_397,In_1072,In_1611);
nor U398 (N_398,In_729,In_420);
or U399 (N_399,In_1901,In_968);
or U400 (N_400,In_497,In_1783);
and U401 (N_401,In_440,In_326);
nand U402 (N_402,In_278,In_1993);
nand U403 (N_403,In_234,In_543);
xnor U404 (N_404,In_682,In_602);
and U405 (N_405,In_305,In_953);
nand U406 (N_406,In_2,In_431);
or U407 (N_407,In_208,In_861);
nor U408 (N_408,In_1381,In_1937);
nand U409 (N_409,In_289,In_355);
nor U410 (N_410,In_1853,In_957);
nor U411 (N_411,In_1117,In_1149);
or U412 (N_412,In_1259,In_1598);
nor U413 (N_413,In_1303,In_60);
nor U414 (N_414,In_1687,In_1847);
nand U415 (N_415,In_86,In_986);
nor U416 (N_416,In_1521,In_1316);
and U417 (N_417,In_604,In_1139);
nand U418 (N_418,In_1263,In_728);
nor U419 (N_419,In_1130,In_244);
xor U420 (N_420,In_973,In_1276);
and U421 (N_421,In_1530,In_1532);
nand U422 (N_422,In_1202,In_1401);
and U423 (N_423,In_68,In_316);
nor U424 (N_424,In_538,In_1821);
nor U425 (N_425,In_1083,In_1208);
and U426 (N_426,In_830,In_1806);
nor U427 (N_427,In_288,In_1319);
or U428 (N_428,In_1476,In_1365);
and U429 (N_429,In_201,In_1207);
and U430 (N_430,In_255,In_509);
nand U431 (N_431,In_1528,In_1245);
nor U432 (N_432,In_1438,In_398);
or U433 (N_433,In_1279,In_1036);
nor U434 (N_434,In_618,In_1606);
or U435 (N_435,In_81,In_755);
or U436 (N_436,In_773,In_356);
nor U437 (N_437,In_1376,In_1003);
or U438 (N_438,In_1882,In_530);
or U439 (N_439,In_1837,In_1198);
nor U440 (N_440,In_822,In_1710);
and U441 (N_441,In_1294,In_934);
nand U442 (N_442,In_142,In_1630);
and U443 (N_443,In_657,In_583);
nand U444 (N_444,In_1608,In_754);
nor U445 (N_445,In_777,In_739);
and U446 (N_446,In_1004,In_1549);
or U447 (N_447,In_1934,In_295);
or U448 (N_448,In_1164,In_1380);
xor U449 (N_449,In_1426,In_1527);
nand U450 (N_450,In_8,In_1131);
and U451 (N_451,In_1642,In_1494);
nor U452 (N_452,In_1590,In_688);
and U453 (N_453,In_3,In_1029);
xor U454 (N_454,In_1491,In_1805);
xnor U455 (N_455,In_1563,In_230);
or U456 (N_456,In_110,In_1811);
nor U457 (N_457,In_131,In_1947);
nand U458 (N_458,In_143,In_66);
nor U459 (N_459,In_835,In_1927);
or U460 (N_460,In_363,In_699);
and U461 (N_461,In_601,In_1);
or U462 (N_462,In_369,In_264);
and U463 (N_463,In_1902,In_1397);
and U464 (N_464,In_770,In_1077);
or U465 (N_465,In_909,In_608);
nor U466 (N_466,In_1385,In_34);
xnor U467 (N_467,In_51,In_1387);
nand U468 (N_468,In_1849,In_1459);
xnor U469 (N_469,In_406,In_629);
and U470 (N_470,In_1073,In_277);
xor U471 (N_471,In_1039,In_899);
or U472 (N_472,In_1571,In_1727);
nor U473 (N_473,In_374,In_912);
xor U474 (N_474,In_1884,In_1185);
and U475 (N_475,In_312,In_1282);
nand U476 (N_476,In_732,In_981);
and U477 (N_477,In_481,In_1560);
nor U478 (N_478,In_387,In_1012);
nand U479 (N_479,In_419,In_48);
nand U480 (N_480,In_551,In_1057);
and U481 (N_481,In_1126,In_160);
or U482 (N_482,In_922,In_857);
and U483 (N_483,In_78,In_303);
or U484 (N_484,In_1091,In_1706);
or U485 (N_485,In_980,In_616);
and U486 (N_486,In_1850,In_552);
and U487 (N_487,In_100,In_1797);
and U488 (N_488,In_1255,In_880);
nor U489 (N_489,In_599,In_814);
and U490 (N_490,In_1775,In_1700);
and U491 (N_491,In_280,In_1949);
xor U492 (N_492,In_877,In_1595);
nor U493 (N_493,In_67,In_1017);
nor U494 (N_494,In_309,In_1446);
nand U495 (N_495,In_565,In_1309);
nand U496 (N_496,In_1639,In_727);
nor U497 (N_497,In_191,In_451);
nand U498 (N_498,In_1053,In_1729);
nand U499 (N_499,In_190,In_1361);
or U500 (N_500,In_570,In_1256);
or U501 (N_501,In_1000,In_640);
and U502 (N_502,In_193,In_170);
and U503 (N_503,In_1042,In_994);
or U504 (N_504,In_54,In_644);
nor U505 (N_505,In_1535,In_1328);
nor U506 (N_506,In_1321,In_1511);
nor U507 (N_507,In_1038,In_308);
nor U508 (N_508,In_1680,In_1790);
nor U509 (N_509,In_1539,In_943);
nor U510 (N_510,In_426,In_1765);
and U511 (N_511,In_1725,In_913);
and U512 (N_512,In_911,In_1177);
nand U513 (N_513,In_789,In_490);
or U514 (N_514,In_1905,In_932);
or U515 (N_515,In_425,In_15);
xnor U516 (N_516,In_364,In_1197);
nor U517 (N_517,In_1586,In_831);
nand U518 (N_518,In_1966,In_866);
nand U519 (N_519,In_502,In_719);
xnor U520 (N_520,In_1526,In_1460);
nor U521 (N_521,In_586,In_388);
nor U522 (N_522,In_1043,In_698);
or U523 (N_523,In_9,In_1518);
and U524 (N_524,In_578,In_1660);
nor U525 (N_525,In_559,In_197);
xnor U526 (N_526,In_428,In_1784);
and U527 (N_527,In_1195,In_1668);
or U528 (N_528,In_483,In_1156);
and U529 (N_529,In_470,In_365);
or U530 (N_530,In_442,In_1178);
nand U531 (N_531,In_1513,In_47);
nand U532 (N_532,In_1114,In_1573);
or U533 (N_533,In_1524,In_1723);
xnor U534 (N_534,In_1266,In_294);
nor U535 (N_535,In_103,In_619);
nor U536 (N_536,In_1914,In_359);
and U537 (N_537,In_702,In_1971);
nor U538 (N_538,In_1009,In_1632);
nand U539 (N_539,In_1481,In_1615);
and U540 (N_540,In_1717,In_1345);
or U541 (N_541,In_1575,In_926);
nand U542 (N_542,In_1299,In_1058);
nor U543 (N_543,In_665,In_105);
and U544 (N_544,In_463,In_1759);
or U545 (N_545,In_1770,In_1478);
nor U546 (N_546,In_495,In_501);
or U547 (N_547,In_914,In_691);
or U548 (N_548,In_1721,In_1933);
nand U549 (N_549,In_281,In_1928);
or U550 (N_550,In_638,In_1188);
and U551 (N_551,In_215,In_1868);
or U552 (N_552,In_684,In_972);
nand U553 (N_553,In_1510,In_1857);
or U554 (N_554,In_225,In_605);
nor U555 (N_555,In_218,In_1506);
or U556 (N_556,In_1619,In_1154);
nor U557 (N_557,In_1144,In_895);
xor U558 (N_558,In_1100,In_1746);
nand U559 (N_559,In_1472,In_633);
or U560 (N_560,In_1599,In_759);
or U561 (N_561,In_82,In_709);
nand U562 (N_562,In_904,In_226);
and U563 (N_563,In_23,In_1219);
and U564 (N_564,In_258,In_474);
or U565 (N_565,In_1984,In_315);
or U566 (N_566,In_156,In_1655);
xor U567 (N_567,In_761,In_158);
nor U568 (N_568,In_205,In_1741);
or U569 (N_569,In_1427,In_1696);
or U570 (N_570,In_1181,In_210);
nor U571 (N_571,In_249,In_1906);
and U572 (N_572,In_1135,In_1843);
nor U573 (N_573,In_679,In_342);
and U574 (N_574,In_503,In_1848);
and U575 (N_575,In_1957,In_1110);
and U576 (N_576,In_1516,In_576);
and U577 (N_577,In_1554,In_1800);
nand U578 (N_578,In_827,In_1789);
or U579 (N_579,In_1895,In_1570);
nor U580 (N_580,In_290,In_1671);
xor U581 (N_581,In_1310,In_1470);
xor U582 (N_582,In_140,In_1467);
nor U583 (N_583,In_562,In_869);
nor U584 (N_584,In_696,In_1339);
and U585 (N_585,In_1090,In_514);
nand U586 (N_586,In_670,In_1536);
nand U587 (N_587,In_1720,In_1952);
nor U588 (N_588,In_1669,In_795);
nand U589 (N_589,In_1712,In_507);
nand U590 (N_590,In_1538,In_1354);
nor U591 (N_591,In_465,In_1752);
or U592 (N_592,In_816,In_135);
nand U593 (N_593,In_839,In_782);
nand U594 (N_594,In_1638,In_438);
nor U595 (N_595,In_1286,In_443);
and U596 (N_596,In_164,In_743);
or U597 (N_597,In_1593,In_569);
nand U598 (N_598,In_1825,In_256);
xor U599 (N_599,In_1751,In_964);
xor U600 (N_600,In_1209,In_1543);
or U601 (N_601,In_1052,In_522);
or U602 (N_602,In_1841,In_385);
nor U603 (N_603,In_1931,In_1618);
nor U604 (N_604,In_1585,In_1682);
nand U605 (N_605,In_1480,In_1343);
and U606 (N_606,In_104,In_1233);
nand U607 (N_607,In_1362,In_982);
nor U608 (N_608,In_1423,In_1089);
nor U609 (N_609,In_1153,In_421);
and U610 (N_610,In_1333,In_320);
and U611 (N_611,In_146,In_43);
and U612 (N_612,In_512,In_1877);
or U613 (N_613,In_1794,In_1148);
and U614 (N_614,In_1355,In_622);
and U615 (N_615,In_1244,In_1776);
nand U616 (N_616,In_1832,In_774);
nor U617 (N_617,In_20,In_853);
nand U618 (N_618,In_1379,In_1287);
nor U619 (N_619,In_475,In_623);
nor U620 (N_620,In_637,In_1964);
or U621 (N_621,In_1429,In_1503);
xnor U622 (N_622,In_1436,In_1274);
nor U623 (N_623,In_184,In_1792);
or U624 (N_624,In_1313,In_106);
xnor U625 (N_625,In_1060,In_1347);
nand U626 (N_626,In_377,In_1604);
xnor U627 (N_627,In_153,In_1292);
or U628 (N_628,In_1870,In_299);
nand U629 (N_629,In_1094,In_1269);
nand U630 (N_630,In_1701,In_1248);
or U631 (N_631,In_1325,In_1612);
or U632 (N_632,In_318,In_1757);
nand U633 (N_633,In_1862,In_24);
nand U634 (N_634,In_1406,In_1229);
and U635 (N_635,In_88,In_874);
and U636 (N_636,In_493,In_174);
and U637 (N_637,In_1622,In_1414);
nand U638 (N_638,In_1587,In_793);
nand U639 (N_639,In_1495,In_1831);
nor U640 (N_640,In_252,In_188);
nand U641 (N_641,In_588,In_1913);
or U642 (N_642,In_313,In_1352);
xnor U643 (N_643,In_1211,In_343);
and U644 (N_644,In_931,In_548);
and U645 (N_645,In_1363,In_798);
nor U646 (N_646,In_1960,In_1265);
nand U647 (N_647,In_1674,In_1275);
or U648 (N_648,In_1559,In_1107);
and U649 (N_649,In_330,In_1672);
nand U650 (N_650,In_843,In_941);
or U651 (N_651,In_971,In_1119);
or U652 (N_652,In_796,In_1922);
or U653 (N_653,In_801,In_1137);
or U654 (N_654,In_1486,In_929);
nor U655 (N_655,In_598,In_744);
and U656 (N_656,In_16,In_1068);
xnor U657 (N_657,In_1817,In_1048);
xor U658 (N_658,In_1173,In_165);
or U659 (N_659,In_1419,In_560);
xor U660 (N_660,In_1364,In_124);
and U661 (N_661,In_1888,In_220);
or U662 (N_662,In_580,In_850);
and U663 (N_663,In_1338,In_1132);
nand U664 (N_664,In_1452,In_311);
or U665 (N_665,In_1603,In_94);
nand U666 (N_666,In_99,In_195);
nand U667 (N_667,In_725,In_1455);
or U668 (N_668,In_1768,In_687);
or U669 (N_669,In_1711,In_1301);
nor U670 (N_670,In_351,In_656);
xor U671 (N_671,In_1159,In_1565);
nor U672 (N_672,In_63,In_521);
nor U673 (N_673,In_947,In_127);
nor U674 (N_674,In_787,In_137);
nand U675 (N_675,In_649,In_1474);
or U676 (N_676,In_219,In_668);
nand U677 (N_677,In_38,In_1675);
or U678 (N_678,In_1171,In_1795);
xnor U679 (N_679,In_1420,In_97);
or U680 (N_680,In_1740,In_722);
nand U681 (N_681,In_154,In_11);
and U682 (N_682,In_1392,In_967);
or U683 (N_683,In_1298,In_1483);
xnor U684 (N_684,In_1912,In_966);
and U685 (N_685,In_1519,In_1187);
xnor U686 (N_686,In_467,In_760);
and U687 (N_687,In_817,In_1935);
nand U688 (N_688,In_35,In_1501);
nor U689 (N_689,In_1155,In_1443);
nand U690 (N_690,In_1975,In_1115);
nand U691 (N_691,In_1070,In_1273);
nor U692 (N_692,In_1498,In_432);
nor U693 (N_693,In_1635,In_52);
and U694 (N_694,In_751,In_325);
nand U695 (N_695,In_1050,In_811);
or U696 (N_696,In_677,In_399);
or U697 (N_697,In_247,In_1739);
xnor U698 (N_698,In_1327,In_1496);
nand U699 (N_699,In_384,In_628);
nor U700 (N_700,In_1340,In_1076);
or U701 (N_701,In_1393,In_1508);
nor U702 (N_702,In_1241,In_1488);
or U703 (N_703,In_714,In_1500);
and U704 (N_704,In_489,In_1021);
nand U705 (N_705,In_1772,In_1415);
or U706 (N_706,In_666,In_519);
nand U707 (N_707,In_1755,In_1490);
nand U708 (N_708,In_1628,In_332);
nor U709 (N_709,In_1442,In_395);
or U710 (N_710,In_1030,In_166);
nand U711 (N_711,In_799,In_1232);
nor U712 (N_712,In_999,In_1551);
xor U713 (N_713,In_1407,In_511);
or U714 (N_714,In_571,In_990);
nor U715 (N_715,In_1690,In_1223);
and U716 (N_716,In_198,In_321);
or U717 (N_717,In_236,In_624);
and U718 (N_718,In_1833,In_1075);
and U719 (N_719,In_669,In_1257);
and U720 (N_720,In_1285,In_1141);
xnor U721 (N_721,In_1240,In_1676);
or U722 (N_722,In_1808,In_1726);
nor U723 (N_723,In_1899,In_1974);
or U724 (N_724,In_42,In_1640);
and U725 (N_725,In_1066,In_1827);
and U726 (N_726,In_1170,In_683);
nand U727 (N_727,In_49,In_1780);
or U728 (N_728,In_1348,In_1475);
or U729 (N_729,In_785,In_1357);
nand U730 (N_730,In_1096,In_1649);
and U731 (N_731,In_62,In_1627);
or U732 (N_732,In_69,In_1791);
and U733 (N_733,In_491,In_891);
nor U734 (N_734,In_157,In_306);
or U735 (N_735,In_85,In_697);
or U736 (N_736,In_730,In_1813);
and U737 (N_737,In_300,In_407);
or U738 (N_738,In_1713,In_371);
nor U739 (N_739,In_79,In_708);
or U740 (N_740,In_889,In_589);
or U741 (N_741,In_1062,In_207);
nor U742 (N_742,In_1331,In_1262);
or U743 (N_743,In_851,In_112);
or U744 (N_744,In_824,In_1728);
nand U745 (N_745,In_1552,In_1673);
nand U746 (N_746,In_930,In_863);
xor U747 (N_747,In_1213,In_345);
nor U748 (N_748,In_1180,In_1522);
xor U749 (N_749,In_783,In_1981);
nand U750 (N_750,In_1812,In_1502);
and U751 (N_751,In_411,In_1230);
nand U752 (N_752,In_664,In_650);
or U753 (N_753,In_1556,In_339);
and U754 (N_754,In_1161,In_126);
or U755 (N_755,In_883,In_265);
or U756 (N_756,In_902,In_1142);
nand U757 (N_757,In_479,In_1193);
or U758 (N_758,In_1756,In_317);
and U759 (N_759,In_918,In_1434);
nor U760 (N_760,In_1863,In_806);
nor U761 (N_761,In_1929,In_724);
nor U762 (N_762,In_695,In_767);
nor U763 (N_763,In_1662,In_788);
or U764 (N_764,In_422,In_1707);
nor U765 (N_765,In_1648,In_98);
nor U766 (N_766,In_1450,In_527);
or U767 (N_767,In_1143,In_516);
xnor U768 (N_768,In_1761,In_961);
or U769 (N_769,In_1412,In_1113);
nor U770 (N_770,In_1664,In_905);
nand U771 (N_771,In_998,In_298);
or U772 (N_772,In_636,In_344);
xnor U773 (N_773,In_661,In_826);
nor U774 (N_774,In_1657,In_246);
nand U775 (N_775,In_1235,In_733);
nor U776 (N_776,In_1835,In_251);
nor U777 (N_777,In_1190,In_1413);
nor U778 (N_778,In_177,In_301);
nor U779 (N_779,In_1602,In_1865);
nand U780 (N_780,In_1212,In_1637);
nand U781 (N_781,In_1471,In_248);
nor U782 (N_782,In_1919,In_1629);
or U783 (N_783,In_1330,In_1851);
nor U784 (N_784,In_1942,In_1332);
and U785 (N_785,In_449,In_1227);
nor U786 (N_786,In_692,In_1228);
nor U787 (N_787,In_1258,In_405);
nand U788 (N_788,In_646,In_1032);
nor U789 (N_789,In_1454,In_1517);
and U790 (N_790,In_136,In_1461);
and U791 (N_791,In_462,In_894);
nor U792 (N_792,In_892,In_1109);
nor U793 (N_793,In_1425,In_4);
nand U794 (N_794,In_643,In_1018);
xor U795 (N_795,In_64,In_1531);
and U796 (N_796,In_1990,In_1324);
nor U797 (N_797,In_804,In_273);
xnor U798 (N_798,In_645,In_557);
or U799 (N_799,In_1105,In_307);
or U800 (N_800,In_954,In_368);
nand U801 (N_801,In_1836,In_1885);
or U802 (N_802,In_523,In_870);
or U803 (N_803,In_17,In_397);
or U804 (N_804,In_1011,In_1082);
nor U805 (N_805,In_132,In_854);
nor U806 (N_806,In_927,In_948);
and U807 (N_807,In_1191,In_515);
or U808 (N_808,In_678,In_700);
nand U809 (N_809,In_386,In_270);
xor U810 (N_810,In_1016,In_654);
xnor U811 (N_811,In_239,In_736);
xor U812 (N_812,In_976,In_1976);
nand U813 (N_813,In_1226,In_1337);
xor U814 (N_814,In_1447,In_452);
nor U815 (N_815,In_212,In_1360);
nand U816 (N_816,In_334,In_189);
and U817 (N_817,In_416,In_1566);
and U818 (N_818,In_1764,In_1855);
nand U819 (N_819,In_1996,In_1945);
and U820 (N_820,In_27,In_1801);
nand U821 (N_821,In_541,In_1270);
nor U822 (N_822,In_1261,In_1568);
and U823 (N_823,In_1715,In_1897);
or U824 (N_824,In_1730,In_257);
xor U825 (N_825,In_92,In_1351);
nand U826 (N_826,In_1965,In_447);
nand U827 (N_827,In_147,In_1968);
or U828 (N_828,In_341,In_77);
and U829 (N_829,In_1607,In_336);
nor U830 (N_830,In_1767,In_1771);
and U831 (N_831,In_1753,In_117);
and U832 (N_832,In_1653,In_450);
and U833 (N_833,In_1054,In_842);
and U834 (N_834,In_1145,In_549);
nand U835 (N_835,In_1074,In_974);
and U836 (N_836,In_1028,In_834);
or U837 (N_837,In_1886,In_182);
nand U838 (N_838,In_1977,In_1605);
and U839 (N_839,In_1714,In_1830);
nand U840 (N_840,In_837,In_1097);
nand U841 (N_841,In_26,In_458);
or U842 (N_842,In_130,In_1625);
and U843 (N_843,In_539,In_1403);
nor U844 (N_844,In_36,In_903);
xor U845 (N_845,In_717,In_1879);
or U846 (N_846,In_1823,In_1204);
or U847 (N_847,In_1579,In_1634);
and U848 (N_848,In_1260,In_167);
or U849 (N_849,In_1306,In_1192);
or U850 (N_850,In_476,In_1588);
nor U851 (N_851,In_1737,In_434);
nor U852 (N_852,In_1875,In_145);
nor U853 (N_853,In_977,In_1147);
or U854 (N_854,In_819,In_829);
and U855 (N_855,In_969,In_983);
nand U856 (N_856,In_53,In_962);
and U857 (N_857,In_1349,In_844);
xnor U858 (N_858,In_1445,In_1200);
and U859 (N_859,In_114,In_1101);
nor U860 (N_860,In_988,In_1453);
and U861 (N_861,In_323,In_1312);
nand U862 (N_862,In_1305,In_18);
and U863 (N_863,In_0,In_613);
and U864 (N_864,In_958,In_737);
nand U865 (N_865,In_1932,In_224);
nand U866 (N_866,In_1084,In_535);
nand U867 (N_867,In_1816,In_1574);
nor U868 (N_868,In_876,In_1163);
nand U869 (N_869,In_410,In_292);
nand U870 (N_870,In_1350,In_1617);
or U871 (N_871,In_750,In_1295);
or U872 (N_872,In_758,In_1372);
or U873 (N_873,In_171,In_595);
and U874 (N_874,In_1982,In_671);
and U875 (N_875,In_72,In_1356);
and U876 (N_876,In_1243,In_1512);
or U877 (N_877,In_1678,In_1025);
or U878 (N_878,In_987,In_1473);
nand U879 (N_879,In_1542,In_1979);
nand U880 (N_880,In_1988,In_1308);
or U881 (N_881,In_1252,In_963);
xnor U882 (N_882,In_1487,In_632);
xor U883 (N_883,In_65,In_148);
or U884 (N_884,In_779,In_1277);
nor U885 (N_885,In_1210,In_1196);
nand U886 (N_886,In_1166,In_547);
or U887 (N_887,In_1854,In_437);
nand U888 (N_888,In_1576,In_1186);
or U889 (N_889,In_1856,In_701);
nor U890 (N_890,In_1264,In_1150);
and U891 (N_891,In_240,In_1924);
xor U892 (N_892,In_659,In_1112);
nand U893 (N_893,In_993,In_478);
xor U894 (N_894,In_1031,In_1724);
nand U895 (N_895,In_261,In_116);
nand U896 (N_896,In_1320,In_1997);
nand U897 (N_897,In_370,In_492);
nor U898 (N_898,In_216,In_496);
nor U899 (N_899,In_1809,In_390);
nor U900 (N_900,In_367,In_951);
nand U901 (N_901,In_896,In_1128);
and U902 (N_902,In_121,In_203);
nor U903 (N_903,In_900,In_849);
nand U904 (N_904,In_404,In_1317);
nor U905 (N_905,In_753,In_1623);
or U906 (N_906,In_159,In_44);
nand U907 (N_907,In_890,In_1218);
or U908 (N_908,In_681,In_1448);
nand U909 (N_909,In_1620,In_1402);
and U910 (N_910,In_1970,In_1544);
nand U911 (N_911,In_1852,In_1111);
or U912 (N_912,In_689,In_271);
and U913 (N_913,In_573,In_90);
nand U914 (N_914,In_91,In_860);
and U915 (N_915,In_302,In_1010);
nand U916 (N_916,In_703,In_821);
and U917 (N_917,In_389,In_178);
xnor U918 (N_918,In_1558,In_1890);
or U919 (N_919,In_1661,In_1430);
xnor U920 (N_920,In_989,In_1910);
and U921 (N_921,In_194,In_268);
and U922 (N_922,In_1395,In_1152);
and U923 (N_923,In_1562,In_942);
nor U924 (N_924,In_1709,In_1873);
nand U925 (N_925,In_1846,In_253);
nor U926 (N_926,In_1026,In_455);
or U927 (N_927,In_716,In_907);
nor U928 (N_928,In_1288,In_933);
nand U929 (N_929,In_227,In_111);
xnor U930 (N_930,In_396,In_1222);
nand U931 (N_931,In_1344,In_1291);
or U932 (N_932,In_965,In_76);
xor U933 (N_933,In_181,In_1708);
and U934 (N_934,In_818,In_1557);
nand U935 (N_935,In_1006,In_1692);
or U936 (N_936,In_1525,In_1214);
or U937 (N_937,In_1024,In_337);
nor U938 (N_938,In_1394,In_1033);
and U939 (N_939,In_872,In_1015);
nor U940 (N_940,In_1433,In_1955);
xor U941 (N_941,In_1880,In_617);
nand U942 (N_942,In_1703,In_887);
nor U943 (N_943,In_985,In_1694);
and U944 (N_944,In_1457,In_1785);
and U945 (N_945,In_1698,In_898);
xor U946 (N_946,In_1045,In_125);
nand U947 (N_947,In_1936,In_1465);
and U948 (N_948,In_1798,In_55);
nand U949 (N_949,In_653,In_477);
or U950 (N_950,In_6,In_429);
nor U951 (N_951,In_1802,In_1418);
and U952 (N_952,In_590,In_923);
nor U953 (N_953,In_712,In_486);
nor U954 (N_954,In_284,In_217);
and U955 (N_955,In_488,In_1659);
xor U956 (N_956,In_591,In_1065);
and U957 (N_957,In_1774,In_1742);
xnor U958 (N_958,In_845,In_563);
or U959 (N_959,In_718,In_403);
nand U960 (N_960,In_1685,In_960);
nand U961 (N_961,In_1237,In_673);
nand U962 (N_962,In_173,In_1383);
or U963 (N_963,In_1103,In_517);
nand U964 (N_964,In_838,In_1878);
nor U965 (N_965,In_506,In_1626);
or U966 (N_966,In_1911,In_1876);
nand U967 (N_967,In_1553,In_879);
or U968 (N_968,In_959,In_297);
nand U969 (N_969,In_89,In_1322);
nor U970 (N_970,In_1766,In_1253);
nor U971 (N_971,In_327,In_952);
xnor U972 (N_972,In_762,In_1702);
or U973 (N_973,In_80,In_453);
or U974 (N_974,In_118,In_75);
nand U975 (N_975,In_484,In_1249);
or U976 (N_976,In_1168,In_444);
xnor U977 (N_977,In_1845,In_1466);
or U978 (N_978,In_1799,In_1231);
and U979 (N_979,In_1973,In_155);
nor U980 (N_980,In_1861,In_888);
nor U981 (N_981,In_781,In_1763);
nor U982 (N_982,In_1297,In_41);
and U983 (N_983,In_524,In_1613);
xnor U984 (N_984,In_1550,In_1652);
xnor U985 (N_985,In_545,In_642);
and U986 (N_986,In_738,In_615);
and U987 (N_987,In_1162,In_1382);
and U988 (N_988,In_1810,In_1547);
and U989 (N_989,In_1366,In_1129);
nand U990 (N_990,In_711,In_138);
or U991 (N_991,In_924,In_1215);
nand U992 (N_992,In_1216,In_1939);
nand U993 (N_993,In_199,In_380);
or U994 (N_994,In_917,In_430);
and U995 (N_995,In_667,In_1373);
nor U996 (N_996,In_291,In_1008);
and U997 (N_997,In_652,In_786);
or U998 (N_998,In_544,In_553);
or U999 (N_999,In_803,In_1829);
or U1000 (N_1000,In_1155,In_969);
and U1001 (N_1001,In_1850,In_1411);
nand U1002 (N_1002,In_1972,In_728);
nor U1003 (N_1003,In_1174,In_783);
nand U1004 (N_1004,In_1263,In_1322);
nand U1005 (N_1005,In_1344,In_72);
nor U1006 (N_1006,In_1244,In_900);
or U1007 (N_1007,In_312,In_1541);
and U1008 (N_1008,In_1334,In_1552);
xnor U1009 (N_1009,In_140,In_198);
xor U1010 (N_1010,In_1479,In_619);
nand U1011 (N_1011,In_1013,In_345);
and U1012 (N_1012,In_146,In_140);
nor U1013 (N_1013,In_408,In_48);
or U1014 (N_1014,In_169,In_658);
or U1015 (N_1015,In_1894,In_1756);
nand U1016 (N_1016,In_452,In_730);
nor U1017 (N_1017,In_1064,In_1897);
nand U1018 (N_1018,In_630,In_1144);
xnor U1019 (N_1019,In_132,In_951);
xor U1020 (N_1020,In_603,In_1823);
nand U1021 (N_1021,In_428,In_1275);
nand U1022 (N_1022,In_617,In_1521);
or U1023 (N_1023,In_855,In_155);
nor U1024 (N_1024,In_299,In_1981);
and U1025 (N_1025,In_1990,In_914);
and U1026 (N_1026,In_878,In_1735);
or U1027 (N_1027,In_54,In_575);
nor U1028 (N_1028,In_1672,In_754);
nand U1029 (N_1029,In_832,In_392);
nor U1030 (N_1030,In_1035,In_888);
nor U1031 (N_1031,In_412,In_16);
nand U1032 (N_1032,In_586,In_1041);
and U1033 (N_1033,In_776,In_1582);
nand U1034 (N_1034,In_778,In_696);
nand U1035 (N_1035,In_1236,In_410);
nand U1036 (N_1036,In_618,In_1706);
nand U1037 (N_1037,In_1296,In_94);
and U1038 (N_1038,In_1012,In_1309);
nor U1039 (N_1039,In_943,In_1349);
nor U1040 (N_1040,In_1981,In_1027);
nand U1041 (N_1041,In_1843,In_1199);
and U1042 (N_1042,In_1448,In_349);
nor U1043 (N_1043,In_1758,In_1109);
or U1044 (N_1044,In_911,In_1766);
nand U1045 (N_1045,In_143,In_552);
nor U1046 (N_1046,In_767,In_712);
nor U1047 (N_1047,In_1584,In_1351);
and U1048 (N_1048,In_985,In_1138);
or U1049 (N_1049,In_943,In_444);
and U1050 (N_1050,In_1029,In_1144);
or U1051 (N_1051,In_853,In_214);
nor U1052 (N_1052,In_151,In_990);
and U1053 (N_1053,In_1939,In_840);
and U1054 (N_1054,In_1550,In_279);
or U1055 (N_1055,In_1524,In_29);
and U1056 (N_1056,In_1216,In_218);
nor U1057 (N_1057,In_1780,In_297);
nand U1058 (N_1058,In_700,In_774);
and U1059 (N_1059,In_377,In_93);
nor U1060 (N_1060,In_1101,In_861);
xor U1061 (N_1061,In_1139,In_1650);
nor U1062 (N_1062,In_1968,In_1360);
nor U1063 (N_1063,In_476,In_236);
or U1064 (N_1064,In_230,In_1975);
nand U1065 (N_1065,In_1155,In_1198);
nor U1066 (N_1066,In_1647,In_1514);
and U1067 (N_1067,In_951,In_1526);
and U1068 (N_1068,In_1968,In_1914);
and U1069 (N_1069,In_448,In_982);
and U1070 (N_1070,In_885,In_216);
nor U1071 (N_1071,In_654,In_187);
nor U1072 (N_1072,In_694,In_1833);
nor U1073 (N_1073,In_854,In_1375);
and U1074 (N_1074,In_759,In_1343);
nor U1075 (N_1075,In_1076,In_1330);
and U1076 (N_1076,In_197,In_1693);
and U1077 (N_1077,In_1723,In_1078);
nor U1078 (N_1078,In_868,In_562);
nand U1079 (N_1079,In_1362,In_92);
nand U1080 (N_1080,In_410,In_800);
and U1081 (N_1081,In_1196,In_877);
nor U1082 (N_1082,In_1506,In_103);
or U1083 (N_1083,In_1964,In_1992);
xor U1084 (N_1084,In_1941,In_7);
nand U1085 (N_1085,In_1534,In_173);
nor U1086 (N_1086,In_897,In_1194);
or U1087 (N_1087,In_1284,In_1858);
or U1088 (N_1088,In_218,In_60);
nand U1089 (N_1089,In_1269,In_578);
or U1090 (N_1090,In_1084,In_1802);
nand U1091 (N_1091,In_1382,In_753);
and U1092 (N_1092,In_1158,In_1653);
nor U1093 (N_1093,In_89,In_630);
nor U1094 (N_1094,In_60,In_1606);
nor U1095 (N_1095,In_1404,In_15);
nor U1096 (N_1096,In_1087,In_581);
nand U1097 (N_1097,In_335,In_691);
or U1098 (N_1098,In_1212,In_1688);
and U1099 (N_1099,In_1384,In_923);
or U1100 (N_1100,In_1051,In_376);
or U1101 (N_1101,In_929,In_1330);
nand U1102 (N_1102,In_1527,In_995);
nor U1103 (N_1103,In_1660,In_351);
nor U1104 (N_1104,In_690,In_391);
nor U1105 (N_1105,In_781,In_613);
or U1106 (N_1106,In_630,In_969);
nand U1107 (N_1107,In_1915,In_819);
and U1108 (N_1108,In_98,In_1054);
nor U1109 (N_1109,In_1021,In_1227);
or U1110 (N_1110,In_1817,In_1680);
or U1111 (N_1111,In_1519,In_976);
or U1112 (N_1112,In_688,In_671);
nand U1113 (N_1113,In_1293,In_914);
nor U1114 (N_1114,In_607,In_1024);
nor U1115 (N_1115,In_1500,In_719);
nor U1116 (N_1116,In_1677,In_695);
and U1117 (N_1117,In_842,In_538);
nor U1118 (N_1118,In_220,In_1301);
nor U1119 (N_1119,In_656,In_965);
nand U1120 (N_1120,In_304,In_1983);
nor U1121 (N_1121,In_535,In_224);
and U1122 (N_1122,In_750,In_1058);
or U1123 (N_1123,In_788,In_782);
or U1124 (N_1124,In_1482,In_849);
nand U1125 (N_1125,In_1986,In_1305);
or U1126 (N_1126,In_1702,In_789);
or U1127 (N_1127,In_273,In_1328);
or U1128 (N_1128,In_1739,In_380);
and U1129 (N_1129,In_172,In_1780);
and U1130 (N_1130,In_1301,In_183);
or U1131 (N_1131,In_953,In_60);
nand U1132 (N_1132,In_184,In_1539);
and U1133 (N_1133,In_1258,In_374);
nand U1134 (N_1134,In_1351,In_1562);
and U1135 (N_1135,In_99,In_1142);
xor U1136 (N_1136,In_1894,In_0);
nand U1137 (N_1137,In_1536,In_1714);
or U1138 (N_1138,In_1958,In_730);
nand U1139 (N_1139,In_1480,In_593);
or U1140 (N_1140,In_1407,In_1832);
and U1141 (N_1141,In_1151,In_1097);
nand U1142 (N_1142,In_1780,In_1182);
xnor U1143 (N_1143,In_244,In_1842);
nand U1144 (N_1144,In_1792,In_1652);
xor U1145 (N_1145,In_813,In_1036);
nand U1146 (N_1146,In_923,In_1744);
and U1147 (N_1147,In_1177,In_1175);
and U1148 (N_1148,In_1859,In_1854);
nor U1149 (N_1149,In_919,In_1506);
nand U1150 (N_1150,In_1164,In_419);
nor U1151 (N_1151,In_66,In_294);
or U1152 (N_1152,In_1778,In_1817);
or U1153 (N_1153,In_1125,In_835);
or U1154 (N_1154,In_1317,In_1844);
nor U1155 (N_1155,In_1688,In_1805);
and U1156 (N_1156,In_1383,In_1049);
nand U1157 (N_1157,In_1700,In_1891);
xnor U1158 (N_1158,In_1305,In_16);
xor U1159 (N_1159,In_1893,In_1);
nand U1160 (N_1160,In_0,In_12);
or U1161 (N_1161,In_63,In_1509);
xnor U1162 (N_1162,In_567,In_1043);
nand U1163 (N_1163,In_1882,In_1637);
xnor U1164 (N_1164,In_1748,In_1672);
and U1165 (N_1165,In_999,In_1224);
and U1166 (N_1166,In_1742,In_770);
and U1167 (N_1167,In_1900,In_102);
nand U1168 (N_1168,In_765,In_977);
or U1169 (N_1169,In_652,In_1782);
nand U1170 (N_1170,In_1191,In_1640);
nor U1171 (N_1171,In_912,In_1699);
nor U1172 (N_1172,In_208,In_920);
nand U1173 (N_1173,In_740,In_473);
and U1174 (N_1174,In_1344,In_445);
and U1175 (N_1175,In_1771,In_334);
nand U1176 (N_1176,In_1299,In_1621);
and U1177 (N_1177,In_529,In_1715);
nand U1178 (N_1178,In_757,In_851);
nor U1179 (N_1179,In_1052,In_112);
nand U1180 (N_1180,In_1279,In_1968);
nor U1181 (N_1181,In_1497,In_1531);
or U1182 (N_1182,In_59,In_1714);
nor U1183 (N_1183,In_1117,In_362);
nor U1184 (N_1184,In_230,In_1519);
nor U1185 (N_1185,In_1568,In_1046);
nand U1186 (N_1186,In_607,In_1546);
nor U1187 (N_1187,In_291,In_1116);
or U1188 (N_1188,In_68,In_296);
xor U1189 (N_1189,In_1117,In_1658);
xnor U1190 (N_1190,In_1354,In_1375);
nand U1191 (N_1191,In_1414,In_360);
nor U1192 (N_1192,In_643,In_201);
nor U1193 (N_1193,In_1707,In_1485);
or U1194 (N_1194,In_91,In_1436);
nand U1195 (N_1195,In_1654,In_1343);
or U1196 (N_1196,In_1039,In_889);
or U1197 (N_1197,In_1746,In_282);
xor U1198 (N_1198,In_312,In_1922);
xor U1199 (N_1199,In_1658,In_1355);
and U1200 (N_1200,In_1763,In_399);
or U1201 (N_1201,In_1701,In_1238);
xor U1202 (N_1202,In_798,In_972);
nor U1203 (N_1203,In_1861,In_310);
nor U1204 (N_1204,In_767,In_759);
or U1205 (N_1205,In_52,In_863);
nor U1206 (N_1206,In_1282,In_1640);
nor U1207 (N_1207,In_491,In_1323);
and U1208 (N_1208,In_330,In_1205);
nor U1209 (N_1209,In_611,In_640);
nand U1210 (N_1210,In_1526,In_843);
or U1211 (N_1211,In_913,In_1749);
nor U1212 (N_1212,In_1689,In_549);
and U1213 (N_1213,In_201,In_1356);
xnor U1214 (N_1214,In_1829,In_121);
nor U1215 (N_1215,In_921,In_1783);
nand U1216 (N_1216,In_272,In_1881);
nand U1217 (N_1217,In_1010,In_1606);
nor U1218 (N_1218,In_1266,In_941);
nor U1219 (N_1219,In_335,In_1938);
nor U1220 (N_1220,In_1453,In_1496);
nor U1221 (N_1221,In_585,In_91);
or U1222 (N_1222,In_876,In_872);
or U1223 (N_1223,In_1035,In_1666);
nand U1224 (N_1224,In_612,In_497);
nand U1225 (N_1225,In_177,In_86);
xor U1226 (N_1226,In_1119,In_858);
or U1227 (N_1227,In_708,In_1206);
and U1228 (N_1228,In_1039,In_252);
nor U1229 (N_1229,In_353,In_368);
nor U1230 (N_1230,In_841,In_963);
and U1231 (N_1231,In_1494,In_1592);
nand U1232 (N_1232,In_8,In_907);
or U1233 (N_1233,In_154,In_1134);
nor U1234 (N_1234,In_279,In_482);
nand U1235 (N_1235,In_1621,In_1065);
nor U1236 (N_1236,In_803,In_676);
nor U1237 (N_1237,In_227,In_65);
nor U1238 (N_1238,In_1107,In_410);
nor U1239 (N_1239,In_169,In_1202);
nand U1240 (N_1240,In_601,In_1266);
xor U1241 (N_1241,In_1301,In_291);
nor U1242 (N_1242,In_1716,In_1914);
or U1243 (N_1243,In_1064,In_792);
or U1244 (N_1244,In_826,In_1537);
nor U1245 (N_1245,In_168,In_1389);
nand U1246 (N_1246,In_1467,In_650);
and U1247 (N_1247,In_1837,In_435);
nand U1248 (N_1248,In_639,In_1496);
and U1249 (N_1249,In_441,In_1147);
nand U1250 (N_1250,In_1100,In_1265);
nand U1251 (N_1251,In_915,In_256);
or U1252 (N_1252,In_134,In_361);
xnor U1253 (N_1253,In_740,In_1222);
nand U1254 (N_1254,In_996,In_190);
or U1255 (N_1255,In_840,In_155);
and U1256 (N_1256,In_988,In_1493);
xnor U1257 (N_1257,In_1057,In_1982);
or U1258 (N_1258,In_947,In_1401);
or U1259 (N_1259,In_754,In_1185);
or U1260 (N_1260,In_100,In_370);
nand U1261 (N_1261,In_1349,In_1134);
nor U1262 (N_1262,In_1992,In_804);
nor U1263 (N_1263,In_160,In_1006);
nor U1264 (N_1264,In_765,In_684);
and U1265 (N_1265,In_541,In_1307);
nor U1266 (N_1266,In_80,In_303);
or U1267 (N_1267,In_194,In_1876);
nor U1268 (N_1268,In_1817,In_793);
nand U1269 (N_1269,In_333,In_386);
or U1270 (N_1270,In_787,In_256);
nand U1271 (N_1271,In_1167,In_691);
xnor U1272 (N_1272,In_628,In_286);
or U1273 (N_1273,In_1788,In_1069);
xnor U1274 (N_1274,In_1423,In_1623);
nand U1275 (N_1275,In_1742,In_734);
or U1276 (N_1276,In_96,In_1981);
nand U1277 (N_1277,In_66,In_1859);
and U1278 (N_1278,In_1937,In_1034);
nor U1279 (N_1279,In_589,In_288);
and U1280 (N_1280,In_56,In_1678);
nand U1281 (N_1281,In_1082,In_1024);
and U1282 (N_1282,In_925,In_1646);
nor U1283 (N_1283,In_168,In_1091);
nand U1284 (N_1284,In_947,In_1331);
nor U1285 (N_1285,In_1483,In_1558);
and U1286 (N_1286,In_1611,In_1371);
and U1287 (N_1287,In_1504,In_1231);
or U1288 (N_1288,In_680,In_1815);
nand U1289 (N_1289,In_1477,In_1160);
nand U1290 (N_1290,In_812,In_1704);
or U1291 (N_1291,In_1292,In_1873);
or U1292 (N_1292,In_1154,In_20);
nand U1293 (N_1293,In_1045,In_1042);
xnor U1294 (N_1294,In_1264,In_693);
and U1295 (N_1295,In_640,In_1777);
nor U1296 (N_1296,In_1006,In_1787);
or U1297 (N_1297,In_327,In_533);
nor U1298 (N_1298,In_106,In_1754);
nand U1299 (N_1299,In_1343,In_1078);
nand U1300 (N_1300,In_1052,In_1747);
or U1301 (N_1301,In_1807,In_1980);
nand U1302 (N_1302,In_1474,In_1435);
nand U1303 (N_1303,In_41,In_364);
and U1304 (N_1304,In_1633,In_184);
nand U1305 (N_1305,In_1862,In_1994);
and U1306 (N_1306,In_187,In_1448);
nand U1307 (N_1307,In_1987,In_1788);
and U1308 (N_1308,In_1650,In_873);
or U1309 (N_1309,In_952,In_1519);
nand U1310 (N_1310,In_907,In_1158);
and U1311 (N_1311,In_1146,In_995);
nor U1312 (N_1312,In_345,In_1497);
xnor U1313 (N_1313,In_710,In_995);
nor U1314 (N_1314,In_883,In_517);
nor U1315 (N_1315,In_935,In_1358);
xnor U1316 (N_1316,In_1282,In_1137);
nor U1317 (N_1317,In_155,In_1555);
nand U1318 (N_1318,In_1690,In_1977);
and U1319 (N_1319,In_661,In_1517);
or U1320 (N_1320,In_271,In_1194);
and U1321 (N_1321,In_92,In_1555);
nand U1322 (N_1322,In_1542,In_883);
nor U1323 (N_1323,In_1187,In_1760);
or U1324 (N_1324,In_767,In_1147);
and U1325 (N_1325,In_1505,In_1770);
nor U1326 (N_1326,In_1239,In_758);
and U1327 (N_1327,In_806,In_1631);
xnor U1328 (N_1328,In_1906,In_110);
nor U1329 (N_1329,In_1326,In_1172);
nand U1330 (N_1330,In_323,In_1587);
nand U1331 (N_1331,In_106,In_1761);
nor U1332 (N_1332,In_371,In_824);
and U1333 (N_1333,In_99,In_516);
nor U1334 (N_1334,In_1368,In_1439);
and U1335 (N_1335,In_1840,In_1579);
nor U1336 (N_1336,In_437,In_1603);
or U1337 (N_1337,In_1356,In_1067);
nor U1338 (N_1338,In_1717,In_34);
nor U1339 (N_1339,In_491,In_201);
nor U1340 (N_1340,In_1906,In_153);
nand U1341 (N_1341,In_1596,In_1288);
and U1342 (N_1342,In_1233,In_387);
or U1343 (N_1343,In_494,In_1138);
xor U1344 (N_1344,In_372,In_1459);
or U1345 (N_1345,In_281,In_1102);
nor U1346 (N_1346,In_928,In_918);
nor U1347 (N_1347,In_494,In_673);
and U1348 (N_1348,In_1176,In_1744);
or U1349 (N_1349,In_116,In_1933);
and U1350 (N_1350,In_812,In_1525);
nor U1351 (N_1351,In_1441,In_1666);
xnor U1352 (N_1352,In_1139,In_1258);
nand U1353 (N_1353,In_1478,In_1877);
xnor U1354 (N_1354,In_1013,In_1606);
xnor U1355 (N_1355,In_1664,In_1711);
nor U1356 (N_1356,In_1794,In_1772);
xor U1357 (N_1357,In_987,In_1678);
or U1358 (N_1358,In_672,In_358);
xor U1359 (N_1359,In_1345,In_738);
nand U1360 (N_1360,In_179,In_1932);
or U1361 (N_1361,In_1445,In_140);
xnor U1362 (N_1362,In_1077,In_1921);
and U1363 (N_1363,In_1754,In_1225);
nand U1364 (N_1364,In_169,In_128);
nand U1365 (N_1365,In_1897,In_1834);
nor U1366 (N_1366,In_819,In_1867);
and U1367 (N_1367,In_858,In_728);
nand U1368 (N_1368,In_1988,In_493);
and U1369 (N_1369,In_883,In_552);
or U1370 (N_1370,In_1434,In_919);
nand U1371 (N_1371,In_1793,In_31);
nor U1372 (N_1372,In_169,In_1661);
nor U1373 (N_1373,In_411,In_140);
xor U1374 (N_1374,In_812,In_1626);
or U1375 (N_1375,In_1365,In_974);
and U1376 (N_1376,In_289,In_685);
or U1377 (N_1377,In_1734,In_926);
xnor U1378 (N_1378,In_26,In_1955);
nor U1379 (N_1379,In_554,In_1600);
nor U1380 (N_1380,In_58,In_698);
nand U1381 (N_1381,In_1491,In_1331);
nand U1382 (N_1382,In_508,In_151);
nor U1383 (N_1383,In_566,In_1299);
or U1384 (N_1384,In_654,In_633);
and U1385 (N_1385,In_1709,In_261);
xor U1386 (N_1386,In_12,In_1429);
or U1387 (N_1387,In_1311,In_164);
nor U1388 (N_1388,In_388,In_916);
nand U1389 (N_1389,In_296,In_1676);
or U1390 (N_1390,In_54,In_105);
or U1391 (N_1391,In_644,In_1603);
nor U1392 (N_1392,In_1405,In_305);
nand U1393 (N_1393,In_458,In_163);
nand U1394 (N_1394,In_786,In_399);
xnor U1395 (N_1395,In_1618,In_562);
nor U1396 (N_1396,In_1553,In_93);
nand U1397 (N_1397,In_305,In_1614);
or U1398 (N_1398,In_1993,In_1451);
and U1399 (N_1399,In_449,In_217);
or U1400 (N_1400,In_257,In_698);
nand U1401 (N_1401,In_267,In_1879);
nor U1402 (N_1402,In_289,In_714);
nor U1403 (N_1403,In_1858,In_1105);
and U1404 (N_1404,In_184,In_1055);
nand U1405 (N_1405,In_1575,In_1788);
nor U1406 (N_1406,In_1916,In_836);
or U1407 (N_1407,In_732,In_178);
or U1408 (N_1408,In_1654,In_1083);
and U1409 (N_1409,In_479,In_427);
and U1410 (N_1410,In_104,In_1278);
or U1411 (N_1411,In_793,In_1632);
or U1412 (N_1412,In_1552,In_1484);
nand U1413 (N_1413,In_809,In_1398);
xnor U1414 (N_1414,In_1677,In_114);
nor U1415 (N_1415,In_1528,In_546);
nand U1416 (N_1416,In_563,In_1604);
xnor U1417 (N_1417,In_1073,In_1694);
or U1418 (N_1418,In_808,In_1183);
and U1419 (N_1419,In_1722,In_1652);
or U1420 (N_1420,In_1333,In_247);
and U1421 (N_1421,In_194,In_1634);
xor U1422 (N_1422,In_85,In_67);
or U1423 (N_1423,In_727,In_1023);
or U1424 (N_1424,In_82,In_1024);
nand U1425 (N_1425,In_955,In_1797);
nor U1426 (N_1426,In_1491,In_1748);
nor U1427 (N_1427,In_981,In_1062);
and U1428 (N_1428,In_872,In_963);
nor U1429 (N_1429,In_872,In_1343);
nor U1430 (N_1430,In_57,In_291);
or U1431 (N_1431,In_633,In_135);
nor U1432 (N_1432,In_1089,In_1185);
and U1433 (N_1433,In_406,In_1168);
and U1434 (N_1434,In_1964,In_1909);
nand U1435 (N_1435,In_1697,In_1892);
nor U1436 (N_1436,In_1273,In_921);
or U1437 (N_1437,In_924,In_1972);
xor U1438 (N_1438,In_241,In_117);
or U1439 (N_1439,In_1224,In_1248);
nand U1440 (N_1440,In_1446,In_238);
or U1441 (N_1441,In_1778,In_795);
nand U1442 (N_1442,In_489,In_1313);
nand U1443 (N_1443,In_1496,In_930);
and U1444 (N_1444,In_1072,In_1707);
nor U1445 (N_1445,In_613,In_190);
nand U1446 (N_1446,In_667,In_434);
xnor U1447 (N_1447,In_1586,In_1133);
nor U1448 (N_1448,In_1802,In_1795);
nand U1449 (N_1449,In_1589,In_1015);
or U1450 (N_1450,In_663,In_574);
or U1451 (N_1451,In_1776,In_1887);
xnor U1452 (N_1452,In_1660,In_800);
xnor U1453 (N_1453,In_709,In_83);
xnor U1454 (N_1454,In_1968,In_361);
or U1455 (N_1455,In_94,In_63);
nor U1456 (N_1456,In_762,In_1513);
or U1457 (N_1457,In_62,In_1206);
nor U1458 (N_1458,In_349,In_1356);
nand U1459 (N_1459,In_1330,In_1792);
nand U1460 (N_1460,In_133,In_1679);
nor U1461 (N_1461,In_178,In_768);
nor U1462 (N_1462,In_727,In_1297);
nand U1463 (N_1463,In_885,In_438);
nor U1464 (N_1464,In_845,In_94);
and U1465 (N_1465,In_65,In_208);
xnor U1466 (N_1466,In_1763,In_1660);
or U1467 (N_1467,In_1312,In_1222);
or U1468 (N_1468,In_255,In_536);
nor U1469 (N_1469,In_1895,In_303);
nor U1470 (N_1470,In_319,In_83);
and U1471 (N_1471,In_340,In_1121);
nand U1472 (N_1472,In_1403,In_1326);
nand U1473 (N_1473,In_1831,In_582);
nor U1474 (N_1474,In_1795,In_395);
nand U1475 (N_1475,In_989,In_973);
nand U1476 (N_1476,In_1641,In_27);
or U1477 (N_1477,In_98,In_285);
or U1478 (N_1478,In_19,In_1319);
or U1479 (N_1479,In_1325,In_602);
or U1480 (N_1480,In_1947,In_615);
and U1481 (N_1481,In_993,In_1252);
nor U1482 (N_1482,In_118,In_804);
and U1483 (N_1483,In_372,In_1325);
and U1484 (N_1484,In_1612,In_1119);
nand U1485 (N_1485,In_366,In_553);
nand U1486 (N_1486,In_1315,In_1469);
nor U1487 (N_1487,In_1230,In_121);
nor U1488 (N_1488,In_66,In_1737);
nor U1489 (N_1489,In_1418,In_342);
and U1490 (N_1490,In_1746,In_248);
nor U1491 (N_1491,In_1723,In_1290);
or U1492 (N_1492,In_34,In_1313);
or U1493 (N_1493,In_965,In_1652);
nor U1494 (N_1494,In_1869,In_689);
nand U1495 (N_1495,In_1529,In_1424);
or U1496 (N_1496,In_1477,In_730);
nand U1497 (N_1497,In_710,In_943);
and U1498 (N_1498,In_578,In_844);
nor U1499 (N_1499,In_1094,In_1107);
and U1500 (N_1500,In_834,In_758);
nor U1501 (N_1501,In_1388,In_565);
nor U1502 (N_1502,In_1605,In_1282);
or U1503 (N_1503,In_888,In_1298);
nor U1504 (N_1504,In_301,In_572);
nand U1505 (N_1505,In_1851,In_679);
and U1506 (N_1506,In_631,In_615);
and U1507 (N_1507,In_1810,In_1334);
nor U1508 (N_1508,In_1043,In_408);
and U1509 (N_1509,In_751,In_1646);
nor U1510 (N_1510,In_859,In_877);
nand U1511 (N_1511,In_1135,In_713);
or U1512 (N_1512,In_841,In_1426);
nand U1513 (N_1513,In_1796,In_189);
xnor U1514 (N_1514,In_1322,In_976);
and U1515 (N_1515,In_316,In_1198);
and U1516 (N_1516,In_1636,In_878);
nand U1517 (N_1517,In_1236,In_659);
or U1518 (N_1518,In_507,In_672);
or U1519 (N_1519,In_1712,In_1303);
or U1520 (N_1520,In_232,In_1871);
nand U1521 (N_1521,In_87,In_1859);
or U1522 (N_1522,In_252,In_1317);
and U1523 (N_1523,In_1891,In_830);
xor U1524 (N_1524,In_1659,In_681);
or U1525 (N_1525,In_1757,In_460);
nand U1526 (N_1526,In_1842,In_351);
or U1527 (N_1527,In_230,In_400);
nor U1528 (N_1528,In_440,In_865);
nand U1529 (N_1529,In_346,In_1191);
nand U1530 (N_1530,In_723,In_525);
and U1531 (N_1531,In_1398,In_1561);
and U1532 (N_1532,In_1571,In_1854);
xor U1533 (N_1533,In_686,In_1684);
xor U1534 (N_1534,In_1296,In_1814);
or U1535 (N_1535,In_1428,In_703);
nand U1536 (N_1536,In_399,In_78);
or U1537 (N_1537,In_1148,In_1901);
nand U1538 (N_1538,In_556,In_1920);
nor U1539 (N_1539,In_768,In_425);
or U1540 (N_1540,In_1303,In_1402);
nor U1541 (N_1541,In_263,In_1849);
nor U1542 (N_1542,In_1134,In_1747);
or U1543 (N_1543,In_1835,In_1932);
nor U1544 (N_1544,In_700,In_1062);
and U1545 (N_1545,In_1853,In_276);
nand U1546 (N_1546,In_1808,In_1530);
xor U1547 (N_1547,In_1291,In_277);
nor U1548 (N_1548,In_568,In_259);
nor U1549 (N_1549,In_1072,In_1632);
nor U1550 (N_1550,In_1546,In_235);
xor U1551 (N_1551,In_1515,In_726);
xor U1552 (N_1552,In_1161,In_628);
or U1553 (N_1553,In_1509,In_672);
and U1554 (N_1554,In_1188,In_897);
and U1555 (N_1555,In_1822,In_312);
nor U1556 (N_1556,In_366,In_1462);
and U1557 (N_1557,In_902,In_317);
or U1558 (N_1558,In_565,In_880);
or U1559 (N_1559,In_653,In_1627);
nand U1560 (N_1560,In_143,In_1378);
and U1561 (N_1561,In_1467,In_565);
and U1562 (N_1562,In_1608,In_1970);
xor U1563 (N_1563,In_284,In_34);
nor U1564 (N_1564,In_1960,In_1432);
xnor U1565 (N_1565,In_341,In_710);
nand U1566 (N_1566,In_444,In_1412);
nand U1567 (N_1567,In_1407,In_175);
nand U1568 (N_1568,In_1755,In_905);
nand U1569 (N_1569,In_1494,In_1134);
and U1570 (N_1570,In_1549,In_691);
xor U1571 (N_1571,In_1695,In_1513);
nor U1572 (N_1572,In_1519,In_1524);
or U1573 (N_1573,In_703,In_1623);
nand U1574 (N_1574,In_65,In_1551);
nor U1575 (N_1575,In_627,In_534);
nand U1576 (N_1576,In_1154,In_955);
or U1577 (N_1577,In_1326,In_1931);
nor U1578 (N_1578,In_875,In_748);
or U1579 (N_1579,In_572,In_480);
and U1580 (N_1580,In_1218,In_1006);
or U1581 (N_1581,In_1180,In_882);
nand U1582 (N_1582,In_1695,In_119);
or U1583 (N_1583,In_550,In_1657);
xnor U1584 (N_1584,In_1351,In_259);
and U1585 (N_1585,In_1311,In_1138);
xor U1586 (N_1586,In_1042,In_256);
nand U1587 (N_1587,In_1698,In_1454);
nand U1588 (N_1588,In_1175,In_1519);
nand U1589 (N_1589,In_1141,In_460);
nor U1590 (N_1590,In_580,In_349);
nand U1591 (N_1591,In_1326,In_97);
or U1592 (N_1592,In_1836,In_1180);
and U1593 (N_1593,In_828,In_619);
nor U1594 (N_1594,In_1075,In_434);
and U1595 (N_1595,In_676,In_1769);
and U1596 (N_1596,In_351,In_459);
and U1597 (N_1597,In_1586,In_1653);
or U1598 (N_1598,In_1092,In_1719);
and U1599 (N_1599,In_745,In_808);
nand U1600 (N_1600,In_805,In_305);
or U1601 (N_1601,In_1529,In_633);
and U1602 (N_1602,In_1936,In_513);
nor U1603 (N_1603,In_937,In_962);
xor U1604 (N_1604,In_1124,In_790);
and U1605 (N_1605,In_905,In_1379);
and U1606 (N_1606,In_230,In_682);
xnor U1607 (N_1607,In_21,In_600);
and U1608 (N_1608,In_1217,In_633);
xor U1609 (N_1609,In_1916,In_649);
or U1610 (N_1610,In_1908,In_1264);
or U1611 (N_1611,In_741,In_54);
nand U1612 (N_1612,In_1983,In_1948);
and U1613 (N_1613,In_1468,In_1530);
nor U1614 (N_1614,In_1225,In_797);
or U1615 (N_1615,In_1584,In_1773);
nor U1616 (N_1616,In_1245,In_431);
nor U1617 (N_1617,In_1718,In_736);
or U1618 (N_1618,In_1231,In_539);
and U1619 (N_1619,In_1037,In_1466);
nor U1620 (N_1620,In_194,In_1254);
or U1621 (N_1621,In_1172,In_1640);
nand U1622 (N_1622,In_1080,In_1698);
or U1623 (N_1623,In_374,In_17);
or U1624 (N_1624,In_1448,In_1880);
or U1625 (N_1625,In_43,In_1824);
nand U1626 (N_1626,In_7,In_1947);
nand U1627 (N_1627,In_175,In_1142);
and U1628 (N_1628,In_1309,In_1924);
nor U1629 (N_1629,In_862,In_424);
nor U1630 (N_1630,In_1323,In_678);
and U1631 (N_1631,In_132,In_324);
nor U1632 (N_1632,In_894,In_1444);
or U1633 (N_1633,In_599,In_482);
xnor U1634 (N_1634,In_1674,In_1387);
nand U1635 (N_1635,In_1787,In_1816);
nand U1636 (N_1636,In_1373,In_331);
or U1637 (N_1637,In_708,In_1336);
or U1638 (N_1638,In_313,In_869);
nor U1639 (N_1639,In_1879,In_659);
nand U1640 (N_1640,In_256,In_120);
or U1641 (N_1641,In_728,In_232);
nor U1642 (N_1642,In_1962,In_825);
nor U1643 (N_1643,In_1732,In_991);
and U1644 (N_1644,In_1161,In_814);
nor U1645 (N_1645,In_672,In_702);
or U1646 (N_1646,In_748,In_1532);
xor U1647 (N_1647,In_593,In_1493);
and U1648 (N_1648,In_796,In_1779);
xnor U1649 (N_1649,In_513,In_1697);
and U1650 (N_1650,In_51,In_1229);
and U1651 (N_1651,In_1789,In_518);
or U1652 (N_1652,In_1404,In_63);
and U1653 (N_1653,In_973,In_59);
or U1654 (N_1654,In_1953,In_610);
nor U1655 (N_1655,In_686,In_866);
and U1656 (N_1656,In_1993,In_769);
nand U1657 (N_1657,In_364,In_1485);
or U1658 (N_1658,In_533,In_768);
nand U1659 (N_1659,In_659,In_1131);
or U1660 (N_1660,In_1861,In_370);
and U1661 (N_1661,In_521,In_1303);
nand U1662 (N_1662,In_803,In_84);
nor U1663 (N_1663,In_514,In_1577);
nor U1664 (N_1664,In_1679,In_1071);
nor U1665 (N_1665,In_1997,In_468);
nand U1666 (N_1666,In_1642,In_1320);
and U1667 (N_1667,In_377,In_235);
nand U1668 (N_1668,In_1643,In_1075);
nor U1669 (N_1669,In_1713,In_1160);
and U1670 (N_1670,In_1439,In_413);
xnor U1671 (N_1671,In_1182,In_320);
or U1672 (N_1672,In_25,In_1108);
or U1673 (N_1673,In_1025,In_130);
nor U1674 (N_1674,In_410,In_1491);
nor U1675 (N_1675,In_434,In_219);
xor U1676 (N_1676,In_333,In_973);
or U1677 (N_1677,In_1128,In_1573);
nand U1678 (N_1678,In_1252,In_691);
and U1679 (N_1679,In_351,In_1342);
nor U1680 (N_1680,In_774,In_400);
nand U1681 (N_1681,In_1809,In_1190);
or U1682 (N_1682,In_158,In_928);
or U1683 (N_1683,In_1026,In_1390);
nor U1684 (N_1684,In_634,In_979);
nand U1685 (N_1685,In_1227,In_1032);
or U1686 (N_1686,In_279,In_1246);
and U1687 (N_1687,In_376,In_1062);
nor U1688 (N_1688,In_1999,In_1148);
nand U1689 (N_1689,In_1901,In_1087);
and U1690 (N_1690,In_919,In_1500);
or U1691 (N_1691,In_650,In_403);
or U1692 (N_1692,In_1655,In_35);
or U1693 (N_1693,In_1298,In_603);
nand U1694 (N_1694,In_1635,In_1413);
or U1695 (N_1695,In_1708,In_1852);
nand U1696 (N_1696,In_391,In_233);
nand U1697 (N_1697,In_987,In_1212);
nand U1698 (N_1698,In_563,In_251);
or U1699 (N_1699,In_1177,In_1820);
or U1700 (N_1700,In_1151,In_262);
nand U1701 (N_1701,In_1481,In_279);
xor U1702 (N_1702,In_1460,In_261);
nand U1703 (N_1703,In_1588,In_1598);
nand U1704 (N_1704,In_1083,In_74);
and U1705 (N_1705,In_1885,In_803);
nor U1706 (N_1706,In_1356,In_228);
nor U1707 (N_1707,In_281,In_1106);
nand U1708 (N_1708,In_1482,In_1283);
or U1709 (N_1709,In_1961,In_204);
nand U1710 (N_1710,In_479,In_198);
nand U1711 (N_1711,In_1334,In_379);
or U1712 (N_1712,In_1309,In_1691);
nand U1713 (N_1713,In_1425,In_1927);
nor U1714 (N_1714,In_1407,In_1979);
xor U1715 (N_1715,In_542,In_475);
and U1716 (N_1716,In_341,In_641);
and U1717 (N_1717,In_246,In_90);
nand U1718 (N_1718,In_1501,In_1938);
or U1719 (N_1719,In_1117,In_100);
nand U1720 (N_1720,In_1992,In_787);
nand U1721 (N_1721,In_1573,In_1126);
xor U1722 (N_1722,In_160,In_1115);
xnor U1723 (N_1723,In_1065,In_1777);
and U1724 (N_1724,In_1413,In_689);
or U1725 (N_1725,In_1647,In_1047);
or U1726 (N_1726,In_1715,In_1792);
and U1727 (N_1727,In_586,In_1318);
nor U1728 (N_1728,In_637,In_1487);
or U1729 (N_1729,In_1762,In_945);
and U1730 (N_1730,In_1673,In_806);
xor U1731 (N_1731,In_1588,In_1019);
nand U1732 (N_1732,In_292,In_1458);
xor U1733 (N_1733,In_1622,In_1733);
nand U1734 (N_1734,In_38,In_26);
nand U1735 (N_1735,In_32,In_990);
nor U1736 (N_1736,In_585,In_873);
or U1737 (N_1737,In_1064,In_1690);
and U1738 (N_1738,In_387,In_1728);
xor U1739 (N_1739,In_182,In_1061);
nor U1740 (N_1740,In_1544,In_1352);
or U1741 (N_1741,In_725,In_1160);
and U1742 (N_1742,In_386,In_431);
and U1743 (N_1743,In_815,In_1950);
nand U1744 (N_1744,In_1199,In_1350);
nor U1745 (N_1745,In_693,In_1054);
xor U1746 (N_1746,In_1337,In_27);
xor U1747 (N_1747,In_1572,In_748);
nand U1748 (N_1748,In_995,In_838);
and U1749 (N_1749,In_1600,In_1030);
nand U1750 (N_1750,In_1254,In_1365);
and U1751 (N_1751,In_291,In_352);
nor U1752 (N_1752,In_371,In_680);
and U1753 (N_1753,In_1409,In_343);
or U1754 (N_1754,In_1641,In_208);
nand U1755 (N_1755,In_1062,In_1776);
nor U1756 (N_1756,In_1174,In_1906);
nor U1757 (N_1757,In_1588,In_610);
nand U1758 (N_1758,In_546,In_1944);
nand U1759 (N_1759,In_614,In_100);
nor U1760 (N_1760,In_1451,In_1067);
xor U1761 (N_1761,In_1587,In_718);
nor U1762 (N_1762,In_1282,In_283);
and U1763 (N_1763,In_582,In_1907);
nor U1764 (N_1764,In_283,In_1451);
and U1765 (N_1765,In_1347,In_1733);
nor U1766 (N_1766,In_1967,In_437);
nor U1767 (N_1767,In_1794,In_1001);
and U1768 (N_1768,In_798,In_97);
nand U1769 (N_1769,In_1319,In_592);
nand U1770 (N_1770,In_1331,In_772);
nor U1771 (N_1771,In_1776,In_1023);
and U1772 (N_1772,In_422,In_1973);
and U1773 (N_1773,In_1376,In_1753);
or U1774 (N_1774,In_1964,In_321);
and U1775 (N_1775,In_235,In_205);
or U1776 (N_1776,In_1756,In_1169);
nor U1777 (N_1777,In_507,In_1126);
and U1778 (N_1778,In_57,In_802);
nor U1779 (N_1779,In_998,In_1037);
nor U1780 (N_1780,In_1462,In_458);
nand U1781 (N_1781,In_113,In_134);
or U1782 (N_1782,In_1451,In_460);
or U1783 (N_1783,In_1252,In_786);
nand U1784 (N_1784,In_1151,In_280);
nand U1785 (N_1785,In_44,In_617);
or U1786 (N_1786,In_1045,In_202);
nor U1787 (N_1787,In_291,In_1341);
or U1788 (N_1788,In_1131,In_116);
and U1789 (N_1789,In_532,In_273);
xor U1790 (N_1790,In_875,In_1961);
nor U1791 (N_1791,In_1927,In_890);
nor U1792 (N_1792,In_1662,In_1138);
and U1793 (N_1793,In_1565,In_123);
nor U1794 (N_1794,In_1660,In_794);
xor U1795 (N_1795,In_181,In_564);
and U1796 (N_1796,In_623,In_917);
xnor U1797 (N_1797,In_484,In_1943);
or U1798 (N_1798,In_514,In_842);
nand U1799 (N_1799,In_1392,In_1369);
and U1800 (N_1800,In_589,In_353);
nor U1801 (N_1801,In_127,In_1287);
nand U1802 (N_1802,In_1979,In_1475);
nand U1803 (N_1803,In_427,In_341);
nand U1804 (N_1804,In_1380,In_1999);
nor U1805 (N_1805,In_1660,In_77);
nor U1806 (N_1806,In_506,In_263);
nor U1807 (N_1807,In_995,In_338);
or U1808 (N_1808,In_1542,In_629);
nand U1809 (N_1809,In_419,In_1172);
nand U1810 (N_1810,In_167,In_100);
nor U1811 (N_1811,In_1718,In_58);
nor U1812 (N_1812,In_820,In_1866);
nand U1813 (N_1813,In_539,In_1576);
and U1814 (N_1814,In_388,In_527);
or U1815 (N_1815,In_1093,In_905);
nor U1816 (N_1816,In_1796,In_904);
and U1817 (N_1817,In_1261,In_163);
and U1818 (N_1818,In_1508,In_1686);
nand U1819 (N_1819,In_647,In_614);
nor U1820 (N_1820,In_444,In_410);
or U1821 (N_1821,In_1903,In_1098);
or U1822 (N_1822,In_826,In_1706);
xor U1823 (N_1823,In_526,In_632);
xnor U1824 (N_1824,In_1565,In_1889);
nor U1825 (N_1825,In_1398,In_1308);
and U1826 (N_1826,In_1680,In_995);
and U1827 (N_1827,In_489,In_856);
xor U1828 (N_1828,In_462,In_1510);
and U1829 (N_1829,In_1155,In_1478);
nor U1830 (N_1830,In_760,In_1465);
or U1831 (N_1831,In_166,In_516);
nor U1832 (N_1832,In_1757,In_1440);
and U1833 (N_1833,In_641,In_272);
nor U1834 (N_1834,In_1425,In_1063);
or U1835 (N_1835,In_534,In_1710);
nand U1836 (N_1836,In_860,In_1380);
nor U1837 (N_1837,In_1446,In_1862);
or U1838 (N_1838,In_1019,In_920);
and U1839 (N_1839,In_668,In_229);
nand U1840 (N_1840,In_1527,In_510);
and U1841 (N_1841,In_763,In_265);
nand U1842 (N_1842,In_1793,In_1693);
and U1843 (N_1843,In_1941,In_1502);
and U1844 (N_1844,In_719,In_1917);
nor U1845 (N_1845,In_1555,In_339);
or U1846 (N_1846,In_876,In_1991);
xor U1847 (N_1847,In_1383,In_741);
nand U1848 (N_1848,In_78,In_41);
nor U1849 (N_1849,In_1120,In_669);
or U1850 (N_1850,In_317,In_909);
nor U1851 (N_1851,In_233,In_60);
and U1852 (N_1852,In_1926,In_485);
or U1853 (N_1853,In_1194,In_1463);
or U1854 (N_1854,In_1092,In_1434);
xnor U1855 (N_1855,In_15,In_1306);
or U1856 (N_1856,In_1888,In_1146);
and U1857 (N_1857,In_211,In_876);
or U1858 (N_1858,In_1589,In_1126);
nand U1859 (N_1859,In_1279,In_1165);
nand U1860 (N_1860,In_431,In_1975);
nor U1861 (N_1861,In_1368,In_557);
nand U1862 (N_1862,In_968,In_479);
xnor U1863 (N_1863,In_721,In_862);
and U1864 (N_1864,In_1720,In_1249);
or U1865 (N_1865,In_1939,In_1543);
xnor U1866 (N_1866,In_1403,In_1786);
xnor U1867 (N_1867,In_999,In_304);
and U1868 (N_1868,In_1734,In_99);
and U1869 (N_1869,In_517,In_1676);
nand U1870 (N_1870,In_702,In_980);
xnor U1871 (N_1871,In_1009,In_1002);
and U1872 (N_1872,In_1727,In_1538);
nor U1873 (N_1873,In_1818,In_102);
and U1874 (N_1874,In_1036,In_640);
xnor U1875 (N_1875,In_370,In_1371);
nand U1876 (N_1876,In_590,In_614);
xnor U1877 (N_1877,In_469,In_1084);
and U1878 (N_1878,In_434,In_815);
nor U1879 (N_1879,In_817,In_1346);
or U1880 (N_1880,In_1882,In_4);
and U1881 (N_1881,In_404,In_1202);
and U1882 (N_1882,In_826,In_1127);
nor U1883 (N_1883,In_1695,In_842);
xor U1884 (N_1884,In_1997,In_1122);
or U1885 (N_1885,In_67,In_1306);
or U1886 (N_1886,In_292,In_875);
or U1887 (N_1887,In_1477,In_75);
xnor U1888 (N_1888,In_1556,In_1904);
or U1889 (N_1889,In_957,In_1128);
or U1890 (N_1890,In_843,In_1970);
nor U1891 (N_1891,In_1911,In_807);
nand U1892 (N_1892,In_1377,In_585);
and U1893 (N_1893,In_985,In_50);
nor U1894 (N_1894,In_1513,In_1432);
and U1895 (N_1895,In_446,In_1029);
or U1896 (N_1896,In_346,In_1391);
nor U1897 (N_1897,In_1639,In_1119);
nor U1898 (N_1898,In_1991,In_1724);
and U1899 (N_1899,In_672,In_1858);
nand U1900 (N_1900,In_1717,In_142);
nor U1901 (N_1901,In_172,In_1723);
or U1902 (N_1902,In_1812,In_1330);
and U1903 (N_1903,In_553,In_1599);
and U1904 (N_1904,In_1566,In_1685);
nand U1905 (N_1905,In_774,In_179);
nor U1906 (N_1906,In_780,In_238);
and U1907 (N_1907,In_18,In_1662);
or U1908 (N_1908,In_1414,In_867);
and U1909 (N_1909,In_1255,In_1921);
nand U1910 (N_1910,In_1406,In_1737);
or U1911 (N_1911,In_861,In_632);
nor U1912 (N_1912,In_211,In_602);
or U1913 (N_1913,In_226,In_717);
and U1914 (N_1914,In_728,In_1704);
nor U1915 (N_1915,In_1438,In_499);
nor U1916 (N_1916,In_874,In_1784);
or U1917 (N_1917,In_105,In_1811);
nor U1918 (N_1918,In_264,In_6);
nand U1919 (N_1919,In_682,In_1008);
or U1920 (N_1920,In_1563,In_754);
nor U1921 (N_1921,In_680,In_726);
nor U1922 (N_1922,In_1337,In_1909);
nand U1923 (N_1923,In_858,In_1483);
and U1924 (N_1924,In_264,In_1651);
nor U1925 (N_1925,In_1784,In_164);
nand U1926 (N_1926,In_150,In_384);
or U1927 (N_1927,In_190,In_115);
xnor U1928 (N_1928,In_922,In_659);
or U1929 (N_1929,In_1382,In_356);
or U1930 (N_1930,In_1611,In_1240);
and U1931 (N_1931,In_374,In_593);
nor U1932 (N_1932,In_308,In_1507);
and U1933 (N_1933,In_1840,In_1251);
nor U1934 (N_1934,In_1187,In_1273);
nand U1935 (N_1935,In_672,In_689);
nand U1936 (N_1936,In_908,In_1983);
nor U1937 (N_1937,In_1001,In_770);
nand U1938 (N_1938,In_1760,In_1018);
nand U1939 (N_1939,In_72,In_1432);
xor U1940 (N_1940,In_685,In_271);
nor U1941 (N_1941,In_1548,In_1542);
nor U1942 (N_1942,In_546,In_807);
nand U1943 (N_1943,In_1857,In_1150);
nor U1944 (N_1944,In_807,In_336);
and U1945 (N_1945,In_800,In_1050);
and U1946 (N_1946,In_1277,In_257);
and U1947 (N_1947,In_1571,In_113);
and U1948 (N_1948,In_1278,In_1048);
and U1949 (N_1949,In_913,In_1989);
or U1950 (N_1950,In_1223,In_814);
and U1951 (N_1951,In_483,In_805);
nand U1952 (N_1952,In_1725,In_1552);
or U1953 (N_1953,In_313,In_424);
and U1954 (N_1954,In_726,In_1960);
nor U1955 (N_1955,In_4,In_848);
or U1956 (N_1956,In_910,In_186);
and U1957 (N_1957,In_1962,In_3);
nand U1958 (N_1958,In_1383,In_1473);
nand U1959 (N_1959,In_407,In_1938);
nand U1960 (N_1960,In_861,In_140);
or U1961 (N_1961,In_851,In_620);
or U1962 (N_1962,In_1501,In_445);
xor U1963 (N_1963,In_1633,In_1638);
nand U1964 (N_1964,In_745,In_1035);
or U1965 (N_1965,In_1178,In_570);
xor U1966 (N_1966,In_1294,In_1198);
and U1967 (N_1967,In_254,In_517);
or U1968 (N_1968,In_120,In_1602);
xor U1969 (N_1969,In_489,In_1053);
nor U1970 (N_1970,In_395,In_1344);
nor U1971 (N_1971,In_1535,In_1576);
and U1972 (N_1972,In_819,In_740);
or U1973 (N_1973,In_1110,In_54);
or U1974 (N_1974,In_89,In_1070);
or U1975 (N_1975,In_488,In_1167);
nand U1976 (N_1976,In_948,In_1299);
nand U1977 (N_1977,In_385,In_464);
nand U1978 (N_1978,In_555,In_72);
nor U1979 (N_1979,In_476,In_597);
nor U1980 (N_1980,In_1970,In_1620);
or U1981 (N_1981,In_1471,In_1283);
nor U1982 (N_1982,In_105,In_328);
and U1983 (N_1983,In_888,In_771);
and U1984 (N_1984,In_185,In_154);
or U1985 (N_1985,In_100,In_1191);
and U1986 (N_1986,In_518,In_1900);
nor U1987 (N_1987,In_1960,In_1169);
nand U1988 (N_1988,In_1274,In_470);
nor U1989 (N_1989,In_788,In_565);
nor U1990 (N_1990,In_440,In_727);
nor U1991 (N_1991,In_1331,In_332);
and U1992 (N_1992,In_1644,In_1670);
xnor U1993 (N_1993,In_697,In_1773);
and U1994 (N_1994,In_42,In_1220);
nor U1995 (N_1995,In_1646,In_483);
or U1996 (N_1996,In_936,In_889);
or U1997 (N_1997,In_538,In_703);
xor U1998 (N_1998,In_1819,In_1320);
xnor U1999 (N_1999,In_713,In_502);
and U2000 (N_2000,In_715,In_1750);
and U2001 (N_2001,In_251,In_845);
xnor U2002 (N_2002,In_1397,In_238);
or U2003 (N_2003,In_1107,In_1896);
nor U2004 (N_2004,In_936,In_1293);
nor U2005 (N_2005,In_1314,In_1818);
and U2006 (N_2006,In_804,In_1342);
and U2007 (N_2007,In_952,In_1941);
nand U2008 (N_2008,In_278,In_138);
or U2009 (N_2009,In_1424,In_87);
or U2010 (N_2010,In_288,In_1461);
nor U2011 (N_2011,In_425,In_993);
nand U2012 (N_2012,In_472,In_1264);
nand U2013 (N_2013,In_1773,In_1635);
nor U2014 (N_2014,In_1339,In_511);
nand U2015 (N_2015,In_1821,In_1225);
nor U2016 (N_2016,In_1127,In_500);
or U2017 (N_2017,In_1696,In_462);
xor U2018 (N_2018,In_1669,In_714);
or U2019 (N_2019,In_1842,In_316);
nor U2020 (N_2020,In_1342,In_1815);
or U2021 (N_2021,In_520,In_1441);
nor U2022 (N_2022,In_1108,In_1341);
nor U2023 (N_2023,In_607,In_1772);
nor U2024 (N_2024,In_510,In_1672);
and U2025 (N_2025,In_493,In_378);
xnor U2026 (N_2026,In_1455,In_1167);
nor U2027 (N_2027,In_644,In_690);
and U2028 (N_2028,In_1492,In_623);
and U2029 (N_2029,In_1726,In_1914);
nor U2030 (N_2030,In_1927,In_1429);
or U2031 (N_2031,In_729,In_1217);
xnor U2032 (N_2032,In_1246,In_627);
and U2033 (N_2033,In_566,In_874);
nor U2034 (N_2034,In_1179,In_1213);
nand U2035 (N_2035,In_1602,In_542);
and U2036 (N_2036,In_878,In_480);
or U2037 (N_2037,In_196,In_647);
or U2038 (N_2038,In_1745,In_885);
or U2039 (N_2039,In_1047,In_1853);
and U2040 (N_2040,In_1998,In_809);
or U2041 (N_2041,In_604,In_1643);
or U2042 (N_2042,In_853,In_1922);
nor U2043 (N_2043,In_1243,In_1641);
xnor U2044 (N_2044,In_1750,In_1183);
nor U2045 (N_2045,In_531,In_1198);
and U2046 (N_2046,In_531,In_1421);
and U2047 (N_2047,In_1731,In_640);
xnor U2048 (N_2048,In_1920,In_369);
and U2049 (N_2049,In_1425,In_1098);
nand U2050 (N_2050,In_1620,In_1861);
nor U2051 (N_2051,In_1482,In_1813);
and U2052 (N_2052,In_169,In_1866);
nand U2053 (N_2053,In_1882,In_395);
and U2054 (N_2054,In_1911,In_1747);
and U2055 (N_2055,In_259,In_1937);
and U2056 (N_2056,In_1456,In_124);
nand U2057 (N_2057,In_1072,In_1429);
nor U2058 (N_2058,In_1286,In_512);
nor U2059 (N_2059,In_1602,In_1452);
or U2060 (N_2060,In_683,In_129);
nand U2061 (N_2061,In_436,In_503);
nor U2062 (N_2062,In_151,In_1651);
nor U2063 (N_2063,In_158,In_1241);
or U2064 (N_2064,In_1018,In_1096);
or U2065 (N_2065,In_158,In_1522);
or U2066 (N_2066,In_655,In_1952);
and U2067 (N_2067,In_1710,In_828);
or U2068 (N_2068,In_169,In_1594);
xnor U2069 (N_2069,In_711,In_575);
xor U2070 (N_2070,In_875,In_985);
nor U2071 (N_2071,In_161,In_1282);
nor U2072 (N_2072,In_1444,In_851);
nand U2073 (N_2073,In_364,In_278);
and U2074 (N_2074,In_1301,In_399);
nand U2075 (N_2075,In_1757,In_1219);
nor U2076 (N_2076,In_1146,In_1340);
nand U2077 (N_2077,In_1362,In_430);
nor U2078 (N_2078,In_967,In_841);
or U2079 (N_2079,In_1737,In_1574);
nor U2080 (N_2080,In_1728,In_589);
and U2081 (N_2081,In_216,In_1801);
or U2082 (N_2082,In_1221,In_160);
and U2083 (N_2083,In_1393,In_1552);
or U2084 (N_2084,In_990,In_781);
or U2085 (N_2085,In_239,In_1969);
or U2086 (N_2086,In_13,In_1316);
nor U2087 (N_2087,In_256,In_1639);
nor U2088 (N_2088,In_1268,In_1116);
and U2089 (N_2089,In_1504,In_1953);
nand U2090 (N_2090,In_1192,In_351);
nand U2091 (N_2091,In_1969,In_1361);
or U2092 (N_2092,In_1252,In_680);
or U2093 (N_2093,In_862,In_744);
or U2094 (N_2094,In_1286,In_650);
or U2095 (N_2095,In_1487,In_877);
nor U2096 (N_2096,In_1505,In_964);
or U2097 (N_2097,In_1945,In_1954);
nor U2098 (N_2098,In_1846,In_1272);
nand U2099 (N_2099,In_1475,In_1252);
xor U2100 (N_2100,In_224,In_1833);
nor U2101 (N_2101,In_181,In_563);
nand U2102 (N_2102,In_46,In_1341);
nand U2103 (N_2103,In_1828,In_1732);
nand U2104 (N_2104,In_1598,In_1017);
and U2105 (N_2105,In_1450,In_1599);
nand U2106 (N_2106,In_1277,In_628);
xor U2107 (N_2107,In_461,In_1932);
nor U2108 (N_2108,In_1859,In_837);
and U2109 (N_2109,In_1959,In_444);
nand U2110 (N_2110,In_1981,In_1428);
nor U2111 (N_2111,In_1246,In_1963);
nand U2112 (N_2112,In_701,In_726);
or U2113 (N_2113,In_1734,In_577);
nand U2114 (N_2114,In_1299,In_1470);
nor U2115 (N_2115,In_1312,In_482);
or U2116 (N_2116,In_159,In_1572);
and U2117 (N_2117,In_255,In_281);
nor U2118 (N_2118,In_404,In_1133);
and U2119 (N_2119,In_1538,In_568);
nand U2120 (N_2120,In_579,In_1216);
and U2121 (N_2121,In_521,In_106);
or U2122 (N_2122,In_89,In_807);
or U2123 (N_2123,In_377,In_1140);
xor U2124 (N_2124,In_1365,In_1437);
nor U2125 (N_2125,In_1832,In_779);
or U2126 (N_2126,In_647,In_290);
nor U2127 (N_2127,In_210,In_975);
and U2128 (N_2128,In_374,In_1103);
and U2129 (N_2129,In_359,In_1022);
nor U2130 (N_2130,In_162,In_1404);
xor U2131 (N_2131,In_606,In_1837);
or U2132 (N_2132,In_1054,In_855);
nor U2133 (N_2133,In_1379,In_586);
and U2134 (N_2134,In_1623,In_440);
and U2135 (N_2135,In_203,In_91);
or U2136 (N_2136,In_1621,In_1233);
nand U2137 (N_2137,In_874,In_1191);
and U2138 (N_2138,In_1420,In_1046);
nand U2139 (N_2139,In_1756,In_175);
nor U2140 (N_2140,In_835,In_842);
or U2141 (N_2141,In_1622,In_411);
and U2142 (N_2142,In_1188,In_867);
nand U2143 (N_2143,In_1659,In_1695);
and U2144 (N_2144,In_889,In_1033);
nand U2145 (N_2145,In_861,In_996);
and U2146 (N_2146,In_1367,In_296);
nand U2147 (N_2147,In_864,In_1635);
and U2148 (N_2148,In_1325,In_812);
and U2149 (N_2149,In_1076,In_2);
or U2150 (N_2150,In_1348,In_1698);
and U2151 (N_2151,In_985,In_1292);
nor U2152 (N_2152,In_1324,In_673);
nor U2153 (N_2153,In_1734,In_1079);
nand U2154 (N_2154,In_1198,In_1982);
nor U2155 (N_2155,In_1917,In_0);
and U2156 (N_2156,In_1099,In_653);
nor U2157 (N_2157,In_1523,In_1796);
or U2158 (N_2158,In_1118,In_1304);
nand U2159 (N_2159,In_299,In_1706);
or U2160 (N_2160,In_1893,In_711);
or U2161 (N_2161,In_382,In_1873);
or U2162 (N_2162,In_1636,In_1158);
nand U2163 (N_2163,In_1507,In_920);
nor U2164 (N_2164,In_1660,In_92);
nand U2165 (N_2165,In_943,In_173);
and U2166 (N_2166,In_752,In_961);
and U2167 (N_2167,In_1821,In_848);
nor U2168 (N_2168,In_795,In_857);
or U2169 (N_2169,In_1510,In_167);
xor U2170 (N_2170,In_1585,In_497);
or U2171 (N_2171,In_727,In_1530);
or U2172 (N_2172,In_1440,In_634);
nor U2173 (N_2173,In_295,In_569);
nor U2174 (N_2174,In_1991,In_372);
and U2175 (N_2175,In_677,In_252);
nor U2176 (N_2176,In_422,In_363);
and U2177 (N_2177,In_981,In_1512);
or U2178 (N_2178,In_1805,In_786);
nand U2179 (N_2179,In_546,In_279);
nor U2180 (N_2180,In_1697,In_1330);
nand U2181 (N_2181,In_171,In_1485);
xnor U2182 (N_2182,In_906,In_1792);
nand U2183 (N_2183,In_1346,In_1731);
and U2184 (N_2184,In_1726,In_392);
nor U2185 (N_2185,In_102,In_798);
nand U2186 (N_2186,In_599,In_622);
or U2187 (N_2187,In_516,In_242);
and U2188 (N_2188,In_1329,In_699);
xor U2189 (N_2189,In_1093,In_1747);
nand U2190 (N_2190,In_1206,In_423);
nand U2191 (N_2191,In_234,In_1401);
nand U2192 (N_2192,In_299,In_661);
nor U2193 (N_2193,In_992,In_1133);
nor U2194 (N_2194,In_1526,In_622);
or U2195 (N_2195,In_310,In_982);
nor U2196 (N_2196,In_1042,In_681);
nor U2197 (N_2197,In_1213,In_1116);
nor U2198 (N_2198,In_422,In_1231);
nor U2199 (N_2199,In_177,In_1340);
nor U2200 (N_2200,In_1610,In_142);
and U2201 (N_2201,In_731,In_825);
nor U2202 (N_2202,In_824,In_494);
and U2203 (N_2203,In_957,In_1658);
and U2204 (N_2204,In_611,In_1608);
nand U2205 (N_2205,In_1522,In_1317);
nand U2206 (N_2206,In_1825,In_903);
nand U2207 (N_2207,In_1714,In_990);
nand U2208 (N_2208,In_1693,In_1561);
nand U2209 (N_2209,In_1243,In_947);
nor U2210 (N_2210,In_459,In_541);
nor U2211 (N_2211,In_1444,In_921);
and U2212 (N_2212,In_443,In_1800);
or U2213 (N_2213,In_593,In_1289);
and U2214 (N_2214,In_722,In_239);
and U2215 (N_2215,In_1104,In_26);
or U2216 (N_2216,In_141,In_599);
nand U2217 (N_2217,In_576,In_1574);
nor U2218 (N_2218,In_305,In_738);
and U2219 (N_2219,In_1842,In_1778);
or U2220 (N_2220,In_1183,In_847);
nand U2221 (N_2221,In_1688,In_765);
and U2222 (N_2222,In_26,In_231);
nor U2223 (N_2223,In_463,In_28);
or U2224 (N_2224,In_1383,In_977);
nor U2225 (N_2225,In_304,In_1518);
nand U2226 (N_2226,In_1890,In_1471);
nand U2227 (N_2227,In_456,In_1783);
nand U2228 (N_2228,In_1095,In_1169);
nor U2229 (N_2229,In_1931,In_781);
nand U2230 (N_2230,In_335,In_371);
and U2231 (N_2231,In_222,In_669);
or U2232 (N_2232,In_1667,In_1829);
or U2233 (N_2233,In_114,In_1244);
nor U2234 (N_2234,In_38,In_1911);
xor U2235 (N_2235,In_564,In_1586);
or U2236 (N_2236,In_1285,In_1011);
nand U2237 (N_2237,In_1060,In_508);
or U2238 (N_2238,In_361,In_80);
nor U2239 (N_2239,In_902,In_444);
or U2240 (N_2240,In_1160,In_1591);
xnor U2241 (N_2241,In_1147,In_1233);
nand U2242 (N_2242,In_1258,In_654);
nor U2243 (N_2243,In_119,In_1136);
and U2244 (N_2244,In_1584,In_750);
nor U2245 (N_2245,In_1092,In_483);
nand U2246 (N_2246,In_71,In_634);
and U2247 (N_2247,In_1092,In_1407);
xor U2248 (N_2248,In_1272,In_1620);
nand U2249 (N_2249,In_85,In_242);
nand U2250 (N_2250,In_1703,In_1767);
nand U2251 (N_2251,In_1555,In_864);
and U2252 (N_2252,In_1885,In_523);
and U2253 (N_2253,In_1894,In_612);
and U2254 (N_2254,In_1675,In_1011);
nor U2255 (N_2255,In_176,In_58);
xnor U2256 (N_2256,In_493,In_1385);
nand U2257 (N_2257,In_716,In_1932);
and U2258 (N_2258,In_102,In_870);
or U2259 (N_2259,In_1306,In_290);
xor U2260 (N_2260,In_1322,In_1803);
nand U2261 (N_2261,In_1787,In_1286);
and U2262 (N_2262,In_1103,In_580);
or U2263 (N_2263,In_1411,In_300);
xor U2264 (N_2264,In_230,In_1268);
nor U2265 (N_2265,In_1803,In_917);
nor U2266 (N_2266,In_1226,In_874);
and U2267 (N_2267,In_489,In_1126);
or U2268 (N_2268,In_437,In_540);
and U2269 (N_2269,In_464,In_976);
or U2270 (N_2270,In_744,In_464);
xor U2271 (N_2271,In_168,In_1708);
nor U2272 (N_2272,In_1138,In_805);
nor U2273 (N_2273,In_660,In_1511);
or U2274 (N_2274,In_262,In_1839);
nand U2275 (N_2275,In_1305,In_221);
or U2276 (N_2276,In_1262,In_142);
and U2277 (N_2277,In_622,In_1680);
nor U2278 (N_2278,In_1378,In_1999);
and U2279 (N_2279,In_667,In_1593);
or U2280 (N_2280,In_540,In_1777);
or U2281 (N_2281,In_486,In_659);
nor U2282 (N_2282,In_1397,In_966);
or U2283 (N_2283,In_558,In_1188);
xor U2284 (N_2284,In_1432,In_3);
and U2285 (N_2285,In_732,In_1535);
nor U2286 (N_2286,In_48,In_328);
or U2287 (N_2287,In_1674,In_1421);
nor U2288 (N_2288,In_1449,In_331);
and U2289 (N_2289,In_1295,In_1032);
and U2290 (N_2290,In_1804,In_516);
nand U2291 (N_2291,In_581,In_15);
nand U2292 (N_2292,In_807,In_1577);
nor U2293 (N_2293,In_1258,In_1455);
nor U2294 (N_2294,In_1921,In_1640);
xor U2295 (N_2295,In_1601,In_1109);
nor U2296 (N_2296,In_1118,In_1269);
or U2297 (N_2297,In_845,In_1576);
nor U2298 (N_2298,In_1088,In_1258);
nand U2299 (N_2299,In_781,In_1394);
xnor U2300 (N_2300,In_1975,In_1264);
nor U2301 (N_2301,In_1284,In_335);
nand U2302 (N_2302,In_155,In_1103);
or U2303 (N_2303,In_1318,In_1670);
nor U2304 (N_2304,In_1663,In_476);
nand U2305 (N_2305,In_1564,In_294);
nor U2306 (N_2306,In_1442,In_840);
nand U2307 (N_2307,In_1925,In_606);
or U2308 (N_2308,In_408,In_1248);
or U2309 (N_2309,In_1958,In_1447);
or U2310 (N_2310,In_405,In_1138);
nor U2311 (N_2311,In_1771,In_1015);
nor U2312 (N_2312,In_1754,In_1921);
nand U2313 (N_2313,In_475,In_958);
and U2314 (N_2314,In_562,In_941);
or U2315 (N_2315,In_1578,In_1933);
and U2316 (N_2316,In_583,In_588);
and U2317 (N_2317,In_1100,In_272);
or U2318 (N_2318,In_911,In_1156);
nor U2319 (N_2319,In_772,In_1317);
and U2320 (N_2320,In_228,In_1633);
or U2321 (N_2321,In_1598,In_473);
nor U2322 (N_2322,In_348,In_1278);
nor U2323 (N_2323,In_1895,In_1923);
nand U2324 (N_2324,In_1195,In_294);
nor U2325 (N_2325,In_862,In_1134);
nor U2326 (N_2326,In_26,In_1203);
and U2327 (N_2327,In_1716,In_1398);
nand U2328 (N_2328,In_782,In_541);
nand U2329 (N_2329,In_807,In_415);
and U2330 (N_2330,In_875,In_54);
and U2331 (N_2331,In_1888,In_261);
nand U2332 (N_2332,In_400,In_472);
and U2333 (N_2333,In_1895,In_1430);
xor U2334 (N_2334,In_263,In_850);
nand U2335 (N_2335,In_1770,In_1147);
nor U2336 (N_2336,In_791,In_891);
and U2337 (N_2337,In_517,In_500);
nand U2338 (N_2338,In_1057,In_452);
or U2339 (N_2339,In_318,In_660);
and U2340 (N_2340,In_1581,In_74);
or U2341 (N_2341,In_499,In_477);
and U2342 (N_2342,In_1345,In_260);
nor U2343 (N_2343,In_1267,In_724);
nor U2344 (N_2344,In_1877,In_1393);
and U2345 (N_2345,In_221,In_398);
and U2346 (N_2346,In_1560,In_630);
or U2347 (N_2347,In_306,In_715);
or U2348 (N_2348,In_1533,In_1222);
nand U2349 (N_2349,In_381,In_1964);
and U2350 (N_2350,In_209,In_331);
or U2351 (N_2351,In_1132,In_1094);
nand U2352 (N_2352,In_1245,In_1284);
nand U2353 (N_2353,In_1689,In_1896);
and U2354 (N_2354,In_1952,In_1770);
and U2355 (N_2355,In_1298,In_409);
nor U2356 (N_2356,In_1171,In_1583);
nor U2357 (N_2357,In_1612,In_1752);
or U2358 (N_2358,In_928,In_208);
nor U2359 (N_2359,In_167,In_850);
or U2360 (N_2360,In_392,In_744);
nor U2361 (N_2361,In_1630,In_1187);
and U2362 (N_2362,In_885,In_332);
nand U2363 (N_2363,In_77,In_750);
nand U2364 (N_2364,In_837,In_226);
and U2365 (N_2365,In_1416,In_519);
xnor U2366 (N_2366,In_620,In_882);
xor U2367 (N_2367,In_570,In_1025);
or U2368 (N_2368,In_790,In_797);
or U2369 (N_2369,In_958,In_1483);
or U2370 (N_2370,In_711,In_1583);
nand U2371 (N_2371,In_1877,In_69);
xor U2372 (N_2372,In_1151,In_859);
nor U2373 (N_2373,In_230,In_591);
and U2374 (N_2374,In_725,In_284);
xnor U2375 (N_2375,In_839,In_1420);
nand U2376 (N_2376,In_1809,In_1402);
nand U2377 (N_2377,In_595,In_696);
nand U2378 (N_2378,In_1739,In_974);
and U2379 (N_2379,In_1473,In_271);
nor U2380 (N_2380,In_1137,In_1671);
nor U2381 (N_2381,In_592,In_753);
nand U2382 (N_2382,In_1137,In_1420);
xnor U2383 (N_2383,In_397,In_993);
or U2384 (N_2384,In_1897,In_250);
nand U2385 (N_2385,In_974,In_1499);
or U2386 (N_2386,In_616,In_1781);
or U2387 (N_2387,In_1482,In_1376);
or U2388 (N_2388,In_1374,In_1348);
nor U2389 (N_2389,In_1729,In_1471);
nor U2390 (N_2390,In_217,In_422);
nand U2391 (N_2391,In_1794,In_1587);
nand U2392 (N_2392,In_1234,In_1324);
xnor U2393 (N_2393,In_441,In_476);
nand U2394 (N_2394,In_381,In_1167);
xnor U2395 (N_2395,In_388,In_1076);
and U2396 (N_2396,In_1205,In_885);
or U2397 (N_2397,In_1318,In_1058);
nand U2398 (N_2398,In_569,In_764);
nor U2399 (N_2399,In_522,In_436);
or U2400 (N_2400,In_879,In_1437);
or U2401 (N_2401,In_1119,In_1107);
nand U2402 (N_2402,In_1269,In_681);
or U2403 (N_2403,In_1484,In_620);
nor U2404 (N_2404,In_1703,In_1217);
and U2405 (N_2405,In_1646,In_627);
or U2406 (N_2406,In_1519,In_895);
nand U2407 (N_2407,In_392,In_105);
or U2408 (N_2408,In_1870,In_507);
or U2409 (N_2409,In_858,In_1373);
xor U2410 (N_2410,In_1,In_908);
and U2411 (N_2411,In_1565,In_171);
or U2412 (N_2412,In_1527,In_673);
or U2413 (N_2413,In_573,In_1851);
nor U2414 (N_2414,In_569,In_24);
and U2415 (N_2415,In_1195,In_434);
or U2416 (N_2416,In_214,In_600);
nor U2417 (N_2417,In_392,In_1581);
nand U2418 (N_2418,In_1514,In_1931);
nand U2419 (N_2419,In_1640,In_329);
xnor U2420 (N_2420,In_107,In_1835);
xnor U2421 (N_2421,In_257,In_1779);
nor U2422 (N_2422,In_334,In_1409);
nor U2423 (N_2423,In_97,In_832);
and U2424 (N_2424,In_1266,In_1349);
or U2425 (N_2425,In_288,In_750);
nor U2426 (N_2426,In_661,In_82);
or U2427 (N_2427,In_1092,In_1954);
and U2428 (N_2428,In_541,In_70);
nor U2429 (N_2429,In_1034,In_1102);
nand U2430 (N_2430,In_1665,In_1909);
and U2431 (N_2431,In_665,In_1614);
or U2432 (N_2432,In_916,In_425);
nand U2433 (N_2433,In_1692,In_426);
xnor U2434 (N_2434,In_1343,In_1010);
and U2435 (N_2435,In_1961,In_146);
nor U2436 (N_2436,In_1035,In_280);
nor U2437 (N_2437,In_1423,In_1140);
nand U2438 (N_2438,In_1907,In_1125);
or U2439 (N_2439,In_1998,In_564);
or U2440 (N_2440,In_499,In_1261);
nand U2441 (N_2441,In_794,In_99);
nand U2442 (N_2442,In_561,In_1624);
nor U2443 (N_2443,In_817,In_293);
and U2444 (N_2444,In_819,In_1384);
nand U2445 (N_2445,In_928,In_1824);
nor U2446 (N_2446,In_1788,In_993);
xnor U2447 (N_2447,In_1307,In_916);
xnor U2448 (N_2448,In_156,In_1739);
nand U2449 (N_2449,In_223,In_1148);
or U2450 (N_2450,In_1267,In_333);
nor U2451 (N_2451,In_801,In_1501);
nand U2452 (N_2452,In_230,In_1377);
or U2453 (N_2453,In_615,In_1698);
and U2454 (N_2454,In_481,In_787);
and U2455 (N_2455,In_1160,In_270);
nor U2456 (N_2456,In_1286,In_1417);
nand U2457 (N_2457,In_709,In_1247);
nand U2458 (N_2458,In_1567,In_729);
nand U2459 (N_2459,In_269,In_1143);
or U2460 (N_2460,In_1467,In_1713);
nor U2461 (N_2461,In_904,In_970);
and U2462 (N_2462,In_345,In_20);
nor U2463 (N_2463,In_789,In_320);
or U2464 (N_2464,In_1877,In_464);
nand U2465 (N_2465,In_1643,In_474);
and U2466 (N_2466,In_1369,In_416);
nand U2467 (N_2467,In_1597,In_323);
or U2468 (N_2468,In_1553,In_868);
and U2469 (N_2469,In_624,In_818);
nor U2470 (N_2470,In_1337,In_367);
or U2471 (N_2471,In_1956,In_1794);
nor U2472 (N_2472,In_1671,In_1067);
nand U2473 (N_2473,In_641,In_1598);
nor U2474 (N_2474,In_286,In_97);
xnor U2475 (N_2475,In_1467,In_752);
nor U2476 (N_2476,In_879,In_1934);
nor U2477 (N_2477,In_148,In_1248);
and U2478 (N_2478,In_1542,In_1802);
and U2479 (N_2479,In_95,In_204);
or U2480 (N_2480,In_1824,In_490);
or U2481 (N_2481,In_1969,In_1698);
nand U2482 (N_2482,In_302,In_349);
and U2483 (N_2483,In_1472,In_402);
nor U2484 (N_2484,In_1955,In_182);
xor U2485 (N_2485,In_135,In_540);
or U2486 (N_2486,In_1135,In_975);
nor U2487 (N_2487,In_1556,In_1634);
nor U2488 (N_2488,In_1323,In_17);
xor U2489 (N_2489,In_1679,In_108);
or U2490 (N_2490,In_1207,In_1741);
nor U2491 (N_2491,In_497,In_542);
or U2492 (N_2492,In_1032,In_1461);
xor U2493 (N_2493,In_1123,In_1115);
nand U2494 (N_2494,In_1275,In_1465);
nand U2495 (N_2495,In_1486,In_1861);
or U2496 (N_2496,In_1213,In_1349);
nand U2497 (N_2497,In_1777,In_180);
xor U2498 (N_2498,In_151,In_1093);
xor U2499 (N_2499,In_28,In_393);
and U2500 (N_2500,In_504,In_502);
nand U2501 (N_2501,In_1460,In_360);
nor U2502 (N_2502,In_50,In_185);
and U2503 (N_2503,In_292,In_1646);
and U2504 (N_2504,In_1253,In_1754);
or U2505 (N_2505,In_47,In_1865);
and U2506 (N_2506,In_393,In_57);
nor U2507 (N_2507,In_231,In_1759);
nand U2508 (N_2508,In_1664,In_1959);
or U2509 (N_2509,In_82,In_1444);
or U2510 (N_2510,In_1157,In_1279);
nor U2511 (N_2511,In_74,In_658);
or U2512 (N_2512,In_1003,In_812);
or U2513 (N_2513,In_717,In_29);
nand U2514 (N_2514,In_1077,In_1518);
and U2515 (N_2515,In_1049,In_461);
and U2516 (N_2516,In_378,In_920);
or U2517 (N_2517,In_275,In_1301);
and U2518 (N_2518,In_1458,In_1418);
nor U2519 (N_2519,In_1299,In_832);
nor U2520 (N_2520,In_1332,In_348);
nor U2521 (N_2521,In_1367,In_1087);
or U2522 (N_2522,In_946,In_336);
and U2523 (N_2523,In_1079,In_1474);
nor U2524 (N_2524,In_189,In_466);
or U2525 (N_2525,In_850,In_892);
and U2526 (N_2526,In_758,In_389);
or U2527 (N_2527,In_1883,In_76);
and U2528 (N_2528,In_1546,In_17);
or U2529 (N_2529,In_1455,In_830);
nand U2530 (N_2530,In_1170,In_522);
and U2531 (N_2531,In_1973,In_1181);
or U2532 (N_2532,In_470,In_1830);
nand U2533 (N_2533,In_508,In_1278);
and U2534 (N_2534,In_396,In_698);
nand U2535 (N_2535,In_1342,In_1212);
or U2536 (N_2536,In_942,In_1602);
nand U2537 (N_2537,In_765,In_1525);
nand U2538 (N_2538,In_217,In_522);
nand U2539 (N_2539,In_193,In_214);
nand U2540 (N_2540,In_1876,In_1341);
nand U2541 (N_2541,In_1131,In_1502);
and U2542 (N_2542,In_792,In_23);
and U2543 (N_2543,In_212,In_996);
nor U2544 (N_2544,In_24,In_220);
nand U2545 (N_2545,In_951,In_1008);
nor U2546 (N_2546,In_847,In_1509);
and U2547 (N_2547,In_1458,In_1019);
nand U2548 (N_2548,In_101,In_203);
nand U2549 (N_2549,In_256,In_103);
xnor U2550 (N_2550,In_1303,In_748);
nor U2551 (N_2551,In_1622,In_1174);
nor U2552 (N_2552,In_187,In_332);
and U2553 (N_2553,In_1513,In_801);
or U2554 (N_2554,In_583,In_849);
xor U2555 (N_2555,In_42,In_650);
nand U2556 (N_2556,In_581,In_1523);
nor U2557 (N_2557,In_557,In_1806);
and U2558 (N_2558,In_1404,In_1626);
xnor U2559 (N_2559,In_934,In_746);
or U2560 (N_2560,In_1479,In_38);
and U2561 (N_2561,In_955,In_120);
xor U2562 (N_2562,In_592,In_661);
nor U2563 (N_2563,In_1668,In_1115);
or U2564 (N_2564,In_132,In_1187);
nand U2565 (N_2565,In_1749,In_374);
or U2566 (N_2566,In_328,In_1598);
nor U2567 (N_2567,In_835,In_158);
nor U2568 (N_2568,In_514,In_824);
or U2569 (N_2569,In_1509,In_1134);
nand U2570 (N_2570,In_1707,In_80);
xnor U2571 (N_2571,In_961,In_776);
nand U2572 (N_2572,In_769,In_1279);
and U2573 (N_2573,In_877,In_219);
nand U2574 (N_2574,In_386,In_1575);
nor U2575 (N_2575,In_695,In_764);
nand U2576 (N_2576,In_1090,In_1360);
xnor U2577 (N_2577,In_1107,In_1718);
and U2578 (N_2578,In_1445,In_1894);
or U2579 (N_2579,In_963,In_1728);
or U2580 (N_2580,In_679,In_292);
xor U2581 (N_2581,In_1858,In_1392);
nor U2582 (N_2582,In_1098,In_1918);
nand U2583 (N_2583,In_1836,In_1401);
nor U2584 (N_2584,In_1093,In_433);
nor U2585 (N_2585,In_1025,In_497);
nor U2586 (N_2586,In_572,In_966);
nor U2587 (N_2587,In_1414,In_1772);
nand U2588 (N_2588,In_979,In_1805);
nand U2589 (N_2589,In_84,In_1608);
or U2590 (N_2590,In_1432,In_1581);
or U2591 (N_2591,In_548,In_520);
and U2592 (N_2592,In_702,In_1696);
nor U2593 (N_2593,In_439,In_768);
nand U2594 (N_2594,In_513,In_1928);
and U2595 (N_2595,In_395,In_245);
nor U2596 (N_2596,In_1537,In_1386);
xnor U2597 (N_2597,In_381,In_339);
nor U2598 (N_2598,In_1721,In_1223);
or U2599 (N_2599,In_1856,In_1787);
nand U2600 (N_2600,In_1184,In_1043);
and U2601 (N_2601,In_1063,In_480);
or U2602 (N_2602,In_221,In_387);
nand U2603 (N_2603,In_1688,In_1519);
or U2604 (N_2604,In_1819,In_1556);
nand U2605 (N_2605,In_888,In_1261);
and U2606 (N_2606,In_1077,In_653);
nand U2607 (N_2607,In_715,In_1057);
nor U2608 (N_2608,In_398,In_1619);
nor U2609 (N_2609,In_1316,In_1566);
nand U2610 (N_2610,In_1045,In_1712);
xor U2611 (N_2611,In_1385,In_1837);
nand U2612 (N_2612,In_953,In_259);
nand U2613 (N_2613,In_464,In_872);
and U2614 (N_2614,In_975,In_400);
or U2615 (N_2615,In_700,In_617);
or U2616 (N_2616,In_577,In_1415);
nand U2617 (N_2617,In_1247,In_656);
nor U2618 (N_2618,In_362,In_1485);
nand U2619 (N_2619,In_150,In_1);
nand U2620 (N_2620,In_1358,In_197);
nand U2621 (N_2621,In_639,In_382);
xnor U2622 (N_2622,In_792,In_1456);
nand U2623 (N_2623,In_994,In_648);
or U2624 (N_2624,In_88,In_1034);
and U2625 (N_2625,In_1176,In_1158);
and U2626 (N_2626,In_656,In_257);
and U2627 (N_2627,In_1428,In_1576);
or U2628 (N_2628,In_1613,In_599);
xnor U2629 (N_2629,In_1823,In_769);
nor U2630 (N_2630,In_1466,In_87);
or U2631 (N_2631,In_868,In_557);
nor U2632 (N_2632,In_329,In_1601);
or U2633 (N_2633,In_1628,In_206);
nand U2634 (N_2634,In_433,In_1078);
nor U2635 (N_2635,In_388,In_944);
or U2636 (N_2636,In_590,In_661);
nand U2637 (N_2637,In_935,In_730);
or U2638 (N_2638,In_143,In_1849);
nor U2639 (N_2639,In_921,In_314);
nand U2640 (N_2640,In_1775,In_1315);
nor U2641 (N_2641,In_1523,In_876);
nand U2642 (N_2642,In_1036,In_822);
or U2643 (N_2643,In_1101,In_644);
xor U2644 (N_2644,In_1850,In_953);
nor U2645 (N_2645,In_1129,In_1204);
nand U2646 (N_2646,In_82,In_1957);
and U2647 (N_2647,In_1799,In_907);
and U2648 (N_2648,In_1431,In_475);
and U2649 (N_2649,In_410,In_626);
nand U2650 (N_2650,In_821,In_423);
and U2651 (N_2651,In_978,In_1899);
xor U2652 (N_2652,In_1785,In_1086);
or U2653 (N_2653,In_909,In_62);
and U2654 (N_2654,In_1570,In_1788);
nand U2655 (N_2655,In_599,In_296);
nor U2656 (N_2656,In_1337,In_215);
nand U2657 (N_2657,In_904,In_757);
xnor U2658 (N_2658,In_34,In_871);
or U2659 (N_2659,In_618,In_161);
and U2660 (N_2660,In_1902,In_1736);
nand U2661 (N_2661,In_916,In_1580);
nor U2662 (N_2662,In_545,In_1452);
and U2663 (N_2663,In_501,In_1);
or U2664 (N_2664,In_218,In_1739);
nand U2665 (N_2665,In_877,In_151);
and U2666 (N_2666,In_109,In_1929);
or U2667 (N_2667,In_1759,In_1143);
xor U2668 (N_2668,In_1353,In_1400);
nor U2669 (N_2669,In_204,In_385);
and U2670 (N_2670,In_621,In_694);
and U2671 (N_2671,In_799,In_1970);
nor U2672 (N_2672,In_1940,In_1553);
nor U2673 (N_2673,In_1988,In_1807);
nand U2674 (N_2674,In_1281,In_550);
nand U2675 (N_2675,In_1901,In_259);
nand U2676 (N_2676,In_316,In_297);
nand U2677 (N_2677,In_667,In_953);
nand U2678 (N_2678,In_1704,In_575);
nand U2679 (N_2679,In_1376,In_240);
nand U2680 (N_2680,In_1135,In_1093);
xor U2681 (N_2681,In_489,In_656);
nor U2682 (N_2682,In_176,In_449);
and U2683 (N_2683,In_603,In_1613);
nand U2684 (N_2684,In_906,In_1762);
or U2685 (N_2685,In_437,In_444);
nand U2686 (N_2686,In_611,In_6);
xor U2687 (N_2687,In_956,In_403);
and U2688 (N_2688,In_732,In_1282);
and U2689 (N_2689,In_1704,In_1959);
or U2690 (N_2690,In_692,In_516);
or U2691 (N_2691,In_1907,In_1104);
nand U2692 (N_2692,In_776,In_1315);
nor U2693 (N_2693,In_1009,In_361);
nor U2694 (N_2694,In_119,In_1619);
nor U2695 (N_2695,In_1366,In_422);
and U2696 (N_2696,In_725,In_1951);
and U2697 (N_2697,In_1072,In_1175);
nand U2698 (N_2698,In_1841,In_688);
xor U2699 (N_2699,In_1224,In_1853);
and U2700 (N_2700,In_1533,In_253);
nand U2701 (N_2701,In_475,In_616);
nor U2702 (N_2702,In_1865,In_775);
and U2703 (N_2703,In_52,In_220);
and U2704 (N_2704,In_1015,In_1344);
nand U2705 (N_2705,In_1552,In_417);
and U2706 (N_2706,In_11,In_1255);
and U2707 (N_2707,In_1975,In_1463);
and U2708 (N_2708,In_723,In_56);
nor U2709 (N_2709,In_1981,In_1918);
xor U2710 (N_2710,In_1067,In_170);
or U2711 (N_2711,In_573,In_1804);
nor U2712 (N_2712,In_1117,In_736);
and U2713 (N_2713,In_541,In_1392);
nand U2714 (N_2714,In_866,In_1710);
or U2715 (N_2715,In_1707,In_758);
nor U2716 (N_2716,In_1475,In_1385);
and U2717 (N_2717,In_1560,In_1229);
nor U2718 (N_2718,In_747,In_1134);
nor U2719 (N_2719,In_1038,In_1106);
nand U2720 (N_2720,In_71,In_1160);
nor U2721 (N_2721,In_714,In_1938);
and U2722 (N_2722,In_169,In_467);
and U2723 (N_2723,In_114,In_1557);
nand U2724 (N_2724,In_683,In_1115);
and U2725 (N_2725,In_252,In_1074);
or U2726 (N_2726,In_761,In_231);
and U2727 (N_2727,In_312,In_153);
or U2728 (N_2728,In_237,In_760);
and U2729 (N_2729,In_869,In_994);
and U2730 (N_2730,In_376,In_565);
nor U2731 (N_2731,In_862,In_1124);
or U2732 (N_2732,In_73,In_103);
xnor U2733 (N_2733,In_1536,In_1803);
and U2734 (N_2734,In_1823,In_1350);
or U2735 (N_2735,In_816,In_695);
nor U2736 (N_2736,In_196,In_1902);
and U2737 (N_2737,In_1534,In_899);
xnor U2738 (N_2738,In_462,In_1677);
nand U2739 (N_2739,In_1027,In_1512);
nor U2740 (N_2740,In_1187,In_856);
nand U2741 (N_2741,In_1573,In_1443);
nor U2742 (N_2742,In_484,In_1568);
nor U2743 (N_2743,In_1969,In_64);
or U2744 (N_2744,In_371,In_1332);
and U2745 (N_2745,In_431,In_1503);
nand U2746 (N_2746,In_1721,In_72);
xor U2747 (N_2747,In_782,In_219);
nand U2748 (N_2748,In_800,In_1009);
or U2749 (N_2749,In_338,In_128);
and U2750 (N_2750,In_135,In_451);
nand U2751 (N_2751,In_1998,In_179);
xor U2752 (N_2752,In_916,In_1741);
and U2753 (N_2753,In_1790,In_381);
or U2754 (N_2754,In_1603,In_1998);
nand U2755 (N_2755,In_510,In_1805);
xnor U2756 (N_2756,In_177,In_293);
nand U2757 (N_2757,In_1283,In_770);
nor U2758 (N_2758,In_1276,In_541);
nand U2759 (N_2759,In_1659,In_190);
nand U2760 (N_2760,In_1820,In_1899);
nor U2761 (N_2761,In_1480,In_1183);
or U2762 (N_2762,In_1432,In_182);
or U2763 (N_2763,In_862,In_815);
or U2764 (N_2764,In_1741,In_1620);
nor U2765 (N_2765,In_18,In_1241);
and U2766 (N_2766,In_532,In_1178);
and U2767 (N_2767,In_1291,In_214);
and U2768 (N_2768,In_1750,In_615);
or U2769 (N_2769,In_1456,In_591);
and U2770 (N_2770,In_621,In_1560);
nor U2771 (N_2771,In_915,In_158);
nor U2772 (N_2772,In_1709,In_506);
nand U2773 (N_2773,In_502,In_1136);
and U2774 (N_2774,In_1816,In_1150);
and U2775 (N_2775,In_1795,In_437);
and U2776 (N_2776,In_707,In_698);
and U2777 (N_2777,In_1383,In_666);
nor U2778 (N_2778,In_921,In_875);
and U2779 (N_2779,In_1252,In_1985);
and U2780 (N_2780,In_1180,In_476);
and U2781 (N_2781,In_285,In_163);
or U2782 (N_2782,In_831,In_1180);
or U2783 (N_2783,In_1725,In_1166);
nand U2784 (N_2784,In_1412,In_671);
and U2785 (N_2785,In_2,In_1052);
xnor U2786 (N_2786,In_574,In_1066);
nor U2787 (N_2787,In_1877,In_1167);
nand U2788 (N_2788,In_185,In_659);
and U2789 (N_2789,In_1390,In_123);
and U2790 (N_2790,In_587,In_299);
nor U2791 (N_2791,In_1610,In_1103);
or U2792 (N_2792,In_1238,In_1979);
or U2793 (N_2793,In_902,In_1185);
nand U2794 (N_2794,In_1104,In_1866);
nand U2795 (N_2795,In_1558,In_320);
and U2796 (N_2796,In_584,In_1245);
or U2797 (N_2797,In_131,In_138);
nor U2798 (N_2798,In_1079,In_1473);
or U2799 (N_2799,In_1086,In_1230);
or U2800 (N_2800,In_1991,In_529);
and U2801 (N_2801,In_1539,In_1676);
nor U2802 (N_2802,In_1616,In_1815);
nor U2803 (N_2803,In_1798,In_405);
nand U2804 (N_2804,In_1462,In_815);
nor U2805 (N_2805,In_56,In_100);
or U2806 (N_2806,In_1302,In_37);
nor U2807 (N_2807,In_1679,In_566);
or U2808 (N_2808,In_1292,In_1908);
xnor U2809 (N_2809,In_349,In_175);
nand U2810 (N_2810,In_1172,In_983);
and U2811 (N_2811,In_1018,In_584);
and U2812 (N_2812,In_1890,In_421);
and U2813 (N_2813,In_1328,In_1889);
and U2814 (N_2814,In_390,In_989);
nand U2815 (N_2815,In_563,In_167);
nand U2816 (N_2816,In_246,In_1988);
nor U2817 (N_2817,In_1893,In_1175);
nand U2818 (N_2818,In_704,In_1541);
or U2819 (N_2819,In_476,In_1608);
nor U2820 (N_2820,In_1535,In_565);
and U2821 (N_2821,In_1201,In_1191);
or U2822 (N_2822,In_1655,In_1699);
nor U2823 (N_2823,In_733,In_1296);
or U2824 (N_2824,In_1775,In_559);
nor U2825 (N_2825,In_702,In_1999);
or U2826 (N_2826,In_196,In_249);
and U2827 (N_2827,In_1282,In_865);
and U2828 (N_2828,In_151,In_840);
nand U2829 (N_2829,In_1320,In_266);
or U2830 (N_2830,In_1201,In_1940);
nand U2831 (N_2831,In_1663,In_895);
nor U2832 (N_2832,In_1240,In_1028);
and U2833 (N_2833,In_1640,In_344);
xnor U2834 (N_2834,In_336,In_1431);
or U2835 (N_2835,In_264,In_599);
xnor U2836 (N_2836,In_557,In_553);
nand U2837 (N_2837,In_199,In_1520);
and U2838 (N_2838,In_1881,In_866);
or U2839 (N_2839,In_1057,In_1322);
nand U2840 (N_2840,In_1080,In_990);
nand U2841 (N_2841,In_1509,In_1963);
nor U2842 (N_2842,In_1784,In_1238);
or U2843 (N_2843,In_1926,In_838);
or U2844 (N_2844,In_939,In_325);
nand U2845 (N_2845,In_1238,In_179);
or U2846 (N_2846,In_1489,In_779);
and U2847 (N_2847,In_1783,In_1893);
nand U2848 (N_2848,In_1936,In_1512);
nor U2849 (N_2849,In_762,In_1222);
nor U2850 (N_2850,In_1051,In_1748);
and U2851 (N_2851,In_1002,In_38);
xor U2852 (N_2852,In_1705,In_142);
nor U2853 (N_2853,In_361,In_919);
and U2854 (N_2854,In_703,In_651);
or U2855 (N_2855,In_1698,In_1363);
nor U2856 (N_2856,In_1193,In_212);
xnor U2857 (N_2857,In_781,In_761);
xor U2858 (N_2858,In_1573,In_616);
nor U2859 (N_2859,In_1688,In_892);
xnor U2860 (N_2860,In_1728,In_745);
or U2861 (N_2861,In_642,In_1446);
nor U2862 (N_2862,In_1375,In_580);
nand U2863 (N_2863,In_866,In_1456);
or U2864 (N_2864,In_1241,In_1057);
nor U2865 (N_2865,In_693,In_712);
or U2866 (N_2866,In_1996,In_1525);
nand U2867 (N_2867,In_700,In_550);
or U2868 (N_2868,In_109,In_857);
nand U2869 (N_2869,In_752,In_281);
nand U2870 (N_2870,In_1203,In_1608);
and U2871 (N_2871,In_852,In_516);
nand U2872 (N_2872,In_175,In_1004);
nor U2873 (N_2873,In_499,In_850);
nand U2874 (N_2874,In_1715,In_1176);
or U2875 (N_2875,In_1006,In_1);
nor U2876 (N_2876,In_1748,In_947);
and U2877 (N_2877,In_146,In_1245);
nand U2878 (N_2878,In_1189,In_1603);
and U2879 (N_2879,In_1277,In_1593);
xor U2880 (N_2880,In_1426,In_1522);
nor U2881 (N_2881,In_881,In_506);
nand U2882 (N_2882,In_287,In_1877);
nor U2883 (N_2883,In_11,In_1925);
xnor U2884 (N_2884,In_120,In_1443);
and U2885 (N_2885,In_837,In_534);
nand U2886 (N_2886,In_969,In_772);
and U2887 (N_2887,In_822,In_486);
nand U2888 (N_2888,In_364,In_1763);
xor U2889 (N_2889,In_3,In_511);
nand U2890 (N_2890,In_569,In_997);
nand U2891 (N_2891,In_985,In_249);
nand U2892 (N_2892,In_1100,In_502);
nor U2893 (N_2893,In_1592,In_448);
nand U2894 (N_2894,In_1818,In_1967);
or U2895 (N_2895,In_521,In_379);
nand U2896 (N_2896,In_1175,In_304);
or U2897 (N_2897,In_1416,In_1569);
nor U2898 (N_2898,In_186,In_374);
and U2899 (N_2899,In_1414,In_255);
and U2900 (N_2900,In_249,In_869);
or U2901 (N_2901,In_1938,In_894);
or U2902 (N_2902,In_661,In_371);
nor U2903 (N_2903,In_1647,In_79);
and U2904 (N_2904,In_1671,In_649);
or U2905 (N_2905,In_1542,In_739);
nor U2906 (N_2906,In_429,In_1877);
nand U2907 (N_2907,In_1333,In_733);
or U2908 (N_2908,In_399,In_1123);
and U2909 (N_2909,In_876,In_1858);
nand U2910 (N_2910,In_1865,In_551);
or U2911 (N_2911,In_1218,In_33);
or U2912 (N_2912,In_845,In_1823);
xnor U2913 (N_2913,In_57,In_1374);
nand U2914 (N_2914,In_715,In_883);
or U2915 (N_2915,In_809,In_1113);
nor U2916 (N_2916,In_1172,In_1155);
nor U2917 (N_2917,In_1628,In_1667);
and U2918 (N_2918,In_272,In_435);
nor U2919 (N_2919,In_239,In_99);
xnor U2920 (N_2920,In_1910,In_1241);
and U2921 (N_2921,In_312,In_1842);
or U2922 (N_2922,In_369,In_1733);
and U2923 (N_2923,In_1339,In_1034);
and U2924 (N_2924,In_1710,In_1484);
nand U2925 (N_2925,In_1458,In_738);
nand U2926 (N_2926,In_1410,In_1696);
nor U2927 (N_2927,In_598,In_1565);
xor U2928 (N_2928,In_1671,In_1894);
nor U2929 (N_2929,In_1241,In_1783);
and U2930 (N_2930,In_1828,In_881);
nor U2931 (N_2931,In_874,In_1173);
and U2932 (N_2932,In_1709,In_1084);
and U2933 (N_2933,In_940,In_1985);
xnor U2934 (N_2934,In_1510,In_619);
nor U2935 (N_2935,In_150,In_1588);
and U2936 (N_2936,In_877,In_1700);
or U2937 (N_2937,In_978,In_68);
xnor U2938 (N_2938,In_909,In_567);
nor U2939 (N_2939,In_1907,In_779);
xor U2940 (N_2940,In_440,In_1573);
nor U2941 (N_2941,In_83,In_1803);
or U2942 (N_2942,In_739,In_1120);
nand U2943 (N_2943,In_1263,In_12);
xor U2944 (N_2944,In_1759,In_743);
or U2945 (N_2945,In_295,In_665);
and U2946 (N_2946,In_1138,In_453);
or U2947 (N_2947,In_1573,In_518);
nor U2948 (N_2948,In_690,In_778);
and U2949 (N_2949,In_1561,In_246);
or U2950 (N_2950,In_1258,In_20);
nand U2951 (N_2951,In_1028,In_1764);
and U2952 (N_2952,In_1018,In_509);
and U2953 (N_2953,In_815,In_206);
xor U2954 (N_2954,In_77,In_217);
nand U2955 (N_2955,In_378,In_256);
xor U2956 (N_2956,In_708,In_1604);
and U2957 (N_2957,In_296,In_1781);
nor U2958 (N_2958,In_126,In_432);
nand U2959 (N_2959,In_1074,In_1127);
xnor U2960 (N_2960,In_1171,In_210);
nand U2961 (N_2961,In_1219,In_1606);
nor U2962 (N_2962,In_142,In_400);
or U2963 (N_2963,In_1216,In_1662);
or U2964 (N_2964,In_143,In_2);
and U2965 (N_2965,In_1388,In_1485);
nand U2966 (N_2966,In_171,In_243);
nand U2967 (N_2967,In_1672,In_309);
xor U2968 (N_2968,In_1631,In_1572);
and U2969 (N_2969,In_1099,In_1381);
nor U2970 (N_2970,In_319,In_527);
or U2971 (N_2971,In_417,In_264);
and U2972 (N_2972,In_876,In_437);
and U2973 (N_2973,In_40,In_30);
nor U2974 (N_2974,In_490,In_1689);
nand U2975 (N_2975,In_143,In_1398);
xor U2976 (N_2976,In_207,In_1864);
nand U2977 (N_2977,In_1050,In_660);
and U2978 (N_2978,In_516,In_1878);
nand U2979 (N_2979,In_754,In_93);
and U2980 (N_2980,In_1292,In_1447);
or U2981 (N_2981,In_1812,In_1317);
nor U2982 (N_2982,In_992,In_374);
and U2983 (N_2983,In_1832,In_387);
and U2984 (N_2984,In_675,In_1471);
or U2985 (N_2985,In_118,In_303);
nor U2986 (N_2986,In_1422,In_491);
nand U2987 (N_2987,In_220,In_393);
nand U2988 (N_2988,In_242,In_1383);
and U2989 (N_2989,In_1770,In_710);
and U2990 (N_2990,In_1781,In_880);
nand U2991 (N_2991,In_250,In_366);
nor U2992 (N_2992,In_1352,In_1894);
xnor U2993 (N_2993,In_1865,In_1334);
or U2994 (N_2994,In_576,In_1383);
nor U2995 (N_2995,In_934,In_1118);
nand U2996 (N_2996,In_854,In_435);
nor U2997 (N_2997,In_1747,In_168);
or U2998 (N_2998,In_1260,In_1571);
and U2999 (N_2999,In_1107,In_1345);
and U3000 (N_3000,In_1447,In_621);
nor U3001 (N_3001,In_1983,In_1051);
and U3002 (N_3002,In_989,In_597);
nand U3003 (N_3003,In_91,In_1374);
or U3004 (N_3004,In_551,In_1222);
or U3005 (N_3005,In_682,In_726);
nor U3006 (N_3006,In_165,In_371);
nor U3007 (N_3007,In_833,In_1930);
xor U3008 (N_3008,In_1398,In_556);
and U3009 (N_3009,In_455,In_188);
nand U3010 (N_3010,In_1208,In_1883);
or U3011 (N_3011,In_290,In_333);
and U3012 (N_3012,In_1415,In_876);
xor U3013 (N_3013,In_439,In_1398);
nor U3014 (N_3014,In_510,In_1181);
and U3015 (N_3015,In_962,In_1053);
nor U3016 (N_3016,In_1089,In_736);
xor U3017 (N_3017,In_1039,In_282);
or U3018 (N_3018,In_617,In_374);
nor U3019 (N_3019,In_1617,In_1717);
nand U3020 (N_3020,In_1000,In_87);
nand U3021 (N_3021,In_398,In_1880);
xnor U3022 (N_3022,In_1846,In_314);
or U3023 (N_3023,In_1260,In_407);
and U3024 (N_3024,In_974,In_1782);
xor U3025 (N_3025,In_370,In_503);
xnor U3026 (N_3026,In_1715,In_1885);
or U3027 (N_3027,In_246,In_238);
nand U3028 (N_3028,In_499,In_1007);
and U3029 (N_3029,In_1022,In_984);
nand U3030 (N_3030,In_1898,In_380);
nand U3031 (N_3031,In_1921,In_1876);
xor U3032 (N_3032,In_676,In_1102);
nor U3033 (N_3033,In_178,In_552);
nand U3034 (N_3034,In_201,In_1525);
or U3035 (N_3035,In_870,In_888);
nor U3036 (N_3036,In_811,In_786);
and U3037 (N_3037,In_1043,In_948);
nand U3038 (N_3038,In_475,In_467);
and U3039 (N_3039,In_1971,In_1174);
or U3040 (N_3040,In_1106,In_1757);
and U3041 (N_3041,In_1545,In_930);
and U3042 (N_3042,In_171,In_1944);
nor U3043 (N_3043,In_317,In_574);
nor U3044 (N_3044,In_426,In_1320);
or U3045 (N_3045,In_787,In_1752);
and U3046 (N_3046,In_465,In_1359);
nor U3047 (N_3047,In_595,In_731);
nand U3048 (N_3048,In_329,In_1489);
or U3049 (N_3049,In_1764,In_1050);
or U3050 (N_3050,In_591,In_17);
or U3051 (N_3051,In_395,In_1651);
nor U3052 (N_3052,In_1806,In_1411);
and U3053 (N_3053,In_282,In_215);
and U3054 (N_3054,In_1673,In_1123);
xor U3055 (N_3055,In_1776,In_789);
nor U3056 (N_3056,In_967,In_941);
and U3057 (N_3057,In_1965,In_968);
nor U3058 (N_3058,In_276,In_1989);
nor U3059 (N_3059,In_1585,In_1736);
or U3060 (N_3060,In_502,In_773);
and U3061 (N_3061,In_460,In_1699);
and U3062 (N_3062,In_1357,In_1004);
nand U3063 (N_3063,In_117,In_1220);
nand U3064 (N_3064,In_56,In_756);
nand U3065 (N_3065,In_1995,In_1322);
nand U3066 (N_3066,In_835,In_1569);
and U3067 (N_3067,In_95,In_504);
and U3068 (N_3068,In_848,In_1372);
nor U3069 (N_3069,In_418,In_1104);
nor U3070 (N_3070,In_174,In_1446);
nor U3071 (N_3071,In_397,In_1231);
nor U3072 (N_3072,In_1992,In_1733);
nor U3073 (N_3073,In_541,In_1807);
or U3074 (N_3074,In_1997,In_994);
nor U3075 (N_3075,In_1315,In_1392);
nor U3076 (N_3076,In_1523,In_1475);
nand U3077 (N_3077,In_45,In_1103);
or U3078 (N_3078,In_1238,In_1838);
and U3079 (N_3079,In_1817,In_1931);
or U3080 (N_3080,In_349,In_255);
and U3081 (N_3081,In_309,In_1035);
or U3082 (N_3082,In_1318,In_1869);
and U3083 (N_3083,In_1364,In_791);
nand U3084 (N_3084,In_85,In_118);
or U3085 (N_3085,In_99,In_1542);
nor U3086 (N_3086,In_167,In_1452);
and U3087 (N_3087,In_332,In_799);
xor U3088 (N_3088,In_243,In_1736);
nand U3089 (N_3089,In_129,In_1621);
nor U3090 (N_3090,In_1784,In_607);
xnor U3091 (N_3091,In_1860,In_759);
nand U3092 (N_3092,In_890,In_1552);
nor U3093 (N_3093,In_860,In_748);
nand U3094 (N_3094,In_1726,In_683);
and U3095 (N_3095,In_1045,In_1350);
nand U3096 (N_3096,In_1118,In_45);
nor U3097 (N_3097,In_1161,In_1430);
xor U3098 (N_3098,In_1668,In_872);
and U3099 (N_3099,In_191,In_1605);
or U3100 (N_3100,In_974,In_1312);
or U3101 (N_3101,In_1344,In_1103);
and U3102 (N_3102,In_1333,In_538);
or U3103 (N_3103,In_839,In_703);
nor U3104 (N_3104,In_750,In_301);
nor U3105 (N_3105,In_142,In_1309);
or U3106 (N_3106,In_21,In_972);
and U3107 (N_3107,In_1893,In_1872);
and U3108 (N_3108,In_149,In_768);
or U3109 (N_3109,In_1512,In_1323);
nor U3110 (N_3110,In_1653,In_210);
nor U3111 (N_3111,In_327,In_1837);
nand U3112 (N_3112,In_87,In_846);
nor U3113 (N_3113,In_1605,In_354);
nor U3114 (N_3114,In_626,In_1002);
xor U3115 (N_3115,In_998,In_586);
nor U3116 (N_3116,In_124,In_456);
and U3117 (N_3117,In_152,In_36);
xnor U3118 (N_3118,In_1283,In_971);
nor U3119 (N_3119,In_1324,In_214);
nand U3120 (N_3120,In_551,In_1551);
or U3121 (N_3121,In_639,In_456);
xnor U3122 (N_3122,In_1996,In_1547);
xnor U3123 (N_3123,In_910,In_1330);
nand U3124 (N_3124,In_1819,In_1844);
nor U3125 (N_3125,In_1057,In_1829);
nand U3126 (N_3126,In_1647,In_1306);
nand U3127 (N_3127,In_826,In_1640);
nand U3128 (N_3128,In_663,In_1375);
nand U3129 (N_3129,In_675,In_140);
xor U3130 (N_3130,In_248,In_200);
nor U3131 (N_3131,In_1023,In_1030);
and U3132 (N_3132,In_736,In_1220);
nand U3133 (N_3133,In_175,In_705);
xor U3134 (N_3134,In_614,In_1511);
nor U3135 (N_3135,In_663,In_87);
or U3136 (N_3136,In_1883,In_27);
nand U3137 (N_3137,In_1458,In_1807);
or U3138 (N_3138,In_1494,In_539);
nand U3139 (N_3139,In_834,In_550);
or U3140 (N_3140,In_1442,In_326);
nor U3141 (N_3141,In_1826,In_1311);
and U3142 (N_3142,In_1161,In_72);
nor U3143 (N_3143,In_95,In_1648);
nand U3144 (N_3144,In_1519,In_1193);
or U3145 (N_3145,In_1887,In_1567);
nand U3146 (N_3146,In_139,In_76);
nor U3147 (N_3147,In_310,In_797);
nor U3148 (N_3148,In_1499,In_1666);
nor U3149 (N_3149,In_1843,In_1425);
or U3150 (N_3150,In_364,In_123);
nand U3151 (N_3151,In_500,In_580);
and U3152 (N_3152,In_678,In_409);
or U3153 (N_3153,In_1404,In_1530);
and U3154 (N_3154,In_366,In_428);
nand U3155 (N_3155,In_73,In_1855);
or U3156 (N_3156,In_599,In_544);
or U3157 (N_3157,In_999,In_1322);
or U3158 (N_3158,In_696,In_363);
and U3159 (N_3159,In_71,In_1139);
nand U3160 (N_3160,In_522,In_793);
nor U3161 (N_3161,In_366,In_388);
nand U3162 (N_3162,In_1313,In_744);
and U3163 (N_3163,In_1526,In_1649);
or U3164 (N_3164,In_353,In_233);
nand U3165 (N_3165,In_593,In_1855);
nand U3166 (N_3166,In_414,In_872);
or U3167 (N_3167,In_1384,In_1672);
nand U3168 (N_3168,In_1056,In_1687);
nand U3169 (N_3169,In_501,In_1470);
and U3170 (N_3170,In_1347,In_1727);
nand U3171 (N_3171,In_1398,In_1211);
or U3172 (N_3172,In_1433,In_1522);
nor U3173 (N_3173,In_1446,In_1651);
or U3174 (N_3174,In_1899,In_1831);
or U3175 (N_3175,In_1903,In_1831);
nand U3176 (N_3176,In_1689,In_1800);
or U3177 (N_3177,In_371,In_1536);
nor U3178 (N_3178,In_1644,In_142);
nor U3179 (N_3179,In_1430,In_1168);
or U3180 (N_3180,In_1468,In_765);
or U3181 (N_3181,In_236,In_1532);
nor U3182 (N_3182,In_1451,In_1727);
nand U3183 (N_3183,In_368,In_1893);
nor U3184 (N_3184,In_1193,In_1453);
nor U3185 (N_3185,In_1863,In_344);
and U3186 (N_3186,In_81,In_1810);
or U3187 (N_3187,In_837,In_669);
or U3188 (N_3188,In_647,In_930);
nor U3189 (N_3189,In_1061,In_1562);
nand U3190 (N_3190,In_1348,In_1858);
nor U3191 (N_3191,In_1986,In_427);
and U3192 (N_3192,In_74,In_138);
nor U3193 (N_3193,In_754,In_1391);
nand U3194 (N_3194,In_1358,In_436);
or U3195 (N_3195,In_527,In_58);
nor U3196 (N_3196,In_1290,In_1849);
and U3197 (N_3197,In_829,In_1169);
xor U3198 (N_3198,In_891,In_178);
xor U3199 (N_3199,In_1999,In_491);
xor U3200 (N_3200,In_1759,In_1370);
and U3201 (N_3201,In_1246,In_1353);
nand U3202 (N_3202,In_161,In_824);
xnor U3203 (N_3203,In_71,In_1780);
or U3204 (N_3204,In_613,In_1995);
nand U3205 (N_3205,In_34,In_1152);
or U3206 (N_3206,In_1817,In_1256);
nor U3207 (N_3207,In_1329,In_157);
nor U3208 (N_3208,In_599,In_503);
and U3209 (N_3209,In_574,In_802);
nor U3210 (N_3210,In_1231,In_876);
or U3211 (N_3211,In_1324,In_785);
and U3212 (N_3212,In_1662,In_1158);
nor U3213 (N_3213,In_1029,In_1686);
nor U3214 (N_3214,In_867,In_1536);
xor U3215 (N_3215,In_1571,In_818);
and U3216 (N_3216,In_502,In_91);
nand U3217 (N_3217,In_733,In_930);
and U3218 (N_3218,In_937,In_66);
or U3219 (N_3219,In_1259,In_714);
or U3220 (N_3220,In_666,In_371);
xor U3221 (N_3221,In_1229,In_1523);
nand U3222 (N_3222,In_841,In_469);
nor U3223 (N_3223,In_54,In_1422);
or U3224 (N_3224,In_1895,In_500);
nor U3225 (N_3225,In_1379,In_1462);
or U3226 (N_3226,In_1778,In_1840);
or U3227 (N_3227,In_236,In_1731);
or U3228 (N_3228,In_1954,In_1231);
or U3229 (N_3229,In_1081,In_855);
nand U3230 (N_3230,In_188,In_1521);
and U3231 (N_3231,In_1540,In_821);
xor U3232 (N_3232,In_916,In_1886);
or U3233 (N_3233,In_609,In_508);
nor U3234 (N_3234,In_293,In_1099);
and U3235 (N_3235,In_1500,In_33);
or U3236 (N_3236,In_660,In_1149);
nor U3237 (N_3237,In_206,In_1677);
and U3238 (N_3238,In_503,In_1669);
nor U3239 (N_3239,In_1078,In_1395);
nor U3240 (N_3240,In_932,In_687);
nor U3241 (N_3241,In_1476,In_1181);
nand U3242 (N_3242,In_1023,In_1223);
or U3243 (N_3243,In_1648,In_68);
and U3244 (N_3244,In_1965,In_1042);
nand U3245 (N_3245,In_1225,In_1370);
or U3246 (N_3246,In_499,In_684);
or U3247 (N_3247,In_518,In_746);
xnor U3248 (N_3248,In_1040,In_1407);
and U3249 (N_3249,In_464,In_793);
nor U3250 (N_3250,In_1637,In_1410);
xnor U3251 (N_3251,In_881,In_1270);
nor U3252 (N_3252,In_1347,In_1467);
or U3253 (N_3253,In_834,In_532);
nand U3254 (N_3254,In_1767,In_1068);
nor U3255 (N_3255,In_397,In_1503);
nand U3256 (N_3256,In_1815,In_1321);
nand U3257 (N_3257,In_349,In_926);
nor U3258 (N_3258,In_138,In_691);
nor U3259 (N_3259,In_1226,In_1829);
xor U3260 (N_3260,In_867,In_1433);
or U3261 (N_3261,In_1636,In_401);
and U3262 (N_3262,In_798,In_1016);
or U3263 (N_3263,In_950,In_233);
and U3264 (N_3264,In_903,In_849);
and U3265 (N_3265,In_151,In_1662);
and U3266 (N_3266,In_608,In_447);
xor U3267 (N_3267,In_1877,In_244);
nand U3268 (N_3268,In_223,In_1700);
nor U3269 (N_3269,In_1745,In_669);
nand U3270 (N_3270,In_1491,In_119);
nand U3271 (N_3271,In_95,In_1158);
nor U3272 (N_3272,In_147,In_465);
and U3273 (N_3273,In_1475,In_383);
nor U3274 (N_3274,In_425,In_1467);
and U3275 (N_3275,In_1367,In_739);
and U3276 (N_3276,In_1100,In_878);
nand U3277 (N_3277,In_1334,In_370);
and U3278 (N_3278,In_1273,In_1491);
nand U3279 (N_3279,In_688,In_64);
xnor U3280 (N_3280,In_941,In_1015);
nor U3281 (N_3281,In_1783,In_884);
and U3282 (N_3282,In_1990,In_1408);
nand U3283 (N_3283,In_494,In_529);
xor U3284 (N_3284,In_190,In_1871);
nand U3285 (N_3285,In_1074,In_1821);
or U3286 (N_3286,In_646,In_265);
or U3287 (N_3287,In_1912,In_634);
and U3288 (N_3288,In_797,In_519);
nor U3289 (N_3289,In_1581,In_659);
or U3290 (N_3290,In_1353,In_1158);
and U3291 (N_3291,In_495,In_664);
nor U3292 (N_3292,In_1491,In_507);
or U3293 (N_3293,In_865,In_1833);
nor U3294 (N_3294,In_1883,In_61);
nand U3295 (N_3295,In_357,In_459);
xnor U3296 (N_3296,In_1133,In_1801);
nor U3297 (N_3297,In_392,In_230);
xnor U3298 (N_3298,In_708,In_181);
xor U3299 (N_3299,In_1105,In_147);
or U3300 (N_3300,In_1389,In_579);
or U3301 (N_3301,In_12,In_993);
or U3302 (N_3302,In_1335,In_115);
nand U3303 (N_3303,In_1987,In_1920);
or U3304 (N_3304,In_240,In_1222);
nor U3305 (N_3305,In_1759,In_1229);
nor U3306 (N_3306,In_903,In_122);
nand U3307 (N_3307,In_342,In_770);
nand U3308 (N_3308,In_1837,In_1772);
nor U3309 (N_3309,In_1176,In_338);
or U3310 (N_3310,In_727,In_799);
or U3311 (N_3311,In_1436,In_854);
and U3312 (N_3312,In_44,In_477);
nand U3313 (N_3313,In_1919,In_659);
and U3314 (N_3314,In_695,In_665);
or U3315 (N_3315,In_1197,In_1467);
nor U3316 (N_3316,In_80,In_62);
and U3317 (N_3317,In_175,In_16);
and U3318 (N_3318,In_993,In_1369);
nand U3319 (N_3319,In_21,In_1383);
nand U3320 (N_3320,In_428,In_952);
nor U3321 (N_3321,In_872,In_191);
or U3322 (N_3322,In_1869,In_1575);
nand U3323 (N_3323,In_1969,In_1036);
and U3324 (N_3324,In_435,In_308);
or U3325 (N_3325,In_1303,In_398);
and U3326 (N_3326,In_1993,In_412);
and U3327 (N_3327,In_796,In_1495);
nor U3328 (N_3328,In_1420,In_879);
and U3329 (N_3329,In_462,In_1735);
and U3330 (N_3330,In_1734,In_1291);
nand U3331 (N_3331,In_1619,In_497);
nand U3332 (N_3332,In_137,In_1010);
nand U3333 (N_3333,In_376,In_1391);
nand U3334 (N_3334,In_1693,In_1582);
nand U3335 (N_3335,In_1639,In_1569);
or U3336 (N_3336,In_449,In_1313);
and U3337 (N_3337,In_1042,In_356);
nor U3338 (N_3338,In_1181,In_572);
nand U3339 (N_3339,In_855,In_1745);
nand U3340 (N_3340,In_457,In_344);
xnor U3341 (N_3341,In_616,In_736);
nand U3342 (N_3342,In_851,In_1894);
nor U3343 (N_3343,In_1376,In_1824);
nor U3344 (N_3344,In_308,In_1424);
xnor U3345 (N_3345,In_1992,In_1846);
nor U3346 (N_3346,In_675,In_1901);
and U3347 (N_3347,In_1719,In_323);
nor U3348 (N_3348,In_1244,In_713);
nor U3349 (N_3349,In_1389,In_1259);
nand U3350 (N_3350,In_1528,In_504);
or U3351 (N_3351,In_1936,In_1193);
and U3352 (N_3352,In_321,In_1911);
nand U3353 (N_3353,In_364,In_813);
nor U3354 (N_3354,In_1345,In_977);
nor U3355 (N_3355,In_171,In_1380);
or U3356 (N_3356,In_1290,In_466);
or U3357 (N_3357,In_1897,In_152);
nand U3358 (N_3358,In_26,In_403);
nor U3359 (N_3359,In_1168,In_1145);
nand U3360 (N_3360,In_781,In_1522);
nor U3361 (N_3361,In_829,In_144);
and U3362 (N_3362,In_1101,In_788);
or U3363 (N_3363,In_619,In_226);
and U3364 (N_3364,In_1742,In_585);
nor U3365 (N_3365,In_307,In_686);
and U3366 (N_3366,In_1544,In_1859);
xor U3367 (N_3367,In_288,In_966);
and U3368 (N_3368,In_100,In_442);
nand U3369 (N_3369,In_659,In_1362);
and U3370 (N_3370,In_135,In_642);
nand U3371 (N_3371,In_1842,In_125);
and U3372 (N_3372,In_671,In_537);
nand U3373 (N_3373,In_1824,In_1066);
and U3374 (N_3374,In_1671,In_1126);
and U3375 (N_3375,In_799,In_1157);
nor U3376 (N_3376,In_958,In_384);
nor U3377 (N_3377,In_1039,In_1202);
nor U3378 (N_3378,In_834,In_1290);
or U3379 (N_3379,In_314,In_1937);
and U3380 (N_3380,In_811,In_950);
and U3381 (N_3381,In_322,In_1749);
or U3382 (N_3382,In_764,In_1468);
xnor U3383 (N_3383,In_660,In_1280);
nor U3384 (N_3384,In_329,In_956);
nor U3385 (N_3385,In_470,In_1729);
nand U3386 (N_3386,In_47,In_1481);
and U3387 (N_3387,In_1349,In_1570);
or U3388 (N_3388,In_788,In_516);
and U3389 (N_3389,In_564,In_1299);
xnor U3390 (N_3390,In_390,In_176);
nor U3391 (N_3391,In_1052,In_1032);
nand U3392 (N_3392,In_523,In_1179);
and U3393 (N_3393,In_260,In_463);
nor U3394 (N_3394,In_1456,In_308);
and U3395 (N_3395,In_608,In_712);
xor U3396 (N_3396,In_1898,In_366);
or U3397 (N_3397,In_165,In_714);
xor U3398 (N_3398,In_1021,In_915);
nor U3399 (N_3399,In_916,In_1535);
or U3400 (N_3400,In_1477,In_966);
and U3401 (N_3401,In_1165,In_65);
and U3402 (N_3402,In_1016,In_1520);
xnor U3403 (N_3403,In_1477,In_699);
xnor U3404 (N_3404,In_1023,In_1530);
xor U3405 (N_3405,In_1247,In_1621);
and U3406 (N_3406,In_954,In_215);
nand U3407 (N_3407,In_243,In_867);
and U3408 (N_3408,In_89,In_312);
nor U3409 (N_3409,In_865,In_1246);
and U3410 (N_3410,In_1127,In_117);
nand U3411 (N_3411,In_1903,In_112);
and U3412 (N_3412,In_163,In_519);
nor U3413 (N_3413,In_1372,In_1726);
or U3414 (N_3414,In_482,In_745);
xnor U3415 (N_3415,In_1273,In_242);
and U3416 (N_3416,In_529,In_1979);
nand U3417 (N_3417,In_1168,In_110);
or U3418 (N_3418,In_1455,In_340);
or U3419 (N_3419,In_1639,In_1899);
xor U3420 (N_3420,In_1104,In_1150);
xnor U3421 (N_3421,In_1069,In_1846);
xor U3422 (N_3422,In_1975,In_1483);
and U3423 (N_3423,In_558,In_1198);
xor U3424 (N_3424,In_1836,In_156);
xor U3425 (N_3425,In_315,In_1393);
and U3426 (N_3426,In_1982,In_810);
nor U3427 (N_3427,In_721,In_522);
nand U3428 (N_3428,In_332,In_1444);
nand U3429 (N_3429,In_1886,In_276);
or U3430 (N_3430,In_1373,In_43);
or U3431 (N_3431,In_961,In_1291);
or U3432 (N_3432,In_34,In_1793);
nor U3433 (N_3433,In_432,In_1630);
nand U3434 (N_3434,In_1763,In_1409);
and U3435 (N_3435,In_612,In_888);
nand U3436 (N_3436,In_627,In_383);
or U3437 (N_3437,In_1680,In_1628);
or U3438 (N_3438,In_1637,In_1004);
and U3439 (N_3439,In_1528,In_1103);
and U3440 (N_3440,In_1454,In_1334);
and U3441 (N_3441,In_1113,In_1319);
and U3442 (N_3442,In_1862,In_1917);
or U3443 (N_3443,In_571,In_685);
nand U3444 (N_3444,In_1314,In_711);
and U3445 (N_3445,In_726,In_734);
nor U3446 (N_3446,In_636,In_547);
nand U3447 (N_3447,In_1832,In_1226);
nor U3448 (N_3448,In_1700,In_1070);
nor U3449 (N_3449,In_439,In_1323);
nor U3450 (N_3450,In_1948,In_1438);
or U3451 (N_3451,In_1789,In_1752);
and U3452 (N_3452,In_1133,In_947);
nand U3453 (N_3453,In_25,In_667);
and U3454 (N_3454,In_471,In_1241);
xnor U3455 (N_3455,In_1180,In_1764);
nor U3456 (N_3456,In_1279,In_208);
or U3457 (N_3457,In_426,In_525);
nor U3458 (N_3458,In_524,In_1261);
nor U3459 (N_3459,In_276,In_1104);
nor U3460 (N_3460,In_1779,In_73);
and U3461 (N_3461,In_1545,In_1575);
nor U3462 (N_3462,In_636,In_1779);
and U3463 (N_3463,In_1423,In_243);
and U3464 (N_3464,In_1760,In_142);
or U3465 (N_3465,In_16,In_351);
or U3466 (N_3466,In_1928,In_1633);
nand U3467 (N_3467,In_1526,In_1519);
nor U3468 (N_3468,In_841,In_576);
nor U3469 (N_3469,In_269,In_443);
and U3470 (N_3470,In_1308,In_589);
xnor U3471 (N_3471,In_853,In_1256);
or U3472 (N_3472,In_838,In_1905);
nor U3473 (N_3473,In_845,In_1675);
and U3474 (N_3474,In_348,In_305);
and U3475 (N_3475,In_1829,In_104);
nand U3476 (N_3476,In_1405,In_732);
or U3477 (N_3477,In_349,In_1644);
nand U3478 (N_3478,In_1146,In_1496);
and U3479 (N_3479,In_1863,In_495);
or U3480 (N_3480,In_86,In_1788);
nand U3481 (N_3481,In_1490,In_1910);
nand U3482 (N_3482,In_1604,In_613);
nand U3483 (N_3483,In_1580,In_634);
nor U3484 (N_3484,In_387,In_1431);
and U3485 (N_3485,In_20,In_1545);
nand U3486 (N_3486,In_131,In_1178);
nand U3487 (N_3487,In_1563,In_328);
nor U3488 (N_3488,In_1722,In_1008);
nand U3489 (N_3489,In_91,In_1867);
and U3490 (N_3490,In_385,In_1100);
nand U3491 (N_3491,In_443,In_844);
and U3492 (N_3492,In_1280,In_1165);
or U3493 (N_3493,In_347,In_1177);
nand U3494 (N_3494,In_617,In_616);
nor U3495 (N_3495,In_1262,In_1915);
nand U3496 (N_3496,In_394,In_1204);
or U3497 (N_3497,In_1602,In_1693);
xnor U3498 (N_3498,In_1366,In_827);
or U3499 (N_3499,In_1834,In_392);
or U3500 (N_3500,In_418,In_1876);
xor U3501 (N_3501,In_1137,In_1060);
and U3502 (N_3502,In_1100,In_1507);
xnor U3503 (N_3503,In_1450,In_1129);
or U3504 (N_3504,In_975,In_577);
or U3505 (N_3505,In_1450,In_482);
or U3506 (N_3506,In_1678,In_433);
xor U3507 (N_3507,In_1649,In_1748);
xor U3508 (N_3508,In_967,In_564);
and U3509 (N_3509,In_1009,In_1084);
nor U3510 (N_3510,In_850,In_1352);
and U3511 (N_3511,In_461,In_901);
and U3512 (N_3512,In_1115,In_1200);
or U3513 (N_3513,In_322,In_914);
and U3514 (N_3514,In_1185,In_1358);
xor U3515 (N_3515,In_1042,In_1855);
nor U3516 (N_3516,In_1229,In_254);
and U3517 (N_3517,In_1498,In_1776);
nand U3518 (N_3518,In_1211,In_896);
or U3519 (N_3519,In_559,In_1080);
nand U3520 (N_3520,In_1689,In_32);
or U3521 (N_3521,In_1609,In_803);
xnor U3522 (N_3522,In_167,In_1296);
and U3523 (N_3523,In_641,In_1266);
nor U3524 (N_3524,In_1874,In_470);
xnor U3525 (N_3525,In_1049,In_209);
and U3526 (N_3526,In_244,In_88);
and U3527 (N_3527,In_1232,In_1714);
nor U3528 (N_3528,In_345,In_1389);
xor U3529 (N_3529,In_1134,In_1647);
nor U3530 (N_3530,In_709,In_36);
xor U3531 (N_3531,In_520,In_1434);
nor U3532 (N_3532,In_1797,In_565);
or U3533 (N_3533,In_983,In_894);
nor U3534 (N_3534,In_1433,In_805);
or U3535 (N_3535,In_741,In_356);
nand U3536 (N_3536,In_1867,In_325);
nand U3537 (N_3537,In_604,In_799);
nand U3538 (N_3538,In_1541,In_1781);
nor U3539 (N_3539,In_544,In_1193);
or U3540 (N_3540,In_900,In_240);
or U3541 (N_3541,In_1896,In_92);
nor U3542 (N_3542,In_258,In_806);
nor U3543 (N_3543,In_1955,In_896);
nand U3544 (N_3544,In_1570,In_1369);
nor U3545 (N_3545,In_1920,In_230);
nand U3546 (N_3546,In_477,In_1663);
or U3547 (N_3547,In_110,In_1588);
nand U3548 (N_3548,In_1194,In_1610);
xor U3549 (N_3549,In_1116,In_1969);
nand U3550 (N_3550,In_1544,In_950);
and U3551 (N_3551,In_1923,In_695);
or U3552 (N_3552,In_1176,In_864);
nand U3553 (N_3553,In_25,In_97);
or U3554 (N_3554,In_363,In_1747);
xnor U3555 (N_3555,In_597,In_1729);
or U3556 (N_3556,In_1557,In_1522);
xor U3557 (N_3557,In_1093,In_1033);
nor U3558 (N_3558,In_934,In_1293);
or U3559 (N_3559,In_535,In_1343);
or U3560 (N_3560,In_1809,In_1507);
nor U3561 (N_3561,In_153,In_1420);
nand U3562 (N_3562,In_42,In_1141);
nand U3563 (N_3563,In_1239,In_1033);
nand U3564 (N_3564,In_883,In_581);
and U3565 (N_3565,In_1878,In_1042);
or U3566 (N_3566,In_745,In_312);
nor U3567 (N_3567,In_609,In_307);
nand U3568 (N_3568,In_928,In_487);
nor U3569 (N_3569,In_872,In_1479);
nand U3570 (N_3570,In_78,In_158);
nand U3571 (N_3571,In_879,In_1903);
nor U3572 (N_3572,In_591,In_921);
nor U3573 (N_3573,In_1959,In_1307);
nor U3574 (N_3574,In_976,In_1052);
nand U3575 (N_3575,In_672,In_237);
or U3576 (N_3576,In_1707,In_1315);
nor U3577 (N_3577,In_794,In_1466);
and U3578 (N_3578,In_706,In_143);
nand U3579 (N_3579,In_779,In_1770);
nor U3580 (N_3580,In_1836,In_1399);
xnor U3581 (N_3581,In_442,In_93);
and U3582 (N_3582,In_1553,In_464);
nor U3583 (N_3583,In_41,In_773);
xnor U3584 (N_3584,In_1616,In_1424);
and U3585 (N_3585,In_1895,In_1122);
or U3586 (N_3586,In_1525,In_421);
nor U3587 (N_3587,In_524,In_907);
nand U3588 (N_3588,In_700,In_715);
or U3589 (N_3589,In_378,In_1509);
nand U3590 (N_3590,In_1509,In_735);
or U3591 (N_3591,In_430,In_38);
xnor U3592 (N_3592,In_1633,In_589);
or U3593 (N_3593,In_424,In_298);
nand U3594 (N_3594,In_889,In_1004);
nor U3595 (N_3595,In_1814,In_1466);
or U3596 (N_3596,In_1361,In_477);
or U3597 (N_3597,In_518,In_981);
and U3598 (N_3598,In_378,In_1260);
nor U3599 (N_3599,In_1214,In_1712);
or U3600 (N_3600,In_1618,In_1957);
xor U3601 (N_3601,In_1902,In_1536);
nand U3602 (N_3602,In_258,In_585);
nand U3603 (N_3603,In_1481,In_313);
or U3604 (N_3604,In_1576,In_1173);
xnor U3605 (N_3605,In_237,In_1980);
and U3606 (N_3606,In_863,In_902);
or U3607 (N_3607,In_1075,In_1568);
or U3608 (N_3608,In_1267,In_1094);
and U3609 (N_3609,In_744,In_751);
and U3610 (N_3610,In_342,In_1735);
and U3611 (N_3611,In_674,In_596);
and U3612 (N_3612,In_1492,In_945);
xor U3613 (N_3613,In_725,In_1227);
nor U3614 (N_3614,In_1357,In_626);
and U3615 (N_3615,In_583,In_1078);
or U3616 (N_3616,In_613,In_1501);
nor U3617 (N_3617,In_283,In_1025);
or U3618 (N_3618,In_217,In_1333);
nor U3619 (N_3619,In_1697,In_0);
nand U3620 (N_3620,In_551,In_759);
nand U3621 (N_3621,In_801,In_1674);
or U3622 (N_3622,In_646,In_1409);
or U3623 (N_3623,In_1873,In_410);
and U3624 (N_3624,In_1532,In_759);
nand U3625 (N_3625,In_781,In_854);
or U3626 (N_3626,In_929,In_286);
or U3627 (N_3627,In_1788,In_1552);
xor U3628 (N_3628,In_1209,In_1494);
nand U3629 (N_3629,In_226,In_1919);
and U3630 (N_3630,In_1568,In_1446);
nor U3631 (N_3631,In_1982,In_82);
xor U3632 (N_3632,In_1919,In_1728);
and U3633 (N_3633,In_360,In_46);
or U3634 (N_3634,In_438,In_1822);
and U3635 (N_3635,In_684,In_4);
nor U3636 (N_3636,In_503,In_1514);
nand U3637 (N_3637,In_62,In_1638);
and U3638 (N_3638,In_323,In_1712);
or U3639 (N_3639,In_343,In_308);
or U3640 (N_3640,In_23,In_193);
nand U3641 (N_3641,In_810,In_1404);
nor U3642 (N_3642,In_299,In_287);
nor U3643 (N_3643,In_1813,In_1290);
and U3644 (N_3644,In_1039,In_1845);
nor U3645 (N_3645,In_1768,In_789);
and U3646 (N_3646,In_1114,In_810);
nand U3647 (N_3647,In_795,In_540);
nand U3648 (N_3648,In_288,In_1630);
and U3649 (N_3649,In_1503,In_709);
or U3650 (N_3650,In_1070,In_1641);
and U3651 (N_3651,In_1310,In_1318);
xor U3652 (N_3652,In_1060,In_1500);
nor U3653 (N_3653,In_1136,In_1497);
nor U3654 (N_3654,In_1534,In_955);
or U3655 (N_3655,In_1014,In_1990);
and U3656 (N_3656,In_208,In_99);
or U3657 (N_3657,In_1945,In_1442);
and U3658 (N_3658,In_1769,In_267);
nor U3659 (N_3659,In_520,In_243);
nand U3660 (N_3660,In_1489,In_1187);
nor U3661 (N_3661,In_1768,In_124);
xor U3662 (N_3662,In_1387,In_648);
or U3663 (N_3663,In_953,In_323);
nor U3664 (N_3664,In_274,In_363);
xor U3665 (N_3665,In_755,In_1989);
nor U3666 (N_3666,In_239,In_1213);
xnor U3667 (N_3667,In_760,In_970);
nor U3668 (N_3668,In_1025,In_1802);
xor U3669 (N_3669,In_1150,In_1335);
nand U3670 (N_3670,In_1087,In_1076);
nand U3671 (N_3671,In_1768,In_1801);
or U3672 (N_3672,In_1017,In_1406);
and U3673 (N_3673,In_869,In_1890);
nand U3674 (N_3674,In_842,In_440);
and U3675 (N_3675,In_1642,In_657);
or U3676 (N_3676,In_639,In_343);
and U3677 (N_3677,In_280,In_1820);
or U3678 (N_3678,In_997,In_1924);
or U3679 (N_3679,In_879,In_1676);
nand U3680 (N_3680,In_1697,In_1291);
and U3681 (N_3681,In_71,In_651);
nand U3682 (N_3682,In_1488,In_188);
nor U3683 (N_3683,In_899,In_547);
nor U3684 (N_3684,In_482,In_1603);
nor U3685 (N_3685,In_406,In_76);
nor U3686 (N_3686,In_332,In_1736);
or U3687 (N_3687,In_319,In_865);
and U3688 (N_3688,In_1979,In_1476);
nand U3689 (N_3689,In_359,In_1716);
nor U3690 (N_3690,In_1340,In_1058);
and U3691 (N_3691,In_782,In_25);
nor U3692 (N_3692,In_708,In_879);
or U3693 (N_3693,In_358,In_373);
nor U3694 (N_3694,In_375,In_1473);
nand U3695 (N_3695,In_1106,In_399);
nor U3696 (N_3696,In_1881,In_668);
and U3697 (N_3697,In_88,In_656);
or U3698 (N_3698,In_850,In_359);
and U3699 (N_3699,In_1881,In_1178);
nor U3700 (N_3700,In_1013,In_1941);
nand U3701 (N_3701,In_660,In_1344);
and U3702 (N_3702,In_1943,In_14);
nor U3703 (N_3703,In_1657,In_1038);
nand U3704 (N_3704,In_786,In_837);
nor U3705 (N_3705,In_565,In_611);
nand U3706 (N_3706,In_390,In_1859);
and U3707 (N_3707,In_1885,In_1770);
nand U3708 (N_3708,In_1029,In_993);
and U3709 (N_3709,In_1257,In_895);
xnor U3710 (N_3710,In_1019,In_982);
nor U3711 (N_3711,In_842,In_891);
or U3712 (N_3712,In_21,In_918);
and U3713 (N_3713,In_1725,In_1951);
and U3714 (N_3714,In_933,In_1961);
or U3715 (N_3715,In_1684,In_1138);
nor U3716 (N_3716,In_1432,In_539);
and U3717 (N_3717,In_668,In_1659);
nor U3718 (N_3718,In_1202,In_43);
nand U3719 (N_3719,In_606,In_1196);
and U3720 (N_3720,In_978,In_344);
nand U3721 (N_3721,In_616,In_1231);
nand U3722 (N_3722,In_874,In_1302);
nand U3723 (N_3723,In_1934,In_1442);
or U3724 (N_3724,In_1876,In_692);
and U3725 (N_3725,In_1242,In_1142);
or U3726 (N_3726,In_84,In_1902);
xnor U3727 (N_3727,In_1105,In_771);
xnor U3728 (N_3728,In_409,In_1951);
nor U3729 (N_3729,In_1768,In_1016);
or U3730 (N_3730,In_1439,In_1872);
or U3731 (N_3731,In_125,In_448);
xor U3732 (N_3732,In_1490,In_1415);
nor U3733 (N_3733,In_1291,In_1860);
nor U3734 (N_3734,In_718,In_1962);
or U3735 (N_3735,In_1869,In_1290);
or U3736 (N_3736,In_1523,In_1897);
and U3737 (N_3737,In_1573,In_264);
nand U3738 (N_3738,In_371,In_561);
or U3739 (N_3739,In_4,In_1551);
and U3740 (N_3740,In_1642,In_971);
and U3741 (N_3741,In_1112,In_1725);
nor U3742 (N_3742,In_1798,In_1931);
or U3743 (N_3743,In_848,In_298);
and U3744 (N_3744,In_149,In_1898);
nor U3745 (N_3745,In_1176,In_487);
and U3746 (N_3746,In_1615,In_1403);
nand U3747 (N_3747,In_144,In_1780);
nor U3748 (N_3748,In_1774,In_1938);
nand U3749 (N_3749,In_1223,In_1128);
and U3750 (N_3750,In_823,In_303);
or U3751 (N_3751,In_1311,In_1159);
nor U3752 (N_3752,In_846,In_1572);
nor U3753 (N_3753,In_740,In_1724);
or U3754 (N_3754,In_1593,In_993);
nand U3755 (N_3755,In_1524,In_600);
nand U3756 (N_3756,In_874,In_652);
nor U3757 (N_3757,In_1308,In_304);
and U3758 (N_3758,In_436,In_632);
xor U3759 (N_3759,In_527,In_592);
nor U3760 (N_3760,In_1225,In_1192);
nor U3761 (N_3761,In_707,In_1634);
xor U3762 (N_3762,In_818,In_1960);
or U3763 (N_3763,In_1054,In_1570);
nand U3764 (N_3764,In_538,In_248);
or U3765 (N_3765,In_1206,In_1863);
or U3766 (N_3766,In_309,In_1707);
xnor U3767 (N_3767,In_26,In_371);
nand U3768 (N_3768,In_1797,In_1985);
and U3769 (N_3769,In_1373,In_1640);
or U3770 (N_3770,In_461,In_652);
xnor U3771 (N_3771,In_724,In_1353);
or U3772 (N_3772,In_1495,In_1719);
xnor U3773 (N_3773,In_1459,In_276);
and U3774 (N_3774,In_1772,In_1438);
nand U3775 (N_3775,In_1166,In_494);
or U3776 (N_3776,In_860,In_332);
or U3777 (N_3777,In_463,In_709);
nand U3778 (N_3778,In_419,In_354);
nand U3779 (N_3779,In_1133,In_319);
and U3780 (N_3780,In_285,In_946);
nand U3781 (N_3781,In_102,In_1115);
and U3782 (N_3782,In_747,In_75);
nor U3783 (N_3783,In_103,In_18);
and U3784 (N_3784,In_929,In_1290);
nor U3785 (N_3785,In_1209,In_1615);
or U3786 (N_3786,In_1881,In_259);
xor U3787 (N_3787,In_1849,In_53);
nor U3788 (N_3788,In_786,In_666);
and U3789 (N_3789,In_1360,In_1990);
nand U3790 (N_3790,In_1503,In_60);
nor U3791 (N_3791,In_891,In_317);
or U3792 (N_3792,In_564,In_11);
or U3793 (N_3793,In_1360,In_678);
or U3794 (N_3794,In_1748,In_473);
or U3795 (N_3795,In_1065,In_1197);
xor U3796 (N_3796,In_1397,In_1565);
or U3797 (N_3797,In_1578,In_1098);
nor U3798 (N_3798,In_172,In_628);
or U3799 (N_3799,In_970,In_1592);
and U3800 (N_3800,In_1639,In_1672);
and U3801 (N_3801,In_1047,In_1672);
nand U3802 (N_3802,In_37,In_1494);
nor U3803 (N_3803,In_830,In_1061);
and U3804 (N_3804,In_871,In_677);
nor U3805 (N_3805,In_1396,In_887);
nor U3806 (N_3806,In_302,In_869);
nand U3807 (N_3807,In_592,In_525);
nor U3808 (N_3808,In_1825,In_826);
nand U3809 (N_3809,In_1630,In_1211);
xnor U3810 (N_3810,In_636,In_1936);
and U3811 (N_3811,In_1388,In_1625);
and U3812 (N_3812,In_1781,In_1695);
nor U3813 (N_3813,In_1208,In_794);
nor U3814 (N_3814,In_569,In_225);
nor U3815 (N_3815,In_1834,In_60);
nor U3816 (N_3816,In_1798,In_769);
and U3817 (N_3817,In_1339,In_566);
or U3818 (N_3818,In_491,In_190);
and U3819 (N_3819,In_1232,In_200);
and U3820 (N_3820,In_997,In_41);
or U3821 (N_3821,In_1852,In_655);
nand U3822 (N_3822,In_1057,In_1938);
or U3823 (N_3823,In_944,In_1292);
nand U3824 (N_3824,In_1068,In_343);
or U3825 (N_3825,In_251,In_1335);
nand U3826 (N_3826,In_1794,In_752);
xor U3827 (N_3827,In_185,In_1958);
nand U3828 (N_3828,In_1527,In_830);
nor U3829 (N_3829,In_1971,In_754);
nor U3830 (N_3830,In_922,In_165);
nand U3831 (N_3831,In_681,In_116);
and U3832 (N_3832,In_29,In_1155);
or U3833 (N_3833,In_1466,In_978);
xor U3834 (N_3834,In_767,In_791);
nor U3835 (N_3835,In_1710,In_1442);
and U3836 (N_3836,In_684,In_411);
nand U3837 (N_3837,In_635,In_1049);
and U3838 (N_3838,In_1108,In_29);
and U3839 (N_3839,In_1644,In_1937);
or U3840 (N_3840,In_778,In_339);
nor U3841 (N_3841,In_451,In_297);
and U3842 (N_3842,In_1653,In_290);
nor U3843 (N_3843,In_568,In_168);
and U3844 (N_3844,In_1617,In_1353);
nand U3845 (N_3845,In_504,In_883);
and U3846 (N_3846,In_406,In_1832);
nand U3847 (N_3847,In_74,In_221);
nor U3848 (N_3848,In_246,In_350);
nor U3849 (N_3849,In_803,In_378);
nor U3850 (N_3850,In_1624,In_467);
xor U3851 (N_3851,In_1488,In_1520);
or U3852 (N_3852,In_1086,In_1087);
nor U3853 (N_3853,In_1107,In_1937);
or U3854 (N_3854,In_155,In_402);
nor U3855 (N_3855,In_426,In_1605);
nand U3856 (N_3856,In_221,In_1368);
or U3857 (N_3857,In_1515,In_1734);
nor U3858 (N_3858,In_1930,In_688);
and U3859 (N_3859,In_1476,In_859);
xor U3860 (N_3860,In_590,In_560);
and U3861 (N_3861,In_969,In_1445);
and U3862 (N_3862,In_1279,In_298);
nand U3863 (N_3863,In_517,In_1357);
and U3864 (N_3864,In_1024,In_986);
nor U3865 (N_3865,In_1359,In_1314);
xnor U3866 (N_3866,In_742,In_541);
or U3867 (N_3867,In_1698,In_1191);
or U3868 (N_3868,In_1120,In_1398);
nor U3869 (N_3869,In_622,In_847);
or U3870 (N_3870,In_487,In_1090);
or U3871 (N_3871,In_604,In_593);
and U3872 (N_3872,In_839,In_238);
nor U3873 (N_3873,In_30,In_7);
nand U3874 (N_3874,In_273,In_1434);
nand U3875 (N_3875,In_232,In_1678);
or U3876 (N_3876,In_1667,In_1836);
nor U3877 (N_3877,In_741,In_1779);
and U3878 (N_3878,In_1735,In_946);
nor U3879 (N_3879,In_372,In_1474);
nor U3880 (N_3880,In_624,In_985);
xnor U3881 (N_3881,In_9,In_1860);
or U3882 (N_3882,In_277,In_174);
xor U3883 (N_3883,In_1146,In_1523);
nand U3884 (N_3884,In_1749,In_134);
and U3885 (N_3885,In_416,In_1038);
and U3886 (N_3886,In_820,In_564);
nand U3887 (N_3887,In_391,In_742);
nand U3888 (N_3888,In_417,In_411);
or U3889 (N_3889,In_736,In_1719);
nor U3890 (N_3890,In_1945,In_1075);
or U3891 (N_3891,In_1565,In_1375);
or U3892 (N_3892,In_1653,In_1882);
nand U3893 (N_3893,In_1505,In_577);
and U3894 (N_3894,In_1629,In_1098);
or U3895 (N_3895,In_911,In_1150);
and U3896 (N_3896,In_1042,In_1758);
and U3897 (N_3897,In_1082,In_1671);
and U3898 (N_3898,In_434,In_1564);
nand U3899 (N_3899,In_819,In_1541);
and U3900 (N_3900,In_1880,In_1719);
nand U3901 (N_3901,In_1757,In_979);
or U3902 (N_3902,In_847,In_585);
nand U3903 (N_3903,In_1472,In_17);
nor U3904 (N_3904,In_1219,In_1736);
and U3905 (N_3905,In_1393,In_1304);
nand U3906 (N_3906,In_1132,In_1707);
nand U3907 (N_3907,In_222,In_434);
xor U3908 (N_3908,In_398,In_407);
nand U3909 (N_3909,In_1448,In_500);
nor U3910 (N_3910,In_1428,In_1140);
and U3911 (N_3911,In_1883,In_895);
nand U3912 (N_3912,In_1430,In_1059);
or U3913 (N_3913,In_1040,In_606);
or U3914 (N_3914,In_370,In_1211);
or U3915 (N_3915,In_10,In_1527);
and U3916 (N_3916,In_1630,In_964);
or U3917 (N_3917,In_320,In_1555);
or U3918 (N_3918,In_1568,In_917);
nor U3919 (N_3919,In_404,In_1288);
nand U3920 (N_3920,In_981,In_112);
nor U3921 (N_3921,In_1081,In_1931);
and U3922 (N_3922,In_84,In_1305);
nand U3923 (N_3923,In_371,In_2);
nand U3924 (N_3924,In_1117,In_754);
xor U3925 (N_3925,In_1596,In_241);
and U3926 (N_3926,In_1662,In_1542);
xor U3927 (N_3927,In_450,In_1393);
nor U3928 (N_3928,In_10,In_1273);
nor U3929 (N_3929,In_752,In_66);
xor U3930 (N_3930,In_824,In_484);
nor U3931 (N_3931,In_1758,In_849);
or U3932 (N_3932,In_1938,In_625);
or U3933 (N_3933,In_141,In_410);
nand U3934 (N_3934,In_478,In_885);
and U3935 (N_3935,In_1112,In_11);
nor U3936 (N_3936,In_1173,In_447);
xnor U3937 (N_3937,In_373,In_1610);
nor U3938 (N_3938,In_639,In_1884);
and U3939 (N_3939,In_1106,In_1935);
nand U3940 (N_3940,In_1762,In_1812);
or U3941 (N_3941,In_1806,In_1765);
nor U3942 (N_3942,In_911,In_1925);
xor U3943 (N_3943,In_231,In_1992);
or U3944 (N_3944,In_1523,In_1853);
and U3945 (N_3945,In_1481,In_696);
or U3946 (N_3946,In_1866,In_599);
and U3947 (N_3947,In_885,In_1489);
or U3948 (N_3948,In_550,In_1938);
nor U3949 (N_3949,In_1370,In_1524);
and U3950 (N_3950,In_1978,In_924);
xor U3951 (N_3951,In_1588,In_28);
and U3952 (N_3952,In_785,In_720);
or U3953 (N_3953,In_992,In_794);
nor U3954 (N_3954,In_967,In_1377);
nand U3955 (N_3955,In_1406,In_384);
or U3956 (N_3956,In_823,In_1872);
nor U3957 (N_3957,In_1258,In_1314);
and U3958 (N_3958,In_1567,In_1550);
xnor U3959 (N_3959,In_491,In_108);
or U3960 (N_3960,In_500,In_179);
xor U3961 (N_3961,In_1778,In_188);
or U3962 (N_3962,In_1662,In_1393);
nor U3963 (N_3963,In_933,In_1085);
nor U3964 (N_3964,In_677,In_403);
and U3965 (N_3965,In_1177,In_1238);
nand U3966 (N_3966,In_872,In_722);
xor U3967 (N_3967,In_1502,In_1097);
or U3968 (N_3968,In_1844,In_526);
nor U3969 (N_3969,In_821,In_313);
and U3970 (N_3970,In_382,In_1479);
nand U3971 (N_3971,In_266,In_618);
nand U3972 (N_3972,In_24,In_761);
or U3973 (N_3973,In_235,In_1684);
nor U3974 (N_3974,In_1350,In_627);
or U3975 (N_3975,In_1104,In_1562);
nand U3976 (N_3976,In_1370,In_1424);
nand U3977 (N_3977,In_575,In_1355);
nor U3978 (N_3978,In_1529,In_161);
nand U3979 (N_3979,In_1219,In_1653);
and U3980 (N_3980,In_1854,In_797);
or U3981 (N_3981,In_467,In_960);
nor U3982 (N_3982,In_462,In_1343);
and U3983 (N_3983,In_747,In_1175);
nor U3984 (N_3984,In_1865,In_1867);
nand U3985 (N_3985,In_793,In_1314);
nand U3986 (N_3986,In_1560,In_10);
nand U3987 (N_3987,In_1416,In_681);
or U3988 (N_3988,In_1362,In_1816);
or U3989 (N_3989,In_1488,In_837);
and U3990 (N_3990,In_1301,In_253);
xor U3991 (N_3991,In_1656,In_965);
xnor U3992 (N_3992,In_1138,In_1479);
or U3993 (N_3993,In_1900,In_196);
nor U3994 (N_3994,In_1478,In_1831);
xor U3995 (N_3995,In_1343,In_617);
or U3996 (N_3996,In_226,In_1608);
and U3997 (N_3997,In_1148,In_374);
or U3998 (N_3998,In_884,In_1281);
or U3999 (N_3999,In_1706,In_767);
or U4000 (N_4000,N_1321,N_2025);
and U4001 (N_4001,N_2994,N_1004);
or U4002 (N_4002,N_3969,N_1879);
and U4003 (N_4003,N_80,N_3613);
nand U4004 (N_4004,N_1048,N_3346);
and U4005 (N_4005,N_903,N_1935);
and U4006 (N_4006,N_141,N_3197);
nand U4007 (N_4007,N_1731,N_179);
nand U4008 (N_4008,N_3411,N_3478);
nand U4009 (N_4009,N_1784,N_3959);
nand U4010 (N_4010,N_738,N_1546);
nand U4011 (N_4011,N_793,N_222);
xnor U4012 (N_4012,N_1076,N_3087);
nor U4013 (N_4013,N_2352,N_610);
nand U4014 (N_4014,N_1122,N_752);
and U4015 (N_4015,N_2164,N_2793);
nor U4016 (N_4016,N_3382,N_2056);
nor U4017 (N_4017,N_770,N_335);
and U4018 (N_4018,N_748,N_3057);
or U4019 (N_4019,N_2970,N_282);
xnor U4020 (N_4020,N_1408,N_686);
nor U4021 (N_4021,N_1206,N_1778);
nor U4022 (N_4022,N_873,N_3585);
and U4023 (N_4023,N_3068,N_1676);
nand U4024 (N_4024,N_110,N_3916);
and U4025 (N_4025,N_236,N_3231);
and U4026 (N_4026,N_2696,N_3279);
or U4027 (N_4027,N_1572,N_123);
nor U4028 (N_4028,N_3256,N_1913);
or U4029 (N_4029,N_2724,N_168);
and U4030 (N_4030,N_594,N_235);
nand U4031 (N_4031,N_1355,N_2374);
nand U4032 (N_4032,N_3958,N_1673);
xor U4033 (N_4033,N_46,N_1767);
nor U4034 (N_4034,N_2776,N_2565);
nor U4035 (N_4035,N_1046,N_263);
and U4036 (N_4036,N_1082,N_219);
nor U4037 (N_4037,N_1325,N_3735);
or U4038 (N_4038,N_1176,N_65);
nor U4039 (N_4039,N_3980,N_3311);
and U4040 (N_4040,N_634,N_2801);
or U4041 (N_4041,N_1818,N_1961);
nor U4042 (N_4042,N_907,N_3862);
and U4043 (N_4043,N_1432,N_356);
nand U4044 (N_4044,N_3496,N_3795);
nor U4045 (N_4045,N_1904,N_3117);
nor U4046 (N_4046,N_290,N_2212);
or U4047 (N_4047,N_2548,N_145);
nor U4048 (N_4048,N_1398,N_3706);
nand U4049 (N_4049,N_2690,N_3334);
xor U4050 (N_4050,N_1967,N_2169);
nand U4051 (N_4051,N_2892,N_3832);
and U4052 (N_4052,N_1926,N_39);
nor U4053 (N_4053,N_3828,N_3244);
or U4054 (N_4054,N_863,N_2803);
and U4055 (N_4055,N_1882,N_3562);
or U4056 (N_4056,N_1244,N_1385);
nand U4057 (N_4057,N_850,N_3645);
or U4058 (N_4058,N_2439,N_2887);
nor U4059 (N_4059,N_2550,N_1171);
nor U4060 (N_4060,N_552,N_3434);
and U4061 (N_4061,N_2507,N_1929);
nand U4062 (N_4062,N_2030,N_2866);
and U4063 (N_4063,N_2980,N_424);
nand U4064 (N_4064,N_3196,N_2356);
nor U4065 (N_4065,N_2010,N_464);
nand U4066 (N_4066,N_171,N_3705);
and U4067 (N_4067,N_2009,N_725);
or U4068 (N_4068,N_573,N_2326);
and U4069 (N_4069,N_1212,N_2131);
and U4070 (N_4070,N_2130,N_3092);
or U4071 (N_4071,N_2218,N_1420);
or U4072 (N_4072,N_718,N_2305);
nand U4073 (N_4073,N_302,N_1607);
nand U4074 (N_4074,N_722,N_2313);
nand U4075 (N_4075,N_1628,N_3631);
nand U4076 (N_4076,N_2713,N_2201);
or U4077 (N_4077,N_1258,N_3050);
or U4078 (N_4078,N_797,N_1109);
xor U4079 (N_4079,N_773,N_375);
nor U4080 (N_4080,N_2469,N_1680);
or U4081 (N_4081,N_104,N_3979);
or U4082 (N_4082,N_1699,N_2271);
nand U4083 (N_4083,N_1378,N_3622);
and U4084 (N_4084,N_2979,N_2945);
or U4085 (N_4085,N_2465,N_3712);
or U4086 (N_4086,N_689,N_369);
and U4087 (N_4087,N_124,N_2826);
and U4088 (N_4088,N_245,N_2380);
nor U4089 (N_4089,N_2828,N_3567);
and U4090 (N_4090,N_451,N_1865);
and U4091 (N_4091,N_1266,N_2347);
and U4092 (N_4092,N_692,N_3161);
or U4093 (N_4093,N_2925,N_212);
xor U4094 (N_4094,N_3599,N_827);
xor U4095 (N_4095,N_1016,N_3544);
or U4096 (N_4096,N_38,N_711);
or U4097 (N_4097,N_1544,N_3282);
nand U4098 (N_4098,N_1028,N_1);
and U4099 (N_4099,N_463,N_2038);
and U4100 (N_4100,N_1468,N_1548);
or U4101 (N_4101,N_361,N_3069);
or U4102 (N_4102,N_2228,N_996);
xor U4103 (N_4103,N_2991,N_3720);
nand U4104 (N_4104,N_1041,N_2244);
nand U4105 (N_4105,N_1257,N_2863);
xor U4106 (N_4106,N_1141,N_3215);
nor U4107 (N_4107,N_2762,N_3875);
or U4108 (N_4108,N_3321,N_2173);
or U4109 (N_4109,N_1602,N_2478);
nor U4110 (N_4110,N_2533,N_980);
or U4111 (N_4111,N_3651,N_240);
nand U4112 (N_4112,N_1578,N_3258);
and U4113 (N_4113,N_3265,N_2922);
nor U4114 (N_4114,N_3404,N_3464);
and U4115 (N_4115,N_1847,N_3878);
nand U4116 (N_4116,N_1391,N_2097);
or U4117 (N_4117,N_408,N_792);
nand U4118 (N_4118,N_2073,N_2425);
nand U4119 (N_4119,N_1466,N_1903);
or U4120 (N_4120,N_681,N_1182);
nand U4121 (N_4121,N_297,N_448);
or U4122 (N_4122,N_1002,N_1438);
or U4123 (N_4123,N_3108,N_1942);
nor U4124 (N_4124,N_3679,N_3836);
xnor U4125 (N_4125,N_3364,N_1284);
or U4126 (N_4126,N_1635,N_3157);
or U4127 (N_4127,N_983,N_2454);
or U4128 (N_4128,N_2032,N_1173);
or U4129 (N_4129,N_579,N_724);
xor U4130 (N_4130,N_2433,N_3417);
and U4131 (N_4131,N_3491,N_1955);
nand U4132 (N_4132,N_1817,N_3486);
nand U4133 (N_4133,N_3426,N_2984);
nor U4134 (N_4134,N_3228,N_596);
or U4135 (N_4135,N_1839,N_1781);
or U4136 (N_4136,N_3280,N_3052);
and U4137 (N_4137,N_1349,N_2785);
and U4138 (N_4138,N_2665,N_842);
nor U4139 (N_4139,N_2282,N_2294);
nand U4140 (N_4140,N_1130,N_3863);
nand U4141 (N_4141,N_2286,N_1744);
xnor U4142 (N_4142,N_2171,N_1019);
and U4143 (N_4143,N_1958,N_2265);
nor U4144 (N_4144,N_2539,N_3275);
nand U4145 (N_4145,N_477,N_326);
xnor U4146 (N_4146,N_3261,N_2728);
and U4147 (N_4147,N_1822,N_3489);
nor U4148 (N_4148,N_1703,N_446);
and U4149 (N_4149,N_0,N_3994);
nor U4150 (N_4150,N_2490,N_1830);
or U4151 (N_4151,N_2018,N_772);
nand U4152 (N_4152,N_1476,N_327);
or U4153 (N_4153,N_1768,N_1064);
nand U4154 (N_4154,N_1045,N_3349);
and U4155 (N_4155,N_2680,N_3109);
and U4156 (N_4156,N_2408,N_2522);
or U4157 (N_4157,N_1639,N_3507);
and U4158 (N_4158,N_2910,N_700);
or U4159 (N_4159,N_1189,N_2328);
nor U4160 (N_4160,N_252,N_407);
or U4161 (N_4161,N_509,N_3656);
nor U4162 (N_4162,N_3472,N_1299);
nand U4163 (N_4163,N_2404,N_760);
nor U4164 (N_4164,N_3596,N_277);
nand U4165 (N_4165,N_3281,N_609);
or U4166 (N_4166,N_2809,N_3754);
xnor U4167 (N_4167,N_591,N_1304);
nand U4168 (N_4168,N_13,N_2068);
and U4169 (N_4169,N_1060,N_668);
nor U4170 (N_4170,N_1196,N_3194);
and U4171 (N_4171,N_309,N_494);
nor U4172 (N_4172,N_2799,N_1871);
nand U4173 (N_4173,N_2476,N_1483);
xor U4174 (N_4174,N_945,N_1588);
and U4175 (N_4175,N_934,N_3377);
nor U4176 (N_4176,N_2114,N_3864);
xor U4177 (N_4177,N_3942,N_1001);
nor U4178 (N_4178,N_1647,N_2702);
or U4179 (N_4179,N_580,N_823);
nor U4180 (N_4180,N_3968,N_1256);
xor U4181 (N_4181,N_1855,N_1282);
nand U4182 (N_4182,N_2575,N_3013);
or U4183 (N_4183,N_3475,N_3744);
nor U4184 (N_4184,N_532,N_3106);
nor U4185 (N_4185,N_3698,N_2111);
or U4186 (N_4186,N_2428,N_2354);
nor U4187 (N_4187,N_1907,N_2623);
and U4188 (N_4188,N_2711,N_2978);
or U4189 (N_4189,N_1663,N_794);
and U4190 (N_4190,N_2930,N_3922);
or U4191 (N_4191,N_1086,N_487);
nand U4192 (N_4192,N_14,N_149);
or U4193 (N_4193,N_1401,N_3753);
or U4194 (N_4194,N_976,N_1869);
or U4195 (N_4195,N_729,N_488);
and U4196 (N_4196,N_1460,N_1192);
nor U4197 (N_4197,N_3722,N_227);
or U4198 (N_4198,N_561,N_1197);
xor U4199 (N_4199,N_430,N_2682);
and U4200 (N_4200,N_111,N_386);
nand U4201 (N_4201,N_2990,N_3331);
nor U4202 (N_4202,N_3771,N_1716);
nand U4203 (N_4203,N_2093,N_2578);
or U4204 (N_4204,N_3127,N_2932);
or U4205 (N_4205,N_1093,N_874);
nor U4206 (N_4206,N_2429,N_3949);
nor U4207 (N_4207,N_3881,N_2914);
nand U4208 (N_4208,N_1362,N_2614);
nand U4209 (N_4209,N_2192,N_2203);
xnor U4210 (N_4210,N_3232,N_3000);
xor U4211 (N_4211,N_501,N_3953);
and U4212 (N_4212,N_1912,N_1027);
nand U4213 (N_4213,N_1318,N_1627);
nor U4214 (N_4214,N_3083,N_3344);
xnor U4215 (N_4215,N_1412,N_2269);
and U4216 (N_4216,N_2086,N_2749);
nor U4217 (N_4217,N_1696,N_2455);
or U4218 (N_4218,N_2783,N_468);
or U4219 (N_4219,N_238,N_2051);
nand U4220 (N_4220,N_3335,N_1096);
or U4221 (N_4221,N_1665,N_2920);
nand U4222 (N_4222,N_3222,N_162);
or U4223 (N_4223,N_2461,N_1311);
and U4224 (N_4224,N_1095,N_1407);
and U4225 (N_4225,N_2243,N_3513);
and U4226 (N_4226,N_3394,N_2502);
or U4227 (N_4227,N_1821,N_2424);
nand U4228 (N_4228,N_916,N_3799);
and U4229 (N_4229,N_3868,N_2570);
nand U4230 (N_4230,N_1536,N_107);
nand U4231 (N_4231,N_1690,N_2035);
nor U4232 (N_4232,N_2880,N_1739);
xnor U4233 (N_4233,N_2733,N_3218);
nor U4234 (N_4234,N_1918,N_2572);
and U4235 (N_4235,N_1779,N_1292);
nor U4236 (N_4236,N_744,N_1145);
nand U4237 (N_4237,N_1714,N_2232);
and U4238 (N_4238,N_1654,N_1146);
nor U4239 (N_4239,N_188,N_777);
xnor U4240 (N_4240,N_1034,N_1344);
and U4241 (N_4241,N_745,N_3471);
nand U4242 (N_4242,N_1606,N_2976);
or U4243 (N_4243,N_28,N_1301);
and U4244 (N_4244,N_1389,N_226);
nand U4245 (N_4245,N_2403,N_2191);
nor U4246 (N_4246,N_3399,N_3607);
xor U4247 (N_4247,N_3427,N_2320);
xor U4248 (N_4248,N_3205,N_1278);
xnor U4249 (N_4249,N_841,N_1488);
or U4250 (N_4250,N_2480,N_1801);
nor U4251 (N_4251,N_3150,N_1701);
nor U4252 (N_4252,N_204,N_2685);
and U4253 (N_4253,N_3251,N_2705);
nand U4254 (N_4254,N_708,N_197);
nand U4255 (N_4255,N_790,N_3152);
xnor U4256 (N_4256,N_3073,N_1477);
xnor U4257 (N_4257,N_768,N_90);
nand U4258 (N_4258,N_3154,N_2481);
and U4259 (N_4259,N_1000,N_1241);
nand U4260 (N_4260,N_1799,N_1185);
xor U4261 (N_4261,N_881,N_714);
nand U4262 (N_4262,N_213,N_17);
nor U4263 (N_4263,N_3664,N_1899);
nor U4264 (N_4264,N_317,N_603);
or U4265 (N_4265,N_2773,N_3879);
xnor U4266 (N_4266,N_3669,N_2784);
or U4267 (N_4267,N_726,N_781);
nor U4268 (N_4268,N_1643,N_3590);
nor U4269 (N_4269,N_2491,N_1294);
nor U4270 (N_4270,N_698,N_19);
nand U4271 (N_4271,N_3522,N_1338);
xor U4272 (N_4272,N_2853,N_1660);
nor U4273 (N_4273,N_1634,N_3580);
nand U4274 (N_4274,N_3717,N_2897);
and U4275 (N_4275,N_938,N_1296);
nand U4276 (N_4276,N_2596,N_1988);
nand U4277 (N_4277,N_2082,N_1623);
and U4278 (N_4278,N_455,N_298);
and U4279 (N_4279,N_626,N_2593);
nor U4280 (N_4280,N_489,N_2398);
nand U4281 (N_4281,N_1062,N_112);
nand U4282 (N_4282,N_342,N_2158);
nor U4283 (N_4283,N_248,N_884);
and U4284 (N_4284,N_3707,N_1646);
or U4285 (N_4285,N_2147,N_258);
nor U4286 (N_4286,N_2715,N_821);
xor U4287 (N_4287,N_1638,N_584);
nor U4288 (N_4288,N_637,N_2759);
nor U4289 (N_4289,N_640,N_647);
nor U4290 (N_4290,N_2662,N_1782);
nand U4291 (N_4291,N_2193,N_2334);
nor U4292 (N_4292,N_1895,N_1564);
nand U4293 (N_4293,N_2797,N_2376);
or U4294 (N_4294,N_3495,N_3313);
nor U4295 (N_4295,N_3120,N_3032);
and U4296 (N_4296,N_3837,N_3571);
nand U4297 (N_4297,N_2775,N_1625);
and U4298 (N_4298,N_527,N_113);
or U4299 (N_4299,N_1126,N_1966);
or U4300 (N_4300,N_2995,N_502);
and U4301 (N_4301,N_3672,N_3220);
xor U4302 (N_4302,N_97,N_1252);
or U4303 (N_4303,N_2867,N_379);
nor U4304 (N_4304,N_2494,N_879);
nand U4305 (N_4305,N_3575,N_1730);
and U4306 (N_4306,N_2007,N_1497);
nand U4307 (N_4307,N_2146,N_384);
nor U4308 (N_4308,N_3686,N_2695);
and U4309 (N_4309,N_1915,N_675);
or U4310 (N_4310,N_568,N_1204);
and U4311 (N_4311,N_1916,N_546);
or U4312 (N_4312,N_128,N_490);
nor U4313 (N_4313,N_1927,N_2024);
and U4314 (N_4314,N_3147,N_2323);
nor U4315 (N_4315,N_1425,N_414);
nor U4316 (N_4316,N_1976,N_2033);
nand U4317 (N_4317,N_3597,N_882);
nor U4318 (N_4318,N_257,N_2556);
nor U4319 (N_4319,N_3768,N_2302);
nand U4320 (N_4320,N_2435,N_1106);
or U4321 (N_4321,N_2971,N_2964);
or U4322 (N_4322,N_998,N_105);
nor U4323 (N_4323,N_1223,N_2220);
and U4324 (N_4324,N_3588,N_3847);
and U4325 (N_4325,N_2876,N_2499);
nor U4326 (N_4326,N_2835,N_592);
nor U4327 (N_4327,N_2573,N_855);
or U4328 (N_4328,N_3971,N_3419);
xor U4329 (N_4329,N_1107,N_1791);
and U4330 (N_4330,N_3249,N_622);
nand U4331 (N_4331,N_1287,N_3777);
or U4332 (N_4332,N_2810,N_2311);
or U4333 (N_4333,N_601,N_3040);
and U4334 (N_4334,N_1891,N_2209);
nor U4335 (N_4335,N_678,N_1520);
xnor U4336 (N_4336,N_2582,N_2726);
xor U4337 (N_4337,N_1137,N_2977);
nor U4338 (N_4338,N_1077,N_313);
nor U4339 (N_4339,N_34,N_2992);
nor U4340 (N_4340,N_2251,N_1552);
nand U4341 (N_4341,N_1575,N_1893);
nor U4342 (N_4342,N_2580,N_2734);
xor U4343 (N_4343,N_1131,N_3418);
and U4344 (N_4344,N_3065,N_1704);
or U4345 (N_4345,N_2020,N_2506);
nor U4346 (N_4346,N_2142,N_2438);
and U4347 (N_4347,N_3165,N_3903);
or U4348 (N_4348,N_2418,N_3762);
and U4349 (N_4349,N_2092,N_2744);
and U4350 (N_4350,N_782,N_595);
xor U4351 (N_4351,N_1764,N_3397);
and U4352 (N_4352,N_3458,N_3051);
nand U4353 (N_4353,N_395,N_2419);
xnor U4354 (N_4354,N_2206,N_2888);
and U4355 (N_4355,N_1218,N_500);
xnor U4356 (N_4356,N_2215,N_3751);
nor U4357 (N_4357,N_51,N_2763);
and U4358 (N_4358,N_3403,N_2255);
nor U4359 (N_4359,N_2878,N_3539);
nand U4360 (N_4360,N_1151,N_3673);
nand U4361 (N_4361,N_3367,N_857);
or U4362 (N_4362,N_3789,N_1377);
nand U4363 (N_4363,N_1169,N_630);
xor U4364 (N_4364,N_1316,N_2997);
nand U4365 (N_4365,N_585,N_3900);
and U4366 (N_4366,N_2249,N_387);
nor U4367 (N_4367,N_969,N_2126);
nor U4368 (N_4368,N_2221,N_1102);
nor U4369 (N_4369,N_201,N_457);
xor U4370 (N_4370,N_537,N_1769);
nand U4371 (N_4371,N_985,N_958);
nand U4372 (N_4372,N_1514,N_1786);
nor U4373 (N_4373,N_3285,N_3175);
nor U4374 (N_4374,N_1043,N_269);
nor U4375 (N_4375,N_2488,N_3520);
xor U4376 (N_4376,N_3337,N_526);
nor U4377 (N_4377,N_2375,N_2242);
and U4378 (N_4378,N_645,N_1090);
nor U4379 (N_4379,N_140,N_2837);
nand U4380 (N_4380,N_899,N_49);
or U4381 (N_4381,N_2153,N_565);
nand U4382 (N_4382,N_3376,N_2022);
nor U4383 (N_4383,N_2520,N_965);
nor U4384 (N_4384,N_2400,N_2864);
nand U4385 (N_4385,N_3430,N_2214);
xnor U4386 (N_4386,N_1110,N_1356);
or U4387 (N_4387,N_2858,N_911);
xor U4388 (N_4388,N_3921,N_955);
nand U4389 (N_4389,N_2697,N_2710);
nor U4390 (N_4390,N_3063,N_435);
nor U4391 (N_4391,N_1422,N_1923);
and U4392 (N_4392,N_2745,N_1533);
nor U4393 (N_4393,N_2371,N_3096);
nor U4394 (N_4394,N_754,N_1314);
or U4395 (N_4395,N_1571,N_679);
and U4396 (N_4396,N_35,N_1614);
nand U4397 (N_4397,N_3917,N_3407);
nor U4398 (N_4398,N_2485,N_1268);
and U4399 (N_4399,N_1247,N_1709);
and U4400 (N_4400,N_3834,N_2462);
or U4401 (N_4401,N_186,N_3423);
and U4402 (N_4402,N_2261,N_260);
xor U4403 (N_4403,N_2679,N_2112);
and U4404 (N_4404,N_2611,N_2771);
nor U4405 (N_4405,N_2437,N_1842);
nor U4406 (N_4406,N_261,N_1957);
or U4407 (N_4407,N_53,N_835);
or U4408 (N_4408,N_33,N_2857);
or U4409 (N_4409,N_3235,N_2752);
nor U4410 (N_4410,N_3927,N_3554);
or U4411 (N_4411,N_554,N_2355);
or U4412 (N_4412,N_3253,N_2150);
or U4413 (N_4413,N_1651,N_454);
or U4414 (N_4414,N_3288,N_1530);
nand U4415 (N_4415,N_2746,N_702);
nand U4416 (N_4416,N_811,N_2196);
nand U4417 (N_4417,N_30,N_2515);
and U4418 (N_4418,N_535,N_787);
and U4419 (N_4419,N_890,N_2811);
and U4420 (N_4420,N_223,N_2337);
or U4421 (N_4421,N_493,N_3779);
and U4422 (N_4422,N_995,N_3355);
or U4423 (N_4423,N_757,N_1860);
or U4424 (N_4424,N_3395,N_1943);
nor U4425 (N_4425,N_858,N_1973);
nor U4426 (N_4426,N_3442,N_1449);
nand U4427 (N_4427,N_2487,N_2591);
and U4428 (N_4428,N_1069,N_37);
xnor U4429 (N_4429,N_3499,N_3904);
nand U4430 (N_4430,N_2,N_2576);
xor U4431 (N_4431,N_705,N_2955);
nand U4432 (N_4432,N_2935,N_2304);
nand U4433 (N_4433,N_129,N_3506);
nand U4434 (N_4434,N_2560,N_3088);
and U4435 (N_4435,N_2276,N_2808);
nor U4436 (N_4436,N_1222,N_3972);
or U4437 (N_4437,N_2152,N_709);
nor U4438 (N_4438,N_2845,N_991);
and U4439 (N_4439,N_3189,N_683);
nand U4440 (N_4440,N_3813,N_1003);
or U4441 (N_4441,N_1450,N_2353);
nand U4442 (N_4442,N_2257,N_1158);
xor U4443 (N_4443,N_3202,N_2227);
or U4444 (N_4444,N_2795,N_1056);
nand U4445 (N_4445,N_363,N_2931);
or U4446 (N_4446,N_1277,N_2890);
xnor U4447 (N_4447,N_1816,N_3966);
or U4448 (N_4448,N_1605,N_5);
nand U4449 (N_4449,N_2350,N_902);
or U4450 (N_4450,N_779,N_564);
or U4451 (N_4451,N_778,N_332);
or U4452 (N_4452,N_2607,N_2444);
and U4453 (N_4453,N_2642,N_2757);
or U4454 (N_4454,N_3605,N_3431);
and U4455 (N_4455,N_2842,N_2238);
or U4456 (N_4456,N_3970,N_321);
and U4457 (N_4457,N_642,N_1962);
nor U4458 (N_4458,N_1458,N_2574);
xor U4459 (N_4459,N_1954,N_2330);
nand U4460 (N_4460,N_479,N_3838);
and U4461 (N_4461,N_2800,N_422);
or U4462 (N_4462,N_735,N_3700);
or U4463 (N_4463,N_923,N_1909);
nor U4464 (N_4464,N_864,N_233);
nand U4465 (N_4465,N_2184,N_2457);
or U4466 (N_4466,N_876,N_1931);
nor U4467 (N_4467,N_2707,N_3238);
nor U4468 (N_4468,N_55,N_1213);
and U4469 (N_4469,N_1862,N_3025);
nand U4470 (N_4470,N_336,N_2034);
or U4471 (N_4471,N_3745,N_1228);
xor U4472 (N_4472,N_2822,N_1760);
nor U4473 (N_4473,N_3726,N_1418);
nand U4474 (N_4474,N_3016,N_3642);
and U4475 (N_4475,N_207,N_2840);
or U4476 (N_4476,N_2412,N_2053);
and U4477 (N_4477,N_1400,N_518);
nand U4478 (N_4478,N_2066,N_1534);
xnor U4479 (N_4479,N_3608,N_1523);
nor U4480 (N_4480,N_2815,N_57);
xnor U4481 (N_4481,N_3634,N_3392);
nand U4482 (N_4482,N_1535,N_1011);
nor U4483 (N_4483,N_3872,N_3448);
xnor U4484 (N_4484,N_2898,N_2751);
and U4485 (N_4485,N_48,N_3001);
and U4486 (N_4486,N_2778,N_497);
nor U4487 (N_4487,N_3037,N_3734);
nor U4488 (N_4488,N_694,N_3998);
xnor U4489 (N_4489,N_3578,N_967);
and U4490 (N_4490,N_87,N_3100);
nand U4491 (N_4491,N_3766,N_230);
nor U4492 (N_4492,N_1910,N_1671);
xor U4493 (N_4493,N_3819,N_2723);
and U4494 (N_4494,N_1889,N_370);
or U4495 (N_4495,N_58,N_2999);
nand U4496 (N_4496,N_1225,N_459);
or U4497 (N_4497,N_220,N_3305);
or U4498 (N_4498,N_2370,N_1516);
xnor U4499 (N_4499,N_3737,N_3286);
and U4500 (N_4500,N_3552,N_901);
or U4501 (N_4501,N_178,N_2615);
nor U4502 (N_4502,N_418,N_549);
nand U4503 (N_4503,N_2956,N_3997);
nand U4504 (N_4504,N_1785,N_139);
or U4505 (N_4505,N_1800,N_951);
nand U4506 (N_4506,N_2941,N_3647);
nand U4507 (N_4507,N_1147,N_1866);
nor U4508 (N_4508,N_2571,N_1724);
xnor U4509 (N_4509,N_3466,N_42);
xnor U4510 (N_4510,N_146,N_307);
or U4511 (N_4511,N_2159,N_1749);
and U4512 (N_4512,N_1068,N_1455);
or U4513 (N_4513,N_3300,N_2510);
and U4514 (N_4514,N_3674,N_2634);
xnor U4515 (N_4515,N_3297,N_3556);
or U4516 (N_4516,N_2902,N_262);
nor U4517 (N_4517,N_3410,N_802);
nor U4518 (N_4518,N_391,N_1710);
and U4519 (N_4519,N_3627,N_1047);
or U4520 (N_4520,N_1156,N_1485);
or U4521 (N_4521,N_2266,N_438);
and U4522 (N_4522,N_1917,N_2782);
xnor U4523 (N_4523,N_3885,N_713);
nand U4524 (N_4524,N_108,N_1340);
xnor U4525 (N_4525,N_250,N_2677);
nand U4526 (N_4526,N_1237,N_530);
or U4527 (N_4527,N_3255,N_3363);
and U4528 (N_4528,N_1977,N_2937);
or U4529 (N_4529,N_1507,N_3594);
nor U4530 (N_4530,N_1459,N_3236);
and U4531 (N_4531,N_1032,N_1933);
nand U4532 (N_4532,N_2868,N_2151);
or U4533 (N_4533,N_2861,N_3151);
or U4534 (N_4534,N_2421,N_3184);
nor U4535 (N_4535,N_3064,N_281);
nor U4536 (N_4536,N_1637,N_2838);
or U4537 (N_4537,N_3713,N_89);
nor U4538 (N_4538,N_401,N_1668);
or U4539 (N_4539,N_2183,N_3931);
nand U4540 (N_4540,N_3260,N_949);
or U4541 (N_4541,N_3465,N_2541);
and U4542 (N_4542,N_3891,N_1150);
nor U4543 (N_4543,N_2601,N_3501);
nor U4544 (N_4544,N_2851,N_2717);
or U4545 (N_4545,N_465,N_21);
and U4546 (N_4546,N_2777,N_570);
or U4547 (N_4547,N_3488,N_3865);
or U4548 (N_4548,N_184,N_2569);
nor U4549 (N_4549,N_1825,N_1366);
xor U4550 (N_4550,N_3003,N_3262);
nor U4551 (N_4551,N_670,N_1285);
and U4552 (N_4552,N_2603,N_2903);
or U4553 (N_4553,N_2383,N_2274);
nor U4554 (N_4554,N_1031,N_3538);
and U4555 (N_4555,N_177,N_95);
nand U4556 (N_4556,N_1841,N_3933);
nor U4557 (N_4557,N_780,N_2430);
nor U4558 (N_4558,N_2789,N_1239);
and U4559 (N_4559,N_3648,N_587);
nor U4560 (N_4560,N_329,N_79);
or U4561 (N_4561,N_3533,N_2176);
and U4562 (N_4562,N_1580,N_1051);
xor U4563 (N_4563,N_676,N_1330);
nor U4564 (N_4564,N_2532,N_1369);
nor U4565 (N_4565,N_3185,N_555);
nor U4566 (N_4566,N_2831,N_1804);
nor U4567 (N_4567,N_2568,N_1140);
and U4568 (N_4568,N_279,N_1928);
xor U4569 (N_4569,N_453,N_1058);
xnor U4570 (N_4570,N_1867,N_2008);
nor U4571 (N_4571,N_3250,N_2381);
xor U4572 (N_4572,N_1787,N_3615);
nand U4573 (N_4573,N_3960,N_2637);
nand U4574 (N_4574,N_1610,N_289);
or U4575 (N_4575,N_2630,N_3541);
or U4576 (N_4576,N_1517,N_1863);
and U4577 (N_4577,N_664,N_155);
nor U4578 (N_4578,N_2417,N_3210);
xnor U4579 (N_4579,N_3172,N_954);
and U4580 (N_4580,N_3490,N_814);
nand U4581 (N_4581,N_1375,N_2252);
and U4582 (N_4582,N_924,N_505);
and U4583 (N_4583,N_2513,N_2640);
nor U4584 (N_4584,N_1858,N_926);
xnor U4585 (N_4585,N_2508,N_1365);
and U4586 (N_4586,N_1772,N_2540);
nor U4587 (N_4587,N_3167,N_1208);
nor U4588 (N_4588,N_2960,N_710);
or U4589 (N_4589,N_1898,N_813);
nor U4590 (N_4590,N_3266,N_3542);
and U4591 (N_4591,N_433,N_2564);
nor U4592 (N_4592,N_1104,N_2040);
or U4593 (N_4593,N_2975,N_1971);
and U4594 (N_4594,N_3089,N_3659);
and U4595 (N_4595,N_3144,N_3206);
nor U4596 (N_4596,N_3156,N_132);
or U4597 (N_4597,N_3637,N_1792);
or U4598 (N_4598,N_1161,N_2889);
nand U4599 (N_4599,N_406,N_3180);
nand U4600 (N_4600,N_2916,N_832);
and U4601 (N_4601,N_3389,N_1220);
or U4602 (N_4602,N_2894,N_613);
nand U4603 (N_4603,N_1376,N_3388);
nor U4604 (N_4604,N_2736,N_81);
and U4605 (N_4605,N_3304,N_1834);
or U4606 (N_4606,N_1326,N_2285);
and U4607 (N_4607,N_1593,N_1896);
xnor U4608 (N_4608,N_3540,N_880);
nand U4609 (N_4609,N_3830,N_1947);
xor U4610 (N_4610,N_182,N_3441);
nand U4611 (N_4611,N_1991,N_1348);
and U4612 (N_4612,N_1443,N_1888);
or U4613 (N_4613,N_3586,N_543);
or U4614 (N_4614,N_1775,N_503);
and U4615 (N_4615,N_352,N_3110);
and U4616 (N_4616,N_1687,N_3243);
nand U4617 (N_4617,N_2368,N_2256);
or U4618 (N_4618,N_3952,N_2846);
nand U4619 (N_4619,N_3320,N_3444);
or U4620 (N_4620,N_2753,N_1656);
and U4621 (N_4621,N_2241,N_2748);
nand U4622 (N_4622,N_2125,N_1255);
and U4623 (N_4623,N_1629,N_1611);
nor U4624 (N_4624,N_3798,N_599);
and U4625 (N_4625,N_3224,N_3005);
or U4626 (N_4626,N_2289,N_88);
nand U4627 (N_4627,N_2676,N_3030);
or U4628 (N_4628,N_3894,N_2624);
and U4629 (N_4629,N_866,N_3564);
nor U4630 (N_4630,N_1600,N_3190);
and U4631 (N_4631,N_3242,N_3118);
nand U4632 (N_4632,N_1324,N_3254);
xnor U4633 (N_4633,N_2058,N_1829);
nor U4634 (N_4634,N_1819,N_121);
nor U4635 (N_4635,N_175,N_3433);
nor U4636 (N_4636,N_930,N_1735);
nand U4637 (N_4637,N_181,N_1334);
nor U4638 (N_4638,N_3169,N_2155);
nor U4639 (N_4639,N_1674,N_3784);
nor U4640 (N_4640,N_1693,N_1329);
xor U4641 (N_4641,N_36,N_1529);
nand U4642 (N_4642,N_3662,N_1682);
nor U4643 (N_4643,N_75,N_1463);
nand U4644 (N_4644,N_2600,N_109);
nand U4645 (N_4645,N_3962,N_1993);
nand U4646 (N_4646,N_2277,N_3617);
nand U4647 (N_4647,N_452,N_960);
nor U4648 (N_4648,N_2985,N_1054);
and U4649 (N_4649,N_3125,N_409);
xnor U4650 (N_4650,N_1952,N_2012);
nand U4651 (N_4651,N_1824,N_2095);
xnor U4652 (N_4652,N_3812,N_1722);
and U4653 (N_4653,N_3711,N_3770);
nor U4654 (N_4654,N_229,N_243);
nor U4655 (N_4655,N_71,N_812);
or U4656 (N_4656,N_997,N_1388);
and U4657 (N_4657,N_1541,N_2659);
and U4658 (N_4658,N_1480,N_878);
and U4659 (N_4659,N_2993,N_3019);
and U4660 (N_4660,N_441,N_753);
nand U4661 (N_4661,N_917,N_936);
nor U4662 (N_4662,N_1644,N_2635);
nor U4663 (N_4663,N_848,N_2714);
nor U4664 (N_4664,N_3233,N_2464);
or U4665 (N_4665,N_3755,N_3623);
xor U4666 (N_4666,N_2456,N_946);
nor U4667 (N_4667,N_1813,N_54);
xor U4668 (N_4668,N_3702,N_344);
nor U4669 (N_4669,N_3806,N_3644);
nor U4670 (N_4670,N_746,N_978);
nand U4671 (N_4671,N_820,N_3369);
and U4672 (N_4672,N_3307,N_3055);
or U4673 (N_4673,N_2299,N_1856);
nand U4674 (N_4674,N_1920,N_305);
and U4675 (N_4675,N_2048,N_3512);
nor U4676 (N_4676,N_2850,N_1951);
nand U4677 (N_4677,N_3691,N_2127);
nand U4678 (N_4678,N_2388,N_1186);
nor U4679 (N_4679,N_3362,N_3119);
and U4680 (N_4680,N_2078,N_3602);
and U4681 (N_4681,N_206,N_474);
or U4682 (N_4682,N_2397,N_156);
nand U4683 (N_4683,N_1194,N_1323);
nand U4684 (N_4684,N_2798,N_784);
xnor U4685 (N_4685,N_3866,N_2604);
nand U4686 (N_4686,N_663,N_1428);
xnor U4687 (N_4687,N_809,N_1846);
and U4688 (N_4688,N_3939,N_3340);
nor U4689 (N_4689,N_3148,N_2059);
nor U4690 (N_4690,N_3529,N_1242);
or U4691 (N_4691,N_1759,N_63);
nand U4692 (N_4692,N_1788,N_1604);
nor U4693 (N_4693,N_3975,N_3521);
or U4694 (N_4694,N_1590,N_2501);
xor U4695 (N_4695,N_3111,N_1584);
nand U4696 (N_4696,N_547,N_1120);
and U4697 (N_4697,N_699,N_193);
nor U4698 (N_4698,N_1802,N_2413);
nand U4699 (N_4699,N_3328,N_286);
and U4700 (N_4700,N_76,N_94);
nor U4701 (N_4701,N_715,N_2770);
or U4702 (N_4702,N_703,N_1945);
nand U4703 (N_4703,N_2727,N_2836);
nand U4704 (N_4704,N_2530,N_2447);
and U4705 (N_4705,N_2466,N_3326);
or U4706 (N_4706,N_655,N_2722);
nor U4707 (N_4707,N_1148,N_649);
or U4708 (N_4708,N_2551,N_2667);
and U4709 (N_4709,N_3467,N_684);
or U4710 (N_4710,N_431,N_701);
or U4711 (N_4711,N_1112,N_3778);
nor U4712 (N_4712,N_1317,N_3825);
xnor U4713 (N_4713,N_2879,N_2672);
nor U4714 (N_4714,N_1880,N_7);
or U4715 (N_4715,N_483,N_2295);
nor U4716 (N_4716,N_3681,N_2598);
nor U4717 (N_4717,N_1965,N_1873);
and U4718 (N_4718,N_2199,N_3414);
nor U4719 (N_4719,N_8,N_3502);
nor U4720 (N_4720,N_952,N_2019);
nand U4721 (N_4721,N_2526,N_513);
nand U4722 (N_4722,N_3171,N_2170);
nor U4723 (N_4723,N_1437,N_2581);
and U4724 (N_4724,N_1423,N_825);
nand U4725 (N_4725,N_1044,N_904);
and U4726 (N_4726,N_3145,N_3849);
or U4727 (N_4727,N_534,N_216);
nor U4728 (N_4728,N_3170,N_1650);
and U4729 (N_4729,N_3988,N_331);
and U4730 (N_4730,N_2774,N_2361);
nand U4731 (N_4731,N_2422,N_2426);
or U4732 (N_4732,N_1964,N_2967);
and U4733 (N_4733,N_1417,N_3387);
nor U4734 (N_4734,N_1946,N_3908);
or U4735 (N_4735,N_3007,N_1447);
or U4736 (N_4736,N_1982,N_3956);
or U4737 (N_4737,N_2531,N_1579);
and U4738 (N_4738,N_1039,N_1207);
nand U4739 (N_4739,N_504,N_3203);
or U4740 (N_4740,N_3469,N_3947);
and U4741 (N_4741,N_2616,N_2737);
nor U4742 (N_4742,N_1490,N_1427);
and U4743 (N_4743,N_2140,N_2652);
or U4744 (N_4744,N_3292,N_3379);
xor U4745 (N_4745,N_118,N_3757);
and U4746 (N_4746,N_3628,N_2904);
nand U4747 (N_4747,N_3081,N_583);
or U4748 (N_4748,N_2262,N_3446);
or U4749 (N_4749,N_2293,N_2790);
nor U4750 (N_4750,N_1307,N_751);
nand U4751 (N_4751,N_2959,N_1662);
or U4752 (N_4752,N_196,N_3887);
xor U4753 (N_4753,N_1621,N_425);
xor U4754 (N_4754,N_3078,N_3102);
xnor U4755 (N_4755,N_2860,N_3168);
and U4756 (N_4756,N_1079,N_3420);
or U4757 (N_4757,N_551,N_2805);
and U4758 (N_4758,N_2719,N_1547);
nor U4759 (N_4759,N_1061,N_1272);
nor U4760 (N_4760,N_2555,N_1410);
or U4761 (N_4761,N_1094,N_2961);
or U4762 (N_4762,N_931,N_1210);
and U4763 (N_4763,N_324,N_3829);
and U4764 (N_4764,N_1370,N_3045);
nor U4765 (N_4765,N_3283,N_1424);
and U4766 (N_4766,N_2284,N_3187);
or U4767 (N_4767,N_627,N_933);
nor U4768 (N_4768,N_1631,N_1098);
nand U4769 (N_4769,N_3701,N_3658);
and U4770 (N_4770,N_2674,N_325);
or U4771 (N_4771,N_3324,N_1890);
nor U4772 (N_4772,N_1981,N_1113);
or U4773 (N_4773,N_982,N_1021);
or U4774 (N_4774,N_2129,N_3246);
xnor U4775 (N_4775,N_643,N_1795);
or U4776 (N_4776,N_1240,N_2534);
and U4777 (N_4777,N_2105,N_3855);
xor U4778 (N_4778,N_1948,N_2869);
or U4779 (N_4779,N_2738,N_1585);
and U4780 (N_4780,N_3274,N_2197);
nor U4781 (N_4781,N_2135,N_1065);
nor U4782 (N_4782,N_355,N_799);
nand U4783 (N_4783,N_1097,N_2944);
and U4784 (N_4784,N_3405,N_2307);
nor U4785 (N_4785,N_3824,N_1914);
nand U4786 (N_4786,N_717,N_354);
and U4787 (N_4787,N_3930,N_1531);
xnor U4788 (N_4788,N_2664,N_1181);
nor U4789 (N_4789,N_147,N_704);
and U4790 (N_4790,N_1386,N_1937);
xnor U4791 (N_4791,N_1167,N_1677);
nor U4792 (N_4792,N_1870,N_2681);
nand U4793 (N_4793,N_837,N_3919);
and U4794 (N_4794,N_2156,N_719);
nor U4795 (N_4795,N_3685,N_3248);
nand U4796 (N_4796,N_2545,N_2405);
and U4797 (N_4797,N_1115,N_3724);
nand U4798 (N_4798,N_2946,N_3213);
or U4799 (N_4799,N_1599,N_3551);
nand U4800 (N_4800,N_817,N_2643);
xor U4801 (N_4801,N_3181,N_2584);
nand U4802 (N_4802,N_1133,N_3668);
or U4803 (N_4803,N_3974,N_1025);
or U4804 (N_4804,N_3760,N_3805);
or U4805 (N_4805,N_3534,N_15);
or U4806 (N_4806,N_944,N_1713);
and U4807 (N_4807,N_1949,N_2002);
and U4808 (N_4808,N_1576,N_795);
and U4809 (N_4809,N_3882,N_1454);
nand U4810 (N_4810,N_3058,N_918);
nand U4811 (N_4811,N_1559,N_2700);
nand U4812 (N_4812,N_604,N_3510);
and U4813 (N_4813,N_3173,N_2395);
nor U4814 (N_4814,N_2163,N_935);
or U4815 (N_4815,N_1059,N_619);
xnor U4816 (N_4816,N_1615,N_2026);
or U4817 (N_4817,N_1953,N_1509);
and U4818 (N_4818,N_99,N_2415);
nor U4819 (N_4819,N_2367,N_2440);
nor U4820 (N_4820,N_919,N_1436);
xnor U4821 (N_4821,N_1469,N_2044);
and U4822 (N_4822,N_3354,N_666);
and U4823 (N_4823,N_3359,N_2083);
nor U4824 (N_4824,N_538,N_3531);
or U4825 (N_4825,N_959,N_1959);
and U4826 (N_4826,N_964,N_3443);
or U4827 (N_4827,N_2505,N_2968);
and U4828 (N_4828,N_2308,N_2363);
nand U4829 (N_4829,N_990,N_3902);
nor U4830 (N_4830,N_1850,N_2099);
and U4831 (N_4831,N_210,N_3727);
nand U4832 (N_4832,N_3264,N_3400);
or U4833 (N_4833,N_3455,N_3626);
or U4834 (N_4834,N_2104,N_690);
xnor U4835 (N_4835,N_897,N_1471);
nor U4836 (N_4836,N_3230,N_1101);
nand U4837 (N_4837,N_1707,N_2021);
nand U4838 (N_4838,N_956,N_69);
or U4839 (N_4839,N_1522,N_1549);
nor U4840 (N_4840,N_3085,N_844);
nand U4841 (N_4841,N_966,N_1036);
and U4842 (N_4842,N_3042,N_638);
nand U4843 (N_4843,N_3155,N_1711);
nor U4844 (N_4844,N_2365,N_843);
or U4845 (N_4845,N_3957,N_3425);
or U4846 (N_4846,N_323,N_1111);
nor U4847 (N_4847,N_2175,N_460);
nor U4848 (N_4848,N_3445,N_2779);
or U4849 (N_4849,N_1551,N_851);
or U4850 (N_4850,N_1905,N_1911);
nor U4851 (N_4851,N_2905,N_972);
nor U4852 (N_4852,N_865,N_1612);
and U4853 (N_4853,N_541,N_2951);
nor U4854 (N_4854,N_1310,N_1777);
nand U4855 (N_4855,N_264,N_3630);
xnor U4856 (N_4856,N_3162,N_135);
nor U4857 (N_4857,N_2210,N_1124);
nor U4858 (N_4858,N_3823,N_2817);
nand U4859 (N_4859,N_1558,N_1636);
and U4860 (N_4860,N_3112,N_806);
or U4861 (N_4861,N_1681,N_3670);
nand U4862 (N_4862,N_2731,N_3229);
or U4863 (N_4863,N_1295,N_2750);
and U4864 (N_4864,N_2651,N_2606);
nor U4865 (N_4865,N_3643,N_3614);
nand U4866 (N_4866,N_3577,N_2594);
nand U4867 (N_4867,N_148,N_3329);
and U4868 (N_4868,N_3289,N_2141);
nand U4869 (N_4869,N_1157,N_840);
and U4870 (N_4870,N_2661,N_330);
or U4871 (N_4871,N_301,N_3950);
or U4872 (N_4872,N_470,N_189);
nand U4873 (N_4873,N_3024,N_1142);
and U4874 (N_4874,N_308,N_62);
nor U4875 (N_4875,N_316,N_3461);
and U4876 (N_4876,N_2553,N_3976);
and U4877 (N_4877,N_3853,N_3240);
or U4878 (N_4878,N_3781,N_2527);
and U4879 (N_4879,N_228,N_3128);
nand U4880 (N_4880,N_2585,N_100);
or U4881 (N_4881,N_2264,N_1188);
or U4882 (N_4882,N_3267,N_2358);
or U4883 (N_4883,N_270,N_1381);
nor U4884 (N_4884,N_2340,N_824);
nand U4885 (N_4885,N_1015,N_3730);
or U4886 (N_4886,N_130,N_2675);
xor U4887 (N_4887,N_2830,N_2883);
nor U4888 (N_4888,N_900,N_1797);
nor U4889 (N_4889,N_1925,N_2620);
nor U4890 (N_4890,N_333,N_769);
nor U4891 (N_4891,N_3398,N_29);
nor U4892 (N_4892,N_3543,N_445);
and U4893 (N_4893,N_3833,N_1227);
nor U4894 (N_4894,N_3375,N_2712);
nor U4895 (N_4895,N_2786,N_1884);
or U4896 (N_4896,N_288,N_120);
nor U4897 (N_4897,N_3782,N_1290);
and U4898 (N_4898,N_733,N_1738);
or U4899 (N_4899,N_2619,N_3481);
and U4900 (N_4900,N_419,N_2202);
or U4901 (N_4901,N_136,N_12);
and U4902 (N_4902,N_1848,N_1193);
nand U4903 (N_4903,N_3356,N_578);
nand U4904 (N_4904,N_1267,N_399);
xnor U4905 (N_4905,N_3046,N_1633);
and U4906 (N_4906,N_1630,N_1897);
or U4907 (N_4907,N_1139,N_3818);
and U4908 (N_4908,N_3484,N_989);
or U4909 (N_4909,N_2108,N_3309);
nor U4910 (N_4910,N_283,N_2226);
or U4911 (N_4911,N_981,N_3869);
or U4912 (N_4912,N_3299,N_2528);
or U4913 (N_4913,N_2909,N_372);
nand U4914 (N_4914,N_1743,N_199);
nand U4915 (N_4915,N_426,N_3791);
and U4916 (N_4916,N_3850,N_473);
nand U4917 (N_4917,N_2766,N_3844);
and U4918 (N_4918,N_3383,N_1202);
nor U4919 (N_4919,N_3652,N_776);
nand U4920 (N_4920,N_1554,N_2613);
nor U4921 (N_4921,N_3990,N_343);
nand U4922 (N_4922,N_285,N_3338);
and U4923 (N_4923,N_558,N_756);
and U4924 (N_4924,N_1669,N_636);
and U4925 (N_4925,N_2186,N_3323);
or U4926 (N_4926,N_2538,N_2915);
nand U4927 (N_4927,N_623,N_2357);
nor U4928 (N_4928,N_2224,N_347);
nand U4929 (N_4929,N_2764,N_563);
and U4930 (N_4930,N_400,N_2704);
nor U4931 (N_4931,N_3107,N_2387);
nor U4932 (N_4932,N_3177,N_3993);
nand U4933 (N_4933,N_3570,N_3029);
xor U4934 (N_4934,N_3163,N_2230);
or U4935 (N_4935,N_383,N_1380);
or U4936 (N_4936,N_3123,N_1877);
or U4937 (N_4937,N_1794,N_1342);
nand U4938 (N_4938,N_1160,N_3485);
nand U4939 (N_4939,N_466,N_2934);
or U4940 (N_4940,N_1881,N_3616);
xnor U4941 (N_4941,N_1499,N_3010);
or U4942 (N_4942,N_2919,N_3725);
xnor U4943 (N_4943,N_2755,N_2627);
and U4944 (N_4944,N_167,N_3708);
and U4945 (N_4945,N_2013,N_2189);
nand U4946 (N_4946,N_180,N_1123);
and U4947 (N_4947,N_1596,N_1099);
nor U4948 (N_4948,N_2546,N_1989);
nor U4949 (N_4949,N_3733,N_2349);
or U4950 (N_4950,N_3339,N_762);
and U4951 (N_4951,N_2076,N_340);
or U4952 (N_4952,N_1518,N_720);
and U4953 (N_4953,N_1657,N_979);
nand U4954 (N_4954,N_1963,N_3817);
and U4955 (N_4955,N_1998,N_1472);
and U4956 (N_4956,N_255,N_3503);
nor U4957 (N_4957,N_3033,N_3696);
and U4958 (N_4958,N_633,N_478);
or U4959 (N_4959,N_170,N_2213);
or U4960 (N_4960,N_2281,N_364);
and U4961 (N_4961,N_2947,N_677);
xnor U4962 (N_4962,N_117,N_1695);
nand U4963 (N_4963,N_3090,N_1752);
nor U4964 (N_4964,N_1372,N_616);
nor U4965 (N_4965,N_3723,N_1303);
or U4966 (N_4966,N_3593,N_1315);
nand U4967 (N_4967,N_2577,N_3483);
or U4968 (N_4968,N_1333,N_1309);
nand U4969 (N_4969,N_22,N_221);
nand U4970 (N_4970,N_614,N_1387);
and U4971 (N_4971,N_617,N_2597);
or U4972 (N_4972,N_553,N_1249);
and U4973 (N_4973,N_2843,N_1080);
or U4974 (N_4974,N_593,N_833);
or U4975 (N_4975,N_2895,N_3139);
or U4976 (N_4976,N_380,N_533);
or U4977 (N_4977,N_1494,N_3973);
nand U4978 (N_4978,N_2854,N_385);
nor U4979 (N_4979,N_1144,N_47);
or U4980 (N_4980,N_2362,N_3839);
nand U4981 (N_4981,N_1231,N_3062);
nand U4982 (N_4982,N_2537,N_3663);
nand U4983 (N_4983,N_2885,N_877);
or U4984 (N_4984,N_20,N_315);
nand U4985 (N_4985,N_2525,N_1812);
and U4986 (N_4986,N_2566,N_2259);
nor U4987 (N_4987,N_271,N_1464);
nor U4988 (N_4988,N_434,N_1705);
and U4989 (N_4989,N_2684,N_566);
and U4990 (N_4990,N_2754,N_3193);
nand U4991 (N_4991,N_144,N_1968);
nor U4992 (N_4992,N_1444,N_3831);
and U4993 (N_4993,N_1919,N_251);
and U4994 (N_4994,N_475,N_2834);
and U4995 (N_4995,N_1810,N_2645);
nand U4996 (N_4996,N_3415,N_1726);
nand U4997 (N_4997,N_2106,N_1430);
or U4998 (N_4998,N_2267,N_412);
or U4999 (N_4999,N_3880,N_2599);
and U5000 (N_5000,N_849,N_3252);
or U5001 (N_5001,N_1975,N_328);
nor U5002 (N_5002,N_1555,N_2896);
and U5003 (N_5003,N_209,N_458);
nor U5004 (N_5004,N_476,N_742);
and U5005 (N_5005,N_763,N_1495);
nand U5006 (N_5006,N_3547,N_174);
and U5007 (N_5007,N_50,N_828);
nor U5008 (N_5008,N_3797,N_2563);
or U5009 (N_5009,N_3191,N_1125);
nor U5010 (N_5010,N_548,N_3892);
or U5011 (N_5011,N_1807,N_1224);
nor U5012 (N_5012,N_52,N_3301);
and U5013 (N_5013,N_1396,N_1403);
nor U5014 (N_5014,N_492,N_818);
or U5015 (N_5015,N_3688,N_1174);
xnor U5016 (N_5016,N_1138,N_3901);
or U5017 (N_5017,N_1421,N_2004);
nor U5018 (N_5018,N_894,N_3138);
and U5019 (N_5019,N_3565,N_706);
or U5020 (N_5020,N_1071,N_1527);
or U5021 (N_5021,N_2119,N_3807);
nor U5022 (N_5022,N_1364,N_1561);
xnor U5023 (N_5023,N_1510,N_291);
or U5024 (N_5024,N_1608,N_3684);
xor U5025 (N_5025,N_3940,N_2512);
nand U5026 (N_5026,N_1694,N_2160);
nand U5027 (N_5027,N_1251,N_2586);
and U5028 (N_5028,N_3943,N_3438);
nor U5029 (N_5029,N_1085,N_1143);
xor U5030 (N_5030,N_1540,N_2966);
nor U5031 (N_5031,N_159,N_1345);
nand U5032 (N_5032,N_940,N_1357);
xnor U5033 (N_5033,N_667,N_559);
or U5034 (N_5034,N_2509,N_687);
or U5035 (N_5035,N_1941,N_1020);
and U5036 (N_5036,N_1776,N_218);
or U5037 (N_5037,N_1688,N_3474);
nor U5038 (N_5038,N_1205,N_796);
and U5039 (N_5039,N_2602,N_1496);
nor U5040 (N_5040,N_3076,N_3857);
nor U5041 (N_5041,N_3028,N_1885);
nand U5042 (N_5042,N_1836,N_3460);
or U5043 (N_5043,N_915,N_1320);
xnor U5044 (N_5044,N_1371,N_2148);
or U5045 (N_5045,N_1771,N_411);
or U5046 (N_5046,N_143,N_2103);
or U5047 (N_5047,N_3536,N_3624);
and U5048 (N_5048,N_691,N_605);
xnor U5049 (N_5049,N_1505,N_1128);
nor U5050 (N_5050,N_2949,N_1512);
nor U5051 (N_5051,N_495,N_1426);
nor U5052 (N_5052,N_1996,N_3332);
and U5053 (N_5053,N_3764,N_521);
and U5054 (N_5054,N_2145,N_217);
nand U5055 (N_5055,N_1155,N_524);
nor U5056 (N_5056,N_2547,N_3790);
nor U5057 (N_5057,N_2341,N_2194);
nand U5058 (N_5058,N_2235,N_3476);
nand U5059 (N_5059,N_3934,N_1838);
nand U5060 (N_5060,N_3920,N_1159);
nand U5061 (N_5061,N_2721,N_3130);
nand U5062 (N_5062,N_2862,N_3272);
nor U5063 (N_5063,N_1587,N_2443);
or U5064 (N_5064,N_1232,N_2706);
and U5065 (N_5065,N_1659,N_920);
and U5066 (N_5066,N_3742,N_1474);
nor U5067 (N_5067,N_2877,N_2802);
or U5068 (N_5068,N_3963,N_367);
and U5069 (N_5069,N_3293,N_2410);
nor U5070 (N_5070,N_2923,N_2943);
and U5071 (N_5071,N_1515,N_1243);
nand U5072 (N_5072,N_846,N_3072);
or U5073 (N_5073,N_639,N_2394);
xnor U5074 (N_5074,N_3131,N_2918);
or U5075 (N_5075,N_472,N_1501);
nand U5076 (N_5076,N_1129,N_845);
or U5077 (N_5077,N_2486,N_2280);
nand U5078 (N_5078,N_3767,N_3316);
nand U5079 (N_5079,N_669,N_3516);
or U5080 (N_5080,N_2110,N_1481);
nor U5081 (N_5081,N_3945,N_3826);
nor U5082 (N_5082,N_3666,N_2335);
nor U5083 (N_5083,N_3965,N_3689);
or U5084 (N_5084,N_1557,N_2969);
nor U5085 (N_5085,N_2182,N_2872);
and U5086 (N_5086,N_2986,N_3548);
xor U5087 (N_5087,N_3424,N_3549);
and U5088 (N_5088,N_3006,N_1853);
and U5089 (N_5089,N_3188,N_1184);
nand U5090 (N_5090,N_2161,N_525);
or U5091 (N_5091,N_2767,N_3710);
or U5092 (N_5092,N_300,N_1748);
and U5093 (N_5093,N_2649,N_562);
and U5094 (N_5094,N_1367,N_2998);
or U5095 (N_5095,N_2187,N_3084);
xnor U5096 (N_5096,N_1234,N_3704);
or U5097 (N_5097,N_3583,N_3296);
nand U5098 (N_5098,N_202,N_1511);
xor U5099 (N_5099,N_577,N_267);
and U5100 (N_5100,N_1983,N_511);
and U5101 (N_5101,N_2741,N_3774);
nor U5102 (N_5102,N_3740,N_3703);
nor U5103 (N_5103,N_3948,N_2011);
xnor U5104 (N_5104,N_2558,N_1803);
or U5105 (N_5105,N_3582,N_3018);
or U5106 (N_5106,N_1997,N_624);
nor U5107 (N_5107,N_1350,N_1279);
or U5108 (N_5108,N_1286,N_2686);
or U5109 (N_5109,N_1203,N_1736);
or U5110 (N_5110,N_1894,N_3066);
or U5111 (N_5111,N_3017,N_1456);
nor U5112 (N_5112,N_1010,N_1165);
and U5113 (N_5113,N_1740,N_1543);
and U5114 (N_5114,N_3287,N_3378);
or U5115 (N_5115,N_3409,N_394);
or U5116 (N_5116,N_922,N_1747);
nand U5117 (N_5117,N_1434,N_1550);
nor U5118 (N_5118,N_3846,N_921);
or U5119 (N_5119,N_3992,N_1994);
and U5120 (N_5120,N_2933,N_3034);
and U5121 (N_5121,N_2865,N_962);
or U5122 (N_5122,N_496,N_173);
xor U5123 (N_5123,N_3985,N_1956);
and U5124 (N_5124,N_3122,N_1715);
nand U5125 (N_5125,N_3886,N_1597);
nor U5126 (N_5126,N_750,N_2069);
nor U5127 (N_5127,N_176,N_654);
xor U5128 (N_5128,N_943,N_2650);
or U5129 (N_5129,N_115,N_1346);
nand U5130 (N_5130,N_560,N_3728);
or U5131 (N_5131,N_1339,N_3883);
nand U5132 (N_5132,N_2638,N_1332);
nor U5133 (N_5133,N_3497,N_2298);
nor U5134 (N_5134,N_3721,N_3926);
nand U5135 (N_5135,N_273,N_2332);
and U5136 (N_5136,N_3537,N_1658);
and U5137 (N_5137,N_1491,N_1831);
and U5138 (N_5138,N_3944,N_2091);
and U5139 (N_5139,N_1179,N_24);
nor U5140 (N_5140,N_1706,N_3911);
nor U5141 (N_5141,N_3211,N_941);
or U5142 (N_5142,N_2165,N_3604);
nand U5143 (N_5143,N_2333,N_1603);
nor U5144 (N_5144,N_1409,N_3893);
and U5145 (N_5145,N_2134,N_608);
and U5146 (N_5146,N_3199,N_3747);
nor U5147 (N_5147,N_540,N_2639);
and U5148 (N_5148,N_1359,N_1868);
nand U5149 (N_5149,N_2420,N_2781);
xnor U5150 (N_5150,N_1008,N_2819);
and U5151 (N_5151,N_1035,N_572);
nand U5152 (N_5152,N_1569,N_3217);
nand U5153 (N_5153,N_1944,N_3002);
nor U5154 (N_5154,N_3428,N_2446);
nand U5155 (N_5155,N_1465,N_461);
or U5156 (N_5156,N_1586,N_1399);
and U5157 (N_5157,N_2472,N_2716);
or U5158 (N_5158,N_620,N_377);
nor U5159 (N_5159,N_1265,N_1328);
nor U5160 (N_5160,N_3408,N_3319);
nand U5161 (N_5161,N_1302,N_3858);
nor U5162 (N_5162,N_2386,N_1617);
nor U5163 (N_5163,N_10,N_908);
nor U5164 (N_5164,N_588,N_2498);
xor U5165 (N_5165,N_3015,N_3526);
and U5166 (N_5166,N_2588,N_3736);
nand U5167 (N_5167,N_353,N_2046);
or U5168 (N_5168,N_2913,N_2407);
or U5169 (N_5169,N_161,N_957);
nor U5170 (N_5170,N_3454,N_397);
nor U5171 (N_5171,N_3047,N_3935);
and U5172 (N_5172,N_660,N_25);
or U5173 (N_5173,N_2917,N_2473);
nor U5174 (N_5174,N_2735,N_1040);
or U5175 (N_5175,N_3996,N_1990);
or U5176 (N_5176,N_1720,N_3174);
and U5177 (N_5177,N_1446,N_2177);
and U5178 (N_5178,N_3598,N_3683);
nor U5179 (N_5179,N_2812,N_3695);
nor U5180 (N_5180,N_3792,N_600);
or U5181 (N_5181,N_3808,N_651);
and U5182 (N_5182,N_9,N_3553);
or U5183 (N_5183,N_3278,N_3995);
nand U5184 (N_5184,N_2204,N_1055);
nor U5185 (N_5185,N_2208,N_2343);
xnor U5186 (N_5186,N_672,N_2167);
nand U5187 (N_5187,N_2174,N_1700);
and U5188 (N_5188,N_423,N_3519);
and U5189 (N_5189,N_2436,N_3014);
nand U5190 (N_5190,N_284,N_3325);
or U5191 (N_5191,N_2450,N_2942);
xor U5192 (N_5192,N_1411,N_2321);
and U5193 (N_5193,N_2028,N_1805);
and U5194 (N_5194,N_183,N_3729);
and U5195 (N_5195,N_3655,N_2936);
nor U5196 (N_5196,N_246,N_3558);
nand U5197 (N_5197,N_2331,N_1500);
and U5198 (N_5198,N_514,N_3550);
and U5199 (N_5199,N_157,N_1808);
or U5200 (N_5200,N_3509,N_1609);
nor U5201 (N_5201,N_249,N_2198);
nor U5202 (N_5202,N_2912,N_2813);
and U5203 (N_5203,N_2117,N_968);
or U5204 (N_5204,N_887,N_3103);
and U5205 (N_5205,N_512,N_950);
nor U5206 (N_5206,N_2618,N_914);
or U5207 (N_5207,N_2926,N_2625);
nor U5208 (N_5208,N_172,N_2314);
nand U5209 (N_5209,N_2849,N_2096);
nor U5210 (N_5210,N_2409,N_3915);
nand U5211 (N_5211,N_1263,N_621);
nand U5212 (N_5212,N_788,N_1233);
nand U5213 (N_5213,N_1814,N_3675);
nor U5214 (N_5214,N_1864,N_3192);
nor U5215 (N_5215,N_2258,N_581);
or U5216 (N_5216,N_2658,N_1081);
or U5217 (N_5217,N_2089,N_3715);
nand U5218 (N_5218,N_3822,N_2544);
nor U5219 (N_5219,N_992,N_791);
and U5220 (N_5220,N_1930,N_92);
nand U5221 (N_5221,N_1661,N_345);
xnor U5222 (N_5222,N_2027,N_3910);
or U5223 (N_5223,N_1273,N_932);
or U5224 (N_5224,N_296,N_2939);
or U5225 (N_5225,N_2666,N_2671);
or U5226 (N_5226,N_659,N_3579);
and U5227 (N_5227,N_3845,N_1921);
or U5228 (N_5228,N_1934,N_3938);
nand U5229 (N_5229,N_3067,N_3786);
and U5230 (N_5230,N_127,N_1670);
or U5231 (N_5231,N_3690,N_1641);
and U5232 (N_5232,N_929,N_2278);
or U5233 (N_5233,N_3345,N_3676);
xor U5234 (N_5234,N_2559,N_2149);
nor U5235 (N_5235,N_2389,N_2239);
nor U5236 (N_5236,N_1195,N_2612);
xor U5237 (N_5237,N_1723,N_3);
nand U5238 (N_5238,N_1211,N_1746);
nand U5239 (N_5239,N_2205,N_1017);
nand U5240 (N_5240,N_2373,N_1702);
or U5241 (N_5241,N_590,N_1275);
and U5242 (N_5242,N_977,N_299);
nand U5243 (N_5243,N_1262,N_349);
or U5244 (N_5244,N_1433,N_3884);
nand U5245 (N_5245,N_1078,N_3178);
and U5246 (N_5246,N_2761,N_2590);
nand U5247 (N_5247,N_3955,N_3487);
nand U5248 (N_5248,N_646,N_3671);
and U5249 (N_5249,N_1525,N_3330);
nand U5250 (N_5250,N_2806,N_3219);
nand U5251 (N_5251,N_942,N_586);
and U5252 (N_5252,N_862,N_1006);
or U5253 (N_5253,N_1470,N_98);
nor U5254 (N_5254,N_3095,N_3141);
or U5255 (N_5255,N_3158,N_1685);
or U5256 (N_5256,N_1851,N_3810);
or U5257 (N_5257,N_3561,N_3743);
xnor U5258 (N_5258,N_64,N_3633);
nand U5259 (N_5259,N_2139,N_2052);
nand U5260 (N_5260,N_1248,N_910);
and U5261 (N_5261,N_693,N_2391);
and U5262 (N_5262,N_994,N_3099);
nor U5263 (N_5263,N_569,N_628);
or U5264 (N_5264,N_2317,N_2245);
or U5265 (N_5265,N_2432,N_382);
or U5266 (N_5266,N_2061,N_3731);
nand U5267 (N_5267,N_2983,N_3094);
and U5268 (N_5268,N_3342,N_739);
nor U5269 (N_5269,N_2441,N_3978);
or U5270 (N_5270,N_1645,N_2470);
or U5271 (N_5271,N_3436,N_1773);
and U5272 (N_5272,N_1300,N_482);
nor U5273 (N_5273,N_3750,N_2401);
and U5274 (N_5274,N_785,N_2172);
or U5275 (N_5275,N_2796,N_653);
nand U5276 (N_5276,N_160,N_1374);
nand U5277 (N_5277,N_3946,N_896);
or U5278 (N_5278,N_3716,N_1462);
xnor U5279 (N_5279,N_2517,N_1780);
nand U5280 (N_5280,N_310,N_2039);
xnor U5281 (N_5281,N_3632,N_3610);
nand U5282 (N_5282,N_3748,N_2718);
and U5283 (N_5283,N_2054,N_3276);
nor U5284 (N_5284,N_241,N_1121);
nand U5285 (N_5285,N_198,N_871);
and U5286 (N_5286,N_440,N_2448);
nand U5287 (N_5287,N_2359,N_3772);
or U5288 (N_5288,N_2399,N_44);
nand U5289 (N_5289,N_2392,N_3693);
nor U5290 (N_5290,N_306,N_3358);
and U5291 (N_5291,N_2157,N_3739);
nand U5292 (N_5292,N_545,N_1221);
or U5293 (N_5293,N_625,N_2338);
and U5294 (N_5294,N_1666,N_1442);
nand U5295 (N_5295,N_134,N_334);
nand U5296 (N_5296,N_1513,N_3080);
and U5297 (N_5297,N_1901,N_211);
or U5298 (N_5298,N_2463,N_1358);
and U5299 (N_5299,N_2067,N_948);
and U5300 (N_5300,N_2788,N_3494);
nor U5301 (N_5301,N_3259,N_2908);
nor U5302 (N_5302,N_1583,N_3113);
and U5303 (N_5303,N_2692,N_1642);
nand U5304 (N_5304,N_1519,N_3687);
and U5305 (N_5305,N_1070,N_3936);
or U5306 (N_5306,N_3093,N_439);
nor U5307 (N_5307,N_2377,N_82);
or U5308 (N_5308,N_3473,N_3153);
nand U5309 (N_5309,N_1728,N_1005);
xor U5310 (N_5310,N_2631,N_3247);
nor U5311 (N_5311,N_3198,N_102);
nor U5312 (N_5312,N_116,N_2708);
nor U5313 (N_5313,N_1498,N_96);
nand U5314 (N_5314,N_421,N_2921);
nand U5315 (N_5315,N_1172,N_3074);
or U5316 (N_5316,N_1363,N_1649);
and U5317 (N_5317,N_3843,N_392);
or U5318 (N_5318,N_3515,N_3606);
and U5319 (N_5319,N_937,N_450);
or U5320 (N_5320,N_417,N_854);
and U5321 (N_5321,N_2833,N_1402);
and U5322 (N_5322,N_3318,N_2287);
and U5323 (N_5323,N_2928,N_3384);
nand U5324 (N_5324,N_3638,N_3937);
nand U5325 (N_5325,N_3225,N_67);
or U5326 (N_5326,N_1811,N_1936);
nand U5327 (N_5327,N_3528,N_3545);
and U5328 (N_5328,N_2379,N_428);
or U5329 (N_5329,N_1397,N_1758);
or U5330 (N_5330,N_3761,N_3555);
and U5331 (N_5331,N_2390,N_1152);
or U5332 (N_5332,N_2552,N_2166);
nand U5333 (N_5333,N_1260,N_3719);
and U5334 (N_5334,N_1254,N_1153);
nand U5335 (N_5335,N_611,N_2641);
or U5336 (N_5336,N_2253,N_697);
nand U5337 (N_5337,N_3273,N_2360);
nand U5338 (N_5338,N_3204,N_72);
and U5339 (N_5339,N_137,N_2015);
xor U5340 (N_5340,N_1354,N_3796);
nand U5341 (N_5341,N_607,N_1745);
nand U5342 (N_5342,N_2064,N_208);
nor U5343 (N_5343,N_2246,N_875);
xor U5344 (N_5344,N_1440,N_3636);
nand U5345 (N_5345,N_3365,N_376);
nor U5346 (N_5346,N_1091,N_165);
and U5347 (N_5347,N_867,N_420);
and U5348 (N_5348,N_1198,N_803);
or U5349 (N_5349,N_1833,N_2953);
and U5350 (N_5350,N_3859,N_3038);
or U5351 (N_5351,N_2272,N_1452);
or U5352 (N_5352,N_2452,N_3105);
nand U5353 (N_5353,N_3788,N_2633);
and U5354 (N_5354,N_3842,N_1132);
or U5355 (N_5355,N_3595,N_3146);
nor U5356 (N_5356,N_1553,N_1539);
nand U5357 (N_5357,N_2518,N_2882);
and U5358 (N_5358,N_2222,N_2691);
nor U5359 (N_5359,N_471,N_1136);
or U5360 (N_5360,N_214,N_1906);
xnor U5361 (N_5361,N_939,N_2617);
and U5362 (N_5362,N_486,N_2747);
and U5363 (N_5363,N_1556,N_3574);
xnor U5364 (N_5364,N_885,N_597);
nand U5365 (N_5365,N_3967,N_2236);
nand U5366 (N_5366,N_1154,N_732);
xor U5367 (N_5367,N_898,N_3041);
nand U5368 (N_5368,N_2107,N_3793);
nand U5369 (N_5369,N_3310,N_3075);
nand U5370 (N_5370,N_999,N_1092);
nand U5371 (N_5371,N_2087,N_1382);
or U5372 (N_5372,N_2881,N_2772);
and U5373 (N_5373,N_2137,N_2938);
nor U5374 (N_5374,N_1216,N_1620);
and U5375 (N_5375,N_3498,N_1684);
nand U5376 (N_5376,N_1281,N_2592);
xor U5377 (N_5377,N_1892,N_2693);
and U5378 (N_5378,N_508,N_416);
nor U5379 (N_5379,N_1532,N_2703);
nor U5380 (N_5380,N_1116,N_2077);
nor U5381 (N_5381,N_1201,N_1191);
nand U5382 (N_5382,N_1475,N_1007);
nand U5383 (N_5383,N_727,N_741);
xor U5384 (N_5384,N_912,N_1026);
and U5385 (N_5385,N_2075,N_2113);
and U5386 (N_5386,N_2839,N_362);
or U5387 (N_5387,N_1861,N_2303);
and U5388 (N_5388,N_1289,N_1236);
nor U5389 (N_5389,N_3386,N_1741);
or U5390 (N_5390,N_3257,N_3984);
and U5391 (N_5391,N_2247,N_631);
xor U5392 (N_5392,N_2911,N_1384);
or U5393 (N_5393,N_1066,N_3877);
nand U5394 (N_5394,N_3371,N_2322);
and U5395 (N_5395,N_1276,N_889);
xnor U5396 (N_5396,N_536,N_3020);
nor U5397 (N_5397,N_1972,N_3873);
nand U5398 (N_5398,N_2043,N_974);
or U5399 (N_5399,N_3214,N_3609);
nor U5400 (N_5400,N_1727,N_2451);
xor U5401 (N_5401,N_2369,N_3514);
or U5402 (N_5402,N_529,N_1114);
or U5403 (N_5403,N_550,N_1351);
and U5404 (N_5404,N_1762,N_276);
or U5405 (N_5405,N_766,N_767);
or U5406 (N_5406,N_2823,N_1461);
nand U5407 (N_5407,N_3140,N_1648);
nor U5408 (N_5408,N_1757,N_2768);
and U5409 (N_5409,N_1562,N_2632);
nor U5410 (N_5410,N_93,N_510);
or U5411 (N_5411,N_759,N_1761);
or U5412 (N_5412,N_3620,N_1486);
or U5413 (N_5413,N_2982,N_1876);
xnor U5414 (N_5414,N_432,N_78);
and U5415 (N_5415,N_169,N_2554);
or U5416 (N_5416,N_2609,N_1269);
nor U5417 (N_5417,N_1809,N_23);
and U5418 (N_5418,N_1084,N_2965);
nor U5419 (N_5419,N_1725,N_2821);
nand U5420 (N_5420,N_3207,N_2589);
nand U5421 (N_5421,N_1331,N_1245);
or U5422 (N_5422,N_1835,N_3895);
nor U5423 (N_5423,N_1560,N_3815);
or U5424 (N_5424,N_3077,N_2453);
nand U5425 (N_5425,N_3133,N_3129);
or U5426 (N_5426,N_1347,N_1404);
nor U5427 (N_5427,N_1526,N_3763);
or U5428 (N_5428,N_1484,N_3463);
and U5429 (N_5429,N_826,N_467);
nor U5430 (N_5430,N_852,N_1770);
nand U5431 (N_5431,N_2511,N_1843);
or U5432 (N_5432,N_3741,N_295);
nor U5433 (N_5433,N_3223,N_2557);
or U5434 (N_5434,N_85,N_2406);
nand U5435 (N_5435,N_1230,N_872);
nand U5436 (N_5436,N_728,N_3159);
nor U5437 (N_5437,N_2031,N_26);
nor U5438 (N_5438,N_1844,N_192);
or U5439 (N_5439,N_1886,N_618);
nand U5440 (N_5440,N_3308,N_1419);
or U5441 (N_5441,N_2325,N_3896);
nor U5442 (N_5442,N_314,N_318);
and U5443 (N_5443,N_164,N_3991);
xor U5444 (N_5444,N_3563,N_1698);
nand U5445 (N_5445,N_2794,N_389);
nor U5446 (N_5446,N_203,N_244);
nor U5447 (N_5447,N_2621,N_1246);
nand U5448 (N_5448,N_2460,N_3907);
nor U5449 (N_5449,N_2101,N_3186);
and U5450 (N_5450,N_191,N_2981);
and U5451 (N_5451,N_2122,N_319);
xor U5452 (N_5452,N_3780,N_673);
and U5453 (N_5453,N_3295,N_2342);
nor U5454 (N_5454,N_1565,N_3591);
nand U5455 (N_5455,N_3412,N_1789);
nor U5456 (N_5456,N_3587,N_1582);
nand U5457 (N_5457,N_1624,N_2442);
or U5458 (N_5458,N_2290,N_2636);
and U5459 (N_5459,N_1504,N_1528);
nor U5460 (N_5460,N_86,N_359);
or U5461 (N_5461,N_2689,N_2315);
and U5462 (N_5462,N_405,N_528);
or U5463 (N_5463,N_131,N_2306);
nand U5464 (N_5464,N_1087,N_3653);
nand U5465 (N_5465,N_1992,N_272);
and U5466 (N_5466,N_1312,N_3500);
and U5467 (N_5467,N_1024,N_2318);
nand U5468 (N_5468,N_1595,N_3060);
or U5469 (N_5469,N_764,N_734);
nand U5470 (N_5470,N_3104,N_3452);
or U5471 (N_5471,N_2100,N_1506);
or U5472 (N_5472,N_1940,N_574);
nor U5473 (N_5473,N_1574,N_612);
nor U5474 (N_5474,N_2060,N_2279);
nor U5475 (N_5475,N_3640,N_1567);
xor U5476 (N_5476,N_2090,N_1908);
nand U5477 (N_5477,N_2207,N_2468);
nand U5478 (N_5478,N_3783,N_3209);
or U5479 (N_5479,N_303,N_2924);
and U5480 (N_5480,N_2482,N_231);
nor U5481 (N_5481,N_1103,N_3981);
nor U5482 (N_5482,N_3803,N_3341);
and U5483 (N_5483,N_3402,N_3905);
xnor U5484 (N_5484,N_2893,N_1686);
nor U5485 (N_5485,N_40,N_1798);
nand U5486 (N_5486,N_358,N_662);
nand U5487 (N_5487,N_3179,N_1733);
nand U5488 (N_5488,N_2240,N_1014);
and U5489 (N_5489,N_3573,N_3101);
nor U5490 (N_5490,N_2870,N_1209);
xnor U5491 (N_5491,N_2396,N_322);
nor U5492 (N_5492,N_2057,N_91);
nor U5493 (N_5493,N_1750,N_3374);
xnor U5494 (N_5494,N_2874,N_3525);
or U5495 (N_5495,N_2382,N_2656);
xnor U5496 (N_5496,N_2561,N_2769);
nor U5497 (N_5497,N_2123,N_2519);
and U5498 (N_5498,N_1383,N_2088);
nand U5499 (N_5499,N_3149,N_913);
and U5500 (N_5500,N_3026,N_1439);
nand U5501 (N_5501,N_1335,N_3048);
and U5502 (N_5502,N_3977,N_378);
nand U5503 (N_5503,N_3396,N_374);
nand U5504 (N_5504,N_3667,N_2372);
and U5505 (N_5505,N_716,N_909);
nand U5506 (N_5506,N_2168,N_3964);
nand U5507 (N_5507,N_194,N_2669);
nand U5508 (N_5508,N_357,N_1053);
and U5509 (N_5509,N_1073,N_2270);
xor U5510 (N_5510,N_3237,N_3336);
and U5511 (N_5511,N_1353,N_2493);
and U5512 (N_5512,N_3380,N_373);
nand U5513 (N_5513,N_891,N_3390);
nand U5514 (N_5514,N_3350,N_6);
nand U5515 (N_5515,N_2940,N_3523);
nand U5516 (N_5516,N_1854,N_3303);
nor U5517 (N_5517,N_522,N_3298);
or U5518 (N_5518,N_1313,N_1134);
and U5519 (N_5519,N_1592,N_1050);
nor U5520 (N_5520,N_3239,N_3776);
and U5521 (N_5521,N_3941,N_1215);
nand U5522 (N_5522,N_2856,N_3897);
or U5523 (N_5523,N_32,N_3660);
xnor U5524 (N_5524,N_2128,N_3036);
and U5525 (N_5525,N_834,N_2855);
nor U5526 (N_5526,N_3241,N_2791);
xor U5527 (N_5527,N_869,N_2516);
and U5528 (N_5528,N_1298,N_480);
nor U5529 (N_5529,N_2115,N_1783);
and U5530 (N_5530,N_3923,N_632);
and U5531 (N_5531,N_2434,N_696);
and U5532 (N_5532,N_737,N_2542);
nand U5533 (N_5533,N_339,N_2016);
or U5534 (N_5534,N_1033,N_892);
nand U5535 (N_5535,N_3468,N_2037);
nor U5536 (N_5536,N_1280,N_1774);
xnor U5537 (N_5537,N_539,N_3650);
nand U5538 (N_5538,N_3518,N_2250);
nor U5539 (N_5539,N_736,N_925);
xor U5540 (N_5540,N_3654,N_366);
and U5541 (N_5541,N_2050,N_1984);
nor U5542 (N_5542,N_2595,N_1127);
and U5543 (N_5543,N_3765,N_396);
nand U5544 (N_5544,N_1170,N_661);
nor U5545 (N_5545,N_2524,N_2962);
nor U5546 (N_5546,N_265,N_2223);
and U5547 (N_5547,N_225,N_1763);
nor U5548 (N_5548,N_1199,N_2605);
and U5549 (N_5549,N_2393,N_775);
nand U5550 (N_5550,N_3368,N_350);
or U5551 (N_5551,N_381,N_1393);
nand U5552 (N_5552,N_2474,N_3746);
and U5553 (N_5553,N_635,N_1613);
or U5554 (N_5554,N_1874,N_1214);
and U5555 (N_5555,N_1083,N_2254);
or U5556 (N_5556,N_2663,N_3271);
nand U5557 (N_5557,N_3391,N_2500);
nand U5558 (N_5558,N_3212,N_3600);
nor U5559 (N_5559,N_2329,N_3852);
xnor U5560 (N_5560,N_3657,N_1392);
and U5561 (N_5561,N_3314,N_3800);
or U5562 (N_5562,N_2668,N_2005);
xnor U5563 (N_5563,N_804,N_3004);
and U5564 (N_5564,N_3011,N_2529);
nand U5565 (N_5565,N_3618,N_74);
nor U5566 (N_5566,N_3035,N_3221);
xor U5567 (N_5567,N_3535,N_2740);
nand U5568 (N_5568,N_1341,N_1521);
or U5569 (N_5569,N_1691,N_1689);
xor U5570 (N_5570,N_3021,N_2758);
nand U5571 (N_5571,N_2489,N_3457);
or U5572 (N_5572,N_3347,N_3759);
nand U5573 (N_5573,N_602,N_2041);
and U5574 (N_5574,N_1652,N_1502);
and U5575 (N_5575,N_1023,N_3692);
and U5576 (N_5576,N_2180,N_674);
nor U5577 (N_5577,N_1732,N_410);
or U5578 (N_5578,N_3769,N_2973);
nand U5579 (N_5579,N_3802,N_292);
nand U5580 (N_5580,N_1030,N_906);
nand U5581 (N_5581,N_606,N_2848);
nand U5582 (N_5582,N_1164,N_1117);
xor U5583 (N_5583,N_1018,N_2503);
and U5584 (N_5584,N_1226,N_3493);
nand U5585 (N_5585,N_1815,N_2292);
nor U5586 (N_5586,N_3527,N_665);
and U5587 (N_5587,N_259,N_2297);
nand U5588 (N_5588,N_2423,N_247);
nand U5589 (N_5589,N_1751,N_2701);
xnor U5590 (N_5590,N_1832,N_154);
nor U5591 (N_5591,N_150,N_2496);
nand U5592 (N_5592,N_280,N_986);
or U5593 (N_5593,N_1979,N_3603);
and U5594 (N_5594,N_3848,N_506);
nor U5595 (N_5595,N_3413,N_2344);
or U5596 (N_5596,N_2829,N_1820);
or U5597 (N_5597,N_1924,N_644);
or U5598 (N_5598,N_2143,N_266);
nor U5599 (N_5599,N_304,N_437);
nand U5600 (N_5600,N_3322,N_1721);
nor U5601 (N_5601,N_2610,N_1985);
nor U5602 (N_5602,N_2042,N_3505);
or U5603 (N_5603,N_1875,N_3876);
xnor U5604 (N_5604,N_2732,N_2987);
and U5605 (N_5605,N_1235,N_3572);
and U5606 (N_5606,N_3517,N_680);
nand U5607 (N_5607,N_576,N_2827);
and U5608 (N_5608,N_2414,N_1187);
nor U5609 (N_5609,N_2416,N_415);
nand U5610 (N_5610,N_1859,N_893);
and U5611 (N_5611,N_2402,N_1653);
nand U5612 (N_5612,N_2720,N_462);
nor U5613 (N_5613,N_556,N_3568);
nand U5614 (N_5614,N_1845,N_3566);
nor U5615 (N_5615,N_3079,N_1100);
nand U5616 (N_5616,N_3816,N_3432);
nor U5617 (N_5617,N_3124,N_41);
or U5618 (N_5618,N_1162,N_3718);
xnor U5619 (N_5619,N_166,N_1108);
and U5620 (N_5620,N_3381,N_393);
nor U5621 (N_5621,N_650,N_61);
nor U5622 (N_5622,N_1878,N_215);
and U5623 (N_5623,N_1719,N_2316);
nor U5624 (N_5624,N_2743,N_2958);
xor U5625 (N_5625,N_3581,N_1840);
and U5626 (N_5626,N_3439,N_2231);
nand U5627 (N_5627,N_2875,N_3201);
nand U5628 (N_5628,N_103,N_1219);
nand U5629 (N_5629,N_888,N_1503);
and U5630 (N_5630,N_1581,N_1524);
nor U5631 (N_5631,N_1379,N_3023);
nand U5632 (N_5632,N_2132,N_3333);
or U5633 (N_5633,N_2698,N_427);
and U5634 (N_5634,N_1577,N_2972);
or U5635 (N_5635,N_1900,N_3216);
nor U5636 (N_5636,N_2483,N_3678);
or U5637 (N_5637,N_575,N_3649);
nor U5638 (N_5638,N_390,N_2471);
nand U5639 (N_5639,N_3682,N_1089);
or U5640 (N_5640,N_3450,N_3801);
or U5641 (N_5641,N_3317,N_2310);
and U5642 (N_5642,N_3416,N_2742);
nand U5643 (N_5643,N_232,N_3451);
and U5644 (N_5644,N_3227,N_1063);
or U5645 (N_5645,N_3091,N_2929);
and U5646 (N_5646,N_2023,N_2729);
nand U5647 (N_5647,N_3954,N_3435);
and U5648 (N_5648,N_3889,N_293);
and U5649 (N_5649,N_101,N_3226);
nor U5650 (N_5650,N_2445,N_1467);
and U5651 (N_5651,N_2351,N_3009);
and U5652 (N_5652,N_2260,N_3366);
nor U5653 (N_5653,N_1828,N_516);
or U5654 (N_5654,N_153,N_2080);
nor U5655 (N_5655,N_615,N_3867);
xnor U5656 (N_5656,N_3480,N_1413);
or U5657 (N_5657,N_557,N_3699);
and U5658 (N_5658,N_151,N_1271);
and U5659 (N_5659,N_1537,N_3353);
or U5660 (N_5660,N_1950,N_1368);
nor U5661 (N_5661,N_3453,N_2859);
nand U5662 (N_5662,N_133,N_544);
nand U5663 (N_5663,N_31,N_2116);
and U5664 (N_5664,N_2484,N_3601);
nand U5665 (N_5665,N_3694,N_1591);
nor U5666 (N_5666,N_1149,N_1029);
or U5667 (N_5667,N_1837,N_1969);
nor U5668 (N_5668,N_685,N_2988);
or U5669 (N_5669,N_2648,N_3532);
or U5670 (N_5670,N_3176,N_1075);
or U5671 (N_5671,N_3284,N_3306);
nand U5672 (N_5672,N_2549,N_571);
nor U5673 (N_5673,N_783,N_294);
xnor U5674 (N_5674,N_4,N_847);
xnor U5675 (N_5675,N_1601,N_1190);
or U5676 (N_5676,N_3732,N_3360);
nand U5677 (N_5677,N_1416,N_747);
and U5678 (N_5678,N_274,N_3421);
and U5679 (N_5679,N_810,N_2339);
or U5680 (N_5680,N_3589,N_905);
nand U5681 (N_5681,N_2003,N_268);
xnor U5682 (N_5682,N_3142,N_2900);
nand U5683 (N_5683,N_1352,N_3932);
and U5684 (N_5684,N_870,N_429);
nor U5685 (N_5685,N_2312,N_3440);
nand U5686 (N_5686,N_3070,N_1067);
xnor U5687 (N_5687,N_1009,N_2608);
or U5688 (N_5688,N_927,N_2467);
or U5689 (N_5689,N_1678,N_816);
nand U5690 (N_5690,N_3749,N_1737);
nand U5691 (N_5691,N_3899,N_1057);
nor U5692 (N_5692,N_723,N_3612);
nor U5693 (N_5693,N_3056,N_1264);
xor U5694 (N_5694,N_1852,N_1568);
nor U5695 (N_5695,N_1755,N_1872);
nor U5696 (N_5696,N_77,N_3773);
and U5697 (N_5697,N_2074,N_2070);
or U5698 (N_5698,N_83,N_3646);
and U5699 (N_5699,N_984,N_3482);
xnor U5700 (N_5700,N_2098,N_2899);
nor U5701 (N_5701,N_320,N_443);
nand U5702 (N_5702,N_3524,N_2006);
and U5703 (N_5703,N_1960,N_2543);
and U5704 (N_5704,N_2300,N_3372);
and U5705 (N_5705,N_1088,N_2291);
nor U5706 (N_5706,N_671,N_3143);
or U5707 (N_5707,N_185,N_971);
nand U5708 (N_5708,N_886,N_481);
and U5709 (N_5709,N_1478,N_3860);
nand U5710 (N_5710,N_3116,N_2283);
and U5711 (N_5711,N_786,N_2780);
or U5712 (N_5712,N_125,N_1012);
nor U5713 (N_5713,N_3208,N_1980);
xor U5714 (N_5714,N_45,N_928);
nor U5715 (N_5715,N_1754,N_657);
or U5716 (N_5716,N_2229,N_2832);
nor U5717 (N_5717,N_442,N_1373);
and U5718 (N_5718,N_2492,N_2449);
nor U5719 (N_5719,N_1922,N_947);
and U5720 (N_5720,N_2709,N_3840);
or U5721 (N_5721,N_485,N_1178);
nor U5722 (N_5722,N_3961,N_2730);
or U5723 (N_5723,N_3898,N_1618);
nor U5724 (N_5724,N_761,N_3086);
nand U5725 (N_5725,N_1013,N_1545);
or U5726 (N_5726,N_2952,N_3462);
nor U5727 (N_5727,N_3592,N_2121);
nor U5728 (N_5728,N_1288,N_973);
xor U5729 (N_5729,N_3082,N_1319);
or U5730 (N_5730,N_1415,N_1566);
and U5731 (N_5731,N_3635,N_2385);
or U5732 (N_5732,N_2957,N_3559);
xor U5733 (N_5733,N_2000,N_1887);
xnor U5734 (N_5734,N_3373,N_3925);
and U5735 (N_5735,N_1395,N_2124);
and U5736 (N_5736,N_1175,N_195);
or U5737 (N_5737,N_3182,N_1482);
nand U5738 (N_5738,N_1394,N_1238);
or U5739 (N_5739,N_2760,N_365);
nor U5740 (N_5740,N_190,N_3856);
and U5741 (N_5741,N_3821,N_3195);
or U5742 (N_5742,N_2787,N_2562);
or U5743 (N_5743,N_1448,N_1987);
nand U5744 (N_5744,N_3511,N_853);
and U5745 (N_5745,N_1037,N_1675);
xnor U5746 (N_5746,N_2907,N_275);
nand U5747 (N_5747,N_2475,N_652);
and U5748 (N_5748,N_3787,N_3183);
nand U5749 (N_5749,N_2071,N_3641);
xnor U5750 (N_5750,N_311,N_3835);
nand U5751 (N_5751,N_2045,N_3752);
and U5752 (N_5752,N_3924,N_2211);
nand U5753 (N_5753,N_1589,N_2756);
nor U5754 (N_5754,N_2154,N_70);
and U5755 (N_5755,N_2653,N_856);
nand U5756 (N_5756,N_3912,N_1074);
nand U5757 (N_5757,N_3677,N_1200);
nor U5758 (N_5758,N_1708,N_1022);
xor U5759 (N_5759,N_3456,N_341);
and U5760 (N_5760,N_743,N_1250);
or U5761 (N_5761,N_2628,N_2587);
or U5762 (N_5762,N_2688,N_2852);
or U5763 (N_5763,N_1542,N_2655);
nor U5764 (N_5764,N_3270,N_456);
or U5765 (N_5765,N_3951,N_2217);
xor U5766 (N_5766,N_3351,N_589);
and U5767 (N_5767,N_2120,N_253);
nand U5768 (N_5768,N_3044,N_2144);
nand U5769 (N_5769,N_2190,N_721);
nand U5770 (N_5770,N_1259,N_1489);
nand U5771 (N_5771,N_2195,N_337);
nand U5772 (N_5772,N_3492,N_838);
and U5773 (N_5773,N_2954,N_2055);
nor U5774 (N_5774,N_2647,N_3854);
xnor U5775 (N_5775,N_498,N_1632);
nand U5776 (N_5776,N_2029,N_1163);
and U5777 (N_5777,N_2065,N_3098);
nor U5778 (N_5778,N_658,N_3059);
nor U5779 (N_5779,N_1718,N_2657);
and U5780 (N_5780,N_567,N_3820);
and U5781 (N_5781,N_2804,N_648);
and U5782 (N_5782,N_371,N_1508);
and U5783 (N_5783,N_798,N_3406);
or U5784 (N_5784,N_2886,N_641);
nand U5785 (N_5785,N_1487,N_1451);
or U5786 (N_5786,N_348,N_2927);
and U5787 (N_5787,N_119,N_1390);
nor U5788 (N_5788,N_3983,N_1978);
nor U5789 (N_5789,N_73,N_2989);
or U5790 (N_5790,N_730,N_1168);
xnor U5791 (N_5791,N_3841,N_2049);
nor U5792 (N_5792,N_895,N_122);
xnor U5793 (N_5793,N_1337,N_3008);
nand U5794 (N_5794,N_2687,N_755);
or U5795 (N_5795,N_758,N_1435);
or U5796 (N_5796,N_2185,N_3890);
nand U5797 (N_5797,N_402,N_2950);
nor U5798 (N_5798,N_519,N_2792);
and U5799 (N_5799,N_1970,N_1616);
or U5800 (N_5800,N_517,N_3914);
nand U5801 (N_5801,N_3031,N_18);
and U5802 (N_5802,N_2974,N_449);
nor U5803 (N_5803,N_1253,N_2225);
nor U5804 (N_5804,N_1697,N_1883);
xor U5805 (N_5805,N_3775,N_883);
nand U5806 (N_5806,N_2622,N_3999);
nand U5807 (N_5807,N_2523,N_2345);
xnor U5808 (N_5808,N_1619,N_3477);
and U5809 (N_5809,N_404,N_59);
and U5810 (N_5810,N_520,N_239);
and U5811 (N_5811,N_3714,N_2579);
and U5812 (N_5812,N_2275,N_3870);
and U5813 (N_5813,N_1640,N_531);
and U5814 (N_5814,N_2181,N_707);
nand U5815 (N_5815,N_2427,N_3508);
nand U5816 (N_5816,N_66,N_1538);
xnor U5817 (N_5817,N_2847,N_2431);
nand U5818 (N_5818,N_800,N_2162);
or U5819 (N_5819,N_3136,N_1790);
nand U5820 (N_5820,N_1274,N_1857);
or U5821 (N_5821,N_152,N_582);
nand U5822 (N_5822,N_2118,N_1664);
nand U5823 (N_5823,N_1291,N_3137);
or U5824 (N_5824,N_2670,N_3827);
or U5825 (N_5825,N_2678,N_1308);
nand U5826 (N_5826,N_3294,N_3504);
and U5827 (N_5827,N_2535,N_338);
and U5828 (N_5828,N_138,N_2504);
and U5829 (N_5829,N_731,N_200);
nand U5830 (N_5830,N_1999,N_2079);
nand U5831 (N_5831,N_3625,N_142);
nand U5832 (N_5832,N_3929,N_2062);
nor U5833 (N_5833,N_3160,N_1431);
nand U5834 (N_5834,N_839,N_1806);
xor U5835 (N_5835,N_3071,N_256);
xor U5836 (N_5836,N_3871,N_68);
nor U5837 (N_5837,N_740,N_953);
or U5838 (N_5838,N_819,N_1938);
nor U5839 (N_5839,N_523,N_3804);
xor U5840 (N_5840,N_1042,N_1766);
and U5841 (N_5841,N_1622,N_3661);
nand U5842 (N_5842,N_2014,N_1297);
xnor U5843 (N_5843,N_2626,N_3437);
or U5844 (N_5844,N_413,N_3315);
or U5845 (N_5845,N_398,N_688);
nand U5846 (N_5846,N_3054,N_3861);
nor U5847 (N_5847,N_2102,N_2996);
nand U5848 (N_5848,N_3913,N_2660);
and U5849 (N_5849,N_3756,N_3906);
nor U5850 (N_5850,N_1594,N_351);
or U5851 (N_5851,N_807,N_3357);
nand U5852 (N_5852,N_163,N_3982);
and U5853 (N_5853,N_2497,N_1473);
and U5854 (N_5854,N_242,N_2814);
nand U5855 (N_5855,N_1679,N_2081);
or U5856 (N_5856,N_3348,N_771);
nor U5857 (N_5857,N_106,N_2891);
or U5858 (N_5858,N_2384,N_444);
or U5859 (N_5859,N_2094,N_3121);
nand U5860 (N_5860,N_3794,N_2694);
nand U5861 (N_5861,N_3027,N_2366);
xnor U5862 (N_5862,N_3560,N_1361);
and U5863 (N_5863,N_1849,N_3234);
nand U5864 (N_5864,N_988,N_3429);
and U5865 (N_5865,N_3277,N_987);
nor U5866 (N_5866,N_830,N_3470);
nor U5867 (N_5867,N_436,N_1406);
and U5868 (N_5868,N_224,N_2567);
xor U5869 (N_5869,N_1563,N_27);
nand U5870 (N_5870,N_3126,N_3987);
nand U5871 (N_5871,N_2654,N_2739);
or U5872 (N_5872,N_3569,N_1118);
or U5873 (N_5873,N_287,N_2495);
and U5874 (N_5874,N_2036,N_656);
nor U5875 (N_5875,N_1796,N_1229);
nor U5876 (N_5876,N_3290,N_3546);
and U5877 (N_5877,N_2477,N_2906);
nor U5878 (N_5878,N_1765,N_3134);
nor U5879 (N_5879,N_1667,N_3584);
xnor U5880 (N_5880,N_3385,N_2319);
and U5881 (N_5881,N_801,N_3269);
or U5882 (N_5882,N_1573,N_629);
nand U5883 (N_5883,N_1742,N_3245);
and U5884 (N_5884,N_3164,N_2296);
or U5885 (N_5885,N_1261,N_3928);
or U5886 (N_5886,N_2699,N_3447);
nand U5887 (N_5887,N_1453,N_3680);
nor U5888 (N_5888,N_3709,N_491);
xor U5889 (N_5889,N_84,N_2411);
nand U5890 (N_5890,N_1932,N_1753);
nor U5891 (N_5891,N_2324,N_126);
nand U5892 (N_5892,N_3459,N_861);
or U5893 (N_5893,N_2901,N_3166);
or U5894 (N_5894,N_368,N_1166);
nor U5895 (N_5895,N_3263,N_1692);
or U5896 (N_5896,N_975,N_2178);
nor U5897 (N_5897,N_1336,N_1492);
nor U5898 (N_5898,N_2458,N_1049);
nand U5899 (N_5899,N_3200,N_1414);
xnor U5900 (N_5900,N_961,N_805);
and U5901 (N_5901,N_3061,N_1360);
xnor U5902 (N_5902,N_2871,N_1105);
and U5903 (N_5903,N_2233,N_3043);
or U5904 (N_5904,N_3811,N_2646);
and U5905 (N_5905,N_469,N_2047);
or U5906 (N_5906,N_237,N_3989);
or U5907 (N_5907,N_2807,N_2336);
and U5908 (N_5908,N_3097,N_815);
nand U5909 (N_5909,N_3611,N_3449);
or U5910 (N_5910,N_2001,N_3039);
and U5911 (N_5911,N_1655,N_3621);
xor U5912 (N_5912,N_187,N_2479);
and U5913 (N_5913,N_808,N_1939);
or U5914 (N_5914,N_1986,N_2963);
nand U5915 (N_5915,N_774,N_1038);
and U5916 (N_5916,N_3530,N_1683);
or U5917 (N_5917,N_2263,N_2301);
and U5918 (N_5918,N_1305,N_2824);
and U5919 (N_5919,N_1405,N_1135);
nor U5920 (N_5920,N_1479,N_3874);
nand U5921 (N_5921,N_3352,N_3114);
xnor U5922 (N_5922,N_1183,N_507);
nor U5923 (N_5923,N_3639,N_2820);
or U5924 (N_5924,N_3576,N_765);
nand U5925 (N_5925,N_403,N_56);
or U5926 (N_5926,N_1902,N_2948);
nand U5927 (N_5927,N_3115,N_2346);
nand U5928 (N_5928,N_2327,N_16);
nor U5929 (N_5929,N_499,N_388);
or U5930 (N_5930,N_1119,N_2017);
nor U5931 (N_5931,N_2216,N_993);
nand U5932 (N_5932,N_2133,N_360);
and U5933 (N_5933,N_1445,N_3758);
or U5934 (N_5934,N_3909,N_3393);
xnor U5935 (N_5935,N_2268,N_749);
or U5936 (N_5936,N_1293,N_3986);
and U5937 (N_5937,N_1217,N_1734);
xnor U5938 (N_5938,N_1327,N_2072);
nand U5939 (N_5939,N_2109,N_831);
nor U5940 (N_5940,N_484,N_3785);
or U5941 (N_5941,N_3022,N_3557);
or U5942 (N_5942,N_1493,N_1270);
or U5943 (N_5943,N_2725,N_3401);
and U5944 (N_5944,N_682,N_1429);
xor U5945 (N_5945,N_1827,N_2818);
nor U5946 (N_5946,N_1306,N_1441);
and U5947 (N_5947,N_2673,N_43);
nand U5948 (N_5948,N_1826,N_3697);
xnor U5949 (N_5949,N_868,N_1729);
and U5950 (N_5950,N_346,N_2521);
nand U5951 (N_5951,N_2629,N_2248);
and U5952 (N_5952,N_158,N_1626);
nor U5953 (N_5953,N_2644,N_254);
and U5954 (N_5954,N_1598,N_2378);
or U5955 (N_5955,N_789,N_2063);
or U5956 (N_5956,N_3343,N_2583);
xnor U5957 (N_5957,N_1672,N_2459);
xor U5958 (N_5958,N_2188,N_2084);
and U5959 (N_5959,N_3738,N_1072);
or U5960 (N_5960,N_2816,N_3012);
and U5961 (N_5961,N_2514,N_829);
nand U5962 (N_5962,N_2273,N_2234);
or U5963 (N_5963,N_2825,N_2200);
xor U5964 (N_5964,N_3619,N_542);
nor U5965 (N_5965,N_3361,N_3422);
nor U5966 (N_5966,N_859,N_2683);
nand U5967 (N_5967,N_3135,N_1712);
nand U5968 (N_5968,N_3291,N_3918);
nand U5969 (N_5969,N_2085,N_234);
nor U5970 (N_5970,N_278,N_11);
or U5971 (N_5971,N_2536,N_1180);
and U5972 (N_5972,N_3053,N_3268);
xnor U5973 (N_5973,N_2841,N_3814);
nor U5974 (N_5974,N_1793,N_712);
and U5975 (N_5975,N_963,N_2309);
nand U5976 (N_5976,N_114,N_2138);
nand U5977 (N_5977,N_836,N_1717);
and U5978 (N_5978,N_1995,N_205);
and U5979 (N_5979,N_1570,N_2884);
or U5980 (N_5980,N_2288,N_970);
nand U5981 (N_5981,N_3370,N_1177);
or U5982 (N_5982,N_3665,N_3851);
nand U5983 (N_5983,N_2873,N_1823);
xnor U5984 (N_5984,N_3888,N_2237);
or U5985 (N_5985,N_1343,N_2179);
nor U5986 (N_5986,N_3327,N_1283);
or U5987 (N_5987,N_2765,N_1974);
and U5988 (N_5988,N_515,N_860);
nor U5989 (N_5989,N_2844,N_695);
nor U5990 (N_5990,N_2364,N_3479);
nand U5991 (N_5991,N_3049,N_822);
and U5992 (N_5992,N_1457,N_3132);
nor U5993 (N_5993,N_1756,N_447);
and U5994 (N_5994,N_2136,N_1052);
nand U5995 (N_5995,N_3809,N_598);
nor U5996 (N_5996,N_3302,N_3629);
nand U5997 (N_5997,N_1322,N_312);
and U5998 (N_5998,N_60,N_2348);
nand U5999 (N_5999,N_3312,N_2219);
nor U6000 (N_6000,N_2409,N_2850);
nor U6001 (N_6001,N_2000,N_2504);
xor U6002 (N_6002,N_207,N_2519);
and U6003 (N_6003,N_1600,N_3123);
nor U6004 (N_6004,N_777,N_1618);
xor U6005 (N_6005,N_1491,N_2232);
nor U6006 (N_6006,N_1612,N_1954);
or U6007 (N_6007,N_969,N_3326);
nor U6008 (N_6008,N_2544,N_3997);
or U6009 (N_6009,N_268,N_3410);
or U6010 (N_6010,N_1056,N_3214);
nor U6011 (N_6011,N_845,N_2687);
nor U6012 (N_6012,N_3213,N_2362);
xnor U6013 (N_6013,N_2686,N_3976);
xnor U6014 (N_6014,N_1719,N_1418);
and U6015 (N_6015,N_2141,N_2904);
nor U6016 (N_6016,N_829,N_2344);
or U6017 (N_6017,N_2200,N_1440);
or U6018 (N_6018,N_3862,N_1000);
nor U6019 (N_6019,N_1169,N_861);
nor U6020 (N_6020,N_1263,N_3567);
nor U6021 (N_6021,N_2709,N_3383);
or U6022 (N_6022,N_2219,N_2026);
xor U6023 (N_6023,N_224,N_826);
or U6024 (N_6024,N_24,N_2064);
nor U6025 (N_6025,N_366,N_1092);
or U6026 (N_6026,N_3728,N_391);
nand U6027 (N_6027,N_1355,N_2687);
nand U6028 (N_6028,N_1977,N_2839);
nand U6029 (N_6029,N_1407,N_1914);
and U6030 (N_6030,N_685,N_1510);
nor U6031 (N_6031,N_3987,N_366);
or U6032 (N_6032,N_2124,N_1919);
and U6033 (N_6033,N_1731,N_3123);
xnor U6034 (N_6034,N_563,N_2354);
nor U6035 (N_6035,N_2931,N_1234);
or U6036 (N_6036,N_3599,N_3387);
or U6037 (N_6037,N_3724,N_3317);
and U6038 (N_6038,N_306,N_3055);
and U6039 (N_6039,N_1899,N_1422);
nor U6040 (N_6040,N_1119,N_1234);
and U6041 (N_6041,N_552,N_1806);
nand U6042 (N_6042,N_1727,N_2706);
xnor U6043 (N_6043,N_2029,N_2035);
nor U6044 (N_6044,N_2122,N_3761);
nand U6045 (N_6045,N_2449,N_3025);
nor U6046 (N_6046,N_2412,N_2689);
nor U6047 (N_6047,N_2015,N_3290);
and U6048 (N_6048,N_3988,N_2302);
or U6049 (N_6049,N_884,N_217);
nand U6050 (N_6050,N_1368,N_1870);
nor U6051 (N_6051,N_3194,N_3227);
nand U6052 (N_6052,N_202,N_2051);
nand U6053 (N_6053,N_684,N_639);
nor U6054 (N_6054,N_3841,N_1954);
or U6055 (N_6055,N_3764,N_1450);
nand U6056 (N_6056,N_3087,N_2734);
nor U6057 (N_6057,N_477,N_615);
or U6058 (N_6058,N_277,N_885);
and U6059 (N_6059,N_3528,N_3805);
or U6060 (N_6060,N_707,N_2045);
and U6061 (N_6061,N_260,N_3895);
nand U6062 (N_6062,N_2536,N_190);
nor U6063 (N_6063,N_2001,N_2361);
and U6064 (N_6064,N_823,N_880);
nand U6065 (N_6065,N_1689,N_3066);
xnor U6066 (N_6066,N_1301,N_3769);
or U6067 (N_6067,N_2627,N_82);
nor U6068 (N_6068,N_1097,N_367);
and U6069 (N_6069,N_1514,N_2737);
xnor U6070 (N_6070,N_317,N_2545);
xor U6071 (N_6071,N_3956,N_950);
nand U6072 (N_6072,N_2867,N_831);
nor U6073 (N_6073,N_3953,N_807);
nor U6074 (N_6074,N_892,N_1706);
nand U6075 (N_6075,N_3882,N_3351);
and U6076 (N_6076,N_2591,N_3906);
nand U6077 (N_6077,N_3363,N_3155);
or U6078 (N_6078,N_2199,N_2919);
nand U6079 (N_6079,N_1425,N_2010);
and U6080 (N_6080,N_1378,N_2452);
or U6081 (N_6081,N_2803,N_2334);
nand U6082 (N_6082,N_3995,N_1314);
nor U6083 (N_6083,N_2094,N_2200);
or U6084 (N_6084,N_230,N_1081);
nand U6085 (N_6085,N_2986,N_419);
and U6086 (N_6086,N_2586,N_1195);
or U6087 (N_6087,N_143,N_1113);
nand U6088 (N_6088,N_2153,N_3208);
or U6089 (N_6089,N_1321,N_1119);
nor U6090 (N_6090,N_3785,N_2461);
or U6091 (N_6091,N_965,N_846);
or U6092 (N_6092,N_1291,N_2236);
nor U6093 (N_6093,N_420,N_2989);
or U6094 (N_6094,N_2775,N_3669);
nor U6095 (N_6095,N_1230,N_344);
nand U6096 (N_6096,N_2442,N_1482);
nand U6097 (N_6097,N_785,N_3515);
or U6098 (N_6098,N_2889,N_3767);
nand U6099 (N_6099,N_2291,N_3185);
and U6100 (N_6100,N_2938,N_3235);
nand U6101 (N_6101,N_23,N_3713);
and U6102 (N_6102,N_2264,N_3503);
xnor U6103 (N_6103,N_2633,N_1270);
and U6104 (N_6104,N_3927,N_2371);
and U6105 (N_6105,N_3958,N_918);
xor U6106 (N_6106,N_993,N_3629);
or U6107 (N_6107,N_3322,N_1707);
and U6108 (N_6108,N_920,N_2735);
nand U6109 (N_6109,N_687,N_2719);
or U6110 (N_6110,N_3411,N_1112);
or U6111 (N_6111,N_374,N_1719);
nor U6112 (N_6112,N_3282,N_779);
nand U6113 (N_6113,N_3397,N_203);
and U6114 (N_6114,N_1239,N_2663);
or U6115 (N_6115,N_3613,N_2287);
or U6116 (N_6116,N_1959,N_473);
nor U6117 (N_6117,N_2679,N_412);
nor U6118 (N_6118,N_760,N_3533);
and U6119 (N_6119,N_2497,N_3399);
xor U6120 (N_6120,N_2164,N_394);
nand U6121 (N_6121,N_3473,N_538);
and U6122 (N_6122,N_3490,N_3528);
nand U6123 (N_6123,N_2259,N_984);
and U6124 (N_6124,N_3478,N_2666);
nand U6125 (N_6125,N_956,N_3657);
nand U6126 (N_6126,N_2960,N_1460);
and U6127 (N_6127,N_3174,N_3945);
or U6128 (N_6128,N_2584,N_2385);
and U6129 (N_6129,N_387,N_1935);
or U6130 (N_6130,N_885,N_1343);
or U6131 (N_6131,N_932,N_886);
xnor U6132 (N_6132,N_1638,N_437);
nor U6133 (N_6133,N_823,N_1327);
and U6134 (N_6134,N_2848,N_3908);
and U6135 (N_6135,N_3243,N_907);
and U6136 (N_6136,N_3872,N_2315);
and U6137 (N_6137,N_3283,N_1187);
or U6138 (N_6138,N_543,N_3320);
nand U6139 (N_6139,N_3158,N_1463);
nand U6140 (N_6140,N_443,N_1512);
or U6141 (N_6141,N_238,N_858);
xnor U6142 (N_6142,N_2805,N_171);
xnor U6143 (N_6143,N_2938,N_2980);
and U6144 (N_6144,N_726,N_95);
or U6145 (N_6145,N_2088,N_3176);
nor U6146 (N_6146,N_2979,N_2317);
and U6147 (N_6147,N_1136,N_2259);
or U6148 (N_6148,N_3344,N_1233);
nor U6149 (N_6149,N_3365,N_1283);
xnor U6150 (N_6150,N_2694,N_1407);
nor U6151 (N_6151,N_2109,N_2099);
or U6152 (N_6152,N_478,N_1550);
nor U6153 (N_6153,N_182,N_899);
nand U6154 (N_6154,N_886,N_1200);
nand U6155 (N_6155,N_1158,N_2845);
xnor U6156 (N_6156,N_2952,N_1751);
nand U6157 (N_6157,N_2261,N_1530);
nor U6158 (N_6158,N_845,N_3796);
and U6159 (N_6159,N_3588,N_3172);
nand U6160 (N_6160,N_1011,N_1046);
or U6161 (N_6161,N_279,N_3288);
nand U6162 (N_6162,N_1291,N_2963);
nor U6163 (N_6163,N_982,N_1151);
or U6164 (N_6164,N_1505,N_3880);
and U6165 (N_6165,N_168,N_3060);
nor U6166 (N_6166,N_2109,N_2028);
xor U6167 (N_6167,N_3177,N_3653);
nor U6168 (N_6168,N_163,N_649);
and U6169 (N_6169,N_2268,N_1593);
and U6170 (N_6170,N_1901,N_2418);
nor U6171 (N_6171,N_54,N_681);
or U6172 (N_6172,N_2681,N_837);
or U6173 (N_6173,N_3443,N_834);
or U6174 (N_6174,N_3422,N_2312);
nor U6175 (N_6175,N_2684,N_886);
nand U6176 (N_6176,N_3472,N_581);
nor U6177 (N_6177,N_1973,N_3262);
nand U6178 (N_6178,N_2010,N_3085);
or U6179 (N_6179,N_2350,N_2433);
and U6180 (N_6180,N_3720,N_2483);
nor U6181 (N_6181,N_3358,N_1934);
nor U6182 (N_6182,N_2353,N_284);
nor U6183 (N_6183,N_253,N_3319);
or U6184 (N_6184,N_79,N_3470);
nor U6185 (N_6185,N_3063,N_3544);
nor U6186 (N_6186,N_2201,N_2345);
nand U6187 (N_6187,N_522,N_2304);
nor U6188 (N_6188,N_2636,N_1159);
xor U6189 (N_6189,N_1435,N_356);
nand U6190 (N_6190,N_2461,N_3011);
or U6191 (N_6191,N_1536,N_2454);
xnor U6192 (N_6192,N_1165,N_2682);
or U6193 (N_6193,N_890,N_2608);
nor U6194 (N_6194,N_2902,N_1397);
and U6195 (N_6195,N_2512,N_2460);
and U6196 (N_6196,N_2002,N_2654);
nor U6197 (N_6197,N_3438,N_1551);
nand U6198 (N_6198,N_190,N_2416);
nor U6199 (N_6199,N_2267,N_1670);
and U6200 (N_6200,N_376,N_3661);
or U6201 (N_6201,N_2678,N_3937);
or U6202 (N_6202,N_782,N_812);
nor U6203 (N_6203,N_3151,N_1674);
nand U6204 (N_6204,N_3573,N_869);
xnor U6205 (N_6205,N_2666,N_3715);
nor U6206 (N_6206,N_2432,N_1671);
xnor U6207 (N_6207,N_2735,N_1821);
and U6208 (N_6208,N_1330,N_2322);
and U6209 (N_6209,N_2156,N_905);
xor U6210 (N_6210,N_619,N_1378);
or U6211 (N_6211,N_777,N_3353);
nor U6212 (N_6212,N_72,N_3548);
nand U6213 (N_6213,N_1860,N_249);
nor U6214 (N_6214,N_862,N_700);
and U6215 (N_6215,N_2611,N_118);
nor U6216 (N_6216,N_3718,N_2850);
xor U6217 (N_6217,N_225,N_2680);
nor U6218 (N_6218,N_1440,N_1250);
nor U6219 (N_6219,N_3818,N_467);
nor U6220 (N_6220,N_414,N_2615);
nand U6221 (N_6221,N_2194,N_1561);
nand U6222 (N_6222,N_3556,N_2944);
nor U6223 (N_6223,N_3711,N_1654);
nor U6224 (N_6224,N_2768,N_3723);
nor U6225 (N_6225,N_3930,N_1784);
nand U6226 (N_6226,N_80,N_674);
nor U6227 (N_6227,N_160,N_731);
and U6228 (N_6228,N_1216,N_2603);
nand U6229 (N_6229,N_721,N_1303);
nor U6230 (N_6230,N_1063,N_1636);
xor U6231 (N_6231,N_2779,N_2821);
or U6232 (N_6232,N_535,N_3565);
or U6233 (N_6233,N_3797,N_2231);
nand U6234 (N_6234,N_1844,N_3607);
and U6235 (N_6235,N_3657,N_2327);
nand U6236 (N_6236,N_1721,N_2518);
nor U6237 (N_6237,N_76,N_1446);
nor U6238 (N_6238,N_2160,N_1053);
or U6239 (N_6239,N_607,N_525);
and U6240 (N_6240,N_2228,N_3608);
and U6241 (N_6241,N_3843,N_2115);
nand U6242 (N_6242,N_1105,N_250);
xor U6243 (N_6243,N_930,N_667);
nor U6244 (N_6244,N_3559,N_1302);
nor U6245 (N_6245,N_2500,N_1601);
nand U6246 (N_6246,N_3595,N_3212);
nor U6247 (N_6247,N_1085,N_686);
and U6248 (N_6248,N_1709,N_655);
nand U6249 (N_6249,N_2494,N_2119);
or U6250 (N_6250,N_3546,N_186);
xnor U6251 (N_6251,N_595,N_2844);
and U6252 (N_6252,N_3294,N_904);
nor U6253 (N_6253,N_2056,N_188);
or U6254 (N_6254,N_621,N_2806);
or U6255 (N_6255,N_2043,N_1532);
nor U6256 (N_6256,N_900,N_3260);
nor U6257 (N_6257,N_1082,N_3841);
nor U6258 (N_6258,N_3695,N_1989);
and U6259 (N_6259,N_2005,N_1628);
and U6260 (N_6260,N_3480,N_2494);
or U6261 (N_6261,N_1807,N_2715);
nand U6262 (N_6262,N_1222,N_3503);
or U6263 (N_6263,N_12,N_3230);
or U6264 (N_6264,N_1308,N_2222);
xor U6265 (N_6265,N_2472,N_1411);
and U6266 (N_6266,N_3407,N_566);
or U6267 (N_6267,N_3665,N_3880);
nand U6268 (N_6268,N_28,N_1419);
and U6269 (N_6269,N_1188,N_3331);
and U6270 (N_6270,N_3025,N_3674);
nor U6271 (N_6271,N_3992,N_1597);
nand U6272 (N_6272,N_871,N_2989);
or U6273 (N_6273,N_1538,N_3699);
xnor U6274 (N_6274,N_2868,N_2967);
or U6275 (N_6275,N_1244,N_1471);
and U6276 (N_6276,N_510,N_220);
nand U6277 (N_6277,N_3046,N_22);
or U6278 (N_6278,N_376,N_1118);
nor U6279 (N_6279,N_1286,N_2810);
or U6280 (N_6280,N_3689,N_907);
and U6281 (N_6281,N_720,N_2017);
or U6282 (N_6282,N_468,N_3809);
or U6283 (N_6283,N_2241,N_101);
nand U6284 (N_6284,N_1373,N_3181);
nand U6285 (N_6285,N_1759,N_1921);
nor U6286 (N_6286,N_1125,N_1920);
or U6287 (N_6287,N_765,N_81);
xnor U6288 (N_6288,N_3630,N_871);
and U6289 (N_6289,N_3389,N_1891);
nand U6290 (N_6290,N_2121,N_3154);
or U6291 (N_6291,N_1364,N_3630);
nand U6292 (N_6292,N_3461,N_1011);
or U6293 (N_6293,N_3167,N_553);
or U6294 (N_6294,N_3043,N_3080);
nand U6295 (N_6295,N_2074,N_3563);
nand U6296 (N_6296,N_696,N_2443);
nor U6297 (N_6297,N_1632,N_1872);
or U6298 (N_6298,N_1436,N_2758);
xnor U6299 (N_6299,N_3535,N_1211);
nor U6300 (N_6300,N_3236,N_3524);
and U6301 (N_6301,N_825,N_3367);
or U6302 (N_6302,N_2915,N_342);
and U6303 (N_6303,N_397,N_2866);
nand U6304 (N_6304,N_325,N_3596);
and U6305 (N_6305,N_1240,N_260);
and U6306 (N_6306,N_2562,N_898);
nand U6307 (N_6307,N_3641,N_2985);
xnor U6308 (N_6308,N_2685,N_1404);
nor U6309 (N_6309,N_2254,N_272);
nor U6310 (N_6310,N_1755,N_3031);
nand U6311 (N_6311,N_2300,N_467);
nand U6312 (N_6312,N_1300,N_1187);
nand U6313 (N_6313,N_406,N_3714);
nor U6314 (N_6314,N_1952,N_2777);
nor U6315 (N_6315,N_2736,N_1348);
or U6316 (N_6316,N_697,N_1542);
and U6317 (N_6317,N_603,N_670);
and U6318 (N_6318,N_1696,N_3767);
or U6319 (N_6319,N_2069,N_332);
xor U6320 (N_6320,N_1083,N_2159);
or U6321 (N_6321,N_2900,N_3739);
nor U6322 (N_6322,N_3739,N_2252);
nand U6323 (N_6323,N_87,N_3321);
nor U6324 (N_6324,N_528,N_1282);
nand U6325 (N_6325,N_228,N_3439);
nand U6326 (N_6326,N_3808,N_738);
nor U6327 (N_6327,N_1567,N_3638);
or U6328 (N_6328,N_508,N_2028);
nand U6329 (N_6329,N_3356,N_3277);
or U6330 (N_6330,N_1204,N_915);
or U6331 (N_6331,N_1034,N_3763);
or U6332 (N_6332,N_2352,N_1553);
or U6333 (N_6333,N_138,N_3091);
and U6334 (N_6334,N_917,N_2065);
nand U6335 (N_6335,N_672,N_3790);
and U6336 (N_6336,N_1758,N_3120);
or U6337 (N_6337,N_1924,N_2557);
nor U6338 (N_6338,N_1312,N_141);
or U6339 (N_6339,N_2186,N_3942);
or U6340 (N_6340,N_1460,N_3484);
xnor U6341 (N_6341,N_2584,N_1719);
nor U6342 (N_6342,N_3802,N_3689);
nand U6343 (N_6343,N_760,N_3617);
or U6344 (N_6344,N_586,N_2445);
nor U6345 (N_6345,N_3588,N_1120);
or U6346 (N_6346,N_1911,N_3694);
nand U6347 (N_6347,N_989,N_2255);
and U6348 (N_6348,N_918,N_191);
and U6349 (N_6349,N_36,N_530);
nand U6350 (N_6350,N_2560,N_217);
nand U6351 (N_6351,N_3069,N_680);
and U6352 (N_6352,N_3452,N_2900);
or U6353 (N_6353,N_3886,N_1072);
nand U6354 (N_6354,N_399,N_1514);
nor U6355 (N_6355,N_904,N_759);
nand U6356 (N_6356,N_1018,N_7);
or U6357 (N_6357,N_547,N_1451);
nand U6358 (N_6358,N_1539,N_1754);
nor U6359 (N_6359,N_359,N_3815);
xor U6360 (N_6360,N_3626,N_163);
nand U6361 (N_6361,N_3112,N_839);
or U6362 (N_6362,N_3352,N_2914);
nand U6363 (N_6363,N_547,N_1942);
xnor U6364 (N_6364,N_653,N_928);
or U6365 (N_6365,N_2779,N_3619);
or U6366 (N_6366,N_97,N_1162);
xor U6367 (N_6367,N_1753,N_301);
and U6368 (N_6368,N_2817,N_1237);
nand U6369 (N_6369,N_2135,N_3318);
and U6370 (N_6370,N_387,N_473);
nand U6371 (N_6371,N_338,N_2557);
and U6372 (N_6372,N_3144,N_239);
or U6373 (N_6373,N_1868,N_3503);
nor U6374 (N_6374,N_3792,N_1689);
xor U6375 (N_6375,N_2421,N_3158);
or U6376 (N_6376,N_278,N_1096);
and U6377 (N_6377,N_403,N_1328);
or U6378 (N_6378,N_2127,N_256);
or U6379 (N_6379,N_3909,N_3452);
or U6380 (N_6380,N_3862,N_3439);
or U6381 (N_6381,N_391,N_1046);
nand U6382 (N_6382,N_1664,N_3435);
and U6383 (N_6383,N_588,N_467);
and U6384 (N_6384,N_3619,N_3500);
nor U6385 (N_6385,N_3330,N_2324);
nand U6386 (N_6386,N_1808,N_226);
nand U6387 (N_6387,N_3791,N_3760);
or U6388 (N_6388,N_3838,N_530);
or U6389 (N_6389,N_3727,N_1011);
xor U6390 (N_6390,N_763,N_1687);
nor U6391 (N_6391,N_3792,N_1056);
or U6392 (N_6392,N_2057,N_3483);
nor U6393 (N_6393,N_89,N_3079);
or U6394 (N_6394,N_3476,N_2106);
or U6395 (N_6395,N_1084,N_1819);
nor U6396 (N_6396,N_1916,N_3824);
nand U6397 (N_6397,N_3738,N_1754);
nor U6398 (N_6398,N_788,N_1312);
nor U6399 (N_6399,N_2608,N_3644);
nand U6400 (N_6400,N_780,N_3421);
and U6401 (N_6401,N_2099,N_3932);
nor U6402 (N_6402,N_3573,N_2298);
nand U6403 (N_6403,N_3104,N_121);
nor U6404 (N_6404,N_3789,N_2647);
and U6405 (N_6405,N_1182,N_1266);
and U6406 (N_6406,N_2072,N_4);
nor U6407 (N_6407,N_957,N_1059);
and U6408 (N_6408,N_1759,N_792);
nor U6409 (N_6409,N_1681,N_3335);
xnor U6410 (N_6410,N_1224,N_467);
nand U6411 (N_6411,N_2124,N_2681);
or U6412 (N_6412,N_3455,N_3638);
and U6413 (N_6413,N_944,N_3805);
nand U6414 (N_6414,N_2203,N_2120);
nor U6415 (N_6415,N_1575,N_961);
nor U6416 (N_6416,N_2233,N_1270);
nor U6417 (N_6417,N_3800,N_1773);
or U6418 (N_6418,N_52,N_3763);
nand U6419 (N_6419,N_3823,N_2016);
and U6420 (N_6420,N_3869,N_3532);
or U6421 (N_6421,N_1407,N_3884);
nor U6422 (N_6422,N_1931,N_2187);
or U6423 (N_6423,N_3876,N_2572);
and U6424 (N_6424,N_1540,N_711);
or U6425 (N_6425,N_243,N_1194);
or U6426 (N_6426,N_233,N_2331);
and U6427 (N_6427,N_1282,N_1590);
and U6428 (N_6428,N_168,N_2551);
or U6429 (N_6429,N_3369,N_1263);
or U6430 (N_6430,N_3025,N_2385);
nor U6431 (N_6431,N_2620,N_1271);
or U6432 (N_6432,N_2861,N_3936);
or U6433 (N_6433,N_3021,N_2285);
xor U6434 (N_6434,N_2872,N_3675);
or U6435 (N_6435,N_1242,N_1636);
or U6436 (N_6436,N_540,N_1532);
and U6437 (N_6437,N_224,N_345);
and U6438 (N_6438,N_642,N_2015);
and U6439 (N_6439,N_2693,N_1607);
and U6440 (N_6440,N_832,N_1317);
or U6441 (N_6441,N_845,N_953);
and U6442 (N_6442,N_924,N_3024);
and U6443 (N_6443,N_2333,N_3563);
nand U6444 (N_6444,N_138,N_2984);
or U6445 (N_6445,N_1295,N_1465);
nor U6446 (N_6446,N_3313,N_1526);
nor U6447 (N_6447,N_2609,N_2042);
nor U6448 (N_6448,N_1772,N_3085);
or U6449 (N_6449,N_3021,N_3180);
or U6450 (N_6450,N_3633,N_2071);
or U6451 (N_6451,N_2344,N_1788);
nand U6452 (N_6452,N_2875,N_2172);
nor U6453 (N_6453,N_192,N_3090);
xnor U6454 (N_6454,N_2918,N_2405);
or U6455 (N_6455,N_683,N_3188);
or U6456 (N_6456,N_1684,N_3377);
or U6457 (N_6457,N_1554,N_1181);
nor U6458 (N_6458,N_1994,N_2807);
nand U6459 (N_6459,N_3616,N_1539);
or U6460 (N_6460,N_2257,N_293);
nor U6461 (N_6461,N_981,N_3549);
xor U6462 (N_6462,N_171,N_1191);
nand U6463 (N_6463,N_3520,N_2716);
and U6464 (N_6464,N_483,N_511);
and U6465 (N_6465,N_468,N_2604);
nor U6466 (N_6466,N_880,N_974);
and U6467 (N_6467,N_2207,N_300);
and U6468 (N_6468,N_3143,N_1129);
nand U6469 (N_6469,N_4,N_1712);
or U6470 (N_6470,N_2556,N_3118);
and U6471 (N_6471,N_1742,N_1958);
or U6472 (N_6472,N_2881,N_2926);
nor U6473 (N_6473,N_3809,N_1293);
and U6474 (N_6474,N_563,N_645);
or U6475 (N_6475,N_1975,N_513);
nor U6476 (N_6476,N_214,N_571);
nand U6477 (N_6477,N_1670,N_3428);
and U6478 (N_6478,N_1123,N_222);
xor U6479 (N_6479,N_2246,N_859);
or U6480 (N_6480,N_541,N_1938);
or U6481 (N_6481,N_3073,N_745);
and U6482 (N_6482,N_1970,N_3597);
nor U6483 (N_6483,N_2445,N_571);
or U6484 (N_6484,N_1185,N_2135);
nand U6485 (N_6485,N_1183,N_126);
and U6486 (N_6486,N_961,N_2100);
nor U6487 (N_6487,N_3135,N_3766);
nor U6488 (N_6488,N_2044,N_441);
or U6489 (N_6489,N_3614,N_3594);
and U6490 (N_6490,N_3595,N_2925);
or U6491 (N_6491,N_3123,N_1525);
nor U6492 (N_6492,N_1609,N_779);
xor U6493 (N_6493,N_764,N_1461);
nand U6494 (N_6494,N_2632,N_3016);
nand U6495 (N_6495,N_3613,N_2018);
or U6496 (N_6496,N_1368,N_2380);
or U6497 (N_6497,N_3014,N_884);
nand U6498 (N_6498,N_708,N_3007);
nor U6499 (N_6499,N_963,N_1301);
xnor U6500 (N_6500,N_1269,N_2535);
and U6501 (N_6501,N_2060,N_3669);
and U6502 (N_6502,N_625,N_1213);
xnor U6503 (N_6503,N_950,N_3049);
and U6504 (N_6504,N_1090,N_3315);
and U6505 (N_6505,N_3107,N_3409);
and U6506 (N_6506,N_832,N_1923);
nand U6507 (N_6507,N_1418,N_2212);
nor U6508 (N_6508,N_3716,N_2210);
nand U6509 (N_6509,N_2654,N_3056);
nor U6510 (N_6510,N_263,N_179);
xor U6511 (N_6511,N_2046,N_3732);
and U6512 (N_6512,N_2797,N_1887);
nor U6513 (N_6513,N_3590,N_3517);
or U6514 (N_6514,N_1055,N_835);
nand U6515 (N_6515,N_1130,N_3162);
and U6516 (N_6516,N_2671,N_3602);
nand U6517 (N_6517,N_1508,N_844);
nor U6518 (N_6518,N_1260,N_3171);
nor U6519 (N_6519,N_1392,N_2560);
nor U6520 (N_6520,N_2693,N_1069);
and U6521 (N_6521,N_2064,N_2467);
xor U6522 (N_6522,N_170,N_245);
xnor U6523 (N_6523,N_1724,N_3782);
xnor U6524 (N_6524,N_1676,N_3405);
nand U6525 (N_6525,N_817,N_3813);
xor U6526 (N_6526,N_1672,N_3776);
nand U6527 (N_6527,N_2105,N_3458);
and U6528 (N_6528,N_1751,N_3937);
or U6529 (N_6529,N_1430,N_586);
nor U6530 (N_6530,N_1755,N_1378);
and U6531 (N_6531,N_2201,N_1959);
or U6532 (N_6532,N_2591,N_2430);
nor U6533 (N_6533,N_213,N_3834);
nor U6534 (N_6534,N_2594,N_128);
nor U6535 (N_6535,N_2026,N_259);
and U6536 (N_6536,N_2791,N_617);
or U6537 (N_6537,N_1961,N_1394);
and U6538 (N_6538,N_1167,N_3144);
nor U6539 (N_6539,N_3693,N_3305);
and U6540 (N_6540,N_2462,N_2501);
nor U6541 (N_6541,N_2830,N_1904);
nor U6542 (N_6542,N_2084,N_3673);
or U6543 (N_6543,N_2855,N_144);
xor U6544 (N_6544,N_663,N_2787);
nor U6545 (N_6545,N_3539,N_2769);
nor U6546 (N_6546,N_911,N_1380);
and U6547 (N_6547,N_42,N_665);
or U6548 (N_6548,N_2032,N_1772);
nand U6549 (N_6549,N_3056,N_2971);
and U6550 (N_6550,N_3817,N_2972);
nand U6551 (N_6551,N_3754,N_3189);
and U6552 (N_6552,N_2283,N_62);
nand U6553 (N_6553,N_1472,N_2049);
and U6554 (N_6554,N_2709,N_1361);
nor U6555 (N_6555,N_1054,N_2778);
and U6556 (N_6556,N_3206,N_2386);
and U6557 (N_6557,N_859,N_560);
nor U6558 (N_6558,N_3791,N_545);
xor U6559 (N_6559,N_792,N_913);
nor U6560 (N_6560,N_2122,N_3196);
and U6561 (N_6561,N_2002,N_1912);
nor U6562 (N_6562,N_3545,N_1886);
nor U6563 (N_6563,N_2481,N_3119);
or U6564 (N_6564,N_3210,N_3474);
nor U6565 (N_6565,N_2883,N_2390);
and U6566 (N_6566,N_5,N_1438);
nor U6567 (N_6567,N_1818,N_2143);
nor U6568 (N_6568,N_2592,N_3094);
xnor U6569 (N_6569,N_3073,N_953);
or U6570 (N_6570,N_1925,N_2924);
and U6571 (N_6571,N_1401,N_926);
xor U6572 (N_6572,N_2727,N_3648);
nand U6573 (N_6573,N_329,N_2901);
and U6574 (N_6574,N_3407,N_306);
nand U6575 (N_6575,N_721,N_417);
nor U6576 (N_6576,N_3143,N_2480);
or U6577 (N_6577,N_1141,N_1495);
or U6578 (N_6578,N_3288,N_60);
or U6579 (N_6579,N_95,N_1020);
nand U6580 (N_6580,N_3398,N_3404);
or U6581 (N_6581,N_1763,N_1249);
or U6582 (N_6582,N_1323,N_2053);
nor U6583 (N_6583,N_2781,N_2439);
or U6584 (N_6584,N_2145,N_3206);
and U6585 (N_6585,N_1076,N_3969);
nand U6586 (N_6586,N_2212,N_1472);
xor U6587 (N_6587,N_2940,N_1824);
xor U6588 (N_6588,N_2364,N_2175);
nor U6589 (N_6589,N_2480,N_1638);
nand U6590 (N_6590,N_462,N_1443);
and U6591 (N_6591,N_3769,N_794);
and U6592 (N_6592,N_608,N_156);
nor U6593 (N_6593,N_60,N_10);
and U6594 (N_6594,N_3487,N_2866);
and U6595 (N_6595,N_1598,N_1891);
and U6596 (N_6596,N_258,N_2714);
nor U6597 (N_6597,N_3040,N_2226);
nor U6598 (N_6598,N_2540,N_1131);
xor U6599 (N_6599,N_1578,N_3931);
nand U6600 (N_6600,N_2356,N_739);
nand U6601 (N_6601,N_1859,N_968);
and U6602 (N_6602,N_937,N_3375);
nor U6603 (N_6603,N_2560,N_665);
or U6604 (N_6604,N_2621,N_3280);
and U6605 (N_6605,N_2032,N_1200);
nand U6606 (N_6606,N_2214,N_1677);
nand U6607 (N_6607,N_797,N_669);
nor U6608 (N_6608,N_2378,N_3917);
and U6609 (N_6609,N_1343,N_827);
or U6610 (N_6610,N_2819,N_3197);
or U6611 (N_6611,N_2818,N_1997);
and U6612 (N_6612,N_3869,N_3893);
and U6613 (N_6613,N_1522,N_197);
nand U6614 (N_6614,N_2965,N_1444);
nor U6615 (N_6615,N_2643,N_77);
and U6616 (N_6616,N_3374,N_242);
nand U6617 (N_6617,N_3406,N_771);
and U6618 (N_6618,N_3425,N_2417);
nor U6619 (N_6619,N_746,N_2282);
or U6620 (N_6620,N_284,N_2087);
or U6621 (N_6621,N_506,N_3867);
nand U6622 (N_6622,N_2332,N_1680);
and U6623 (N_6623,N_1079,N_2536);
or U6624 (N_6624,N_1714,N_125);
nor U6625 (N_6625,N_1275,N_3322);
xor U6626 (N_6626,N_2184,N_3926);
and U6627 (N_6627,N_619,N_2318);
and U6628 (N_6628,N_3769,N_2622);
nor U6629 (N_6629,N_1808,N_3323);
and U6630 (N_6630,N_2197,N_1430);
nor U6631 (N_6631,N_3851,N_175);
nor U6632 (N_6632,N_2539,N_190);
nand U6633 (N_6633,N_1801,N_3883);
nand U6634 (N_6634,N_2083,N_1274);
nor U6635 (N_6635,N_3187,N_1654);
or U6636 (N_6636,N_1421,N_2099);
or U6637 (N_6637,N_1928,N_1423);
and U6638 (N_6638,N_2904,N_2784);
nand U6639 (N_6639,N_1877,N_3280);
nand U6640 (N_6640,N_1558,N_316);
nand U6641 (N_6641,N_2849,N_2487);
nor U6642 (N_6642,N_2116,N_3047);
or U6643 (N_6643,N_106,N_1556);
nand U6644 (N_6644,N_3700,N_2239);
nand U6645 (N_6645,N_1555,N_892);
or U6646 (N_6646,N_3807,N_3176);
nor U6647 (N_6647,N_677,N_3505);
and U6648 (N_6648,N_3167,N_741);
and U6649 (N_6649,N_2115,N_3952);
or U6650 (N_6650,N_3317,N_300);
nor U6651 (N_6651,N_3411,N_1387);
and U6652 (N_6652,N_653,N_843);
nor U6653 (N_6653,N_2268,N_2172);
or U6654 (N_6654,N_2650,N_3977);
nand U6655 (N_6655,N_1444,N_416);
nor U6656 (N_6656,N_3826,N_3250);
and U6657 (N_6657,N_3530,N_3109);
and U6658 (N_6658,N_601,N_3396);
and U6659 (N_6659,N_2783,N_709);
nor U6660 (N_6660,N_2361,N_528);
xor U6661 (N_6661,N_3689,N_3414);
and U6662 (N_6662,N_2678,N_2304);
xor U6663 (N_6663,N_134,N_459);
or U6664 (N_6664,N_175,N_1951);
or U6665 (N_6665,N_3540,N_1762);
and U6666 (N_6666,N_51,N_3569);
or U6667 (N_6667,N_416,N_2099);
nor U6668 (N_6668,N_3769,N_684);
or U6669 (N_6669,N_3053,N_837);
and U6670 (N_6670,N_2530,N_194);
xnor U6671 (N_6671,N_2380,N_1203);
nor U6672 (N_6672,N_1394,N_3302);
and U6673 (N_6673,N_1631,N_3598);
or U6674 (N_6674,N_912,N_33);
and U6675 (N_6675,N_553,N_1888);
or U6676 (N_6676,N_2300,N_3001);
and U6677 (N_6677,N_191,N_2652);
or U6678 (N_6678,N_448,N_2429);
nand U6679 (N_6679,N_1195,N_930);
and U6680 (N_6680,N_362,N_3464);
nand U6681 (N_6681,N_1844,N_2208);
and U6682 (N_6682,N_2575,N_408);
nor U6683 (N_6683,N_2795,N_1549);
or U6684 (N_6684,N_1162,N_2273);
nand U6685 (N_6685,N_1165,N_664);
nand U6686 (N_6686,N_483,N_2500);
or U6687 (N_6687,N_1323,N_2808);
or U6688 (N_6688,N_682,N_2752);
nor U6689 (N_6689,N_2053,N_650);
nand U6690 (N_6690,N_392,N_1116);
or U6691 (N_6691,N_908,N_1411);
and U6692 (N_6692,N_2534,N_3322);
nand U6693 (N_6693,N_1216,N_3275);
nor U6694 (N_6694,N_2713,N_425);
and U6695 (N_6695,N_1063,N_2697);
nand U6696 (N_6696,N_1421,N_1711);
nand U6697 (N_6697,N_1589,N_2021);
xor U6698 (N_6698,N_1389,N_3626);
xor U6699 (N_6699,N_2656,N_87);
nand U6700 (N_6700,N_571,N_1343);
nand U6701 (N_6701,N_702,N_961);
and U6702 (N_6702,N_1084,N_1519);
or U6703 (N_6703,N_2283,N_241);
and U6704 (N_6704,N_3521,N_68);
nand U6705 (N_6705,N_2260,N_835);
nand U6706 (N_6706,N_3142,N_1509);
or U6707 (N_6707,N_2416,N_1418);
nand U6708 (N_6708,N_2814,N_676);
nor U6709 (N_6709,N_3225,N_907);
and U6710 (N_6710,N_2224,N_82);
nand U6711 (N_6711,N_1912,N_1365);
nor U6712 (N_6712,N_3187,N_3471);
nor U6713 (N_6713,N_1494,N_3954);
nand U6714 (N_6714,N_966,N_3175);
or U6715 (N_6715,N_2354,N_694);
or U6716 (N_6716,N_3234,N_2308);
nand U6717 (N_6717,N_123,N_1714);
nand U6718 (N_6718,N_3218,N_1291);
or U6719 (N_6719,N_608,N_641);
nor U6720 (N_6720,N_3599,N_26);
xor U6721 (N_6721,N_671,N_1071);
xnor U6722 (N_6722,N_2110,N_2529);
xor U6723 (N_6723,N_2080,N_2040);
nor U6724 (N_6724,N_2508,N_912);
nor U6725 (N_6725,N_156,N_2435);
nor U6726 (N_6726,N_2539,N_1757);
nor U6727 (N_6727,N_1130,N_2204);
nand U6728 (N_6728,N_132,N_3690);
or U6729 (N_6729,N_277,N_2356);
or U6730 (N_6730,N_285,N_147);
or U6731 (N_6731,N_3666,N_3044);
nor U6732 (N_6732,N_2568,N_1059);
nor U6733 (N_6733,N_3632,N_2951);
xnor U6734 (N_6734,N_902,N_1054);
nor U6735 (N_6735,N_379,N_3030);
and U6736 (N_6736,N_1879,N_687);
or U6737 (N_6737,N_296,N_907);
nand U6738 (N_6738,N_1829,N_3931);
nand U6739 (N_6739,N_1285,N_3243);
nand U6740 (N_6740,N_1749,N_3760);
nand U6741 (N_6741,N_1564,N_2314);
and U6742 (N_6742,N_860,N_1447);
nor U6743 (N_6743,N_3965,N_3147);
nor U6744 (N_6744,N_165,N_980);
nand U6745 (N_6745,N_2043,N_1639);
xor U6746 (N_6746,N_2746,N_1271);
or U6747 (N_6747,N_840,N_2655);
nand U6748 (N_6748,N_1735,N_3374);
or U6749 (N_6749,N_807,N_3195);
and U6750 (N_6750,N_998,N_3177);
nand U6751 (N_6751,N_186,N_1192);
xor U6752 (N_6752,N_666,N_2596);
and U6753 (N_6753,N_2501,N_2739);
nand U6754 (N_6754,N_439,N_123);
nor U6755 (N_6755,N_469,N_1044);
or U6756 (N_6756,N_1433,N_567);
or U6757 (N_6757,N_2148,N_2714);
or U6758 (N_6758,N_594,N_1190);
nor U6759 (N_6759,N_736,N_978);
and U6760 (N_6760,N_3111,N_972);
xnor U6761 (N_6761,N_3313,N_3471);
nor U6762 (N_6762,N_3185,N_2276);
nand U6763 (N_6763,N_3970,N_519);
nand U6764 (N_6764,N_209,N_3695);
or U6765 (N_6765,N_1142,N_486);
nand U6766 (N_6766,N_2392,N_3413);
and U6767 (N_6767,N_900,N_1034);
or U6768 (N_6768,N_1068,N_3589);
nand U6769 (N_6769,N_1951,N_128);
and U6770 (N_6770,N_1241,N_2876);
or U6771 (N_6771,N_281,N_2530);
or U6772 (N_6772,N_2688,N_1075);
nand U6773 (N_6773,N_3621,N_1991);
and U6774 (N_6774,N_2013,N_1894);
xnor U6775 (N_6775,N_3934,N_2124);
and U6776 (N_6776,N_532,N_163);
xor U6777 (N_6777,N_403,N_2604);
and U6778 (N_6778,N_702,N_2814);
and U6779 (N_6779,N_1867,N_376);
nor U6780 (N_6780,N_1955,N_3429);
nor U6781 (N_6781,N_2403,N_337);
nand U6782 (N_6782,N_3635,N_3426);
or U6783 (N_6783,N_3613,N_2481);
or U6784 (N_6784,N_2022,N_73);
or U6785 (N_6785,N_224,N_3575);
nand U6786 (N_6786,N_894,N_1432);
or U6787 (N_6787,N_2849,N_2049);
and U6788 (N_6788,N_3070,N_1566);
or U6789 (N_6789,N_1601,N_2581);
nand U6790 (N_6790,N_651,N_358);
nand U6791 (N_6791,N_1070,N_3256);
and U6792 (N_6792,N_2904,N_3023);
or U6793 (N_6793,N_104,N_45);
xor U6794 (N_6794,N_1251,N_2096);
or U6795 (N_6795,N_2976,N_3584);
or U6796 (N_6796,N_3624,N_499);
and U6797 (N_6797,N_510,N_187);
nand U6798 (N_6798,N_2706,N_578);
and U6799 (N_6799,N_1332,N_389);
nor U6800 (N_6800,N_1800,N_3615);
nand U6801 (N_6801,N_3932,N_2537);
xor U6802 (N_6802,N_1304,N_210);
nor U6803 (N_6803,N_3261,N_3028);
nand U6804 (N_6804,N_1825,N_1528);
nand U6805 (N_6805,N_2456,N_2100);
or U6806 (N_6806,N_1663,N_2860);
xnor U6807 (N_6807,N_507,N_3432);
nand U6808 (N_6808,N_3602,N_311);
or U6809 (N_6809,N_3976,N_2959);
nand U6810 (N_6810,N_2773,N_2276);
or U6811 (N_6811,N_2339,N_422);
and U6812 (N_6812,N_3351,N_452);
xor U6813 (N_6813,N_1279,N_1452);
nor U6814 (N_6814,N_552,N_79);
nor U6815 (N_6815,N_3402,N_2060);
nor U6816 (N_6816,N_1518,N_135);
nor U6817 (N_6817,N_3620,N_3334);
nand U6818 (N_6818,N_2379,N_1108);
nor U6819 (N_6819,N_120,N_3065);
nand U6820 (N_6820,N_3516,N_138);
nor U6821 (N_6821,N_914,N_2470);
nor U6822 (N_6822,N_918,N_976);
nand U6823 (N_6823,N_898,N_3971);
nor U6824 (N_6824,N_3910,N_812);
nor U6825 (N_6825,N_1024,N_2267);
or U6826 (N_6826,N_961,N_1284);
nor U6827 (N_6827,N_224,N_2060);
or U6828 (N_6828,N_298,N_233);
xnor U6829 (N_6829,N_1870,N_1354);
or U6830 (N_6830,N_1757,N_2514);
nor U6831 (N_6831,N_1203,N_713);
nand U6832 (N_6832,N_2198,N_9);
nor U6833 (N_6833,N_1270,N_299);
nand U6834 (N_6834,N_1914,N_3114);
nor U6835 (N_6835,N_2384,N_3728);
or U6836 (N_6836,N_594,N_1381);
nand U6837 (N_6837,N_1801,N_614);
or U6838 (N_6838,N_2543,N_829);
xnor U6839 (N_6839,N_3635,N_1581);
or U6840 (N_6840,N_541,N_150);
nand U6841 (N_6841,N_908,N_879);
nand U6842 (N_6842,N_2578,N_1399);
or U6843 (N_6843,N_2841,N_1688);
or U6844 (N_6844,N_2305,N_3265);
nand U6845 (N_6845,N_2117,N_570);
nand U6846 (N_6846,N_1181,N_1573);
or U6847 (N_6847,N_1886,N_3678);
nand U6848 (N_6848,N_2185,N_3652);
nand U6849 (N_6849,N_1773,N_469);
or U6850 (N_6850,N_881,N_3856);
nor U6851 (N_6851,N_799,N_396);
nor U6852 (N_6852,N_2155,N_1065);
nand U6853 (N_6853,N_2556,N_3270);
and U6854 (N_6854,N_3827,N_1829);
and U6855 (N_6855,N_2596,N_574);
or U6856 (N_6856,N_1420,N_2060);
nand U6857 (N_6857,N_1068,N_1849);
nor U6858 (N_6858,N_195,N_1136);
and U6859 (N_6859,N_3460,N_2194);
and U6860 (N_6860,N_3138,N_3227);
and U6861 (N_6861,N_2052,N_2658);
and U6862 (N_6862,N_1387,N_967);
nor U6863 (N_6863,N_1910,N_2568);
nor U6864 (N_6864,N_3829,N_2434);
nor U6865 (N_6865,N_3882,N_3726);
nor U6866 (N_6866,N_367,N_3762);
and U6867 (N_6867,N_3862,N_2875);
or U6868 (N_6868,N_717,N_826);
nand U6869 (N_6869,N_2754,N_2849);
nor U6870 (N_6870,N_2377,N_1303);
xor U6871 (N_6871,N_515,N_3247);
nand U6872 (N_6872,N_167,N_1846);
nor U6873 (N_6873,N_110,N_1146);
and U6874 (N_6874,N_3,N_2784);
nand U6875 (N_6875,N_232,N_1644);
nand U6876 (N_6876,N_2584,N_3491);
and U6877 (N_6877,N_92,N_2003);
and U6878 (N_6878,N_3425,N_3774);
or U6879 (N_6879,N_1660,N_1266);
nor U6880 (N_6880,N_2649,N_2120);
nand U6881 (N_6881,N_613,N_1738);
nand U6882 (N_6882,N_1372,N_3713);
nand U6883 (N_6883,N_1166,N_661);
or U6884 (N_6884,N_1589,N_3206);
nand U6885 (N_6885,N_3712,N_1133);
or U6886 (N_6886,N_2297,N_2056);
nand U6887 (N_6887,N_735,N_1353);
nor U6888 (N_6888,N_3020,N_3590);
and U6889 (N_6889,N_187,N_3576);
nand U6890 (N_6890,N_3063,N_1334);
xor U6891 (N_6891,N_2692,N_1326);
nand U6892 (N_6892,N_3981,N_532);
nor U6893 (N_6893,N_2909,N_3629);
or U6894 (N_6894,N_1813,N_2716);
nand U6895 (N_6895,N_3057,N_2379);
nor U6896 (N_6896,N_3122,N_3601);
xor U6897 (N_6897,N_3778,N_3138);
or U6898 (N_6898,N_2650,N_3903);
and U6899 (N_6899,N_1380,N_896);
and U6900 (N_6900,N_3130,N_2844);
or U6901 (N_6901,N_150,N_3344);
or U6902 (N_6902,N_1547,N_1407);
nor U6903 (N_6903,N_1805,N_1596);
nand U6904 (N_6904,N_897,N_2696);
nor U6905 (N_6905,N_1783,N_2156);
and U6906 (N_6906,N_1696,N_2727);
nor U6907 (N_6907,N_2179,N_1843);
and U6908 (N_6908,N_605,N_389);
and U6909 (N_6909,N_3419,N_3239);
and U6910 (N_6910,N_3464,N_2182);
nor U6911 (N_6911,N_2246,N_2184);
nand U6912 (N_6912,N_3395,N_1158);
or U6913 (N_6913,N_25,N_3120);
and U6914 (N_6914,N_3995,N_280);
and U6915 (N_6915,N_1108,N_3478);
xor U6916 (N_6916,N_639,N_799);
nor U6917 (N_6917,N_1913,N_1604);
nand U6918 (N_6918,N_2935,N_3924);
or U6919 (N_6919,N_2160,N_758);
or U6920 (N_6920,N_2811,N_1586);
nor U6921 (N_6921,N_200,N_1177);
nand U6922 (N_6922,N_2397,N_3321);
nand U6923 (N_6923,N_3505,N_2926);
or U6924 (N_6924,N_174,N_970);
or U6925 (N_6925,N_3250,N_54);
nand U6926 (N_6926,N_491,N_1106);
nor U6927 (N_6927,N_442,N_3038);
nor U6928 (N_6928,N_1273,N_1751);
or U6929 (N_6929,N_1131,N_3673);
nand U6930 (N_6930,N_716,N_2868);
nand U6931 (N_6931,N_781,N_3384);
nor U6932 (N_6932,N_2238,N_117);
and U6933 (N_6933,N_2231,N_257);
nor U6934 (N_6934,N_810,N_473);
or U6935 (N_6935,N_2922,N_1510);
xnor U6936 (N_6936,N_685,N_194);
nand U6937 (N_6937,N_1890,N_3507);
nor U6938 (N_6938,N_2656,N_783);
xor U6939 (N_6939,N_631,N_684);
nor U6940 (N_6940,N_404,N_172);
nor U6941 (N_6941,N_656,N_3738);
or U6942 (N_6942,N_805,N_2605);
or U6943 (N_6943,N_681,N_3836);
and U6944 (N_6944,N_1094,N_3933);
xnor U6945 (N_6945,N_3887,N_1715);
and U6946 (N_6946,N_2208,N_1801);
nor U6947 (N_6947,N_459,N_2398);
nor U6948 (N_6948,N_2051,N_1568);
and U6949 (N_6949,N_1251,N_2375);
nand U6950 (N_6950,N_2126,N_3);
nor U6951 (N_6951,N_1285,N_2147);
and U6952 (N_6952,N_517,N_1851);
nor U6953 (N_6953,N_465,N_1214);
nor U6954 (N_6954,N_3512,N_518);
nand U6955 (N_6955,N_80,N_3837);
or U6956 (N_6956,N_6,N_478);
nor U6957 (N_6957,N_1022,N_1204);
or U6958 (N_6958,N_2381,N_1090);
and U6959 (N_6959,N_1980,N_3016);
or U6960 (N_6960,N_2469,N_3748);
or U6961 (N_6961,N_1009,N_3651);
or U6962 (N_6962,N_2100,N_1018);
or U6963 (N_6963,N_2526,N_2043);
and U6964 (N_6964,N_1129,N_2619);
nand U6965 (N_6965,N_1766,N_330);
nand U6966 (N_6966,N_2695,N_2209);
nor U6967 (N_6967,N_764,N_3210);
nor U6968 (N_6968,N_2012,N_3800);
and U6969 (N_6969,N_2082,N_734);
nor U6970 (N_6970,N_307,N_2921);
nor U6971 (N_6971,N_2960,N_3279);
and U6972 (N_6972,N_2967,N_431);
nand U6973 (N_6973,N_3418,N_1825);
and U6974 (N_6974,N_1035,N_2383);
and U6975 (N_6975,N_959,N_1026);
or U6976 (N_6976,N_1667,N_2832);
nor U6977 (N_6977,N_3070,N_3990);
nor U6978 (N_6978,N_3859,N_2143);
or U6979 (N_6979,N_2330,N_1470);
nand U6980 (N_6980,N_2657,N_926);
and U6981 (N_6981,N_213,N_934);
nor U6982 (N_6982,N_1517,N_3809);
nand U6983 (N_6983,N_2014,N_57);
nor U6984 (N_6984,N_2421,N_3952);
xor U6985 (N_6985,N_711,N_1835);
nand U6986 (N_6986,N_3408,N_2070);
nor U6987 (N_6987,N_3573,N_25);
xnor U6988 (N_6988,N_1868,N_3325);
nand U6989 (N_6989,N_3804,N_1886);
nand U6990 (N_6990,N_1615,N_761);
nand U6991 (N_6991,N_3516,N_185);
and U6992 (N_6992,N_209,N_3025);
and U6993 (N_6993,N_2939,N_3223);
or U6994 (N_6994,N_871,N_3166);
nor U6995 (N_6995,N_3533,N_1993);
and U6996 (N_6996,N_2763,N_2511);
and U6997 (N_6997,N_3565,N_3197);
nor U6998 (N_6998,N_2794,N_1929);
xnor U6999 (N_6999,N_2634,N_3246);
or U7000 (N_7000,N_2720,N_3557);
nor U7001 (N_7001,N_927,N_797);
and U7002 (N_7002,N_348,N_3642);
nor U7003 (N_7003,N_2039,N_2713);
nand U7004 (N_7004,N_35,N_696);
and U7005 (N_7005,N_3679,N_460);
xnor U7006 (N_7006,N_1597,N_806);
nand U7007 (N_7007,N_2584,N_2803);
xnor U7008 (N_7008,N_2685,N_2795);
or U7009 (N_7009,N_773,N_1058);
nor U7010 (N_7010,N_3786,N_165);
nand U7011 (N_7011,N_1370,N_417);
xor U7012 (N_7012,N_2473,N_3032);
nor U7013 (N_7013,N_383,N_557);
nand U7014 (N_7014,N_885,N_3712);
nor U7015 (N_7015,N_2182,N_1687);
or U7016 (N_7016,N_3992,N_1041);
or U7017 (N_7017,N_815,N_1119);
nor U7018 (N_7018,N_3807,N_2923);
and U7019 (N_7019,N_3585,N_2394);
nor U7020 (N_7020,N_516,N_213);
xnor U7021 (N_7021,N_3826,N_3286);
nor U7022 (N_7022,N_383,N_2355);
nand U7023 (N_7023,N_1762,N_2173);
or U7024 (N_7024,N_1996,N_1998);
or U7025 (N_7025,N_1711,N_1353);
and U7026 (N_7026,N_2174,N_1214);
or U7027 (N_7027,N_2005,N_1486);
or U7028 (N_7028,N_3046,N_3878);
xnor U7029 (N_7029,N_1035,N_2993);
or U7030 (N_7030,N_512,N_2094);
xor U7031 (N_7031,N_2543,N_835);
or U7032 (N_7032,N_3357,N_147);
nor U7033 (N_7033,N_2719,N_3252);
and U7034 (N_7034,N_1638,N_208);
and U7035 (N_7035,N_3887,N_2049);
nand U7036 (N_7036,N_2820,N_1656);
and U7037 (N_7037,N_1865,N_2937);
nor U7038 (N_7038,N_1364,N_206);
and U7039 (N_7039,N_1249,N_3576);
nor U7040 (N_7040,N_1724,N_1000);
or U7041 (N_7041,N_57,N_1703);
or U7042 (N_7042,N_2430,N_2210);
xnor U7043 (N_7043,N_1736,N_1434);
nand U7044 (N_7044,N_1905,N_3443);
nand U7045 (N_7045,N_2574,N_1626);
nor U7046 (N_7046,N_3987,N_1097);
nand U7047 (N_7047,N_1660,N_724);
or U7048 (N_7048,N_1468,N_1560);
or U7049 (N_7049,N_1882,N_1409);
nor U7050 (N_7050,N_233,N_333);
nand U7051 (N_7051,N_3156,N_3911);
nor U7052 (N_7052,N_3984,N_3693);
and U7053 (N_7053,N_3167,N_3170);
or U7054 (N_7054,N_3475,N_3355);
nand U7055 (N_7055,N_3352,N_1108);
or U7056 (N_7056,N_978,N_1610);
nor U7057 (N_7057,N_1372,N_1124);
nand U7058 (N_7058,N_1481,N_85);
and U7059 (N_7059,N_3118,N_3974);
or U7060 (N_7060,N_3396,N_460);
nand U7061 (N_7061,N_3992,N_1781);
or U7062 (N_7062,N_1698,N_3537);
and U7063 (N_7063,N_746,N_199);
nor U7064 (N_7064,N_1976,N_907);
nor U7065 (N_7065,N_3903,N_3727);
xor U7066 (N_7066,N_875,N_3469);
nor U7067 (N_7067,N_2685,N_2643);
xor U7068 (N_7068,N_850,N_3714);
xor U7069 (N_7069,N_2432,N_1508);
nor U7070 (N_7070,N_2993,N_2803);
and U7071 (N_7071,N_3045,N_2631);
nand U7072 (N_7072,N_1454,N_905);
xor U7073 (N_7073,N_3301,N_2652);
and U7074 (N_7074,N_1325,N_3505);
nand U7075 (N_7075,N_3748,N_1828);
nand U7076 (N_7076,N_3405,N_1582);
nor U7077 (N_7077,N_1165,N_483);
nor U7078 (N_7078,N_1482,N_1801);
nand U7079 (N_7079,N_2243,N_2527);
nor U7080 (N_7080,N_980,N_3048);
and U7081 (N_7081,N_1510,N_616);
nor U7082 (N_7082,N_527,N_1529);
or U7083 (N_7083,N_3856,N_1156);
or U7084 (N_7084,N_446,N_1562);
nor U7085 (N_7085,N_907,N_3530);
or U7086 (N_7086,N_1442,N_1111);
or U7087 (N_7087,N_1261,N_3770);
or U7088 (N_7088,N_744,N_3766);
nand U7089 (N_7089,N_3631,N_1675);
and U7090 (N_7090,N_1001,N_69);
and U7091 (N_7091,N_2764,N_2782);
nand U7092 (N_7092,N_1304,N_407);
and U7093 (N_7093,N_3341,N_1629);
nor U7094 (N_7094,N_3558,N_2810);
nand U7095 (N_7095,N_627,N_1201);
or U7096 (N_7096,N_772,N_3171);
nand U7097 (N_7097,N_2816,N_3548);
and U7098 (N_7098,N_3899,N_2886);
or U7099 (N_7099,N_302,N_2401);
nor U7100 (N_7100,N_1555,N_1686);
or U7101 (N_7101,N_947,N_549);
or U7102 (N_7102,N_173,N_61);
xor U7103 (N_7103,N_220,N_2801);
nand U7104 (N_7104,N_1521,N_1380);
nand U7105 (N_7105,N_3316,N_1827);
nor U7106 (N_7106,N_3591,N_2510);
nor U7107 (N_7107,N_2334,N_3320);
nand U7108 (N_7108,N_2928,N_1220);
and U7109 (N_7109,N_2975,N_285);
and U7110 (N_7110,N_106,N_2485);
nor U7111 (N_7111,N_1647,N_773);
or U7112 (N_7112,N_2847,N_1715);
and U7113 (N_7113,N_626,N_1964);
or U7114 (N_7114,N_76,N_3917);
and U7115 (N_7115,N_2539,N_1138);
nor U7116 (N_7116,N_2439,N_3926);
and U7117 (N_7117,N_2364,N_990);
or U7118 (N_7118,N_3674,N_248);
nand U7119 (N_7119,N_2663,N_3840);
or U7120 (N_7120,N_621,N_1937);
or U7121 (N_7121,N_3580,N_2234);
nand U7122 (N_7122,N_2274,N_2609);
and U7123 (N_7123,N_1943,N_2658);
nor U7124 (N_7124,N_3863,N_3094);
nand U7125 (N_7125,N_1029,N_3353);
nand U7126 (N_7126,N_2343,N_1577);
nor U7127 (N_7127,N_1499,N_156);
and U7128 (N_7128,N_1756,N_667);
or U7129 (N_7129,N_2147,N_1510);
and U7130 (N_7130,N_3701,N_2833);
nand U7131 (N_7131,N_109,N_1013);
nor U7132 (N_7132,N_2513,N_2264);
and U7133 (N_7133,N_902,N_1097);
or U7134 (N_7134,N_264,N_599);
nand U7135 (N_7135,N_3039,N_3018);
xor U7136 (N_7136,N_3897,N_586);
nand U7137 (N_7137,N_722,N_3783);
or U7138 (N_7138,N_176,N_1180);
nor U7139 (N_7139,N_3043,N_2028);
and U7140 (N_7140,N_72,N_3945);
xor U7141 (N_7141,N_607,N_2018);
or U7142 (N_7142,N_2419,N_2607);
nor U7143 (N_7143,N_1877,N_2584);
nor U7144 (N_7144,N_2988,N_2287);
nor U7145 (N_7145,N_170,N_2745);
nor U7146 (N_7146,N_3698,N_2175);
nor U7147 (N_7147,N_745,N_179);
and U7148 (N_7148,N_3504,N_464);
or U7149 (N_7149,N_2801,N_357);
nor U7150 (N_7150,N_609,N_2903);
and U7151 (N_7151,N_963,N_867);
and U7152 (N_7152,N_2302,N_1488);
nor U7153 (N_7153,N_1274,N_3023);
and U7154 (N_7154,N_3049,N_1623);
and U7155 (N_7155,N_3468,N_2154);
nor U7156 (N_7156,N_1068,N_3816);
and U7157 (N_7157,N_111,N_2208);
nor U7158 (N_7158,N_3555,N_2606);
nand U7159 (N_7159,N_1660,N_458);
and U7160 (N_7160,N_1387,N_2039);
or U7161 (N_7161,N_2754,N_1424);
nor U7162 (N_7162,N_267,N_3045);
or U7163 (N_7163,N_3923,N_2472);
or U7164 (N_7164,N_2137,N_3758);
nand U7165 (N_7165,N_1744,N_3254);
nand U7166 (N_7166,N_22,N_325);
nand U7167 (N_7167,N_597,N_298);
or U7168 (N_7168,N_2999,N_716);
and U7169 (N_7169,N_1299,N_1269);
nor U7170 (N_7170,N_1235,N_3979);
nor U7171 (N_7171,N_644,N_332);
or U7172 (N_7172,N_2102,N_2521);
and U7173 (N_7173,N_981,N_2195);
nor U7174 (N_7174,N_120,N_1488);
and U7175 (N_7175,N_253,N_2423);
or U7176 (N_7176,N_3928,N_3039);
nand U7177 (N_7177,N_1126,N_3762);
nand U7178 (N_7178,N_2211,N_3865);
nand U7179 (N_7179,N_1710,N_1192);
and U7180 (N_7180,N_1944,N_324);
nand U7181 (N_7181,N_209,N_514);
nand U7182 (N_7182,N_619,N_30);
nand U7183 (N_7183,N_3116,N_3811);
nand U7184 (N_7184,N_1204,N_2132);
nor U7185 (N_7185,N_2089,N_3407);
and U7186 (N_7186,N_2000,N_1118);
xnor U7187 (N_7187,N_484,N_3637);
or U7188 (N_7188,N_3613,N_244);
xor U7189 (N_7189,N_1185,N_486);
nor U7190 (N_7190,N_965,N_2802);
nand U7191 (N_7191,N_1969,N_3296);
nor U7192 (N_7192,N_1236,N_2426);
nand U7193 (N_7193,N_920,N_1736);
nand U7194 (N_7194,N_3374,N_1644);
or U7195 (N_7195,N_2999,N_1852);
or U7196 (N_7196,N_3679,N_2473);
nor U7197 (N_7197,N_2715,N_747);
xnor U7198 (N_7198,N_23,N_2745);
or U7199 (N_7199,N_1013,N_8);
nand U7200 (N_7200,N_1672,N_1795);
nand U7201 (N_7201,N_2876,N_861);
nand U7202 (N_7202,N_394,N_3604);
or U7203 (N_7203,N_1028,N_3653);
and U7204 (N_7204,N_3450,N_869);
and U7205 (N_7205,N_2481,N_2569);
and U7206 (N_7206,N_2315,N_74);
nand U7207 (N_7207,N_2757,N_775);
or U7208 (N_7208,N_3795,N_3689);
and U7209 (N_7209,N_2465,N_894);
or U7210 (N_7210,N_2879,N_99);
and U7211 (N_7211,N_1332,N_159);
or U7212 (N_7212,N_1914,N_3680);
nor U7213 (N_7213,N_2108,N_3016);
and U7214 (N_7214,N_104,N_249);
nor U7215 (N_7215,N_1633,N_1653);
nand U7216 (N_7216,N_1035,N_2906);
and U7217 (N_7217,N_914,N_1757);
and U7218 (N_7218,N_858,N_2293);
or U7219 (N_7219,N_2621,N_2422);
and U7220 (N_7220,N_1165,N_1541);
nand U7221 (N_7221,N_3446,N_2057);
nand U7222 (N_7222,N_3250,N_1194);
or U7223 (N_7223,N_3868,N_527);
and U7224 (N_7224,N_3197,N_246);
or U7225 (N_7225,N_2194,N_3743);
or U7226 (N_7226,N_2794,N_2010);
and U7227 (N_7227,N_3789,N_3644);
nand U7228 (N_7228,N_3015,N_1085);
nor U7229 (N_7229,N_863,N_3225);
nand U7230 (N_7230,N_3119,N_565);
or U7231 (N_7231,N_3027,N_3182);
nor U7232 (N_7232,N_3626,N_2272);
nor U7233 (N_7233,N_2344,N_315);
or U7234 (N_7234,N_34,N_2095);
and U7235 (N_7235,N_108,N_3991);
nor U7236 (N_7236,N_3495,N_2517);
and U7237 (N_7237,N_574,N_2673);
xor U7238 (N_7238,N_1482,N_1955);
or U7239 (N_7239,N_2907,N_1516);
xnor U7240 (N_7240,N_2019,N_2517);
xnor U7241 (N_7241,N_2359,N_2533);
or U7242 (N_7242,N_2329,N_2313);
or U7243 (N_7243,N_3402,N_167);
and U7244 (N_7244,N_2779,N_1000);
or U7245 (N_7245,N_1357,N_1715);
nand U7246 (N_7246,N_3677,N_3009);
and U7247 (N_7247,N_1373,N_1362);
or U7248 (N_7248,N_1492,N_1484);
or U7249 (N_7249,N_974,N_1979);
nor U7250 (N_7250,N_1,N_3426);
nand U7251 (N_7251,N_1240,N_2164);
or U7252 (N_7252,N_1755,N_2498);
and U7253 (N_7253,N_2549,N_3742);
nand U7254 (N_7254,N_473,N_3455);
nor U7255 (N_7255,N_3512,N_3827);
or U7256 (N_7256,N_551,N_2669);
nor U7257 (N_7257,N_3032,N_1688);
nand U7258 (N_7258,N_2222,N_1219);
nand U7259 (N_7259,N_224,N_2726);
nand U7260 (N_7260,N_439,N_1862);
or U7261 (N_7261,N_3967,N_26);
nand U7262 (N_7262,N_2714,N_2691);
and U7263 (N_7263,N_3594,N_3481);
and U7264 (N_7264,N_3601,N_2042);
xor U7265 (N_7265,N_2903,N_1977);
or U7266 (N_7266,N_422,N_2019);
xnor U7267 (N_7267,N_1915,N_929);
or U7268 (N_7268,N_1549,N_1065);
nand U7269 (N_7269,N_3455,N_2876);
nor U7270 (N_7270,N_2735,N_1937);
nand U7271 (N_7271,N_1670,N_3976);
and U7272 (N_7272,N_3693,N_3569);
nor U7273 (N_7273,N_1800,N_809);
or U7274 (N_7274,N_2589,N_1666);
and U7275 (N_7275,N_2066,N_1649);
xnor U7276 (N_7276,N_3447,N_1097);
nand U7277 (N_7277,N_3280,N_1157);
or U7278 (N_7278,N_1027,N_261);
or U7279 (N_7279,N_470,N_963);
and U7280 (N_7280,N_677,N_2803);
xor U7281 (N_7281,N_1964,N_3244);
nand U7282 (N_7282,N_3167,N_3646);
xnor U7283 (N_7283,N_2670,N_2154);
and U7284 (N_7284,N_895,N_1321);
xor U7285 (N_7285,N_2864,N_1374);
or U7286 (N_7286,N_3222,N_3757);
or U7287 (N_7287,N_2259,N_3468);
nand U7288 (N_7288,N_3357,N_2655);
or U7289 (N_7289,N_2670,N_452);
nor U7290 (N_7290,N_2256,N_3411);
or U7291 (N_7291,N_2535,N_491);
nor U7292 (N_7292,N_1318,N_1749);
nand U7293 (N_7293,N_2040,N_3030);
nor U7294 (N_7294,N_1324,N_3319);
and U7295 (N_7295,N_1977,N_2896);
nor U7296 (N_7296,N_1919,N_1609);
and U7297 (N_7297,N_3356,N_1909);
nor U7298 (N_7298,N_1289,N_2457);
nor U7299 (N_7299,N_2476,N_2959);
and U7300 (N_7300,N_3738,N_1865);
xnor U7301 (N_7301,N_3168,N_3859);
or U7302 (N_7302,N_774,N_1225);
nor U7303 (N_7303,N_43,N_2607);
or U7304 (N_7304,N_1182,N_1630);
nand U7305 (N_7305,N_1152,N_3406);
and U7306 (N_7306,N_3835,N_3356);
or U7307 (N_7307,N_311,N_1709);
and U7308 (N_7308,N_870,N_2162);
and U7309 (N_7309,N_2902,N_1205);
xor U7310 (N_7310,N_1506,N_3245);
or U7311 (N_7311,N_2743,N_2133);
nor U7312 (N_7312,N_3469,N_390);
nor U7313 (N_7313,N_99,N_2753);
xor U7314 (N_7314,N_1521,N_3285);
nor U7315 (N_7315,N_2851,N_3890);
nor U7316 (N_7316,N_3904,N_549);
xor U7317 (N_7317,N_3892,N_2942);
nand U7318 (N_7318,N_2648,N_2343);
nor U7319 (N_7319,N_3150,N_3452);
and U7320 (N_7320,N_2443,N_1499);
nor U7321 (N_7321,N_3913,N_639);
nor U7322 (N_7322,N_3199,N_864);
nor U7323 (N_7323,N_548,N_2902);
or U7324 (N_7324,N_2570,N_3974);
or U7325 (N_7325,N_168,N_3708);
nand U7326 (N_7326,N_1295,N_374);
or U7327 (N_7327,N_848,N_1305);
or U7328 (N_7328,N_1295,N_2502);
and U7329 (N_7329,N_1222,N_524);
nor U7330 (N_7330,N_260,N_3491);
nand U7331 (N_7331,N_2654,N_179);
xnor U7332 (N_7332,N_789,N_3857);
and U7333 (N_7333,N_120,N_225);
and U7334 (N_7334,N_2392,N_624);
or U7335 (N_7335,N_2657,N_114);
and U7336 (N_7336,N_2141,N_2739);
or U7337 (N_7337,N_3512,N_860);
nor U7338 (N_7338,N_1018,N_2123);
and U7339 (N_7339,N_2234,N_1125);
nor U7340 (N_7340,N_2150,N_316);
nor U7341 (N_7341,N_3506,N_3850);
nand U7342 (N_7342,N_432,N_3989);
nand U7343 (N_7343,N_2683,N_3623);
and U7344 (N_7344,N_211,N_534);
nor U7345 (N_7345,N_1340,N_3957);
xor U7346 (N_7346,N_3023,N_3472);
xnor U7347 (N_7347,N_1769,N_2272);
nor U7348 (N_7348,N_1321,N_512);
nand U7349 (N_7349,N_1484,N_338);
nand U7350 (N_7350,N_306,N_2874);
or U7351 (N_7351,N_3211,N_2150);
or U7352 (N_7352,N_1826,N_3120);
and U7353 (N_7353,N_2642,N_330);
nor U7354 (N_7354,N_999,N_1743);
nor U7355 (N_7355,N_937,N_3908);
nand U7356 (N_7356,N_1359,N_2271);
xnor U7357 (N_7357,N_2843,N_681);
and U7358 (N_7358,N_2041,N_2533);
and U7359 (N_7359,N_1485,N_1030);
or U7360 (N_7360,N_3326,N_3683);
nand U7361 (N_7361,N_2335,N_575);
nor U7362 (N_7362,N_36,N_2851);
xnor U7363 (N_7363,N_344,N_749);
or U7364 (N_7364,N_3979,N_1077);
nand U7365 (N_7365,N_2561,N_2983);
nor U7366 (N_7366,N_2366,N_3795);
nor U7367 (N_7367,N_3496,N_1118);
nor U7368 (N_7368,N_2960,N_1874);
or U7369 (N_7369,N_586,N_689);
nand U7370 (N_7370,N_1111,N_1213);
nor U7371 (N_7371,N_3700,N_986);
and U7372 (N_7372,N_3245,N_1276);
and U7373 (N_7373,N_3015,N_2764);
nand U7374 (N_7374,N_478,N_706);
and U7375 (N_7375,N_3697,N_589);
nand U7376 (N_7376,N_3372,N_2984);
nand U7377 (N_7377,N_724,N_986);
xnor U7378 (N_7378,N_1758,N_2441);
nand U7379 (N_7379,N_801,N_1327);
nor U7380 (N_7380,N_3770,N_3607);
nand U7381 (N_7381,N_272,N_2625);
and U7382 (N_7382,N_2970,N_3794);
and U7383 (N_7383,N_953,N_3991);
and U7384 (N_7384,N_2621,N_1581);
nand U7385 (N_7385,N_2170,N_1844);
nand U7386 (N_7386,N_2113,N_1861);
nand U7387 (N_7387,N_3876,N_452);
and U7388 (N_7388,N_506,N_1634);
and U7389 (N_7389,N_71,N_2912);
nand U7390 (N_7390,N_530,N_1360);
nand U7391 (N_7391,N_2569,N_1057);
xor U7392 (N_7392,N_1829,N_2961);
xnor U7393 (N_7393,N_2655,N_1512);
nor U7394 (N_7394,N_3005,N_2646);
nor U7395 (N_7395,N_50,N_3364);
xor U7396 (N_7396,N_984,N_1105);
xnor U7397 (N_7397,N_3082,N_98);
nand U7398 (N_7398,N_3453,N_825);
and U7399 (N_7399,N_3184,N_2720);
or U7400 (N_7400,N_1836,N_1783);
nand U7401 (N_7401,N_2977,N_3318);
and U7402 (N_7402,N_526,N_3541);
nor U7403 (N_7403,N_1393,N_2844);
nor U7404 (N_7404,N_2555,N_1006);
or U7405 (N_7405,N_1370,N_2044);
nand U7406 (N_7406,N_2348,N_1991);
and U7407 (N_7407,N_3176,N_3629);
or U7408 (N_7408,N_1810,N_2620);
nor U7409 (N_7409,N_898,N_2929);
nor U7410 (N_7410,N_1290,N_159);
xor U7411 (N_7411,N_88,N_2045);
nor U7412 (N_7412,N_2853,N_769);
nor U7413 (N_7413,N_3490,N_3286);
nand U7414 (N_7414,N_601,N_2902);
and U7415 (N_7415,N_3543,N_2503);
nor U7416 (N_7416,N_2594,N_1793);
or U7417 (N_7417,N_710,N_1886);
or U7418 (N_7418,N_1986,N_1691);
nor U7419 (N_7419,N_3852,N_295);
nand U7420 (N_7420,N_3747,N_859);
nand U7421 (N_7421,N_1222,N_1412);
nand U7422 (N_7422,N_794,N_1871);
nand U7423 (N_7423,N_2925,N_1024);
xor U7424 (N_7424,N_2759,N_3424);
or U7425 (N_7425,N_2771,N_253);
or U7426 (N_7426,N_2211,N_283);
and U7427 (N_7427,N_2383,N_3710);
xnor U7428 (N_7428,N_1355,N_2351);
or U7429 (N_7429,N_2814,N_604);
nor U7430 (N_7430,N_1731,N_967);
or U7431 (N_7431,N_441,N_56);
and U7432 (N_7432,N_2063,N_1620);
and U7433 (N_7433,N_407,N_2395);
or U7434 (N_7434,N_523,N_2099);
nand U7435 (N_7435,N_1504,N_287);
nor U7436 (N_7436,N_1347,N_3772);
nand U7437 (N_7437,N_2597,N_2503);
nor U7438 (N_7438,N_2384,N_148);
nand U7439 (N_7439,N_3972,N_83);
and U7440 (N_7440,N_500,N_2581);
and U7441 (N_7441,N_2874,N_3015);
and U7442 (N_7442,N_266,N_1533);
nor U7443 (N_7443,N_3226,N_1589);
nor U7444 (N_7444,N_1919,N_3574);
and U7445 (N_7445,N_1070,N_3369);
or U7446 (N_7446,N_301,N_1605);
nor U7447 (N_7447,N_322,N_3057);
or U7448 (N_7448,N_2263,N_1357);
nor U7449 (N_7449,N_817,N_1142);
nor U7450 (N_7450,N_3677,N_1382);
xnor U7451 (N_7451,N_3320,N_3064);
or U7452 (N_7452,N_3897,N_3802);
nand U7453 (N_7453,N_2083,N_2230);
nand U7454 (N_7454,N_3680,N_1853);
nand U7455 (N_7455,N_23,N_1636);
and U7456 (N_7456,N_1570,N_863);
nor U7457 (N_7457,N_55,N_295);
and U7458 (N_7458,N_298,N_957);
or U7459 (N_7459,N_52,N_1463);
xor U7460 (N_7460,N_1826,N_2022);
nand U7461 (N_7461,N_3233,N_3357);
nand U7462 (N_7462,N_3973,N_1882);
nor U7463 (N_7463,N_1592,N_2715);
xnor U7464 (N_7464,N_2032,N_148);
or U7465 (N_7465,N_2543,N_119);
xor U7466 (N_7466,N_2151,N_1027);
nand U7467 (N_7467,N_1865,N_1847);
nand U7468 (N_7468,N_1009,N_3522);
or U7469 (N_7469,N_1506,N_1035);
xnor U7470 (N_7470,N_1514,N_3348);
and U7471 (N_7471,N_33,N_1428);
nor U7472 (N_7472,N_3619,N_468);
or U7473 (N_7473,N_1669,N_3623);
nand U7474 (N_7474,N_1911,N_2068);
or U7475 (N_7475,N_1286,N_1666);
xnor U7476 (N_7476,N_1310,N_2998);
nor U7477 (N_7477,N_1197,N_1626);
nand U7478 (N_7478,N_2442,N_18);
nor U7479 (N_7479,N_223,N_229);
nand U7480 (N_7480,N_3534,N_1282);
nor U7481 (N_7481,N_1545,N_809);
nand U7482 (N_7482,N_1801,N_2036);
nor U7483 (N_7483,N_2885,N_1609);
or U7484 (N_7484,N_3799,N_3033);
or U7485 (N_7485,N_2095,N_648);
nor U7486 (N_7486,N_3575,N_3583);
or U7487 (N_7487,N_3671,N_3274);
or U7488 (N_7488,N_3073,N_2245);
and U7489 (N_7489,N_1576,N_3326);
and U7490 (N_7490,N_1732,N_3956);
or U7491 (N_7491,N_2457,N_3329);
or U7492 (N_7492,N_1010,N_3210);
or U7493 (N_7493,N_3954,N_2340);
nand U7494 (N_7494,N_433,N_3835);
and U7495 (N_7495,N_383,N_1223);
and U7496 (N_7496,N_112,N_796);
nor U7497 (N_7497,N_2981,N_1834);
nor U7498 (N_7498,N_571,N_3071);
nor U7499 (N_7499,N_3620,N_2377);
nor U7500 (N_7500,N_1384,N_2023);
and U7501 (N_7501,N_3419,N_3854);
nor U7502 (N_7502,N_3759,N_1969);
and U7503 (N_7503,N_2178,N_3090);
xor U7504 (N_7504,N_1827,N_2484);
nand U7505 (N_7505,N_1271,N_3190);
xor U7506 (N_7506,N_3983,N_3125);
nor U7507 (N_7507,N_2264,N_464);
nor U7508 (N_7508,N_1478,N_271);
nor U7509 (N_7509,N_989,N_2640);
or U7510 (N_7510,N_3333,N_2741);
nor U7511 (N_7511,N_3079,N_3456);
nand U7512 (N_7512,N_3033,N_2740);
and U7513 (N_7513,N_2026,N_3311);
or U7514 (N_7514,N_1755,N_925);
xor U7515 (N_7515,N_1444,N_803);
nor U7516 (N_7516,N_2624,N_1906);
and U7517 (N_7517,N_847,N_2643);
nand U7518 (N_7518,N_3787,N_2458);
and U7519 (N_7519,N_1698,N_3919);
nand U7520 (N_7520,N_1438,N_1761);
nor U7521 (N_7521,N_1454,N_2860);
nand U7522 (N_7522,N_448,N_3327);
or U7523 (N_7523,N_3096,N_2893);
nor U7524 (N_7524,N_729,N_3405);
or U7525 (N_7525,N_2943,N_916);
and U7526 (N_7526,N_1192,N_1908);
or U7527 (N_7527,N_2828,N_1521);
and U7528 (N_7528,N_570,N_20);
xnor U7529 (N_7529,N_801,N_2242);
or U7530 (N_7530,N_1440,N_3517);
and U7531 (N_7531,N_2088,N_1186);
or U7532 (N_7532,N_1543,N_160);
nand U7533 (N_7533,N_2096,N_2840);
or U7534 (N_7534,N_2096,N_3932);
nor U7535 (N_7535,N_3943,N_2428);
nor U7536 (N_7536,N_3582,N_2131);
xor U7537 (N_7537,N_2731,N_2778);
and U7538 (N_7538,N_3238,N_344);
nand U7539 (N_7539,N_3177,N_280);
nor U7540 (N_7540,N_1435,N_2094);
nor U7541 (N_7541,N_1733,N_22);
nand U7542 (N_7542,N_1853,N_2063);
and U7543 (N_7543,N_898,N_2270);
and U7544 (N_7544,N_916,N_2844);
nor U7545 (N_7545,N_3595,N_533);
xor U7546 (N_7546,N_715,N_2446);
and U7547 (N_7547,N_3016,N_1555);
nand U7548 (N_7548,N_3022,N_2116);
xor U7549 (N_7549,N_4,N_2656);
or U7550 (N_7550,N_3297,N_2065);
or U7551 (N_7551,N_2525,N_1631);
and U7552 (N_7552,N_2407,N_1837);
and U7553 (N_7553,N_88,N_3289);
and U7554 (N_7554,N_1124,N_812);
nor U7555 (N_7555,N_1904,N_547);
and U7556 (N_7556,N_1297,N_3924);
nand U7557 (N_7557,N_2218,N_751);
and U7558 (N_7558,N_230,N_1515);
nor U7559 (N_7559,N_2623,N_3963);
and U7560 (N_7560,N_3573,N_246);
or U7561 (N_7561,N_3826,N_791);
nor U7562 (N_7562,N_329,N_3991);
and U7563 (N_7563,N_1476,N_3471);
xnor U7564 (N_7564,N_1235,N_554);
xnor U7565 (N_7565,N_3506,N_2941);
and U7566 (N_7566,N_3148,N_3041);
nand U7567 (N_7567,N_2623,N_192);
or U7568 (N_7568,N_2402,N_2304);
nor U7569 (N_7569,N_2933,N_3755);
xor U7570 (N_7570,N_2367,N_190);
or U7571 (N_7571,N_1290,N_3549);
nor U7572 (N_7572,N_1225,N_2597);
and U7573 (N_7573,N_959,N_3648);
or U7574 (N_7574,N_3499,N_3234);
nor U7575 (N_7575,N_889,N_3853);
nor U7576 (N_7576,N_1632,N_2867);
and U7577 (N_7577,N_2902,N_341);
and U7578 (N_7578,N_3644,N_1748);
and U7579 (N_7579,N_257,N_3036);
or U7580 (N_7580,N_140,N_2508);
nor U7581 (N_7581,N_949,N_1592);
and U7582 (N_7582,N_214,N_184);
nand U7583 (N_7583,N_922,N_3066);
and U7584 (N_7584,N_3517,N_408);
or U7585 (N_7585,N_3841,N_1923);
and U7586 (N_7586,N_2889,N_2893);
and U7587 (N_7587,N_1860,N_2347);
xor U7588 (N_7588,N_1586,N_269);
or U7589 (N_7589,N_83,N_2427);
and U7590 (N_7590,N_843,N_855);
nand U7591 (N_7591,N_2150,N_1208);
xnor U7592 (N_7592,N_2444,N_3943);
or U7593 (N_7593,N_3985,N_1345);
nand U7594 (N_7594,N_966,N_68);
nor U7595 (N_7595,N_2407,N_3402);
xor U7596 (N_7596,N_2138,N_1746);
nand U7597 (N_7597,N_500,N_3700);
or U7598 (N_7598,N_1905,N_158);
nor U7599 (N_7599,N_773,N_1691);
and U7600 (N_7600,N_1937,N_947);
or U7601 (N_7601,N_1117,N_3570);
or U7602 (N_7602,N_1134,N_662);
xor U7603 (N_7603,N_3079,N_1234);
nand U7604 (N_7604,N_998,N_1983);
nand U7605 (N_7605,N_1978,N_3300);
and U7606 (N_7606,N_1660,N_1600);
and U7607 (N_7607,N_2714,N_3765);
or U7608 (N_7608,N_1383,N_3673);
or U7609 (N_7609,N_3667,N_2782);
or U7610 (N_7610,N_810,N_3405);
or U7611 (N_7611,N_2083,N_3724);
nand U7612 (N_7612,N_3852,N_325);
xor U7613 (N_7613,N_2456,N_203);
and U7614 (N_7614,N_1619,N_2964);
or U7615 (N_7615,N_2059,N_567);
nor U7616 (N_7616,N_3462,N_2496);
nand U7617 (N_7617,N_2173,N_880);
nand U7618 (N_7618,N_3655,N_41);
or U7619 (N_7619,N_341,N_3772);
or U7620 (N_7620,N_1827,N_2519);
nor U7621 (N_7621,N_2305,N_2185);
nand U7622 (N_7622,N_469,N_2504);
or U7623 (N_7623,N_3153,N_2116);
or U7624 (N_7624,N_594,N_2660);
and U7625 (N_7625,N_482,N_3782);
or U7626 (N_7626,N_81,N_336);
and U7627 (N_7627,N_1284,N_2262);
nor U7628 (N_7628,N_183,N_3811);
xnor U7629 (N_7629,N_1336,N_342);
and U7630 (N_7630,N_3263,N_1925);
xor U7631 (N_7631,N_2395,N_1165);
and U7632 (N_7632,N_3897,N_3622);
xor U7633 (N_7633,N_2906,N_2616);
and U7634 (N_7634,N_1134,N_1764);
or U7635 (N_7635,N_1641,N_2411);
nand U7636 (N_7636,N_2595,N_1957);
nor U7637 (N_7637,N_3664,N_3409);
and U7638 (N_7638,N_1626,N_1324);
or U7639 (N_7639,N_1825,N_1463);
and U7640 (N_7640,N_3913,N_2334);
nor U7641 (N_7641,N_3489,N_1212);
nand U7642 (N_7642,N_278,N_3817);
and U7643 (N_7643,N_2037,N_1606);
and U7644 (N_7644,N_3646,N_2598);
and U7645 (N_7645,N_319,N_696);
and U7646 (N_7646,N_3520,N_3732);
and U7647 (N_7647,N_2807,N_495);
nor U7648 (N_7648,N_2950,N_3558);
nand U7649 (N_7649,N_2425,N_1992);
and U7650 (N_7650,N_3222,N_3035);
and U7651 (N_7651,N_1273,N_3265);
or U7652 (N_7652,N_568,N_928);
and U7653 (N_7653,N_1766,N_2653);
or U7654 (N_7654,N_248,N_2112);
and U7655 (N_7655,N_379,N_550);
nor U7656 (N_7656,N_1306,N_452);
nand U7657 (N_7657,N_3718,N_1666);
nand U7658 (N_7658,N_2860,N_812);
and U7659 (N_7659,N_1626,N_2883);
or U7660 (N_7660,N_622,N_402);
nand U7661 (N_7661,N_3416,N_3693);
and U7662 (N_7662,N_2448,N_2385);
nor U7663 (N_7663,N_2110,N_1156);
nand U7664 (N_7664,N_1107,N_1220);
and U7665 (N_7665,N_1640,N_1312);
or U7666 (N_7666,N_516,N_2955);
nand U7667 (N_7667,N_1604,N_2733);
or U7668 (N_7668,N_2333,N_3434);
or U7669 (N_7669,N_757,N_3485);
nor U7670 (N_7670,N_2299,N_1359);
and U7671 (N_7671,N_3201,N_3956);
xnor U7672 (N_7672,N_3142,N_3828);
nor U7673 (N_7673,N_1512,N_1544);
or U7674 (N_7674,N_2665,N_1731);
or U7675 (N_7675,N_2152,N_2294);
or U7676 (N_7676,N_2977,N_3690);
nand U7677 (N_7677,N_3197,N_1841);
or U7678 (N_7678,N_648,N_3277);
nor U7679 (N_7679,N_1818,N_1017);
nor U7680 (N_7680,N_2614,N_278);
or U7681 (N_7681,N_2003,N_1825);
nor U7682 (N_7682,N_2535,N_124);
or U7683 (N_7683,N_2605,N_3794);
and U7684 (N_7684,N_2546,N_127);
xor U7685 (N_7685,N_3514,N_1140);
or U7686 (N_7686,N_374,N_2036);
nor U7687 (N_7687,N_2044,N_14);
nor U7688 (N_7688,N_580,N_2723);
or U7689 (N_7689,N_2426,N_1733);
nor U7690 (N_7690,N_844,N_3609);
xor U7691 (N_7691,N_246,N_2348);
and U7692 (N_7692,N_2117,N_79);
or U7693 (N_7693,N_3024,N_370);
xnor U7694 (N_7694,N_1486,N_2952);
nor U7695 (N_7695,N_3424,N_1168);
or U7696 (N_7696,N_3524,N_3383);
nand U7697 (N_7697,N_554,N_1451);
or U7698 (N_7698,N_1134,N_3334);
and U7699 (N_7699,N_1318,N_1349);
and U7700 (N_7700,N_1085,N_3816);
nand U7701 (N_7701,N_3508,N_2152);
nand U7702 (N_7702,N_119,N_2977);
or U7703 (N_7703,N_1621,N_2320);
and U7704 (N_7704,N_2524,N_167);
or U7705 (N_7705,N_105,N_3980);
xor U7706 (N_7706,N_1759,N_2535);
nand U7707 (N_7707,N_2516,N_879);
nor U7708 (N_7708,N_2237,N_3295);
nor U7709 (N_7709,N_1292,N_3455);
nor U7710 (N_7710,N_3264,N_153);
nor U7711 (N_7711,N_901,N_2812);
nor U7712 (N_7712,N_3145,N_1053);
nand U7713 (N_7713,N_42,N_2447);
nor U7714 (N_7714,N_2938,N_2184);
or U7715 (N_7715,N_2446,N_354);
and U7716 (N_7716,N_483,N_526);
nand U7717 (N_7717,N_92,N_2868);
nor U7718 (N_7718,N_2008,N_1830);
and U7719 (N_7719,N_188,N_1563);
or U7720 (N_7720,N_2243,N_2158);
nand U7721 (N_7721,N_3777,N_212);
nor U7722 (N_7722,N_3882,N_2720);
or U7723 (N_7723,N_1967,N_102);
or U7724 (N_7724,N_2284,N_2773);
nand U7725 (N_7725,N_2984,N_703);
and U7726 (N_7726,N_1415,N_3188);
and U7727 (N_7727,N_731,N_505);
xnor U7728 (N_7728,N_3077,N_2851);
or U7729 (N_7729,N_3038,N_1858);
nor U7730 (N_7730,N_3226,N_1833);
nand U7731 (N_7731,N_2043,N_308);
and U7732 (N_7732,N_3595,N_2307);
or U7733 (N_7733,N_3325,N_1403);
nor U7734 (N_7734,N_673,N_2435);
nand U7735 (N_7735,N_2202,N_2815);
nand U7736 (N_7736,N_2845,N_675);
and U7737 (N_7737,N_1624,N_1254);
or U7738 (N_7738,N_1120,N_253);
nor U7739 (N_7739,N_223,N_2276);
nand U7740 (N_7740,N_1497,N_490);
and U7741 (N_7741,N_728,N_3839);
xnor U7742 (N_7742,N_952,N_954);
nor U7743 (N_7743,N_1022,N_2679);
and U7744 (N_7744,N_262,N_3020);
xnor U7745 (N_7745,N_871,N_2831);
nor U7746 (N_7746,N_1374,N_286);
nor U7747 (N_7747,N_3965,N_1293);
nand U7748 (N_7748,N_508,N_2483);
nand U7749 (N_7749,N_2370,N_2371);
nor U7750 (N_7750,N_2101,N_3454);
or U7751 (N_7751,N_986,N_629);
nor U7752 (N_7752,N_1036,N_983);
or U7753 (N_7753,N_3083,N_3758);
or U7754 (N_7754,N_3959,N_2146);
and U7755 (N_7755,N_974,N_551);
nand U7756 (N_7756,N_2586,N_867);
and U7757 (N_7757,N_3521,N_1679);
and U7758 (N_7758,N_501,N_717);
nor U7759 (N_7759,N_3282,N_2409);
and U7760 (N_7760,N_528,N_3772);
nand U7761 (N_7761,N_661,N_424);
xnor U7762 (N_7762,N_7,N_22);
nand U7763 (N_7763,N_3848,N_3953);
or U7764 (N_7764,N_20,N_2198);
nor U7765 (N_7765,N_1011,N_1017);
nand U7766 (N_7766,N_615,N_499);
or U7767 (N_7767,N_2068,N_3702);
or U7768 (N_7768,N_2264,N_1163);
nand U7769 (N_7769,N_685,N_3353);
nand U7770 (N_7770,N_1674,N_2547);
or U7771 (N_7771,N_2191,N_3325);
and U7772 (N_7772,N_2722,N_510);
nor U7773 (N_7773,N_1602,N_3649);
nand U7774 (N_7774,N_3093,N_2993);
nor U7775 (N_7775,N_840,N_386);
nand U7776 (N_7776,N_2509,N_173);
and U7777 (N_7777,N_1075,N_1247);
xnor U7778 (N_7778,N_2481,N_3023);
or U7779 (N_7779,N_2176,N_3219);
and U7780 (N_7780,N_2123,N_189);
and U7781 (N_7781,N_1016,N_3223);
nor U7782 (N_7782,N_31,N_3868);
nand U7783 (N_7783,N_2531,N_1953);
or U7784 (N_7784,N_2145,N_3430);
or U7785 (N_7785,N_255,N_517);
or U7786 (N_7786,N_1052,N_3618);
nor U7787 (N_7787,N_456,N_213);
or U7788 (N_7788,N_1302,N_2719);
and U7789 (N_7789,N_736,N_2693);
nand U7790 (N_7790,N_1214,N_682);
nand U7791 (N_7791,N_2739,N_1182);
xnor U7792 (N_7792,N_531,N_343);
nor U7793 (N_7793,N_833,N_3700);
or U7794 (N_7794,N_3992,N_1529);
or U7795 (N_7795,N_2715,N_3941);
and U7796 (N_7796,N_2390,N_2725);
and U7797 (N_7797,N_2675,N_506);
and U7798 (N_7798,N_2669,N_3135);
nor U7799 (N_7799,N_3025,N_349);
and U7800 (N_7800,N_3594,N_493);
or U7801 (N_7801,N_3328,N_3699);
xor U7802 (N_7802,N_1190,N_3038);
nand U7803 (N_7803,N_3780,N_1363);
nor U7804 (N_7804,N_3637,N_2117);
xnor U7805 (N_7805,N_1693,N_3450);
and U7806 (N_7806,N_3330,N_1721);
nor U7807 (N_7807,N_15,N_1674);
or U7808 (N_7808,N_1711,N_409);
and U7809 (N_7809,N_357,N_914);
and U7810 (N_7810,N_2908,N_1380);
and U7811 (N_7811,N_3953,N_417);
nor U7812 (N_7812,N_952,N_3106);
and U7813 (N_7813,N_901,N_1545);
and U7814 (N_7814,N_2628,N_3607);
xor U7815 (N_7815,N_2410,N_1919);
nand U7816 (N_7816,N_2520,N_692);
or U7817 (N_7817,N_3742,N_1817);
nor U7818 (N_7818,N_2071,N_3529);
nor U7819 (N_7819,N_2064,N_3994);
nand U7820 (N_7820,N_224,N_258);
or U7821 (N_7821,N_805,N_2932);
nand U7822 (N_7822,N_1513,N_709);
nor U7823 (N_7823,N_2496,N_3761);
nand U7824 (N_7824,N_385,N_3851);
or U7825 (N_7825,N_1613,N_2936);
nor U7826 (N_7826,N_1823,N_150);
or U7827 (N_7827,N_1777,N_2178);
and U7828 (N_7828,N_94,N_2444);
xnor U7829 (N_7829,N_3814,N_673);
or U7830 (N_7830,N_2782,N_2868);
nand U7831 (N_7831,N_1791,N_2465);
nand U7832 (N_7832,N_1758,N_1104);
nand U7833 (N_7833,N_2852,N_2317);
nor U7834 (N_7834,N_2689,N_3786);
and U7835 (N_7835,N_1117,N_1595);
nand U7836 (N_7836,N_3651,N_2719);
nor U7837 (N_7837,N_1244,N_2922);
xor U7838 (N_7838,N_3119,N_3257);
nand U7839 (N_7839,N_382,N_2144);
xor U7840 (N_7840,N_2773,N_3768);
nor U7841 (N_7841,N_1403,N_3639);
or U7842 (N_7842,N_214,N_3662);
xnor U7843 (N_7843,N_2509,N_2837);
or U7844 (N_7844,N_2640,N_2778);
nor U7845 (N_7845,N_3954,N_471);
or U7846 (N_7846,N_495,N_1543);
nand U7847 (N_7847,N_3954,N_2923);
nor U7848 (N_7848,N_1933,N_1294);
nand U7849 (N_7849,N_1158,N_3725);
and U7850 (N_7850,N_1170,N_282);
nor U7851 (N_7851,N_395,N_767);
nand U7852 (N_7852,N_3717,N_991);
or U7853 (N_7853,N_2766,N_1408);
nor U7854 (N_7854,N_3745,N_919);
nand U7855 (N_7855,N_1637,N_427);
and U7856 (N_7856,N_2056,N_624);
and U7857 (N_7857,N_2756,N_1733);
or U7858 (N_7858,N_221,N_558);
or U7859 (N_7859,N_2243,N_881);
and U7860 (N_7860,N_2291,N_2743);
nand U7861 (N_7861,N_3676,N_2143);
nor U7862 (N_7862,N_1855,N_2439);
or U7863 (N_7863,N_375,N_676);
and U7864 (N_7864,N_2892,N_3426);
xnor U7865 (N_7865,N_3690,N_2408);
nand U7866 (N_7866,N_1150,N_1082);
nand U7867 (N_7867,N_3937,N_2096);
or U7868 (N_7868,N_3159,N_935);
and U7869 (N_7869,N_26,N_474);
or U7870 (N_7870,N_2879,N_2471);
or U7871 (N_7871,N_257,N_2805);
nand U7872 (N_7872,N_34,N_2598);
or U7873 (N_7873,N_3648,N_507);
nor U7874 (N_7874,N_2684,N_1281);
nand U7875 (N_7875,N_245,N_2618);
or U7876 (N_7876,N_1524,N_381);
nand U7877 (N_7877,N_1981,N_2411);
or U7878 (N_7878,N_2078,N_632);
nand U7879 (N_7879,N_482,N_620);
or U7880 (N_7880,N_2694,N_1499);
and U7881 (N_7881,N_2378,N_2706);
nand U7882 (N_7882,N_1987,N_3600);
nor U7883 (N_7883,N_1997,N_870);
xnor U7884 (N_7884,N_3516,N_3667);
xnor U7885 (N_7885,N_3053,N_2558);
nand U7886 (N_7886,N_2690,N_1619);
nand U7887 (N_7887,N_1020,N_3414);
and U7888 (N_7888,N_1071,N_3362);
or U7889 (N_7889,N_3435,N_375);
and U7890 (N_7890,N_3575,N_3476);
and U7891 (N_7891,N_774,N_2947);
nand U7892 (N_7892,N_178,N_932);
nand U7893 (N_7893,N_1684,N_3487);
nand U7894 (N_7894,N_2787,N_3041);
nand U7895 (N_7895,N_43,N_3503);
and U7896 (N_7896,N_2556,N_276);
nand U7897 (N_7897,N_196,N_670);
xnor U7898 (N_7898,N_93,N_415);
and U7899 (N_7899,N_3976,N_515);
xor U7900 (N_7900,N_2375,N_181);
xnor U7901 (N_7901,N_1305,N_115);
nand U7902 (N_7902,N_335,N_2221);
and U7903 (N_7903,N_960,N_1247);
nor U7904 (N_7904,N_3783,N_2131);
and U7905 (N_7905,N_3385,N_821);
nand U7906 (N_7906,N_1196,N_1996);
xor U7907 (N_7907,N_1906,N_432);
or U7908 (N_7908,N_2235,N_1260);
nand U7909 (N_7909,N_1829,N_711);
nand U7910 (N_7910,N_37,N_2742);
nand U7911 (N_7911,N_3475,N_2729);
nand U7912 (N_7912,N_314,N_2210);
and U7913 (N_7913,N_332,N_3770);
or U7914 (N_7914,N_2984,N_719);
or U7915 (N_7915,N_728,N_3605);
nor U7916 (N_7916,N_16,N_3891);
nor U7917 (N_7917,N_1368,N_1767);
nand U7918 (N_7918,N_860,N_3484);
nand U7919 (N_7919,N_2404,N_3101);
nand U7920 (N_7920,N_1257,N_523);
nand U7921 (N_7921,N_638,N_289);
nand U7922 (N_7922,N_1987,N_2489);
nor U7923 (N_7923,N_2397,N_3148);
nor U7924 (N_7924,N_620,N_2775);
nor U7925 (N_7925,N_1524,N_1151);
or U7926 (N_7926,N_2234,N_2276);
nor U7927 (N_7927,N_1808,N_3674);
or U7928 (N_7928,N_3956,N_519);
and U7929 (N_7929,N_1566,N_1824);
or U7930 (N_7930,N_1041,N_909);
and U7931 (N_7931,N_809,N_3112);
and U7932 (N_7932,N_2175,N_3877);
nand U7933 (N_7933,N_2784,N_3826);
nor U7934 (N_7934,N_2185,N_3070);
nor U7935 (N_7935,N_2985,N_304);
xor U7936 (N_7936,N_1441,N_352);
nand U7937 (N_7937,N_2054,N_1028);
or U7938 (N_7938,N_424,N_3813);
and U7939 (N_7939,N_2589,N_2032);
xor U7940 (N_7940,N_3429,N_1283);
nand U7941 (N_7941,N_770,N_2234);
nor U7942 (N_7942,N_1972,N_1990);
nor U7943 (N_7943,N_1699,N_1840);
nand U7944 (N_7944,N_2761,N_3846);
nand U7945 (N_7945,N_1006,N_1922);
or U7946 (N_7946,N_1308,N_3317);
nand U7947 (N_7947,N_840,N_3496);
nand U7948 (N_7948,N_3081,N_3425);
nand U7949 (N_7949,N_1045,N_1310);
xor U7950 (N_7950,N_1354,N_1454);
or U7951 (N_7951,N_465,N_719);
nor U7952 (N_7952,N_435,N_777);
or U7953 (N_7953,N_1290,N_211);
nor U7954 (N_7954,N_41,N_116);
xor U7955 (N_7955,N_2848,N_3788);
or U7956 (N_7956,N_3720,N_3102);
nand U7957 (N_7957,N_2665,N_2949);
and U7958 (N_7958,N_1577,N_2476);
and U7959 (N_7959,N_3705,N_3417);
and U7960 (N_7960,N_1232,N_572);
or U7961 (N_7961,N_1694,N_3668);
nand U7962 (N_7962,N_1257,N_2728);
or U7963 (N_7963,N_2572,N_1370);
nand U7964 (N_7964,N_3747,N_430);
nand U7965 (N_7965,N_2552,N_1457);
nor U7966 (N_7966,N_63,N_3835);
nand U7967 (N_7967,N_3601,N_598);
or U7968 (N_7968,N_275,N_945);
and U7969 (N_7969,N_2722,N_3487);
nor U7970 (N_7970,N_3696,N_2031);
and U7971 (N_7971,N_1051,N_1271);
and U7972 (N_7972,N_3578,N_3590);
or U7973 (N_7973,N_3942,N_390);
nand U7974 (N_7974,N_3800,N_2079);
nand U7975 (N_7975,N_3015,N_517);
nand U7976 (N_7976,N_3731,N_1154);
nand U7977 (N_7977,N_3118,N_2171);
nand U7978 (N_7978,N_1449,N_2810);
or U7979 (N_7979,N_1422,N_40);
nand U7980 (N_7980,N_3322,N_1975);
xor U7981 (N_7981,N_660,N_778);
nand U7982 (N_7982,N_3523,N_1342);
nand U7983 (N_7983,N_1664,N_1624);
nand U7984 (N_7984,N_1060,N_760);
nor U7985 (N_7985,N_3532,N_2017);
or U7986 (N_7986,N_2754,N_102);
or U7987 (N_7987,N_2932,N_2164);
xnor U7988 (N_7988,N_1897,N_2173);
and U7989 (N_7989,N_1078,N_1496);
nor U7990 (N_7990,N_3680,N_3438);
or U7991 (N_7991,N_3142,N_442);
or U7992 (N_7992,N_3758,N_1352);
nor U7993 (N_7993,N_939,N_3542);
nor U7994 (N_7994,N_3076,N_2388);
xor U7995 (N_7995,N_3943,N_3296);
and U7996 (N_7996,N_457,N_261);
nor U7997 (N_7997,N_2711,N_1945);
nor U7998 (N_7998,N_2869,N_3348);
nor U7999 (N_7999,N_3479,N_3761);
nand U8000 (N_8000,N_5712,N_7321);
nand U8001 (N_8001,N_4548,N_5865);
and U8002 (N_8002,N_6261,N_4260);
nor U8003 (N_8003,N_4246,N_7594);
nand U8004 (N_8004,N_6477,N_7922);
nand U8005 (N_8005,N_6746,N_4638);
and U8006 (N_8006,N_5192,N_5351);
or U8007 (N_8007,N_4608,N_6404);
or U8008 (N_8008,N_7012,N_6945);
or U8009 (N_8009,N_4201,N_5056);
or U8010 (N_8010,N_7401,N_7505);
nand U8011 (N_8011,N_4499,N_4739);
or U8012 (N_8012,N_5738,N_4685);
nand U8013 (N_8013,N_5264,N_5105);
and U8014 (N_8014,N_7875,N_6664);
nor U8015 (N_8015,N_7059,N_6509);
and U8016 (N_8016,N_4082,N_4004);
nand U8017 (N_8017,N_6081,N_6745);
and U8018 (N_8018,N_4288,N_5224);
nor U8019 (N_8019,N_4470,N_6764);
or U8020 (N_8020,N_4182,N_7013);
nand U8021 (N_8021,N_4071,N_5500);
nand U8022 (N_8022,N_5068,N_6326);
or U8023 (N_8023,N_4196,N_5281);
nand U8024 (N_8024,N_5615,N_5377);
nor U8025 (N_8025,N_4407,N_7710);
or U8026 (N_8026,N_6559,N_4338);
nand U8027 (N_8027,N_7280,N_7530);
and U8028 (N_8028,N_6085,N_6075);
nor U8029 (N_8029,N_5783,N_5528);
or U8030 (N_8030,N_5510,N_6990);
nor U8031 (N_8031,N_4994,N_6044);
nor U8032 (N_8032,N_7291,N_7999);
nor U8033 (N_8033,N_4213,N_7735);
or U8034 (N_8034,N_5019,N_4653);
nand U8035 (N_8035,N_6388,N_7090);
nand U8036 (N_8036,N_4589,N_4275);
nor U8037 (N_8037,N_7623,N_6293);
nand U8038 (N_8038,N_7770,N_6489);
and U8039 (N_8039,N_6137,N_7340);
nor U8040 (N_8040,N_4403,N_4237);
xnor U8041 (N_8041,N_5532,N_5853);
or U8042 (N_8042,N_5075,N_6316);
or U8043 (N_8043,N_4755,N_5246);
nand U8044 (N_8044,N_4840,N_4610);
nand U8045 (N_8045,N_5529,N_4358);
nor U8046 (N_8046,N_5168,N_7435);
xor U8047 (N_8047,N_6178,N_4846);
or U8048 (N_8048,N_7158,N_6063);
and U8049 (N_8049,N_6949,N_4981);
xnor U8050 (N_8050,N_5496,N_5256);
xnor U8051 (N_8051,N_4224,N_6280);
nand U8052 (N_8052,N_6049,N_6046);
nand U8053 (N_8053,N_4666,N_5342);
xnor U8054 (N_8054,N_7440,N_7602);
nor U8055 (N_8055,N_4208,N_7124);
or U8056 (N_8056,N_5521,N_5164);
and U8057 (N_8057,N_6629,N_5597);
and U8058 (N_8058,N_5625,N_6740);
and U8059 (N_8059,N_7860,N_4335);
nor U8060 (N_8060,N_6970,N_4724);
nor U8061 (N_8061,N_4423,N_7891);
nand U8062 (N_8062,N_7094,N_7589);
xnor U8063 (N_8063,N_7600,N_6121);
nor U8064 (N_8064,N_5462,N_7498);
or U8065 (N_8065,N_7266,N_4058);
and U8066 (N_8066,N_4662,N_4342);
nand U8067 (N_8067,N_5209,N_7077);
nand U8068 (N_8068,N_4329,N_5405);
nand U8069 (N_8069,N_7564,N_6129);
and U8070 (N_8070,N_7842,N_6573);
or U8071 (N_8071,N_4523,N_6311);
or U8072 (N_8072,N_5852,N_7264);
nor U8073 (N_8073,N_7986,N_7847);
nand U8074 (N_8074,N_5727,N_7822);
nor U8075 (N_8075,N_4787,N_5449);
or U8076 (N_8076,N_7328,N_7753);
and U8077 (N_8077,N_6766,N_7349);
and U8078 (N_8078,N_6038,N_5763);
and U8079 (N_8079,N_4028,N_7415);
nand U8080 (N_8080,N_6636,N_6959);
and U8081 (N_8081,N_6184,N_4131);
nor U8082 (N_8082,N_5686,N_5578);
and U8083 (N_8083,N_7631,N_6756);
nor U8084 (N_8084,N_4216,N_5034);
and U8085 (N_8085,N_7980,N_6267);
or U8086 (N_8086,N_4581,N_6268);
or U8087 (N_8087,N_4207,N_6774);
nor U8088 (N_8088,N_7320,N_4868);
and U8089 (N_8089,N_5593,N_5653);
or U8090 (N_8090,N_7252,N_4545);
nor U8091 (N_8091,N_5459,N_6017);
and U8092 (N_8092,N_7299,N_5990);
and U8093 (N_8093,N_5309,N_4247);
nand U8094 (N_8094,N_6103,N_4191);
nand U8095 (N_8095,N_7899,N_7816);
nor U8096 (N_8096,N_7987,N_6929);
or U8097 (N_8097,N_5797,N_4178);
nand U8098 (N_8098,N_6466,N_5822);
nor U8099 (N_8099,N_4331,N_7197);
nor U8100 (N_8100,N_5675,N_5910);
nand U8101 (N_8101,N_4042,N_5243);
nor U8102 (N_8102,N_7443,N_6961);
or U8103 (N_8103,N_7595,N_4929);
or U8104 (N_8104,N_5298,N_6066);
nor U8105 (N_8105,N_7040,N_6521);
nand U8106 (N_8106,N_6177,N_6741);
or U8107 (N_8107,N_4026,N_4534);
nor U8108 (N_8108,N_6626,N_6885);
and U8109 (N_8109,N_5173,N_7927);
nand U8110 (N_8110,N_4007,N_6158);
nand U8111 (N_8111,N_4549,N_6187);
and U8112 (N_8112,N_7356,N_7783);
xnor U8113 (N_8113,N_7955,N_5607);
nor U8114 (N_8114,N_7615,N_5466);
nand U8115 (N_8115,N_7931,N_5894);
nand U8116 (N_8116,N_6455,N_5965);
and U8117 (N_8117,N_5713,N_4038);
and U8118 (N_8118,N_5219,N_4965);
nand U8119 (N_8119,N_5914,N_5308);
or U8120 (N_8120,N_6068,N_6878);
nor U8121 (N_8121,N_4832,N_6348);
and U8122 (N_8122,N_7620,N_5217);
nor U8123 (N_8123,N_5488,N_7430);
and U8124 (N_8124,N_4629,N_5334);
or U8125 (N_8125,N_7640,N_7337);
nor U8126 (N_8126,N_4798,N_6433);
nor U8127 (N_8127,N_4094,N_7063);
nand U8128 (N_8128,N_7103,N_5489);
nor U8129 (N_8129,N_7400,N_7871);
and U8130 (N_8130,N_7187,N_5268);
and U8131 (N_8131,N_7684,N_5467);
nand U8132 (N_8132,N_6880,N_5533);
nor U8133 (N_8133,N_4886,N_6033);
or U8134 (N_8134,N_6580,N_5670);
xnor U8135 (N_8135,N_4673,N_6381);
nor U8136 (N_8136,N_4044,N_7976);
and U8137 (N_8137,N_5399,N_7627);
nand U8138 (N_8138,N_5933,N_4463);
and U8139 (N_8139,N_4884,N_7186);
nand U8140 (N_8140,N_7593,N_5674);
or U8141 (N_8141,N_6804,N_4343);
and U8142 (N_8142,N_6201,N_4993);
or U8143 (N_8143,N_6667,N_6142);
and U8144 (N_8144,N_5960,N_6834);
nand U8145 (N_8145,N_7730,N_6993);
nand U8146 (N_8146,N_7511,N_6550);
nor U8147 (N_8147,N_5747,N_6757);
nor U8148 (N_8148,N_5288,N_5958);
nand U8149 (N_8149,N_6242,N_4823);
and U8150 (N_8150,N_6452,N_5320);
nor U8151 (N_8151,N_6493,N_7675);
nand U8152 (N_8152,N_5723,N_4515);
and U8153 (N_8153,N_5983,N_7000);
nand U8154 (N_8154,N_4264,N_4458);
or U8155 (N_8155,N_4778,N_4544);
xnor U8156 (N_8156,N_5296,N_7901);
and U8157 (N_8157,N_5711,N_4507);
nor U8158 (N_8158,N_7765,N_6344);
or U8159 (N_8159,N_4771,N_7062);
nand U8160 (N_8160,N_4266,N_6064);
and U8161 (N_8161,N_5354,N_6868);
or U8162 (N_8162,N_4114,N_7178);
nor U8163 (N_8163,N_5913,N_4604);
nor U8164 (N_8164,N_7801,N_6045);
or U8165 (N_8165,N_5031,N_5132);
nor U8166 (N_8166,N_7236,N_5680);
nand U8167 (N_8167,N_5574,N_5795);
nand U8168 (N_8168,N_4133,N_5819);
xnor U8169 (N_8169,N_6728,N_7874);
nand U8170 (N_8170,N_6875,N_7611);
xor U8171 (N_8171,N_7935,N_7778);
or U8172 (N_8172,N_4256,N_5641);
or U8173 (N_8173,N_5315,N_6445);
and U8174 (N_8174,N_7429,N_4424);
nor U8175 (N_8175,N_6652,N_5370);
nand U8176 (N_8176,N_6405,N_5906);
nand U8177 (N_8177,N_4913,N_5468);
or U8178 (N_8178,N_7669,N_6974);
and U8179 (N_8179,N_4933,N_6671);
or U8180 (N_8180,N_7172,N_5773);
nand U8181 (N_8181,N_7231,N_4811);
and U8182 (N_8182,N_5430,N_5474);
or U8183 (N_8183,N_4102,N_7664);
and U8184 (N_8184,N_5052,N_7348);
nand U8185 (N_8185,N_7475,N_4719);
nor U8186 (N_8186,N_5194,N_6858);
nor U8187 (N_8187,N_6851,N_7542);
nand U8188 (N_8188,N_5142,N_5411);
and U8189 (N_8189,N_7395,N_4992);
and U8190 (N_8190,N_5935,N_5427);
or U8191 (N_8191,N_7943,N_7466);
and U8192 (N_8192,N_7556,N_7764);
or U8193 (N_8193,N_5214,N_5276);
nor U8194 (N_8194,N_4824,N_4974);
nand U8195 (N_8195,N_6313,N_6659);
nor U8196 (N_8196,N_6727,N_4030);
xnor U8197 (N_8197,N_6004,N_6911);
xor U8198 (N_8198,N_7306,N_6128);
or U8199 (N_8199,N_4002,N_5972);
xor U8200 (N_8200,N_4758,N_5051);
or U8201 (N_8201,N_7723,N_7112);
and U8202 (N_8202,N_7016,N_6848);
or U8203 (N_8203,N_5361,N_6801);
nand U8204 (N_8204,N_7212,N_5606);
xnor U8205 (N_8205,N_7681,N_4128);
and U8206 (N_8206,N_4779,N_4391);
or U8207 (N_8207,N_4437,N_4351);
or U8208 (N_8208,N_7536,N_5678);
or U8209 (N_8209,N_4144,N_4495);
nand U8210 (N_8210,N_7362,N_6341);
xnor U8211 (N_8211,N_6503,N_6333);
and U8212 (N_8212,N_6428,N_6748);
nand U8213 (N_8213,N_7833,N_4226);
or U8214 (N_8214,N_4000,N_6174);
and U8215 (N_8215,N_4326,N_4765);
and U8216 (N_8216,N_6853,N_5555);
and U8217 (N_8217,N_7119,N_7687);
nand U8218 (N_8218,N_7984,N_4177);
and U8219 (N_8219,N_5832,N_5324);
or U8220 (N_8220,N_5175,N_4679);
nand U8221 (N_8221,N_4878,N_6214);
xor U8222 (N_8222,N_4921,N_5321);
xnor U8223 (N_8223,N_7583,N_6950);
nor U8224 (N_8224,N_7581,N_6586);
or U8225 (N_8225,N_6170,N_5450);
xor U8226 (N_8226,N_6546,N_6976);
and U8227 (N_8227,N_6624,N_7422);
xor U8228 (N_8228,N_4917,N_5022);
and U8229 (N_8229,N_6207,N_6401);
or U8230 (N_8230,N_7585,N_7323);
nand U8231 (N_8231,N_4530,N_5242);
and U8232 (N_8232,N_5486,N_7128);
and U8233 (N_8233,N_5750,N_5921);
or U8234 (N_8234,N_6013,N_7161);
nand U8235 (N_8235,N_5305,N_7192);
nand U8236 (N_8236,N_5098,N_6031);
nand U8237 (N_8237,N_4942,N_5067);
nand U8238 (N_8238,N_6377,N_4429);
nor U8239 (N_8239,N_6930,N_7480);
nor U8240 (N_8240,N_7707,N_5721);
and U8241 (N_8241,N_6903,N_5918);
xnor U8242 (N_8242,N_5250,N_7477);
or U8243 (N_8243,N_4257,N_4928);
and U8244 (N_8244,N_5543,N_4242);
nand U8245 (N_8245,N_4789,N_4962);
nand U8246 (N_8246,N_6818,N_6233);
nor U8247 (N_8247,N_5801,N_5549);
and U8248 (N_8248,N_6844,N_5681);
or U8249 (N_8249,N_6651,N_7425);
nor U8250 (N_8250,N_5930,N_7274);
nand U8251 (N_8251,N_5915,N_4215);
or U8252 (N_8252,N_7727,N_4672);
or U8253 (N_8253,N_7771,N_5538);
nor U8254 (N_8254,N_5688,N_7529);
nor U8255 (N_8255,N_7567,N_7642);
nand U8256 (N_8256,N_6159,N_4436);
nand U8257 (N_8257,N_6850,N_4756);
nand U8258 (N_8258,N_4899,N_4217);
nand U8259 (N_8259,N_7363,N_5603);
nor U8260 (N_8260,N_4946,N_6355);
or U8261 (N_8261,N_6827,N_5041);
nand U8262 (N_8262,N_7796,N_4788);
and U8263 (N_8263,N_6361,N_5842);
nor U8264 (N_8264,N_4931,N_7700);
and U8265 (N_8265,N_5338,N_6935);
and U8266 (N_8266,N_4891,N_4851);
nor U8267 (N_8267,N_5698,N_4912);
or U8268 (N_8268,N_5774,N_7919);
or U8269 (N_8269,N_7933,N_7058);
nand U8270 (N_8270,N_7882,N_6977);
or U8271 (N_8271,N_7867,N_5900);
nand U8272 (N_8272,N_5493,N_7499);
xnor U8273 (N_8273,N_7702,N_7939);
nor U8274 (N_8274,N_5277,N_5248);
nor U8275 (N_8275,N_5078,N_6135);
and U8276 (N_8276,N_6524,N_4564);
nor U8277 (N_8277,N_6857,N_5882);
nor U8278 (N_8278,N_4949,N_6003);
nand U8279 (N_8279,N_7590,N_6584);
or U8280 (N_8280,N_6587,N_5089);
nor U8281 (N_8281,N_4618,N_5013);
nand U8282 (N_8282,N_5151,N_5285);
or U8283 (N_8283,N_7985,N_6092);
nand U8284 (N_8284,N_5981,N_7803);
nor U8285 (N_8285,N_4444,N_5854);
nand U8286 (N_8286,N_6471,N_6581);
nor U8287 (N_8287,N_4095,N_5350);
nand U8288 (N_8288,N_5835,N_7402);
or U8289 (N_8289,N_5456,N_5708);
nand U8290 (N_8290,N_4076,N_6676);
or U8291 (N_8291,N_7247,N_5509);
and U8292 (N_8292,N_6026,N_4220);
nor U8293 (N_8293,N_7731,N_7864);
nor U8294 (N_8294,N_4729,N_4843);
and U8295 (N_8295,N_4790,N_5647);
nor U8296 (N_8296,N_5109,N_7513);
and U8297 (N_8297,N_5352,N_7746);
xor U8298 (N_8298,N_6492,N_5153);
and U8299 (N_8299,N_4100,N_5679);
nor U8300 (N_8300,N_6653,N_5663);
nand U8301 (N_8301,N_4054,N_6001);
nand U8302 (N_8302,N_4737,N_4218);
and U8303 (N_8303,N_6924,N_6324);
nor U8304 (N_8304,N_4117,N_6702);
nor U8305 (N_8305,N_6752,N_5064);
xor U8306 (N_8306,N_4035,N_7944);
or U8307 (N_8307,N_5279,N_5623);
nor U8308 (N_8308,N_5416,N_7175);
nor U8309 (N_8309,N_5793,N_4835);
and U8310 (N_8310,N_6148,N_7827);
nand U8311 (N_8311,N_7526,N_4193);
xor U8312 (N_8312,N_6622,N_6803);
or U8313 (N_8313,N_7460,N_4920);
and U8314 (N_8314,N_7390,N_5152);
xnor U8315 (N_8315,N_6419,N_4171);
and U8316 (N_8316,N_6271,N_7879);
or U8317 (N_8317,N_6755,N_6450);
or U8318 (N_8318,N_5568,N_4289);
nor U8319 (N_8319,N_6287,N_5146);
or U8320 (N_8320,N_5785,N_6206);
nand U8321 (N_8321,N_7146,N_4483);
or U8322 (N_8322,N_7651,N_4923);
nor U8323 (N_8323,N_5760,N_7004);
nor U8324 (N_8324,N_7223,N_7292);
nor U8325 (N_8325,N_4582,N_5612);
or U8326 (N_8326,N_4613,N_6320);
nor U8327 (N_8327,N_5886,N_4097);
or U8328 (N_8328,N_7504,N_7604);
nand U8329 (N_8329,N_7653,N_7745);
xor U8330 (N_8330,N_5552,N_5107);
nand U8331 (N_8331,N_4989,N_4579);
xnor U8332 (N_8332,N_7354,N_5563);
or U8333 (N_8333,N_4172,N_5779);
or U8334 (N_8334,N_5893,N_6500);
nor U8335 (N_8335,N_5630,N_6364);
or U8336 (N_8336,N_5683,N_7289);
nand U8337 (N_8337,N_7497,N_6809);
and U8338 (N_8338,N_6558,N_5622);
nor U8339 (N_8339,N_6086,N_4195);
and U8340 (N_8340,N_7371,N_7540);
xnor U8341 (N_8341,N_4990,N_6495);
nor U8342 (N_8342,N_4657,N_6883);
nand U8343 (N_8343,N_5008,N_4278);
nor U8344 (N_8344,N_7085,N_4211);
or U8345 (N_8345,N_4733,N_4497);
and U8346 (N_8346,N_6016,N_6519);
or U8347 (N_8347,N_7450,N_4656);
nand U8348 (N_8348,N_6513,N_4893);
xor U8349 (N_8349,N_6877,N_6838);
or U8350 (N_8350,N_7311,N_7397);
xor U8351 (N_8351,N_7137,N_7160);
nor U8352 (N_8352,N_4642,N_7574);
or U8353 (N_8353,N_7331,N_5984);
xor U8354 (N_8354,N_5860,N_5764);
and U8355 (N_8355,N_4651,N_4048);
and U8356 (N_8356,N_7408,N_5048);
or U8357 (N_8357,N_4572,N_6662);
or U8358 (N_8358,N_5782,N_5085);
nor U8359 (N_8359,N_4189,N_6527);
nor U8360 (N_8360,N_6354,N_7214);
and U8361 (N_8361,N_4454,N_6856);
nor U8362 (N_8362,N_4438,N_5436);
nand U8363 (N_8363,N_7147,N_5551);
nor U8364 (N_8364,N_4556,N_5083);
and U8365 (N_8365,N_5144,N_5768);
nor U8366 (N_8366,N_5699,N_5891);
xnor U8367 (N_8367,N_5955,N_5505);
nand U8368 (N_8368,N_6528,N_5881);
and U8369 (N_8369,N_7367,N_4230);
or U8370 (N_8370,N_4286,N_6946);
and U8371 (N_8371,N_6523,N_5762);
and U8372 (N_8372,N_5252,N_5344);
nor U8373 (N_8373,N_6685,N_6988);
or U8374 (N_8374,N_4587,N_5635);
nand U8375 (N_8375,N_4456,N_6269);
and U8376 (N_8376,N_4280,N_7206);
nand U8377 (N_8377,N_6152,N_4379);
and U8378 (N_8378,N_7720,N_7238);
nand U8379 (N_8379,N_5788,N_6772);
nor U8380 (N_8380,N_5043,N_5957);
and U8381 (N_8381,N_4713,N_5439);
nand U8382 (N_8382,N_5784,N_6094);
xor U8383 (N_8383,N_4064,N_7350);
nor U8384 (N_8384,N_5627,N_4809);
nand U8385 (N_8385,N_5070,N_7992);
nand U8386 (N_8386,N_6231,N_4939);
xnor U8387 (N_8387,N_6140,N_5617);
nand U8388 (N_8388,N_4982,N_7237);
nand U8389 (N_8389,N_5885,N_7414);
or U8390 (N_8390,N_4205,N_7619);
or U8391 (N_8391,N_6413,N_6424);
and U8392 (N_8392,N_6668,N_5827);
or U8393 (N_8393,N_5204,N_6821);
nand U8394 (N_8394,N_7195,N_6356);
or U8395 (N_8395,N_6021,N_5065);
nor U8396 (N_8396,N_7938,N_6539);
or U8397 (N_8397,N_4732,N_7960);
nor U8398 (N_8398,N_4304,N_7934);
nor U8399 (N_8399,N_6778,N_4032);
nand U8400 (N_8400,N_6458,N_6327);
nor U8401 (N_8401,N_4985,N_4187);
or U8402 (N_8402,N_6340,N_4011);
xor U8403 (N_8403,N_6125,N_5407);
nand U8404 (N_8404,N_6217,N_6494);
and U8405 (N_8405,N_5452,N_4793);
and U8406 (N_8406,N_4726,N_5263);
nor U8407 (N_8407,N_7189,N_6947);
and U8408 (N_8408,N_6904,N_6788);
or U8409 (N_8409,N_6347,N_6808);
nor U8410 (N_8410,N_4493,N_6371);
and U8411 (N_8411,N_5036,N_4911);
xor U8412 (N_8412,N_7857,N_5304);
or U8413 (N_8413,N_7277,N_4950);
and U8414 (N_8414,N_7257,N_6162);
and U8415 (N_8415,N_4759,N_6249);
nor U8416 (N_8416,N_7767,N_7445);
nand U8417 (N_8417,N_7045,N_7819);
or U8418 (N_8418,N_5421,N_7483);
nor U8419 (N_8419,N_4749,N_6087);
nor U8420 (N_8420,N_4705,N_6168);
nand U8421 (N_8421,N_4780,N_7145);
nor U8422 (N_8422,N_4001,N_4448);
nor U8423 (N_8423,N_5471,N_6266);
or U8424 (N_8424,N_6093,N_5804);
nor U8425 (N_8425,N_5483,N_7133);
or U8426 (N_8426,N_4668,N_5870);
nor U8427 (N_8427,N_7033,N_7517);
xor U8428 (N_8428,N_7817,N_6897);
xor U8429 (N_8429,N_5463,N_6056);
nor U8430 (N_8430,N_5072,N_6035);
nand U8431 (N_8431,N_7728,N_7772);
and U8432 (N_8432,N_6108,N_4966);
nor U8433 (N_8433,N_6510,N_7360);
nand U8434 (N_8434,N_6015,N_6180);
or U8435 (N_8435,N_7557,N_7449);
nor U8436 (N_8436,N_7918,N_5948);
nand U8437 (N_8437,N_4777,N_6717);
or U8438 (N_8438,N_4163,N_7351);
nor U8439 (N_8439,N_7578,N_7151);
and U8440 (N_8440,N_6270,N_6608);
xor U8441 (N_8441,N_4664,N_7926);
and U8442 (N_8442,N_7246,N_6039);
or U8443 (N_8443,N_6363,N_5969);
or U8444 (N_8444,N_4876,N_5247);
and U8445 (N_8445,N_5582,N_7650);
or U8446 (N_8446,N_4800,N_4181);
nand U8447 (N_8447,N_5709,N_5063);
nor U8448 (N_8448,N_5476,N_4748);
or U8449 (N_8449,N_6606,N_5672);
nor U8450 (N_8450,N_4400,N_5267);
nand U8451 (N_8451,N_6790,N_4746);
nand U8452 (N_8452,N_7853,N_5403);
nor U8453 (N_8453,N_7163,N_5831);
or U8454 (N_8454,N_4111,N_5047);
xor U8455 (N_8455,N_6545,N_7658);
nor U8456 (N_8456,N_6654,N_5049);
and U8457 (N_8457,N_7873,N_7895);
or U8458 (N_8458,N_5671,N_6005);
xnor U8459 (N_8459,N_6609,N_4791);
and U8460 (N_8460,N_4482,N_7794);
or U8461 (N_8461,N_4369,N_7506);
or U8462 (N_8462,N_6576,N_7129);
and U8463 (N_8463,N_6783,N_4015);
nand U8464 (N_8464,N_4339,N_7203);
or U8465 (N_8465,N_4816,N_7598);
nand U8466 (N_8466,N_7198,N_5038);
and U8467 (N_8467,N_6127,N_6952);
nor U8468 (N_8468,N_6058,N_7263);
nand U8469 (N_8469,N_6516,N_4754);
and U8470 (N_8470,N_4362,N_7296);
nand U8471 (N_8471,N_6010,N_4807);
xnor U8472 (N_8472,N_7607,N_6175);
nand U8473 (N_8473,N_5238,N_6585);
and U8474 (N_8474,N_6720,N_4644);
nand U8475 (N_8475,N_5585,N_6724);
and U8476 (N_8476,N_4873,N_7486);
and U8477 (N_8477,N_7271,N_7758);
or U8478 (N_8478,N_6318,N_5758);
nor U8479 (N_8479,N_7152,N_6050);
or U8480 (N_8480,N_6711,N_6597);
or U8481 (N_8481,N_7659,N_7314);
xnor U8482 (N_8482,N_7208,N_4970);
or U8483 (N_8483,N_4055,N_7887);
nand U8484 (N_8484,N_4248,N_5249);
xor U8485 (N_8485,N_4874,N_7005);
nor U8486 (N_8486,N_6973,N_7890);
nor U8487 (N_8487,N_6053,N_6688);
and U8488 (N_8488,N_5447,N_6721);
nor U8489 (N_8489,N_5702,N_6866);
or U8490 (N_8490,N_5824,N_6379);
and U8491 (N_8491,N_4848,N_7714);
xnor U8492 (N_8492,N_7718,N_7079);
or U8493 (N_8493,N_7057,N_5943);
or U8494 (N_8494,N_4730,N_6917);
or U8495 (N_8495,N_5260,N_4822);
and U8496 (N_8496,N_7126,N_6637);
nand U8497 (N_8497,N_5490,N_6060);
nor U8498 (N_8498,N_5274,N_5970);
xnor U8499 (N_8499,N_6157,N_5556);
or U8500 (N_8500,N_6847,N_6700);
nor U8501 (N_8501,N_4442,N_7821);
nand U8502 (N_8502,N_4586,N_7267);
nor U8503 (N_8503,N_5689,N_4374);
nand U8504 (N_8504,N_7020,N_7806);
and U8505 (N_8505,N_5851,N_5134);
nand U8506 (N_8506,N_6468,N_6518);
and U8507 (N_8507,N_5733,N_7240);
or U8508 (N_8508,N_5423,N_6963);
nand U8509 (N_8509,N_4605,N_5618);
nand U8510 (N_8510,N_4504,N_7521);
nand U8511 (N_8511,N_4080,N_7878);
nand U8512 (N_8512,N_7643,N_7648);
or U8513 (N_8513,N_6426,N_5290);
nor U8514 (N_8514,N_4595,N_7761);
nor U8515 (N_8515,N_4623,N_6512);
nand U8516 (N_8516,N_7672,N_6762);
and U8517 (N_8517,N_7222,N_4494);
nor U8518 (N_8518,N_4795,N_5364);
and U8519 (N_8519,N_7464,N_5327);
and U8520 (N_8520,N_6234,N_6018);
and U8521 (N_8521,N_4479,N_6623);
or U8522 (N_8522,N_4892,N_7674);
xnor U8523 (N_8523,N_6384,N_4694);
nor U8524 (N_8524,N_4150,N_6467);
nor U8525 (N_8525,N_4696,N_5514);
or U8526 (N_8526,N_5378,N_7885);
nor U8527 (N_8527,N_6984,N_7582);
nand U8528 (N_8528,N_7940,N_7473);
or U8529 (N_8529,N_4075,N_6743);
nor U8530 (N_8530,N_5158,N_7951);
or U8531 (N_8531,N_4558,N_7716);
or U8532 (N_8532,N_6421,N_7793);
and U8533 (N_8533,N_4984,N_7325);
nand U8534 (N_8534,N_5292,N_4432);
and U8535 (N_8535,N_6439,N_7456);
or U8536 (N_8536,N_7113,N_7327);
or U8537 (N_8537,N_4236,N_7888);
xnor U8538 (N_8538,N_7164,N_4802);
and U8539 (N_8539,N_4706,N_4743);
and U8540 (N_8540,N_5477,N_7157);
nor U8541 (N_8541,N_5156,N_4017);
nor U8542 (N_8542,N_7162,N_4637);
and U8543 (N_8543,N_4745,N_4952);
nand U8544 (N_8544,N_4121,N_5283);
and U8545 (N_8545,N_5113,N_7549);
nor U8546 (N_8546,N_4542,N_6395);
nor U8547 (N_8547,N_7964,N_4460);
or U8548 (N_8548,N_7883,N_6082);
nand U8549 (N_8549,N_6104,N_7592);
nor U8550 (N_8550,N_7807,N_6954);
nand U8551 (N_8551,N_4488,N_7073);
or U8552 (N_8552,N_6908,N_6686);
or U8553 (N_8553,N_7234,N_6620);
xnor U8554 (N_8554,N_6474,N_4915);
or U8555 (N_8555,N_5343,N_4692);
nor U8556 (N_8556,N_6628,N_5103);
and U8557 (N_8557,N_7855,N_7584);
nand U8558 (N_8558,N_4474,N_6392);
or U8559 (N_8559,N_6096,N_5081);
nor U8560 (N_8560,N_6899,N_7990);
and U8561 (N_8561,N_4318,N_7019);
nand U8562 (N_8562,N_5461,N_4269);
and U8563 (N_8563,N_4136,N_5908);
xor U8564 (N_8564,N_6195,N_6561);
or U8565 (N_8565,N_4661,N_5029);
and U8566 (N_8566,N_6716,N_5736);
and U8567 (N_8567,N_4820,N_7524);
and U8568 (N_8568,N_5964,N_4935);
or U8569 (N_8569,N_4412,N_6696);
nand U8570 (N_8570,N_5431,N_4925);
or U8571 (N_8571,N_5179,N_4113);
nor U8572 (N_8572,N_4366,N_4297);
nor U8573 (N_8573,N_4066,N_7032);
and U8574 (N_8574,N_4258,N_7712);
nand U8575 (N_8575,N_5867,N_4634);
or U8576 (N_8576,N_6487,N_5319);
or U8577 (N_8577,N_4227,N_5588);
nor U8578 (N_8578,N_4684,N_6120);
nand U8579 (N_8579,N_6694,N_7127);
nand U8580 (N_8580,N_6109,N_6002);
and U8581 (N_8581,N_7239,N_6193);
or U8582 (N_8582,N_5642,N_7176);
and U8583 (N_8583,N_5464,N_4049);
and U8584 (N_8584,N_6505,N_7996);
nor U8585 (N_8585,N_5237,N_4522);
and U8586 (N_8586,N_6274,N_4654);
xnor U8587 (N_8587,N_7039,N_6566);
xnor U8588 (N_8588,N_5602,N_5752);
and U8589 (N_8589,N_5880,N_4197);
and U8590 (N_8590,N_6220,N_5810);
and U8591 (N_8591,N_5759,N_4203);
or U8592 (N_8592,N_4910,N_6029);
xor U8593 (N_8593,N_7225,N_7150);
nand U8594 (N_8594,N_5731,N_5554);
or U8595 (N_8595,N_6633,N_5371);
or U8596 (N_8596,N_5201,N_4022);
and U8597 (N_8597,N_7558,N_4519);
nand U8598 (N_8598,N_5222,N_5492);
nor U8599 (N_8599,N_5748,N_6981);
nor U8600 (N_8600,N_7546,N_6223);
xnor U8601 (N_8601,N_6806,N_5655);
or U8602 (N_8602,N_7491,N_4239);
xnor U8603 (N_8603,N_5143,N_7114);
and U8604 (N_8604,N_5005,N_5188);
nor U8605 (N_8605,N_5262,N_6779);
and U8606 (N_8606,N_6726,N_6683);
nand U8607 (N_8607,N_5323,N_7869);
and U8608 (N_8608,N_7722,N_5728);
nor U8609 (N_8609,N_4360,N_4550);
or U8610 (N_8610,N_7319,N_6131);
or U8611 (N_8611,N_7101,N_5130);
nand U8612 (N_8612,N_6909,N_4068);
nand U8613 (N_8613,N_5876,N_7089);
or U8614 (N_8614,N_4413,N_7553);
nand U8615 (N_8615,N_6331,N_5245);
or U8616 (N_8616,N_6607,N_5775);
or U8617 (N_8617,N_4574,N_6396);
or U8618 (N_8618,N_7988,N_4430);
xnor U8619 (N_8619,N_6777,N_7135);
nand U8620 (N_8620,N_6943,N_5772);
and U8621 (N_8621,N_4089,N_4593);
xor U8622 (N_8622,N_4842,N_4417);
and U8623 (N_8623,N_4650,N_5902);
or U8624 (N_8624,N_5947,N_7125);
and U8625 (N_8625,N_6964,N_4079);
or U8626 (N_8626,N_7110,N_7838);
and U8627 (N_8627,N_7393,N_6329);
nor U8628 (N_8628,N_7965,N_7006);
or U8629 (N_8629,N_4821,N_5565);
or U8630 (N_8630,N_4869,N_7193);
xor U8631 (N_8631,N_5258,N_7696);
and U8632 (N_8632,N_5437,N_6596);
or U8633 (N_8633,N_6887,N_7523);
and U8634 (N_8634,N_6101,N_4986);
nor U8635 (N_8635,N_7748,N_5996);
nand U8636 (N_8636,N_6936,N_6958);
or U8637 (N_8637,N_5682,N_5751);
nor U8638 (N_8638,N_6669,N_4639);
and U8639 (N_8639,N_6376,N_6831);
nand U8640 (N_8640,N_6643,N_7957);
and U8641 (N_8641,N_7322,N_7616);
nor U8642 (N_8642,N_4158,N_6453);
nor U8643 (N_8643,N_5926,N_7601);
and U8644 (N_8644,N_4419,N_6613);
and U8645 (N_8645,N_7202,N_7762);
nand U8646 (N_8646,N_7898,N_7034);
and U8647 (N_8647,N_6473,N_7799);
nor U8648 (N_8648,N_6353,N_4881);
and U8649 (N_8649,N_4074,N_6410);
nand U8650 (N_8650,N_6257,N_4861);
or U8651 (N_8651,N_7784,N_5061);
or U8652 (N_8652,N_7115,N_4462);
nand U8653 (N_8653,N_6310,N_7647);
or U8654 (N_8654,N_7353,N_6130);
or U8655 (N_8655,N_5503,N_5718);
or U8656 (N_8656,N_6009,N_5223);
nand U8657 (N_8657,N_5090,N_5724);
and U8658 (N_8658,N_4699,N_7385);
nand U8659 (N_8659,N_6955,N_4296);
nand U8660 (N_8660,N_6083,N_4640);
or U8661 (N_8661,N_5975,N_5030);
nor U8662 (N_8662,N_7398,N_7387);
nor U8663 (N_8663,N_7610,N_7682);
nand U8664 (N_8664,N_4914,N_6497);
and U8665 (N_8665,N_5742,N_4168);
and U8666 (N_8666,N_7141,N_7250);
xnor U8667 (N_8667,N_7382,N_4728);
nor U8668 (N_8668,N_4954,N_6572);
nor U8669 (N_8669,N_6674,N_4397);
or U8670 (N_8670,N_7269,N_4212);
or U8671 (N_8671,N_6718,N_6432);
or U8672 (N_8672,N_6744,N_6677);
nor U8673 (N_8673,N_6248,N_6239);
and U8674 (N_8674,N_5954,N_6932);
and U8675 (N_8675,N_6071,N_5730);
and U8676 (N_8676,N_5383,N_7043);
and U8677 (N_8677,N_4371,N_6434);
nor U8678 (N_8678,N_4406,N_7453);
or U8679 (N_8679,N_5055,N_6107);
and U8680 (N_8680,N_5613,N_5390);
nor U8681 (N_8681,N_4622,N_4781);
nand U8682 (N_8682,N_7457,N_6116);
nor U8683 (N_8683,N_5368,N_7573);
and U8684 (N_8684,N_4760,N_7302);
or U8685 (N_8685,N_4169,N_7276);
and U8686 (N_8686,N_5306,N_6544);
nand U8687 (N_8687,N_4120,N_7913);
nor U8688 (N_8688,N_5301,N_7220);
nor U8689 (N_8689,N_6383,N_4901);
or U8690 (N_8690,N_5695,N_4021);
nor U8691 (N_8691,N_4206,N_6338);
nand U8692 (N_8692,N_7035,N_4710);
nor U8693 (N_8693,N_7142,N_6975);
or U8694 (N_8694,N_7199,N_6143);
and U8695 (N_8695,N_5167,N_7841);
nor U8696 (N_8696,N_4782,N_7446);
or U8697 (N_8697,N_6095,N_7974);
and U8698 (N_8698,N_4894,N_7537);
and U8699 (N_8699,N_7975,N_4877);
or U8700 (N_8700,N_4336,N_4819);
nor U8701 (N_8701,N_6461,N_7575);
nand U8702 (N_8702,N_6709,N_4088);
xor U8703 (N_8703,N_4667,N_4092);
or U8704 (N_8704,N_4827,N_6861);
or U8705 (N_8705,N_6812,N_4741);
or U8706 (N_8706,N_6731,N_7338);
and U8707 (N_8707,N_6784,N_7886);
or U8708 (N_8708,N_6186,N_5725);
nand U8709 (N_8709,N_4138,N_7489);
or U8710 (N_8710,N_4389,N_6701);
and U8711 (N_8711,N_4200,N_5904);
nor U8712 (N_8712,N_6618,N_4505);
nand U8713 (N_8713,N_5363,N_4533);
xnor U8714 (N_8714,N_7946,N_4775);
and U8715 (N_8715,N_4231,N_4972);
and U8716 (N_8716,N_7066,N_4971);
xnor U8717 (N_8717,N_7143,N_5690);
or U8718 (N_8718,N_7279,N_6000);
and U8719 (N_8719,N_6925,N_4398);
and U8720 (N_8720,N_4531,N_6385);
or U8721 (N_8721,N_5392,N_5202);
nor U8722 (N_8722,N_7431,N_7268);
nand U8723 (N_8723,N_7412,N_6479);
nand U8724 (N_8724,N_7704,N_5207);
nand U8725 (N_8725,N_7774,N_5621);
nor U8726 (N_8726,N_6564,N_5203);
nor U8727 (N_8727,N_5897,N_4599);
or U8728 (N_8728,N_7865,N_4955);
xor U8729 (N_8729,N_4799,N_5646);
nand U8730 (N_8730,N_5924,N_5187);
nor U8731 (N_8731,N_7516,N_5811);
nor U8732 (N_8732,N_4305,N_6161);
xor U8733 (N_8733,N_6118,N_4126);
xor U8734 (N_8734,N_7810,N_4090);
or U8735 (N_8735,N_4508,N_7389);
nand U8736 (N_8736,N_6910,N_7973);
nor U8737 (N_8737,N_4520,N_6454);
nor U8738 (N_8738,N_7636,N_7868);
nor U8739 (N_8739,N_5453,N_4784);
nor U8740 (N_8740,N_6598,N_5261);
nand U8741 (N_8741,N_7352,N_7185);
nand U8742 (N_8742,N_4689,N_6994);
or U8743 (N_8743,N_6279,N_7733);
and U8744 (N_8744,N_7906,N_6956);
or U8745 (N_8745,N_6188,N_4166);
and U8746 (N_8746,N_7686,N_6167);
nand U8747 (N_8747,N_7538,N_5084);
nor U8748 (N_8748,N_6146,N_7165);
or U8749 (N_8749,N_5189,N_4941);
nor U8750 (N_8750,N_7153,N_7394);
nor U8751 (N_8751,N_5629,N_6264);
and U8752 (N_8752,N_7182,N_5927);
nand U8753 (N_8753,N_6616,N_7293);
nor U8754 (N_8754,N_6867,N_4850);
nand U8755 (N_8755,N_5413,N_6486);
or U8756 (N_8756,N_7297,N_6942);
or U8757 (N_8757,N_7872,N_7078);
nor U8758 (N_8758,N_6872,N_4880);
or U8759 (N_8759,N_4624,N_5544);
and U8760 (N_8760,N_7782,N_4521);
nand U8761 (N_8761,N_7587,N_6533);
or U8762 (N_8762,N_7916,N_4561);
nand U8763 (N_8763,N_5226,N_5346);
nand U8764 (N_8764,N_7002,N_7968);
or U8765 (N_8765,N_6828,N_5211);
nand U8766 (N_8766,N_7031,N_6308);
xor U8767 (N_8767,N_5949,N_4233);
nor U8768 (N_8768,N_6951,N_7562);
or U8769 (N_8769,N_6967,N_4188);
nand U8770 (N_8770,N_7342,N_6641);
nand U8771 (N_8771,N_7470,N_4222);
nor U8772 (N_8772,N_7436,N_7630);
nor U8773 (N_8773,N_7074,N_4447);
nor U8774 (N_8774,N_4281,N_5208);
nor U8775 (N_8775,N_5393,N_4223);
nand U8776 (N_8776,N_5410,N_4062);
and U8777 (N_8777,N_5215,N_6845);
xnor U8778 (N_8778,N_5572,N_7937);
xnor U8779 (N_8779,N_7694,N_4135);
or U8780 (N_8780,N_6065,N_7433);
nor U8781 (N_8781,N_7003,N_6871);
nor U8782 (N_8782,N_4353,N_5482);
nand U8783 (N_8783,N_6230,N_5454);
and U8784 (N_8784,N_5438,N_5542);
or U8785 (N_8785,N_4484,N_7755);
nor U8786 (N_8786,N_5767,N_7649);
and U8787 (N_8787,N_4686,N_4979);
or U8788 (N_8788,N_6548,N_6678);
and U8789 (N_8789,N_7358,N_4645);
nand U8790 (N_8790,N_6884,N_5938);
or U8791 (N_8791,N_7329,N_5172);
nand U8792 (N_8792,N_4023,N_7295);
and U8793 (N_8793,N_7586,N_4426);
or U8794 (N_8794,N_7166,N_4776);
or U8795 (N_8795,N_5180,N_6940);
nor U8796 (N_8796,N_4895,N_6603);
and U8797 (N_8797,N_5362,N_5523);
and U8798 (N_8798,N_6747,N_4578);
or U8799 (N_8799,N_6285,N_7335);
or U8800 (N_8800,N_7050,N_5023);
nor U8801 (N_8801,N_6281,N_7029);
and U8802 (N_8802,N_7304,N_4711);
xnor U8803 (N_8803,N_5967,N_7849);
nand U8804 (N_8804,N_7467,N_7318);
or U8805 (N_8805,N_7792,N_4043);
xnor U8806 (N_8806,N_6415,N_5905);
or U8807 (N_8807,N_4047,N_6819);
nand U8808 (N_8808,N_7472,N_7705);
or U8809 (N_8809,N_7942,N_6611);
and U8810 (N_8810,N_6182,N_4130);
and U8811 (N_8811,N_4927,N_4161);
and U8812 (N_8812,N_5987,N_4443);
nand U8813 (N_8813,N_5701,N_4633);
or U8814 (N_8814,N_4332,N_6789);
or U8815 (N_8815,N_5859,N_6569);
and U8816 (N_8816,N_5406,N_5050);
nand U8817 (N_8817,N_4630,N_6169);
nand U8818 (N_8818,N_4801,N_6916);
or U8819 (N_8819,N_4715,N_4018);
or U8820 (N_8820,N_6189,N_5460);
nand U8821 (N_8821,N_6814,N_4421);
and U8822 (N_8822,N_6440,N_4404);
or U8823 (N_8823,N_4467,N_5901);
nand U8824 (N_8824,N_4378,N_7481);
xor U8825 (N_8825,N_7815,N_7671);
and U8826 (N_8826,N_5857,N_5559);
and U8827 (N_8827,N_6771,N_5340);
or U8828 (N_8828,N_6089,N_5009);
or U8829 (N_8829,N_7249,N_5212);
or U8830 (N_8830,N_6714,N_6530);
or U8831 (N_8831,N_7326,N_5633);
or U8832 (N_8832,N_6881,N_7365);
or U8833 (N_8833,N_4722,N_5332);
nand U8834 (N_8834,N_6644,N_5257);
nor U8835 (N_8835,N_5704,N_4009);
nor U8836 (N_8836,N_4372,N_5080);
or U8837 (N_8837,N_4767,N_6672);
xor U8838 (N_8838,N_7966,N_6735);
xor U8839 (N_8839,N_5911,N_7495);
nand U8840 (N_8840,N_4936,N_7566);
nor U8841 (N_8841,N_4948,N_5592);
nor U8842 (N_8842,N_5524,N_5353);
and U8843 (N_8843,N_6164,N_6782);
nor U8844 (N_8844,N_7027,N_4024);
nand U8845 (N_8845,N_6097,N_5548);
or U8846 (N_8846,N_5118,N_7420);
xnor U8847 (N_8847,N_6796,N_6407);
nor U8848 (N_8848,N_5147,N_4959);
nor U8849 (N_8849,N_5020,N_4720);
xor U8850 (N_8850,N_6478,N_6681);
or U8851 (N_8851,N_5210,N_7554);
nand U8852 (N_8852,N_7184,N_5959);
nor U8853 (N_8853,N_5185,N_7963);
xnor U8854 (N_8854,N_5799,N_6250);
nand U8855 (N_8855,N_5837,N_4900);
and U8856 (N_8856,N_5826,N_4409);
nor U8857 (N_8857,N_6240,N_7309);
or U8858 (N_8858,N_4384,N_6794);
xor U8859 (N_8859,N_4688,N_7177);
xor U8860 (N_8860,N_6837,N_5191);
nor U8861 (N_8861,N_5769,N_4446);
nor U8862 (N_8862,N_5269,N_4277);
nor U8863 (N_8863,N_5841,N_6582);
nand U8864 (N_8864,N_4073,N_5316);
nor U8865 (N_8865,N_5444,N_6054);
xnor U8866 (N_8866,N_6807,N_7386);
or U8867 (N_8867,N_4439,N_7285);
xor U8868 (N_8868,N_5878,N_6816);
and U8869 (N_8869,N_6699,N_4052);
and U8870 (N_8870,N_6173,N_5418);
and U8871 (N_8871,N_4317,N_4245);
and U8872 (N_8872,N_7482,N_5550);
and U8873 (N_8873,N_6321,N_6055);
and U8874 (N_8874,N_5515,N_6091);
nand U8875 (N_8875,N_6197,N_7854);
nor U8876 (N_8876,N_5576,N_4600);
nand U8877 (N_8877,N_7288,N_6560);
nor U8878 (N_8878,N_6589,N_7149);
nand U8879 (N_8879,N_7978,N_6914);
nand U8880 (N_8880,N_4804,N_6194);
nor U8881 (N_8881,N_7880,N_5235);
and U8882 (N_8882,N_4887,N_4451);
nor U8883 (N_8883,N_6425,N_6430);
nor U8884 (N_8884,N_7282,N_5808);
or U8885 (N_8885,N_5737,N_6591);
or U8886 (N_8886,N_7970,N_7201);
nor U8887 (N_8887,N_4267,N_5435);
and U8888 (N_8888,N_6823,N_5575);
or U8889 (N_8889,N_5170,N_5534);
nor U8890 (N_8890,N_7122,N_5384);
and U8891 (N_8891,N_6715,N_4511);
or U8892 (N_8892,N_6499,N_5117);
nor U8893 (N_8893,N_7242,N_5001);
or U8894 (N_8894,N_5650,N_7417);
nand U8895 (N_8895,N_4453,N_4571);
or U8896 (N_8896,N_5169,N_7219);
or U8897 (N_8897,N_4290,N_4768);
xnor U8898 (N_8898,N_5424,N_7995);
nor U8899 (N_8899,N_6057,N_6219);
nor U8900 (N_8900,N_5121,N_5213);
nand U8901 (N_8901,N_5286,N_6926);
nor U8902 (N_8902,N_5570,N_6299);
nor U8903 (N_8903,N_4466,N_4380);
nor U8904 (N_8904,N_6708,N_7979);
nand U8905 (N_8905,N_5385,N_4477);
nor U8906 (N_8906,N_6222,N_5166);
xnor U8907 (N_8907,N_7454,N_5003);
and U8908 (N_8908,N_6457,N_4697);
nor U8909 (N_8909,N_5805,N_4148);
nand U8910 (N_8910,N_5806,N_5059);
nor U8911 (N_8911,N_7075,N_5526);
or U8912 (N_8912,N_4411,N_4553);
or U8913 (N_8913,N_6792,N_6705);
nor U8914 (N_8914,N_4860,N_7708);
nor U8915 (N_8915,N_7605,N_5006);
nor U8916 (N_8916,N_5786,N_4858);
or U8917 (N_8917,N_5159,N_4602);
xor U8918 (N_8918,N_5787,N_4098);
xor U8919 (N_8919,N_4324,N_4951);
or U8920 (N_8920,N_4998,N_4736);
and U8921 (N_8921,N_6382,N_4830);
nor U8922 (N_8922,N_5912,N_5873);
xnor U8923 (N_8923,N_6275,N_7346);
xnor U8924 (N_8924,N_7426,N_5726);
nor U8925 (N_8925,N_5953,N_4879);
nand U8926 (N_8926,N_7028,N_7972);
nand U8927 (N_8927,N_6244,N_6575);
nor U8928 (N_8928,N_6088,N_6588);
or U8929 (N_8929,N_5251,N_7923);
nor U8930 (N_8930,N_4938,N_7917);
and U8931 (N_8931,N_6166,N_6665);
nand U8932 (N_8932,N_7448,N_5928);
nor U8933 (N_8933,N_6179,N_4480);
or U8934 (N_8934,N_6100,N_5977);
and U8935 (N_8935,N_4159,N_5497);
nand U8936 (N_8936,N_6391,N_6022);
and U8937 (N_8937,N_4234,N_5883);
nand U8938 (N_8938,N_6625,N_7629);
nor U8939 (N_8939,N_7909,N_5000);
nor U8940 (N_8940,N_4792,N_5148);
and U8941 (N_8941,N_6542,N_6563);
xor U8942 (N_8942,N_5703,N_6854);
or U8943 (N_8943,N_6552,N_6833);
nor U8944 (N_8944,N_4487,N_7776);
or U8945 (N_8945,N_5190,N_6879);
nor U8946 (N_8946,N_5445,N_5599);
nand U8947 (N_8947,N_5330,N_6515);
xnor U8948 (N_8948,N_6446,N_4687);
nand U8949 (N_8949,N_4678,N_4723);
or U8950 (N_8950,N_7211,N_5216);
nor U8951 (N_8951,N_5687,N_7908);
and U8952 (N_8952,N_7844,N_5896);
nand U8953 (N_8953,N_6387,N_5093);
nor U8954 (N_8954,N_7652,N_4344);
xor U8955 (N_8955,N_5478,N_6294);
xnor U8956 (N_8956,N_4674,N_4402);
and U8957 (N_8957,N_7915,N_5026);
nand U8958 (N_8958,N_4340,N_4156);
and U8959 (N_8959,N_6398,N_4116);
or U8960 (N_8960,N_7463,N_7155);
nor U8961 (N_8961,N_7026,N_4302);
and U8962 (N_8962,N_7655,N_5807);
nand U8963 (N_8963,N_6359,N_7777);
nor U8964 (N_8964,N_4810,N_5856);
and U8965 (N_8965,N_5066,N_7685);
xor U8966 (N_8966,N_7565,N_6754);
and U8967 (N_8967,N_5386,N_6380);
nand U8968 (N_8968,N_4244,N_7967);
or U8969 (N_8969,N_5951,N_6334);
and U8970 (N_8970,N_6218,N_7754);
and U8971 (N_8971,N_7088,N_5163);
nand U8972 (N_8972,N_5137,N_4376);
nand U8973 (N_8973,N_5271,N_7752);
or U8974 (N_8974,N_6076,N_4747);
or U8975 (N_8975,N_4041,N_5241);
and U8976 (N_8976,N_6902,N_5923);
and U8977 (N_8977,N_5982,N_5666);
nor U8978 (N_8978,N_7478,N_6781);
nor U8979 (N_8979,N_7461,N_5253);
and U8980 (N_8980,N_5171,N_5501);
nor U8981 (N_8981,N_5934,N_5302);
nor U8982 (N_8982,N_6488,N_6614);
and U8983 (N_8983,N_4890,N_4859);
nor U8984 (N_8984,N_4383,N_6966);
nor U8985 (N_8985,N_6444,N_5796);
nand U8986 (N_8986,N_5348,N_6070);
nor U8987 (N_8987,N_5669,N_6139);
nand U8988 (N_8988,N_5451,N_4255);
nor U8989 (N_8989,N_5817,N_7493);
or U8990 (N_8990,N_4518,N_7048);
and U8991 (N_8991,N_7531,N_5183);
and U8992 (N_8992,N_7379,N_4763);
nand U8993 (N_8993,N_4870,N_7894);
nor U8994 (N_8994,N_4445,N_6619);
and U8995 (N_8995,N_4149,N_4096);
or U8996 (N_8996,N_5126,N_4857);
and U8997 (N_8997,N_7049,N_7121);
and U8998 (N_8998,N_7484,N_6181);
and U8999 (N_8999,N_5259,N_4420);
nand U9000 (N_9000,N_6639,N_7725);
nand U9001 (N_9001,N_5971,N_4926);
nand U9002 (N_9002,N_7496,N_5999);
xnor U9003 (N_9003,N_5589,N_4839);
nor U9004 (N_9004,N_5746,N_6397);
nor U9005 (N_9005,N_5553,N_4875);
or U9006 (N_9006,N_5355,N_6894);
nand U9007 (N_9007,N_4395,N_7030);
and U9008 (N_9008,N_7547,N_5614);
xnor U9009 (N_9009,N_6941,N_4157);
or U9010 (N_9010,N_6309,N_5749);
and U9011 (N_9011,N_5527,N_5944);
nor U9012 (N_9012,N_4037,N_7808);
or U9013 (N_9013,N_6541,N_6111);
nor U9014 (N_9014,N_4320,N_5099);
or U9015 (N_9015,N_4845,N_5499);
nor U9016 (N_9016,N_5766,N_4347);
nand U9017 (N_9017,N_5382,N_7375);
or U9018 (N_9018,N_6490,N_5858);
nor U9019 (N_9019,N_6780,N_7210);
nand U9020 (N_9020,N_7618,N_4770);
or U9021 (N_9021,N_4491,N_7055);
nor U9022 (N_9022,N_7539,N_7001);
or U9023 (N_9023,N_4510,N_4349);
xnor U9024 (N_9024,N_4167,N_7948);
nand U9025 (N_9025,N_4872,N_7852);
xor U9026 (N_9026,N_6890,N_6006);
nor U9027 (N_9027,N_6763,N_5404);
or U9028 (N_9028,N_7775,N_6995);
or U9029 (N_9029,N_5339,N_7876);
nor U9030 (N_9030,N_7010,N_7698);
xnor U9031 (N_9031,N_5925,N_5102);
nor U9032 (N_9032,N_7527,N_7076);
and U9033 (N_9033,N_7315,N_7545);
nor U9034 (N_9034,N_7954,N_5945);
nand U9035 (N_9035,N_7552,N_4418);
or U9036 (N_9036,N_6939,N_4410);
xor U9037 (N_9037,N_6506,N_5843);
or U9038 (N_9038,N_4132,N_6706);
or U9039 (N_9039,N_4031,N_7333);
nand U9040 (N_9040,N_4364,N_6339);
nor U9041 (N_9041,N_6144,N_7097);
nor U9042 (N_9042,N_6163,N_6437);
xnor U9043 (N_9043,N_6431,N_4968);
nor U9044 (N_9044,N_5012,N_4573);
nand U9045 (N_9045,N_7503,N_7637);
nand U9046 (N_9046,N_4478,N_6041);
xnor U9047 (N_9047,N_4590,N_5336);
nand U9048 (N_9048,N_4005,N_5649);
nand U9049 (N_9049,N_6825,N_4057);
or U9050 (N_9050,N_7416,N_6011);
nand U9051 (N_9051,N_5356,N_5922);
and U9052 (N_9052,N_7579,N_7233);
and U9053 (N_9053,N_4119,N_4253);
and U9054 (N_9054,N_7863,N_5402);
nand U9055 (N_9055,N_6992,N_5033);
xor U9056 (N_9056,N_5284,N_4864);
xnor U9057 (N_9057,N_7228,N_4053);
nand U9058 (N_9058,N_6697,N_6570);
nor U9059 (N_9059,N_7200,N_6742);
and U9060 (N_9060,N_4352,N_6888);
nor U9061 (N_9061,N_7324,N_7091);
or U9062 (N_9062,N_6427,N_7699);
nor U9063 (N_9063,N_4828,N_7111);
nor U9064 (N_9064,N_4625,N_6028);
nand U9065 (N_9065,N_6839,N_5697);
or U9066 (N_9066,N_4937,N_4902);
or U9067 (N_9067,N_6402,N_6375);
or U9068 (N_9068,N_5771,N_7756);
nand U9069 (N_9069,N_5420,N_5743);
nor U9070 (N_9070,N_4753,N_4575);
or U9071 (N_9071,N_7459,N_5366);
and U9072 (N_9072,N_7661,N_5015);
and U9073 (N_9073,N_4265,N_7900);
or U9074 (N_9074,N_7087,N_5639);
xnor U9075 (N_9075,N_7991,N_4153);
and U9076 (N_9076,N_6390,N_6416);
or U9077 (N_9077,N_6295,N_6124);
or U9078 (N_9078,N_7850,N_7645);
nor U9079 (N_9079,N_7275,N_6155);
nand U9080 (N_9080,N_5604,N_6110);
nand U9081 (N_9081,N_4509,N_4742);
nand U9082 (N_9082,N_6052,N_6978);
and U9083 (N_9083,N_5218,N_7406);
xor U9084 (N_9084,N_4069,N_6251);
nor U9085 (N_9085,N_6122,N_4295);
xor U9086 (N_9086,N_5094,N_5376);
nand U9087 (N_9087,N_7692,N_4251);
and U9088 (N_9088,N_6346,N_7889);
or U9089 (N_9089,N_5178,N_5694);
or U9090 (N_9090,N_5517,N_6459);
nand U9091 (N_9091,N_6775,N_4885);
and U9092 (N_9092,N_4580,N_4072);
and U9093 (N_9093,N_5129,N_5198);
and U9094 (N_9094,N_6737,N_4808);
nor U9095 (N_9095,N_4228,N_7998);
nor U9096 (N_9096,N_5729,N_4261);
and U9097 (N_9097,N_4769,N_4498);
xor U9098 (N_9098,N_4794,N_7788);
or U9099 (N_9099,N_5270,N_6864);
or U9100 (N_9100,N_5868,N_5594);
or U9101 (N_9101,N_4147,N_7877);
and U9102 (N_9102,N_6522,N_4174);
nor U9103 (N_9103,N_4862,N_7100);
and U9104 (N_9104,N_6835,N_6019);
and U9105 (N_9105,N_4337,N_7779);
and U9106 (N_9106,N_7294,N_5705);
nor U9107 (N_9107,N_4975,N_6208);
and U9108 (N_9108,N_6198,N_7308);
nand U9109 (N_9109,N_4905,N_7568);
nand U9110 (N_9110,N_5136,N_6319);
nor U9111 (N_9111,N_7588,N_7042);
and U9112 (N_9112,N_6507,N_4546);
nand U9113 (N_9113,N_5479,N_7548);
nor U9114 (N_9114,N_7763,N_6928);
or U9115 (N_9115,N_7227,N_6209);
nand U9116 (N_9116,N_4285,N_5676);
nand U9117 (N_9117,N_6829,N_7823);
or U9118 (N_9118,N_5632,N_4486);
and U9119 (N_9119,N_6335,N_4270);
nor U9120 (N_9120,N_5890,N_7407);
nor U9121 (N_9121,N_6918,N_6481);
or U9122 (N_9122,N_7800,N_4457);
nor U9123 (N_9123,N_5161,N_4489);
or U9124 (N_9124,N_6859,N_7181);
or U9125 (N_9125,N_5300,N_4606);
and U9126 (N_9126,N_6722,N_4727);
nand U9127 (N_9127,N_5275,N_4170);
nor U9128 (N_9128,N_7654,N_7518);
and U9129 (N_9129,N_6891,N_7444);
xor U9130 (N_9130,N_5184,N_7543);
and U9131 (N_9131,N_5266,N_4152);
or U9132 (N_9132,N_5076,N_7508);
and U9133 (N_9133,N_7286,N_4173);
and U9134 (N_9134,N_6343,N_4655);
nand U9135 (N_9135,N_6491,N_6769);
and U9136 (N_9136,N_7571,N_7232);
and U9137 (N_9137,N_6798,N_4060);
nand U9138 (N_9138,N_5637,N_5776);
and U9139 (N_9139,N_4309,N_6126);
nor U9140 (N_9140,N_4866,N_7082);
or U9141 (N_9141,N_5299,N_7805);
and U9142 (N_9142,N_4888,N_7829);
or U9143 (N_9143,N_7834,N_7797);
and U9144 (N_9144,N_6350,N_6296);
nor U9145 (N_9145,N_6215,N_6695);
and U9146 (N_9146,N_7635,N_7205);
nor U9147 (N_9147,N_4341,N_4660);
and U9148 (N_9148,N_4263,N_7502);
or U9149 (N_9149,N_6660,N_7747);
and U9150 (N_9150,N_6462,N_5100);
xnor U9151 (N_9151,N_5638,N_4399);
or U9152 (N_9152,N_5976,N_7307);
or U9153 (N_9153,N_4896,N_4310);
or U9154 (N_9154,N_4210,N_5535);
xor U9155 (N_9155,N_6113,N_6480);
nand U9156 (N_9156,N_5401,N_5475);
and U9157 (N_9157,N_5504,N_7945);
nand U9158 (N_9158,N_4061,N_5128);
or U9159 (N_9159,N_5155,N_4919);
and U9160 (N_9160,N_7924,N_5700);
nand U9161 (N_9161,N_5531,N_6937);
nand U9162 (N_9162,N_5375,N_5608);
nand U9163 (N_9163,N_4658,N_7953);
or U9164 (N_9164,N_6042,N_7442);
nand U9165 (N_9165,N_5507,N_7392);
and U9166 (N_9166,N_7683,N_4155);
nor U9167 (N_9167,N_5863,N_4243);
nand U9168 (N_9168,N_4214,N_6289);
nor U9169 (N_9169,N_4803,N_6263);
nor U9170 (N_9170,N_4924,N_5829);
and U9171 (N_9171,N_7781,N_7832);
and U9172 (N_9172,N_7469,N_4356);
nor U9173 (N_9173,N_7740,N_4298);
nand U9174 (N_9174,N_7343,N_7920);
and U9175 (N_9175,N_7561,N_6971);
or U9176 (N_9176,N_5567,N_4940);
or U9177 (N_9177,N_6237,N_6855);
or U9178 (N_9178,N_6204,N_7434);
xor U9179 (N_9179,N_6436,N_6216);
and U9180 (N_9180,N_5087,N_7840);
and U9181 (N_9181,N_5963,N_6768);
and U9182 (N_9182,N_7438,N_4740);
or U9183 (N_9183,N_5619,N_6255);
nor U9184 (N_9184,N_6642,N_4631);
or U9185 (N_9185,N_7260,N_5396);
or U9186 (N_9186,N_5941,N_7369);
or U9187 (N_9187,N_6934,N_7053);
nand U9188 (N_9188,N_4194,N_7824);
or U9189 (N_9189,N_5004,N_4099);
or U9190 (N_9190,N_5053,N_5326);
nor U9191 (N_9191,N_6863,N_7912);
nor U9192 (N_9192,N_7492,N_4583);
or U9193 (N_9193,N_4704,N_4554);
and U9194 (N_9194,N_4503,N_7670);
or U9195 (N_9195,N_4772,N_7341);
or U9196 (N_9196,N_5440,N_6525);
and U9197 (N_9197,N_7591,N_4620);
xnor U9198 (N_9198,N_5112,N_6760);
xnor U9199 (N_9199,N_4086,N_4825);
or U9200 (N_9200,N_4455,N_4871);
nor U9201 (N_9201,N_6273,N_7140);
and U9202 (N_9202,N_6422,N_7789);
nor U9203 (N_9203,N_5820,N_4294);
nand U9204 (N_9204,N_4552,N_5487);
nand U9205 (N_9205,N_7896,N_7662);
or U9206 (N_9206,N_7345,N_6535);
xor U9207 (N_9207,N_6332,N_4034);
nand U9208 (N_9208,N_7828,N_5716);
and U9209 (N_9209,N_4311,N_7528);
or U9210 (N_9210,N_5016,N_4431);
nand U9211 (N_9211,N_4646,N_4434);
nand U9212 (N_9212,N_4773,N_6399);
nand U9213 (N_9213,N_5741,N_6684);
and U9214 (N_9214,N_4287,N_5273);
nand U9215 (N_9215,N_4922,N_6927);
or U9216 (N_9216,N_5744,N_4669);
nor U9217 (N_9217,N_6635,N_5519);
xnor U9218 (N_9218,N_6115,N_6256);
nor U9219 (N_9219,N_7080,N_5206);
or U9220 (N_9220,N_7638,N_5739);
xnor U9221 (N_9221,N_5127,N_4980);
nor U9222 (N_9222,N_6024,N_6351);
or U9223 (N_9223,N_7154,N_7044);
xnor U9224 (N_9224,N_4204,N_4192);
or U9225 (N_9225,N_5502,N_5294);
xor U9226 (N_9226,N_7597,N_6765);
or U9227 (N_9227,N_7099,N_5412);
xor U9228 (N_9228,N_6534,N_6317);
nand U9229 (N_9229,N_6556,N_6810);
or U9230 (N_9230,N_5398,N_6590);
or U9231 (N_9231,N_4229,N_5888);
nand U9232 (N_9232,N_7576,N_7070);
nand U9233 (N_9233,N_5379,N_4354);
nand U9234 (N_9234,N_7136,N_6032);
or U9235 (N_9235,N_4179,N_6403);
nand U9236 (N_9236,N_4199,N_4570);
nor U9237 (N_9237,N_6312,N_5611);
and U9238 (N_9238,N_6134,N_4906);
nand U9239 (N_9239,N_4141,N_7677);
and U9240 (N_9240,N_4078,N_4083);
nor U9241 (N_9241,N_5761,N_4735);
nor U9242 (N_9242,N_7383,N_6414);
or U9243 (N_9243,N_5313,N_6460);
and U9244 (N_9244,N_4958,N_4738);
and U9245 (N_9245,N_5929,N_5991);
xnor U9246 (N_9246,N_7191,N_4997);
nand U9247 (N_9247,N_7424,N_4250);
nor U9248 (N_9248,N_7633,N_5397);
nor U9249 (N_9249,N_4774,N_7474);
or U9250 (N_9250,N_4611,N_6358);
and U9251 (N_9251,N_6567,N_6117);
and U9252 (N_9252,N_7666,N_6112);
xor U9253 (N_9253,N_6147,N_7634);
xnor U9254 (N_9254,N_4815,N_7609);
and U9255 (N_9255,N_5394,N_5798);
nand U9256 (N_9256,N_5014,N_5530);
or U9257 (N_9257,N_5571,N_6176);
nand U9258 (N_9258,N_4591,N_5830);
nor U9259 (N_9259,N_5322,N_7930);
and U9260 (N_9260,N_5441,N_4852);
nand U9261 (N_9261,N_5255,N_7848);
or U9262 (N_9262,N_7067,N_5287);
or U9263 (N_9263,N_6553,N_7116);
nand U9264 (N_9264,N_4143,N_6802);
nand U9265 (N_9265,N_6972,N_6776);
nand U9266 (N_9266,N_5874,N_7441);
and U9267 (N_9267,N_4836,N_5380);
nor U9268 (N_9268,N_4361,N_7830);
and U9269 (N_9269,N_7278,N_5989);
nor U9270 (N_9270,N_4315,N_7646);
and U9271 (N_9271,N_4091,N_5088);
or U9272 (N_9272,N_7313,N_5988);
nor U9273 (N_9273,N_7244,N_7690);
nor U9274 (N_9274,N_6719,N_5903);
and U9275 (N_9275,N_4433,N_7717);
nor U9276 (N_9276,N_6650,N_6090);
and U9277 (N_9277,N_5429,N_5978);
and U9278 (N_9278,N_4056,N_5409);
or U9279 (N_9279,N_5469,N_7679);
nand U9280 (N_9280,N_6595,N_7628);
or U9281 (N_9281,N_6759,N_6876);
or U9282 (N_9282,N_5473,N_6483);
or U9283 (N_9283,N_6368,N_5667);
nand U9284 (N_9284,N_7243,N_4988);
nor U9285 (N_9285,N_5895,N_4496);
nor U9286 (N_9286,N_4853,N_4616);
and U9287 (N_9287,N_5395,N_5836);
and U9288 (N_9288,N_5777,N_5513);
xor U9289 (N_9289,N_4615,N_4040);
nand U9290 (N_9290,N_5869,N_7550);
nand U9291 (N_9291,N_4649,N_5060);
nand U9292 (N_9292,N_7715,N_7139);
nor U9293 (N_9293,N_4964,N_7977);
or U9294 (N_9294,N_5317,N_5595);
and U9295 (N_9295,N_5839,N_6982);
nor U9296 (N_9296,N_7812,N_6265);
nand U9297 (N_9297,N_6185,N_7196);
and U9298 (N_9298,N_7509,N_4717);
and U9299 (N_9299,N_7703,N_4987);
nand U9300 (N_9300,N_6577,N_5966);
and U9301 (N_9301,N_6360,N_7903);
and U9302 (N_9302,N_7814,N_4930);
nand U9303 (N_9303,N_4103,N_6931);
xnor U9304 (N_9304,N_6138,N_5472);
and U9305 (N_9305,N_5849,N_4357);
nor U9306 (N_9306,N_6689,N_5044);
and U9307 (N_9307,N_6406,N_6547);
and U9308 (N_9308,N_6238,N_7599);
nor U9309 (N_9309,N_4541,N_5220);
and U9310 (N_9310,N_7316,N_4259);
or U9311 (N_9311,N_4834,N_4635);
and U9312 (N_9312,N_4865,N_6172);
xor U9313 (N_9313,N_4659,N_4676);
nand U9314 (N_9314,N_6451,N_7226);
nand U9315 (N_9315,N_4137,N_7660);
xor U9316 (N_9316,N_4293,N_6627);
or U9317 (N_9317,N_7798,N_6484);
nor U9318 (N_9318,N_6901,N_5898);
or U9319 (N_9319,N_6805,N_4814);
and U9320 (N_9320,N_5979,N_4414);
nor U9321 (N_9321,N_6725,N_6862);
nor U9322 (N_9322,N_7096,N_6638);
nand U9323 (N_9323,N_5601,N_4325);
nand U9324 (N_9324,N_6156,N_5310);
or U9325 (N_9325,N_7069,N_4108);
nand U9326 (N_9326,N_4563,N_7109);
and U9327 (N_9327,N_7023,N_5221);
xor U9328 (N_9328,N_5131,N_7281);
nand U9329 (N_9329,N_4567,N_7893);
nand U9330 (N_9330,N_7259,N_7381);
or U9331 (N_9331,N_7215,N_4221);
nand U9332 (N_9332,N_7551,N_5193);
and U9333 (N_9333,N_4313,N_4619);
or U9334 (N_9334,N_5181,N_6571);
nand U9335 (N_9335,N_7218,N_6698);
or U9336 (N_9336,N_4565,N_7904);
nand U9337 (N_9337,N_7766,N_5391);
and U9338 (N_9338,N_4976,N_5845);
or U9339 (N_9339,N_7015,N_6301);
and U9340 (N_9340,N_4381,N_5426);
or U9341 (N_9341,N_6171,N_5125);
nand U9342 (N_9342,N_7384,N_7462);
xnor U9343 (N_9343,N_4670,N_5186);
and U9344 (N_9344,N_7421,N_4225);
or U9345 (N_9345,N_5569,N_7458);
or U9346 (N_9346,N_6630,N_7171);
and U9347 (N_9347,N_4140,N_5042);
nor U9348 (N_9348,N_4469,N_7476);
and U9349 (N_9349,N_6482,N_4601);
or U9350 (N_9350,N_5640,N_4105);
or U9351 (N_9351,N_5195,N_5021);
nor U9352 (N_9352,N_6084,N_5007);
nand U9353 (N_9353,N_7344,N_6447);
xor U9354 (N_9354,N_6228,N_6373);
and U9355 (N_9355,N_4525,N_6841);
and U9356 (N_9356,N_7911,N_7366);
and U9357 (N_9357,N_5579,N_5116);
and U9358 (N_9358,N_7108,N_5314);
nor U9359 (N_9359,N_7639,N_4101);
or U9360 (N_9360,N_6051,N_6703);
nor U9361 (N_9361,N_7287,N_4408);
nand U9362 (N_9362,N_6649,N_6508);
or U9363 (N_9363,N_6793,N_4416);
and U9364 (N_9364,N_6661,N_6286);
nand U9365 (N_9365,N_7515,N_6648);
nor U9366 (N_9366,N_6602,N_4956);
nor U9367 (N_9367,N_6919,N_6183);
nand U9368 (N_9368,N_7962,N_7107);
nor U9369 (N_9369,N_6145,N_5919);
or U9370 (N_9370,N_7465,N_6980);
nand U9371 (N_9371,N_5303,N_5481);
or U9372 (N_9372,N_5506,N_6393);
or U9373 (N_9373,N_7858,N_4330);
nand U9374 (N_9374,N_6886,N_6860);
and U9375 (N_9375,N_6800,N_6290);
nor U9376 (N_9376,N_5879,N_5297);
or U9377 (N_9377,N_5974,N_6555);
and U9378 (N_9378,N_4405,N_6983);
xnor U9379 (N_9379,N_7106,N_4527);
nand U9380 (N_9380,N_4314,N_4882);
nor U9381 (N_9381,N_6073,N_6357);
or U9382 (N_9382,N_4276,N_4129);
nand U9383 (N_9383,N_6969,N_7437);
nand U9384 (N_9384,N_6246,N_4070);
or U9385 (N_9385,N_6149,N_5145);
or U9386 (N_9386,N_6723,N_6229);
and U9387 (N_9387,N_7804,N_6734);
and U9388 (N_9388,N_4712,N_4016);
nor U9389 (N_9389,N_5278,N_6923);
or U9390 (N_9390,N_4175,N_5620);
xor U9391 (N_9391,N_4485,N_6865);
nor U9392 (N_9392,N_6501,N_4757);
or U9393 (N_9393,N_4046,N_4299);
nand U9394 (N_9394,N_5037,N_5328);
or U9395 (N_9395,N_5465,N_4569);
nand U9396 (N_9396,N_6824,N_4146);
nor U9397 (N_9397,N_5498,N_7544);
or U9398 (N_9398,N_6476,N_4514);
nand U9399 (N_9399,N_5986,N_5939);
and U9400 (N_9400,N_6394,N_4472);
nor U9401 (N_9401,N_5046,N_7859);
and U9402 (N_9402,N_4401,N_6791);
or U9403 (N_9403,N_5558,N_7391);
or U9404 (N_9404,N_4855,N_4818);
nand U9405 (N_9405,N_7284,N_4435);
nor U9406 (N_9406,N_7614,N_6423);
nor U9407 (N_9407,N_5657,N_7334);
and U9408 (N_9408,N_6448,N_4535);
nor U9409 (N_9409,N_7021,N_4388);
nand U9410 (N_9410,N_7051,N_5115);
or U9411 (N_9411,N_4812,N_7399);
and U9412 (N_9412,N_6079,N_7856);
and U9413 (N_9413,N_5141,N_5685);
or U9414 (N_9414,N_6298,N_5634);
nand U9415 (N_9415,N_4008,N_7144);
nor U9416 (N_9416,N_4020,N_6132);
nand U9417 (N_9417,N_5864,N_4903);
nor U9418 (N_9418,N_4045,N_4883);
nor U9419 (N_9419,N_5062,N_4983);
and U9420 (N_9420,N_4731,N_5381);
and U9421 (N_9421,N_6739,N_6417);
or U9422 (N_9422,N_4960,N_6098);
nor U9423 (N_9423,N_7956,N_7820);
nand U9424 (N_9424,N_4334,N_7713);
xnor U9425 (N_9425,N_6895,N_6514);
or U9426 (N_9426,N_5225,N_4785);
or U9427 (N_9427,N_7994,N_4909);
nor U9428 (N_9428,N_4198,N_6786);
nand U9429 (N_9429,N_6852,N_5584);
nand U9430 (N_9430,N_6557,N_4273);
nand U9431 (N_9431,N_5174,N_5135);
or U9432 (N_9432,N_5717,N_4695);
nor U9433 (N_9433,N_5347,N_6205);
nand U9434 (N_9434,N_5032,N_7018);
nor U9435 (N_9435,N_5101,N_4889);
nand U9436 (N_9436,N_6957,N_5710);
nor U9437 (N_9437,N_5596,N_6944);
nor U9438 (N_9438,N_5230,N_5139);
or U9439 (N_9439,N_5054,N_6811);
and U9440 (N_9440,N_5862,N_6693);
nor U9441 (N_9441,N_5648,N_4863);
or U9442 (N_9442,N_5834,N_5039);
nor U9443 (N_9443,N_7736,N_5887);
nor U9444 (N_9444,N_4709,N_6920);
or U9445 (N_9445,N_6673,N_7982);
or U9446 (N_9446,N_7255,N_6640);
or U9447 (N_9447,N_6621,N_7488);
nor U9448 (N_9448,N_5707,N_6733);
or U9449 (N_9449,N_7559,N_4450);
or U9450 (N_9450,N_4576,N_4663);
and U9451 (N_9451,N_6999,N_7092);
xnor U9452 (N_9452,N_7411,N_6795);
or U9453 (N_9453,N_7750,N_5196);
xnor U9454 (N_9454,N_4854,N_5656);
nor U9455 (N_9455,N_4904,N_5644);
nor U9456 (N_9456,N_6254,N_7921);
nor U9457 (N_9457,N_6882,N_6372);
or U9458 (N_9458,N_7625,N_7221);
or U9459 (N_9459,N_4190,N_4327);
and U9460 (N_9460,N_4716,N_4249);
and U9461 (N_9461,N_5889,N_7760);
nand U9462 (N_9462,N_7230,N_6061);
and U9463 (N_9463,N_4328,N_4907);
nand U9464 (N_9464,N_4012,N_7046);
or U9465 (N_9465,N_5756,N_5800);
or U9466 (N_9466,N_6578,N_7928);
xor U9467 (N_9467,N_4396,N_4084);
nor U9468 (N_9468,N_7455,N_5325);
nor U9469 (N_9469,N_6366,N_6979);
and U9470 (N_9470,N_7757,N_7068);
nand U9471 (N_9471,N_6292,N_5470);
nor U9472 (N_9472,N_6679,N_6826);
nand U9473 (N_9473,N_7216,N_4826);
nor U9474 (N_9474,N_7751,N_5566);
and U9475 (N_9475,N_5157,N_5358);
and U9476 (N_9476,N_6732,N_4500);
nand U9477 (N_9477,N_7428,N_4566);
nand U9478 (N_9478,N_6211,N_5414);
xnor U9479 (N_9479,N_5652,N_5909);
nor U9480 (N_9480,N_6463,N_4609);
or U9481 (N_9481,N_4607,N_5821);
or U9482 (N_9482,N_7622,N_7768);
nor U9483 (N_9483,N_7041,N_5095);
or U9484 (N_9484,N_6617,N_4350);
and U9485 (N_9485,N_7881,N_6315);
or U9486 (N_9486,N_6043,N_7300);
nand U9487 (N_9487,N_7330,N_6682);
nor U9488 (N_9488,N_7156,N_6540);
and U9489 (N_9489,N_4363,N_6235);
and U9490 (N_9490,N_4536,N_6059);
nor U9491 (N_9491,N_5058,N_4647);
or U9492 (N_9492,N_7168,N_6245);
nand U9493 (N_9493,N_5586,N_6276);
nor U9494 (N_9494,N_5754,N_5765);
and U9495 (N_9495,N_7056,N_7843);
nor U9496 (N_9496,N_5295,N_5123);
and U9497 (N_9497,N_5591,N_4112);
nand U9498 (N_9498,N_4106,N_5165);
and U9499 (N_9499,N_7310,N_7795);
and U9500 (N_9500,N_5318,N_5980);
nor U9501 (N_9501,N_5236,N_7060);
nand U9502 (N_9502,N_6922,N_5916);
nand U9503 (N_9503,N_7102,N_7501);
and U9504 (N_9504,N_6014,N_5541);
nand U9505 (N_9505,N_7826,N_4151);
and U9506 (N_9506,N_5176,N_5040);
or U9507 (N_9507,N_4104,N_6593);
or U9508 (N_9508,N_6418,N_4125);
nor U9509 (N_9509,N_5443,N_4300);
and U9510 (N_9510,N_4124,N_7813);
nand U9511 (N_9511,N_5790,N_5573);
or U9512 (N_9512,N_6150,N_5661);
or U9513 (N_9513,N_4934,N_5659);
or U9514 (N_9514,N_6998,N_7357);
nand U9515 (N_9515,N_7959,N_6713);
or U9516 (N_9516,N_6907,N_7721);
or U9517 (N_9517,N_6386,N_5590);
or U9518 (N_9518,N_5815,N_4813);
nor U9519 (N_9519,N_7011,N_5092);
and U9520 (N_9520,N_4427,N_5160);
nand U9521 (N_9521,N_6036,N_7298);
or U9522 (N_9522,N_7596,N_5082);
nor U9523 (N_9523,N_6203,N_7447);
nand U9524 (N_9524,N_6429,N_5636);
xnor U9525 (N_9525,N_4691,N_5104);
or U9526 (N_9526,N_5875,N_7993);
nor U9527 (N_9527,N_7024,N_4123);
or U9528 (N_9528,N_6896,N_4468);
nand U9529 (N_9529,N_6210,N_5520);
and U9530 (N_9530,N_6905,N_7118);
nor U9531 (N_9531,N_5446,N_4978);
nor U9532 (N_9532,N_6307,N_7064);
or U9533 (N_9533,N_5823,N_4750);
or U9534 (N_9534,N_7409,N_5780);
and U9535 (N_9535,N_6225,N_7697);
nand U9536 (N_9536,N_5289,N_5993);
nand U9537 (N_9537,N_4751,N_6062);
or U9538 (N_9538,N_4272,N_5946);
and U9539 (N_9539,N_5973,N_7405);
xor U9540 (N_9540,N_7617,N_6692);
or U9541 (N_9541,N_7626,N_4513);
and U9542 (N_9542,N_5794,N_4963);
or U9543 (N_9543,N_4977,N_4683);
nand U9544 (N_9544,N_7861,N_4856);
and U9545 (N_9545,N_6968,N_7418);
nand U9546 (N_9546,N_4999,N_7608);
nand U9547 (N_9547,N_4019,N_4292);
or U9548 (N_9548,N_4817,N_4957);
nor U9549 (N_9549,N_7037,N_6378);
and U9550 (N_9550,N_6675,N_6658);
nor U9551 (N_9551,N_5400,N_6799);
nor U9552 (N_9552,N_5495,N_5560);
nor U9553 (N_9553,N_4284,N_5540);
nor U9554 (N_9554,N_7866,N_5664);
nand U9555 (N_9555,N_6753,N_5522);
xor U9556 (N_9556,N_6102,N_5789);
nand U9557 (N_9557,N_4365,N_5415);
and U9558 (N_9558,N_7902,N_6199);
nor U9559 (N_9559,N_6749,N_4065);
xor U9560 (N_9560,N_7061,N_5057);
xor U9561 (N_9561,N_7261,N_7701);
nand U9562 (N_9562,N_4680,N_5111);
or U9563 (N_9563,N_5341,N_7014);
or U9564 (N_9564,N_5091,N_7818);
and U9565 (N_9565,N_6435,N_5877);
and U9566 (N_9566,N_7373,N_5994);
nor U9567 (N_9567,N_4528,N_5628);
nor U9568 (N_9568,N_6870,N_7148);
nor U9569 (N_9569,N_4543,N_4145);
nand U9570 (N_9570,N_5734,N_4764);
nand U9571 (N_9571,N_5484,N_7380);
xnor U9572 (N_9572,N_4301,N_6047);
nand U9573 (N_9573,N_4202,N_7936);
nand U9574 (N_9574,N_6464,N_5516);
nor U9575 (N_9575,N_6906,N_4142);
and U9576 (N_9576,N_7656,N_6710);
nand U9577 (N_9577,N_7580,N_6260);
or U9578 (N_9578,N_5525,N_6190);
or U9579 (N_9579,N_5069,N_4947);
nor U9580 (N_9580,N_4559,N_6074);
xnor U9581 (N_9581,N_4077,N_6212);
nor U9582 (N_9582,N_4665,N_6960);
nor U9583 (N_9583,N_6472,N_5077);
xnor U9584 (N_9584,N_5182,N_6987);
or U9585 (N_9585,N_6119,N_4991);
or U9586 (N_9586,N_6815,N_6365);
or U9587 (N_9587,N_4373,N_4718);
nor U9588 (N_9588,N_5645,N_4240);
or U9589 (N_9589,N_7093,N_4838);
or U9590 (N_9590,N_7709,N_7413);
nand U9591 (N_9591,N_7025,N_5508);
nor U9592 (N_9592,N_6691,N_7932);
nor U9593 (N_9593,N_5228,N_7839);
nand U9594 (N_9594,N_5234,N_5205);
and U9595 (N_9595,N_5840,N_4283);
nand U9596 (N_9596,N_6574,N_6443);
nor U9597 (N_9597,N_6258,N_5838);
nand U9598 (N_9598,N_4449,N_7846);
and U9599 (N_9599,N_4847,N_5114);
and U9600 (N_9600,N_4185,N_5333);
xnor U9601 (N_9601,N_7169,N_6551);
and U9602 (N_9602,N_7054,N_5937);
nor U9603 (N_9603,N_7305,N_5605);
nand U9604 (N_9604,N_7130,N_5331);
nand U9605 (N_9605,N_5714,N_5442);
or U9606 (N_9606,N_6072,N_7665);
or U9607 (N_9607,N_7676,N_7897);
or U9608 (N_9608,N_6283,N_4025);
xor U9609 (N_9609,N_7188,N_7811);
nand U9610 (N_9610,N_6511,N_4714);
nand U9611 (N_9611,N_7270,N_6330);
nor U9612 (N_9612,N_6889,N_5846);
nand U9613 (N_9613,N_7167,N_4829);
nand U9614 (N_9614,N_7009,N_7131);
and U9615 (N_9615,N_5124,N_7081);
nand U9616 (N_9616,N_7071,N_6656);
nand U9617 (N_9617,N_7283,N_4051);
xor U9618 (N_9618,N_4786,N_7719);
nand U9619 (N_9619,N_7680,N_5434);
and U9620 (N_9620,N_4490,N_6893);
nand U9621 (N_9621,N_5587,N_5950);
nor U9622 (N_9622,N_6153,N_4370);
and U9623 (N_9623,N_6832,N_4252);
xnor U9624 (N_9624,N_6106,N_5942);
nand U9625 (N_9625,N_4805,N_5812);
nand U9626 (N_9626,N_4612,N_4626);
and U9627 (N_9627,N_6820,N_6037);
and U9628 (N_9628,N_5422,N_6048);
nor U9629 (N_9629,N_6288,N_7120);
xor U9630 (N_9630,N_5740,N_4180);
and U9631 (N_9631,N_4698,N_5311);
xor U9632 (N_9632,N_6830,N_5227);
or U9633 (N_9633,N_4708,N_4440);
or U9634 (N_9634,N_5936,N_6297);
or U9635 (N_9635,N_5753,N_4033);
or U9636 (N_9636,N_5899,N_7245);
and U9637 (N_9637,N_5494,N_7862);
nor U9638 (N_9638,N_5419,N_7265);
and U9639 (N_9639,N_6900,N_6583);
or U9640 (N_9640,N_7657,N_6191);
nor U9641 (N_9641,N_7533,N_4652);
xnor U9642 (N_9642,N_4614,N_7570);
nor U9643 (N_9643,N_5802,N_5120);
or U9644 (N_9644,N_7332,N_6869);
or U9645 (N_9645,N_4597,N_5197);
or U9646 (N_9646,N_5372,N_6034);
nor U9647 (N_9647,N_5365,N_5518);
nand U9648 (N_9648,N_7791,N_6475);
xnor U9649 (N_9649,N_5265,N_6123);
nand U9650 (N_9650,N_5828,N_4734);
nand U9651 (N_9651,N_7355,N_6282);
nand U9652 (N_9652,N_6154,N_5684);
or U9653 (N_9653,N_4464,N_7534);
and U9654 (N_9654,N_7372,N_4682);
nand U9655 (N_9655,N_5809,N_5814);
nand U9656 (N_9656,N_6836,N_4898);
xnor U9657 (N_9657,N_7668,N_4598);
and U9658 (N_9658,N_4752,N_4394);
and U9659 (N_9659,N_7451,N_5359);
nand U9660 (N_9660,N_5280,N_5122);
or U9661 (N_9661,N_5995,N_6817);
nand U9662 (N_9662,N_5665,N_5177);
and U9663 (N_9663,N_6770,N_6252);
or U9664 (N_9664,N_4029,N_5491);
nor U9665 (N_9665,N_5932,N_5956);
xor U9666 (N_9666,N_4165,N_6517);
and U9667 (N_9667,N_4585,N_5329);
nor U9668 (N_9668,N_6729,N_6502);
xnor U9669 (N_9669,N_4796,N_6704);
or U9670 (N_9670,N_7947,N_7737);
nand U9671 (N_9671,N_5715,N_4867);
and U9672 (N_9672,N_6601,N_7825);
or U9673 (N_9673,N_6680,N_6562);
and U9674 (N_9674,N_4944,N_7134);
or U9675 (N_9675,N_5417,N_6666);
or U9676 (N_9676,N_6543,N_5373);
nor U9677 (N_9677,N_7905,N_5677);
nor U9678 (N_9678,N_6996,N_5546);
or U9679 (N_9679,N_5940,N_6938);
and U9680 (N_9680,N_4461,N_4367);
nand U9681 (N_9681,N_5010,N_4348);
or U9682 (N_9682,N_6202,N_5631);
or U9683 (N_9683,N_6605,N_5931);
nor U9684 (N_9684,N_7535,N_4636);
nor U9685 (N_9685,N_5557,N_7180);
xor U9686 (N_9686,N_5985,N_5307);
nor U9687 (N_9687,N_4333,N_7364);
xor U9688 (N_9688,N_6241,N_6007);
nor U9689 (N_9689,N_6236,N_4322);
nand U9690 (N_9690,N_7510,N_6874);
nor U9691 (N_9691,N_7949,N_4118);
nand U9692 (N_9692,N_4473,N_4063);
nand U9693 (N_9693,N_5992,N_7952);
nor U9694 (N_9694,N_7706,N_7072);
nor U9695 (N_9695,N_4588,N_7729);
xnor U9696 (N_9696,N_5511,N_6921);
and U9697 (N_9697,N_5035,N_5002);
nor U9698 (N_9698,N_5884,N_7086);
nand U9699 (N_9699,N_7910,N_7083);
or U9700 (N_9700,N_6751,N_7845);
and U9701 (N_9701,N_5017,N_5074);
xnor U9702 (N_9702,N_6989,N_4562);
or U9703 (N_9703,N_5349,N_4701);
nand U9704 (N_9704,N_7929,N_6913);
xnor U9705 (N_9705,N_7301,N_5872);
or U9706 (N_9706,N_5312,N_6099);
nor U9707 (N_9707,N_7235,N_6272);
nor U9708 (N_9708,N_6986,N_5583);
nor U9709 (N_9709,N_6409,N_4945);
xnor U9710 (N_9710,N_4232,N_6532);
nor U9711 (N_9711,N_6962,N_7739);
nand U9712 (N_9712,N_7500,N_4115);
nor U9713 (N_9713,N_7632,N_6400);
and U9714 (N_9714,N_4368,N_4603);
or U9715 (N_9715,N_4154,N_5997);
nor U9716 (N_9716,N_5577,N_5357);
and U9717 (N_9717,N_5660,N_4584);
xor U9718 (N_9718,N_5537,N_6730);
and U9719 (N_9719,N_5755,N_4557);
xnor U9720 (N_9720,N_7179,N_5337);
and U9721 (N_9721,N_5654,N_4127);
nor U9722 (N_9722,N_7606,N_6411);
or U9723 (N_9723,N_5662,N_6631);
and U9724 (N_9724,N_6787,N_6069);
and U9725 (N_9725,N_4183,N_5998);
or U9726 (N_9726,N_7432,N_5600);
nand U9727 (N_9727,N_7780,N_4355);
and U9728 (N_9728,N_6151,N_4797);
nand U9729 (N_9729,N_6040,N_4262);
xnor U9730 (N_9730,N_4539,N_5643);
nand U9731 (N_9731,N_4677,N_6892);
nor U9732 (N_9732,N_7950,N_5233);
or U9733 (N_9733,N_6670,N_5071);
and U9734 (N_9734,N_4506,N_4459);
xnor U9735 (N_9735,N_7790,N_7347);
nand U9736 (N_9736,N_4693,N_5745);
xnor U9737 (N_9737,N_7749,N_6707);
nand U9738 (N_9738,N_5855,N_7065);
nand U9739 (N_9739,N_4897,N_5025);
nor U9740 (N_9740,N_5624,N_4059);
nand U9741 (N_9741,N_6221,N_6687);
or U9742 (N_9742,N_7724,N_6278);
nand U9743 (N_9743,N_4806,N_4087);
or U9744 (N_9744,N_4721,N_6485);
or U9745 (N_9745,N_7376,N_4517);
nor U9746 (N_9746,N_6030,N_6469);
nor U9747 (N_9747,N_4036,N_7981);
or U9748 (N_9748,N_5293,N_7663);
nand U9749 (N_9749,N_7404,N_6612);
or U9750 (N_9750,N_6813,N_4551);
or U9751 (N_9751,N_4027,N_5200);
nand U9752 (N_9752,N_6253,N_5432);
nand U9753 (N_9753,N_7138,N_5106);
xor U9754 (N_9754,N_5458,N_4393);
or U9755 (N_9755,N_4109,N_6160);
nand U9756 (N_9756,N_6314,N_7173);
or U9757 (N_9757,N_7370,N_7787);
or U9758 (N_9758,N_7744,N_7569);
nand U9759 (N_9759,N_7541,N_4681);
or U9760 (N_9760,N_5952,N_7229);
and U9761 (N_9761,N_6647,N_5598);
nand U9762 (N_9762,N_7052,N_4013);
or U9763 (N_9763,N_5581,N_5651);
and U9764 (N_9764,N_7907,N_7248);
nand U9765 (N_9765,N_7183,N_7759);
and U9766 (N_9766,N_4916,N_5110);
nor U9767 (N_9767,N_4014,N_7667);
nand U9768 (N_9768,N_6736,N_6526);
nand U9769 (N_9769,N_6105,N_6690);
nor U9770 (N_9770,N_4134,N_4107);
and U9771 (N_9771,N_4291,N_4219);
or U9772 (N_9772,N_6537,N_4377);
xnor U9773 (N_9773,N_5833,N_5866);
nor U9774 (N_9774,N_6080,N_4932);
nand U9775 (N_9775,N_5735,N_6898);
or U9776 (N_9776,N_7507,N_6657);
and U9777 (N_9777,N_6165,N_5722);
and U9778 (N_9778,N_6610,N_5850);
and U9779 (N_9779,N_7008,N_7742);
nand U9780 (N_9780,N_5150,N_6133);
or U9781 (N_9781,N_7624,N_5668);
and U9782 (N_9782,N_5917,N_5545);
nand U9783 (N_9783,N_6200,N_7241);
nor U9784 (N_9784,N_5254,N_5229);
nor U9785 (N_9785,N_7738,N_6328);
nor U9786 (N_9786,N_5539,N_6604);
nor U9787 (N_9787,N_5140,N_6842);
or U9788 (N_9788,N_4254,N_6077);
nand U9789 (N_9789,N_6915,N_4849);
nand U9790 (N_9790,N_5792,N_7961);
and U9791 (N_9791,N_7532,N_6374);
or U9792 (N_9792,N_4555,N_4241);
or U9793 (N_9793,N_4160,N_4346);
nand U9794 (N_9794,N_6247,N_7258);
or U9795 (N_9795,N_6594,N_7339);
and U9796 (N_9796,N_7555,N_5162);
nand U9797 (N_9797,N_4003,N_7644);
or U9798 (N_9798,N_6758,N_5961);
or U9799 (N_9799,N_6438,N_5962);
or U9800 (N_9800,N_7997,N_5149);
nand U9801 (N_9801,N_5803,N_7688);
nand U9802 (N_9802,N_7941,N_7378);
nor U9803 (N_9803,N_5564,N_5448);
xor U9804 (N_9804,N_6873,N_6498);
or U9805 (N_9805,N_7272,N_4690);
and U9806 (N_9806,N_4538,N_4481);
nand U9807 (N_9807,N_4139,N_4547);
and U9808 (N_9808,N_5408,N_6712);
nor U9809 (N_9809,N_7485,N_5108);
nand U9810 (N_9810,N_7925,N_4050);
and U9811 (N_9811,N_7726,N_6345);
and U9812 (N_9812,N_4359,N_4282);
and U9813 (N_9813,N_4441,N_4010);
nor U9814 (N_9814,N_5825,N_7439);
or U9815 (N_9815,N_6262,N_4093);
xnor U9816 (N_9816,N_5369,N_5673);
nor U9817 (N_9817,N_7572,N_7732);
nor U9818 (N_9818,N_5696,N_7377);
nor U9819 (N_9819,N_7403,N_5335);
xor U9820 (N_9820,N_6291,N_4323);
nor U9821 (N_9821,N_7520,N_5818);
nor U9822 (N_9822,N_5154,N_4184);
nand U9823 (N_9823,N_6634,N_4725);
xor U9824 (N_9824,N_6912,N_7673);
nand U9825 (N_9825,N_4039,N_7132);
nand U9826 (N_9826,N_4537,N_6408);
and U9827 (N_9827,N_4996,N_5282);
nor U9828 (N_9828,N_7419,N_5692);
xor U9829 (N_9829,N_4973,N_5387);
and U9830 (N_9830,N_7254,N_6599);
nor U9831 (N_9831,N_6342,N_5861);
nand U9832 (N_9832,N_5360,N_5616);
nand U9833 (N_9833,N_4382,N_4465);
nand U9834 (N_9834,N_4492,N_4592);
nor U9835 (N_9835,N_6305,N_4122);
or U9836 (N_9836,N_6389,N_4235);
nand U9837 (N_9837,N_4908,N_6953);
or U9838 (N_9838,N_5658,N_7396);
nor U9839 (N_9839,N_4274,N_6012);
and U9840 (N_9840,N_4761,N_7410);
nand U9841 (N_9841,N_7836,N_6600);
nand U9842 (N_9842,N_7273,N_6322);
and U9843 (N_9843,N_5133,N_4577);
nor U9844 (N_9844,N_6192,N_6592);
or U9845 (N_9845,N_6496,N_6646);
or U9846 (N_9846,N_5239,N_4675);
nor U9847 (N_9847,N_7098,N_6277);
or U9848 (N_9848,N_7514,N_7490);
nor U9849 (N_9849,N_4385,N_6504);
and U9850 (N_9850,N_6531,N_7621);
nand U9851 (N_9851,N_5480,N_7047);
or U9852 (N_9852,N_4475,N_5096);
nand U9853 (N_9853,N_4844,N_6750);
nor U9854 (N_9854,N_6965,N_5706);
xnor U9855 (N_9855,N_7388,N_6336);
and U9856 (N_9856,N_5720,N_5512);
nand U9857 (N_9857,N_7971,N_4621);
and U9858 (N_9858,N_4502,N_6529);
and U9859 (N_9859,N_7769,N_7577);
nand U9860 (N_9860,N_7468,N_5086);
xor U9861 (N_9861,N_5244,N_6554);
xnor U9862 (N_9862,N_6767,N_7512);
and U9863 (N_9863,N_4632,N_7741);
or U9864 (N_9864,N_4271,N_5580);
and U9865 (N_9865,N_4918,N_7479);
nor U9866 (N_9866,N_5770,N_4707);
nand U9867 (N_9867,N_7017,N_6520);
nor U9868 (N_9868,N_7253,N_4387);
or U9869 (N_9869,N_6232,N_6645);
nand U9870 (N_9870,N_5719,N_6141);
or U9871 (N_9871,N_7969,N_6997);
or U9872 (N_9872,N_6849,N_6549);
nand U9873 (N_9873,N_6797,N_5920);
nand U9874 (N_9874,N_7117,N_7209);
and U9875 (N_9875,N_5561,N_5433);
xnor U9876 (N_9876,N_5847,N_5455);
or U9877 (N_9877,N_5907,N_4596);
and U9878 (N_9878,N_4345,N_4238);
nand U9879 (N_9879,N_4321,N_4540);
nor U9880 (N_9880,N_5388,N_7427);
and U9881 (N_9881,N_5367,N_4308);
nand U9882 (N_9882,N_4162,N_5609);
nor U9883 (N_9883,N_7773,N_7159);
nand U9884 (N_9884,N_4319,N_6224);
nor U9885 (N_9885,N_5757,N_4831);
and U9886 (N_9886,N_5138,N_5199);
nor U9887 (N_9887,N_7190,N_7983);
nor U9888 (N_9888,N_7213,N_6259);
nand U9889 (N_9889,N_6300,N_6441);
or U9890 (N_9890,N_4176,N_4476);
nand U9891 (N_9891,N_7312,N_5232);
nor U9892 (N_9892,N_7487,N_6442);
or U9893 (N_9893,N_5562,N_6008);
nand U9894 (N_9894,N_4312,N_6303);
nand U9895 (N_9895,N_4516,N_4833);
nand U9896 (N_9896,N_4969,N_7224);
or U9897 (N_9897,N_4837,N_4643);
nor U9898 (N_9898,N_6370,N_6843);
and U9899 (N_9899,N_6023,N_4425);
or U9900 (N_9900,N_6337,N_6067);
and U9901 (N_9901,N_4390,N_6349);
or U9902 (N_9902,N_7471,N_6284);
nor U9903 (N_9903,N_4783,N_7786);
nand U9904 (N_9904,N_7693,N_6196);
or U9905 (N_9905,N_4006,N_5871);
or U9906 (N_9906,N_6773,N_5231);
nor U9907 (N_9907,N_6985,N_4386);
and U9908 (N_9908,N_6412,N_7870);
and U9909 (N_9909,N_4268,N_7494);
or U9910 (N_9910,N_7368,N_7170);
nand U9911 (N_9911,N_6020,N_6663);
nand U9912 (N_9912,N_7038,N_6565);
xnor U9913 (N_9913,N_4671,N_7563);
and U9914 (N_9914,N_7194,N_6449);
nor U9915 (N_9915,N_7522,N_5345);
or U9916 (N_9916,N_4943,N_5732);
nor U9917 (N_9917,N_4512,N_6465);
xnor U9918 (N_9918,N_7711,N_4110);
nand U9919 (N_9919,N_4594,N_5781);
and U9920 (N_9920,N_5626,N_4085);
and U9921 (N_9921,N_5610,N_6470);
nand U9922 (N_9922,N_7837,N_6991);
nand U9923 (N_9923,N_5892,N_5848);
nor U9924 (N_9924,N_6846,N_7884);
nand U9925 (N_9925,N_7084,N_5291);
and U9926 (N_9926,N_7802,N_7603);
nand U9927 (N_9927,N_4415,N_5778);
nand U9928 (N_9928,N_4303,N_7734);
nand U9929 (N_9929,N_5119,N_7785);
or U9930 (N_9930,N_7958,N_5011);
or U9931 (N_9931,N_5791,N_5691);
or U9932 (N_9932,N_7105,N_6025);
and U9933 (N_9933,N_4617,N_4164);
nor U9934 (N_9934,N_7525,N_4501);
nor U9935 (N_9935,N_4306,N_4307);
nor U9936 (N_9936,N_5097,N_7251);
nor U9937 (N_9937,N_7689,N_7612);
xor U9938 (N_9938,N_4526,N_7262);
or U9939 (N_9939,N_7989,N_4279);
nor U9940 (N_9940,N_6114,N_7303);
and U9941 (N_9941,N_4209,N_6367);
nand U9942 (N_9942,N_5485,N_5536);
or U9943 (N_9943,N_7835,N_5028);
nand U9944 (N_9944,N_5425,N_5693);
or U9945 (N_9945,N_4529,N_4532);
and U9946 (N_9946,N_4392,N_7851);
xor U9947 (N_9947,N_6420,N_7641);
nand U9948 (N_9948,N_6738,N_5079);
and U9949 (N_9949,N_7256,N_4471);
nand U9950 (N_9950,N_7452,N_6325);
nor U9951 (N_9951,N_4961,N_5968);
or U9952 (N_9952,N_6227,N_4641);
nand U9953 (N_9953,N_6369,N_6761);
or U9954 (N_9954,N_7095,N_7519);
nor U9955 (N_9955,N_7007,N_6948);
nand U9956 (N_9956,N_7207,N_5374);
or U9957 (N_9957,N_6822,N_4452);
nor U9958 (N_9958,N_7374,N_7691);
nor U9959 (N_9959,N_6785,N_4524);
and U9960 (N_9960,N_6078,N_7914);
nand U9961 (N_9961,N_4560,N_7336);
and U9962 (N_9962,N_6304,N_7892);
and U9963 (N_9963,N_7423,N_4995);
or U9964 (N_9964,N_6306,N_6579);
or U9965 (N_9965,N_7290,N_4744);
nor U9966 (N_9966,N_7361,N_7678);
nand U9967 (N_9967,N_5024,N_6538);
or U9968 (N_9968,N_6655,N_5389);
or U9969 (N_9969,N_7695,N_6027);
nand U9970 (N_9970,N_4081,N_4703);
nor U9971 (N_9971,N_5045,N_5018);
and U9972 (N_9972,N_4702,N_6568);
and U9973 (N_9973,N_5844,N_4766);
xor U9974 (N_9974,N_5457,N_4627);
nand U9975 (N_9975,N_6352,N_6243);
nand U9976 (N_9976,N_4186,N_4568);
nor U9977 (N_9977,N_5073,N_4375);
or U9978 (N_9978,N_6362,N_7831);
xnor U9979 (N_9979,N_6840,N_5027);
or U9980 (N_9980,N_4316,N_7359);
or U9981 (N_9981,N_6213,N_6226);
and U9982 (N_9982,N_4067,N_6456);
or U9983 (N_9983,N_5272,N_7036);
and U9984 (N_9984,N_4422,N_4700);
nand U9985 (N_9985,N_6536,N_6933);
nand U9986 (N_9986,N_6136,N_7022);
xnor U9987 (N_9987,N_4428,N_5240);
or U9988 (N_9988,N_7560,N_6323);
or U9989 (N_9989,N_7123,N_5813);
nand U9990 (N_9990,N_4628,N_4762);
nand U9991 (N_9991,N_6632,N_4648);
and U9992 (N_9992,N_5428,N_6615);
nor U9993 (N_9993,N_6302,N_5816);
nor U9994 (N_9994,N_7217,N_7104);
xnor U9995 (N_9995,N_4967,N_7809);
nor U9996 (N_9996,N_7317,N_4841);
or U9997 (N_9997,N_7613,N_4953);
nor U9998 (N_9998,N_5547,N_7743);
nand U9999 (N_9999,N_7174,N_7204);
and U10000 (N_10000,N_5803,N_6498);
nand U10001 (N_10001,N_4502,N_7058);
and U10002 (N_10002,N_4742,N_4324);
nand U10003 (N_10003,N_6003,N_7455);
and U10004 (N_10004,N_7551,N_5174);
and U10005 (N_10005,N_5791,N_6153);
or U10006 (N_10006,N_4286,N_6247);
and U10007 (N_10007,N_4654,N_6627);
nand U10008 (N_10008,N_7820,N_6372);
nor U10009 (N_10009,N_4574,N_4945);
or U10010 (N_10010,N_7156,N_4769);
nor U10011 (N_10011,N_6139,N_4570);
nand U10012 (N_10012,N_6219,N_5488);
or U10013 (N_10013,N_5335,N_5356);
nand U10014 (N_10014,N_4532,N_5459);
or U10015 (N_10015,N_7493,N_6253);
or U10016 (N_10016,N_6563,N_4466);
or U10017 (N_10017,N_4842,N_7544);
or U10018 (N_10018,N_5174,N_7301);
and U10019 (N_10019,N_4720,N_7846);
and U10020 (N_10020,N_4154,N_5832);
nor U10021 (N_10021,N_6928,N_4587);
nand U10022 (N_10022,N_5931,N_4205);
or U10023 (N_10023,N_5056,N_5225);
and U10024 (N_10024,N_7965,N_7045);
nand U10025 (N_10025,N_4863,N_7283);
nand U10026 (N_10026,N_5819,N_7068);
or U10027 (N_10027,N_5833,N_7015);
nand U10028 (N_10028,N_7451,N_6623);
nor U10029 (N_10029,N_5948,N_7370);
nor U10030 (N_10030,N_4602,N_6082);
nand U10031 (N_10031,N_5012,N_4547);
xor U10032 (N_10032,N_5793,N_4640);
nor U10033 (N_10033,N_6893,N_6035);
nor U10034 (N_10034,N_4463,N_5410);
nand U10035 (N_10035,N_7611,N_5846);
nand U10036 (N_10036,N_5461,N_7013);
or U10037 (N_10037,N_5799,N_6274);
nor U10038 (N_10038,N_5744,N_4243);
nor U10039 (N_10039,N_6965,N_5937);
nand U10040 (N_10040,N_5265,N_6792);
nand U10041 (N_10041,N_5808,N_4750);
nor U10042 (N_10042,N_4906,N_4205);
or U10043 (N_10043,N_6987,N_4214);
nand U10044 (N_10044,N_7820,N_7504);
nor U10045 (N_10045,N_5038,N_7726);
nand U10046 (N_10046,N_7109,N_4512);
nor U10047 (N_10047,N_4424,N_4356);
nor U10048 (N_10048,N_6412,N_4990);
and U10049 (N_10049,N_6269,N_5471);
nand U10050 (N_10050,N_6968,N_5403);
nor U10051 (N_10051,N_7406,N_5434);
nor U10052 (N_10052,N_4729,N_5384);
and U10053 (N_10053,N_6619,N_4707);
nor U10054 (N_10054,N_4427,N_6804);
nor U10055 (N_10055,N_5325,N_4418);
and U10056 (N_10056,N_5174,N_6033);
and U10057 (N_10057,N_7712,N_7105);
or U10058 (N_10058,N_7991,N_4977);
and U10059 (N_10059,N_4968,N_6642);
nor U10060 (N_10060,N_7527,N_7541);
and U10061 (N_10061,N_7861,N_4944);
or U10062 (N_10062,N_6867,N_6600);
and U10063 (N_10063,N_6822,N_7934);
and U10064 (N_10064,N_4138,N_7688);
nand U10065 (N_10065,N_7356,N_6011);
nand U10066 (N_10066,N_6078,N_7975);
or U10067 (N_10067,N_7590,N_4448);
xor U10068 (N_10068,N_6761,N_4630);
or U10069 (N_10069,N_5923,N_4546);
and U10070 (N_10070,N_5957,N_7571);
nand U10071 (N_10071,N_6235,N_5146);
nand U10072 (N_10072,N_5957,N_5715);
and U10073 (N_10073,N_6990,N_4573);
nand U10074 (N_10074,N_5341,N_5798);
xnor U10075 (N_10075,N_7553,N_7579);
and U10076 (N_10076,N_4872,N_6567);
and U10077 (N_10077,N_4625,N_5011);
or U10078 (N_10078,N_6507,N_7413);
or U10079 (N_10079,N_5928,N_7077);
nor U10080 (N_10080,N_5599,N_7299);
and U10081 (N_10081,N_4493,N_4768);
or U10082 (N_10082,N_4271,N_4910);
nand U10083 (N_10083,N_6087,N_7564);
nor U10084 (N_10084,N_4326,N_7410);
nand U10085 (N_10085,N_4574,N_6069);
or U10086 (N_10086,N_5791,N_7068);
or U10087 (N_10087,N_5000,N_7459);
and U10088 (N_10088,N_5609,N_4340);
nor U10089 (N_10089,N_4246,N_5862);
nor U10090 (N_10090,N_4927,N_4239);
or U10091 (N_10091,N_6241,N_7811);
nand U10092 (N_10092,N_6277,N_6442);
and U10093 (N_10093,N_6918,N_7192);
or U10094 (N_10094,N_7413,N_5151);
nand U10095 (N_10095,N_5103,N_7324);
xnor U10096 (N_10096,N_6219,N_4245);
nor U10097 (N_10097,N_5350,N_7674);
or U10098 (N_10098,N_5112,N_5389);
and U10099 (N_10099,N_7300,N_7842);
nor U10100 (N_10100,N_7248,N_4092);
nand U10101 (N_10101,N_4231,N_4514);
nor U10102 (N_10102,N_5832,N_5464);
nor U10103 (N_10103,N_6453,N_4429);
or U10104 (N_10104,N_7360,N_7521);
and U10105 (N_10105,N_6291,N_5948);
or U10106 (N_10106,N_5244,N_4876);
nor U10107 (N_10107,N_7182,N_7691);
and U10108 (N_10108,N_6030,N_6098);
and U10109 (N_10109,N_7697,N_6718);
nand U10110 (N_10110,N_7900,N_7215);
nand U10111 (N_10111,N_6283,N_5426);
xnor U10112 (N_10112,N_5942,N_7933);
and U10113 (N_10113,N_7746,N_6523);
nor U10114 (N_10114,N_5429,N_7065);
or U10115 (N_10115,N_5953,N_6917);
and U10116 (N_10116,N_6525,N_6685);
or U10117 (N_10117,N_7764,N_5983);
nand U10118 (N_10118,N_7556,N_5184);
nand U10119 (N_10119,N_6621,N_5852);
nor U10120 (N_10120,N_6235,N_6640);
xnor U10121 (N_10121,N_5586,N_7646);
xnor U10122 (N_10122,N_4908,N_4801);
nand U10123 (N_10123,N_5592,N_6411);
nor U10124 (N_10124,N_6328,N_5229);
nand U10125 (N_10125,N_6709,N_6817);
xor U10126 (N_10126,N_7612,N_4122);
or U10127 (N_10127,N_5977,N_4694);
and U10128 (N_10128,N_7659,N_5482);
or U10129 (N_10129,N_7926,N_7900);
or U10130 (N_10130,N_5085,N_5347);
and U10131 (N_10131,N_7923,N_5807);
or U10132 (N_10132,N_5505,N_5525);
and U10133 (N_10133,N_7001,N_5500);
nor U10134 (N_10134,N_5611,N_4913);
nand U10135 (N_10135,N_7456,N_6478);
nand U10136 (N_10136,N_6808,N_5198);
and U10137 (N_10137,N_5952,N_7209);
and U10138 (N_10138,N_4381,N_6763);
nand U10139 (N_10139,N_7879,N_4046);
nand U10140 (N_10140,N_6417,N_5873);
nor U10141 (N_10141,N_4740,N_6747);
or U10142 (N_10142,N_5585,N_6637);
or U10143 (N_10143,N_5993,N_5070);
or U10144 (N_10144,N_7968,N_6794);
nand U10145 (N_10145,N_4703,N_4259);
and U10146 (N_10146,N_5186,N_7521);
or U10147 (N_10147,N_6052,N_5621);
nand U10148 (N_10148,N_4224,N_4899);
or U10149 (N_10149,N_4885,N_5007);
nand U10150 (N_10150,N_7307,N_4182);
nand U10151 (N_10151,N_4586,N_5097);
nand U10152 (N_10152,N_4504,N_6717);
nand U10153 (N_10153,N_5406,N_4593);
nor U10154 (N_10154,N_5878,N_5943);
or U10155 (N_10155,N_5564,N_6877);
or U10156 (N_10156,N_4487,N_4433);
nor U10157 (N_10157,N_6039,N_7295);
nand U10158 (N_10158,N_6549,N_5280);
nand U10159 (N_10159,N_6067,N_6379);
or U10160 (N_10160,N_4990,N_7833);
or U10161 (N_10161,N_6154,N_6888);
or U10162 (N_10162,N_5165,N_7744);
nor U10163 (N_10163,N_5428,N_6241);
xnor U10164 (N_10164,N_7776,N_4910);
and U10165 (N_10165,N_6887,N_7439);
nand U10166 (N_10166,N_7955,N_7272);
and U10167 (N_10167,N_6035,N_7875);
nor U10168 (N_10168,N_5294,N_6286);
and U10169 (N_10169,N_5104,N_5761);
nor U10170 (N_10170,N_7398,N_7527);
nor U10171 (N_10171,N_4504,N_6223);
nand U10172 (N_10172,N_5503,N_4049);
and U10173 (N_10173,N_7573,N_6131);
nand U10174 (N_10174,N_4296,N_6743);
or U10175 (N_10175,N_5853,N_7155);
nand U10176 (N_10176,N_5031,N_7290);
nand U10177 (N_10177,N_5169,N_4645);
or U10178 (N_10178,N_4370,N_5356);
and U10179 (N_10179,N_5448,N_6727);
nor U10180 (N_10180,N_6021,N_6762);
and U10181 (N_10181,N_7218,N_7949);
nand U10182 (N_10182,N_5635,N_7796);
xor U10183 (N_10183,N_5920,N_4399);
nor U10184 (N_10184,N_7410,N_5486);
or U10185 (N_10185,N_7241,N_5627);
xor U10186 (N_10186,N_4777,N_6914);
xor U10187 (N_10187,N_6079,N_7833);
nor U10188 (N_10188,N_7744,N_6363);
xor U10189 (N_10189,N_4811,N_6916);
and U10190 (N_10190,N_7154,N_4393);
or U10191 (N_10191,N_6385,N_6350);
xor U10192 (N_10192,N_5183,N_6291);
and U10193 (N_10193,N_5515,N_5101);
and U10194 (N_10194,N_7665,N_6967);
or U10195 (N_10195,N_6811,N_4388);
or U10196 (N_10196,N_6348,N_7820);
nor U10197 (N_10197,N_6980,N_5234);
and U10198 (N_10198,N_7918,N_5516);
or U10199 (N_10199,N_6435,N_7437);
nand U10200 (N_10200,N_7436,N_6277);
or U10201 (N_10201,N_7523,N_4722);
nor U10202 (N_10202,N_7214,N_6717);
nor U10203 (N_10203,N_5768,N_6088);
and U10204 (N_10204,N_6339,N_4563);
nor U10205 (N_10205,N_4219,N_6327);
or U10206 (N_10206,N_7004,N_7884);
or U10207 (N_10207,N_5816,N_4173);
nand U10208 (N_10208,N_7412,N_7535);
nand U10209 (N_10209,N_7148,N_7968);
xnor U10210 (N_10210,N_4960,N_4778);
nand U10211 (N_10211,N_4606,N_7657);
nor U10212 (N_10212,N_4102,N_6135);
or U10213 (N_10213,N_6544,N_5226);
nor U10214 (N_10214,N_7204,N_4768);
nand U10215 (N_10215,N_7569,N_7179);
or U10216 (N_10216,N_5326,N_5484);
xnor U10217 (N_10217,N_5434,N_5152);
and U10218 (N_10218,N_7037,N_6960);
nor U10219 (N_10219,N_5465,N_5259);
and U10220 (N_10220,N_5700,N_5122);
nor U10221 (N_10221,N_5173,N_4683);
xor U10222 (N_10222,N_6682,N_6888);
or U10223 (N_10223,N_5867,N_5971);
nand U10224 (N_10224,N_6768,N_5343);
nor U10225 (N_10225,N_6064,N_7444);
nand U10226 (N_10226,N_6231,N_5835);
and U10227 (N_10227,N_7299,N_6040);
and U10228 (N_10228,N_4727,N_7359);
nor U10229 (N_10229,N_6558,N_5389);
and U10230 (N_10230,N_4216,N_4563);
and U10231 (N_10231,N_5420,N_7593);
nor U10232 (N_10232,N_6865,N_7935);
nand U10233 (N_10233,N_4271,N_4064);
and U10234 (N_10234,N_5587,N_4253);
nand U10235 (N_10235,N_7344,N_5813);
nand U10236 (N_10236,N_6704,N_4784);
nand U10237 (N_10237,N_4025,N_6458);
and U10238 (N_10238,N_6872,N_4495);
nor U10239 (N_10239,N_7793,N_4298);
and U10240 (N_10240,N_5607,N_7279);
nand U10241 (N_10241,N_5748,N_4549);
or U10242 (N_10242,N_7328,N_4368);
nand U10243 (N_10243,N_6640,N_5603);
or U10244 (N_10244,N_7705,N_6196);
or U10245 (N_10245,N_7466,N_5359);
or U10246 (N_10246,N_5315,N_5973);
nor U10247 (N_10247,N_6029,N_5741);
nor U10248 (N_10248,N_7497,N_7095);
or U10249 (N_10249,N_5034,N_7081);
or U10250 (N_10250,N_4621,N_6900);
nor U10251 (N_10251,N_7276,N_6454);
or U10252 (N_10252,N_4352,N_4032);
nand U10253 (N_10253,N_7491,N_6697);
or U10254 (N_10254,N_5436,N_4296);
and U10255 (N_10255,N_6641,N_7282);
and U10256 (N_10256,N_4193,N_5853);
and U10257 (N_10257,N_6955,N_4819);
and U10258 (N_10258,N_4845,N_7563);
nand U10259 (N_10259,N_6228,N_6751);
and U10260 (N_10260,N_5061,N_5578);
xnor U10261 (N_10261,N_7592,N_7293);
xor U10262 (N_10262,N_4840,N_4001);
xnor U10263 (N_10263,N_6262,N_4041);
nand U10264 (N_10264,N_5619,N_7077);
xor U10265 (N_10265,N_5435,N_4002);
and U10266 (N_10266,N_6317,N_6586);
and U10267 (N_10267,N_4919,N_5101);
nor U10268 (N_10268,N_6127,N_6148);
and U10269 (N_10269,N_6065,N_7983);
nand U10270 (N_10270,N_4661,N_7754);
or U10271 (N_10271,N_7390,N_5891);
xor U10272 (N_10272,N_7302,N_7202);
nor U10273 (N_10273,N_5504,N_4534);
and U10274 (N_10274,N_4869,N_5990);
or U10275 (N_10275,N_5079,N_5127);
or U10276 (N_10276,N_4085,N_7923);
nor U10277 (N_10277,N_4242,N_4191);
nand U10278 (N_10278,N_4867,N_4574);
or U10279 (N_10279,N_5181,N_5368);
or U10280 (N_10280,N_7272,N_6473);
or U10281 (N_10281,N_5579,N_7454);
nor U10282 (N_10282,N_7554,N_4101);
xnor U10283 (N_10283,N_4493,N_7227);
or U10284 (N_10284,N_6518,N_5535);
nand U10285 (N_10285,N_7704,N_7871);
or U10286 (N_10286,N_4968,N_5934);
xnor U10287 (N_10287,N_7503,N_4764);
nand U10288 (N_10288,N_4038,N_6703);
nor U10289 (N_10289,N_7869,N_5016);
or U10290 (N_10290,N_6460,N_7608);
nor U10291 (N_10291,N_6056,N_4643);
and U10292 (N_10292,N_6995,N_6128);
nor U10293 (N_10293,N_4329,N_4203);
nand U10294 (N_10294,N_6863,N_7152);
or U10295 (N_10295,N_7958,N_6066);
or U10296 (N_10296,N_6331,N_4172);
nand U10297 (N_10297,N_5238,N_6508);
nor U10298 (N_10298,N_4653,N_5010);
and U10299 (N_10299,N_6570,N_4387);
or U10300 (N_10300,N_7746,N_4651);
or U10301 (N_10301,N_7307,N_5545);
and U10302 (N_10302,N_5754,N_6910);
and U10303 (N_10303,N_5510,N_6140);
and U10304 (N_10304,N_4383,N_7431);
and U10305 (N_10305,N_5704,N_4469);
or U10306 (N_10306,N_7308,N_6919);
and U10307 (N_10307,N_5562,N_7103);
nand U10308 (N_10308,N_6009,N_7886);
nand U10309 (N_10309,N_7660,N_5314);
or U10310 (N_10310,N_7625,N_5822);
nor U10311 (N_10311,N_4209,N_6287);
or U10312 (N_10312,N_7216,N_4886);
and U10313 (N_10313,N_4420,N_7342);
or U10314 (N_10314,N_5066,N_5616);
nand U10315 (N_10315,N_6090,N_7365);
nand U10316 (N_10316,N_4004,N_4470);
or U10317 (N_10317,N_7605,N_6118);
nor U10318 (N_10318,N_6712,N_5782);
or U10319 (N_10319,N_5541,N_4573);
nor U10320 (N_10320,N_4922,N_5179);
and U10321 (N_10321,N_4190,N_6781);
or U10322 (N_10322,N_6834,N_4278);
and U10323 (N_10323,N_7337,N_5161);
nand U10324 (N_10324,N_5608,N_5828);
nor U10325 (N_10325,N_4080,N_5533);
nor U10326 (N_10326,N_6325,N_5302);
nor U10327 (N_10327,N_6275,N_4244);
nand U10328 (N_10328,N_6002,N_7675);
xnor U10329 (N_10329,N_6769,N_6114);
nor U10330 (N_10330,N_5947,N_4725);
nor U10331 (N_10331,N_5865,N_6134);
or U10332 (N_10332,N_6093,N_4941);
nor U10333 (N_10333,N_7285,N_7355);
or U10334 (N_10334,N_7786,N_6226);
nand U10335 (N_10335,N_6182,N_6071);
nor U10336 (N_10336,N_4096,N_6783);
nor U10337 (N_10337,N_7594,N_4274);
and U10338 (N_10338,N_6588,N_7096);
nand U10339 (N_10339,N_5326,N_5160);
xor U10340 (N_10340,N_5909,N_7576);
and U10341 (N_10341,N_7992,N_6943);
xor U10342 (N_10342,N_6087,N_4410);
or U10343 (N_10343,N_6664,N_5057);
or U10344 (N_10344,N_6990,N_5663);
and U10345 (N_10345,N_5811,N_4574);
nand U10346 (N_10346,N_5236,N_5214);
nand U10347 (N_10347,N_4409,N_6992);
nand U10348 (N_10348,N_6729,N_6022);
and U10349 (N_10349,N_6335,N_4306);
and U10350 (N_10350,N_5374,N_6530);
nor U10351 (N_10351,N_7530,N_6261);
nand U10352 (N_10352,N_5298,N_7083);
or U10353 (N_10353,N_7177,N_5175);
nor U10354 (N_10354,N_6882,N_4669);
and U10355 (N_10355,N_7056,N_5370);
or U10356 (N_10356,N_7266,N_5551);
nand U10357 (N_10357,N_4854,N_5222);
nand U10358 (N_10358,N_6412,N_6773);
and U10359 (N_10359,N_5574,N_5645);
or U10360 (N_10360,N_4425,N_5811);
or U10361 (N_10361,N_4301,N_7459);
nand U10362 (N_10362,N_7216,N_6597);
nor U10363 (N_10363,N_4370,N_6189);
nand U10364 (N_10364,N_5703,N_4985);
nand U10365 (N_10365,N_6902,N_7481);
nor U10366 (N_10366,N_6842,N_7884);
nand U10367 (N_10367,N_6436,N_6493);
and U10368 (N_10368,N_4806,N_7271);
or U10369 (N_10369,N_7302,N_5903);
xnor U10370 (N_10370,N_7009,N_6937);
or U10371 (N_10371,N_7742,N_4299);
or U10372 (N_10372,N_6081,N_6909);
or U10373 (N_10373,N_7309,N_4148);
and U10374 (N_10374,N_5325,N_5940);
or U10375 (N_10375,N_7668,N_4334);
or U10376 (N_10376,N_4459,N_5731);
and U10377 (N_10377,N_7940,N_5243);
nor U10378 (N_10378,N_6543,N_4160);
nand U10379 (N_10379,N_4805,N_7427);
or U10380 (N_10380,N_6267,N_7796);
xnor U10381 (N_10381,N_6723,N_5413);
nor U10382 (N_10382,N_5539,N_6371);
nand U10383 (N_10383,N_5494,N_4490);
nor U10384 (N_10384,N_6484,N_7367);
or U10385 (N_10385,N_4030,N_4250);
nor U10386 (N_10386,N_5056,N_7774);
nand U10387 (N_10387,N_6469,N_6938);
or U10388 (N_10388,N_6915,N_5989);
nand U10389 (N_10389,N_7101,N_7035);
nor U10390 (N_10390,N_6318,N_7175);
nor U10391 (N_10391,N_4949,N_5684);
nor U10392 (N_10392,N_7813,N_4187);
nand U10393 (N_10393,N_4001,N_7475);
nand U10394 (N_10394,N_7510,N_4222);
nor U10395 (N_10395,N_7865,N_7864);
xor U10396 (N_10396,N_7579,N_6158);
or U10397 (N_10397,N_4006,N_4091);
and U10398 (N_10398,N_4954,N_7373);
nand U10399 (N_10399,N_7159,N_4428);
nand U10400 (N_10400,N_7524,N_7358);
or U10401 (N_10401,N_5764,N_7314);
nand U10402 (N_10402,N_4720,N_7976);
nand U10403 (N_10403,N_4259,N_7686);
xnor U10404 (N_10404,N_7248,N_4860);
nor U10405 (N_10405,N_7904,N_4954);
and U10406 (N_10406,N_6236,N_6946);
or U10407 (N_10407,N_4156,N_5464);
and U10408 (N_10408,N_5096,N_4646);
nand U10409 (N_10409,N_6632,N_4365);
or U10410 (N_10410,N_7104,N_4959);
or U10411 (N_10411,N_4914,N_6681);
and U10412 (N_10412,N_7821,N_6929);
nand U10413 (N_10413,N_7495,N_5762);
nand U10414 (N_10414,N_4958,N_6566);
and U10415 (N_10415,N_5242,N_4497);
xor U10416 (N_10416,N_5163,N_6789);
xnor U10417 (N_10417,N_5578,N_4642);
or U10418 (N_10418,N_5357,N_4836);
nor U10419 (N_10419,N_7504,N_6582);
xor U10420 (N_10420,N_7958,N_4706);
or U10421 (N_10421,N_7062,N_5324);
nor U10422 (N_10422,N_4735,N_6043);
and U10423 (N_10423,N_7514,N_4830);
nand U10424 (N_10424,N_6122,N_5458);
nor U10425 (N_10425,N_5733,N_5669);
nor U10426 (N_10426,N_7011,N_7799);
and U10427 (N_10427,N_6684,N_4555);
nand U10428 (N_10428,N_6659,N_6914);
and U10429 (N_10429,N_4862,N_4189);
nor U10430 (N_10430,N_5903,N_6098);
or U10431 (N_10431,N_6399,N_6781);
xor U10432 (N_10432,N_6491,N_7383);
xnor U10433 (N_10433,N_7047,N_7938);
nor U10434 (N_10434,N_7120,N_4487);
or U10435 (N_10435,N_4534,N_7980);
nor U10436 (N_10436,N_6199,N_6090);
nor U10437 (N_10437,N_7902,N_7799);
nor U10438 (N_10438,N_6370,N_7724);
nand U10439 (N_10439,N_7163,N_5353);
xnor U10440 (N_10440,N_5373,N_7734);
and U10441 (N_10441,N_4578,N_5489);
nand U10442 (N_10442,N_4623,N_6037);
or U10443 (N_10443,N_7535,N_6293);
nor U10444 (N_10444,N_5324,N_7734);
nand U10445 (N_10445,N_6139,N_7895);
nand U10446 (N_10446,N_5046,N_5514);
nand U10447 (N_10447,N_7833,N_6474);
and U10448 (N_10448,N_4958,N_7040);
nor U10449 (N_10449,N_6735,N_6929);
or U10450 (N_10450,N_5831,N_4551);
and U10451 (N_10451,N_5520,N_6475);
nor U10452 (N_10452,N_7054,N_4290);
nor U10453 (N_10453,N_7884,N_5236);
or U10454 (N_10454,N_4522,N_4772);
xnor U10455 (N_10455,N_6272,N_4007);
and U10456 (N_10456,N_5915,N_5973);
nor U10457 (N_10457,N_7210,N_4274);
nor U10458 (N_10458,N_4433,N_7016);
and U10459 (N_10459,N_5222,N_7469);
nor U10460 (N_10460,N_7052,N_4522);
and U10461 (N_10461,N_7015,N_5190);
xor U10462 (N_10462,N_6050,N_4214);
nand U10463 (N_10463,N_5181,N_6113);
and U10464 (N_10464,N_7130,N_5746);
or U10465 (N_10465,N_6970,N_5441);
or U10466 (N_10466,N_7570,N_6920);
nor U10467 (N_10467,N_7374,N_5393);
nand U10468 (N_10468,N_7354,N_7655);
nor U10469 (N_10469,N_7847,N_7430);
xnor U10470 (N_10470,N_5231,N_5193);
nand U10471 (N_10471,N_4124,N_6037);
xor U10472 (N_10472,N_6276,N_5023);
nand U10473 (N_10473,N_6325,N_6435);
nor U10474 (N_10474,N_4168,N_6062);
and U10475 (N_10475,N_7599,N_5831);
and U10476 (N_10476,N_5918,N_7979);
nand U10477 (N_10477,N_7552,N_5937);
and U10478 (N_10478,N_5564,N_6477);
and U10479 (N_10479,N_5015,N_6892);
and U10480 (N_10480,N_6340,N_4463);
or U10481 (N_10481,N_7772,N_6579);
nor U10482 (N_10482,N_7924,N_5482);
or U10483 (N_10483,N_7652,N_4264);
nor U10484 (N_10484,N_4241,N_5204);
nand U10485 (N_10485,N_7693,N_6574);
nor U10486 (N_10486,N_6803,N_5950);
nor U10487 (N_10487,N_6491,N_5896);
or U10488 (N_10488,N_4322,N_7044);
and U10489 (N_10489,N_4765,N_7307);
nor U10490 (N_10490,N_4029,N_5412);
nor U10491 (N_10491,N_6955,N_7911);
or U10492 (N_10492,N_5199,N_6281);
xor U10493 (N_10493,N_4061,N_6884);
and U10494 (N_10494,N_6799,N_7644);
nor U10495 (N_10495,N_4493,N_7444);
and U10496 (N_10496,N_7667,N_7005);
or U10497 (N_10497,N_6985,N_7652);
nor U10498 (N_10498,N_4726,N_7581);
nor U10499 (N_10499,N_7893,N_4659);
and U10500 (N_10500,N_7046,N_4873);
nor U10501 (N_10501,N_5385,N_6669);
nand U10502 (N_10502,N_5543,N_4862);
or U10503 (N_10503,N_4353,N_6491);
nor U10504 (N_10504,N_4840,N_6574);
nor U10505 (N_10505,N_6073,N_7616);
and U10506 (N_10506,N_6350,N_4271);
and U10507 (N_10507,N_5664,N_5770);
nor U10508 (N_10508,N_5625,N_6722);
nand U10509 (N_10509,N_5118,N_7790);
or U10510 (N_10510,N_5851,N_6410);
nand U10511 (N_10511,N_4159,N_7615);
and U10512 (N_10512,N_4638,N_5138);
or U10513 (N_10513,N_4222,N_6984);
and U10514 (N_10514,N_5771,N_7978);
nand U10515 (N_10515,N_7822,N_5691);
nand U10516 (N_10516,N_6625,N_4578);
nor U10517 (N_10517,N_4437,N_4887);
nand U10518 (N_10518,N_7599,N_6921);
or U10519 (N_10519,N_5420,N_6598);
or U10520 (N_10520,N_6696,N_5836);
and U10521 (N_10521,N_7168,N_4558);
and U10522 (N_10522,N_6727,N_4642);
nand U10523 (N_10523,N_7367,N_7337);
or U10524 (N_10524,N_4608,N_4336);
nand U10525 (N_10525,N_6100,N_6503);
nor U10526 (N_10526,N_7228,N_7631);
nand U10527 (N_10527,N_6212,N_5149);
nand U10528 (N_10528,N_4051,N_6777);
nor U10529 (N_10529,N_6328,N_6786);
and U10530 (N_10530,N_5751,N_5320);
nor U10531 (N_10531,N_5636,N_7351);
xnor U10532 (N_10532,N_7537,N_5682);
nor U10533 (N_10533,N_6255,N_7267);
nand U10534 (N_10534,N_4207,N_6239);
and U10535 (N_10535,N_4414,N_4272);
nand U10536 (N_10536,N_7702,N_4431);
or U10537 (N_10537,N_6808,N_4232);
or U10538 (N_10538,N_6469,N_4988);
nor U10539 (N_10539,N_5671,N_7393);
nor U10540 (N_10540,N_6016,N_7295);
and U10541 (N_10541,N_4126,N_7256);
or U10542 (N_10542,N_6299,N_4511);
or U10543 (N_10543,N_6733,N_5580);
nand U10544 (N_10544,N_7344,N_7316);
nor U10545 (N_10545,N_4348,N_6133);
or U10546 (N_10546,N_6070,N_7483);
or U10547 (N_10547,N_7368,N_7906);
or U10548 (N_10548,N_5781,N_4044);
nand U10549 (N_10549,N_6052,N_4454);
nand U10550 (N_10550,N_6882,N_6078);
nor U10551 (N_10551,N_6223,N_4122);
or U10552 (N_10552,N_5786,N_7475);
nand U10553 (N_10553,N_5017,N_4413);
nand U10554 (N_10554,N_4093,N_5927);
and U10555 (N_10555,N_5141,N_7578);
nor U10556 (N_10556,N_7815,N_4741);
or U10557 (N_10557,N_5724,N_5021);
and U10558 (N_10558,N_6156,N_5558);
nor U10559 (N_10559,N_5446,N_7432);
nand U10560 (N_10560,N_6853,N_4270);
or U10561 (N_10561,N_5448,N_4976);
or U10562 (N_10562,N_7584,N_7138);
nand U10563 (N_10563,N_6573,N_4475);
nand U10564 (N_10564,N_6702,N_6392);
xnor U10565 (N_10565,N_7918,N_6848);
nand U10566 (N_10566,N_7251,N_6748);
nand U10567 (N_10567,N_7638,N_6657);
and U10568 (N_10568,N_4265,N_7002);
and U10569 (N_10569,N_6090,N_4957);
and U10570 (N_10570,N_5676,N_5747);
xor U10571 (N_10571,N_4119,N_4984);
and U10572 (N_10572,N_4349,N_5431);
or U10573 (N_10573,N_4494,N_6910);
nand U10574 (N_10574,N_5567,N_6288);
nor U10575 (N_10575,N_5889,N_5578);
or U10576 (N_10576,N_5092,N_6367);
and U10577 (N_10577,N_6655,N_6834);
or U10578 (N_10578,N_6929,N_6320);
nand U10579 (N_10579,N_7991,N_4313);
xor U10580 (N_10580,N_6327,N_7945);
nand U10581 (N_10581,N_4199,N_4036);
and U10582 (N_10582,N_4683,N_6432);
nand U10583 (N_10583,N_7543,N_4619);
or U10584 (N_10584,N_6888,N_4963);
and U10585 (N_10585,N_7636,N_4807);
or U10586 (N_10586,N_7145,N_4729);
nand U10587 (N_10587,N_6068,N_5263);
or U10588 (N_10588,N_4398,N_7109);
nand U10589 (N_10589,N_6506,N_5013);
and U10590 (N_10590,N_4530,N_4050);
or U10591 (N_10591,N_4432,N_5224);
or U10592 (N_10592,N_6460,N_7120);
nand U10593 (N_10593,N_6277,N_6856);
and U10594 (N_10594,N_5319,N_7003);
nand U10595 (N_10595,N_4670,N_5059);
nand U10596 (N_10596,N_4815,N_5207);
and U10597 (N_10597,N_4459,N_6387);
or U10598 (N_10598,N_4833,N_4069);
nor U10599 (N_10599,N_6830,N_5859);
nor U10600 (N_10600,N_7128,N_4364);
nor U10601 (N_10601,N_7344,N_6747);
or U10602 (N_10602,N_4499,N_7009);
or U10603 (N_10603,N_7497,N_4703);
nand U10604 (N_10604,N_7133,N_7983);
nand U10605 (N_10605,N_5306,N_4123);
xor U10606 (N_10606,N_7262,N_4621);
or U10607 (N_10607,N_6661,N_4178);
or U10608 (N_10608,N_6122,N_5033);
or U10609 (N_10609,N_7302,N_7183);
xnor U10610 (N_10610,N_7349,N_6536);
nor U10611 (N_10611,N_7307,N_7239);
xor U10612 (N_10612,N_5847,N_4124);
and U10613 (N_10613,N_6232,N_4773);
nand U10614 (N_10614,N_7400,N_7908);
nor U10615 (N_10615,N_6745,N_6314);
nor U10616 (N_10616,N_7972,N_6633);
nand U10617 (N_10617,N_6804,N_4359);
nor U10618 (N_10618,N_5257,N_6924);
or U10619 (N_10619,N_5382,N_4814);
and U10620 (N_10620,N_7436,N_4088);
nor U10621 (N_10621,N_5752,N_5022);
and U10622 (N_10622,N_4965,N_4207);
or U10623 (N_10623,N_5827,N_6005);
xor U10624 (N_10624,N_6956,N_4481);
or U10625 (N_10625,N_4861,N_4722);
or U10626 (N_10626,N_6719,N_6499);
or U10627 (N_10627,N_4989,N_5966);
nor U10628 (N_10628,N_5352,N_6888);
nor U10629 (N_10629,N_5056,N_5287);
nor U10630 (N_10630,N_5772,N_7796);
and U10631 (N_10631,N_7653,N_6950);
nand U10632 (N_10632,N_7950,N_5724);
nor U10633 (N_10633,N_5318,N_6741);
or U10634 (N_10634,N_7806,N_4998);
and U10635 (N_10635,N_6346,N_4411);
and U10636 (N_10636,N_7543,N_7805);
xor U10637 (N_10637,N_6165,N_6211);
and U10638 (N_10638,N_4031,N_5384);
nor U10639 (N_10639,N_7007,N_6108);
and U10640 (N_10640,N_5532,N_6369);
or U10641 (N_10641,N_5385,N_7559);
and U10642 (N_10642,N_4001,N_6191);
and U10643 (N_10643,N_6846,N_5348);
or U10644 (N_10644,N_7298,N_7555);
nor U10645 (N_10645,N_7179,N_6599);
nand U10646 (N_10646,N_4112,N_5910);
and U10647 (N_10647,N_7558,N_4359);
nor U10648 (N_10648,N_5246,N_4190);
nand U10649 (N_10649,N_4757,N_7179);
nand U10650 (N_10650,N_6540,N_4018);
or U10651 (N_10651,N_7818,N_4177);
and U10652 (N_10652,N_4727,N_7652);
and U10653 (N_10653,N_4040,N_5328);
or U10654 (N_10654,N_5665,N_5367);
nor U10655 (N_10655,N_6630,N_7166);
nor U10656 (N_10656,N_6035,N_5704);
and U10657 (N_10657,N_5529,N_5535);
or U10658 (N_10658,N_7913,N_5893);
nor U10659 (N_10659,N_6041,N_4293);
xor U10660 (N_10660,N_6643,N_6186);
or U10661 (N_10661,N_5539,N_6042);
or U10662 (N_10662,N_4419,N_4693);
or U10663 (N_10663,N_6894,N_7328);
or U10664 (N_10664,N_7171,N_6469);
nand U10665 (N_10665,N_6943,N_4267);
and U10666 (N_10666,N_6449,N_7851);
nor U10667 (N_10667,N_5006,N_6911);
and U10668 (N_10668,N_4888,N_4894);
nand U10669 (N_10669,N_7135,N_6352);
nor U10670 (N_10670,N_7426,N_6140);
nand U10671 (N_10671,N_4904,N_4812);
nor U10672 (N_10672,N_4551,N_6136);
nor U10673 (N_10673,N_7337,N_6945);
or U10674 (N_10674,N_6895,N_7799);
and U10675 (N_10675,N_4527,N_5559);
and U10676 (N_10676,N_6756,N_7306);
or U10677 (N_10677,N_6327,N_6801);
nand U10678 (N_10678,N_4096,N_5005);
xor U10679 (N_10679,N_5176,N_6254);
and U10680 (N_10680,N_5271,N_4477);
and U10681 (N_10681,N_5023,N_4900);
nor U10682 (N_10682,N_6558,N_4742);
nand U10683 (N_10683,N_7248,N_7156);
or U10684 (N_10684,N_4069,N_7869);
or U10685 (N_10685,N_6087,N_6697);
and U10686 (N_10686,N_4713,N_7826);
or U10687 (N_10687,N_6782,N_5856);
and U10688 (N_10688,N_6381,N_7161);
and U10689 (N_10689,N_5235,N_5154);
or U10690 (N_10690,N_7475,N_7449);
and U10691 (N_10691,N_7428,N_4890);
nand U10692 (N_10692,N_7182,N_6232);
nor U10693 (N_10693,N_5227,N_5361);
nand U10694 (N_10694,N_6360,N_6544);
nand U10695 (N_10695,N_7278,N_7408);
and U10696 (N_10696,N_6717,N_6512);
nor U10697 (N_10697,N_6336,N_5518);
or U10698 (N_10698,N_5372,N_5977);
nor U10699 (N_10699,N_5341,N_5491);
nor U10700 (N_10700,N_7793,N_4444);
nand U10701 (N_10701,N_5822,N_7267);
and U10702 (N_10702,N_6831,N_5901);
and U10703 (N_10703,N_7608,N_5600);
nor U10704 (N_10704,N_7886,N_4142);
or U10705 (N_10705,N_5990,N_6032);
or U10706 (N_10706,N_6926,N_4893);
nor U10707 (N_10707,N_6068,N_6430);
nor U10708 (N_10708,N_6001,N_6629);
and U10709 (N_10709,N_6934,N_6889);
nor U10710 (N_10710,N_5061,N_6753);
and U10711 (N_10711,N_4610,N_4295);
nor U10712 (N_10712,N_7724,N_4740);
xnor U10713 (N_10713,N_5753,N_4386);
xnor U10714 (N_10714,N_6588,N_7927);
or U10715 (N_10715,N_4783,N_5621);
or U10716 (N_10716,N_5098,N_7216);
nor U10717 (N_10717,N_4239,N_4019);
and U10718 (N_10718,N_7297,N_4432);
and U10719 (N_10719,N_5317,N_5683);
nand U10720 (N_10720,N_4372,N_7383);
nand U10721 (N_10721,N_7985,N_5673);
and U10722 (N_10722,N_4168,N_5975);
and U10723 (N_10723,N_6973,N_7673);
and U10724 (N_10724,N_7793,N_6715);
nand U10725 (N_10725,N_4761,N_7957);
nand U10726 (N_10726,N_6014,N_4920);
nor U10727 (N_10727,N_4628,N_7028);
xnor U10728 (N_10728,N_7266,N_6913);
or U10729 (N_10729,N_7288,N_7357);
nor U10730 (N_10730,N_6935,N_7716);
nand U10731 (N_10731,N_7215,N_5543);
xor U10732 (N_10732,N_7761,N_5483);
or U10733 (N_10733,N_6525,N_5713);
and U10734 (N_10734,N_6266,N_7127);
and U10735 (N_10735,N_5916,N_4671);
nand U10736 (N_10736,N_6077,N_6102);
nor U10737 (N_10737,N_6234,N_5252);
nand U10738 (N_10738,N_7566,N_6908);
or U10739 (N_10739,N_7393,N_5022);
nor U10740 (N_10740,N_5414,N_4647);
nand U10741 (N_10741,N_7510,N_5222);
nor U10742 (N_10742,N_7788,N_6319);
nor U10743 (N_10743,N_7806,N_4656);
and U10744 (N_10744,N_7552,N_6256);
nor U10745 (N_10745,N_4465,N_6208);
and U10746 (N_10746,N_4623,N_5838);
nand U10747 (N_10747,N_6004,N_4895);
xnor U10748 (N_10748,N_4228,N_6631);
or U10749 (N_10749,N_4790,N_7436);
nand U10750 (N_10750,N_4936,N_4409);
or U10751 (N_10751,N_4137,N_6556);
xnor U10752 (N_10752,N_6019,N_4373);
nand U10753 (N_10753,N_6067,N_7944);
nor U10754 (N_10754,N_6997,N_6122);
nand U10755 (N_10755,N_6814,N_5524);
nand U10756 (N_10756,N_5464,N_6859);
and U10757 (N_10757,N_7532,N_6132);
and U10758 (N_10758,N_5236,N_4764);
and U10759 (N_10759,N_4492,N_7899);
nor U10760 (N_10760,N_4085,N_4293);
and U10761 (N_10761,N_4306,N_6441);
nor U10762 (N_10762,N_7837,N_6989);
nor U10763 (N_10763,N_7583,N_6816);
or U10764 (N_10764,N_6118,N_6667);
or U10765 (N_10765,N_7330,N_7711);
or U10766 (N_10766,N_7771,N_5486);
and U10767 (N_10767,N_4561,N_5971);
xor U10768 (N_10768,N_7664,N_6119);
and U10769 (N_10769,N_4845,N_7911);
and U10770 (N_10770,N_6861,N_4541);
or U10771 (N_10771,N_4407,N_5922);
or U10772 (N_10772,N_6331,N_7493);
and U10773 (N_10773,N_7669,N_7287);
and U10774 (N_10774,N_6496,N_6008);
or U10775 (N_10775,N_4589,N_4208);
nand U10776 (N_10776,N_4645,N_5370);
nor U10777 (N_10777,N_5057,N_5522);
xor U10778 (N_10778,N_4940,N_7404);
nor U10779 (N_10779,N_5890,N_7280);
nor U10780 (N_10780,N_7867,N_4864);
nor U10781 (N_10781,N_5654,N_6745);
xor U10782 (N_10782,N_7523,N_6943);
nand U10783 (N_10783,N_6054,N_4138);
nor U10784 (N_10784,N_6012,N_6465);
nor U10785 (N_10785,N_5164,N_4956);
nor U10786 (N_10786,N_5450,N_4048);
nor U10787 (N_10787,N_6372,N_7965);
and U10788 (N_10788,N_5784,N_5448);
or U10789 (N_10789,N_6771,N_7776);
nor U10790 (N_10790,N_7933,N_7237);
or U10791 (N_10791,N_6659,N_7830);
or U10792 (N_10792,N_6667,N_5910);
nand U10793 (N_10793,N_4286,N_4774);
nand U10794 (N_10794,N_4583,N_4554);
or U10795 (N_10795,N_4001,N_5038);
nand U10796 (N_10796,N_7571,N_6082);
or U10797 (N_10797,N_4966,N_4090);
xnor U10798 (N_10798,N_5579,N_6615);
nand U10799 (N_10799,N_5861,N_5965);
nor U10800 (N_10800,N_4615,N_4160);
or U10801 (N_10801,N_6915,N_4295);
and U10802 (N_10802,N_6392,N_5831);
or U10803 (N_10803,N_5194,N_5410);
xnor U10804 (N_10804,N_6855,N_4817);
and U10805 (N_10805,N_4060,N_7695);
nor U10806 (N_10806,N_6630,N_5610);
nor U10807 (N_10807,N_7058,N_7674);
or U10808 (N_10808,N_4174,N_6932);
nor U10809 (N_10809,N_4390,N_7834);
xor U10810 (N_10810,N_6579,N_4912);
nor U10811 (N_10811,N_5838,N_6383);
and U10812 (N_10812,N_6481,N_5571);
nor U10813 (N_10813,N_5016,N_4066);
nand U10814 (N_10814,N_7681,N_5721);
nand U10815 (N_10815,N_6914,N_4524);
xor U10816 (N_10816,N_7003,N_5991);
nor U10817 (N_10817,N_4089,N_6464);
nand U10818 (N_10818,N_6208,N_5407);
nor U10819 (N_10819,N_7554,N_4466);
xor U10820 (N_10820,N_6270,N_7200);
and U10821 (N_10821,N_4685,N_5820);
or U10822 (N_10822,N_6244,N_7401);
and U10823 (N_10823,N_5168,N_6258);
nand U10824 (N_10824,N_6700,N_7135);
nand U10825 (N_10825,N_6310,N_7158);
nand U10826 (N_10826,N_7173,N_4314);
nand U10827 (N_10827,N_7623,N_6819);
xor U10828 (N_10828,N_7578,N_5118);
nor U10829 (N_10829,N_4868,N_6591);
nand U10830 (N_10830,N_4039,N_7669);
nand U10831 (N_10831,N_4243,N_6723);
and U10832 (N_10832,N_4560,N_7326);
nand U10833 (N_10833,N_7602,N_7560);
nor U10834 (N_10834,N_7983,N_6923);
nand U10835 (N_10835,N_7069,N_6460);
and U10836 (N_10836,N_7549,N_4452);
nor U10837 (N_10837,N_7595,N_7888);
nor U10838 (N_10838,N_6287,N_6355);
xor U10839 (N_10839,N_5892,N_7513);
xor U10840 (N_10840,N_6454,N_4535);
xor U10841 (N_10841,N_4273,N_6322);
nand U10842 (N_10842,N_7707,N_6880);
or U10843 (N_10843,N_4199,N_5788);
or U10844 (N_10844,N_7797,N_6242);
nand U10845 (N_10845,N_4685,N_4066);
and U10846 (N_10846,N_7530,N_5449);
nor U10847 (N_10847,N_6378,N_4961);
or U10848 (N_10848,N_6398,N_5527);
or U10849 (N_10849,N_4593,N_4577);
nand U10850 (N_10850,N_5025,N_5442);
or U10851 (N_10851,N_6698,N_4414);
and U10852 (N_10852,N_6542,N_4030);
xor U10853 (N_10853,N_5032,N_6329);
nor U10854 (N_10854,N_6293,N_7263);
nor U10855 (N_10855,N_4940,N_7406);
nand U10856 (N_10856,N_7345,N_6203);
nor U10857 (N_10857,N_5251,N_5229);
xnor U10858 (N_10858,N_5131,N_7959);
and U10859 (N_10859,N_7967,N_4385);
nand U10860 (N_10860,N_5704,N_7014);
xnor U10861 (N_10861,N_7392,N_5417);
nor U10862 (N_10862,N_5850,N_7441);
nand U10863 (N_10863,N_7160,N_7642);
and U10864 (N_10864,N_7708,N_6309);
nand U10865 (N_10865,N_4602,N_7862);
nor U10866 (N_10866,N_7262,N_7188);
or U10867 (N_10867,N_5656,N_7373);
nand U10868 (N_10868,N_5244,N_6889);
nand U10869 (N_10869,N_4674,N_5443);
or U10870 (N_10870,N_6155,N_5435);
and U10871 (N_10871,N_6590,N_6885);
and U10872 (N_10872,N_6653,N_4430);
or U10873 (N_10873,N_5339,N_4845);
nand U10874 (N_10874,N_4836,N_4383);
xor U10875 (N_10875,N_4123,N_6317);
and U10876 (N_10876,N_4725,N_7606);
and U10877 (N_10877,N_7680,N_5445);
and U10878 (N_10878,N_4465,N_7107);
nor U10879 (N_10879,N_4869,N_7863);
or U10880 (N_10880,N_4440,N_7580);
nor U10881 (N_10881,N_7208,N_7149);
nand U10882 (N_10882,N_4457,N_6370);
or U10883 (N_10883,N_6596,N_6889);
nand U10884 (N_10884,N_4620,N_6899);
nand U10885 (N_10885,N_5430,N_6295);
or U10886 (N_10886,N_7615,N_4794);
nand U10887 (N_10887,N_6583,N_5205);
nand U10888 (N_10888,N_6596,N_4334);
nand U10889 (N_10889,N_6697,N_5763);
xnor U10890 (N_10890,N_5469,N_7480);
nor U10891 (N_10891,N_6829,N_5933);
and U10892 (N_10892,N_4852,N_4950);
nand U10893 (N_10893,N_4955,N_7938);
or U10894 (N_10894,N_7624,N_7076);
nand U10895 (N_10895,N_4201,N_7629);
and U10896 (N_10896,N_4258,N_5064);
and U10897 (N_10897,N_4634,N_4660);
nand U10898 (N_10898,N_7617,N_6594);
and U10899 (N_10899,N_5502,N_5623);
nand U10900 (N_10900,N_5373,N_7883);
and U10901 (N_10901,N_5342,N_4832);
nand U10902 (N_10902,N_7227,N_6743);
and U10903 (N_10903,N_5251,N_6498);
and U10904 (N_10904,N_5009,N_6863);
and U10905 (N_10905,N_5354,N_6566);
and U10906 (N_10906,N_4623,N_4328);
nand U10907 (N_10907,N_7380,N_7862);
or U10908 (N_10908,N_5205,N_7480);
nand U10909 (N_10909,N_6243,N_6042);
nand U10910 (N_10910,N_5096,N_6328);
nand U10911 (N_10911,N_5959,N_4272);
or U10912 (N_10912,N_4947,N_5202);
nor U10913 (N_10913,N_4020,N_4885);
and U10914 (N_10914,N_5944,N_4720);
or U10915 (N_10915,N_6983,N_6550);
xor U10916 (N_10916,N_6190,N_4494);
or U10917 (N_10917,N_6782,N_7064);
xor U10918 (N_10918,N_7742,N_7182);
nor U10919 (N_10919,N_4525,N_7640);
nor U10920 (N_10920,N_5138,N_4125);
nand U10921 (N_10921,N_5019,N_7941);
nand U10922 (N_10922,N_4084,N_6306);
and U10923 (N_10923,N_4377,N_7907);
nand U10924 (N_10924,N_7190,N_6317);
nand U10925 (N_10925,N_6899,N_6403);
and U10926 (N_10926,N_7699,N_6871);
or U10927 (N_10927,N_6978,N_5718);
nand U10928 (N_10928,N_4543,N_5455);
nor U10929 (N_10929,N_5251,N_7161);
or U10930 (N_10930,N_5546,N_4250);
nor U10931 (N_10931,N_6239,N_4430);
or U10932 (N_10932,N_7519,N_4005);
or U10933 (N_10933,N_4805,N_4206);
nand U10934 (N_10934,N_5117,N_6087);
xnor U10935 (N_10935,N_6071,N_7964);
and U10936 (N_10936,N_5938,N_5137);
or U10937 (N_10937,N_7569,N_4322);
or U10938 (N_10938,N_7151,N_5181);
or U10939 (N_10939,N_4093,N_7403);
nor U10940 (N_10940,N_7469,N_4414);
or U10941 (N_10941,N_5026,N_5100);
nand U10942 (N_10942,N_4067,N_7697);
nor U10943 (N_10943,N_4715,N_5145);
nor U10944 (N_10944,N_6228,N_4533);
xnor U10945 (N_10945,N_4829,N_7029);
nand U10946 (N_10946,N_5584,N_7600);
and U10947 (N_10947,N_5914,N_6119);
nor U10948 (N_10948,N_4425,N_7293);
xnor U10949 (N_10949,N_5643,N_5352);
nand U10950 (N_10950,N_4173,N_5051);
nand U10951 (N_10951,N_6516,N_4279);
nand U10952 (N_10952,N_5296,N_7245);
nor U10953 (N_10953,N_4636,N_7523);
and U10954 (N_10954,N_5916,N_7180);
xor U10955 (N_10955,N_5400,N_5601);
xor U10956 (N_10956,N_6563,N_4243);
or U10957 (N_10957,N_4399,N_4971);
and U10958 (N_10958,N_4726,N_5947);
and U10959 (N_10959,N_6630,N_5649);
nor U10960 (N_10960,N_6318,N_7621);
nor U10961 (N_10961,N_5726,N_7327);
nor U10962 (N_10962,N_5697,N_5080);
and U10963 (N_10963,N_5864,N_5268);
nand U10964 (N_10964,N_7244,N_7781);
nand U10965 (N_10965,N_5124,N_7060);
or U10966 (N_10966,N_4620,N_6855);
nor U10967 (N_10967,N_4047,N_6803);
or U10968 (N_10968,N_6931,N_5295);
or U10969 (N_10969,N_6729,N_7301);
or U10970 (N_10970,N_4641,N_4385);
nand U10971 (N_10971,N_7798,N_5262);
nand U10972 (N_10972,N_4861,N_7533);
nand U10973 (N_10973,N_4323,N_6126);
and U10974 (N_10974,N_4992,N_5381);
and U10975 (N_10975,N_7896,N_4375);
and U10976 (N_10976,N_5675,N_4925);
nand U10977 (N_10977,N_7639,N_5212);
and U10978 (N_10978,N_4547,N_6747);
or U10979 (N_10979,N_7378,N_6598);
nand U10980 (N_10980,N_4153,N_7293);
nand U10981 (N_10981,N_4339,N_5108);
or U10982 (N_10982,N_5520,N_6202);
and U10983 (N_10983,N_5590,N_5230);
or U10984 (N_10984,N_6272,N_7786);
or U10985 (N_10985,N_4780,N_7254);
nand U10986 (N_10986,N_7341,N_7232);
xor U10987 (N_10987,N_5007,N_6873);
nand U10988 (N_10988,N_7248,N_5378);
nand U10989 (N_10989,N_7134,N_6140);
xor U10990 (N_10990,N_6553,N_5013);
nand U10991 (N_10991,N_4354,N_6295);
or U10992 (N_10992,N_5794,N_4946);
nor U10993 (N_10993,N_7914,N_7840);
xor U10994 (N_10994,N_4669,N_7484);
or U10995 (N_10995,N_5726,N_6003);
nor U10996 (N_10996,N_7232,N_6549);
and U10997 (N_10997,N_5052,N_6427);
nand U10998 (N_10998,N_6823,N_4836);
or U10999 (N_10999,N_6905,N_7253);
xnor U11000 (N_11000,N_5269,N_4484);
or U11001 (N_11001,N_4582,N_6965);
nand U11002 (N_11002,N_6303,N_6846);
nand U11003 (N_11003,N_5603,N_6677);
nor U11004 (N_11004,N_4660,N_6271);
or U11005 (N_11005,N_4361,N_4808);
nor U11006 (N_11006,N_6197,N_6771);
or U11007 (N_11007,N_7721,N_7457);
nand U11008 (N_11008,N_4468,N_7058);
nand U11009 (N_11009,N_5545,N_5072);
and U11010 (N_11010,N_4767,N_4348);
nor U11011 (N_11011,N_5723,N_5921);
nor U11012 (N_11012,N_6659,N_7151);
or U11013 (N_11013,N_4898,N_5612);
nor U11014 (N_11014,N_5759,N_4575);
nand U11015 (N_11015,N_6228,N_7568);
or U11016 (N_11016,N_4024,N_5657);
nor U11017 (N_11017,N_6184,N_7524);
and U11018 (N_11018,N_7279,N_6333);
nand U11019 (N_11019,N_7242,N_7383);
and U11020 (N_11020,N_4833,N_6716);
or U11021 (N_11021,N_5834,N_6876);
and U11022 (N_11022,N_4307,N_6503);
nand U11023 (N_11023,N_6836,N_4515);
and U11024 (N_11024,N_7300,N_6094);
or U11025 (N_11025,N_5379,N_4398);
and U11026 (N_11026,N_4276,N_4181);
xor U11027 (N_11027,N_5388,N_6635);
nand U11028 (N_11028,N_6826,N_7584);
or U11029 (N_11029,N_5551,N_5235);
xnor U11030 (N_11030,N_7586,N_4711);
and U11031 (N_11031,N_5350,N_6946);
nor U11032 (N_11032,N_7843,N_6182);
nand U11033 (N_11033,N_4008,N_4187);
or U11034 (N_11034,N_7154,N_4789);
nand U11035 (N_11035,N_6569,N_5104);
and U11036 (N_11036,N_7887,N_6432);
and U11037 (N_11037,N_5764,N_7951);
nand U11038 (N_11038,N_4506,N_7943);
and U11039 (N_11039,N_6532,N_5181);
nand U11040 (N_11040,N_5084,N_5068);
or U11041 (N_11041,N_4318,N_4989);
nand U11042 (N_11042,N_5147,N_5902);
nor U11043 (N_11043,N_7589,N_7273);
or U11044 (N_11044,N_5071,N_4995);
xnor U11045 (N_11045,N_4914,N_6248);
nor U11046 (N_11046,N_4580,N_7846);
and U11047 (N_11047,N_7649,N_6870);
nand U11048 (N_11048,N_5238,N_5897);
nand U11049 (N_11049,N_6251,N_6816);
nand U11050 (N_11050,N_7584,N_7255);
xor U11051 (N_11051,N_6552,N_6533);
or U11052 (N_11052,N_6612,N_5076);
and U11053 (N_11053,N_7334,N_6334);
or U11054 (N_11054,N_6873,N_7596);
and U11055 (N_11055,N_7433,N_5586);
nand U11056 (N_11056,N_6451,N_4884);
nor U11057 (N_11057,N_5635,N_5289);
nand U11058 (N_11058,N_6738,N_4865);
nor U11059 (N_11059,N_7062,N_7616);
and U11060 (N_11060,N_5166,N_4919);
and U11061 (N_11061,N_4943,N_7241);
and U11062 (N_11062,N_4967,N_7384);
and U11063 (N_11063,N_6591,N_5843);
or U11064 (N_11064,N_7118,N_7672);
nor U11065 (N_11065,N_6127,N_4167);
or U11066 (N_11066,N_6636,N_7161);
or U11067 (N_11067,N_5737,N_5202);
nor U11068 (N_11068,N_5992,N_7319);
and U11069 (N_11069,N_6281,N_5706);
nand U11070 (N_11070,N_4184,N_5086);
xor U11071 (N_11071,N_6768,N_7534);
xor U11072 (N_11072,N_4763,N_6427);
and U11073 (N_11073,N_5676,N_7771);
nor U11074 (N_11074,N_4091,N_6229);
nor U11075 (N_11075,N_6628,N_7099);
nor U11076 (N_11076,N_7845,N_7722);
or U11077 (N_11077,N_7675,N_5147);
or U11078 (N_11078,N_5635,N_4497);
or U11079 (N_11079,N_7766,N_5258);
or U11080 (N_11080,N_6728,N_6244);
nor U11081 (N_11081,N_4197,N_7965);
nand U11082 (N_11082,N_7015,N_4043);
or U11083 (N_11083,N_4685,N_4547);
nand U11084 (N_11084,N_5232,N_6377);
nand U11085 (N_11085,N_7669,N_4318);
nand U11086 (N_11086,N_5258,N_4425);
nand U11087 (N_11087,N_4362,N_6185);
xnor U11088 (N_11088,N_7352,N_4708);
and U11089 (N_11089,N_6091,N_5996);
or U11090 (N_11090,N_5754,N_7924);
nor U11091 (N_11091,N_4011,N_7118);
and U11092 (N_11092,N_7109,N_4298);
or U11093 (N_11093,N_7900,N_4944);
nand U11094 (N_11094,N_7891,N_5054);
or U11095 (N_11095,N_6204,N_4519);
or U11096 (N_11096,N_7695,N_5046);
xnor U11097 (N_11097,N_5159,N_7680);
and U11098 (N_11098,N_4159,N_6689);
or U11099 (N_11099,N_4431,N_4913);
nor U11100 (N_11100,N_6689,N_5450);
nor U11101 (N_11101,N_7948,N_7210);
and U11102 (N_11102,N_7199,N_6959);
and U11103 (N_11103,N_6563,N_6999);
or U11104 (N_11104,N_5062,N_6369);
or U11105 (N_11105,N_4734,N_4587);
nand U11106 (N_11106,N_4032,N_7105);
and U11107 (N_11107,N_4419,N_5774);
and U11108 (N_11108,N_5124,N_5744);
nor U11109 (N_11109,N_6981,N_6724);
nand U11110 (N_11110,N_4392,N_6914);
and U11111 (N_11111,N_4149,N_5328);
nand U11112 (N_11112,N_7739,N_7150);
nor U11113 (N_11113,N_5600,N_6129);
nand U11114 (N_11114,N_4739,N_4709);
nor U11115 (N_11115,N_5121,N_7205);
nand U11116 (N_11116,N_5779,N_5346);
or U11117 (N_11117,N_5730,N_5168);
nor U11118 (N_11118,N_5792,N_6064);
nor U11119 (N_11119,N_6293,N_5215);
nor U11120 (N_11120,N_4926,N_5408);
nand U11121 (N_11121,N_5446,N_5228);
nor U11122 (N_11122,N_5452,N_7181);
nor U11123 (N_11123,N_5461,N_5914);
and U11124 (N_11124,N_4974,N_7184);
xor U11125 (N_11125,N_7909,N_6509);
and U11126 (N_11126,N_7726,N_4996);
xnor U11127 (N_11127,N_7106,N_6975);
nor U11128 (N_11128,N_5826,N_7264);
nand U11129 (N_11129,N_7966,N_7783);
xnor U11130 (N_11130,N_5940,N_5538);
nand U11131 (N_11131,N_5268,N_5595);
and U11132 (N_11132,N_6960,N_7348);
nand U11133 (N_11133,N_6581,N_4284);
or U11134 (N_11134,N_6966,N_4829);
xor U11135 (N_11135,N_4667,N_7100);
or U11136 (N_11136,N_5994,N_7088);
nand U11137 (N_11137,N_4639,N_6106);
nand U11138 (N_11138,N_6004,N_7348);
and U11139 (N_11139,N_5827,N_5698);
nand U11140 (N_11140,N_7850,N_6796);
and U11141 (N_11141,N_6000,N_6832);
and U11142 (N_11142,N_6935,N_4180);
or U11143 (N_11143,N_7196,N_6870);
or U11144 (N_11144,N_6229,N_4238);
and U11145 (N_11145,N_6183,N_4223);
nor U11146 (N_11146,N_5594,N_7109);
and U11147 (N_11147,N_6629,N_7234);
xor U11148 (N_11148,N_6114,N_6065);
and U11149 (N_11149,N_5949,N_5745);
or U11150 (N_11150,N_5805,N_4970);
and U11151 (N_11151,N_7192,N_4561);
nor U11152 (N_11152,N_5320,N_7994);
or U11153 (N_11153,N_5785,N_6212);
and U11154 (N_11154,N_5621,N_6274);
nor U11155 (N_11155,N_6488,N_6595);
or U11156 (N_11156,N_7329,N_7249);
nand U11157 (N_11157,N_6594,N_4635);
or U11158 (N_11158,N_6231,N_6893);
nand U11159 (N_11159,N_6316,N_7344);
nor U11160 (N_11160,N_7744,N_4267);
and U11161 (N_11161,N_5531,N_4579);
or U11162 (N_11162,N_5961,N_7285);
nand U11163 (N_11163,N_6579,N_5742);
and U11164 (N_11164,N_7813,N_5206);
nand U11165 (N_11165,N_6322,N_7666);
nor U11166 (N_11166,N_7731,N_7460);
nand U11167 (N_11167,N_4594,N_7393);
and U11168 (N_11168,N_4624,N_4086);
and U11169 (N_11169,N_6236,N_6752);
or U11170 (N_11170,N_7828,N_6892);
nor U11171 (N_11171,N_6506,N_4414);
nand U11172 (N_11172,N_7036,N_5972);
xor U11173 (N_11173,N_5550,N_4721);
and U11174 (N_11174,N_5644,N_7531);
and U11175 (N_11175,N_4871,N_7103);
or U11176 (N_11176,N_4112,N_6794);
nor U11177 (N_11177,N_6147,N_6132);
xor U11178 (N_11178,N_5755,N_4762);
nor U11179 (N_11179,N_6437,N_7000);
nand U11180 (N_11180,N_6249,N_7201);
and U11181 (N_11181,N_6915,N_5431);
nand U11182 (N_11182,N_6828,N_5812);
or U11183 (N_11183,N_7357,N_4790);
and U11184 (N_11184,N_6544,N_5669);
nor U11185 (N_11185,N_6486,N_4140);
nand U11186 (N_11186,N_6491,N_4387);
or U11187 (N_11187,N_7449,N_6925);
or U11188 (N_11188,N_6840,N_6524);
nor U11189 (N_11189,N_7717,N_6765);
or U11190 (N_11190,N_6066,N_5356);
nand U11191 (N_11191,N_5055,N_4422);
nor U11192 (N_11192,N_4911,N_6023);
nor U11193 (N_11193,N_5541,N_6114);
and U11194 (N_11194,N_4872,N_5493);
nand U11195 (N_11195,N_4498,N_7608);
or U11196 (N_11196,N_5656,N_7405);
or U11197 (N_11197,N_4967,N_4345);
xor U11198 (N_11198,N_5221,N_4517);
or U11199 (N_11199,N_5610,N_7565);
nand U11200 (N_11200,N_7431,N_4205);
or U11201 (N_11201,N_6075,N_6753);
or U11202 (N_11202,N_7327,N_6822);
xnor U11203 (N_11203,N_7464,N_6961);
nand U11204 (N_11204,N_7642,N_4250);
nor U11205 (N_11205,N_4953,N_5014);
nand U11206 (N_11206,N_4911,N_4075);
nor U11207 (N_11207,N_7921,N_4287);
and U11208 (N_11208,N_4354,N_7018);
or U11209 (N_11209,N_5508,N_6738);
nor U11210 (N_11210,N_7971,N_4432);
and U11211 (N_11211,N_4750,N_7615);
nand U11212 (N_11212,N_5764,N_6657);
and U11213 (N_11213,N_6356,N_7554);
nor U11214 (N_11214,N_5919,N_7223);
and U11215 (N_11215,N_7748,N_5853);
or U11216 (N_11216,N_6495,N_5690);
or U11217 (N_11217,N_6401,N_4699);
or U11218 (N_11218,N_5595,N_4668);
and U11219 (N_11219,N_4586,N_5206);
nand U11220 (N_11220,N_7878,N_7913);
nand U11221 (N_11221,N_7007,N_6699);
and U11222 (N_11222,N_5963,N_6618);
and U11223 (N_11223,N_6476,N_5660);
or U11224 (N_11224,N_4398,N_6322);
xnor U11225 (N_11225,N_4871,N_7318);
or U11226 (N_11226,N_5384,N_5219);
nand U11227 (N_11227,N_5371,N_6371);
and U11228 (N_11228,N_4447,N_4217);
nand U11229 (N_11229,N_7649,N_6624);
and U11230 (N_11230,N_7681,N_4463);
xnor U11231 (N_11231,N_4498,N_6566);
nor U11232 (N_11232,N_7940,N_5745);
or U11233 (N_11233,N_6657,N_4483);
and U11234 (N_11234,N_5107,N_7216);
nor U11235 (N_11235,N_5710,N_4403);
and U11236 (N_11236,N_5756,N_7873);
nor U11237 (N_11237,N_6788,N_6632);
and U11238 (N_11238,N_5812,N_7231);
xor U11239 (N_11239,N_4977,N_5420);
and U11240 (N_11240,N_4023,N_4730);
nor U11241 (N_11241,N_5319,N_6995);
nand U11242 (N_11242,N_6427,N_6295);
xor U11243 (N_11243,N_4531,N_5769);
xnor U11244 (N_11244,N_5563,N_4891);
or U11245 (N_11245,N_6721,N_6393);
nor U11246 (N_11246,N_6240,N_7029);
nand U11247 (N_11247,N_7035,N_6761);
nor U11248 (N_11248,N_7250,N_4054);
xnor U11249 (N_11249,N_5265,N_7782);
xor U11250 (N_11250,N_6139,N_4966);
or U11251 (N_11251,N_6657,N_5463);
nor U11252 (N_11252,N_4038,N_6240);
nor U11253 (N_11253,N_5468,N_5752);
and U11254 (N_11254,N_7442,N_4944);
nand U11255 (N_11255,N_4608,N_7519);
and U11256 (N_11256,N_6100,N_5147);
nor U11257 (N_11257,N_7496,N_4337);
and U11258 (N_11258,N_4513,N_4840);
nand U11259 (N_11259,N_7457,N_7531);
nand U11260 (N_11260,N_5448,N_6985);
nor U11261 (N_11261,N_5622,N_5131);
nand U11262 (N_11262,N_5153,N_5395);
nor U11263 (N_11263,N_4126,N_6088);
nand U11264 (N_11264,N_5164,N_6017);
or U11265 (N_11265,N_5482,N_6318);
nand U11266 (N_11266,N_7255,N_7428);
nor U11267 (N_11267,N_5282,N_7639);
nor U11268 (N_11268,N_6728,N_7525);
nor U11269 (N_11269,N_6450,N_5023);
or U11270 (N_11270,N_6236,N_5949);
xnor U11271 (N_11271,N_6675,N_7294);
or U11272 (N_11272,N_6092,N_7748);
and U11273 (N_11273,N_4839,N_4421);
nand U11274 (N_11274,N_6706,N_7110);
or U11275 (N_11275,N_7075,N_7444);
and U11276 (N_11276,N_4181,N_7942);
xnor U11277 (N_11277,N_4738,N_4594);
nor U11278 (N_11278,N_7504,N_6450);
nand U11279 (N_11279,N_4501,N_6450);
xor U11280 (N_11280,N_5261,N_7631);
nor U11281 (N_11281,N_6098,N_7657);
or U11282 (N_11282,N_5415,N_7844);
or U11283 (N_11283,N_7256,N_4602);
or U11284 (N_11284,N_5473,N_5765);
or U11285 (N_11285,N_6154,N_7061);
or U11286 (N_11286,N_5652,N_7559);
and U11287 (N_11287,N_4577,N_5082);
nor U11288 (N_11288,N_4748,N_5329);
nand U11289 (N_11289,N_4653,N_6119);
nand U11290 (N_11290,N_7537,N_4710);
and U11291 (N_11291,N_4849,N_5411);
nor U11292 (N_11292,N_6146,N_4203);
or U11293 (N_11293,N_6084,N_6918);
or U11294 (N_11294,N_5960,N_7926);
xor U11295 (N_11295,N_6793,N_5659);
xnor U11296 (N_11296,N_4967,N_5372);
and U11297 (N_11297,N_7812,N_4486);
and U11298 (N_11298,N_4049,N_4463);
and U11299 (N_11299,N_5869,N_4352);
nor U11300 (N_11300,N_4944,N_6763);
or U11301 (N_11301,N_7437,N_7101);
and U11302 (N_11302,N_7449,N_4507);
or U11303 (N_11303,N_5613,N_7966);
nor U11304 (N_11304,N_5544,N_4504);
or U11305 (N_11305,N_4617,N_4394);
nor U11306 (N_11306,N_4019,N_6589);
or U11307 (N_11307,N_5359,N_7970);
or U11308 (N_11308,N_7397,N_7910);
and U11309 (N_11309,N_5862,N_5211);
nand U11310 (N_11310,N_4798,N_7558);
xnor U11311 (N_11311,N_5367,N_6814);
nor U11312 (N_11312,N_6168,N_7195);
and U11313 (N_11313,N_6293,N_5546);
or U11314 (N_11314,N_6740,N_6777);
nand U11315 (N_11315,N_7667,N_7295);
nor U11316 (N_11316,N_7834,N_7690);
or U11317 (N_11317,N_6010,N_6888);
or U11318 (N_11318,N_5248,N_7557);
xnor U11319 (N_11319,N_6461,N_4857);
or U11320 (N_11320,N_4587,N_5350);
or U11321 (N_11321,N_4668,N_7497);
xor U11322 (N_11322,N_6100,N_5705);
or U11323 (N_11323,N_7044,N_5908);
or U11324 (N_11324,N_4744,N_6490);
nand U11325 (N_11325,N_4493,N_5941);
and U11326 (N_11326,N_7397,N_5488);
and U11327 (N_11327,N_5110,N_7552);
or U11328 (N_11328,N_7702,N_5394);
nor U11329 (N_11329,N_4402,N_7876);
nand U11330 (N_11330,N_6362,N_6051);
nand U11331 (N_11331,N_7020,N_7239);
xor U11332 (N_11332,N_4882,N_5606);
or U11333 (N_11333,N_7521,N_6365);
nor U11334 (N_11334,N_5775,N_6157);
and U11335 (N_11335,N_6802,N_6715);
nand U11336 (N_11336,N_7536,N_4617);
nand U11337 (N_11337,N_5302,N_5923);
and U11338 (N_11338,N_7904,N_6971);
nand U11339 (N_11339,N_4521,N_6463);
nor U11340 (N_11340,N_7128,N_5503);
or U11341 (N_11341,N_7729,N_5187);
and U11342 (N_11342,N_5905,N_6090);
and U11343 (N_11343,N_6380,N_7391);
nand U11344 (N_11344,N_4946,N_4514);
or U11345 (N_11345,N_7056,N_4356);
xor U11346 (N_11346,N_5191,N_6140);
nor U11347 (N_11347,N_6372,N_4792);
nand U11348 (N_11348,N_5993,N_7239);
nor U11349 (N_11349,N_6764,N_5753);
nor U11350 (N_11350,N_7730,N_6488);
and U11351 (N_11351,N_7864,N_6177);
and U11352 (N_11352,N_7887,N_7171);
and U11353 (N_11353,N_6376,N_6627);
nand U11354 (N_11354,N_6206,N_5230);
nor U11355 (N_11355,N_6159,N_6299);
xnor U11356 (N_11356,N_6599,N_7099);
or U11357 (N_11357,N_7073,N_6553);
and U11358 (N_11358,N_6191,N_5882);
nand U11359 (N_11359,N_7307,N_6726);
nor U11360 (N_11360,N_7997,N_5371);
nand U11361 (N_11361,N_7327,N_4989);
xnor U11362 (N_11362,N_5992,N_5079);
nor U11363 (N_11363,N_4667,N_5717);
xnor U11364 (N_11364,N_5808,N_7634);
nor U11365 (N_11365,N_6856,N_4649);
and U11366 (N_11366,N_7824,N_7439);
nand U11367 (N_11367,N_6457,N_4738);
and U11368 (N_11368,N_6433,N_7891);
and U11369 (N_11369,N_6255,N_5819);
xnor U11370 (N_11370,N_4868,N_6325);
or U11371 (N_11371,N_5250,N_6576);
xor U11372 (N_11372,N_6970,N_6049);
xnor U11373 (N_11373,N_4487,N_4401);
nand U11374 (N_11374,N_4163,N_6999);
xnor U11375 (N_11375,N_6556,N_4843);
nor U11376 (N_11376,N_5928,N_4741);
and U11377 (N_11377,N_4693,N_6236);
or U11378 (N_11378,N_5048,N_5258);
nor U11379 (N_11379,N_4360,N_4446);
and U11380 (N_11380,N_7857,N_5145);
nor U11381 (N_11381,N_6573,N_6673);
or U11382 (N_11382,N_6681,N_4543);
or U11383 (N_11383,N_6617,N_5803);
nor U11384 (N_11384,N_4254,N_5172);
nand U11385 (N_11385,N_5769,N_6009);
nand U11386 (N_11386,N_4901,N_4741);
nor U11387 (N_11387,N_7621,N_5154);
nor U11388 (N_11388,N_6524,N_5371);
or U11389 (N_11389,N_7315,N_4692);
nor U11390 (N_11390,N_5604,N_4624);
nand U11391 (N_11391,N_6113,N_6490);
nand U11392 (N_11392,N_7048,N_4092);
xnor U11393 (N_11393,N_4309,N_7595);
nor U11394 (N_11394,N_7349,N_4556);
nand U11395 (N_11395,N_5166,N_6398);
nand U11396 (N_11396,N_6185,N_5542);
nand U11397 (N_11397,N_4719,N_6881);
or U11398 (N_11398,N_7500,N_4141);
nor U11399 (N_11399,N_7183,N_4246);
or U11400 (N_11400,N_5788,N_7266);
nand U11401 (N_11401,N_6809,N_7590);
and U11402 (N_11402,N_4493,N_4699);
or U11403 (N_11403,N_5232,N_7714);
or U11404 (N_11404,N_7128,N_6772);
or U11405 (N_11405,N_5234,N_5947);
and U11406 (N_11406,N_4855,N_4787);
or U11407 (N_11407,N_7991,N_5771);
nand U11408 (N_11408,N_4888,N_6538);
nor U11409 (N_11409,N_6383,N_4880);
and U11410 (N_11410,N_6598,N_4223);
and U11411 (N_11411,N_7861,N_6374);
nor U11412 (N_11412,N_6390,N_6843);
nand U11413 (N_11413,N_4531,N_4882);
or U11414 (N_11414,N_6200,N_5385);
or U11415 (N_11415,N_4767,N_7956);
or U11416 (N_11416,N_6788,N_6802);
nor U11417 (N_11417,N_5941,N_6329);
or U11418 (N_11418,N_7695,N_6184);
nand U11419 (N_11419,N_4128,N_7150);
and U11420 (N_11420,N_7214,N_5970);
and U11421 (N_11421,N_7414,N_5123);
or U11422 (N_11422,N_4752,N_7139);
nand U11423 (N_11423,N_6788,N_7900);
nand U11424 (N_11424,N_5281,N_5889);
and U11425 (N_11425,N_5446,N_6712);
nand U11426 (N_11426,N_5850,N_6819);
nand U11427 (N_11427,N_4975,N_6881);
nand U11428 (N_11428,N_5976,N_5203);
and U11429 (N_11429,N_5153,N_6998);
and U11430 (N_11430,N_4555,N_4985);
and U11431 (N_11431,N_5669,N_6169);
and U11432 (N_11432,N_5913,N_4278);
and U11433 (N_11433,N_7114,N_4514);
nand U11434 (N_11434,N_7530,N_4056);
and U11435 (N_11435,N_6715,N_6840);
nor U11436 (N_11436,N_7936,N_7318);
or U11437 (N_11437,N_5261,N_7010);
or U11438 (N_11438,N_7188,N_4038);
and U11439 (N_11439,N_7863,N_5388);
nand U11440 (N_11440,N_7246,N_5458);
or U11441 (N_11441,N_4288,N_5742);
or U11442 (N_11442,N_4247,N_6876);
and U11443 (N_11443,N_4666,N_5282);
nor U11444 (N_11444,N_7886,N_5262);
or U11445 (N_11445,N_6347,N_5331);
or U11446 (N_11446,N_7857,N_6807);
or U11447 (N_11447,N_7667,N_5468);
nor U11448 (N_11448,N_6317,N_4606);
nor U11449 (N_11449,N_5550,N_7633);
or U11450 (N_11450,N_4882,N_5226);
or U11451 (N_11451,N_6079,N_4721);
or U11452 (N_11452,N_4004,N_7956);
xnor U11453 (N_11453,N_4157,N_5992);
xor U11454 (N_11454,N_7081,N_7273);
and U11455 (N_11455,N_5611,N_4487);
nand U11456 (N_11456,N_5927,N_4974);
xor U11457 (N_11457,N_7922,N_7357);
nor U11458 (N_11458,N_7346,N_4326);
and U11459 (N_11459,N_4066,N_6400);
or U11460 (N_11460,N_6400,N_7033);
nor U11461 (N_11461,N_4720,N_5790);
nor U11462 (N_11462,N_5165,N_5086);
and U11463 (N_11463,N_7628,N_7794);
or U11464 (N_11464,N_5211,N_5788);
nor U11465 (N_11465,N_6246,N_6773);
or U11466 (N_11466,N_5869,N_6423);
or U11467 (N_11467,N_6889,N_7747);
and U11468 (N_11468,N_6392,N_7734);
nor U11469 (N_11469,N_6176,N_6203);
nand U11470 (N_11470,N_4565,N_5992);
nand U11471 (N_11471,N_6126,N_6586);
nor U11472 (N_11472,N_7549,N_6805);
and U11473 (N_11473,N_6304,N_7022);
or U11474 (N_11474,N_5854,N_4468);
nor U11475 (N_11475,N_7132,N_5543);
nand U11476 (N_11476,N_6451,N_5497);
nor U11477 (N_11477,N_4076,N_6928);
and U11478 (N_11478,N_4730,N_6322);
xnor U11479 (N_11479,N_6610,N_4408);
nand U11480 (N_11480,N_6626,N_5922);
or U11481 (N_11481,N_5798,N_4289);
nand U11482 (N_11482,N_6235,N_4659);
xor U11483 (N_11483,N_7329,N_5390);
nand U11484 (N_11484,N_4458,N_6412);
or U11485 (N_11485,N_5051,N_5349);
or U11486 (N_11486,N_4416,N_4118);
and U11487 (N_11487,N_7319,N_6015);
or U11488 (N_11488,N_6738,N_7000);
nor U11489 (N_11489,N_6153,N_4421);
nor U11490 (N_11490,N_7914,N_6212);
and U11491 (N_11491,N_5891,N_4168);
nor U11492 (N_11492,N_6960,N_7706);
and U11493 (N_11493,N_6111,N_5536);
nand U11494 (N_11494,N_7939,N_4454);
or U11495 (N_11495,N_4875,N_7326);
nand U11496 (N_11496,N_7285,N_4901);
or U11497 (N_11497,N_5296,N_7051);
nor U11498 (N_11498,N_7250,N_6721);
xor U11499 (N_11499,N_5114,N_4908);
nand U11500 (N_11500,N_4987,N_7837);
nand U11501 (N_11501,N_7039,N_6254);
nor U11502 (N_11502,N_6171,N_5029);
nand U11503 (N_11503,N_4895,N_6262);
nor U11504 (N_11504,N_4331,N_6544);
xnor U11505 (N_11505,N_6979,N_4607);
nand U11506 (N_11506,N_5104,N_6190);
nor U11507 (N_11507,N_4806,N_7074);
nor U11508 (N_11508,N_6052,N_5397);
and U11509 (N_11509,N_6206,N_7151);
nand U11510 (N_11510,N_5487,N_6763);
and U11511 (N_11511,N_7521,N_4772);
and U11512 (N_11512,N_6881,N_7660);
xor U11513 (N_11513,N_4394,N_7032);
nand U11514 (N_11514,N_5574,N_5963);
and U11515 (N_11515,N_5852,N_6992);
or U11516 (N_11516,N_4226,N_4872);
nor U11517 (N_11517,N_6302,N_5517);
nor U11518 (N_11518,N_6991,N_7506);
nor U11519 (N_11519,N_6894,N_5846);
nand U11520 (N_11520,N_6348,N_5401);
nand U11521 (N_11521,N_6781,N_7006);
nor U11522 (N_11522,N_4586,N_5153);
nor U11523 (N_11523,N_6232,N_6079);
nand U11524 (N_11524,N_7047,N_5472);
nor U11525 (N_11525,N_7887,N_7088);
or U11526 (N_11526,N_7550,N_5972);
nor U11527 (N_11527,N_5978,N_6321);
nor U11528 (N_11528,N_6326,N_4883);
nand U11529 (N_11529,N_5505,N_5177);
and U11530 (N_11530,N_6504,N_4554);
nand U11531 (N_11531,N_7656,N_7379);
nand U11532 (N_11532,N_7705,N_5931);
xnor U11533 (N_11533,N_4604,N_5356);
nor U11534 (N_11534,N_4063,N_5385);
nand U11535 (N_11535,N_6531,N_5247);
or U11536 (N_11536,N_7463,N_4758);
and U11537 (N_11537,N_6594,N_4958);
nor U11538 (N_11538,N_4994,N_4352);
or U11539 (N_11539,N_4348,N_7417);
and U11540 (N_11540,N_7135,N_5949);
xor U11541 (N_11541,N_5410,N_4941);
nand U11542 (N_11542,N_7607,N_6566);
and U11543 (N_11543,N_6840,N_4176);
nand U11544 (N_11544,N_7542,N_4625);
and U11545 (N_11545,N_4135,N_5392);
nor U11546 (N_11546,N_4095,N_7239);
nand U11547 (N_11547,N_7618,N_5239);
nor U11548 (N_11548,N_6310,N_7474);
xnor U11549 (N_11549,N_7526,N_5376);
and U11550 (N_11550,N_4361,N_6958);
nor U11551 (N_11551,N_5716,N_5919);
nor U11552 (N_11552,N_4844,N_5106);
nor U11553 (N_11553,N_4689,N_4341);
nor U11554 (N_11554,N_5497,N_4113);
and U11555 (N_11555,N_7889,N_5680);
nand U11556 (N_11556,N_4744,N_5599);
and U11557 (N_11557,N_7158,N_7769);
nor U11558 (N_11558,N_6886,N_7215);
nand U11559 (N_11559,N_7940,N_6423);
and U11560 (N_11560,N_4215,N_4716);
nor U11561 (N_11561,N_6737,N_6185);
and U11562 (N_11562,N_6167,N_4415);
nor U11563 (N_11563,N_5168,N_4636);
xnor U11564 (N_11564,N_6319,N_4765);
nand U11565 (N_11565,N_7896,N_5940);
nor U11566 (N_11566,N_4259,N_6116);
or U11567 (N_11567,N_7867,N_4258);
nor U11568 (N_11568,N_5852,N_6135);
nand U11569 (N_11569,N_7334,N_7771);
nor U11570 (N_11570,N_7666,N_5457);
nand U11571 (N_11571,N_6133,N_5776);
nor U11572 (N_11572,N_6528,N_6342);
or U11573 (N_11573,N_6426,N_5875);
nand U11574 (N_11574,N_7632,N_6966);
nand U11575 (N_11575,N_6731,N_5359);
or U11576 (N_11576,N_6686,N_4025);
nand U11577 (N_11577,N_4133,N_4023);
nor U11578 (N_11578,N_6023,N_4932);
or U11579 (N_11579,N_5468,N_5660);
or U11580 (N_11580,N_4397,N_4487);
or U11581 (N_11581,N_5747,N_4725);
or U11582 (N_11582,N_7640,N_5555);
nor U11583 (N_11583,N_6284,N_5745);
nor U11584 (N_11584,N_5615,N_7498);
and U11585 (N_11585,N_5605,N_4627);
and U11586 (N_11586,N_5167,N_7679);
nor U11587 (N_11587,N_6438,N_6336);
and U11588 (N_11588,N_4605,N_7291);
nand U11589 (N_11589,N_6998,N_5783);
nor U11590 (N_11590,N_7213,N_5552);
nand U11591 (N_11591,N_6308,N_7669);
nand U11592 (N_11592,N_7943,N_5620);
and U11593 (N_11593,N_7300,N_6394);
and U11594 (N_11594,N_7213,N_6768);
and U11595 (N_11595,N_7403,N_6216);
nand U11596 (N_11596,N_6397,N_6099);
nor U11597 (N_11597,N_6757,N_6645);
xnor U11598 (N_11598,N_4035,N_7877);
nor U11599 (N_11599,N_5580,N_6055);
nor U11600 (N_11600,N_6898,N_4059);
nor U11601 (N_11601,N_4472,N_5233);
or U11602 (N_11602,N_4949,N_5386);
nand U11603 (N_11603,N_7045,N_5166);
or U11604 (N_11604,N_5945,N_4441);
or U11605 (N_11605,N_5128,N_7620);
nor U11606 (N_11606,N_7286,N_5381);
or U11607 (N_11607,N_6162,N_5476);
and U11608 (N_11608,N_5629,N_7886);
or U11609 (N_11609,N_5473,N_7037);
and U11610 (N_11610,N_7012,N_5734);
and U11611 (N_11611,N_4127,N_4134);
and U11612 (N_11612,N_5620,N_7728);
nor U11613 (N_11613,N_6466,N_6004);
nand U11614 (N_11614,N_5427,N_6436);
nand U11615 (N_11615,N_4205,N_6431);
or U11616 (N_11616,N_6755,N_5104);
xnor U11617 (N_11617,N_5967,N_6599);
and U11618 (N_11618,N_5764,N_5593);
nand U11619 (N_11619,N_5757,N_4509);
xor U11620 (N_11620,N_4379,N_4771);
or U11621 (N_11621,N_7901,N_7255);
nand U11622 (N_11622,N_7106,N_5673);
and U11623 (N_11623,N_5280,N_4344);
nand U11624 (N_11624,N_4688,N_6958);
and U11625 (N_11625,N_7581,N_7254);
and U11626 (N_11626,N_5149,N_4360);
nand U11627 (N_11627,N_6283,N_7723);
nor U11628 (N_11628,N_4179,N_7078);
and U11629 (N_11629,N_6643,N_4210);
nor U11630 (N_11630,N_7594,N_4115);
nand U11631 (N_11631,N_7059,N_6601);
nor U11632 (N_11632,N_6845,N_4697);
nand U11633 (N_11633,N_4346,N_5592);
and U11634 (N_11634,N_4450,N_6448);
and U11635 (N_11635,N_7447,N_4489);
and U11636 (N_11636,N_4505,N_6036);
or U11637 (N_11637,N_6606,N_6588);
nand U11638 (N_11638,N_4214,N_6340);
nor U11639 (N_11639,N_5837,N_5431);
xnor U11640 (N_11640,N_4764,N_5604);
nand U11641 (N_11641,N_6857,N_6683);
nand U11642 (N_11642,N_5258,N_5558);
nor U11643 (N_11643,N_5528,N_5664);
and U11644 (N_11644,N_5345,N_7371);
or U11645 (N_11645,N_5110,N_7901);
and U11646 (N_11646,N_4080,N_6702);
and U11647 (N_11647,N_4353,N_4144);
nor U11648 (N_11648,N_5750,N_5300);
xor U11649 (N_11649,N_7779,N_4320);
nand U11650 (N_11650,N_6139,N_6457);
or U11651 (N_11651,N_5756,N_5761);
nor U11652 (N_11652,N_5584,N_4050);
or U11653 (N_11653,N_5470,N_4357);
nor U11654 (N_11654,N_7807,N_5262);
xor U11655 (N_11655,N_4008,N_4313);
nand U11656 (N_11656,N_7047,N_5421);
and U11657 (N_11657,N_7538,N_5346);
and U11658 (N_11658,N_6531,N_5674);
or U11659 (N_11659,N_5030,N_5818);
and U11660 (N_11660,N_6100,N_5752);
nand U11661 (N_11661,N_6614,N_5811);
and U11662 (N_11662,N_7937,N_5215);
and U11663 (N_11663,N_7247,N_4961);
and U11664 (N_11664,N_6642,N_7564);
and U11665 (N_11665,N_6697,N_7126);
and U11666 (N_11666,N_5239,N_6050);
or U11667 (N_11667,N_5990,N_6598);
and U11668 (N_11668,N_4813,N_6936);
nand U11669 (N_11669,N_4119,N_4634);
or U11670 (N_11670,N_7267,N_4270);
nor U11671 (N_11671,N_6534,N_5901);
or U11672 (N_11672,N_6765,N_6849);
nand U11673 (N_11673,N_6199,N_6051);
nand U11674 (N_11674,N_5324,N_6781);
or U11675 (N_11675,N_4705,N_5073);
or U11676 (N_11676,N_5330,N_6258);
and U11677 (N_11677,N_4931,N_7804);
and U11678 (N_11678,N_7149,N_5049);
nor U11679 (N_11679,N_7922,N_4676);
or U11680 (N_11680,N_4696,N_4326);
and U11681 (N_11681,N_7189,N_7554);
nand U11682 (N_11682,N_5261,N_6836);
or U11683 (N_11683,N_4530,N_6714);
nand U11684 (N_11684,N_6276,N_6633);
nand U11685 (N_11685,N_6117,N_4555);
nor U11686 (N_11686,N_6686,N_5824);
or U11687 (N_11687,N_7192,N_7693);
and U11688 (N_11688,N_4692,N_4691);
or U11689 (N_11689,N_4915,N_7788);
and U11690 (N_11690,N_7510,N_5404);
nor U11691 (N_11691,N_6266,N_6245);
nor U11692 (N_11692,N_6707,N_7499);
xor U11693 (N_11693,N_6102,N_6791);
or U11694 (N_11694,N_7299,N_4146);
nand U11695 (N_11695,N_6018,N_5477);
or U11696 (N_11696,N_4925,N_5249);
xnor U11697 (N_11697,N_6052,N_7479);
nand U11698 (N_11698,N_5082,N_4757);
or U11699 (N_11699,N_6262,N_7599);
nand U11700 (N_11700,N_4024,N_7711);
and U11701 (N_11701,N_5449,N_6715);
nand U11702 (N_11702,N_7364,N_4975);
or U11703 (N_11703,N_4752,N_7578);
nor U11704 (N_11704,N_6908,N_7490);
or U11705 (N_11705,N_5038,N_6385);
and U11706 (N_11706,N_6255,N_7665);
xor U11707 (N_11707,N_5151,N_6002);
xnor U11708 (N_11708,N_7251,N_4953);
and U11709 (N_11709,N_4388,N_5256);
and U11710 (N_11710,N_5935,N_4630);
and U11711 (N_11711,N_5591,N_5802);
nand U11712 (N_11712,N_6858,N_4790);
or U11713 (N_11713,N_7672,N_7318);
nand U11714 (N_11714,N_4134,N_6911);
xnor U11715 (N_11715,N_4583,N_7038);
nand U11716 (N_11716,N_5709,N_4789);
nand U11717 (N_11717,N_7999,N_4504);
nor U11718 (N_11718,N_6862,N_6164);
nand U11719 (N_11719,N_5100,N_5759);
nor U11720 (N_11720,N_4283,N_5502);
nand U11721 (N_11721,N_7011,N_7481);
nand U11722 (N_11722,N_7480,N_7836);
nor U11723 (N_11723,N_5849,N_4632);
and U11724 (N_11724,N_5785,N_6766);
nor U11725 (N_11725,N_6901,N_7866);
nand U11726 (N_11726,N_4412,N_5414);
nand U11727 (N_11727,N_6704,N_7490);
and U11728 (N_11728,N_4615,N_5756);
or U11729 (N_11729,N_6589,N_6848);
and U11730 (N_11730,N_5515,N_7728);
and U11731 (N_11731,N_5414,N_6820);
xnor U11732 (N_11732,N_6873,N_4865);
or U11733 (N_11733,N_7512,N_7858);
and U11734 (N_11734,N_6407,N_7951);
or U11735 (N_11735,N_5578,N_5048);
and U11736 (N_11736,N_4170,N_5993);
and U11737 (N_11737,N_7782,N_6567);
and U11738 (N_11738,N_4257,N_4522);
or U11739 (N_11739,N_6914,N_7322);
xor U11740 (N_11740,N_6563,N_7603);
nor U11741 (N_11741,N_4861,N_7234);
nor U11742 (N_11742,N_7637,N_4740);
and U11743 (N_11743,N_4126,N_6377);
and U11744 (N_11744,N_4367,N_6566);
nor U11745 (N_11745,N_5615,N_6835);
and U11746 (N_11746,N_5879,N_6710);
xor U11747 (N_11747,N_4792,N_5690);
or U11748 (N_11748,N_4508,N_6226);
nor U11749 (N_11749,N_6887,N_7415);
nor U11750 (N_11750,N_6105,N_4950);
nand U11751 (N_11751,N_5103,N_4249);
xor U11752 (N_11752,N_5481,N_4957);
or U11753 (N_11753,N_7480,N_6038);
nand U11754 (N_11754,N_7482,N_5827);
xor U11755 (N_11755,N_6799,N_6597);
nand U11756 (N_11756,N_6798,N_6029);
and U11757 (N_11757,N_6710,N_7378);
nand U11758 (N_11758,N_4524,N_4551);
nor U11759 (N_11759,N_4824,N_4999);
nor U11760 (N_11760,N_4420,N_7666);
xor U11761 (N_11761,N_7550,N_5599);
and U11762 (N_11762,N_6241,N_6714);
nor U11763 (N_11763,N_6226,N_6025);
and U11764 (N_11764,N_4743,N_5126);
and U11765 (N_11765,N_5769,N_5729);
nor U11766 (N_11766,N_4517,N_5175);
nand U11767 (N_11767,N_7927,N_5420);
and U11768 (N_11768,N_6049,N_7528);
nand U11769 (N_11769,N_7071,N_7742);
nand U11770 (N_11770,N_5070,N_6428);
or U11771 (N_11771,N_4201,N_7932);
or U11772 (N_11772,N_5043,N_6413);
nand U11773 (N_11773,N_4396,N_6259);
and U11774 (N_11774,N_4978,N_4378);
or U11775 (N_11775,N_4357,N_4898);
nor U11776 (N_11776,N_4465,N_6390);
or U11777 (N_11777,N_6602,N_5734);
nand U11778 (N_11778,N_6665,N_5934);
and U11779 (N_11779,N_4492,N_5580);
and U11780 (N_11780,N_7985,N_6318);
nor U11781 (N_11781,N_5707,N_5383);
or U11782 (N_11782,N_7338,N_6094);
xnor U11783 (N_11783,N_4212,N_7384);
or U11784 (N_11784,N_6704,N_6645);
nand U11785 (N_11785,N_7740,N_6668);
and U11786 (N_11786,N_6232,N_7978);
and U11787 (N_11787,N_7664,N_5869);
nand U11788 (N_11788,N_4822,N_6294);
or U11789 (N_11789,N_5169,N_7190);
nand U11790 (N_11790,N_4878,N_4053);
nand U11791 (N_11791,N_6255,N_4107);
xor U11792 (N_11792,N_6349,N_7914);
and U11793 (N_11793,N_5778,N_7599);
nand U11794 (N_11794,N_4992,N_6004);
or U11795 (N_11795,N_5902,N_7455);
or U11796 (N_11796,N_6524,N_5429);
or U11797 (N_11797,N_6421,N_4114);
or U11798 (N_11798,N_7410,N_6276);
nor U11799 (N_11799,N_6521,N_6952);
or U11800 (N_11800,N_5539,N_5876);
and U11801 (N_11801,N_4709,N_6816);
nor U11802 (N_11802,N_5816,N_7711);
nand U11803 (N_11803,N_7552,N_7714);
nand U11804 (N_11804,N_4230,N_7769);
or U11805 (N_11805,N_4538,N_4925);
and U11806 (N_11806,N_6529,N_4631);
or U11807 (N_11807,N_4756,N_7186);
nand U11808 (N_11808,N_5181,N_6362);
nor U11809 (N_11809,N_4173,N_7252);
nor U11810 (N_11810,N_6918,N_7887);
xnor U11811 (N_11811,N_7342,N_4508);
or U11812 (N_11812,N_6468,N_5627);
or U11813 (N_11813,N_5581,N_5208);
or U11814 (N_11814,N_6058,N_4140);
nor U11815 (N_11815,N_7170,N_4377);
nand U11816 (N_11816,N_7458,N_4532);
or U11817 (N_11817,N_7282,N_5355);
nor U11818 (N_11818,N_5739,N_5143);
nand U11819 (N_11819,N_6315,N_4611);
or U11820 (N_11820,N_5905,N_6628);
or U11821 (N_11821,N_5844,N_4668);
nor U11822 (N_11822,N_4916,N_5113);
xnor U11823 (N_11823,N_5262,N_4182);
xnor U11824 (N_11824,N_6393,N_7823);
nand U11825 (N_11825,N_4089,N_5802);
xor U11826 (N_11826,N_6450,N_6284);
or U11827 (N_11827,N_4249,N_6589);
and U11828 (N_11828,N_6785,N_5864);
or U11829 (N_11829,N_6890,N_4338);
nor U11830 (N_11830,N_6401,N_5754);
or U11831 (N_11831,N_5743,N_5316);
nand U11832 (N_11832,N_5969,N_6087);
and U11833 (N_11833,N_5235,N_6716);
nor U11834 (N_11834,N_7220,N_6390);
and U11835 (N_11835,N_4119,N_7227);
nor U11836 (N_11836,N_4114,N_4687);
nor U11837 (N_11837,N_4699,N_6727);
nand U11838 (N_11838,N_4540,N_7684);
nand U11839 (N_11839,N_4034,N_6733);
nor U11840 (N_11840,N_4480,N_4482);
nor U11841 (N_11841,N_7517,N_5618);
and U11842 (N_11842,N_7673,N_4102);
and U11843 (N_11843,N_6023,N_5019);
nand U11844 (N_11844,N_7539,N_4820);
nand U11845 (N_11845,N_5434,N_5793);
and U11846 (N_11846,N_6407,N_6974);
xnor U11847 (N_11847,N_4749,N_5976);
and U11848 (N_11848,N_4391,N_5972);
or U11849 (N_11849,N_5818,N_5564);
nor U11850 (N_11850,N_6581,N_4164);
nor U11851 (N_11851,N_4372,N_7144);
nand U11852 (N_11852,N_6822,N_7734);
nor U11853 (N_11853,N_7112,N_6033);
nand U11854 (N_11854,N_7058,N_7022);
or U11855 (N_11855,N_6103,N_6782);
nor U11856 (N_11856,N_7911,N_6134);
or U11857 (N_11857,N_4095,N_4741);
nor U11858 (N_11858,N_5093,N_4772);
nand U11859 (N_11859,N_7408,N_6748);
or U11860 (N_11860,N_5884,N_7528);
and U11861 (N_11861,N_6459,N_4976);
nand U11862 (N_11862,N_5493,N_6626);
xnor U11863 (N_11863,N_5152,N_4816);
xor U11864 (N_11864,N_4292,N_7806);
nand U11865 (N_11865,N_6826,N_7609);
or U11866 (N_11866,N_5031,N_5731);
or U11867 (N_11867,N_6086,N_7849);
nor U11868 (N_11868,N_6766,N_5139);
and U11869 (N_11869,N_5198,N_5650);
nor U11870 (N_11870,N_7033,N_6328);
nand U11871 (N_11871,N_6772,N_5711);
nor U11872 (N_11872,N_6217,N_5331);
or U11873 (N_11873,N_4154,N_6859);
and U11874 (N_11874,N_7585,N_6421);
nor U11875 (N_11875,N_4469,N_7531);
or U11876 (N_11876,N_6145,N_5763);
or U11877 (N_11877,N_4324,N_7621);
and U11878 (N_11878,N_7979,N_6253);
and U11879 (N_11879,N_4584,N_6848);
or U11880 (N_11880,N_4066,N_5664);
nand U11881 (N_11881,N_6497,N_7825);
and U11882 (N_11882,N_4092,N_4933);
or U11883 (N_11883,N_6008,N_6478);
xnor U11884 (N_11884,N_6461,N_6368);
nor U11885 (N_11885,N_6066,N_6653);
nor U11886 (N_11886,N_5778,N_6986);
nor U11887 (N_11887,N_4866,N_6703);
or U11888 (N_11888,N_6570,N_7702);
or U11889 (N_11889,N_5275,N_6772);
nand U11890 (N_11890,N_5618,N_6090);
and U11891 (N_11891,N_7063,N_5222);
and U11892 (N_11892,N_7236,N_4228);
xor U11893 (N_11893,N_7505,N_7703);
and U11894 (N_11894,N_5256,N_7184);
or U11895 (N_11895,N_5425,N_7449);
xnor U11896 (N_11896,N_7685,N_6025);
or U11897 (N_11897,N_6515,N_4295);
and U11898 (N_11898,N_5449,N_7278);
or U11899 (N_11899,N_4252,N_4807);
nor U11900 (N_11900,N_4512,N_5708);
xor U11901 (N_11901,N_7622,N_5304);
nand U11902 (N_11902,N_5090,N_5558);
or U11903 (N_11903,N_4658,N_5696);
nor U11904 (N_11904,N_5292,N_4184);
or U11905 (N_11905,N_4186,N_7492);
and U11906 (N_11906,N_5996,N_7152);
nand U11907 (N_11907,N_7989,N_7661);
nand U11908 (N_11908,N_4673,N_6126);
and U11909 (N_11909,N_6328,N_5550);
nor U11910 (N_11910,N_4064,N_7272);
nand U11911 (N_11911,N_7351,N_6114);
nor U11912 (N_11912,N_7513,N_6019);
and U11913 (N_11913,N_5071,N_5382);
or U11914 (N_11914,N_4220,N_6755);
nand U11915 (N_11915,N_6449,N_6981);
nor U11916 (N_11916,N_4886,N_7362);
and U11917 (N_11917,N_5586,N_6144);
nand U11918 (N_11918,N_5211,N_4687);
and U11919 (N_11919,N_7934,N_5248);
xnor U11920 (N_11920,N_4722,N_5692);
and U11921 (N_11921,N_7046,N_7186);
and U11922 (N_11922,N_5132,N_5147);
nor U11923 (N_11923,N_5458,N_6770);
or U11924 (N_11924,N_7544,N_7389);
nand U11925 (N_11925,N_7339,N_4172);
or U11926 (N_11926,N_6595,N_5020);
or U11927 (N_11927,N_4250,N_5302);
nor U11928 (N_11928,N_4747,N_5886);
and U11929 (N_11929,N_4008,N_5492);
nand U11930 (N_11930,N_7165,N_6163);
nand U11931 (N_11931,N_5384,N_6064);
and U11932 (N_11932,N_4713,N_4367);
nand U11933 (N_11933,N_5358,N_5586);
and U11934 (N_11934,N_5874,N_7420);
or U11935 (N_11935,N_4612,N_4097);
nor U11936 (N_11936,N_7489,N_4000);
and U11937 (N_11937,N_5574,N_6015);
and U11938 (N_11938,N_7744,N_5097);
nand U11939 (N_11939,N_4012,N_4382);
xor U11940 (N_11940,N_7286,N_4451);
nand U11941 (N_11941,N_4117,N_6855);
or U11942 (N_11942,N_7498,N_7425);
nor U11943 (N_11943,N_5467,N_5204);
nand U11944 (N_11944,N_7340,N_5576);
and U11945 (N_11945,N_4561,N_4610);
or U11946 (N_11946,N_5242,N_6096);
or U11947 (N_11947,N_4885,N_4870);
and U11948 (N_11948,N_4776,N_7318);
xnor U11949 (N_11949,N_5606,N_6626);
nor U11950 (N_11950,N_6616,N_6391);
nand U11951 (N_11951,N_4664,N_4319);
and U11952 (N_11952,N_5662,N_7367);
and U11953 (N_11953,N_5714,N_7384);
or U11954 (N_11954,N_6249,N_5591);
or U11955 (N_11955,N_4704,N_7018);
nand U11956 (N_11956,N_7807,N_4512);
nor U11957 (N_11957,N_7394,N_6339);
nor U11958 (N_11958,N_6244,N_5735);
nand U11959 (N_11959,N_5138,N_4329);
and U11960 (N_11960,N_5424,N_7748);
nand U11961 (N_11961,N_5080,N_5049);
or U11962 (N_11962,N_4091,N_5820);
xor U11963 (N_11963,N_4248,N_6907);
and U11964 (N_11964,N_7590,N_4017);
nor U11965 (N_11965,N_5800,N_6549);
nor U11966 (N_11966,N_4280,N_4176);
or U11967 (N_11967,N_6905,N_6283);
nor U11968 (N_11968,N_7356,N_7761);
or U11969 (N_11969,N_4320,N_5525);
or U11970 (N_11970,N_4715,N_6170);
and U11971 (N_11971,N_6414,N_4584);
nand U11972 (N_11972,N_6252,N_5683);
nand U11973 (N_11973,N_4574,N_7263);
and U11974 (N_11974,N_4462,N_6784);
nor U11975 (N_11975,N_5162,N_6337);
and U11976 (N_11976,N_4872,N_4100);
or U11977 (N_11977,N_7024,N_5746);
nand U11978 (N_11978,N_6205,N_6232);
nor U11979 (N_11979,N_7203,N_5712);
or U11980 (N_11980,N_7244,N_7919);
nand U11981 (N_11981,N_7130,N_7918);
and U11982 (N_11982,N_4078,N_6764);
and U11983 (N_11983,N_7326,N_7026);
xor U11984 (N_11984,N_6356,N_7882);
or U11985 (N_11985,N_7910,N_5638);
nand U11986 (N_11986,N_4500,N_6804);
nor U11987 (N_11987,N_6914,N_5652);
and U11988 (N_11988,N_5180,N_5181);
or U11989 (N_11989,N_7965,N_7758);
nand U11990 (N_11990,N_7747,N_5151);
nor U11991 (N_11991,N_4515,N_6040);
xnor U11992 (N_11992,N_5248,N_6843);
and U11993 (N_11993,N_4315,N_7054);
nor U11994 (N_11994,N_6184,N_7372);
nand U11995 (N_11995,N_4185,N_4425);
and U11996 (N_11996,N_7233,N_7491);
xnor U11997 (N_11997,N_6681,N_7152);
or U11998 (N_11998,N_6128,N_7903);
xor U11999 (N_11999,N_7338,N_5687);
or U12000 (N_12000,N_9228,N_9369);
nand U12001 (N_12001,N_11407,N_8222);
nand U12002 (N_12002,N_10749,N_8974);
and U12003 (N_12003,N_11273,N_10941);
nor U12004 (N_12004,N_8921,N_10835);
or U12005 (N_12005,N_8212,N_8582);
or U12006 (N_12006,N_9265,N_10585);
and U12007 (N_12007,N_8016,N_8751);
or U12008 (N_12008,N_11835,N_10610);
or U12009 (N_12009,N_11982,N_11399);
nor U12010 (N_12010,N_11760,N_8736);
or U12011 (N_12011,N_10712,N_10188);
nand U12012 (N_12012,N_11465,N_10074);
nor U12013 (N_12013,N_11627,N_8643);
nor U12014 (N_12014,N_9580,N_11496);
or U12015 (N_12015,N_11227,N_8127);
or U12016 (N_12016,N_8721,N_9170);
and U12017 (N_12017,N_11703,N_8515);
or U12018 (N_12018,N_10760,N_8350);
and U12019 (N_12019,N_8288,N_11120);
and U12020 (N_12020,N_8714,N_10916);
nand U12021 (N_12021,N_10391,N_11722);
xor U12022 (N_12022,N_11172,N_8894);
or U12023 (N_12023,N_10522,N_10840);
and U12024 (N_12024,N_9291,N_8730);
nand U12025 (N_12025,N_11428,N_10015);
and U12026 (N_12026,N_10626,N_10934);
xor U12027 (N_12027,N_9384,N_11926);
nor U12028 (N_12028,N_10380,N_9778);
nand U12029 (N_12029,N_10078,N_8346);
and U12030 (N_12030,N_10530,N_10531);
or U12031 (N_12031,N_9518,N_11584);
nor U12032 (N_12032,N_8740,N_11395);
nand U12033 (N_12033,N_10133,N_8103);
xor U12034 (N_12034,N_10359,N_8844);
or U12035 (N_12035,N_10955,N_9623);
nand U12036 (N_12036,N_10839,N_10231);
xor U12037 (N_12037,N_10647,N_10874);
nand U12038 (N_12038,N_11095,N_9978);
nand U12039 (N_12039,N_9264,N_11024);
nand U12040 (N_12040,N_10121,N_11951);
or U12041 (N_12041,N_10731,N_9593);
nor U12042 (N_12042,N_11650,N_11681);
nor U12043 (N_12043,N_10292,N_8654);
and U12044 (N_12044,N_10014,N_8951);
or U12045 (N_12045,N_9312,N_10221);
or U12046 (N_12046,N_9278,N_9124);
nor U12047 (N_12047,N_8939,N_9025);
nand U12048 (N_12048,N_8846,N_9241);
and U12049 (N_12049,N_8551,N_9434);
and U12050 (N_12050,N_9438,N_8697);
nand U12051 (N_12051,N_9780,N_11676);
xor U12052 (N_12052,N_9202,N_11664);
and U12053 (N_12053,N_9368,N_9811);
and U12054 (N_12054,N_11727,N_8683);
or U12055 (N_12055,N_9327,N_8649);
nand U12056 (N_12056,N_11740,N_10478);
and U12057 (N_12057,N_10498,N_10191);
and U12058 (N_12058,N_8702,N_10897);
nand U12059 (N_12059,N_11839,N_11992);
nor U12060 (N_12060,N_8457,N_9709);
nor U12061 (N_12061,N_9388,N_9948);
and U12062 (N_12062,N_11252,N_10118);
or U12063 (N_12063,N_10947,N_11777);
nor U12064 (N_12064,N_8087,N_8512);
xnor U12065 (N_12065,N_9804,N_8318);
nand U12066 (N_12066,N_10108,N_11006);
and U12067 (N_12067,N_11848,N_11483);
nand U12068 (N_12068,N_10989,N_8991);
nand U12069 (N_12069,N_8419,N_8597);
or U12070 (N_12070,N_8246,N_11343);
nand U12071 (N_12071,N_9850,N_9561);
nor U12072 (N_12072,N_11797,N_9942);
nor U12073 (N_12073,N_11861,N_9796);
xnor U12074 (N_12074,N_9949,N_8647);
nor U12075 (N_12075,N_11271,N_10907);
or U12076 (N_12076,N_11813,N_8373);
nand U12077 (N_12077,N_9958,N_10476);
nand U12078 (N_12078,N_10434,N_8653);
nand U12079 (N_12079,N_9827,N_11278);
and U12080 (N_12080,N_11738,N_10379);
nor U12081 (N_12081,N_8577,N_9238);
nor U12082 (N_12082,N_10335,N_8453);
nand U12083 (N_12083,N_11964,N_10643);
nand U12084 (N_12084,N_10573,N_10136);
and U12085 (N_12085,N_9073,N_8100);
and U12086 (N_12086,N_10737,N_10253);
and U12087 (N_12087,N_9766,N_9122);
nand U12088 (N_12088,N_9716,N_9583);
nand U12089 (N_12089,N_11834,N_10879);
nand U12090 (N_12090,N_8726,N_8251);
nand U12091 (N_12091,N_11542,N_8285);
nor U12092 (N_12092,N_9159,N_8628);
nor U12093 (N_12093,N_8341,N_10134);
nand U12094 (N_12094,N_9431,N_8106);
nand U12095 (N_12095,N_9531,N_11218);
and U12096 (N_12096,N_8078,N_8071);
nand U12097 (N_12097,N_11558,N_11036);
or U12098 (N_12098,N_8493,N_9450);
and U12099 (N_12099,N_10742,N_11642);
nand U12100 (N_12100,N_11795,N_9281);
or U12101 (N_12101,N_8096,N_8933);
nand U12102 (N_12102,N_9986,N_10356);
and U12103 (N_12103,N_10795,N_9971);
or U12104 (N_12104,N_10022,N_11305);
nand U12105 (N_12105,N_8445,N_9497);
nor U12106 (N_12106,N_8215,N_10666);
nor U12107 (N_12107,N_10618,N_9868);
and U12108 (N_12108,N_9755,N_9399);
nor U12109 (N_12109,N_9220,N_10741);
and U12110 (N_12110,N_8172,N_11893);
and U12111 (N_12111,N_10200,N_10197);
or U12112 (N_12112,N_10606,N_8990);
and U12113 (N_12113,N_11934,N_8710);
and U12114 (N_12114,N_8830,N_9364);
nand U12115 (N_12115,N_8323,N_9818);
nor U12116 (N_12116,N_8422,N_10347);
and U12117 (N_12117,N_11240,N_8541);
nor U12118 (N_12118,N_9671,N_9663);
and U12119 (N_12119,N_10710,N_10398);
and U12120 (N_12120,N_10541,N_10894);
and U12121 (N_12121,N_9582,N_10295);
or U12122 (N_12122,N_11264,N_9000);
nand U12123 (N_12123,N_10457,N_8178);
xnor U12124 (N_12124,N_9683,N_8790);
nand U12125 (N_12125,N_9690,N_8755);
nor U12126 (N_12126,N_9395,N_10829);
xnor U12127 (N_12127,N_11393,N_10613);
and U12128 (N_12128,N_9039,N_8182);
nor U12129 (N_12129,N_11942,N_8104);
nor U12130 (N_12130,N_10405,N_10274);
nor U12131 (N_12131,N_11787,N_10285);
and U12132 (N_12132,N_10538,N_8188);
and U12133 (N_12133,N_9844,N_8042);
xnor U12134 (N_12134,N_9062,N_8009);
xnor U12135 (N_12135,N_11699,N_8336);
or U12136 (N_12136,N_8584,N_11220);
nand U12137 (N_12137,N_11749,N_11160);
or U12138 (N_12138,N_11648,N_8191);
or U12139 (N_12139,N_10755,N_10848);
nor U12140 (N_12140,N_10272,N_9400);
nand U12141 (N_12141,N_10492,N_8248);
or U12142 (N_12142,N_10901,N_10583);
xnor U12143 (N_12143,N_8829,N_10066);
and U12144 (N_12144,N_11471,N_8081);
nor U12145 (N_12145,N_8559,N_11451);
nor U12146 (N_12146,N_10519,N_10466);
or U12147 (N_12147,N_9102,N_10709);
nor U12148 (N_12148,N_10876,N_9689);
nor U12149 (N_12149,N_10552,N_9240);
and U12150 (N_12150,N_11728,N_11423);
or U12151 (N_12151,N_11838,N_11279);
nor U12152 (N_12152,N_10609,N_11513);
and U12153 (N_12153,N_8168,N_11157);
nor U12154 (N_12154,N_11463,N_10770);
nor U12155 (N_12155,N_10301,N_10058);
nand U12156 (N_12156,N_9514,N_10224);
nor U12157 (N_12157,N_11309,N_9767);
or U12158 (N_12158,N_11236,N_10338);
xor U12159 (N_12159,N_8332,N_9317);
and U12160 (N_12160,N_11411,N_11497);
and U12161 (N_12161,N_11198,N_10497);
and U12162 (N_12162,N_8851,N_10308);
and U12163 (N_12163,N_10238,N_9157);
and U12164 (N_12164,N_8136,N_8708);
nand U12165 (N_12165,N_10304,N_8057);
nand U12166 (N_12166,N_11621,N_8499);
or U12167 (N_12167,N_8214,N_11166);
and U12168 (N_12168,N_8548,N_8496);
nor U12169 (N_12169,N_9807,N_9425);
or U12170 (N_12170,N_10496,N_8902);
or U12171 (N_12171,N_10079,N_9307);
nand U12172 (N_12172,N_10441,N_10184);
or U12173 (N_12173,N_11444,N_8865);
nor U12174 (N_12174,N_10299,N_10411);
and U12175 (N_12175,N_10378,N_9888);
or U12176 (N_12176,N_9511,N_8839);
or U12177 (N_12177,N_11800,N_9776);
xnor U12178 (N_12178,N_9866,N_9253);
and U12179 (N_12179,N_10882,N_9761);
and U12180 (N_12180,N_9218,N_11080);
and U12181 (N_12181,N_9254,N_8429);
xnor U12182 (N_12182,N_11223,N_11832);
or U12183 (N_12183,N_8281,N_11689);
and U12184 (N_12184,N_9084,N_8623);
or U12185 (N_12185,N_8473,N_8211);
nor U12186 (N_12186,N_10604,N_8195);
and U12187 (N_12187,N_9640,N_10766);
nand U12188 (N_12188,N_11469,N_9275);
nand U12189 (N_12189,N_8513,N_9939);
and U12190 (N_12190,N_11091,N_8528);
nor U12191 (N_12191,N_10454,N_11314);
and U12192 (N_12192,N_11665,N_11563);
xnor U12193 (N_12193,N_8900,N_11477);
nor U12194 (N_12194,N_9493,N_8811);
and U12195 (N_12195,N_10801,N_9429);
and U12196 (N_12196,N_11219,N_10319);
nand U12197 (N_12197,N_9851,N_8271);
xnor U12198 (N_12198,N_8502,N_9647);
nand U12199 (N_12199,N_9309,N_8053);
nand U12200 (N_12200,N_8770,N_11801);
or U12201 (N_12201,N_9193,N_10664);
nand U12202 (N_12202,N_9350,N_11806);
nor U12203 (N_12203,N_8298,N_8561);
and U12204 (N_12204,N_10919,N_11456);
or U12205 (N_12205,N_8669,N_10781);
xor U12206 (N_12206,N_9462,N_10089);
and U12207 (N_12207,N_9287,N_9797);
or U12208 (N_12208,N_11420,N_10355);
or U12209 (N_12209,N_9311,N_9417);
nor U12210 (N_12210,N_8012,N_9562);
nand U12211 (N_12211,N_10008,N_9565);
or U12212 (N_12212,N_9374,N_10678);
nand U12213 (N_12213,N_8937,N_11545);
xnor U12214 (N_12214,N_8718,N_9831);
and U12215 (N_12215,N_9167,N_10268);
and U12216 (N_12216,N_11057,N_11031);
nand U12217 (N_12217,N_10908,N_9319);
nand U12218 (N_12218,N_8064,N_8032);
and U12219 (N_12219,N_8901,N_8370);
nor U12220 (N_12220,N_11818,N_8060);
xor U12221 (N_12221,N_11882,N_10258);
nand U12222 (N_12222,N_10122,N_11377);
and U12223 (N_12223,N_10462,N_8870);
nand U12224 (N_12224,N_10322,N_8772);
nor U12225 (N_12225,N_10991,N_9981);
or U12226 (N_12226,N_9294,N_9702);
xor U12227 (N_12227,N_10461,N_10427);
and U12228 (N_12228,N_10433,N_8992);
and U12229 (N_12229,N_10679,N_8689);
nand U12230 (N_12230,N_11492,N_10085);
nand U12231 (N_12231,N_11662,N_11318);
or U12232 (N_12232,N_8908,N_11906);
nand U12233 (N_12233,N_8014,N_8166);
nand U12234 (N_12234,N_10521,N_11661);
xnor U12235 (N_12235,N_9096,N_8923);
nand U12236 (N_12236,N_9829,N_8297);
and U12237 (N_12237,N_8793,N_10768);
or U12238 (N_12238,N_10579,N_9624);
and U12239 (N_12239,N_8389,N_10414);
nor U12240 (N_12240,N_11557,N_11762);
and U12241 (N_12241,N_11506,N_9943);
or U12242 (N_12242,N_10520,N_9370);
or U12243 (N_12243,N_10255,N_8677);
and U12244 (N_12244,N_10192,N_11412);
or U12245 (N_12245,N_10365,N_9605);
and U12246 (N_12246,N_8241,N_11405);
and U12247 (N_12247,N_8880,N_9917);
or U12248 (N_12248,N_9828,N_10107);
and U12249 (N_12249,N_9701,N_11347);
xor U12250 (N_12250,N_9970,N_11002);
or U12251 (N_12251,N_9083,N_8126);
nor U12252 (N_12252,N_8219,N_10649);
and U12253 (N_12253,N_9478,N_8996);
and U12254 (N_12254,N_11546,N_9197);
nor U12255 (N_12255,N_10037,N_9236);
or U12256 (N_12256,N_8668,N_8075);
nor U12257 (N_12257,N_9487,N_11780);
nand U12258 (N_12258,N_9026,N_8632);
nand U12259 (N_12259,N_9688,N_11410);
or U12260 (N_12260,N_9321,N_9610);
xor U12261 (N_12261,N_10569,N_10262);
nor U12262 (N_12262,N_11603,N_8265);
and U12263 (N_12263,N_8269,N_11379);
and U12264 (N_12264,N_10963,N_11698);
nor U12265 (N_12265,N_11782,N_8437);
nor U12266 (N_12266,N_11671,N_10254);
or U12267 (N_12267,N_8885,N_11173);
nor U12268 (N_12268,N_9907,N_9789);
and U12269 (N_12269,N_10309,N_9656);
nand U12270 (N_12270,N_9335,N_8920);
nor U12271 (N_12271,N_8270,N_8759);
nand U12272 (N_12272,N_10448,N_11324);
and U12273 (N_12273,N_11179,N_10748);
nand U12274 (N_12274,N_8912,N_10185);
and U12275 (N_12275,N_10542,N_11487);
nor U12276 (N_12276,N_11589,N_11065);
and U12277 (N_12277,N_11328,N_11628);
and U12278 (N_12278,N_8511,N_10269);
or U12279 (N_12279,N_10648,N_11739);
nor U12280 (N_12280,N_8919,N_8769);
xor U12281 (N_12281,N_8159,N_11015);
nand U12282 (N_12282,N_8746,N_8181);
nor U12283 (N_12283,N_9775,N_9224);
and U12284 (N_12284,N_9256,N_10743);
nor U12285 (N_12285,N_11927,N_10999);
nor U12286 (N_12286,N_10844,N_11097);
or U12287 (N_12287,N_9152,N_8129);
nor U12288 (N_12288,N_10658,N_10921);
or U12289 (N_12289,N_8569,N_11680);
and U12290 (N_12290,N_9921,N_10445);
or U12291 (N_12291,N_10446,N_9505);
nor U12292 (N_12292,N_10716,N_10241);
and U12293 (N_12293,N_8595,N_11018);
and U12294 (N_12294,N_11960,N_11802);
or U12295 (N_12295,N_8006,N_8925);
and U12296 (N_12296,N_9460,N_10633);
and U12297 (N_12297,N_9235,N_9955);
and U12298 (N_12298,N_8462,N_9628);
nand U12299 (N_12299,N_8757,N_9210);
xor U12300 (N_12300,N_9172,N_9817);
nand U12301 (N_12301,N_11997,N_11550);
nor U12302 (N_12302,N_11498,N_10501);
and U12303 (N_12303,N_10399,N_8508);
and U12304 (N_12304,N_11235,N_8537);
or U12305 (N_12305,N_11099,N_8845);
nand U12306 (N_12306,N_11216,N_10518);
or U12307 (N_12307,N_11453,N_9185);
nand U12308 (N_12308,N_10597,N_8801);
or U12309 (N_12309,N_11148,N_9573);
or U12310 (N_12310,N_10036,N_10788);
nor U12311 (N_12311,N_9894,N_11745);
nor U12312 (N_12312,N_11586,N_8095);
nor U12313 (N_12313,N_9128,N_10543);
nand U12314 (N_12314,N_8066,N_11985);
nor U12315 (N_12315,N_8640,N_9244);
or U12316 (N_12316,N_9262,N_10333);
and U12317 (N_12317,N_10546,N_8286);
xnor U12318 (N_12318,N_10611,N_10437);
or U12319 (N_12319,N_8624,N_8224);
and U12320 (N_12320,N_10870,N_10053);
or U12321 (N_12321,N_11983,N_11862);
or U12322 (N_12322,N_10953,N_11955);
xor U12323 (N_12323,N_8238,N_10983);
xor U12324 (N_12324,N_8343,N_9198);
xnor U12325 (N_12325,N_9551,N_8555);
or U12326 (N_12326,N_9024,N_10313);
nand U12327 (N_12327,N_8744,N_10169);
nor U12328 (N_12328,N_11730,N_8564);
nand U12329 (N_12329,N_8538,N_8748);
nand U12330 (N_12330,N_11679,N_8633);
xnor U12331 (N_12331,N_9937,N_11617);
xor U12332 (N_12332,N_9289,N_8884);
and U12333 (N_12333,N_8447,N_11261);
nand U12334 (N_12334,N_9738,N_8401);
or U12335 (N_12335,N_8853,N_9534);
nor U12336 (N_12336,N_8626,N_9510);
and U12337 (N_12337,N_8068,N_8897);
nand U12338 (N_12338,N_8326,N_10063);
or U12339 (N_12339,N_11084,N_8662);
xor U12340 (N_12340,N_8890,N_10463);
nand U12341 (N_12341,N_10578,N_10003);
nand U12342 (N_12342,N_11635,N_11161);
nand U12343 (N_12343,N_11989,N_8590);
and U12344 (N_12344,N_10951,N_11707);
or U12345 (N_12345,N_10957,N_10850);
and U12346 (N_12346,N_10390,N_10413);
nand U12347 (N_12347,N_9972,N_10728);
and U12348 (N_12348,N_8691,N_9156);
nor U12349 (N_12349,N_11247,N_9279);
or U12350 (N_12350,N_9132,N_8122);
or U12351 (N_12351,N_11063,N_8613);
or U12352 (N_12352,N_9316,N_11638);
nand U12353 (N_12353,N_9536,N_10420);
or U12354 (N_12354,N_10034,N_9858);
and U12355 (N_12355,N_9875,N_9589);
nand U12356 (N_12356,N_9477,N_8079);
nor U12357 (N_12357,N_10673,N_11479);
xnor U12358 (N_12358,N_11943,N_10039);
nand U12359 (N_12359,N_9303,N_10720);
or U12360 (N_12360,N_8152,N_9737);
and U12361 (N_12361,N_10704,N_11724);
or U12362 (N_12362,N_9023,N_9773);
nor U12363 (N_12363,N_8715,N_11280);
xor U12364 (N_12364,N_8099,N_10902);
or U12365 (N_12365,N_8418,N_10928);
nor U12366 (N_12366,N_8956,N_8121);
or U12367 (N_12367,N_9239,N_8587);
nor U12368 (N_12368,N_10923,N_10425);
nand U12369 (N_12369,N_11784,N_11958);
or U12370 (N_12370,N_10650,N_9414);
or U12371 (N_12371,N_9560,N_11899);
nand U12372 (N_12372,N_8158,N_10959);
and U12373 (N_12373,N_8774,N_10106);
nor U12374 (N_12374,N_8678,N_11809);
and U12375 (N_12375,N_11076,N_11337);
or U12376 (N_12376,N_10562,N_9657);
nor U12377 (N_12377,N_9598,N_8444);
xnor U12378 (N_12378,N_10789,N_9543);
or U12379 (N_12379,N_10846,N_9838);
or U12380 (N_12380,N_11928,N_9246);
or U12381 (N_12381,N_9104,N_9923);
or U12382 (N_12382,N_10857,N_8354);
and U12383 (N_12383,N_10337,N_11569);
nor U12384 (N_12384,N_10315,N_8477);
nor U12385 (N_12385,N_9087,N_8245);
nor U12386 (N_12386,N_9140,N_9134);
nor U12387 (N_12387,N_10240,N_11770);
or U12388 (N_12388,N_9208,N_11375);
or U12389 (N_12389,N_11885,N_11109);
and U12390 (N_12390,N_9045,N_11098);
nor U12391 (N_12391,N_9464,N_10297);
and U12392 (N_12392,N_8945,N_9322);
nand U12393 (N_12393,N_9799,N_11733);
nor U12394 (N_12394,N_10627,N_9847);
nand U12395 (N_12395,N_10150,N_10205);
and U12396 (N_12396,N_8328,N_9064);
and U12397 (N_12397,N_9173,N_11041);
and U12398 (N_12398,N_10084,N_11244);
or U12399 (N_12399,N_10290,N_9017);
or U12400 (N_12400,N_8509,N_11941);
xor U12401 (N_12401,N_9604,N_11092);
and U12402 (N_12402,N_9225,N_11446);
nor U12403 (N_12403,N_8601,N_9976);
and U12404 (N_12404,N_10625,N_10995);
or U12405 (N_12405,N_11517,N_9138);
and U12406 (N_12406,N_9661,N_10558);
nand U12407 (N_12407,N_9528,N_8641);
nand U12408 (N_12408,N_10212,N_11228);
and U12409 (N_12409,N_8478,N_11027);
xnor U12410 (N_12410,N_10777,N_11887);
nand U12411 (N_12411,N_10276,N_11349);
or U12412 (N_12412,N_9398,N_10363);
nor U12413 (N_12413,N_9670,N_9496);
xnor U12414 (N_12414,N_8289,N_9150);
or U12415 (N_12415,N_11156,N_11003);
or U12416 (N_12416,N_10910,N_8824);
or U12417 (N_12417,N_9304,N_8474);
nand U12418 (N_12418,N_8593,N_11089);
and U12419 (N_12419,N_11512,N_9795);
nand U12420 (N_12420,N_11898,N_11189);
nand U12421 (N_12421,N_9394,N_11987);
or U12422 (N_12422,N_11133,N_10261);
nor U12423 (N_12423,N_8118,N_9343);
and U12424 (N_12424,N_9862,N_11323);
xnor U12425 (N_12425,N_9996,N_10988);
and U12426 (N_12426,N_11599,N_11275);
nand U12427 (N_12427,N_8260,N_10932);
or U12428 (N_12428,N_10830,N_11397);
or U12429 (N_12429,N_11302,N_10431);
nor U12430 (N_12430,N_11493,N_9861);
nand U12431 (N_12431,N_9521,N_10772);
nor U12432 (N_12432,N_8093,N_9905);
nor U12433 (N_12433,N_10087,N_8797);
and U12434 (N_12434,N_9061,N_11077);
and U12435 (N_12435,N_10971,N_8335);
nand U12436 (N_12436,N_10641,N_8406);
and U12437 (N_12437,N_11759,N_9823);
xor U12438 (N_12438,N_10732,N_10582);
or U12439 (N_12439,N_9001,N_11445);
nand U12440 (N_12440,N_9344,N_9612);
nand U12441 (N_12441,N_9930,N_10278);
or U12442 (N_12442,N_9199,N_8680);
and U12443 (N_12443,N_9579,N_11953);
or U12444 (N_12444,N_9712,N_9339);
nand U12445 (N_12445,N_8517,N_10909);
nand U12446 (N_12446,N_8156,N_9544);
and U12447 (N_12447,N_8969,N_9008);
nand U12448 (N_12448,N_11583,N_9871);
or U12449 (N_12449,N_11931,N_10170);
and U12450 (N_12450,N_10080,N_11540);
and U12451 (N_12451,N_9472,N_9479);
and U12452 (N_12452,N_11267,N_9678);
nand U12453 (N_12453,N_10888,N_9979);
and U12454 (N_12454,N_8130,N_10128);
xnor U12455 (N_12455,N_11805,N_10097);
nor U12456 (N_12456,N_11744,N_11028);
or U12457 (N_12457,N_9704,N_10306);
and U12458 (N_12458,N_9574,N_10807);
or U12459 (N_12459,N_9853,N_8592);
nor U12460 (N_12460,N_8507,N_8637);
xor U12461 (N_12461,N_9732,N_9808);
and U12462 (N_12462,N_9361,N_11436);
nor U12463 (N_12463,N_8239,N_9735);
or U12464 (N_12464,N_10616,N_8621);
and U12465 (N_12465,N_11081,N_8922);
or U12466 (N_12466,N_11153,N_8021);
nor U12467 (N_12467,N_11340,N_9860);
or U12468 (N_12468,N_11214,N_10836);
nor U12469 (N_12469,N_8927,N_9461);
or U12470 (N_12470,N_11585,N_8781);
or U12471 (N_12471,N_10473,N_8023);
or U12472 (N_12472,N_9115,N_8430);
nor U12473 (N_12473,N_9163,N_9100);
or U12474 (N_12474,N_11536,N_10554);
nand U12475 (N_12475,N_11310,N_9268);
or U12476 (N_12476,N_10670,N_8028);
nor U12477 (N_12477,N_9741,N_11345);
nand U12478 (N_12478,N_10342,N_9845);
or U12479 (N_12479,N_10581,N_9836);
nand U12480 (N_12480,N_8972,N_11306);
nand U12481 (N_12481,N_11685,N_8411);
or U12482 (N_12482,N_9047,N_10402);
and U12483 (N_12483,N_9591,N_9506);
and U12484 (N_12484,N_8109,N_9255);
nand U12485 (N_12485,N_8388,N_10256);
and U12486 (N_12486,N_10283,N_9397);
xnor U12487 (N_12487,N_11946,N_9569);
or U12488 (N_12488,N_9934,N_11562);
and U12489 (N_12489,N_8931,N_9248);
nand U12490 (N_12490,N_8938,N_9031);
xor U12491 (N_12491,N_9600,N_11115);
nand U12492 (N_12492,N_8552,N_10186);
nor U12493 (N_12493,N_8739,N_8142);
nand U12494 (N_12494,N_10539,N_10102);
nor U12495 (N_12495,N_11535,N_11718);
nor U12496 (N_12496,N_10472,N_8864);
and U12497 (N_12497,N_10249,N_8791);
nor U12498 (N_12498,N_9125,N_9118);
and U12499 (N_12499,N_11573,N_9044);
nor U12500 (N_12500,N_8775,N_8723);
xnor U12501 (N_12501,N_10061,N_8000);
nand U12502 (N_12502,N_10528,N_10385);
nor U12503 (N_12503,N_11804,N_9998);
or U12504 (N_12504,N_11012,N_9390);
or U12505 (N_12505,N_9613,N_11390);
xnor U12506 (N_12506,N_8918,N_9575);
and U12507 (N_12507,N_11771,N_11154);
nor U12508 (N_12508,N_9874,N_10394);
xnor U12509 (N_12509,N_11342,N_9523);
xnor U12510 (N_12510,N_11765,N_11243);
nand U12511 (N_12511,N_8796,N_11248);
nor U12512 (N_12512,N_9145,N_8300);
nor U12513 (N_12513,N_10140,N_11268);
xnor U12514 (N_12514,N_11640,N_11304);
xor U12515 (N_12515,N_11167,N_11525);
xnor U12516 (N_12516,N_10806,N_9620);
nand U12517 (N_12517,N_10565,N_10040);
nor U12518 (N_12518,N_8727,N_9230);
nor U12519 (N_12519,N_10813,N_10271);
nand U12520 (N_12520,N_10044,N_10175);
nand U12521 (N_12521,N_9091,N_8661);
nand U12522 (N_12522,N_10688,N_9404);
or U12523 (N_12523,N_10114,N_11067);
nand U12524 (N_12524,N_9086,N_9771);
nand U12525 (N_12525,N_11991,N_8644);
nand U12526 (N_12526,N_8380,N_11604);
nor U12527 (N_12527,N_8971,N_11523);
or U12528 (N_12528,N_8510,N_8877);
nand U12529 (N_12529,N_11969,N_8230);
and U12530 (N_12530,N_11623,N_9703);
and U12531 (N_12531,N_11697,N_11449);
and U12532 (N_12532,N_9237,N_8261);
nand U12533 (N_12533,N_11786,N_11203);
nand U12534 (N_12534,N_10395,N_11692);
and U12535 (N_12535,N_9722,N_11910);
nor U12536 (N_12536,N_10288,N_11435);
and U12537 (N_12537,N_11774,N_10396);
nor U12538 (N_12538,N_8650,N_9896);
nand U12539 (N_12539,N_10368,N_11826);
xor U12540 (N_12540,N_11865,N_10904);
xor U12541 (N_12541,N_11008,N_11933);
nand U12542 (N_12542,N_10126,N_11262);
nand U12543 (N_12543,N_8934,N_11502);
or U12544 (N_12544,N_8518,N_11670);
nor U12545 (N_12545,N_9405,N_8606);
nand U12546 (N_12546,N_10852,N_10364);
and U12547 (N_12547,N_10404,N_11594);
or U12548 (N_12548,N_9920,N_9476);
nor U12549 (N_12549,N_10873,N_10819);
or U12550 (N_12550,N_10467,N_8685);
nor U12551 (N_12551,N_11966,N_11396);
nand U12552 (N_12552,N_10477,N_11641);
xor U12553 (N_12553,N_8361,N_10490);
nor U12554 (N_12554,N_8596,N_8352);
xnor U12555 (N_12555,N_8169,N_9490);
nand U12556 (N_12556,N_8110,N_10314);
xor U12557 (N_12557,N_8657,N_11221);
nand U12558 (N_12558,N_10451,N_11889);
and U12559 (N_12559,N_11597,N_11674);
or U12560 (N_12560,N_9919,N_11767);
or U12561 (N_12561,N_11821,N_10636);
xnor U12562 (N_12562,N_9806,N_8840);
xnor U12563 (N_12563,N_9975,N_9359);
nand U12564 (N_12564,N_9577,N_9112);
nor U12565 (N_12565,N_8725,N_11439);
nor U12566 (N_12566,N_8420,N_9774);
nand U12567 (N_12567,N_10556,N_9649);
and U12568 (N_12568,N_8227,N_11281);
nand U12569 (N_12569,N_8194,N_8960);
xor U12570 (N_12570,N_11678,N_11505);
nand U12571 (N_12571,N_11852,N_10432);
or U12572 (N_12572,N_11352,N_11769);
nand U12573 (N_12573,N_11791,N_8225);
nor U12574 (N_12574,N_8903,N_11136);
nand U12575 (N_12575,N_8107,N_10973);
or U12576 (N_12576,N_11491,N_11677);
nor U12577 (N_12577,N_11117,N_8315);
nand U12578 (N_12578,N_9337,N_8754);
or U12579 (N_12579,N_8985,N_10350);
or U12580 (N_12580,N_9819,N_10330);
or U12581 (N_12581,N_11182,N_11011);
or U12582 (N_12582,N_10568,N_9352);
or U12583 (N_12583,N_11532,N_10219);
and U12584 (N_12584,N_8174,N_8008);
nand U12585 (N_12585,N_11462,N_10802);
or U12586 (N_12586,N_8728,N_10596);
xnor U12587 (N_12587,N_9297,N_11311);
nor U12588 (N_12588,N_11030,N_10042);
nand U12589 (N_12589,N_9884,N_11624);
and U12590 (N_12590,N_11432,N_8961);
xnor U12591 (N_12591,N_8134,N_10864);
or U12592 (N_12592,N_8385,N_10922);
and U12593 (N_12593,N_11757,N_10302);
nand U12594 (N_12594,N_8716,N_11100);
nand U12595 (N_12595,N_8321,N_8586);
and U12596 (N_12596,N_8402,N_8011);
nor U12597 (N_12597,N_9902,N_11144);
nor U12598 (N_12598,N_8184,N_11424);
or U12599 (N_12599,N_9618,N_10747);
nand U12600 (N_12600,N_8133,N_8287);
xnor U12601 (N_12601,N_11970,N_10282);
nand U12602 (N_12602,N_10550,N_10035);
and U12603 (N_12603,N_10028,N_10294);
nand U12604 (N_12604,N_8256,N_9985);
and U12605 (N_12605,N_9284,N_9068);
and U12606 (N_12606,N_10164,N_11591);
xor U12607 (N_12607,N_8396,N_8916);
nor U12608 (N_12608,N_11124,N_10936);
and U12609 (N_12609,N_10729,N_8558);
xnor U12610 (N_12610,N_11963,N_9938);
or U12611 (N_12611,N_10702,N_9314);
and U12612 (N_12612,N_9906,N_10157);
nand U12613 (N_12613,N_8879,N_9426);
nor U12614 (N_12614,N_9572,N_10719);
and U12615 (N_12615,N_11870,N_10619);
and U12616 (N_12616,N_8196,N_11949);
and U12617 (N_12617,N_11849,N_8849);
nand U12618 (N_12618,N_10341,N_11355);
nand U12619 (N_12619,N_8583,N_10527);
or U12620 (N_12620,N_8976,N_11807);
xnor U12621 (N_12621,N_8600,N_8675);
nand U12622 (N_12622,N_8591,N_10529);
xnor U12623 (N_12623,N_8799,N_8108);
nor U12624 (N_12624,N_9502,N_9527);
nand U12625 (N_12625,N_8489,N_9727);
or U12626 (N_12626,N_10064,N_11122);
or U12627 (N_12627,N_11217,N_10016);
nor U12628 (N_12628,N_11331,N_10586);
xnor U12629 (N_12629,N_9877,N_9707);
nor U12630 (N_12630,N_9548,N_11858);
or U12631 (N_12631,N_10489,N_9922);
nor U12632 (N_12632,N_11042,N_11068);
nor U12633 (N_12633,N_9837,N_8494);
and U12634 (N_12634,N_10764,N_11593);
nor U12635 (N_12635,N_9728,N_11929);
and U12636 (N_12636,N_8198,N_10438);
nor U12637 (N_12637,N_10194,N_9219);
or U12638 (N_12638,N_10523,N_10310);
or U12639 (N_12639,N_11007,N_11962);
or U12640 (N_12640,N_8898,N_10148);
nor U12641 (N_12641,N_9665,N_11211);
nor U12642 (N_12642,N_9504,N_10885);
or U12643 (N_12643,N_11110,N_10939);
nand U12644 (N_12644,N_10228,N_8186);
nor U12645 (N_12645,N_8425,N_11684);
nand U12646 (N_12646,N_8773,N_10590);
nand U12647 (N_12647,N_9108,N_9857);
nand U12648 (N_12648,N_11206,N_8762);
and U12649 (N_12649,N_10099,N_11868);
nand U12650 (N_12650,N_10805,N_8819);
nand U12651 (N_12651,N_8896,N_10436);
or U12652 (N_12652,N_9048,N_11440);
and U12653 (N_12653,N_11317,N_8783);
and U12654 (N_12654,N_8472,N_8692);
xor U12655 (N_12655,N_8123,N_10361);
nor U12656 (N_12656,N_10895,N_10151);
and U12657 (N_12657,N_11087,N_9662);
nand U12658 (N_12658,N_9825,N_11534);
nor U12659 (N_12659,N_8594,N_9468);
nor U12660 (N_12660,N_9679,N_9015);
nand U12661 (N_12661,N_9341,N_11066);
nand U12662 (N_12662,N_11325,N_9331);
nand U12663 (N_12663,N_10858,N_8454);
xor U12664 (N_12664,N_8374,N_11297);
or U12665 (N_12665,N_10632,N_10767);
or U12666 (N_12666,N_8519,N_8975);
nor U12667 (N_12667,N_9009,N_11168);
nor U12668 (N_12668,N_9557,N_8292);
nor U12669 (N_12669,N_10123,N_9883);
nor U12670 (N_12670,N_10311,N_8568);
and U12671 (N_12671,N_9158,N_10841);
nor U12672 (N_12672,N_10911,N_8616);
nor U12673 (N_12673,N_9346,N_10145);
and U12674 (N_12674,N_9298,N_8247);
nand U12675 (N_12675,N_10101,N_11233);
nor U12676 (N_12676,N_8325,N_11488);
xnor U12677 (N_12677,N_11812,N_11329);
nand U12678 (N_12678,N_9820,N_8235);
nand U12679 (N_12679,N_10407,N_8794);
nand U12680 (N_12680,N_10471,N_11316);
and U12681 (N_12681,N_8035,N_8612);
nor U12682 (N_12682,N_11196,N_10000);
or U12683 (N_12683,N_11719,N_9074);
nand U12684 (N_12684,N_8554,N_9277);
nor U12685 (N_12685,N_8426,N_8242);
nand U12686 (N_12686,N_8155,N_8722);
nor U12687 (N_12687,N_9099,N_9899);
nand U12688 (N_12688,N_8428,N_8069);
and U12689 (N_12689,N_8067,N_9482);
nand U12690 (N_12690,N_8666,N_10624);
and U12691 (N_12691,N_11796,N_10639);
or U12692 (N_12692,N_9285,N_11052);
nor U12693 (N_12693,N_9597,N_8455);
nor U12694 (N_12694,N_11330,N_9873);
nand U12695 (N_12695,N_9079,N_9379);
or U12696 (N_12696,N_10450,N_10235);
or U12697 (N_12697,N_9340,N_8019);
nand U12698 (N_12698,N_8145,N_9622);
nor U12699 (N_12699,N_9078,N_10001);
xor U12700 (N_12700,N_10524,N_11129);
nand U12701 (N_12701,N_11714,N_11315);
nor U12702 (N_12702,N_10326,N_11263);
nor U12703 (N_12703,N_8795,N_10726);
or U12704 (N_12704,N_9056,N_8404);
or U12705 (N_12705,N_10642,N_8400);
or U12706 (N_12706,N_9320,N_11705);
and U12707 (N_12707,N_8565,N_10149);
or U12708 (N_12708,N_11171,N_8828);
nand U12709 (N_12709,N_9957,N_10575);
or U12710 (N_12710,N_9222,N_10045);
nand U12711 (N_12711,N_8193,N_11164);
and U12712 (N_12712,N_9280,N_9067);
and U12713 (N_12713,N_11972,N_10257);
nor U12714 (N_12714,N_11819,N_11504);
nor U12715 (N_12715,N_8482,N_9136);
and U12716 (N_12716,N_10945,N_8752);
and U12717 (N_12717,N_11202,N_10986);
nand U12718 (N_12718,N_10116,N_10680);
nor U12719 (N_12719,N_9174,N_11241);
or U12720 (N_12720,N_9673,N_8345);
or U12721 (N_12721,N_9456,N_8415);
or U12722 (N_12722,N_10465,N_11470);
or U12723 (N_12723,N_8676,N_11897);
or U12724 (N_12724,N_8382,N_9787);
or U12725 (N_12725,N_9481,N_8475);
xor U12726 (N_12726,N_9513,N_11040);
nand U12727 (N_12727,N_11014,N_10890);
and U12728 (N_12728,N_10487,N_9977);
or U12729 (N_12729,N_8378,N_10695);
nand U12730 (N_12730,N_11693,N_8434);
and U12731 (N_12731,N_9681,N_11378);
and U12732 (N_12732,N_8372,N_9676);
nor U12733 (N_12733,N_8205,N_11061);
nand U12734 (N_12734,N_9733,N_10357);
or U12735 (N_12735,N_10937,N_9537);
nor U12736 (N_12736,N_11155,N_8316);
or U12737 (N_12737,N_11231,N_8116);
and U12738 (N_12738,N_10623,N_10903);
nor U12739 (N_12739,N_11509,N_10849);
and U12740 (N_12740,N_8257,N_8233);
xor U12741 (N_12741,N_10180,N_9012);
or U12742 (N_12742,N_11215,N_9660);
or U12743 (N_12743,N_10900,N_8450);
or U12744 (N_12744,N_9731,N_9123);
xnor U12745 (N_12745,N_10092,N_9301);
nand U12746 (N_12746,N_8146,N_10832);
or U12747 (N_12747,N_9803,N_9967);
or U12748 (N_12748,N_9849,N_11073);
nand U12749 (N_12749,N_10112,N_9990);
xnor U12750 (N_12750,N_8501,N_11614);
nor U12751 (N_12751,N_9006,N_9432);
or U12752 (N_12752,N_8377,N_11021);
nor U12753 (N_12753,N_11853,N_10020);
nand U12754 (N_12754,N_10202,N_9492);
nor U12755 (N_12755,N_10245,N_11494);
and U12756 (N_12756,N_8049,N_11876);
and U12757 (N_12757,N_8882,N_9153);
or U12758 (N_12758,N_10701,N_8814);
nand U12759 (N_12759,N_10449,N_8317);
and U12760 (N_12760,N_10750,N_8914);
or U12761 (N_12761,N_9770,N_9036);
nor U12762 (N_12762,N_11086,N_11764);
or U12763 (N_12763,N_11609,N_11060);
nor U12764 (N_12764,N_10981,N_11135);
or U12765 (N_12765,N_8337,N_11704);
or U12766 (N_12766,N_11053,N_8579);
or U12767 (N_12767,N_10203,N_9987);
nor U12768 (N_12768,N_8547,N_8539);
nor U12769 (N_12769,N_11631,N_8826);
nor U12770 (N_12770,N_11923,N_10567);
and U12771 (N_12771,N_11967,N_8304);
and U12772 (N_12772,N_8605,N_8203);
and U12773 (N_12773,N_9793,N_9470);
and U12774 (N_12774,N_9962,N_9687);
nand U12775 (N_12775,N_10593,N_10880);
or U12776 (N_12776,N_11111,N_11074);
nand U12777 (N_12777,N_9376,N_8854);
nor U12778 (N_12778,N_9925,N_9192);
or U12779 (N_12779,N_11803,N_8039);
nor U12780 (N_12780,N_11134,N_9995);
nor U12781 (N_12781,N_8137,N_9076);
and U12782 (N_12782,N_11118,N_10775);
nor U12783 (N_12783,N_8815,N_9391);
nor U12784 (N_12784,N_9447,N_10771);
nand U12785 (N_12785,N_8563,N_10935);
or U12786 (N_12786,N_8139,N_11472);
or U12787 (N_12787,N_8128,N_10862);
nor U12788 (N_12788,N_10686,N_9201);
xnor U12789 (N_12789,N_11867,N_11924);
nand U12790 (N_12790,N_9360,N_10082);
or U12791 (N_12791,N_8293,N_8005);
or U12792 (N_12792,N_11551,N_11398);
and U12793 (N_12793,N_11106,N_10744);
or U12794 (N_12794,N_9872,N_8670);
nor U12795 (N_12795,N_9296,N_11590);
xor U12796 (N_12796,N_8362,N_9585);
and U12797 (N_12797,N_9720,N_8311);
or U12798 (N_12798,N_11696,N_11956);
nor U12799 (N_12799,N_11475,N_10886);
nor U12800 (N_12800,N_8197,N_11957);
nand U12801 (N_12801,N_10386,N_9900);
or U12802 (N_12802,N_11779,N_8785);
and U12803 (N_12803,N_11418,N_11365);
nor U12804 (N_12804,N_10759,N_8868);
nor U12805 (N_12805,N_9674,N_11308);
nand U12806 (N_12806,N_8483,N_8386);
and U12807 (N_12807,N_11503,N_9127);
or U12808 (N_12808,N_9956,N_10735);
or U12809 (N_12809,N_9430,N_10866);
or U12810 (N_12810,N_10351,N_10834);
nor U12811 (N_12811,N_11177,N_8738);
or U12812 (N_12812,N_9541,N_8946);
xnor U12813 (N_12813,N_9403,N_10577);
and U12814 (N_12814,N_11335,N_11713);
or U12815 (N_12815,N_10174,N_11560);
nor U12816 (N_12816,N_9042,N_8448);
nor U12817 (N_12817,N_11457,N_8414);
nand U12818 (N_12818,N_8303,N_11636);
nor U12819 (N_12819,N_10693,N_9446);
and U12820 (N_12820,N_11709,N_11723);
nor U12821 (N_12821,N_10815,N_11766);
nor U12822 (N_12822,N_9554,N_11113);
nor U12823 (N_12823,N_10843,N_9913);
or U12824 (N_12824,N_10799,N_8278);
or U12825 (N_12825,N_8185,N_10495);
or U12826 (N_12826,N_10204,N_11184);
or U12827 (N_12827,N_8761,N_11448);
and U12828 (N_12828,N_10757,N_10430);
xnor U12829 (N_12829,N_8250,N_8443);
nand U12830 (N_12830,N_8891,N_8439);
nor U12831 (N_12831,N_8610,N_8698);
or U12832 (N_12832,N_10098,N_10109);
xor U12833 (N_12833,N_8506,N_10065);
and U12834 (N_12834,N_11515,N_10452);
nand U12835 (N_12835,N_9334,N_10948);
nand U12836 (N_12836,N_8549,N_8369);
nand U12837 (N_12837,N_9615,N_11307);
and U12838 (N_12838,N_8074,N_11285);
or U12839 (N_12839,N_11200,N_11464);
xor U12840 (N_12840,N_10711,N_8484);
or U12841 (N_12841,N_9954,N_8812);
xnor U12842 (N_12842,N_8705,N_10054);
nand U12843 (N_12843,N_8572,N_11431);
or U12844 (N_12844,N_11841,N_9992);
and U12845 (N_12845,N_8878,N_8798);
nor U12846 (N_12846,N_8098,N_11790);
nand U12847 (N_12847,N_8243,N_8465);
or U12848 (N_12848,N_10141,N_11139);
or U12849 (N_12849,N_10733,N_8324);
nand U12850 (N_12850,N_10804,N_8742);
or U12851 (N_12851,N_10931,N_10217);
and U12852 (N_12852,N_9651,N_10793);
xor U12853 (N_12853,N_11715,N_9375);
or U12854 (N_12854,N_8917,N_9328);
or U12855 (N_12855,N_11754,N_11646);
xor U12856 (N_12856,N_9055,N_8629);
nor U12857 (N_12857,N_11911,N_8700);
and U12858 (N_12858,N_8038,N_8210);
xnor U12859 (N_12859,N_8082,N_10181);
or U12860 (N_12860,N_11283,N_8982);
xnor U12861 (N_12861,N_8217,N_10177);
or U12862 (N_12862,N_10871,N_8979);
nand U12863 (N_12863,N_9085,N_11903);
and U12864 (N_12864,N_10198,N_8872);
nand U12865 (N_12865,N_9040,N_8530);
nor U12866 (N_12866,N_10195,N_8161);
or U12867 (N_12867,N_8077,N_10331);
or U12868 (N_12868,N_10893,N_8526);
and U12869 (N_12869,N_9555,N_8704);
nand U12870 (N_12870,N_9846,N_8763);
and U12871 (N_12871,N_11341,N_9387);
nor U12872 (N_12872,N_10826,N_10440);
nand U12873 (N_12873,N_8267,N_11291);
or U12874 (N_12874,N_8431,N_8907);
nand U12875 (N_12875,N_11121,N_11357);
nand U12876 (N_12876,N_8832,N_9148);
and U12877 (N_12877,N_8803,N_9559);
nand U12878 (N_12878,N_9441,N_8207);
nor U12879 (N_12879,N_10172,N_10412);
nand U12880 (N_12880,N_11195,N_11039);
or U12881 (N_12881,N_9503,N_11810);
and U12882 (N_12882,N_8782,N_9764);
nor U12883 (N_12883,N_9194,N_10965);
xor U12884 (N_12884,N_9336,N_8962);
or U12885 (N_12885,N_10725,N_10485);
or U12886 (N_12886,N_10470,N_11128);
nand U12887 (N_12887,N_9168,N_9614);
nor U12888 (N_12888,N_8611,N_8228);
or U12889 (N_12889,N_9594,N_10952);
nor U12890 (N_12890,N_11169,N_9550);
and U12891 (N_12891,N_9037,N_11409);
nor U12892 (N_12892,N_8807,N_10925);
nand U12893 (N_12893,N_9353,N_11427);
and U12894 (N_12894,N_11392,N_11829);
and U12895 (N_12895,N_11939,N_10316);
or U12896 (N_12896,N_9736,N_11372);
and U12897 (N_12897,N_11274,N_9105);
or U12898 (N_12898,N_11763,N_8280);
xor U12899 (N_12899,N_10071,N_10734);
or U12900 (N_12900,N_8859,N_9362);
and U12901 (N_12901,N_8062,N_11572);
nor U12902 (N_12902,N_8756,N_10924);
and U12903 (N_12903,N_11596,N_11468);
nand U12904 (N_12904,N_10814,N_11374);
and U12905 (N_12905,N_9418,N_8451);
and U12906 (N_12906,N_10086,N_8200);
and U12907 (N_12907,N_9744,N_11484);
or U12908 (N_12908,N_10416,N_11478);
nor U12909 (N_12909,N_8338,N_11874);
nand U12910 (N_12910,N_9165,N_11598);
or U12911 (N_12911,N_10920,N_8699);
nand U12912 (N_12912,N_9552,N_8153);
or U12913 (N_12913,N_8684,N_10421);
and U12914 (N_12914,N_10754,N_9864);
nand U12915 (N_12915,N_11847,N_10713);
nor U12916 (N_12916,N_9603,N_11104);
nor U12917 (N_12917,N_11059,N_9982);
nand U12918 (N_12918,N_9436,N_8604);
nor U12919 (N_12919,N_9454,N_8983);
nand U12920 (N_12920,N_9854,N_11556);
nor U12921 (N_12921,N_9435,N_11312);
xor U12922 (N_12922,N_8866,N_9519);
nand U12923 (N_12923,N_11046,N_10517);
nand U12924 (N_12924,N_9019,N_10124);
or U12925 (N_12925,N_9750,N_11675);
and U12926 (N_12926,N_9276,N_9950);
nor U12927 (N_12927,N_11666,N_8874);
and U12928 (N_12928,N_11032,N_9119);
and U12929 (N_12929,N_8307,N_8745);
and U12930 (N_12930,N_10602,N_9821);
nor U12931 (N_12931,N_10332,N_11592);
or U12932 (N_12932,N_10560,N_8709);
nor U12933 (N_12933,N_11185,N_8342);
nor U12934 (N_12934,N_11150,N_8351);
xor U12935 (N_12935,N_8743,N_11326);
and U12936 (N_12936,N_10975,N_11454);
nand U12937 (N_12937,N_9881,N_8800);
and U12938 (N_12938,N_9177,N_10329);
and U12939 (N_12939,N_11276,N_10004);
nor U12940 (N_12940,N_10669,N_10601);
nor U12941 (N_12941,N_8112,N_9188);
nand U12942 (N_12942,N_8440,N_11165);
nand U12943 (N_12943,N_8703,N_11524);
nand U12944 (N_12944,N_11152,N_9355);
nor U12945 (N_12945,N_8391,N_8026);
and U12946 (N_12946,N_11237,N_8364);
xor U12947 (N_12947,N_9973,N_10488);
or U12948 (N_12948,N_9200,N_8486);
nor U12949 (N_12949,N_9223,N_8602);
and U12950 (N_12950,N_10640,N_10362);
and U12951 (N_12951,N_8111,N_10152);
nor U12952 (N_12952,N_9832,N_8306);
nand U12953 (N_12953,N_9323,N_8277);
and U12954 (N_12954,N_9189,N_8575);
and U12955 (N_12955,N_8091,N_8964);
nand U12956 (N_12956,N_11907,N_8886);
or U12957 (N_12957,N_9677,N_8567);
and U12958 (N_12958,N_10051,N_11455);
and U12959 (N_12959,N_8576,N_8627);
and U12960 (N_12960,N_11712,N_11799);
nand U12961 (N_12961,N_10024,N_8994);
nor U12962 (N_12962,N_10435,N_11450);
and U12963 (N_12963,N_9229,N_11078);
nand U12964 (N_12964,N_9269,N_10095);
xnor U12965 (N_12965,N_8379,N_8266);
nand U12966 (N_12966,N_10179,N_8163);
nor U12967 (N_12967,N_11417,N_8344);
nand U12968 (N_12968,N_10030,N_11406);
and U12969 (N_12969,N_10631,N_8686);
nand U12970 (N_12970,N_10595,N_8737);
and U12971 (N_12971,N_11857,N_9745);
xor U12972 (N_12972,N_9263,N_8468);
nor U12973 (N_12973,N_11553,N_11541);
nor U12974 (N_12974,N_8822,N_9693);
or U12975 (N_12975,N_10672,N_9354);
and U12976 (N_12976,N_10842,N_8030);
nand U12977 (N_12977,N_9581,N_11389);
nand U12978 (N_12978,N_9166,N_11499);
nor U12979 (N_12979,N_9988,N_8376);
nor U12980 (N_12980,N_8258,N_11344);
or U12981 (N_12981,N_10727,N_10837);
and U12982 (N_12982,N_11751,N_8092);
and U12983 (N_12983,N_9684,N_10745);
and U12984 (N_12984,N_11752,N_10792);
and U12985 (N_12985,N_8957,N_11851);
nor U12986 (N_12986,N_11606,N_9306);
or U12987 (N_12987,N_10656,N_11029);
or U12988 (N_12988,N_9608,N_10960);
or U12989 (N_12989,N_10809,N_8952);
or U12990 (N_12990,N_11204,N_10566);
or U12991 (N_12991,N_9348,N_9221);
and U12992 (N_12992,N_8978,N_11668);
nand U12993 (N_12993,N_9984,N_10484);
xor U12994 (N_12994,N_11403,N_11973);
nor U12995 (N_12995,N_8357,N_8221);
nor U12996 (N_12996,N_10409,N_11746);
xnor U12997 (N_12997,N_10060,N_10753);
and U12998 (N_12998,N_9095,N_11825);
and U12999 (N_12999,N_11778,N_9824);
and U13000 (N_13000,N_8170,N_10216);
nor U13001 (N_13001,N_11878,N_9946);
and U13002 (N_13002,N_8690,N_8220);
nor U13003 (N_13003,N_8423,N_9409);
nand U13004 (N_13004,N_11434,N_8977);
xor U13005 (N_13005,N_9699,N_8639);
nor U13006 (N_13006,N_11295,N_9959);
and U13007 (N_13007,N_9964,N_9072);
or U13008 (N_13008,N_10927,N_9195);
nor U13009 (N_13009,N_10048,N_10692);
and U13010 (N_13010,N_8648,N_8693);
and U13011 (N_13011,N_8660,N_8176);
nand U13012 (N_13012,N_10868,N_10993);
nand U13013 (N_13013,N_11529,N_10774);
nand U13014 (N_13014,N_9752,N_8149);
nor U13015 (N_13015,N_8063,N_11413);
and U13016 (N_13016,N_10091,N_8664);
nand U13017 (N_13017,N_9090,N_9742);
nand U13018 (N_13018,N_8999,N_10166);
nand U13019 (N_13019,N_8365,N_9106);
nor U13020 (N_13020,N_11612,N_9928);
nor U13021 (N_13021,N_9433,N_9634);
nand U13022 (N_13022,N_9448,N_8679);
and U13023 (N_13023,N_8747,N_10119);
and U13024 (N_13024,N_10171,N_8835);
nand U13025 (N_13025,N_9754,N_11986);
or U13026 (N_13026,N_8570,N_9474);
nand U13027 (N_13027,N_11735,N_11669);
nand U13028 (N_13028,N_8818,N_8932);
or U13029 (N_13029,N_10072,N_9029);
xor U13030 (N_13030,N_10803,N_9259);
or U13031 (N_13031,N_8407,N_9184);
and U13032 (N_13032,N_11672,N_10324);
nand U13033 (N_13033,N_9867,N_9077);
or U13034 (N_13034,N_9131,N_9212);
xor U13035 (N_13035,N_8881,N_10913);
nand U13036 (N_13036,N_10453,N_8860);
xnor U13037 (N_13037,N_11366,N_9520);
xor U13038 (N_13038,N_11026,N_11965);
and U13039 (N_13039,N_10023,N_9310);
and U13040 (N_13040,N_11690,N_9114);
nand U13041 (N_13041,N_9473,N_10137);
and U13042 (N_13042,N_10223,N_8131);
xor U13043 (N_13043,N_9160,N_10574);
xor U13044 (N_13044,N_8481,N_8456);
nor U13045 (N_13045,N_8778,N_11292);
and U13046 (N_13046,N_9895,N_10275);
nor U13047 (N_13047,N_9659,N_10117);
and U13048 (N_13048,N_8138,N_10160);
nand U13049 (N_13049,N_10077,N_10950);
nor U13050 (N_13050,N_9272,N_10591);
nor U13051 (N_13051,N_10861,N_8147);
nor U13052 (N_13052,N_8719,N_9103);
nand U13053 (N_13053,N_8764,N_8065);
nand U13054 (N_13054,N_9129,N_8463);
or U13055 (N_13055,N_8941,N_9180);
and U13056 (N_13056,N_9209,N_10088);
xnor U13057 (N_13057,N_9705,N_8562);
or U13058 (N_13058,N_9142,N_10698);
and U13059 (N_13059,N_9288,N_11575);
or U13060 (N_13060,N_11447,N_9570);
or U13061 (N_13061,N_9422,N_11998);
nand U13062 (N_13062,N_10589,N_11846);
nor U13063 (N_13063,N_9018,N_10377);
nand U13064 (N_13064,N_10382,N_8308);
nand U13065 (N_13065,N_10668,N_11564);
nor U13066 (N_13066,N_11514,N_8873);
or U13067 (N_13067,N_11313,N_11788);
nor U13068 (N_13068,N_11266,N_11201);
and U13069 (N_13069,N_10723,N_9332);
nand U13070 (N_13070,N_10621,N_10422);
and U13071 (N_13071,N_8713,N_9383);
or U13072 (N_13072,N_8371,N_11561);
and U13073 (N_13073,N_11915,N_8500);
nor U13074 (N_13074,N_8027,N_10645);
nor U13075 (N_13075,N_9926,N_8542);
nor U13076 (N_13076,N_8272,N_8910);
and U13077 (N_13077,N_11643,N_11510);
nor U13078 (N_13078,N_9203,N_10424);
and U13079 (N_13079,N_9389,N_10244);
nor U13080 (N_13080,N_10784,N_11269);
nand U13081 (N_13081,N_9859,N_10296);
nand U13082 (N_13082,N_8089,N_10388);
or U13083 (N_13083,N_9644,N_9547);
nand U13084 (N_13084,N_8585,N_10682);
nand U13085 (N_13085,N_11729,N_8167);
or U13086 (N_13086,N_11149,N_11755);
nor U13087 (N_13087,N_10652,N_9739);
xnor U13088 (N_13088,N_9252,N_10387);
and U13089 (N_13089,N_11338,N_9813);
nor U13090 (N_13090,N_10214,N_11683);
or U13091 (N_13091,N_11652,N_11119);
or U13092 (N_13092,N_10323,N_10557);
nand U13093 (N_13093,N_11495,N_9117);
and U13094 (N_13094,N_10383,N_10544);
xnor U13095 (N_13095,N_11288,N_10563);
nand U13096 (N_13096,N_10442,N_10794);
nand U13097 (N_13097,N_9629,N_11146);
and U13098 (N_13098,N_10994,N_9929);
nand U13099 (N_13099,N_8294,N_10155);
and U13100 (N_13100,N_11798,N_10962);
or U13101 (N_13101,N_9843,N_8199);
or U13102 (N_13102,N_11384,N_9983);
and U13103 (N_13103,N_9013,N_10287);
or U13104 (N_13104,N_10354,N_11108);
and U13105 (N_13105,N_9522,N_9242);
nor U13106 (N_13106,N_9516,N_9333);
nor U13107 (N_13107,N_10511,N_9692);
nand U13108 (N_13108,N_10778,N_10393);
nand U13109 (N_13109,N_8531,N_10005);
nor U13110 (N_13110,N_10374,N_11695);
or U13111 (N_13111,N_11916,N_8061);
nand U13112 (N_13112,N_8953,N_9625);
and U13113 (N_13113,N_10827,N_11836);
and U13114 (N_13114,N_8805,N_8836);
or U13115 (N_13115,N_11380,N_11656);
nor U13116 (N_13116,N_10018,N_8201);
xnor U13117 (N_13117,N_10073,N_9302);
and U13118 (N_13118,N_9653,N_9075);
nor U13119 (N_13119,N_9458,N_11388);
nand U13120 (N_13120,N_11010,N_10676);
nor U13121 (N_13121,N_10279,N_8720);
and U13122 (N_13122,N_10982,N_9642);
and U13123 (N_13123,N_9762,N_9993);
nor U13124 (N_13124,N_8143,N_8329);
nand U13125 (N_13125,N_11250,N_11945);
or U13126 (N_13126,N_11577,N_8119);
or U13127 (N_13127,N_9440,N_8522);
nor U13128 (N_13128,N_8218,N_10344);
nor U13129 (N_13129,N_10818,N_10942);
or U13130 (N_13130,N_11837,N_9110);
nor U13131 (N_13131,N_9809,N_9500);
xor U13132 (N_13132,N_8788,N_11050);
nand U13133 (N_13133,N_8262,N_8658);
xnor U13134 (N_13134,N_9082,N_8802);
nand U13135 (N_13135,N_10055,N_9161);
nand U13136 (N_13136,N_11253,N_11284);
and U13137 (N_13137,N_11320,N_8397);
nand U13138 (N_13138,N_9812,N_11855);
nand U13139 (N_13139,N_11935,N_8875);
nor U13140 (N_13140,N_8331,N_11629);
and U13141 (N_13141,N_9126,N_8237);
nand U13142 (N_13142,N_11143,N_11576);
nand U13143 (N_13143,N_9507,N_8905);
nand U13144 (N_13144,N_11234,N_8987);
xor U13145 (N_13145,N_11637,N_11112);
nand U13146 (N_13146,N_10423,N_10415);
nand U13147 (N_13147,N_9267,N_11522);
nor U13148 (N_13148,N_8663,N_10780);
or U13149 (N_13149,N_11845,N_8787);
nand U13150 (N_13150,N_10985,N_9885);
and U13151 (N_13151,N_10736,N_9183);
or U13152 (N_13152,N_11360,N_8015);
or U13153 (N_13153,N_8909,N_8216);
nand U13154 (N_13154,N_10494,N_11101);
nand U13155 (N_13155,N_8498,N_10009);
nand U13156 (N_13156,N_8821,N_11213);
nand U13157 (N_13157,N_10677,N_11055);
nand U13158 (N_13158,N_8458,N_9590);
nand U13159 (N_13159,N_8655,N_11538);
nand U13160 (N_13160,N_11183,N_11270);
xnor U13161 (N_13161,N_9903,N_11866);
nand U13162 (N_13162,N_8847,N_10629);
nor U13163 (N_13163,N_11667,N_10372);
and U13164 (N_13164,N_8892,N_8557);
or U13165 (N_13165,N_10429,N_10075);
xor U13166 (N_13166,N_10250,N_11137);
nor U13167 (N_13167,N_8634,N_9879);
nor U13168 (N_13168,N_8940,N_9207);
or U13169 (N_13169,N_8013,N_8412);
and U13170 (N_13170,N_11896,N_10689);
nand U13171 (N_13171,N_9270,N_10878);
or U13172 (N_13172,N_10049,N_9402);
and U13173 (N_13173,N_11520,N_8135);
nor U13174 (N_13174,N_10977,N_9030);
nor U13175 (N_13175,N_11421,N_10358);
nand U13176 (N_13176,N_8037,N_10183);
nor U13177 (N_13177,N_11358,N_8861);
or U13178 (N_13178,N_11930,N_9786);
nor U13179 (N_13179,N_11582,N_9980);
or U13180 (N_13180,N_10944,N_8735);
nor U13181 (N_13181,N_10367,N_10859);
nor U13182 (N_13182,N_10328,N_10348);
and U13183 (N_13183,N_9116,N_11999);
or U13184 (N_13184,N_8665,N_9729);
nor U13185 (N_13185,N_10113,N_9232);
nor U13186 (N_13186,N_8516,N_9911);
nand U13187 (N_13187,N_9187,N_9999);
and U13188 (N_13188,N_8024,N_9151);
or U13189 (N_13189,N_11976,N_10312);
nand U13190 (N_13190,N_10969,N_11753);
nand U13191 (N_13191,N_10161,N_8438);
nor U13192 (N_13192,N_9717,N_9234);
and U13193 (N_13193,N_9179,N_11387);
and U13194 (N_13194,N_11178,N_8040);
nand U13195 (N_13195,N_9749,N_11543);
nand U13196 (N_13196,N_11251,N_8780);
or U13197 (N_13197,N_10320,N_11549);
nor U13198 (N_13198,N_8432,N_8367);
nand U13199 (N_13199,N_9186,N_9410);
and U13200 (N_13200,N_8712,N_8302);
nand U13201 (N_13201,N_9810,N_11959);
and U13202 (N_13202,N_9756,N_9539);
nand U13203 (N_13203,N_10142,N_8441);
nand U13204 (N_13204,N_11595,N_10940);
nor U13205 (N_13205,N_9330,N_9965);
nand U13206 (N_13206,N_9927,N_11741);
nand U13207 (N_13207,N_9162,N_8175);
or U13208 (N_13208,N_8656,N_10968);
or U13209 (N_13209,N_10865,N_10132);
nor U13210 (N_13210,N_8051,N_8603);
and U13211 (N_13211,N_10110,N_11630);
and U13212 (N_13212,N_10021,N_9070);
nor U13213 (N_13213,N_8809,N_8521);
or U13214 (N_13214,N_9887,N_10334);
xor U13215 (N_13215,N_10081,N_9338);
or U13216 (N_13216,N_9367,N_11651);
or U13217 (N_13217,N_10659,N_11079);
nand U13218 (N_13218,N_9034,N_10500);
nand U13219 (N_13219,N_9509,N_11226);
nand U13220 (N_13220,N_10176,N_8234);
xnor U13221 (N_13221,N_8358,N_11371);
xnor U13222 (N_13222,N_8928,N_9800);
xnor U13223 (N_13223,N_8322,N_11105);
or U13224 (N_13224,N_9951,N_9016);
xnor U13225 (N_13225,N_11408,N_10259);
nand U13226 (N_13226,N_10032,N_8503);
or U13227 (N_13227,N_11990,N_11442);
or U13228 (N_13228,N_11193,N_9378);
xor U13229 (N_13229,N_9616,N_8636);
nand U13230 (N_13230,N_11721,N_8615);
nor U13231 (N_13231,N_10260,N_8179);
nor U13232 (N_13232,N_8550,N_9038);
nand U13233 (N_13233,N_9530,N_11145);
or U13234 (N_13234,N_11952,N_8753);
and U13235 (N_13235,N_8842,N_9542);
or U13236 (N_13236,N_11519,N_9392);
nand U13237 (N_13237,N_8020,N_9371);
and U13238 (N_13238,N_8360,N_10615);
nand U13239 (N_13239,N_10428,N_10056);
and U13240 (N_13240,N_8276,N_11854);
xnor U13241 (N_13241,N_10267,N_10211);
nor U13242 (N_13242,N_9595,N_9308);
or U13243 (N_13243,N_10469,N_9685);
nand U13244 (N_13244,N_8862,N_9974);
or U13245 (N_13245,N_11879,N_8080);
nand U13246 (N_13246,N_8617,N_10503);
xnor U13247 (N_13247,N_10193,N_11197);
xnor U13248 (N_13248,N_8827,N_8359);
xor U13249 (N_13249,N_9007,N_10851);
nor U13250 (N_13250,N_10252,N_8333);
nand U13251 (N_13251,N_8858,N_8771);
nor U13252 (N_13252,N_11950,N_8955);
or U13253 (N_13253,N_9171,N_9486);
and U13254 (N_13254,N_10208,N_8034);
nand U13255 (N_13255,N_10545,N_9596);
and U13256 (N_13256,N_10505,N_9002);
and U13257 (N_13257,N_10588,N_10168);
nor U13258 (N_13258,N_11940,N_10277);
xor U13259 (N_13259,N_10233,N_11900);
xor U13260 (N_13260,N_11660,N_11914);
or U13261 (N_13261,N_11579,N_9407);
nor U13262 (N_13262,N_8806,N_10617);
nand U13263 (N_13263,N_10138,N_8433);
and U13264 (N_13264,N_8413,N_8701);
and U13265 (N_13265,N_11984,N_10782);
nor U13266 (N_13266,N_9621,N_9329);
xnor U13267 (N_13267,N_8192,N_9182);
or U13268 (N_13268,N_11376,N_10376);
nor U13269 (N_13269,N_10439,N_11083);
nor U13270 (N_13270,N_8571,N_9769);
and U13271 (N_13271,N_9205,N_11130);
or U13272 (N_13272,N_10525,N_10655);
nand U13273 (N_13273,N_11634,N_11605);
nand U13274 (N_13274,N_11632,N_9377);
nor U13275 (N_13275,N_11386,N_10662);
or U13276 (N_13276,N_9363,N_8706);
xor U13277 (N_13277,N_11369,N_10587);
nand U13278 (N_13278,N_9870,N_10206);
nand U13279 (N_13279,N_9667,N_11781);
nand U13280 (N_13280,N_10526,N_8164);
and U13281 (N_13281,N_8574,N_11125);
nor U13282 (N_13282,N_10182,N_8981);
nand U13283 (N_13283,N_8825,N_11971);
nor U13284 (N_13284,N_10459,N_8857);
nand U13285 (N_13285,N_9427,N_8741);
or U13286 (N_13286,N_11047,N_9451);
xnor U13287 (N_13287,N_8823,N_11711);
or U13288 (N_13288,N_10533,N_10043);
nand U13289 (N_13289,N_11655,N_9463);
nor U13290 (N_13290,N_11968,N_11301);
nor U13291 (N_13291,N_8291,N_9020);
and U13292 (N_13292,N_11072,N_8410);
nor U13293 (N_13293,N_11554,N_11222);
nor U13294 (N_13294,N_9632,N_8813);
and U13295 (N_13295,N_9814,N_9021);
xnor U13296 (N_13296,N_8004,N_10997);
xor U13297 (N_13297,N_8480,N_10100);
or U13298 (N_13298,N_8556,N_11333);
xnor U13299 (N_13299,N_8766,N_8929);
nor U13300 (N_13300,N_9576,N_11048);
xor U13301 (N_13301,N_10776,N_8301);
nand U13302 (N_13302,N_10555,N_9071);
nor U13303 (N_13303,N_10856,N_11613);
nand U13304 (N_13304,N_9178,N_9865);
nand U13305 (N_13305,N_9947,N_9805);
or U13306 (N_13306,N_10189,N_11555);
nor U13307 (N_13307,N_11140,N_8240);
nand U13308 (N_13308,N_10906,N_10458);
or U13309 (N_13309,N_9401,N_10990);
nor U13310 (N_13310,N_9723,N_9424);
nor U13311 (N_13311,N_10828,N_10103);
nand U13312 (N_13312,N_10339,N_9782);
nand U13313 (N_13313,N_11192,N_11938);
nand U13314 (N_13314,N_10551,N_9607);
nand U13315 (N_13315,N_10242,N_9935);
nand U13316 (N_13316,N_9498,N_11174);
and U13317 (N_13317,N_8915,N_8838);
nand U13318 (N_13318,N_10220,N_9711);
nor U13319 (N_13319,N_8533,N_9415);
xnor U13320 (N_13320,N_11356,N_10293);
xor U13321 (N_13321,N_11265,N_8274);
nor U13322 (N_13322,N_9726,N_9483);
and U13323 (N_13323,N_11808,N_9801);
nand U13324 (N_13324,N_10660,N_9412);
and U13325 (N_13325,N_9066,N_8290);
nand U13326 (N_13326,N_11830,N_8467);
or U13327 (N_13327,N_11460,N_8883);
or U13328 (N_13328,N_11954,N_11069);
and U13329 (N_13329,N_8349,N_8296);
and U13330 (N_13330,N_9295,N_9991);
or U13331 (N_13331,N_8056,N_9718);
and U13332 (N_13332,N_10129,N_8383);
nand U13333 (N_13333,N_11937,N_11611);
nand U13334 (N_13334,N_11186,N_10929);
and U13335 (N_13335,N_9892,N_11792);
nand U13336 (N_13336,N_10974,N_9508);
or U13337 (N_13337,N_10289,N_8305);
or U13338 (N_13338,N_8213,N_11567);
nand U13339 (N_13339,N_8749,N_11385);
or U13340 (N_13340,N_9816,N_9216);
or U13341 (N_13341,N_8497,N_10025);
nor U13342 (N_13342,N_11151,N_9092);
nand U13343 (N_13343,N_11880,N_9586);
and U13344 (N_13344,N_9053,N_9419);
nor U13345 (N_13345,N_9147,N_9093);
and U13346 (N_13346,N_8017,N_10707);
nand U13347 (N_13347,N_8673,N_9058);
and U13348 (N_13348,N_9247,N_11716);
and U13349 (N_13349,N_8926,N_11610);
and U13350 (N_13350,N_8792,N_11009);
and U13351 (N_13351,N_8630,N_9396);
nor U13352 (N_13352,N_10236,N_10229);
xor U13353 (N_13353,N_11644,N_11443);
or U13354 (N_13354,N_8837,N_8608);
nor U13355 (N_13355,N_10047,N_10104);
nand U13356 (N_13356,N_10456,N_11093);
nand U13357 (N_13357,N_11618,N_11742);
nand U13358 (N_13358,N_10006,N_11242);
and U13359 (N_13359,N_8399,N_11881);
or U13360 (N_13360,N_9994,N_9231);
nand U13361 (N_13361,N_10738,N_11574);
and U13362 (N_13362,N_11772,N_9652);
nor U13363 (N_13363,N_8232,N_10881);
or U13364 (N_13364,N_11361,N_10218);
and U13365 (N_13365,N_10482,N_8765);
or U13366 (N_13366,N_9763,N_11905);
and U13367 (N_13367,N_8050,N_10502);
nand U13368 (N_13368,N_10635,N_10027);
and U13369 (N_13369,N_11518,N_8487);
and U13370 (N_13370,N_11016,N_10509);
and U13371 (N_13371,N_11552,N_8543);
and U13372 (N_13372,N_11038,N_10002);
nand U13373 (N_13373,N_9924,N_9113);
or U13374 (N_13374,N_10345,N_8514);
nor U13375 (N_13375,N_11287,N_10535);
nor U13376 (N_13376,N_11426,N_11034);
or U13377 (N_13377,N_11581,N_10594);
nand U13378 (N_13378,N_8767,N_8993);
nor U13379 (N_13379,N_9357,N_9815);
nor U13380 (N_13380,N_8177,N_8033);
and U13381 (N_13381,N_10630,N_10549);
nand U13382 (N_13382,N_10291,N_10510);
nand U13383 (N_13383,N_9740,N_8942);
or U13384 (N_13384,N_8491,N_9826);
and U13385 (N_13385,N_11225,N_10120);
xor U13386 (N_13386,N_9848,N_9641);
or U13387 (N_13387,N_11071,N_10887);
nor U13388 (N_13388,N_9251,N_11473);
or U13389 (N_13389,N_9283,N_9292);
or U13390 (N_13390,N_9611,N_8273);
xor U13391 (N_13391,N_9636,N_11622);
nand U13392 (N_13392,N_10717,N_10553);
or U13393 (N_13393,N_8236,N_9109);
and U13394 (N_13394,N_11402,N_8820);
or U13395 (N_13395,N_9260,N_11229);
and U13396 (N_13396,N_11490,N_10751);
and U13397 (N_13397,N_9556,N_10570);
or U13398 (N_13398,N_8893,N_9088);
nand U13399 (N_13399,N_10938,N_9633);
or U13400 (N_13400,N_9467,N_11382);
and U13401 (N_13401,N_11725,N_11415);
nor U13402 (N_13402,N_11537,N_11416);
and U13403 (N_13403,N_8148,N_11869);
and U13404 (N_13404,N_9495,N_9963);
nand U13405 (N_13405,N_10603,N_10232);
xnor U13406 (N_13406,N_8667,N_10083);
nor U13407 (N_13407,N_8187,N_10773);
nor U13408 (N_13408,N_8206,N_9841);
nand U13409 (N_13409,N_11918,N_11654);
and U13410 (N_13410,N_11013,N_9059);
nand U13411 (N_13411,N_8157,N_10371);
or U13412 (N_13412,N_11114,N_8527);
nand U13413 (N_13413,N_10699,N_11658);
nor U13414 (N_13414,N_10130,N_9748);
nor U13415 (N_13415,N_8980,N_11023);
nor U13416 (N_13416,N_11925,N_8036);
and U13417 (N_13417,N_9599,N_8102);
and U13418 (N_13418,N_10634,N_9880);
or U13419 (N_13419,N_9638,N_9743);
and U13420 (N_13420,N_10251,N_8416);
or U13421 (N_13421,N_8776,N_9700);
and U13422 (N_13422,N_9214,N_10196);
or U13423 (N_13423,N_8989,N_10651);
or U13424 (N_13424,N_9630,N_8889);
or U13425 (N_13425,N_8696,N_10419);
nand U13426 (N_13426,N_10845,N_11913);
or U13427 (N_13427,N_9747,N_10564);
nor U13428 (N_13428,N_8580,N_11833);
or U13429 (N_13429,N_11731,N_8581);
xnor U13430 (N_13430,N_8958,N_9886);
nor U13431 (N_13431,N_9549,N_10918);
nand U13432 (N_13432,N_8959,N_9715);
and U13433 (N_13433,N_10665,N_11891);
and U13434 (N_13434,N_10300,N_10144);
nand U13435 (N_13435,N_10779,N_8334);
nand U13436 (N_13436,N_10867,N_8264);
or U13437 (N_13437,N_9546,N_8631);
or U13438 (N_13438,N_10162,N_8779);
xor U13439 (N_13439,N_10105,N_11748);
nand U13440 (N_13440,N_10653,N_10684);
or U13441 (N_13441,N_10392,N_11132);
nand U13442 (N_13442,N_11056,N_8312);
nand U13443 (N_13443,N_10352,N_11974);
and U13444 (N_13444,N_11353,N_11521);
nor U13445 (N_13445,N_10891,N_10400);
or U13446 (N_13446,N_10824,N_9785);
nand U13447 (N_13447,N_11944,N_9890);
nor U13448 (N_13448,N_8954,N_8895);
xor U13449 (N_13449,N_11917,N_9069);
nor U13450 (N_13450,N_11282,N_9176);
or U13451 (N_13451,N_10190,N_10165);
nand U13452 (N_13452,N_10769,N_11820);
xnor U13453 (N_13453,N_11045,N_11107);
xor U13454 (N_13454,N_9326,N_11871);
nor U13455 (N_13455,N_11441,N_11017);
or U13456 (N_13456,N_10756,N_9940);
or U13457 (N_13457,N_11303,N_8442);
nor U13458 (N_13458,N_9325,N_10763);
nand U13459 (N_13459,N_8777,N_10761);
nor U13460 (N_13460,N_8495,N_11904);
and U13461 (N_13461,N_10810,N_11294);
and U13462 (N_13462,N_11239,N_9563);
xor U13463 (N_13463,N_8622,N_11570);
nor U13464 (N_13464,N_9876,N_11350);
nand U13465 (N_13465,N_9457,N_10514);
and U13466 (N_13466,N_9758,N_10031);
nor U13467 (N_13467,N_8259,N_8646);
or U13468 (N_13468,N_11401,N_11615);
and U13469 (N_13469,N_9003,N_11035);
xnor U13470 (N_13470,N_10068,N_8492);
nand U13471 (N_13471,N_8614,N_11811);
and U13472 (N_13472,N_8906,N_9453);
nor U13473 (N_13473,N_11756,N_8417);
nor U13474 (N_13474,N_10046,N_8083);
or U13475 (N_13475,N_9535,N_10992);
nand U13476 (N_13476,N_8540,N_9882);
and U13477 (N_13477,N_8132,N_9139);
or U13478 (N_13478,N_11840,N_8115);
nor U13479 (N_13479,N_8249,N_11996);
or U13480 (N_13480,N_8671,N_8113);
nor U13481 (N_13481,N_11533,N_8165);
xor U13482 (N_13482,N_8097,N_8310);
nand U13483 (N_13483,N_10143,N_9578);
nand U13484 (N_13484,N_10375,N_9028);
and U13485 (N_13485,N_11037,N_8151);
nand U13486 (N_13486,N_10026,N_8054);
and U13487 (N_13487,N_11977,N_11626);
and U13488 (N_13488,N_8002,N_9730);
xnor U13489 (N_13489,N_11688,N_8279);
or U13490 (N_13490,N_8944,N_11327);
and U13491 (N_13491,N_8073,N_10280);
nor U13492 (N_13492,N_11750,N_9760);
and U13493 (N_13493,N_11601,N_11566);
or U13494 (N_13494,N_10346,N_8052);
nor U13495 (N_13495,N_8384,N_9617);
nor U13496 (N_13496,N_8140,N_9351);
nor U13497 (N_13497,N_8254,N_10674);
xor U13498 (N_13498,N_8283,N_8599);
or U13499 (N_13499,N_11706,N_8263);
or U13500 (N_13500,N_8180,N_9668);
nand U13501 (N_13501,N_10657,N_10915);
nor U13502 (N_13502,N_11147,N_8652);
nand U13503 (N_13503,N_11482,N_11332);
or U13504 (N_13504,N_9098,N_10943);
or U13505 (N_13505,N_11793,N_9706);
xor U13506 (N_13506,N_10933,N_11461);
nor U13507 (N_13507,N_9408,N_8041);
nor U13508 (N_13508,N_8850,N_10480);
nor U13509 (N_13509,N_9558,N_9215);
and U13510 (N_13510,N_11775,N_8424);
and U13511 (N_13511,N_11033,N_8529);
and U13512 (N_13512,N_9005,N_9428);
nand U13513 (N_13513,N_11480,N_9941);
and U13514 (N_13514,N_9835,N_9914);
or U13515 (N_13515,N_11367,N_11170);
nand U13516 (N_13516,N_11004,N_11773);
and U13517 (N_13517,N_11909,N_8950);
nand U13518 (N_13518,N_10273,N_9833);
or U13519 (N_13519,N_10721,N_10946);
and U13520 (N_13520,N_10547,N_10752);
xor U13521 (N_13521,N_8045,N_10671);
xor U13522 (N_13522,N_8523,N_9133);
or U13523 (N_13523,N_11544,N_9386);
nand U13524 (N_13524,N_8076,N_11863);
and U13525 (N_13525,N_8573,N_9680);
nor U13526 (N_13526,N_11368,N_9347);
or U13527 (N_13527,N_8117,N_10154);
xor U13528 (N_13528,N_9484,N_10384);
xor U13529 (N_13529,N_11348,N_8876);
or U13530 (N_13530,N_9725,N_10281);
nor U13531 (N_13531,N_9602,N_9856);
nor U13532 (N_13532,N_9130,N_10265);
nor U13533 (N_13533,N_10912,N_9587);
and U13534 (N_13534,N_11922,N_9471);
nor U13535 (N_13535,N_9961,N_11359);
xor U13536 (N_13536,N_11064,N_11430);
nor U13537 (N_13537,N_11452,N_8995);
or U13538 (N_13538,N_8299,N_10475);
nand U13539 (N_13539,N_9855,N_8831);
nand U13540 (N_13540,N_8046,N_9783);
nand U13541 (N_13541,N_10984,N_11334);
and U13542 (N_13542,N_9413,N_8786);
and U13543 (N_13543,N_8863,N_8949);
nor U13544 (N_13544,N_11321,N_11979);
or U13545 (N_13545,N_8553,N_11961);
xor U13546 (N_13546,N_9908,N_8150);
nand U13547 (N_13547,N_9233,N_8488);
xor U13548 (N_13548,N_11176,N_9734);
nand U13549 (N_13549,N_11051,N_10860);
or U13550 (N_13550,N_8834,N_11259);
nand U13551 (N_13551,N_10783,N_9358);
or U13552 (N_13552,N_9893,N_11090);
and U13553 (N_13553,N_9101,N_9349);
and U13554 (N_13554,N_10654,N_10808);
xor U13555 (N_13555,N_8284,N_10366);
xor U13556 (N_13556,N_8395,N_9724);
or U13557 (N_13557,N_9916,N_8695);
nor U13558 (N_13558,N_11020,N_9465);
nor U13559 (N_13559,N_8968,N_9051);
nor U13560 (N_13560,N_8532,N_10976);
xnor U13561 (N_13561,N_8070,N_10011);
and U13562 (N_13562,N_11843,N_10694);
or U13563 (N_13563,N_10967,N_11438);
or U13564 (N_13564,N_9443,N_11188);
or U13565 (N_13565,N_9654,N_10158);
and U13566 (N_13566,N_10426,N_11659);
or U13567 (N_13567,N_10724,N_9931);
nand U13568 (N_13568,N_10958,N_8154);
and U13569 (N_13569,N_8505,N_11673);
or U13570 (N_13570,N_10070,N_11548);
and U13571 (N_13571,N_8711,N_10548);
or U13572 (N_13572,N_8984,N_9584);
and U13573 (N_13573,N_10872,N_9501);
or U13574 (N_13574,N_11710,N_11102);
or U13575 (N_13575,N_9751,N_11062);
nor U13576 (N_13576,N_10628,N_9839);
xnor U13577 (N_13577,N_8398,N_11831);
nor U13578 (N_13578,N_9834,N_9891);
xor U13579 (N_13579,N_9533,N_11419);
nor U13580 (N_13580,N_11508,N_8651);
nor U13581 (N_13581,N_10691,N_9406);
nand U13582 (N_13582,N_11131,N_9571);
or U13583 (N_13583,N_10017,N_8688);
and U13584 (N_13584,N_11886,N_9553);
nor U13585 (N_13585,N_8466,N_11230);
nand U13586 (N_13586,N_10622,N_8947);
nor U13587 (N_13587,N_10612,N_9601);
or U13588 (N_13588,N_10898,N_10111);
and U13589 (N_13589,N_9944,N_8566);
nand U13590 (N_13590,N_10373,N_10406);
or U13591 (N_13591,N_8943,N_8314);
or U13592 (N_13592,N_9459,N_11433);
and U13593 (N_13593,N_8887,N_11877);
nand U13594 (N_13594,N_10246,N_8282);
and U13595 (N_13595,N_11908,N_11187);
or U13596 (N_13596,N_11649,N_8578);
xor U13597 (N_13597,N_8936,N_10796);
or U13598 (N_13598,N_8808,N_10513);
or U13599 (N_13599,N_11691,N_10209);
nor U13600 (N_13600,N_11096,N_10317);
nor U13601 (N_13601,N_11789,N_10966);
nand U13602 (N_13602,N_9606,N_11232);
nand U13603 (N_13603,N_8997,N_8173);
nand U13604 (N_13604,N_11001,N_10638);
xor U13605 (N_13605,N_11747,N_11768);
or U13606 (N_13606,N_11000,N_10135);
nand U13607 (N_13607,N_11864,N_10248);
or U13608 (N_13608,N_11043,N_9191);
or U13609 (N_13609,N_9494,N_10418);
nor U13610 (N_13610,N_9290,N_10318);
and U13611 (N_13611,N_10012,N_9545);
nand U13612 (N_13612,N_8589,N_10270);
nand U13613 (N_13613,N_11559,N_8105);
xnor U13614 (N_13614,N_10746,N_8355);
nand U13615 (N_13615,N_10608,N_8001);
nand U13616 (N_13616,N_9568,N_8560);
nor U13617 (N_13617,N_10646,N_8408);
xnor U13618 (N_13618,N_11025,N_8869);
and U13619 (N_13619,N_11141,N_10798);
nand U13620 (N_13620,N_8366,N_11286);
nand U13621 (N_13621,N_9698,N_11616);
or U13622 (N_13622,N_9912,N_10614);
nand U13623 (N_13623,N_9863,N_10447);
and U13624 (N_13624,N_10847,N_8055);
nand U13625 (N_13625,N_8659,N_10349);
xnor U13626 (N_13626,N_11138,N_8022);
or U13627 (N_13627,N_8760,N_9206);
and U13628 (N_13628,N_9366,N_8904);
nand U13629 (N_13629,N_9293,N_10683);
and U13630 (N_13630,N_10790,N_10822);
nor U13631 (N_13631,N_9299,N_9146);
or U13632 (N_13632,N_10343,N_9989);
nand U13633 (N_13633,N_10620,N_10210);
or U13634 (N_13634,N_8202,N_11647);
and U13635 (N_13635,N_10820,N_10298);
or U13636 (N_13636,N_9282,N_8620);
and U13637 (N_13637,N_8810,N_10247);
or U13638 (N_13638,N_9765,N_10584);
nor U13639 (N_13639,N_10637,N_9027);
or U13640 (N_13640,N_9666,N_11842);
nor U13641 (N_13641,N_8545,N_8967);
and U13642 (N_13642,N_11794,N_11022);
nor U13643 (N_13643,N_10230,N_9190);
nand U13644 (N_13644,N_8973,N_10914);
xnor U13645 (N_13645,N_10838,N_9499);
or U13646 (N_13646,N_11894,N_11088);
nand U13647 (N_13647,N_10263,N_10515);
nand U13648 (N_13648,N_10327,N_10644);
xor U13649 (N_13649,N_11645,N_8930);
or U13650 (N_13650,N_11511,N_10491);
and U13651 (N_13651,N_11116,N_11657);
nor U13652 (N_13652,N_10883,N_8086);
nand U13653 (N_13653,N_10786,N_11500);
nand U13654 (N_13654,N_9592,N_9211);
nor U13655 (N_13655,N_10817,N_10507);
and U13656 (N_13656,N_11827,N_9393);
nor U13657 (N_13657,N_11936,N_11912);
nand U13658 (N_13658,N_9772,N_9798);
or U13659 (N_13659,N_11726,N_8085);
and U13660 (N_13660,N_11528,N_8048);
and U13661 (N_13661,N_10156,N_11602);
or U13662 (N_13662,N_11816,N_11296);
nor U13663 (N_13663,N_10041,N_9564);
and U13664 (N_13664,N_10069,N_8965);
nand U13665 (N_13665,N_8309,N_8043);
nor U13666 (N_13666,N_11988,N_9960);
nand U13667 (N_13667,N_9675,N_8010);
nand U13668 (N_13668,N_10173,N_11892);
or U13669 (N_13669,N_8144,N_9619);
nand U13670 (N_13670,N_8452,N_8275);
nor U13671 (N_13671,N_11414,N_11700);
nor U13672 (N_13672,N_9566,N_10706);
xnor U13673 (N_13673,N_10892,N_11210);
nor U13674 (N_13674,N_10889,N_11070);
or U13675 (N_13675,N_9324,N_9121);
nor U13676 (N_13676,N_9682,N_8855);
nor U13677 (N_13677,N_8231,N_8029);
nor U13678 (N_13678,N_11736,N_8833);
nand U13679 (N_13679,N_10147,N_10093);
nand U13680 (N_13680,N_9694,N_10930);
nor U13681 (N_13681,N_10115,N_9532);
nand U13682 (N_13682,N_9149,N_9901);
xor U13683 (N_13683,N_9664,N_10536);
nor U13684 (N_13684,N_11370,N_8368);
xnor U13685 (N_13685,N_9753,N_9274);
xnor U13686 (N_13686,N_11336,N_11289);
and U13687 (N_13687,N_9439,N_9356);
or U13688 (N_13688,N_9953,N_8485);
and U13689 (N_13689,N_10972,N_9217);
and U13690 (N_13690,N_10410,N_8536);
and U13691 (N_13691,N_9714,N_10512);
and U13692 (N_13692,N_11884,N_10059);
nand U13693 (N_13693,N_9889,N_10540);
or U13694 (N_13694,N_11180,N_10561);
and U13695 (N_13695,N_10444,N_8546);
or U13696 (N_13696,N_9155,N_9449);
and U13697 (N_13697,N_11245,N_8729);
and U13698 (N_13698,N_8295,N_11694);
or U13699 (N_13699,N_10685,N_9802);
nor U13700 (N_13700,N_9181,N_11516);
and U13701 (N_13701,N_11300,N_9672);
nor U13702 (N_13702,N_11207,N_9626);
nand U13703 (N_13703,N_8226,N_11322);
xnor U13704 (N_13704,N_8750,N_10758);
nor U13705 (N_13705,N_9137,N_9213);
and U13706 (N_13706,N_8018,N_8125);
xnor U13707 (N_13707,N_9143,N_10187);
nor U13708 (N_13708,N_8471,N_8913);
nor U13709 (N_13709,N_11489,N_10956);
nor U13710 (N_13710,N_9033,N_8124);
nand U13711 (N_13711,N_9169,N_10961);
or U13712 (N_13712,N_10146,N_8852);
nor U13713 (N_13713,N_11205,N_11823);
xnor U13714 (N_13714,N_8446,N_8253);
nor U13715 (N_13715,N_11980,N_9655);
or U13716 (N_13716,N_11981,N_11607);
and U13717 (N_13717,N_11351,N_10823);
or U13718 (N_13718,N_10019,N_9696);
nand U13719 (N_13719,N_10740,N_9097);
nand U13720 (N_13720,N_10821,N_10417);
nand U13721 (N_13721,N_9057,N_10303);
xor U13722 (N_13722,N_10690,N_8183);
nand U13723 (N_13723,N_10222,N_9710);
nor U13724 (N_13724,N_10816,N_8340);
nor U13725 (N_13725,N_10076,N_8072);
and U13726 (N_13726,N_11404,N_11547);
and U13727 (N_13727,N_9777,N_11127);
and U13728 (N_13728,N_11256,N_10508);
nor U13729 (N_13729,N_8642,N_9475);
nor U13730 (N_13730,N_9300,N_10370);
nor U13731 (N_13731,N_9757,N_9489);
nor U13732 (N_13732,N_8381,N_9878);
and U13733 (N_13733,N_10264,N_9918);
nor U13734 (N_13734,N_8101,N_8356);
or U13735 (N_13735,N_8229,N_9840);
and U13736 (N_13736,N_11422,N_10730);
and U13737 (N_13737,N_8353,N_10321);
nand U13738 (N_13738,N_10516,N_9144);
or U13739 (N_13739,N_9250,N_8460);
or U13740 (N_13740,N_10029,N_10284);
and U13741 (N_13741,N_11466,N_9381);
nand U13742 (N_13742,N_11400,N_8520);
nand U13743 (N_13743,N_10499,N_11530);
nor U13744 (N_13744,N_10899,N_9708);
nand U13745 (N_13745,N_9517,N_10096);
nor U13746 (N_13746,N_11094,N_11902);
xor U13747 (N_13747,N_9697,N_9691);
nor U13748 (N_13748,N_8707,N_11814);
nand U13749 (N_13749,N_11875,N_9645);
nand U13750 (N_13750,N_9639,N_10199);
nand U13751 (N_13751,N_9305,N_9515);
nand U13752 (N_13752,N_8911,N_9719);
nand U13753 (N_13753,N_8031,N_10703);
or U13754 (N_13754,N_8717,N_9650);
and U13755 (N_13755,N_9631,N_11425);
nor U13756 (N_13756,N_8694,N_9609);
and U13757 (N_13757,N_9411,N_11058);
nand U13758 (N_13758,N_10167,N_10464);
xor U13759 (N_13759,N_9713,N_11458);
and U13760 (N_13760,N_10201,N_10592);
or U13761 (N_13761,N_9746,N_11844);
and U13762 (N_13762,N_11373,N_11633);
or U13763 (N_13763,N_10286,N_8088);
or U13764 (N_13764,N_10714,N_11005);
nor U13765 (N_13765,N_8007,N_11254);
or U13766 (N_13766,N_8435,N_8899);
xnor U13767 (N_13767,N_11260,N_11054);
nand U13768 (N_13768,N_9792,N_11682);
and U13769 (N_13769,N_11527,N_10381);
nor U13770 (N_13770,N_9830,N_8588);
nor U13771 (N_13771,N_9442,N_10483);
nand U13772 (N_13772,N_10853,N_8393);
nand U13773 (N_13773,N_9063,N_9054);
and U13774 (N_13774,N_9420,N_8635);
nand U13775 (N_13775,N_8189,N_8524);
or U13776 (N_13776,N_9257,N_8619);
and U13777 (N_13777,N_8966,N_10739);
nor U13778 (N_13778,N_11298,N_11588);
nor U13779 (N_13779,N_9469,N_10708);
nand U13780 (N_13780,N_10833,N_11701);
nor U13781 (N_13781,N_10863,N_11082);
nand U13782 (N_13782,N_9794,N_10559);
and U13783 (N_13783,N_11539,N_11364);
nand U13784 (N_13784,N_9141,N_10401);
or U13785 (N_13785,N_9373,N_10237);
xnor U13786 (N_13786,N_10094,N_9094);
or U13787 (N_13787,N_10987,N_10607);
nand U13788 (N_13788,N_10534,N_9385);
and U13789 (N_13789,N_9842,N_8490);
or U13790 (N_13790,N_11190,N_11126);
and U13791 (N_13791,N_10090,N_8963);
and U13792 (N_13792,N_10360,N_11485);
nand U13793 (N_13793,N_8058,N_9120);
or U13794 (N_13794,N_10493,N_11459);
nand U13795 (N_13795,N_9081,N_9342);
or U13796 (N_13796,N_11526,N_9627);
and U13797 (N_13797,N_11123,N_9488);
nor U13798 (N_13798,N_11873,N_10884);
nand U13799 (N_13799,N_10791,N_8687);
xnor U13800 (N_13800,N_9050,N_11257);
nand U13801 (N_13801,N_11888,N_10239);
nor U13802 (N_13802,N_11860,N_11568);
xor U13803 (N_13803,N_8848,N_8090);
nand U13804 (N_13804,N_11191,N_9380);
and U13805 (N_13805,N_8141,N_9635);
nor U13806 (N_13806,N_11995,N_8405);
nor U13807 (N_13807,N_11159,N_10705);
xnor U13808 (N_13808,N_9227,N_11044);
and U13809 (N_13809,N_10599,N_9313);
nand U13810 (N_13810,N_11859,N_9969);
nor U13811 (N_13811,N_8734,N_10667);
and U13812 (N_13812,N_8816,N_10980);
and U13813 (N_13813,N_11019,N_8223);
nand U13814 (N_13814,N_11175,N_11049);
nor U13815 (N_13815,N_8525,N_8724);
nand U13816 (N_13816,N_11394,N_8044);
or U13817 (N_13817,N_8461,N_11687);
xor U13818 (N_13818,N_10998,N_11249);
nand U13819 (N_13819,N_9768,N_10580);
or U13820 (N_13820,N_9721,N_8731);
xnor U13821 (N_13821,N_8856,N_10163);
and U13822 (N_13822,N_10127,N_10389);
nand U13823 (N_13823,N_11391,N_9897);
or U13824 (N_13824,N_8204,N_11429);
nand U13825 (N_13825,N_9643,N_9637);
xnor U13826 (N_13826,N_10869,N_8888);
xor U13827 (N_13827,N_10762,N_8047);
and U13828 (N_13828,N_8025,N_9107);
or U13829 (N_13829,N_11299,N_11238);
nand U13830 (N_13830,N_8171,N_8674);
and U13831 (N_13831,N_11920,N_10266);
or U13832 (N_13832,N_8162,N_11194);
nand U13833 (N_13833,N_8160,N_11758);
and U13834 (N_13834,N_11437,N_9485);
nor U13835 (N_13835,N_10479,N_10234);
nand U13836 (N_13836,N_9052,N_8504);
nand U13837 (N_13837,N_10896,N_10905);
or U13838 (N_13838,N_11246,N_10207);
xnor U13839 (N_13839,N_8682,N_10403);
and U13840 (N_13840,N_8209,N_9437);
or U13841 (N_13841,N_8935,N_10226);
nor U13842 (N_13842,N_11209,N_11620);
nor U13843 (N_13843,N_10038,N_8190);
and U13844 (N_13844,N_8970,N_9204);
and U13845 (N_13845,N_10787,N_9080);
nand U13846 (N_13846,N_9196,N_9526);
nor U13847 (N_13847,N_11578,N_10877);
nand U13848 (N_13848,N_9245,N_8841);
or U13849 (N_13849,N_8535,N_9529);
xnor U13850 (N_13850,N_9135,N_11199);
nor U13851 (N_13851,N_9273,N_10506);
nor U13852 (N_13852,N_8618,N_9936);
nor U13853 (N_13853,N_11978,N_8469);
nor U13854 (N_13854,N_10052,N_10227);
and U13855 (N_13855,N_8470,N_11817);
nand U13856 (N_13856,N_8208,N_8449);
nor U13857 (N_13857,N_8817,N_9226);
and U13858 (N_13858,N_8403,N_11608);
nand U13859 (N_13859,N_11571,N_11822);
xnor U13860 (N_13860,N_10681,N_11383);
nor U13861 (N_13861,N_11290,N_8390);
or U13862 (N_13862,N_8768,N_8784);
nor U13863 (N_13863,N_9175,N_11600);
nor U13864 (N_13864,N_9466,N_9421);
nand U13865 (N_13865,N_10696,N_9286);
nor U13866 (N_13866,N_8387,N_8375);
or U13867 (N_13867,N_9646,N_11163);
and U13868 (N_13868,N_10305,N_9669);
nand U13869 (N_13869,N_10831,N_11702);
xnor U13870 (N_13870,N_10340,N_9372);
nand U13871 (N_13871,N_9538,N_11901);
nor U13872 (N_13872,N_8732,N_10243);
nand U13873 (N_13873,N_9822,N_10854);
nand U13874 (N_13874,N_10675,N_10033);
and U13875 (N_13875,N_9154,N_10571);
nor U13876 (N_13876,N_10050,N_11208);
and U13877 (N_13877,N_10722,N_11293);
and U13878 (N_13878,N_11783,N_11158);
or U13879 (N_13879,N_9455,N_8339);
nand U13880 (N_13880,N_9423,N_11319);
or U13881 (N_13881,N_11947,N_9065);
or U13882 (N_13882,N_8348,N_9784);
nor U13883 (N_13883,N_10336,N_10007);
or U13884 (N_13884,N_9898,N_9791);
nand U13885 (N_13885,N_11639,N_10600);
nand U13886 (N_13886,N_11103,N_8319);
nor U13887 (N_13887,N_11895,N_8681);
and U13888 (N_13888,N_9243,N_11381);
nand U13889 (N_13889,N_10067,N_9759);
and U13890 (N_13890,N_11580,N_9512);
and U13891 (N_13891,N_11481,N_10532);
and U13892 (N_13892,N_8084,N_9258);
nand U13893 (N_13893,N_8330,N_10013);
nor U13894 (N_13894,N_10468,N_8789);
nand U13895 (N_13895,N_8843,N_8871);
or U13896 (N_13896,N_8534,N_8392);
or U13897 (N_13897,N_9997,N_11919);
and U13898 (N_13898,N_10978,N_9525);
xnor U13899 (N_13899,N_10605,N_8421);
and U13900 (N_13900,N_11255,N_11734);
nor U13901 (N_13901,N_11565,N_11856);
and U13902 (N_13902,N_11717,N_10225);
and U13903 (N_13903,N_8988,N_9952);
and U13904 (N_13904,N_8645,N_8255);
or U13905 (N_13905,N_9658,N_11476);
or U13906 (N_13906,N_9452,N_8459);
or U13907 (N_13907,N_11587,N_9869);
nor U13908 (N_13908,N_10785,N_10369);
and U13909 (N_13909,N_11501,N_10598);
and U13910 (N_13910,N_9004,N_10697);
or U13911 (N_13911,N_11224,N_8804);
xor U13912 (N_13912,N_9049,N_9491);
xor U13913 (N_13913,N_10800,N_11708);
nor U13914 (N_13914,N_9910,N_8268);
xor U13915 (N_13915,N_11346,N_11828);
nor U13916 (N_13916,N_11890,N_11181);
or U13917 (N_13917,N_11737,N_10159);
xnor U13918 (N_13918,N_10954,N_10825);
and U13919 (N_13919,N_8479,N_8758);
nand U13920 (N_13920,N_11732,N_9781);
or U13921 (N_13921,N_9089,N_10153);
nand U13922 (N_13922,N_10700,N_10537);
nand U13923 (N_13923,N_10917,N_10062);
nor U13924 (N_13924,N_9588,N_11994);
and U13925 (N_13925,N_10408,N_8609);
and U13926 (N_13926,N_9416,N_9010);
nor U13927 (N_13927,N_9046,N_11883);
and U13928 (N_13928,N_8427,N_9790);
nor U13929 (N_13929,N_9567,N_10663);
nand U13930 (N_13930,N_8464,N_11625);
nand U13931 (N_13931,N_9060,N_11085);
or U13932 (N_13932,N_9648,N_10125);
and U13933 (N_13933,N_10215,N_8347);
and U13934 (N_13934,N_11277,N_10504);
xor U13935 (N_13935,N_10812,N_11474);
or U13936 (N_13936,N_10926,N_8544);
nand U13937 (N_13937,N_9852,N_11142);
nand U13938 (N_13938,N_9966,N_9445);
or U13939 (N_13939,N_10765,N_9318);
and U13940 (N_13940,N_9014,N_11872);
nand U13941 (N_13941,N_10718,N_8638);
nand U13942 (N_13942,N_10460,N_8998);
nor U13943 (N_13943,N_10979,N_9968);
nor U13944 (N_13944,N_10687,N_8625);
nor U13945 (N_13945,N_9043,N_8436);
or U13946 (N_13946,N_8409,N_9904);
xor U13947 (N_13947,N_11850,N_11824);
nor U13948 (N_13948,N_10455,N_10855);
nand U13949 (N_13949,N_8476,N_11720);
or U13950 (N_13950,N_10797,N_8394);
or U13951 (N_13951,N_10443,N_9271);
nor U13952 (N_13952,N_10307,N_10353);
and U13953 (N_13953,N_10811,N_10397);
nand U13954 (N_13954,N_11531,N_9249);
nand U13955 (N_13955,N_11162,N_9695);
nor U13956 (N_13956,N_11467,N_11921);
nand U13957 (N_13957,N_9382,N_9011);
xor U13958 (N_13958,N_8986,N_8327);
xor U13959 (N_13959,N_9035,N_11486);
or U13960 (N_13960,N_9032,N_9365);
nand U13961 (N_13961,N_10486,N_11212);
nand U13962 (N_13962,N_11776,N_8059);
and U13963 (N_13963,N_9540,N_8313);
and U13964 (N_13964,N_9686,N_10325);
nand U13965 (N_13965,N_11815,N_10481);
nand U13966 (N_13966,N_9345,N_11272);
or U13967 (N_13967,N_11354,N_9480);
nor U13968 (N_13968,N_9315,N_8244);
xor U13969 (N_13969,N_8672,N_11785);
nand U13970 (N_13970,N_11686,N_8607);
nor U13971 (N_13971,N_9909,N_9933);
nand U13972 (N_13972,N_8598,N_8120);
nand U13973 (N_13973,N_10572,N_11075);
nand U13974 (N_13974,N_9266,N_8363);
nand U13975 (N_13975,N_9779,N_8948);
xnor U13976 (N_13976,N_8320,N_10970);
nand U13977 (N_13977,N_8114,N_11932);
nor U13978 (N_13978,N_10996,N_8733);
and U13979 (N_13979,N_9524,N_10875);
nand U13980 (N_13980,N_11653,N_11363);
nor U13981 (N_13981,N_10964,N_9111);
or U13982 (N_13982,N_10010,N_10661);
nor U13983 (N_13983,N_8252,N_11507);
and U13984 (N_13984,N_9444,N_11948);
or U13985 (N_13985,N_11619,N_8867);
xor U13986 (N_13986,N_11362,N_9915);
and U13987 (N_13987,N_8924,N_11743);
or U13988 (N_13988,N_11258,N_10131);
xnor U13989 (N_13989,N_9261,N_10139);
or U13990 (N_13990,N_11993,N_9041);
and U13991 (N_13991,N_8094,N_11761);
nand U13992 (N_13992,N_8003,N_10178);
nor U13993 (N_13993,N_9164,N_10715);
nor U13994 (N_13994,N_10213,N_11663);
nor U13995 (N_13995,N_9945,N_10474);
nand U13996 (N_13996,N_9788,N_11339);
nor U13997 (N_13997,N_11975,N_9022);
nand U13998 (N_13998,N_10949,N_9932);
nand U13999 (N_13999,N_10576,N_10057);
and U14000 (N_14000,N_10054,N_9616);
or U14001 (N_14001,N_10689,N_8358);
xor U14002 (N_14002,N_8826,N_10224);
nor U14003 (N_14003,N_9739,N_11232);
nand U14004 (N_14004,N_11267,N_8867);
nor U14005 (N_14005,N_11363,N_8491);
or U14006 (N_14006,N_10319,N_8051);
and U14007 (N_14007,N_8860,N_9857);
nand U14008 (N_14008,N_10390,N_10282);
and U14009 (N_14009,N_9139,N_9796);
nand U14010 (N_14010,N_10868,N_9167);
or U14011 (N_14011,N_8433,N_11760);
and U14012 (N_14012,N_11946,N_9123);
xnor U14013 (N_14013,N_11459,N_9913);
or U14014 (N_14014,N_8279,N_11822);
or U14015 (N_14015,N_11956,N_11018);
nor U14016 (N_14016,N_11544,N_10508);
or U14017 (N_14017,N_8445,N_8612);
and U14018 (N_14018,N_8267,N_10063);
or U14019 (N_14019,N_11928,N_9916);
nor U14020 (N_14020,N_11490,N_11492);
and U14021 (N_14021,N_8925,N_8882);
or U14022 (N_14022,N_8259,N_11725);
or U14023 (N_14023,N_9219,N_10578);
nor U14024 (N_14024,N_9928,N_11839);
or U14025 (N_14025,N_11790,N_10279);
or U14026 (N_14026,N_11721,N_8291);
or U14027 (N_14027,N_10990,N_8459);
or U14028 (N_14028,N_9901,N_11700);
or U14029 (N_14029,N_8212,N_11939);
nand U14030 (N_14030,N_11877,N_9958);
xnor U14031 (N_14031,N_9080,N_10226);
nor U14032 (N_14032,N_10276,N_11249);
or U14033 (N_14033,N_8914,N_9475);
nand U14034 (N_14034,N_11023,N_10676);
nor U14035 (N_14035,N_9838,N_10508);
nor U14036 (N_14036,N_9488,N_10300);
nor U14037 (N_14037,N_10265,N_10930);
nand U14038 (N_14038,N_8363,N_11184);
nor U14039 (N_14039,N_11278,N_10394);
and U14040 (N_14040,N_9724,N_10473);
and U14041 (N_14041,N_11367,N_11674);
nor U14042 (N_14042,N_9787,N_11048);
and U14043 (N_14043,N_8042,N_9114);
nand U14044 (N_14044,N_10148,N_8872);
or U14045 (N_14045,N_11409,N_10070);
nor U14046 (N_14046,N_11799,N_11824);
nor U14047 (N_14047,N_9328,N_10984);
or U14048 (N_14048,N_10654,N_9611);
nand U14049 (N_14049,N_11257,N_8891);
and U14050 (N_14050,N_10266,N_8701);
nor U14051 (N_14051,N_11043,N_8244);
nand U14052 (N_14052,N_8975,N_9131);
nand U14053 (N_14053,N_9294,N_9387);
nand U14054 (N_14054,N_10944,N_11658);
or U14055 (N_14055,N_8788,N_11268);
nand U14056 (N_14056,N_10122,N_11139);
nor U14057 (N_14057,N_11669,N_10858);
xor U14058 (N_14058,N_10665,N_8250);
nor U14059 (N_14059,N_8958,N_8601);
or U14060 (N_14060,N_11262,N_9878);
or U14061 (N_14061,N_10254,N_11900);
xor U14062 (N_14062,N_11149,N_11250);
nor U14063 (N_14063,N_9539,N_8106);
or U14064 (N_14064,N_9030,N_10577);
nand U14065 (N_14065,N_10631,N_10814);
or U14066 (N_14066,N_10750,N_9446);
nand U14067 (N_14067,N_8067,N_11414);
nand U14068 (N_14068,N_8072,N_10318);
xnor U14069 (N_14069,N_8684,N_9900);
nor U14070 (N_14070,N_8584,N_11971);
and U14071 (N_14071,N_8833,N_10753);
xor U14072 (N_14072,N_10156,N_8259);
nor U14073 (N_14073,N_8706,N_8358);
or U14074 (N_14074,N_10575,N_9578);
nand U14075 (N_14075,N_9196,N_9053);
nor U14076 (N_14076,N_10863,N_9747);
nand U14077 (N_14077,N_10108,N_8400);
or U14078 (N_14078,N_9871,N_8279);
and U14079 (N_14079,N_8623,N_9817);
nor U14080 (N_14080,N_8547,N_8248);
nand U14081 (N_14081,N_11099,N_8912);
xnor U14082 (N_14082,N_11165,N_8785);
and U14083 (N_14083,N_8034,N_10167);
nor U14084 (N_14084,N_11691,N_9499);
nand U14085 (N_14085,N_10391,N_9063);
nand U14086 (N_14086,N_8566,N_8118);
and U14087 (N_14087,N_8497,N_9464);
nand U14088 (N_14088,N_9434,N_8187);
nand U14089 (N_14089,N_10394,N_9953);
nor U14090 (N_14090,N_11329,N_10118);
nand U14091 (N_14091,N_8118,N_11812);
xnor U14092 (N_14092,N_8810,N_11744);
nand U14093 (N_14093,N_10729,N_10744);
xnor U14094 (N_14094,N_8342,N_11337);
nand U14095 (N_14095,N_9398,N_11873);
or U14096 (N_14096,N_11812,N_11411);
nor U14097 (N_14097,N_11152,N_10727);
nor U14098 (N_14098,N_10195,N_11832);
nand U14099 (N_14099,N_11606,N_8981);
and U14100 (N_14100,N_8380,N_11893);
and U14101 (N_14101,N_11928,N_8492);
and U14102 (N_14102,N_8060,N_9048);
and U14103 (N_14103,N_10912,N_9035);
and U14104 (N_14104,N_8653,N_9027);
and U14105 (N_14105,N_8857,N_10152);
nor U14106 (N_14106,N_11736,N_11875);
or U14107 (N_14107,N_9357,N_8474);
nor U14108 (N_14108,N_11904,N_9324);
nand U14109 (N_14109,N_9254,N_9749);
or U14110 (N_14110,N_8788,N_8724);
xor U14111 (N_14111,N_8835,N_8833);
nor U14112 (N_14112,N_10494,N_8301);
xnor U14113 (N_14113,N_10382,N_11671);
nand U14114 (N_14114,N_8351,N_11430);
nor U14115 (N_14115,N_8218,N_8696);
or U14116 (N_14116,N_10411,N_8637);
or U14117 (N_14117,N_10565,N_10038);
nand U14118 (N_14118,N_8758,N_11868);
and U14119 (N_14119,N_8590,N_11622);
or U14120 (N_14120,N_10538,N_9545);
nor U14121 (N_14121,N_11707,N_8096);
nor U14122 (N_14122,N_11620,N_10983);
or U14123 (N_14123,N_8920,N_10806);
nand U14124 (N_14124,N_8075,N_11760);
nor U14125 (N_14125,N_9690,N_10813);
or U14126 (N_14126,N_8790,N_9353);
or U14127 (N_14127,N_9195,N_11230);
and U14128 (N_14128,N_9526,N_10354);
nor U14129 (N_14129,N_10719,N_10415);
nor U14130 (N_14130,N_11675,N_11348);
or U14131 (N_14131,N_8764,N_11795);
nand U14132 (N_14132,N_11929,N_11259);
xor U14133 (N_14133,N_10952,N_8337);
and U14134 (N_14134,N_8478,N_11615);
or U14135 (N_14135,N_8411,N_11588);
nand U14136 (N_14136,N_9349,N_9616);
nand U14137 (N_14137,N_10369,N_8857);
nor U14138 (N_14138,N_9978,N_9751);
nand U14139 (N_14139,N_8041,N_8046);
and U14140 (N_14140,N_9257,N_10226);
nand U14141 (N_14141,N_10588,N_11508);
nand U14142 (N_14142,N_10709,N_8135);
or U14143 (N_14143,N_10874,N_10643);
nand U14144 (N_14144,N_10429,N_9864);
nor U14145 (N_14145,N_8056,N_9894);
nand U14146 (N_14146,N_9224,N_8937);
nor U14147 (N_14147,N_8631,N_10797);
nor U14148 (N_14148,N_9513,N_10906);
nor U14149 (N_14149,N_10366,N_11648);
nand U14150 (N_14150,N_9429,N_8532);
and U14151 (N_14151,N_8691,N_8304);
or U14152 (N_14152,N_10805,N_9230);
nand U14153 (N_14153,N_10728,N_9400);
and U14154 (N_14154,N_9647,N_9795);
nand U14155 (N_14155,N_9533,N_11566);
or U14156 (N_14156,N_9871,N_8311);
and U14157 (N_14157,N_10599,N_10921);
nand U14158 (N_14158,N_8424,N_9101);
and U14159 (N_14159,N_11686,N_11767);
and U14160 (N_14160,N_9994,N_10919);
or U14161 (N_14161,N_8262,N_9782);
nor U14162 (N_14162,N_10771,N_10806);
xnor U14163 (N_14163,N_9525,N_8899);
nor U14164 (N_14164,N_8545,N_9142);
nor U14165 (N_14165,N_9213,N_10851);
and U14166 (N_14166,N_8394,N_8370);
or U14167 (N_14167,N_9261,N_10390);
nor U14168 (N_14168,N_10160,N_8486);
and U14169 (N_14169,N_10297,N_9295);
and U14170 (N_14170,N_8003,N_10188);
nand U14171 (N_14171,N_9169,N_8736);
nor U14172 (N_14172,N_8988,N_8736);
and U14173 (N_14173,N_9485,N_9620);
or U14174 (N_14174,N_10687,N_8061);
or U14175 (N_14175,N_10546,N_10198);
or U14176 (N_14176,N_8843,N_10091);
xnor U14177 (N_14177,N_9762,N_9801);
nor U14178 (N_14178,N_11886,N_10606);
nand U14179 (N_14179,N_9255,N_8814);
nor U14180 (N_14180,N_11544,N_10476);
xnor U14181 (N_14181,N_10255,N_11198);
nor U14182 (N_14182,N_10050,N_9091);
nor U14183 (N_14183,N_9358,N_10899);
xnor U14184 (N_14184,N_8676,N_8108);
or U14185 (N_14185,N_10163,N_11590);
and U14186 (N_14186,N_9652,N_11277);
and U14187 (N_14187,N_9025,N_9185);
or U14188 (N_14188,N_11033,N_11070);
and U14189 (N_14189,N_9394,N_9581);
nor U14190 (N_14190,N_10781,N_9508);
nor U14191 (N_14191,N_8706,N_9441);
nand U14192 (N_14192,N_11576,N_8611);
nand U14193 (N_14193,N_8943,N_10927);
nand U14194 (N_14194,N_9186,N_8874);
nor U14195 (N_14195,N_8601,N_8881);
or U14196 (N_14196,N_10632,N_11013);
xor U14197 (N_14197,N_8431,N_10173);
nand U14198 (N_14198,N_11829,N_8838);
nand U14199 (N_14199,N_11555,N_8846);
xnor U14200 (N_14200,N_11064,N_9668);
nand U14201 (N_14201,N_11210,N_8629);
nand U14202 (N_14202,N_10965,N_11680);
nand U14203 (N_14203,N_8281,N_11746);
xnor U14204 (N_14204,N_9407,N_8043);
and U14205 (N_14205,N_11250,N_8309);
and U14206 (N_14206,N_11042,N_11316);
or U14207 (N_14207,N_10445,N_8473);
and U14208 (N_14208,N_8654,N_9036);
nor U14209 (N_14209,N_11551,N_9750);
nand U14210 (N_14210,N_9342,N_11973);
nor U14211 (N_14211,N_8206,N_10829);
nand U14212 (N_14212,N_10596,N_11877);
or U14213 (N_14213,N_9790,N_10619);
or U14214 (N_14214,N_9562,N_8074);
nand U14215 (N_14215,N_10436,N_9710);
xor U14216 (N_14216,N_11603,N_8745);
nand U14217 (N_14217,N_11290,N_10298);
nor U14218 (N_14218,N_9729,N_9827);
and U14219 (N_14219,N_10127,N_11783);
and U14220 (N_14220,N_11988,N_10607);
or U14221 (N_14221,N_10475,N_8298);
and U14222 (N_14222,N_8686,N_8773);
nor U14223 (N_14223,N_9676,N_8588);
or U14224 (N_14224,N_11894,N_11562);
nor U14225 (N_14225,N_9807,N_8214);
and U14226 (N_14226,N_11453,N_9156);
nand U14227 (N_14227,N_8293,N_8285);
nor U14228 (N_14228,N_10677,N_11841);
nor U14229 (N_14229,N_11582,N_11471);
nor U14230 (N_14230,N_11967,N_11197);
nand U14231 (N_14231,N_11057,N_10999);
nand U14232 (N_14232,N_8601,N_10153);
nand U14233 (N_14233,N_9447,N_8965);
xnor U14234 (N_14234,N_9688,N_11509);
nor U14235 (N_14235,N_11510,N_8217);
nor U14236 (N_14236,N_11349,N_9791);
nor U14237 (N_14237,N_8128,N_11750);
nor U14238 (N_14238,N_11275,N_9276);
nand U14239 (N_14239,N_11430,N_10129);
nor U14240 (N_14240,N_10892,N_9707);
nand U14241 (N_14241,N_8530,N_10598);
nor U14242 (N_14242,N_11483,N_9948);
and U14243 (N_14243,N_11724,N_8327);
nand U14244 (N_14244,N_8924,N_11905);
or U14245 (N_14245,N_10521,N_8224);
nand U14246 (N_14246,N_11908,N_10631);
nand U14247 (N_14247,N_8071,N_11447);
nor U14248 (N_14248,N_11837,N_11822);
xnor U14249 (N_14249,N_10224,N_8068);
xor U14250 (N_14250,N_8651,N_10465);
and U14251 (N_14251,N_9589,N_11932);
nor U14252 (N_14252,N_10244,N_9351);
nand U14253 (N_14253,N_10382,N_8409);
xor U14254 (N_14254,N_11204,N_11775);
and U14255 (N_14255,N_9499,N_10490);
nor U14256 (N_14256,N_11653,N_9376);
nor U14257 (N_14257,N_9061,N_9956);
nand U14258 (N_14258,N_9535,N_10217);
nor U14259 (N_14259,N_10008,N_9938);
nand U14260 (N_14260,N_11258,N_10017);
and U14261 (N_14261,N_11773,N_11283);
or U14262 (N_14262,N_10021,N_10428);
nor U14263 (N_14263,N_11478,N_11201);
xor U14264 (N_14264,N_11671,N_8859);
nand U14265 (N_14265,N_10799,N_8697);
nor U14266 (N_14266,N_10074,N_9220);
or U14267 (N_14267,N_8284,N_8978);
and U14268 (N_14268,N_10514,N_10808);
and U14269 (N_14269,N_10903,N_8739);
and U14270 (N_14270,N_8144,N_8224);
nand U14271 (N_14271,N_8124,N_8678);
nor U14272 (N_14272,N_11122,N_9241);
or U14273 (N_14273,N_9523,N_9745);
or U14274 (N_14274,N_11698,N_9522);
nor U14275 (N_14275,N_8219,N_11721);
and U14276 (N_14276,N_10531,N_10580);
and U14277 (N_14277,N_9060,N_8022);
nor U14278 (N_14278,N_9641,N_10744);
and U14279 (N_14279,N_11272,N_8818);
xnor U14280 (N_14280,N_9205,N_11111);
nand U14281 (N_14281,N_8925,N_8487);
and U14282 (N_14282,N_11256,N_8541);
xnor U14283 (N_14283,N_9584,N_11507);
nand U14284 (N_14284,N_11767,N_11224);
nor U14285 (N_14285,N_10956,N_9106);
and U14286 (N_14286,N_10214,N_11827);
nor U14287 (N_14287,N_9290,N_11467);
or U14288 (N_14288,N_10249,N_10046);
nor U14289 (N_14289,N_11694,N_10301);
nand U14290 (N_14290,N_9556,N_11771);
nor U14291 (N_14291,N_9731,N_11129);
nor U14292 (N_14292,N_10907,N_11770);
xor U14293 (N_14293,N_8713,N_8083);
xnor U14294 (N_14294,N_9192,N_9686);
nand U14295 (N_14295,N_11898,N_10341);
and U14296 (N_14296,N_10234,N_10082);
nand U14297 (N_14297,N_8375,N_8578);
nand U14298 (N_14298,N_8575,N_9716);
and U14299 (N_14299,N_10323,N_10519);
or U14300 (N_14300,N_11121,N_8228);
and U14301 (N_14301,N_8668,N_9753);
nand U14302 (N_14302,N_8729,N_11765);
xor U14303 (N_14303,N_9782,N_11900);
nand U14304 (N_14304,N_10821,N_11708);
and U14305 (N_14305,N_11336,N_9542);
nor U14306 (N_14306,N_8821,N_10519);
nand U14307 (N_14307,N_11052,N_9597);
or U14308 (N_14308,N_10902,N_9814);
nand U14309 (N_14309,N_8725,N_10448);
xnor U14310 (N_14310,N_8460,N_8038);
or U14311 (N_14311,N_8635,N_9174);
or U14312 (N_14312,N_9270,N_10451);
or U14313 (N_14313,N_11983,N_9064);
or U14314 (N_14314,N_9920,N_10319);
or U14315 (N_14315,N_9016,N_10046);
and U14316 (N_14316,N_8363,N_8496);
or U14317 (N_14317,N_10709,N_8436);
nor U14318 (N_14318,N_10643,N_10699);
or U14319 (N_14319,N_10645,N_11396);
or U14320 (N_14320,N_11993,N_8600);
nor U14321 (N_14321,N_8687,N_11427);
nand U14322 (N_14322,N_10707,N_8530);
and U14323 (N_14323,N_10728,N_8001);
nor U14324 (N_14324,N_11785,N_9415);
and U14325 (N_14325,N_8130,N_11993);
or U14326 (N_14326,N_10360,N_10793);
and U14327 (N_14327,N_8106,N_9885);
xnor U14328 (N_14328,N_10372,N_10203);
nor U14329 (N_14329,N_9480,N_10473);
nor U14330 (N_14330,N_11988,N_11617);
nand U14331 (N_14331,N_10551,N_11619);
nor U14332 (N_14332,N_11184,N_9431);
or U14333 (N_14333,N_9124,N_11325);
nand U14334 (N_14334,N_9601,N_11838);
and U14335 (N_14335,N_10899,N_11082);
nor U14336 (N_14336,N_8251,N_8926);
or U14337 (N_14337,N_11824,N_8277);
nand U14338 (N_14338,N_10872,N_10437);
and U14339 (N_14339,N_10328,N_10227);
and U14340 (N_14340,N_9253,N_9104);
and U14341 (N_14341,N_10472,N_9961);
and U14342 (N_14342,N_11587,N_8432);
or U14343 (N_14343,N_11496,N_9435);
and U14344 (N_14344,N_10362,N_11552);
or U14345 (N_14345,N_11243,N_10251);
or U14346 (N_14346,N_8461,N_9956);
xnor U14347 (N_14347,N_9729,N_8644);
and U14348 (N_14348,N_9512,N_10896);
nor U14349 (N_14349,N_8263,N_11131);
and U14350 (N_14350,N_11690,N_10673);
nand U14351 (N_14351,N_10836,N_9156);
nor U14352 (N_14352,N_8405,N_9686);
and U14353 (N_14353,N_9350,N_8691);
or U14354 (N_14354,N_9180,N_9779);
nand U14355 (N_14355,N_10018,N_10789);
or U14356 (N_14356,N_9672,N_11852);
nor U14357 (N_14357,N_10800,N_10701);
nand U14358 (N_14358,N_8028,N_10069);
or U14359 (N_14359,N_8383,N_8561);
and U14360 (N_14360,N_8500,N_10848);
nor U14361 (N_14361,N_9841,N_9941);
nand U14362 (N_14362,N_10814,N_11509);
nand U14363 (N_14363,N_11952,N_10259);
nor U14364 (N_14364,N_9347,N_10818);
or U14365 (N_14365,N_8376,N_8909);
and U14366 (N_14366,N_10475,N_8648);
nand U14367 (N_14367,N_11750,N_10477);
nand U14368 (N_14368,N_11759,N_8589);
nand U14369 (N_14369,N_11115,N_11168);
and U14370 (N_14370,N_9462,N_8718);
nand U14371 (N_14371,N_8682,N_10213);
nand U14372 (N_14372,N_10363,N_8421);
or U14373 (N_14373,N_8089,N_8368);
nand U14374 (N_14374,N_9324,N_9140);
and U14375 (N_14375,N_11872,N_9574);
or U14376 (N_14376,N_11143,N_8050);
nand U14377 (N_14377,N_8748,N_9452);
and U14378 (N_14378,N_8049,N_10948);
nor U14379 (N_14379,N_11536,N_11299);
nand U14380 (N_14380,N_11126,N_11948);
nor U14381 (N_14381,N_11796,N_8663);
or U14382 (N_14382,N_9398,N_11583);
nor U14383 (N_14383,N_9193,N_8955);
or U14384 (N_14384,N_8883,N_8238);
nor U14385 (N_14385,N_10504,N_8676);
xor U14386 (N_14386,N_8968,N_8487);
nand U14387 (N_14387,N_8373,N_8839);
nand U14388 (N_14388,N_9888,N_11481);
nand U14389 (N_14389,N_11893,N_8203);
or U14390 (N_14390,N_10596,N_9559);
and U14391 (N_14391,N_11358,N_11270);
xor U14392 (N_14392,N_8124,N_11850);
xnor U14393 (N_14393,N_9073,N_11648);
or U14394 (N_14394,N_9052,N_10886);
or U14395 (N_14395,N_10055,N_8921);
nand U14396 (N_14396,N_10876,N_8681);
or U14397 (N_14397,N_9101,N_10642);
or U14398 (N_14398,N_10121,N_11780);
and U14399 (N_14399,N_11930,N_11338);
nand U14400 (N_14400,N_9534,N_10309);
or U14401 (N_14401,N_11732,N_8143);
and U14402 (N_14402,N_9898,N_9989);
or U14403 (N_14403,N_8551,N_9252);
and U14404 (N_14404,N_9677,N_10141);
nor U14405 (N_14405,N_8692,N_11449);
and U14406 (N_14406,N_10164,N_11069);
and U14407 (N_14407,N_10039,N_9046);
nor U14408 (N_14408,N_9798,N_10764);
and U14409 (N_14409,N_8194,N_10426);
or U14410 (N_14410,N_8272,N_8878);
and U14411 (N_14411,N_8235,N_10714);
xnor U14412 (N_14412,N_10953,N_8512);
nand U14413 (N_14413,N_10399,N_9006);
nor U14414 (N_14414,N_10338,N_10280);
nor U14415 (N_14415,N_10227,N_8701);
or U14416 (N_14416,N_10796,N_8247);
and U14417 (N_14417,N_9098,N_11610);
and U14418 (N_14418,N_9322,N_8066);
nand U14419 (N_14419,N_9174,N_9499);
nand U14420 (N_14420,N_10176,N_10504);
or U14421 (N_14421,N_10804,N_9592);
and U14422 (N_14422,N_10207,N_8707);
nand U14423 (N_14423,N_9677,N_10414);
and U14424 (N_14424,N_9009,N_8964);
nand U14425 (N_14425,N_10634,N_9416);
and U14426 (N_14426,N_10189,N_10526);
or U14427 (N_14427,N_8942,N_11776);
xor U14428 (N_14428,N_10870,N_11356);
or U14429 (N_14429,N_11652,N_9032);
nor U14430 (N_14430,N_8159,N_10907);
nor U14431 (N_14431,N_10439,N_8369);
nor U14432 (N_14432,N_9503,N_8017);
or U14433 (N_14433,N_8912,N_9042);
and U14434 (N_14434,N_10069,N_11751);
or U14435 (N_14435,N_11040,N_9465);
and U14436 (N_14436,N_9285,N_10076);
xnor U14437 (N_14437,N_11995,N_8480);
and U14438 (N_14438,N_8840,N_9981);
nor U14439 (N_14439,N_11171,N_11610);
xor U14440 (N_14440,N_10239,N_11867);
nand U14441 (N_14441,N_9812,N_9406);
nand U14442 (N_14442,N_10823,N_9084);
nor U14443 (N_14443,N_11174,N_10973);
and U14444 (N_14444,N_11244,N_8032);
nand U14445 (N_14445,N_10524,N_9867);
and U14446 (N_14446,N_8096,N_10934);
nand U14447 (N_14447,N_11386,N_9145);
and U14448 (N_14448,N_11717,N_9754);
xnor U14449 (N_14449,N_8220,N_9857);
nor U14450 (N_14450,N_9571,N_10816);
xor U14451 (N_14451,N_11954,N_10375);
and U14452 (N_14452,N_11079,N_8841);
and U14453 (N_14453,N_10124,N_11592);
nor U14454 (N_14454,N_10405,N_10636);
and U14455 (N_14455,N_11686,N_8420);
nor U14456 (N_14456,N_11122,N_11808);
or U14457 (N_14457,N_11333,N_10591);
xor U14458 (N_14458,N_10853,N_10908);
or U14459 (N_14459,N_10614,N_8495);
and U14460 (N_14460,N_8656,N_8941);
nand U14461 (N_14461,N_9292,N_11578);
and U14462 (N_14462,N_11135,N_11780);
nor U14463 (N_14463,N_11079,N_9200);
nand U14464 (N_14464,N_8221,N_11424);
and U14465 (N_14465,N_10914,N_10800);
nor U14466 (N_14466,N_10210,N_9480);
or U14467 (N_14467,N_10048,N_8852);
and U14468 (N_14468,N_8611,N_10717);
nand U14469 (N_14469,N_8650,N_11542);
nor U14470 (N_14470,N_9789,N_11562);
nand U14471 (N_14471,N_9577,N_8615);
xnor U14472 (N_14472,N_9171,N_10139);
or U14473 (N_14473,N_10168,N_10589);
or U14474 (N_14474,N_10195,N_11942);
or U14475 (N_14475,N_9452,N_11505);
or U14476 (N_14476,N_9291,N_10598);
and U14477 (N_14477,N_9343,N_11628);
nor U14478 (N_14478,N_10008,N_8661);
xnor U14479 (N_14479,N_10346,N_11421);
and U14480 (N_14480,N_11386,N_10757);
nor U14481 (N_14481,N_10719,N_8448);
or U14482 (N_14482,N_11198,N_9692);
xor U14483 (N_14483,N_11056,N_9703);
nor U14484 (N_14484,N_9763,N_10323);
or U14485 (N_14485,N_11617,N_8961);
or U14486 (N_14486,N_11823,N_9794);
nand U14487 (N_14487,N_9025,N_10047);
nor U14488 (N_14488,N_9683,N_8507);
nor U14489 (N_14489,N_8789,N_11662);
or U14490 (N_14490,N_9101,N_11548);
nor U14491 (N_14491,N_10258,N_10719);
or U14492 (N_14492,N_8023,N_11308);
or U14493 (N_14493,N_8606,N_9875);
or U14494 (N_14494,N_9742,N_10069);
nand U14495 (N_14495,N_8775,N_9127);
or U14496 (N_14496,N_9596,N_8533);
nor U14497 (N_14497,N_8979,N_9894);
nor U14498 (N_14498,N_11148,N_9474);
nand U14499 (N_14499,N_9808,N_8537);
nand U14500 (N_14500,N_11653,N_8307);
nor U14501 (N_14501,N_10882,N_8515);
and U14502 (N_14502,N_8633,N_10931);
nor U14503 (N_14503,N_8815,N_10467);
or U14504 (N_14504,N_8801,N_9459);
nand U14505 (N_14505,N_11194,N_11475);
and U14506 (N_14506,N_9532,N_8797);
nor U14507 (N_14507,N_9116,N_11062);
xnor U14508 (N_14508,N_8875,N_11943);
nand U14509 (N_14509,N_10989,N_10325);
nand U14510 (N_14510,N_8269,N_10330);
and U14511 (N_14511,N_9113,N_11073);
nor U14512 (N_14512,N_8154,N_8758);
and U14513 (N_14513,N_10905,N_10535);
nand U14514 (N_14514,N_9443,N_9227);
nand U14515 (N_14515,N_10599,N_9888);
or U14516 (N_14516,N_9130,N_10700);
or U14517 (N_14517,N_8129,N_8500);
xnor U14518 (N_14518,N_11305,N_11588);
or U14519 (N_14519,N_11013,N_8515);
or U14520 (N_14520,N_8421,N_11355);
nor U14521 (N_14521,N_10393,N_10977);
and U14522 (N_14522,N_10861,N_8759);
nor U14523 (N_14523,N_8211,N_9584);
xnor U14524 (N_14524,N_8400,N_9227);
and U14525 (N_14525,N_10113,N_10972);
xnor U14526 (N_14526,N_8690,N_8079);
nand U14527 (N_14527,N_11429,N_10404);
or U14528 (N_14528,N_10585,N_8082);
xor U14529 (N_14529,N_11366,N_9121);
and U14530 (N_14530,N_11513,N_8634);
nand U14531 (N_14531,N_10746,N_11257);
nand U14532 (N_14532,N_9300,N_9608);
xnor U14533 (N_14533,N_8202,N_11870);
nand U14534 (N_14534,N_10552,N_11017);
or U14535 (N_14535,N_11439,N_10843);
or U14536 (N_14536,N_11092,N_11562);
and U14537 (N_14537,N_8672,N_8442);
nand U14538 (N_14538,N_8616,N_9800);
nor U14539 (N_14539,N_8376,N_9263);
and U14540 (N_14540,N_11081,N_9795);
xor U14541 (N_14541,N_9367,N_8549);
or U14542 (N_14542,N_10822,N_8893);
or U14543 (N_14543,N_11320,N_10853);
xnor U14544 (N_14544,N_11684,N_9090);
or U14545 (N_14545,N_11392,N_10677);
or U14546 (N_14546,N_10514,N_9307);
and U14547 (N_14547,N_10413,N_10715);
xnor U14548 (N_14548,N_11265,N_8661);
nand U14549 (N_14549,N_11824,N_10148);
nor U14550 (N_14550,N_11755,N_11300);
or U14551 (N_14551,N_9969,N_9116);
nand U14552 (N_14552,N_10549,N_8729);
or U14553 (N_14553,N_10840,N_9521);
nor U14554 (N_14554,N_9871,N_10607);
xnor U14555 (N_14555,N_10788,N_11910);
or U14556 (N_14556,N_9848,N_9831);
nor U14557 (N_14557,N_11720,N_10283);
and U14558 (N_14558,N_8977,N_10755);
nand U14559 (N_14559,N_10991,N_11811);
or U14560 (N_14560,N_9277,N_11633);
xor U14561 (N_14561,N_11704,N_8090);
nand U14562 (N_14562,N_8394,N_9880);
nor U14563 (N_14563,N_10616,N_10656);
nand U14564 (N_14564,N_10363,N_8232);
nor U14565 (N_14565,N_9958,N_11355);
or U14566 (N_14566,N_8173,N_8036);
nor U14567 (N_14567,N_11814,N_10662);
and U14568 (N_14568,N_11200,N_10082);
nor U14569 (N_14569,N_8736,N_10856);
and U14570 (N_14570,N_9768,N_10191);
nor U14571 (N_14571,N_9784,N_11641);
nand U14572 (N_14572,N_10846,N_9721);
nand U14573 (N_14573,N_10746,N_11587);
or U14574 (N_14574,N_11932,N_11925);
nand U14575 (N_14575,N_10840,N_9886);
nor U14576 (N_14576,N_11725,N_8738);
or U14577 (N_14577,N_9996,N_10677);
nand U14578 (N_14578,N_10218,N_10133);
nor U14579 (N_14579,N_11221,N_10632);
nor U14580 (N_14580,N_9242,N_10073);
nor U14581 (N_14581,N_9094,N_9811);
or U14582 (N_14582,N_10882,N_11606);
nor U14583 (N_14583,N_11685,N_9698);
nand U14584 (N_14584,N_8075,N_10443);
and U14585 (N_14585,N_9247,N_9108);
and U14586 (N_14586,N_11307,N_8429);
nand U14587 (N_14587,N_8912,N_8958);
or U14588 (N_14588,N_9395,N_9374);
or U14589 (N_14589,N_11473,N_10000);
xnor U14590 (N_14590,N_10072,N_10164);
nand U14591 (N_14591,N_11283,N_11399);
or U14592 (N_14592,N_8482,N_9988);
nor U14593 (N_14593,N_11845,N_11792);
and U14594 (N_14594,N_10693,N_11247);
nand U14595 (N_14595,N_9078,N_9104);
nand U14596 (N_14596,N_11852,N_10869);
or U14597 (N_14597,N_9497,N_11814);
xnor U14598 (N_14598,N_8567,N_9681);
nor U14599 (N_14599,N_11519,N_10860);
nand U14600 (N_14600,N_8990,N_9843);
xnor U14601 (N_14601,N_11469,N_10517);
nor U14602 (N_14602,N_9442,N_11858);
and U14603 (N_14603,N_8379,N_11783);
and U14604 (N_14604,N_8841,N_8719);
or U14605 (N_14605,N_11007,N_8968);
or U14606 (N_14606,N_10121,N_9950);
and U14607 (N_14607,N_10159,N_11085);
nand U14608 (N_14608,N_8520,N_11256);
xor U14609 (N_14609,N_10157,N_11886);
xnor U14610 (N_14610,N_8727,N_11971);
nor U14611 (N_14611,N_10074,N_10107);
or U14612 (N_14612,N_10724,N_10554);
nand U14613 (N_14613,N_9294,N_10467);
or U14614 (N_14614,N_11969,N_11195);
or U14615 (N_14615,N_11516,N_8059);
nor U14616 (N_14616,N_11184,N_11248);
xor U14617 (N_14617,N_8021,N_8933);
and U14618 (N_14618,N_10413,N_10754);
and U14619 (N_14619,N_11627,N_11135);
nor U14620 (N_14620,N_8103,N_9799);
xor U14621 (N_14621,N_8489,N_8281);
nor U14622 (N_14622,N_11874,N_8723);
nand U14623 (N_14623,N_8863,N_10167);
nand U14624 (N_14624,N_8058,N_8477);
nand U14625 (N_14625,N_10994,N_9031);
and U14626 (N_14626,N_8239,N_11218);
nor U14627 (N_14627,N_9099,N_11814);
nand U14628 (N_14628,N_9497,N_10304);
or U14629 (N_14629,N_11162,N_9203);
and U14630 (N_14630,N_11901,N_11428);
and U14631 (N_14631,N_9168,N_11460);
or U14632 (N_14632,N_8747,N_8596);
or U14633 (N_14633,N_8714,N_8375);
and U14634 (N_14634,N_11966,N_9502);
and U14635 (N_14635,N_8970,N_11404);
nor U14636 (N_14636,N_9160,N_8100);
nor U14637 (N_14637,N_8762,N_10821);
nor U14638 (N_14638,N_10153,N_10665);
xor U14639 (N_14639,N_10693,N_9179);
or U14640 (N_14640,N_10439,N_10945);
nand U14641 (N_14641,N_11348,N_8390);
or U14642 (N_14642,N_9242,N_11755);
nand U14643 (N_14643,N_9749,N_9647);
nand U14644 (N_14644,N_9765,N_11944);
nand U14645 (N_14645,N_10094,N_10591);
or U14646 (N_14646,N_9817,N_8715);
and U14647 (N_14647,N_11905,N_8237);
xnor U14648 (N_14648,N_8641,N_10387);
nor U14649 (N_14649,N_9125,N_10121);
or U14650 (N_14650,N_10672,N_10287);
and U14651 (N_14651,N_10344,N_9818);
nor U14652 (N_14652,N_11153,N_11096);
or U14653 (N_14653,N_9637,N_9354);
and U14654 (N_14654,N_9644,N_11738);
xnor U14655 (N_14655,N_9847,N_10482);
or U14656 (N_14656,N_9056,N_8832);
nand U14657 (N_14657,N_11631,N_8691);
nand U14658 (N_14658,N_11386,N_8505);
or U14659 (N_14659,N_10585,N_11143);
xor U14660 (N_14660,N_11584,N_11734);
and U14661 (N_14661,N_10470,N_10048);
or U14662 (N_14662,N_8801,N_10269);
or U14663 (N_14663,N_9177,N_8325);
and U14664 (N_14664,N_8919,N_8872);
or U14665 (N_14665,N_8976,N_11024);
and U14666 (N_14666,N_9485,N_10022);
and U14667 (N_14667,N_11601,N_9158);
xnor U14668 (N_14668,N_9899,N_10063);
and U14669 (N_14669,N_8318,N_10140);
nand U14670 (N_14670,N_9528,N_11904);
nand U14671 (N_14671,N_11952,N_11490);
and U14672 (N_14672,N_10243,N_10525);
or U14673 (N_14673,N_11038,N_9326);
nor U14674 (N_14674,N_8075,N_10094);
or U14675 (N_14675,N_8501,N_8562);
and U14676 (N_14676,N_9434,N_11295);
nor U14677 (N_14677,N_10910,N_11685);
and U14678 (N_14678,N_9465,N_11709);
and U14679 (N_14679,N_9671,N_8507);
xor U14680 (N_14680,N_8144,N_10053);
nor U14681 (N_14681,N_10118,N_10662);
nand U14682 (N_14682,N_8654,N_8927);
or U14683 (N_14683,N_10452,N_9344);
nor U14684 (N_14684,N_11362,N_9406);
nand U14685 (N_14685,N_9278,N_11916);
nand U14686 (N_14686,N_10293,N_8317);
and U14687 (N_14687,N_11354,N_10330);
nand U14688 (N_14688,N_11082,N_10380);
nand U14689 (N_14689,N_11959,N_9278);
and U14690 (N_14690,N_8963,N_10085);
nand U14691 (N_14691,N_11973,N_11767);
nand U14692 (N_14692,N_11198,N_11082);
nor U14693 (N_14693,N_9211,N_8555);
nand U14694 (N_14694,N_9344,N_8040);
xor U14695 (N_14695,N_9648,N_9730);
and U14696 (N_14696,N_9764,N_8658);
nor U14697 (N_14697,N_9483,N_11683);
nand U14698 (N_14698,N_9301,N_10740);
and U14699 (N_14699,N_10740,N_11864);
and U14700 (N_14700,N_9617,N_9138);
or U14701 (N_14701,N_10899,N_8446);
and U14702 (N_14702,N_8226,N_10275);
and U14703 (N_14703,N_10270,N_10481);
nand U14704 (N_14704,N_9974,N_9257);
nor U14705 (N_14705,N_11299,N_10192);
and U14706 (N_14706,N_11942,N_9192);
or U14707 (N_14707,N_10041,N_10891);
nand U14708 (N_14708,N_11073,N_9944);
nand U14709 (N_14709,N_11231,N_9551);
nand U14710 (N_14710,N_11613,N_8870);
nand U14711 (N_14711,N_10232,N_9893);
nor U14712 (N_14712,N_8732,N_10241);
and U14713 (N_14713,N_9157,N_8252);
and U14714 (N_14714,N_11711,N_11062);
xnor U14715 (N_14715,N_8513,N_11716);
nand U14716 (N_14716,N_11799,N_11429);
nor U14717 (N_14717,N_10015,N_9495);
or U14718 (N_14718,N_10616,N_9371);
nor U14719 (N_14719,N_10476,N_9353);
and U14720 (N_14720,N_11775,N_9809);
nor U14721 (N_14721,N_8853,N_8386);
nand U14722 (N_14722,N_10349,N_11162);
nor U14723 (N_14723,N_11745,N_11566);
and U14724 (N_14724,N_9241,N_9190);
or U14725 (N_14725,N_10651,N_11732);
nand U14726 (N_14726,N_8017,N_10307);
nor U14727 (N_14727,N_10226,N_9010);
nor U14728 (N_14728,N_11935,N_8042);
nor U14729 (N_14729,N_11219,N_8130);
nand U14730 (N_14730,N_9079,N_11089);
and U14731 (N_14731,N_9268,N_8050);
and U14732 (N_14732,N_10060,N_9230);
and U14733 (N_14733,N_8749,N_11662);
xor U14734 (N_14734,N_9739,N_9735);
and U14735 (N_14735,N_9271,N_10045);
nor U14736 (N_14736,N_10137,N_9590);
nor U14737 (N_14737,N_8215,N_8021);
nor U14738 (N_14738,N_11037,N_8611);
and U14739 (N_14739,N_10550,N_9556);
nor U14740 (N_14740,N_10472,N_8570);
nor U14741 (N_14741,N_9990,N_11913);
and U14742 (N_14742,N_11827,N_10134);
and U14743 (N_14743,N_9965,N_10354);
and U14744 (N_14744,N_10801,N_10399);
or U14745 (N_14745,N_8028,N_9454);
and U14746 (N_14746,N_11310,N_8192);
or U14747 (N_14747,N_10162,N_10630);
nand U14748 (N_14748,N_10322,N_10579);
or U14749 (N_14749,N_8494,N_8776);
nand U14750 (N_14750,N_8262,N_9174);
and U14751 (N_14751,N_8023,N_9069);
and U14752 (N_14752,N_11037,N_11867);
xor U14753 (N_14753,N_10230,N_11099);
nand U14754 (N_14754,N_9649,N_8299);
nor U14755 (N_14755,N_10764,N_9836);
and U14756 (N_14756,N_10062,N_9577);
xnor U14757 (N_14757,N_8350,N_11974);
or U14758 (N_14758,N_9675,N_8016);
nor U14759 (N_14759,N_9101,N_9456);
nor U14760 (N_14760,N_8065,N_11898);
xor U14761 (N_14761,N_10180,N_11753);
and U14762 (N_14762,N_9347,N_11236);
or U14763 (N_14763,N_11802,N_10360);
or U14764 (N_14764,N_11941,N_11268);
nand U14765 (N_14765,N_8169,N_8261);
nor U14766 (N_14766,N_11512,N_8122);
and U14767 (N_14767,N_11470,N_8671);
nor U14768 (N_14768,N_10441,N_9133);
nor U14769 (N_14769,N_8025,N_11878);
nor U14770 (N_14770,N_8820,N_11286);
or U14771 (N_14771,N_8458,N_9361);
nand U14772 (N_14772,N_8108,N_11658);
nor U14773 (N_14773,N_11245,N_10924);
nor U14774 (N_14774,N_11622,N_8857);
nor U14775 (N_14775,N_11168,N_11692);
and U14776 (N_14776,N_9037,N_11548);
nor U14777 (N_14777,N_8297,N_8500);
nand U14778 (N_14778,N_8103,N_11879);
or U14779 (N_14779,N_11141,N_9984);
nand U14780 (N_14780,N_10224,N_10783);
and U14781 (N_14781,N_11939,N_10945);
and U14782 (N_14782,N_9826,N_9032);
xnor U14783 (N_14783,N_11726,N_8132);
xnor U14784 (N_14784,N_10886,N_11276);
nand U14785 (N_14785,N_10724,N_10638);
and U14786 (N_14786,N_9944,N_9688);
and U14787 (N_14787,N_10928,N_8665);
xnor U14788 (N_14788,N_11542,N_10963);
nand U14789 (N_14789,N_8723,N_8964);
nand U14790 (N_14790,N_8323,N_9798);
nor U14791 (N_14791,N_10298,N_8587);
nand U14792 (N_14792,N_10992,N_8857);
nor U14793 (N_14793,N_11092,N_10980);
and U14794 (N_14794,N_11290,N_9539);
or U14795 (N_14795,N_10586,N_10451);
or U14796 (N_14796,N_10553,N_9841);
or U14797 (N_14797,N_9005,N_10681);
and U14798 (N_14798,N_9576,N_11965);
and U14799 (N_14799,N_10896,N_10761);
and U14800 (N_14800,N_10977,N_9946);
xnor U14801 (N_14801,N_10710,N_11958);
nand U14802 (N_14802,N_11924,N_9877);
nor U14803 (N_14803,N_8254,N_9377);
and U14804 (N_14804,N_9297,N_9356);
xnor U14805 (N_14805,N_9852,N_9936);
and U14806 (N_14806,N_9830,N_9586);
nor U14807 (N_14807,N_9259,N_9366);
nand U14808 (N_14808,N_10076,N_11561);
or U14809 (N_14809,N_9119,N_11522);
nand U14810 (N_14810,N_9624,N_8127);
nand U14811 (N_14811,N_11309,N_9314);
nand U14812 (N_14812,N_11646,N_9320);
nand U14813 (N_14813,N_9563,N_9996);
nand U14814 (N_14814,N_8391,N_8980);
or U14815 (N_14815,N_8128,N_9569);
or U14816 (N_14816,N_8395,N_8292);
nand U14817 (N_14817,N_8594,N_11286);
xnor U14818 (N_14818,N_11538,N_11475);
or U14819 (N_14819,N_8212,N_11238);
or U14820 (N_14820,N_10565,N_11660);
nor U14821 (N_14821,N_10913,N_8164);
xor U14822 (N_14822,N_9946,N_11462);
nor U14823 (N_14823,N_9726,N_9258);
or U14824 (N_14824,N_8419,N_9503);
or U14825 (N_14825,N_9685,N_10348);
and U14826 (N_14826,N_10113,N_10200);
or U14827 (N_14827,N_8516,N_10170);
or U14828 (N_14828,N_9056,N_11089);
nor U14829 (N_14829,N_9856,N_11855);
or U14830 (N_14830,N_8364,N_11731);
nor U14831 (N_14831,N_9609,N_9691);
or U14832 (N_14832,N_9990,N_10871);
and U14833 (N_14833,N_9197,N_11843);
and U14834 (N_14834,N_9789,N_9113);
or U14835 (N_14835,N_11110,N_9178);
xor U14836 (N_14836,N_10707,N_10839);
or U14837 (N_14837,N_10326,N_8009);
nor U14838 (N_14838,N_9661,N_10239);
and U14839 (N_14839,N_9994,N_9935);
nand U14840 (N_14840,N_8537,N_9918);
or U14841 (N_14841,N_10079,N_11521);
nand U14842 (N_14842,N_9590,N_8000);
xor U14843 (N_14843,N_8800,N_11678);
xor U14844 (N_14844,N_9547,N_11266);
and U14845 (N_14845,N_10225,N_9678);
nor U14846 (N_14846,N_8511,N_8929);
nand U14847 (N_14847,N_9047,N_10171);
or U14848 (N_14848,N_8509,N_10898);
nand U14849 (N_14849,N_11688,N_11063);
nand U14850 (N_14850,N_8831,N_10802);
xor U14851 (N_14851,N_8569,N_9991);
nor U14852 (N_14852,N_11379,N_8866);
and U14853 (N_14853,N_8555,N_10156);
nor U14854 (N_14854,N_10994,N_9103);
or U14855 (N_14855,N_11441,N_9909);
nand U14856 (N_14856,N_10384,N_11140);
nor U14857 (N_14857,N_11367,N_8761);
nand U14858 (N_14858,N_11676,N_8839);
nand U14859 (N_14859,N_11392,N_8661);
xor U14860 (N_14860,N_11073,N_10328);
or U14861 (N_14861,N_11511,N_9389);
and U14862 (N_14862,N_8552,N_11464);
nor U14863 (N_14863,N_8690,N_8558);
nand U14864 (N_14864,N_8903,N_9129);
xnor U14865 (N_14865,N_9990,N_8874);
nand U14866 (N_14866,N_10162,N_10547);
nand U14867 (N_14867,N_8450,N_10515);
nor U14868 (N_14868,N_8573,N_10831);
or U14869 (N_14869,N_9645,N_11548);
xor U14870 (N_14870,N_8088,N_8003);
nor U14871 (N_14871,N_8536,N_11320);
and U14872 (N_14872,N_9988,N_10705);
and U14873 (N_14873,N_8043,N_11651);
and U14874 (N_14874,N_10019,N_9746);
and U14875 (N_14875,N_8405,N_11755);
and U14876 (N_14876,N_11420,N_11665);
or U14877 (N_14877,N_10796,N_11819);
nand U14878 (N_14878,N_8033,N_10458);
nand U14879 (N_14879,N_10106,N_9359);
or U14880 (N_14880,N_11594,N_9754);
and U14881 (N_14881,N_10470,N_9060);
and U14882 (N_14882,N_9715,N_9913);
or U14883 (N_14883,N_8329,N_8700);
nand U14884 (N_14884,N_11678,N_10798);
nand U14885 (N_14885,N_10426,N_11003);
and U14886 (N_14886,N_8035,N_11505);
or U14887 (N_14887,N_10148,N_11256);
and U14888 (N_14888,N_9124,N_11869);
or U14889 (N_14889,N_10510,N_10516);
and U14890 (N_14890,N_11470,N_8382);
nand U14891 (N_14891,N_9579,N_8527);
and U14892 (N_14892,N_10463,N_11753);
xor U14893 (N_14893,N_10609,N_10979);
nand U14894 (N_14894,N_11601,N_8742);
nand U14895 (N_14895,N_8277,N_11686);
xor U14896 (N_14896,N_9374,N_10339);
xor U14897 (N_14897,N_9867,N_8497);
nor U14898 (N_14898,N_10435,N_9659);
xnor U14899 (N_14899,N_10534,N_11354);
nand U14900 (N_14900,N_10918,N_8926);
nor U14901 (N_14901,N_10905,N_10746);
nor U14902 (N_14902,N_10459,N_9487);
xor U14903 (N_14903,N_10598,N_8469);
nor U14904 (N_14904,N_11694,N_11396);
nor U14905 (N_14905,N_11428,N_10921);
or U14906 (N_14906,N_8898,N_11799);
and U14907 (N_14907,N_8656,N_10454);
or U14908 (N_14908,N_9084,N_9747);
or U14909 (N_14909,N_9553,N_11404);
nand U14910 (N_14910,N_10264,N_11053);
and U14911 (N_14911,N_8730,N_11246);
or U14912 (N_14912,N_11967,N_10595);
nor U14913 (N_14913,N_9076,N_8499);
or U14914 (N_14914,N_8615,N_10783);
nor U14915 (N_14915,N_11474,N_8801);
or U14916 (N_14916,N_10367,N_10435);
xor U14917 (N_14917,N_11923,N_10436);
nor U14918 (N_14918,N_11250,N_8968);
nor U14919 (N_14919,N_10262,N_9518);
nor U14920 (N_14920,N_8789,N_8573);
nor U14921 (N_14921,N_10149,N_10711);
nor U14922 (N_14922,N_8324,N_11607);
nor U14923 (N_14923,N_9864,N_8867);
and U14924 (N_14924,N_9088,N_9586);
nor U14925 (N_14925,N_9947,N_9730);
xnor U14926 (N_14926,N_11985,N_11129);
xnor U14927 (N_14927,N_9174,N_8877);
nand U14928 (N_14928,N_9773,N_9615);
or U14929 (N_14929,N_10723,N_8044);
or U14930 (N_14930,N_10205,N_9561);
nand U14931 (N_14931,N_11849,N_9248);
and U14932 (N_14932,N_11315,N_9231);
or U14933 (N_14933,N_9918,N_11722);
nand U14934 (N_14934,N_9002,N_9450);
nand U14935 (N_14935,N_8039,N_8474);
or U14936 (N_14936,N_8497,N_10288);
or U14937 (N_14937,N_8541,N_8547);
nor U14938 (N_14938,N_11697,N_10875);
or U14939 (N_14939,N_9131,N_8381);
nand U14940 (N_14940,N_11268,N_10441);
or U14941 (N_14941,N_11874,N_8758);
xnor U14942 (N_14942,N_11679,N_9823);
or U14943 (N_14943,N_11399,N_8303);
or U14944 (N_14944,N_10551,N_9363);
or U14945 (N_14945,N_8389,N_10814);
and U14946 (N_14946,N_11622,N_8097);
and U14947 (N_14947,N_9411,N_9873);
nor U14948 (N_14948,N_11136,N_11168);
or U14949 (N_14949,N_11562,N_9948);
or U14950 (N_14950,N_11758,N_11268);
nand U14951 (N_14951,N_11971,N_9082);
or U14952 (N_14952,N_10692,N_11294);
and U14953 (N_14953,N_11816,N_11910);
nor U14954 (N_14954,N_10450,N_11247);
nand U14955 (N_14955,N_9824,N_11642);
nand U14956 (N_14956,N_10902,N_8968);
or U14957 (N_14957,N_8568,N_10038);
or U14958 (N_14958,N_9236,N_9814);
or U14959 (N_14959,N_10937,N_11446);
nor U14960 (N_14960,N_9004,N_8373);
nand U14961 (N_14961,N_8279,N_9338);
and U14962 (N_14962,N_9745,N_8093);
nand U14963 (N_14963,N_8186,N_8842);
nor U14964 (N_14964,N_11388,N_10393);
or U14965 (N_14965,N_11737,N_11086);
and U14966 (N_14966,N_8193,N_9125);
nand U14967 (N_14967,N_11670,N_8236);
nor U14968 (N_14968,N_10534,N_10450);
or U14969 (N_14969,N_8044,N_8332);
xor U14970 (N_14970,N_9677,N_10125);
xnor U14971 (N_14971,N_10563,N_10836);
or U14972 (N_14972,N_9106,N_11677);
nor U14973 (N_14973,N_9727,N_8580);
xor U14974 (N_14974,N_11948,N_9686);
or U14975 (N_14975,N_9058,N_8950);
and U14976 (N_14976,N_10021,N_10070);
or U14977 (N_14977,N_8461,N_9044);
nor U14978 (N_14978,N_10296,N_9706);
nand U14979 (N_14979,N_8556,N_10594);
nor U14980 (N_14980,N_10026,N_10198);
or U14981 (N_14981,N_11034,N_9517);
nand U14982 (N_14982,N_8604,N_11017);
xnor U14983 (N_14983,N_10765,N_8717);
nor U14984 (N_14984,N_10976,N_11661);
and U14985 (N_14985,N_11527,N_8264);
nand U14986 (N_14986,N_10310,N_8261);
or U14987 (N_14987,N_9140,N_10710);
and U14988 (N_14988,N_9704,N_8455);
xnor U14989 (N_14989,N_8511,N_11191);
or U14990 (N_14990,N_11931,N_11218);
nand U14991 (N_14991,N_10677,N_10878);
nor U14992 (N_14992,N_10227,N_11409);
and U14993 (N_14993,N_10291,N_10630);
and U14994 (N_14994,N_8053,N_9440);
nor U14995 (N_14995,N_11832,N_8821);
and U14996 (N_14996,N_10820,N_11937);
nand U14997 (N_14997,N_11888,N_8780);
and U14998 (N_14998,N_10926,N_9288);
nand U14999 (N_14999,N_11276,N_8245);
or U15000 (N_15000,N_9901,N_11562);
or U15001 (N_15001,N_11330,N_8499);
nand U15002 (N_15002,N_9758,N_10371);
and U15003 (N_15003,N_8173,N_11571);
or U15004 (N_15004,N_11987,N_10660);
nand U15005 (N_15005,N_8733,N_10213);
xor U15006 (N_15006,N_8446,N_11057);
nor U15007 (N_15007,N_10144,N_10245);
and U15008 (N_15008,N_8999,N_10526);
or U15009 (N_15009,N_8891,N_9191);
or U15010 (N_15010,N_11431,N_11309);
or U15011 (N_15011,N_11938,N_9322);
and U15012 (N_15012,N_10871,N_9230);
nor U15013 (N_15013,N_11808,N_9402);
and U15014 (N_15014,N_10843,N_8006);
or U15015 (N_15015,N_10481,N_8100);
xnor U15016 (N_15016,N_8894,N_10927);
or U15017 (N_15017,N_10990,N_9622);
or U15018 (N_15018,N_11759,N_9781);
and U15019 (N_15019,N_9824,N_10633);
xnor U15020 (N_15020,N_8738,N_11764);
or U15021 (N_15021,N_11559,N_11855);
nand U15022 (N_15022,N_8120,N_11661);
nor U15023 (N_15023,N_8385,N_9040);
xnor U15024 (N_15024,N_9773,N_11589);
nor U15025 (N_15025,N_11633,N_9120);
or U15026 (N_15026,N_11343,N_10918);
and U15027 (N_15027,N_11760,N_9675);
xor U15028 (N_15028,N_10669,N_10379);
nor U15029 (N_15029,N_10929,N_8798);
or U15030 (N_15030,N_9539,N_9834);
or U15031 (N_15031,N_8518,N_8069);
nor U15032 (N_15032,N_9751,N_8344);
or U15033 (N_15033,N_8971,N_10497);
and U15034 (N_15034,N_9230,N_9040);
nand U15035 (N_15035,N_11130,N_11847);
nor U15036 (N_15036,N_8426,N_10639);
or U15037 (N_15037,N_11816,N_11206);
xor U15038 (N_15038,N_11954,N_9036);
or U15039 (N_15039,N_9927,N_9632);
nand U15040 (N_15040,N_8116,N_8028);
nand U15041 (N_15041,N_11804,N_8291);
or U15042 (N_15042,N_8361,N_10418);
nand U15043 (N_15043,N_11447,N_10115);
or U15044 (N_15044,N_8050,N_9640);
nand U15045 (N_15045,N_9155,N_8986);
or U15046 (N_15046,N_8038,N_11217);
nand U15047 (N_15047,N_11137,N_8204);
or U15048 (N_15048,N_10643,N_10329);
nand U15049 (N_15049,N_10213,N_10497);
or U15050 (N_15050,N_10647,N_9175);
nand U15051 (N_15051,N_8306,N_11215);
and U15052 (N_15052,N_8752,N_11320);
nor U15053 (N_15053,N_8593,N_9172);
and U15054 (N_15054,N_9982,N_8314);
nand U15055 (N_15055,N_8710,N_10644);
and U15056 (N_15056,N_9814,N_11649);
or U15057 (N_15057,N_10096,N_10300);
nand U15058 (N_15058,N_11120,N_10971);
nand U15059 (N_15059,N_9176,N_8552);
nand U15060 (N_15060,N_11601,N_11221);
or U15061 (N_15061,N_8634,N_9738);
nand U15062 (N_15062,N_8490,N_11929);
and U15063 (N_15063,N_9313,N_10045);
and U15064 (N_15064,N_9210,N_10093);
and U15065 (N_15065,N_10565,N_9151);
nand U15066 (N_15066,N_10680,N_10016);
and U15067 (N_15067,N_9537,N_11700);
nor U15068 (N_15068,N_10275,N_10796);
nor U15069 (N_15069,N_11891,N_8177);
or U15070 (N_15070,N_9907,N_11550);
or U15071 (N_15071,N_11748,N_9521);
nor U15072 (N_15072,N_8188,N_9970);
xor U15073 (N_15073,N_8256,N_8848);
nor U15074 (N_15074,N_11857,N_11822);
nor U15075 (N_15075,N_9132,N_11337);
nor U15076 (N_15076,N_11212,N_10286);
nand U15077 (N_15077,N_10277,N_9987);
or U15078 (N_15078,N_9679,N_10514);
or U15079 (N_15079,N_10739,N_8549);
or U15080 (N_15080,N_9391,N_11326);
nand U15081 (N_15081,N_11805,N_11618);
nand U15082 (N_15082,N_8869,N_9513);
nor U15083 (N_15083,N_9703,N_10326);
nor U15084 (N_15084,N_9688,N_10360);
or U15085 (N_15085,N_9259,N_9660);
nor U15086 (N_15086,N_9088,N_11535);
xnor U15087 (N_15087,N_10627,N_9182);
nand U15088 (N_15088,N_8158,N_8271);
nand U15089 (N_15089,N_8910,N_8959);
and U15090 (N_15090,N_11205,N_8040);
xnor U15091 (N_15091,N_11315,N_8213);
or U15092 (N_15092,N_10493,N_8197);
nor U15093 (N_15093,N_10224,N_11248);
nor U15094 (N_15094,N_8682,N_10027);
nand U15095 (N_15095,N_10146,N_8020);
xnor U15096 (N_15096,N_10846,N_9179);
nor U15097 (N_15097,N_11171,N_10001);
or U15098 (N_15098,N_9778,N_10664);
and U15099 (N_15099,N_9197,N_11512);
or U15100 (N_15100,N_8076,N_8810);
nand U15101 (N_15101,N_9860,N_10810);
xnor U15102 (N_15102,N_9121,N_9002);
xnor U15103 (N_15103,N_11850,N_11405);
xnor U15104 (N_15104,N_11106,N_11675);
nor U15105 (N_15105,N_10640,N_9094);
or U15106 (N_15106,N_9099,N_11021);
or U15107 (N_15107,N_10432,N_10930);
nor U15108 (N_15108,N_8094,N_10052);
nor U15109 (N_15109,N_10724,N_8839);
or U15110 (N_15110,N_8716,N_11248);
or U15111 (N_15111,N_9727,N_9825);
nor U15112 (N_15112,N_10452,N_10309);
xor U15113 (N_15113,N_11990,N_10750);
or U15114 (N_15114,N_10764,N_8458);
nor U15115 (N_15115,N_10541,N_9053);
nand U15116 (N_15116,N_10550,N_11399);
nand U15117 (N_15117,N_11313,N_10674);
or U15118 (N_15118,N_11072,N_8205);
nand U15119 (N_15119,N_11554,N_10908);
and U15120 (N_15120,N_9811,N_9819);
and U15121 (N_15121,N_11642,N_8575);
or U15122 (N_15122,N_11851,N_11695);
nor U15123 (N_15123,N_11279,N_8099);
and U15124 (N_15124,N_9319,N_9791);
nor U15125 (N_15125,N_8236,N_10352);
nand U15126 (N_15126,N_9072,N_10326);
nor U15127 (N_15127,N_10756,N_10063);
nand U15128 (N_15128,N_10340,N_10922);
xnor U15129 (N_15129,N_8775,N_10550);
nor U15130 (N_15130,N_9301,N_11515);
or U15131 (N_15131,N_9130,N_8728);
or U15132 (N_15132,N_10272,N_9579);
or U15133 (N_15133,N_10457,N_9745);
nand U15134 (N_15134,N_9705,N_10325);
nand U15135 (N_15135,N_10624,N_10589);
and U15136 (N_15136,N_11264,N_8009);
or U15137 (N_15137,N_8408,N_10873);
nand U15138 (N_15138,N_9652,N_11731);
xor U15139 (N_15139,N_8362,N_11432);
nand U15140 (N_15140,N_8688,N_9617);
nor U15141 (N_15141,N_8423,N_11000);
and U15142 (N_15142,N_10362,N_10699);
nor U15143 (N_15143,N_11601,N_10511);
xor U15144 (N_15144,N_10544,N_8490);
or U15145 (N_15145,N_9596,N_9873);
or U15146 (N_15146,N_9981,N_11774);
nand U15147 (N_15147,N_8503,N_10487);
and U15148 (N_15148,N_10152,N_8856);
xnor U15149 (N_15149,N_11346,N_10425);
nor U15150 (N_15150,N_9332,N_8696);
or U15151 (N_15151,N_8097,N_9720);
xnor U15152 (N_15152,N_8342,N_9506);
or U15153 (N_15153,N_9138,N_9472);
or U15154 (N_15154,N_8918,N_8224);
nand U15155 (N_15155,N_8877,N_9302);
or U15156 (N_15156,N_10994,N_10734);
nand U15157 (N_15157,N_11150,N_8857);
nor U15158 (N_15158,N_9337,N_11155);
nor U15159 (N_15159,N_9155,N_9893);
nor U15160 (N_15160,N_9097,N_11102);
nand U15161 (N_15161,N_8679,N_8013);
and U15162 (N_15162,N_10345,N_8639);
or U15163 (N_15163,N_10523,N_11508);
and U15164 (N_15164,N_9564,N_10293);
or U15165 (N_15165,N_10690,N_8473);
xnor U15166 (N_15166,N_8638,N_8317);
nand U15167 (N_15167,N_11892,N_10482);
nor U15168 (N_15168,N_11123,N_10927);
nand U15169 (N_15169,N_11845,N_8854);
nor U15170 (N_15170,N_8311,N_8476);
nand U15171 (N_15171,N_11049,N_8135);
xor U15172 (N_15172,N_11072,N_10401);
or U15173 (N_15173,N_10596,N_10778);
and U15174 (N_15174,N_8509,N_10694);
or U15175 (N_15175,N_8284,N_9844);
nor U15176 (N_15176,N_11243,N_11745);
nor U15177 (N_15177,N_9465,N_10749);
nor U15178 (N_15178,N_8932,N_9899);
nand U15179 (N_15179,N_11397,N_10022);
and U15180 (N_15180,N_10974,N_9871);
nand U15181 (N_15181,N_11395,N_8866);
and U15182 (N_15182,N_11371,N_8885);
nand U15183 (N_15183,N_11799,N_10127);
nand U15184 (N_15184,N_10088,N_8214);
or U15185 (N_15185,N_10370,N_9959);
or U15186 (N_15186,N_8709,N_11661);
and U15187 (N_15187,N_9539,N_8988);
nand U15188 (N_15188,N_9768,N_8391);
nand U15189 (N_15189,N_9966,N_10963);
or U15190 (N_15190,N_11256,N_8025);
or U15191 (N_15191,N_8264,N_8112);
and U15192 (N_15192,N_9078,N_8264);
and U15193 (N_15193,N_11579,N_11321);
and U15194 (N_15194,N_8320,N_8888);
nor U15195 (N_15195,N_11824,N_10149);
nor U15196 (N_15196,N_11911,N_10476);
xor U15197 (N_15197,N_11646,N_9914);
nand U15198 (N_15198,N_9589,N_11080);
or U15199 (N_15199,N_11011,N_11291);
and U15200 (N_15200,N_11466,N_8615);
nand U15201 (N_15201,N_9331,N_11925);
nor U15202 (N_15202,N_9342,N_11734);
nand U15203 (N_15203,N_11869,N_8312);
nand U15204 (N_15204,N_8388,N_11163);
and U15205 (N_15205,N_9237,N_11183);
nand U15206 (N_15206,N_9338,N_10888);
nor U15207 (N_15207,N_9185,N_9825);
xor U15208 (N_15208,N_11050,N_10203);
and U15209 (N_15209,N_8943,N_10242);
or U15210 (N_15210,N_9892,N_10595);
nor U15211 (N_15211,N_8161,N_11565);
nand U15212 (N_15212,N_9757,N_10927);
and U15213 (N_15213,N_8686,N_11763);
nand U15214 (N_15214,N_10644,N_9133);
nor U15215 (N_15215,N_11279,N_8675);
or U15216 (N_15216,N_9976,N_9338);
nand U15217 (N_15217,N_8928,N_10667);
or U15218 (N_15218,N_9593,N_10977);
nand U15219 (N_15219,N_11907,N_10986);
nand U15220 (N_15220,N_11312,N_11041);
or U15221 (N_15221,N_9952,N_8689);
and U15222 (N_15222,N_11773,N_9315);
and U15223 (N_15223,N_9661,N_11708);
nand U15224 (N_15224,N_9844,N_11726);
nand U15225 (N_15225,N_11643,N_11178);
and U15226 (N_15226,N_8056,N_8740);
or U15227 (N_15227,N_9806,N_8513);
xor U15228 (N_15228,N_11245,N_8467);
nor U15229 (N_15229,N_9651,N_10824);
or U15230 (N_15230,N_11746,N_10106);
nand U15231 (N_15231,N_10940,N_8635);
xnor U15232 (N_15232,N_11268,N_10949);
xnor U15233 (N_15233,N_10211,N_10724);
or U15234 (N_15234,N_9812,N_9650);
nand U15235 (N_15235,N_8921,N_11963);
xor U15236 (N_15236,N_11985,N_9512);
or U15237 (N_15237,N_9787,N_9341);
and U15238 (N_15238,N_9693,N_8397);
nand U15239 (N_15239,N_9080,N_9316);
and U15240 (N_15240,N_8246,N_10520);
nand U15241 (N_15241,N_10578,N_9056);
nand U15242 (N_15242,N_9240,N_9631);
nor U15243 (N_15243,N_8585,N_8594);
nor U15244 (N_15244,N_11048,N_8114);
nor U15245 (N_15245,N_10215,N_10733);
nor U15246 (N_15246,N_10098,N_9228);
xnor U15247 (N_15247,N_11921,N_9293);
or U15248 (N_15248,N_8689,N_11378);
nor U15249 (N_15249,N_9142,N_9776);
or U15250 (N_15250,N_10077,N_10187);
nor U15251 (N_15251,N_11047,N_11241);
nor U15252 (N_15252,N_10736,N_10157);
and U15253 (N_15253,N_8474,N_10548);
or U15254 (N_15254,N_10640,N_8553);
nor U15255 (N_15255,N_10347,N_8952);
or U15256 (N_15256,N_9836,N_11766);
or U15257 (N_15257,N_11940,N_8266);
or U15258 (N_15258,N_11858,N_9066);
nor U15259 (N_15259,N_8990,N_11280);
nand U15260 (N_15260,N_9883,N_11660);
xnor U15261 (N_15261,N_8615,N_10882);
or U15262 (N_15262,N_11467,N_8360);
nand U15263 (N_15263,N_8086,N_11006);
or U15264 (N_15264,N_8425,N_8150);
and U15265 (N_15265,N_8354,N_10908);
nor U15266 (N_15266,N_11720,N_11357);
or U15267 (N_15267,N_8414,N_9940);
or U15268 (N_15268,N_9733,N_10341);
nor U15269 (N_15269,N_11106,N_10584);
nor U15270 (N_15270,N_8483,N_8036);
nand U15271 (N_15271,N_10287,N_9787);
and U15272 (N_15272,N_8977,N_11408);
or U15273 (N_15273,N_8591,N_10216);
nand U15274 (N_15274,N_11338,N_8297);
nand U15275 (N_15275,N_8298,N_10203);
xnor U15276 (N_15276,N_8823,N_9659);
or U15277 (N_15277,N_9237,N_9762);
nand U15278 (N_15278,N_11443,N_9523);
and U15279 (N_15279,N_10032,N_9161);
nand U15280 (N_15280,N_9224,N_10168);
nor U15281 (N_15281,N_11470,N_10267);
nand U15282 (N_15282,N_10148,N_9769);
nand U15283 (N_15283,N_11931,N_11734);
and U15284 (N_15284,N_9058,N_8158);
or U15285 (N_15285,N_10321,N_9548);
and U15286 (N_15286,N_10403,N_11618);
and U15287 (N_15287,N_8706,N_11148);
and U15288 (N_15288,N_11348,N_10332);
nand U15289 (N_15289,N_10627,N_8684);
and U15290 (N_15290,N_9546,N_11340);
nor U15291 (N_15291,N_9384,N_8636);
and U15292 (N_15292,N_10570,N_11615);
nor U15293 (N_15293,N_9158,N_10295);
nand U15294 (N_15294,N_11973,N_11646);
and U15295 (N_15295,N_11117,N_11804);
nand U15296 (N_15296,N_11766,N_10257);
nor U15297 (N_15297,N_8934,N_11810);
and U15298 (N_15298,N_9387,N_8082);
nor U15299 (N_15299,N_11721,N_9689);
nor U15300 (N_15300,N_10869,N_10410);
or U15301 (N_15301,N_9167,N_11285);
nand U15302 (N_15302,N_9460,N_11977);
xor U15303 (N_15303,N_8721,N_9513);
and U15304 (N_15304,N_11491,N_9036);
nand U15305 (N_15305,N_9124,N_9325);
or U15306 (N_15306,N_8898,N_9085);
nor U15307 (N_15307,N_9872,N_10360);
nor U15308 (N_15308,N_11930,N_8465);
nor U15309 (N_15309,N_11764,N_11582);
and U15310 (N_15310,N_8271,N_10841);
and U15311 (N_15311,N_8834,N_9095);
xor U15312 (N_15312,N_11344,N_11991);
nor U15313 (N_15313,N_11495,N_9122);
nor U15314 (N_15314,N_9717,N_11161);
and U15315 (N_15315,N_10573,N_9547);
and U15316 (N_15316,N_11695,N_9588);
and U15317 (N_15317,N_8584,N_8669);
nand U15318 (N_15318,N_8628,N_8144);
and U15319 (N_15319,N_11785,N_10784);
nor U15320 (N_15320,N_11773,N_8237);
and U15321 (N_15321,N_9811,N_10394);
nand U15322 (N_15322,N_8579,N_9743);
nand U15323 (N_15323,N_9014,N_10410);
nand U15324 (N_15324,N_11156,N_10829);
nand U15325 (N_15325,N_8247,N_9127);
nor U15326 (N_15326,N_8710,N_10330);
and U15327 (N_15327,N_10814,N_10501);
or U15328 (N_15328,N_11113,N_9957);
and U15329 (N_15329,N_8471,N_9395);
nand U15330 (N_15330,N_9696,N_8787);
nor U15331 (N_15331,N_11753,N_9683);
and U15332 (N_15332,N_10416,N_9847);
nand U15333 (N_15333,N_9452,N_9139);
nand U15334 (N_15334,N_11504,N_11920);
and U15335 (N_15335,N_11275,N_8256);
nand U15336 (N_15336,N_8472,N_8689);
nand U15337 (N_15337,N_11223,N_9368);
nand U15338 (N_15338,N_10667,N_10765);
nand U15339 (N_15339,N_8331,N_10070);
nand U15340 (N_15340,N_10107,N_8771);
and U15341 (N_15341,N_8882,N_9906);
or U15342 (N_15342,N_9318,N_8676);
xnor U15343 (N_15343,N_11007,N_11219);
nand U15344 (N_15344,N_9670,N_10316);
or U15345 (N_15345,N_8449,N_11376);
or U15346 (N_15346,N_9080,N_8736);
nand U15347 (N_15347,N_10111,N_9664);
nand U15348 (N_15348,N_11610,N_11908);
nand U15349 (N_15349,N_8586,N_8506);
nor U15350 (N_15350,N_8344,N_11861);
nor U15351 (N_15351,N_9978,N_9849);
xor U15352 (N_15352,N_8076,N_8105);
nand U15353 (N_15353,N_10168,N_8699);
xnor U15354 (N_15354,N_8767,N_10696);
or U15355 (N_15355,N_11743,N_11278);
nand U15356 (N_15356,N_10839,N_8316);
nor U15357 (N_15357,N_10035,N_11348);
or U15358 (N_15358,N_11375,N_11306);
nand U15359 (N_15359,N_8307,N_8245);
nand U15360 (N_15360,N_8228,N_11488);
nand U15361 (N_15361,N_9011,N_10571);
nand U15362 (N_15362,N_11324,N_11385);
and U15363 (N_15363,N_10724,N_10087);
and U15364 (N_15364,N_11024,N_9209);
and U15365 (N_15365,N_11228,N_10742);
nor U15366 (N_15366,N_10190,N_10117);
and U15367 (N_15367,N_8710,N_8966);
xor U15368 (N_15368,N_10085,N_11932);
nor U15369 (N_15369,N_11207,N_8640);
and U15370 (N_15370,N_11664,N_8025);
nor U15371 (N_15371,N_11088,N_11671);
nor U15372 (N_15372,N_8806,N_11433);
and U15373 (N_15373,N_10091,N_10912);
and U15374 (N_15374,N_11319,N_11181);
nor U15375 (N_15375,N_10340,N_8218);
nand U15376 (N_15376,N_8085,N_8571);
or U15377 (N_15377,N_10867,N_11347);
and U15378 (N_15378,N_11381,N_11342);
nor U15379 (N_15379,N_9726,N_9275);
nor U15380 (N_15380,N_8989,N_10140);
nor U15381 (N_15381,N_8864,N_11220);
or U15382 (N_15382,N_10834,N_9962);
or U15383 (N_15383,N_10314,N_8547);
and U15384 (N_15384,N_10830,N_8199);
and U15385 (N_15385,N_11110,N_8177);
nand U15386 (N_15386,N_8426,N_11930);
nor U15387 (N_15387,N_9514,N_9440);
xnor U15388 (N_15388,N_8168,N_9697);
and U15389 (N_15389,N_11071,N_8172);
nand U15390 (N_15390,N_10224,N_10140);
nand U15391 (N_15391,N_11679,N_11049);
nor U15392 (N_15392,N_9300,N_9373);
nand U15393 (N_15393,N_8724,N_9750);
or U15394 (N_15394,N_11032,N_11829);
and U15395 (N_15395,N_11229,N_9201);
or U15396 (N_15396,N_9781,N_8879);
or U15397 (N_15397,N_11586,N_8383);
nor U15398 (N_15398,N_11642,N_10089);
and U15399 (N_15399,N_9069,N_9891);
or U15400 (N_15400,N_9144,N_8519);
and U15401 (N_15401,N_10257,N_10527);
or U15402 (N_15402,N_10793,N_8245);
nand U15403 (N_15403,N_10460,N_11798);
and U15404 (N_15404,N_9864,N_9807);
or U15405 (N_15405,N_8538,N_11518);
and U15406 (N_15406,N_9960,N_8797);
and U15407 (N_15407,N_8589,N_8273);
xor U15408 (N_15408,N_11490,N_10988);
xor U15409 (N_15409,N_10518,N_9975);
nand U15410 (N_15410,N_11181,N_11538);
nand U15411 (N_15411,N_9505,N_10830);
xnor U15412 (N_15412,N_10125,N_9578);
or U15413 (N_15413,N_8876,N_9556);
nor U15414 (N_15414,N_10101,N_8569);
nor U15415 (N_15415,N_9584,N_11006);
nor U15416 (N_15416,N_8026,N_8305);
nand U15417 (N_15417,N_9470,N_9523);
or U15418 (N_15418,N_11753,N_11706);
or U15419 (N_15419,N_10922,N_11397);
xor U15420 (N_15420,N_11845,N_10029);
nor U15421 (N_15421,N_8078,N_11761);
and U15422 (N_15422,N_9659,N_9352);
and U15423 (N_15423,N_9964,N_9996);
nor U15424 (N_15424,N_11812,N_10516);
nor U15425 (N_15425,N_10394,N_8327);
nand U15426 (N_15426,N_11237,N_8155);
xor U15427 (N_15427,N_8222,N_8231);
nor U15428 (N_15428,N_11329,N_8643);
nand U15429 (N_15429,N_10148,N_9416);
nor U15430 (N_15430,N_11267,N_10799);
xnor U15431 (N_15431,N_8823,N_11589);
nand U15432 (N_15432,N_9070,N_8743);
nand U15433 (N_15433,N_10092,N_9230);
and U15434 (N_15434,N_8490,N_11112);
xor U15435 (N_15435,N_9912,N_10342);
and U15436 (N_15436,N_9178,N_9730);
nand U15437 (N_15437,N_9941,N_9232);
and U15438 (N_15438,N_9025,N_8120);
xor U15439 (N_15439,N_8170,N_9858);
and U15440 (N_15440,N_11555,N_10813);
and U15441 (N_15441,N_10460,N_10404);
nor U15442 (N_15442,N_9377,N_11528);
and U15443 (N_15443,N_11812,N_9878);
or U15444 (N_15444,N_11336,N_8651);
xor U15445 (N_15445,N_11125,N_11781);
nand U15446 (N_15446,N_10751,N_11547);
or U15447 (N_15447,N_10439,N_8881);
nor U15448 (N_15448,N_11509,N_11589);
xnor U15449 (N_15449,N_11033,N_10450);
and U15450 (N_15450,N_9474,N_11094);
nor U15451 (N_15451,N_9601,N_9494);
or U15452 (N_15452,N_11273,N_11449);
or U15453 (N_15453,N_8710,N_10124);
nand U15454 (N_15454,N_11993,N_11565);
and U15455 (N_15455,N_11006,N_9605);
or U15456 (N_15456,N_10801,N_10580);
nor U15457 (N_15457,N_11384,N_11845);
or U15458 (N_15458,N_8341,N_9105);
nor U15459 (N_15459,N_11826,N_10074);
xor U15460 (N_15460,N_11551,N_9246);
and U15461 (N_15461,N_9600,N_9990);
nor U15462 (N_15462,N_8710,N_8767);
xor U15463 (N_15463,N_10484,N_11233);
and U15464 (N_15464,N_8907,N_9699);
nor U15465 (N_15465,N_9432,N_10090);
and U15466 (N_15466,N_8971,N_10637);
nand U15467 (N_15467,N_8855,N_10468);
nor U15468 (N_15468,N_11522,N_11855);
or U15469 (N_15469,N_9448,N_9493);
and U15470 (N_15470,N_10007,N_11254);
nor U15471 (N_15471,N_10113,N_11196);
nand U15472 (N_15472,N_10757,N_10575);
and U15473 (N_15473,N_10605,N_11302);
nand U15474 (N_15474,N_8617,N_10253);
or U15475 (N_15475,N_9181,N_10284);
or U15476 (N_15476,N_11062,N_8663);
xor U15477 (N_15477,N_10687,N_10245);
nor U15478 (N_15478,N_8578,N_8493);
xor U15479 (N_15479,N_9824,N_8800);
and U15480 (N_15480,N_11857,N_10226);
nand U15481 (N_15481,N_9820,N_8731);
xor U15482 (N_15482,N_11283,N_10195);
nand U15483 (N_15483,N_9433,N_10546);
nand U15484 (N_15484,N_9347,N_11788);
or U15485 (N_15485,N_9946,N_9013);
xnor U15486 (N_15486,N_8704,N_8961);
nor U15487 (N_15487,N_8492,N_11321);
or U15488 (N_15488,N_10440,N_11837);
xor U15489 (N_15489,N_11007,N_8992);
nand U15490 (N_15490,N_11800,N_9320);
or U15491 (N_15491,N_8388,N_9909);
or U15492 (N_15492,N_9123,N_9275);
nand U15493 (N_15493,N_11736,N_11880);
nand U15494 (N_15494,N_10667,N_11765);
nor U15495 (N_15495,N_11880,N_9498);
xor U15496 (N_15496,N_9393,N_8822);
and U15497 (N_15497,N_11084,N_8068);
xor U15498 (N_15498,N_10234,N_11649);
and U15499 (N_15499,N_8579,N_8631);
and U15500 (N_15500,N_9329,N_8735);
or U15501 (N_15501,N_10039,N_8914);
xor U15502 (N_15502,N_11875,N_8699);
or U15503 (N_15503,N_9252,N_9276);
and U15504 (N_15504,N_10873,N_11549);
nand U15505 (N_15505,N_8135,N_8200);
and U15506 (N_15506,N_11520,N_10907);
and U15507 (N_15507,N_8534,N_10893);
nor U15508 (N_15508,N_11486,N_9585);
and U15509 (N_15509,N_9389,N_8509);
nor U15510 (N_15510,N_9625,N_10321);
and U15511 (N_15511,N_8060,N_9598);
xor U15512 (N_15512,N_9571,N_10532);
and U15513 (N_15513,N_8757,N_8424);
and U15514 (N_15514,N_9501,N_8665);
or U15515 (N_15515,N_8312,N_8750);
nor U15516 (N_15516,N_8073,N_10676);
nor U15517 (N_15517,N_11743,N_9691);
nor U15518 (N_15518,N_9797,N_9185);
or U15519 (N_15519,N_10778,N_10236);
nor U15520 (N_15520,N_9859,N_11491);
nor U15521 (N_15521,N_8155,N_11143);
nor U15522 (N_15522,N_9584,N_9875);
or U15523 (N_15523,N_11406,N_8244);
and U15524 (N_15524,N_8808,N_9403);
nor U15525 (N_15525,N_11054,N_8762);
or U15526 (N_15526,N_9560,N_8623);
and U15527 (N_15527,N_9572,N_11534);
nand U15528 (N_15528,N_11923,N_8922);
or U15529 (N_15529,N_8417,N_11932);
xor U15530 (N_15530,N_9790,N_10057);
nand U15531 (N_15531,N_10526,N_8018);
or U15532 (N_15532,N_8385,N_8729);
or U15533 (N_15533,N_10396,N_10708);
nand U15534 (N_15534,N_11289,N_11898);
and U15535 (N_15535,N_8926,N_11466);
or U15536 (N_15536,N_8511,N_9277);
nor U15537 (N_15537,N_8960,N_9901);
nor U15538 (N_15538,N_11278,N_10348);
nand U15539 (N_15539,N_8612,N_8661);
nor U15540 (N_15540,N_8800,N_10690);
nand U15541 (N_15541,N_11998,N_8346);
nor U15542 (N_15542,N_8870,N_11641);
nand U15543 (N_15543,N_11130,N_10240);
nor U15544 (N_15544,N_8982,N_8692);
nand U15545 (N_15545,N_11800,N_8033);
and U15546 (N_15546,N_10294,N_11477);
nor U15547 (N_15547,N_11245,N_8850);
xnor U15548 (N_15548,N_8709,N_9790);
and U15549 (N_15549,N_8851,N_10675);
nor U15550 (N_15550,N_10982,N_9635);
xnor U15551 (N_15551,N_9150,N_10676);
nand U15552 (N_15552,N_11434,N_11461);
and U15553 (N_15553,N_11657,N_10610);
and U15554 (N_15554,N_10357,N_11572);
xor U15555 (N_15555,N_10887,N_8073);
nor U15556 (N_15556,N_11226,N_11830);
or U15557 (N_15557,N_8834,N_10998);
and U15558 (N_15558,N_11086,N_10842);
nand U15559 (N_15559,N_10913,N_8282);
xnor U15560 (N_15560,N_10470,N_8855);
and U15561 (N_15561,N_10029,N_11230);
nand U15562 (N_15562,N_11910,N_8411);
or U15563 (N_15563,N_10630,N_10569);
nor U15564 (N_15564,N_11199,N_10996);
and U15565 (N_15565,N_8888,N_11682);
or U15566 (N_15566,N_9062,N_9977);
and U15567 (N_15567,N_11843,N_10199);
or U15568 (N_15568,N_8199,N_10166);
or U15569 (N_15569,N_8936,N_8379);
nand U15570 (N_15570,N_10225,N_11438);
and U15571 (N_15571,N_9132,N_10293);
nor U15572 (N_15572,N_11742,N_11319);
or U15573 (N_15573,N_11211,N_11593);
nor U15574 (N_15574,N_10594,N_8641);
and U15575 (N_15575,N_10820,N_9371);
nor U15576 (N_15576,N_8090,N_10889);
or U15577 (N_15577,N_8148,N_11527);
nand U15578 (N_15578,N_11076,N_10808);
or U15579 (N_15579,N_10349,N_10828);
or U15580 (N_15580,N_9341,N_11570);
nor U15581 (N_15581,N_11025,N_10597);
nand U15582 (N_15582,N_11065,N_10901);
nand U15583 (N_15583,N_10067,N_11218);
nand U15584 (N_15584,N_11721,N_11407);
nor U15585 (N_15585,N_11734,N_11148);
nor U15586 (N_15586,N_11450,N_8492);
nor U15587 (N_15587,N_8094,N_11915);
and U15588 (N_15588,N_8369,N_10162);
nor U15589 (N_15589,N_11629,N_8888);
nand U15590 (N_15590,N_10491,N_10563);
or U15591 (N_15591,N_9677,N_11810);
or U15592 (N_15592,N_10919,N_8266);
and U15593 (N_15593,N_9110,N_11314);
nand U15594 (N_15594,N_11462,N_11176);
nand U15595 (N_15595,N_8386,N_11233);
and U15596 (N_15596,N_11057,N_9034);
nor U15597 (N_15597,N_11092,N_8307);
or U15598 (N_15598,N_8361,N_10192);
xor U15599 (N_15599,N_10941,N_11377);
nor U15600 (N_15600,N_8571,N_11853);
nand U15601 (N_15601,N_10142,N_10081);
and U15602 (N_15602,N_8016,N_11647);
or U15603 (N_15603,N_8647,N_8490);
nor U15604 (N_15604,N_8462,N_11980);
or U15605 (N_15605,N_10485,N_11163);
nand U15606 (N_15606,N_11574,N_10132);
and U15607 (N_15607,N_9163,N_9858);
nand U15608 (N_15608,N_8347,N_11615);
and U15609 (N_15609,N_10638,N_9177);
and U15610 (N_15610,N_9499,N_8385);
and U15611 (N_15611,N_8180,N_9823);
nor U15612 (N_15612,N_9847,N_11744);
nand U15613 (N_15613,N_9962,N_9358);
nor U15614 (N_15614,N_10152,N_9977);
or U15615 (N_15615,N_11242,N_8434);
xnor U15616 (N_15616,N_10942,N_10196);
nor U15617 (N_15617,N_11788,N_10101);
nand U15618 (N_15618,N_11750,N_10515);
and U15619 (N_15619,N_8933,N_8616);
nor U15620 (N_15620,N_10158,N_11631);
or U15621 (N_15621,N_11681,N_10141);
nand U15622 (N_15622,N_9435,N_11612);
nor U15623 (N_15623,N_10131,N_8930);
xnor U15624 (N_15624,N_10021,N_9261);
xnor U15625 (N_15625,N_11774,N_8140);
xnor U15626 (N_15626,N_11699,N_11972);
nor U15627 (N_15627,N_9437,N_10240);
nand U15628 (N_15628,N_10248,N_10525);
nor U15629 (N_15629,N_9420,N_10096);
nand U15630 (N_15630,N_10051,N_11391);
and U15631 (N_15631,N_11529,N_11029);
nor U15632 (N_15632,N_11068,N_10338);
nor U15633 (N_15633,N_11289,N_11175);
nor U15634 (N_15634,N_9860,N_10638);
or U15635 (N_15635,N_10965,N_11712);
or U15636 (N_15636,N_8131,N_9409);
and U15637 (N_15637,N_8975,N_8029);
and U15638 (N_15638,N_11077,N_8776);
and U15639 (N_15639,N_9389,N_9824);
or U15640 (N_15640,N_9962,N_10293);
xor U15641 (N_15641,N_8407,N_10738);
or U15642 (N_15642,N_8709,N_9173);
or U15643 (N_15643,N_9536,N_8215);
or U15644 (N_15644,N_8623,N_10328);
xnor U15645 (N_15645,N_11614,N_8870);
or U15646 (N_15646,N_9209,N_10423);
or U15647 (N_15647,N_11288,N_11444);
and U15648 (N_15648,N_9203,N_11109);
nand U15649 (N_15649,N_11782,N_8097);
or U15650 (N_15650,N_11249,N_9557);
nand U15651 (N_15651,N_9546,N_10044);
nand U15652 (N_15652,N_9267,N_9753);
nor U15653 (N_15653,N_11937,N_8742);
or U15654 (N_15654,N_11639,N_9353);
and U15655 (N_15655,N_8828,N_10027);
nand U15656 (N_15656,N_8684,N_8731);
nor U15657 (N_15657,N_10165,N_8378);
or U15658 (N_15658,N_9606,N_11424);
nor U15659 (N_15659,N_11601,N_8713);
nand U15660 (N_15660,N_10381,N_10179);
or U15661 (N_15661,N_9232,N_8834);
or U15662 (N_15662,N_11143,N_11790);
and U15663 (N_15663,N_9272,N_9000);
and U15664 (N_15664,N_10456,N_9679);
xnor U15665 (N_15665,N_8671,N_9711);
xnor U15666 (N_15666,N_9480,N_8637);
nor U15667 (N_15667,N_9137,N_8963);
and U15668 (N_15668,N_11187,N_11431);
and U15669 (N_15669,N_9975,N_10647);
and U15670 (N_15670,N_10801,N_10722);
nor U15671 (N_15671,N_10608,N_10598);
or U15672 (N_15672,N_8565,N_10443);
nor U15673 (N_15673,N_11116,N_8826);
or U15674 (N_15674,N_10966,N_11959);
nor U15675 (N_15675,N_11776,N_10366);
xor U15676 (N_15676,N_8628,N_10702);
nor U15677 (N_15677,N_9415,N_8134);
or U15678 (N_15678,N_8017,N_8779);
nand U15679 (N_15679,N_10126,N_8171);
nor U15680 (N_15680,N_9917,N_9375);
xor U15681 (N_15681,N_10322,N_9303);
and U15682 (N_15682,N_9358,N_11119);
and U15683 (N_15683,N_9572,N_10169);
nor U15684 (N_15684,N_8834,N_11661);
or U15685 (N_15685,N_8768,N_8352);
nor U15686 (N_15686,N_11461,N_8170);
nor U15687 (N_15687,N_11967,N_9828);
nand U15688 (N_15688,N_11348,N_8531);
nand U15689 (N_15689,N_11086,N_10227);
or U15690 (N_15690,N_10857,N_10162);
or U15691 (N_15691,N_8867,N_9546);
nor U15692 (N_15692,N_10509,N_8374);
xnor U15693 (N_15693,N_11555,N_9616);
or U15694 (N_15694,N_8945,N_8302);
nand U15695 (N_15695,N_8268,N_9059);
nand U15696 (N_15696,N_11707,N_9126);
nor U15697 (N_15697,N_8773,N_10042);
nand U15698 (N_15698,N_9795,N_11170);
or U15699 (N_15699,N_11442,N_10238);
nand U15700 (N_15700,N_9650,N_8681);
xor U15701 (N_15701,N_11818,N_11744);
and U15702 (N_15702,N_9519,N_11662);
nor U15703 (N_15703,N_11010,N_9814);
or U15704 (N_15704,N_8142,N_9680);
or U15705 (N_15705,N_9106,N_8476);
and U15706 (N_15706,N_8097,N_8510);
or U15707 (N_15707,N_11865,N_10505);
or U15708 (N_15708,N_8473,N_8604);
and U15709 (N_15709,N_8948,N_8093);
and U15710 (N_15710,N_8099,N_11298);
nor U15711 (N_15711,N_11420,N_8509);
nand U15712 (N_15712,N_11379,N_10339);
and U15713 (N_15713,N_9603,N_11161);
or U15714 (N_15714,N_8125,N_10525);
and U15715 (N_15715,N_9311,N_10546);
nor U15716 (N_15716,N_9209,N_10389);
and U15717 (N_15717,N_8088,N_10071);
xor U15718 (N_15718,N_10931,N_9421);
nor U15719 (N_15719,N_9731,N_9465);
and U15720 (N_15720,N_9382,N_11462);
or U15721 (N_15721,N_10446,N_10665);
and U15722 (N_15722,N_8162,N_10802);
and U15723 (N_15723,N_9855,N_8427);
nor U15724 (N_15724,N_10584,N_11802);
nor U15725 (N_15725,N_10060,N_11568);
nand U15726 (N_15726,N_11997,N_10059);
xor U15727 (N_15727,N_10066,N_11974);
nor U15728 (N_15728,N_9640,N_8765);
nand U15729 (N_15729,N_11572,N_8766);
or U15730 (N_15730,N_11875,N_11122);
nor U15731 (N_15731,N_10634,N_9539);
and U15732 (N_15732,N_9145,N_10978);
xnor U15733 (N_15733,N_11571,N_9813);
nand U15734 (N_15734,N_8878,N_9561);
nand U15735 (N_15735,N_9407,N_9003);
nor U15736 (N_15736,N_11912,N_11600);
nor U15737 (N_15737,N_9298,N_9538);
nor U15738 (N_15738,N_8911,N_10170);
and U15739 (N_15739,N_9104,N_8434);
xnor U15740 (N_15740,N_9621,N_11920);
nand U15741 (N_15741,N_10081,N_11172);
and U15742 (N_15742,N_9486,N_9476);
or U15743 (N_15743,N_11334,N_11017);
xnor U15744 (N_15744,N_9881,N_10832);
nor U15745 (N_15745,N_8978,N_9034);
nand U15746 (N_15746,N_9307,N_8518);
or U15747 (N_15747,N_10341,N_8770);
and U15748 (N_15748,N_10163,N_9296);
and U15749 (N_15749,N_8120,N_8275);
nand U15750 (N_15750,N_8366,N_10995);
or U15751 (N_15751,N_10506,N_11093);
xnor U15752 (N_15752,N_10173,N_8429);
and U15753 (N_15753,N_9654,N_9277);
or U15754 (N_15754,N_11680,N_11896);
nor U15755 (N_15755,N_10759,N_10551);
nand U15756 (N_15756,N_9334,N_11124);
nor U15757 (N_15757,N_10011,N_10530);
or U15758 (N_15758,N_10448,N_8615);
nor U15759 (N_15759,N_11339,N_11545);
nor U15760 (N_15760,N_9776,N_10503);
nor U15761 (N_15761,N_9626,N_9889);
nand U15762 (N_15762,N_9404,N_9169);
nand U15763 (N_15763,N_9897,N_10663);
xnor U15764 (N_15764,N_9523,N_10320);
nor U15765 (N_15765,N_11280,N_8215);
and U15766 (N_15766,N_9894,N_9197);
or U15767 (N_15767,N_10860,N_11430);
nand U15768 (N_15768,N_10846,N_10870);
and U15769 (N_15769,N_8964,N_10278);
nand U15770 (N_15770,N_8793,N_10265);
nor U15771 (N_15771,N_9428,N_8849);
nand U15772 (N_15772,N_9826,N_11327);
nor U15773 (N_15773,N_10868,N_10839);
and U15774 (N_15774,N_10927,N_8983);
and U15775 (N_15775,N_11602,N_11566);
nand U15776 (N_15776,N_8470,N_10156);
nor U15777 (N_15777,N_11281,N_8914);
nand U15778 (N_15778,N_10376,N_10488);
nand U15779 (N_15779,N_11012,N_9290);
xor U15780 (N_15780,N_10766,N_8360);
or U15781 (N_15781,N_8521,N_9573);
nor U15782 (N_15782,N_11568,N_9256);
or U15783 (N_15783,N_11936,N_11324);
or U15784 (N_15784,N_9144,N_10779);
and U15785 (N_15785,N_8759,N_11431);
nand U15786 (N_15786,N_11600,N_8559);
and U15787 (N_15787,N_9714,N_11852);
nor U15788 (N_15788,N_9129,N_10627);
or U15789 (N_15789,N_11673,N_10705);
nand U15790 (N_15790,N_9039,N_10680);
nand U15791 (N_15791,N_8088,N_10015);
nand U15792 (N_15792,N_8689,N_9398);
xor U15793 (N_15793,N_10339,N_8424);
nand U15794 (N_15794,N_9877,N_10814);
and U15795 (N_15795,N_9697,N_8152);
nand U15796 (N_15796,N_9147,N_9823);
nand U15797 (N_15797,N_9585,N_11535);
nand U15798 (N_15798,N_11057,N_8881);
nand U15799 (N_15799,N_9169,N_11333);
or U15800 (N_15800,N_11038,N_9140);
nand U15801 (N_15801,N_9367,N_10897);
and U15802 (N_15802,N_11886,N_9695);
nor U15803 (N_15803,N_9479,N_10829);
nand U15804 (N_15804,N_10328,N_9183);
or U15805 (N_15805,N_11508,N_8946);
or U15806 (N_15806,N_9526,N_11393);
nor U15807 (N_15807,N_10104,N_8496);
nor U15808 (N_15808,N_11646,N_9753);
xnor U15809 (N_15809,N_8701,N_8206);
nand U15810 (N_15810,N_11388,N_10807);
nor U15811 (N_15811,N_8893,N_10167);
and U15812 (N_15812,N_11439,N_8319);
nand U15813 (N_15813,N_8139,N_8142);
nor U15814 (N_15814,N_11666,N_9966);
and U15815 (N_15815,N_9570,N_11719);
nor U15816 (N_15816,N_11891,N_10949);
nor U15817 (N_15817,N_8145,N_8661);
nor U15818 (N_15818,N_8881,N_11751);
nor U15819 (N_15819,N_10166,N_9657);
or U15820 (N_15820,N_11948,N_11616);
nor U15821 (N_15821,N_9857,N_11732);
xnor U15822 (N_15822,N_8999,N_9788);
and U15823 (N_15823,N_8937,N_9739);
xnor U15824 (N_15824,N_8420,N_8392);
or U15825 (N_15825,N_10249,N_8957);
xnor U15826 (N_15826,N_8698,N_8689);
and U15827 (N_15827,N_10116,N_9162);
xor U15828 (N_15828,N_9787,N_8104);
or U15829 (N_15829,N_9996,N_11520);
nor U15830 (N_15830,N_8891,N_11882);
and U15831 (N_15831,N_9955,N_9660);
nor U15832 (N_15832,N_9783,N_9977);
nand U15833 (N_15833,N_11650,N_8430);
and U15834 (N_15834,N_10952,N_11373);
nor U15835 (N_15835,N_8753,N_9077);
and U15836 (N_15836,N_10161,N_9292);
and U15837 (N_15837,N_9372,N_11943);
nand U15838 (N_15838,N_11958,N_9822);
and U15839 (N_15839,N_9087,N_8129);
and U15840 (N_15840,N_11547,N_9614);
nor U15841 (N_15841,N_11608,N_11160);
nor U15842 (N_15842,N_10175,N_9678);
or U15843 (N_15843,N_8696,N_9625);
or U15844 (N_15844,N_9983,N_9628);
nand U15845 (N_15845,N_11479,N_8935);
or U15846 (N_15846,N_8710,N_8844);
and U15847 (N_15847,N_9191,N_8075);
xor U15848 (N_15848,N_10503,N_10221);
or U15849 (N_15849,N_10850,N_11919);
nand U15850 (N_15850,N_9149,N_9336);
or U15851 (N_15851,N_9915,N_11595);
or U15852 (N_15852,N_8573,N_8234);
and U15853 (N_15853,N_8665,N_8292);
nor U15854 (N_15854,N_8656,N_8235);
nor U15855 (N_15855,N_11860,N_11471);
nand U15856 (N_15856,N_9610,N_11925);
nor U15857 (N_15857,N_11115,N_11277);
or U15858 (N_15858,N_9612,N_10386);
and U15859 (N_15859,N_8547,N_11593);
or U15860 (N_15860,N_8178,N_11741);
and U15861 (N_15861,N_11201,N_10301);
nor U15862 (N_15862,N_8785,N_9193);
or U15863 (N_15863,N_10468,N_8834);
or U15864 (N_15864,N_11127,N_11843);
nor U15865 (N_15865,N_11573,N_11719);
nand U15866 (N_15866,N_11268,N_10847);
nor U15867 (N_15867,N_9663,N_10924);
and U15868 (N_15868,N_8764,N_9875);
and U15869 (N_15869,N_10899,N_8942);
and U15870 (N_15870,N_8053,N_8253);
or U15871 (N_15871,N_11855,N_11450);
and U15872 (N_15872,N_8593,N_11954);
and U15873 (N_15873,N_11975,N_9028);
xnor U15874 (N_15874,N_11554,N_10287);
or U15875 (N_15875,N_11220,N_10535);
or U15876 (N_15876,N_11544,N_8004);
nor U15877 (N_15877,N_9341,N_9725);
or U15878 (N_15878,N_8329,N_10037);
nand U15879 (N_15879,N_9501,N_11951);
and U15880 (N_15880,N_8397,N_8540);
xor U15881 (N_15881,N_11626,N_11832);
nand U15882 (N_15882,N_9943,N_8474);
or U15883 (N_15883,N_9115,N_11552);
nor U15884 (N_15884,N_9146,N_10310);
or U15885 (N_15885,N_10076,N_11814);
or U15886 (N_15886,N_9989,N_8275);
or U15887 (N_15887,N_8906,N_11960);
nand U15888 (N_15888,N_11419,N_11824);
or U15889 (N_15889,N_8753,N_8390);
nand U15890 (N_15890,N_11130,N_11409);
nor U15891 (N_15891,N_8324,N_10041);
or U15892 (N_15892,N_8292,N_10231);
and U15893 (N_15893,N_10145,N_10118);
nor U15894 (N_15894,N_11615,N_9702);
and U15895 (N_15895,N_8017,N_9759);
and U15896 (N_15896,N_10741,N_8613);
nand U15897 (N_15897,N_11787,N_10893);
or U15898 (N_15898,N_9100,N_8805);
and U15899 (N_15899,N_8944,N_9139);
nor U15900 (N_15900,N_9414,N_10909);
or U15901 (N_15901,N_8308,N_10408);
nand U15902 (N_15902,N_10635,N_8559);
nand U15903 (N_15903,N_11635,N_9615);
or U15904 (N_15904,N_8875,N_9888);
nand U15905 (N_15905,N_10806,N_8144);
nor U15906 (N_15906,N_10224,N_11922);
or U15907 (N_15907,N_10472,N_9056);
or U15908 (N_15908,N_11055,N_8191);
or U15909 (N_15909,N_10211,N_8240);
and U15910 (N_15910,N_9831,N_8956);
or U15911 (N_15911,N_9949,N_9205);
xnor U15912 (N_15912,N_10550,N_10136);
and U15913 (N_15913,N_9995,N_9495);
nand U15914 (N_15914,N_10785,N_8317);
nor U15915 (N_15915,N_10420,N_11332);
nand U15916 (N_15916,N_11780,N_11282);
or U15917 (N_15917,N_9554,N_11745);
nor U15918 (N_15918,N_8690,N_11604);
nand U15919 (N_15919,N_9484,N_9218);
or U15920 (N_15920,N_10222,N_11455);
nor U15921 (N_15921,N_8048,N_10228);
nand U15922 (N_15922,N_8062,N_11420);
nor U15923 (N_15923,N_10930,N_11267);
nand U15924 (N_15924,N_9067,N_9982);
or U15925 (N_15925,N_8329,N_9465);
and U15926 (N_15926,N_8404,N_11958);
nor U15927 (N_15927,N_10452,N_11702);
and U15928 (N_15928,N_10854,N_11360);
or U15929 (N_15929,N_11371,N_10346);
nor U15930 (N_15930,N_11748,N_9930);
and U15931 (N_15931,N_11211,N_11239);
and U15932 (N_15932,N_11692,N_9959);
xor U15933 (N_15933,N_8377,N_9611);
and U15934 (N_15934,N_8548,N_11523);
or U15935 (N_15935,N_11423,N_8168);
nand U15936 (N_15936,N_11798,N_8745);
or U15937 (N_15937,N_8548,N_10297);
and U15938 (N_15938,N_10491,N_11939);
nor U15939 (N_15939,N_9905,N_10071);
xnor U15940 (N_15940,N_9548,N_8806);
xor U15941 (N_15941,N_8705,N_10922);
nand U15942 (N_15942,N_8002,N_11219);
or U15943 (N_15943,N_11497,N_9167);
nor U15944 (N_15944,N_10904,N_9653);
and U15945 (N_15945,N_9542,N_10133);
nand U15946 (N_15946,N_10393,N_9730);
or U15947 (N_15947,N_10080,N_9335);
nor U15948 (N_15948,N_8250,N_8360);
xnor U15949 (N_15949,N_9198,N_8107);
nor U15950 (N_15950,N_9294,N_10747);
or U15951 (N_15951,N_10979,N_10776);
nor U15952 (N_15952,N_9242,N_9818);
and U15953 (N_15953,N_8060,N_8049);
and U15954 (N_15954,N_11103,N_11045);
nand U15955 (N_15955,N_8914,N_9426);
and U15956 (N_15956,N_8248,N_8947);
or U15957 (N_15957,N_10851,N_8395);
nand U15958 (N_15958,N_8229,N_8841);
nand U15959 (N_15959,N_11288,N_10782);
and U15960 (N_15960,N_11097,N_8903);
and U15961 (N_15961,N_8853,N_10373);
and U15962 (N_15962,N_10710,N_11946);
xor U15963 (N_15963,N_11172,N_11013);
and U15964 (N_15964,N_9150,N_9596);
or U15965 (N_15965,N_11744,N_8903);
nor U15966 (N_15966,N_11838,N_8839);
or U15967 (N_15967,N_11958,N_9697);
or U15968 (N_15968,N_9687,N_11971);
nand U15969 (N_15969,N_8781,N_11299);
xnor U15970 (N_15970,N_8731,N_11980);
and U15971 (N_15971,N_9191,N_8503);
xnor U15972 (N_15972,N_9846,N_10779);
and U15973 (N_15973,N_9405,N_11185);
nand U15974 (N_15974,N_11759,N_10987);
nor U15975 (N_15975,N_9501,N_8527);
and U15976 (N_15976,N_9842,N_11592);
and U15977 (N_15977,N_11028,N_8143);
nor U15978 (N_15978,N_8744,N_9783);
nand U15979 (N_15979,N_8843,N_10530);
and U15980 (N_15980,N_10206,N_8587);
or U15981 (N_15981,N_8753,N_11829);
or U15982 (N_15982,N_11521,N_8822);
nor U15983 (N_15983,N_9110,N_8356);
or U15984 (N_15984,N_9181,N_11998);
nor U15985 (N_15985,N_9971,N_8152);
and U15986 (N_15986,N_9803,N_8490);
nand U15987 (N_15987,N_8543,N_10764);
nor U15988 (N_15988,N_9008,N_10873);
and U15989 (N_15989,N_9048,N_10154);
and U15990 (N_15990,N_9231,N_11208);
nor U15991 (N_15991,N_9173,N_10404);
and U15992 (N_15992,N_9798,N_8081);
or U15993 (N_15993,N_9932,N_9489);
or U15994 (N_15994,N_9577,N_8146);
nand U15995 (N_15995,N_8253,N_9217);
and U15996 (N_15996,N_10929,N_11723);
and U15997 (N_15997,N_10268,N_8518);
and U15998 (N_15998,N_9507,N_10805);
and U15999 (N_15999,N_9534,N_11980);
and U16000 (N_16000,N_13262,N_15555);
and U16001 (N_16001,N_14214,N_12687);
and U16002 (N_16002,N_15642,N_12293);
nor U16003 (N_16003,N_12879,N_12655);
nor U16004 (N_16004,N_13475,N_12104);
xor U16005 (N_16005,N_12114,N_15855);
nor U16006 (N_16006,N_12565,N_13708);
or U16007 (N_16007,N_15711,N_13014);
nand U16008 (N_16008,N_13560,N_15184);
and U16009 (N_16009,N_14169,N_13462);
nor U16010 (N_16010,N_14476,N_14581);
nand U16011 (N_16011,N_15636,N_12092);
and U16012 (N_16012,N_15274,N_15540);
nor U16013 (N_16013,N_12700,N_13709);
nand U16014 (N_16014,N_12434,N_13960);
nor U16015 (N_16015,N_15394,N_13276);
nand U16016 (N_16016,N_15254,N_15877);
and U16017 (N_16017,N_12238,N_15099);
and U16018 (N_16018,N_15885,N_12040);
nor U16019 (N_16019,N_14350,N_14210);
nand U16020 (N_16020,N_12373,N_13627);
and U16021 (N_16021,N_14399,N_12986);
nor U16022 (N_16022,N_14614,N_12522);
and U16023 (N_16023,N_12850,N_14437);
or U16024 (N_16024,N_13691,N_12997);
nand U16025 (N_16025,N_15998,N_15217);
nand U16026 (N_16026,N_12983,N_12604);
nand U16027 (N_16027,N_13530,N_14044);
or U16028 (N_16028,N_12017,N_13765);
or U16029 (N_16029,N_12798,N_14973);
or U16030 (N_16030,N_12710,N_12322);
nand U16031 (N_16031,N_15926,N_15708);
and U16032 (N_16032,N_13211,N_15668);
and U16033 (N_16033,N_13865,N_13784);
nor U16034 (N_16034,N_15408,N_13194);
and U16035 (N_16035,N_12306,N_13569);
nand U16036 (N_16036,N_12985,N_14424);
and U16037 (N_16037,N_13048,N_15065);
nand U16038 (N_16038,N_14982,N_15537);
xor U16039 (N_16039,N_14294,N_15581);
and U16040 (N_16040,N_12180,N_12623);
and U16041 (N_16041,N_15045,N_14160);
nor U16042 (N_16042,N_12569,N_12628);
nor U16043 (N_16043,N_15612,N_15559);
nand U16044 (N_16044,N_13458,N_12724);
nand U16045 (N_16045,N_12036,N_14524);
nor U16046 (N_16046,N_13077,N_12935);
and U16047 (N_16047,N_12463,N_13750);
nor U16048 (N_16048,N_12384,N_14019);
or U16049 (N_16049,N_12122,N_12493);
nand U16050 (N_16050,N_15155,N_13093);
nor U16051 (N_16051,N_15019,N_15788);
or U16052 (N_16052,N_15063,N_13221);
nor U16053 (N_16053,N_12508,N_15978);
nand U16054 (N_16054,N_14027,N_14124);
and U16055 (N_16055,N_12491,N_12460);
nor U16056 (N_16056,N_13894,N_15989);
and U16057 (N_16057,N_14251,N_14109);
xor U16058 (N_16058,N_13380,N_15759);
and U16059 (N_16059,N_14777,N_13264);
xnor U16060 (N_16060,N_14232,N_13736);
nor U16061 (N_16061,N_14346,N_14332);
or U16062 (N_16062,N_14235,N_12324);
and U16063 (N_16063,N_13630,N_12366);
or U16064 (N_16064,N_14444,N_13634);
and U16065 (N_16065,N_14937,N_14928);
nand U16066 (N_16066,N_14551,N_15143);
xor U16067 (N_16067,N_13416,N_12679);
nand U16068 (N_16068,N_13557,N_14688);
nor U16069 (N_16069,N_15638,N_15084);
or U16070 (N_16070,N_12130,N_15589);
nand U16071 (N_16071,N_12099,N_12530);
nand U16072 (N_16072,N_15398,N_14113);
or U16073 (N_16073,N_15022,N_12119);
nor U16074 (N_16074,N_12657,N_15532);
nand U16075 (N_16075,N_14296,N_12572);
nand U16076 (N_16076,N_14366,N_15734);
and U16077 (N_16077,N_12450,N_12472);
or U16078 (N_16078,N_12312,N_15837);
or U16079 (N_16079,N_14550,N_14541);
or U16080 (N_16080,N_14188,N_13379);
nor U16081 (N_16081,N_12348,N_13995);
and U16082 (N_16082,N_14539,N_14711);
nor U16083 (N_16083,N_13711,N_13354);
or U16084 (N_16084,N_14778,N_15058);
or U16085 (N_16085,N_13689,N_12617);
or U16086 (N_16086,N_13655,N_12898);
and U16087 (N_16087,N_15324,N_12095);
or U16088 (N_16088,N_15874,N_15516);
or U16089 (N_16089,N_15320,N_13695);
nand U16090 (N_16090,N_15315,N_14261);
or U16091 (N_16091,N_13968,N_15384);
xnor U16092 (N_16092,N_15270,N_15088);
xnor U16093 (N_16093,N_13269,N_14940);
nand U16094 (N_16094,N_13386,N_13152);
nor U16095 (N_16095,N_12506,N_13028);
and U16096 (N_16096,N_12371,N_13374);
and U16097 (N_16097,N_13329,N_15296);
or U16098 (N_16098,N_15517,N_13297);
and U16099 (N_16099,N_14662,N_15769);
or U16100 (N_16100,N_15389,N_14475);
or U16101 (N_16101,N_15493,N_14865);
nor U16102 (N_16102,N_14193,N_15629);
and U16103 (N_16103,N_14872,N_13722);
and U16104 (N_16104,N_12631,N_15796);
nor U16105 (N_16105,N_15829,N_15840);
nor U16106 (N_16106,N_12034,N_12905);
nand U16107 (N_16107,N_14743,N_13767);
or U16108 (N_16108,N_12767,N_15042);
nor U16109 (N_16109,N_12200,N_14736);
nor U16110 (N_16110,N_14587,N_13710);
nand U16111 (N_16111,N_15003,N_15945);
or U16112 (N_16112,N_14664,N_13758);
or U16113 (N_16113,N_13472,N_12599);
nor U16114 (N_16114,N_13464,N_15176);
or U16115 (N_16115,N_13398,N_15204);
and U16116 (N_16116,N_14230,N_15691);
xnor U16117 (N_16117,N_13236,N_15325);
nor U16118 (N_16118,N_14754,N_12302);
and U16119 (N_16119,N_14161,N_15287);
and U16120 (N_16120,N_14801,N_13017);
and U16121 (N_16121,N_12896,N_12964);
nand U16122 (N_16122,N_15776,N_15009);
nor U16123 (N_16123,N_14384,N_15294);
nand U16124 (N_16124,N_15103,N_15451);
and U16125 (N_16125,N_12390,N_13666);
nor U16126 (N_16126,N_14843,N_15064);
and U16127 (N_16127,N_13195,N_13799);
or U16128 (N_16128,N_12732,N_15562);
or U16129 (N_16129,N_13579,N_15651);
xnor U16130 (N_16130,N_15105,N_14836);
and U16131 (N_16131,N_13278,N_12882);
or U16132 (N_16132,N_12151,N_14717);
nand U16133 (N_16133,N_12581,N_15900);
nor U16134 (N_16134,N_14225,N_12266);
nor U16135 (N_16135,N_14407,N_14381);
and U16136 (N_16136,N_12598,N_15180);
and U16137 (N_16137,N_14927,N_15928);
nor U16138 (N_16138,N_15104,N_14988);
or U16139 (N_16139,N_15052,N_15085);
xor U16140 (N_16140,N_15136,N_13050);
xor U16141 (N_16141,N_14680,N_13690);
and U16142 (N_16142,N_14626,N_15601);
and U16143 (N_16143,N_14157,N_15725);
nor U16144 (N_16144,N_13538,N_15539);
and U16145 (N_16145,N_15054,N_14888);
nand U16146 (N_16146,N_12789,N_13171);
xor U16147 (N_16147,N_14723,N_13218);
or U16148 (N_16148,N_14187,N_14395);
nor U16149 (N_16149,N_14572,N_13571);
and U16150 (N_16150,N_13324,N_14555);
nand U16151 (N_16151,N_14439,N_14410);
or U16152 (N_16152,N_13332,N_12664);
and U16153 (N_16153,N_12795,N_14816);
nand U16154 (N_16154,N_12564,N_14067);
or U16155 (N_16155,N_12072,N_14315);
or U16156 (N_16156,N_13769,N_15605);
and U16157 (N_16157,N_12396,N_15610);
nand U16158 (N_16158,N_12108,N_13613);
or U16159 (N_16159,N_13544,N_12287);
or U16160 (N_16160,N_12411,N_14039);
or U16161 (N_16161,N_14004,N_14164);
and U16162 (N_16162,N_13346,N_12494);
nor U16163 (N_16163,N_15810,N_15674);
nand U16164 (N_16164,N_15859,N_13866);
nand U16165 (N_16165,N_15005,N_13364);
nor U16166 (N_16166,N_13820,N_13284);
xor U16167 (N_16167,N_15972,N_13745);
or U16168 (N_16168,N_14033,N_13577);
nand U16169 (N_16169,N_13759,N_15479);
or U16170 (N_16170,N_12856,N_14518);
nand U16171 (N_16171,N_12006,N_12889);
or U16172 (N_16172,N_12261,N_12027);
nor U16173 (N_16173,N_15750,N_13921);
or U16174 (N_16174,N_15038,N_13441);
or U16175 (N_16175,N_14460,N_14750);
nand U16176 (N_16176,N_14716,N_13053);
xor U16177 (N_16177,N_12961,N_12003);
and U16178 (N_16178,N_13805,N_12298);
xnor U16179 (N_16179,N_15513,N_12982);
and U16180 (N_16180,N_12131,N_12154);
or U16181 (N_16181,N_12023,N_13940);
xor U16182 (N_16182,N_13804,N_13790);
nand U16183 (N_16183,N_13562,N_12519);
nand U16184 (N_16184,N_12821,N_15604);
xor U16185 (N_16185,N_12759,N_12216);
nand U16186 (N_16186,N_12064,N_14172);
nor U16187 (N_16187,N_14922,N_15399);
nand U16188 (N_16188,N_14564,N_14771);
or U16189 (N_16189,N_13643,N_15223);
and U16190 (N_16190,N_14672,N_14069);
or U16191 (N_16191,N_14668,N_15391);
or U16192 (N_16192,N_14563,N_15962);
nand U16193 (N_16193,N_14725,N_12652);
and U16194 (N_16194,N_14738,N_12651);
or U16195 (N_16195,N_13319,N_12280);
and U16196 (N_16196,N_14012,N_14337);
and U16197 (N_16197,N_14496,N_12164);
or U16198 (N_16198,N_13636,N_15069);
nor U16199 (N_16199,N_12041,N_14180);
nand U16200 (N_16200,N_15994,N_15682);
and U16201 (N_16201,N_13788,N_15904);
or U16202 (N_16202,N_14241,N_15655);
nor U16203 (N_16203,N_13253,N_14628);
nand U16204 (N_16204,N_13594,N_12977);
and U16205 (N_16205,N_14093,N_15309);
nand U16206 (N_16206,N_14755,N_13372);
nand U16207 (N_16207,N_13725,N_15806);
xnor U16208 (N_16208,N_13556,N_12193);
nand U16209 (N_16209,N_13434,N_13282);
nand U16210 (N_16210,N_15158,N_13138);
or U16211 (N_16211,N_12455,N_15449);
or U16212 (N_16212,N_15663,N_12816);
nor U16213 (N_16213,N_12735,N_15492);
nand U16214 (N_16214,N_13308,N_14594);
and U16215 (N_16215,N_14154,N_12536);
or U16216 (N_16216,N_12362,N_15267);
nand U16217 (N_16217,N_13299,N_12634);
nor U16218 (N_16218,N_13825,N_12296);
nor U16219 (N_16219,N_15372,N_14508);
nor U16220 (N_16220,N_13290,N_12842);
nor U16221 (N_16221,N_13624,N_13220);
nor U16222 (N_16222,N_15529,N_12899);
and U16223 (N_16223,N_14657,N_13295);
or U16224 (N_16224,N_12421,N_14600);
or U16225 (N_16225,N_12190,N_13701);
nand U16226 (N_16226,N_15863,N_15355);
nand U16227 (N_16227,N_14175,N_12517);
nand U16228 (N_16228,N_13522,N_13687);
xor U16229 (N_16229,N_12205,N_14696);
or U16230 (N_16230,N_13776,N_14469);
xnor U16231 (N_16231,N_12063,N_15758);
nor U16232 (N_16232,N_15474,N_15654);
and U16233 (N_16233,N_15279,N_12400);
xnor U16234 (N_16234,N_14867,N_12538);
xor U16235 (N_16235,N_15293,N_12333);
nand U16236 (N_16236,N_14629,N_13589);
or U16237 (N_16237,N_13551,N_14698);
or U16238 (N_16238,N_12458,N_12911);
nand U16239 (N_16239,N_15077,N_15377);
nor U16240 (N_16240,N_13174,N_14844);
and U16241 (N_16241,N_14009,N_14758);
nor U16242 (N_16242,N_15277,N_15896);
nor U16243 (N_16243,N_14284,N_14719);
nand U16244 (N_16244,N_12271,N_14431);
or U16245 (N_16245,N_14890,N_15114);
or U16246 (N_16246,N_15177,N_15478);
nand U16247 (N_16247,N_14152,N_13659);
or U16248 (N_16248,N_14445,N_15809);
nand U16249 (N_16249,N_14312,N_14921);
or U16250 (N_16250,N_15831,N_12320);
or U16251 (N_16251,N_15603,N_14860);
or U16252 (N_16252,N_13548,N_13239);
or U16253 (N_16253,N_13490,N_15422);
and U16254 (N_16254,N_15954,N_14082);
nand U16255 (N_16255,N_13049,N_15232);
nand U16256 (N_16256,N_14279,N_14919);
xnor U16257 (N_16257,N_14603,N_15059);
nor U16258 (N_16258,N_13588,N_14025);
and U16259 (N_16259,N_14493,N_12738);
xor U16260 (N_16260,N_15801,N_12250);
xor U16261 (N_16261,N_13059,N_12885);
xnor U16262 (N_16262,N_15870,N_14499);
xor U16263 (N_16263,N_14257,N_13073);
or U16264 (N_16264,N_15897,N_14854);
or U16265 (N_16265,N_12689,N_13519);
and U16266 (N_16266,N_14545,N_15000);
nor U16267 (N_16267,N_12674,N_13012);
xnor U16268 (N_16268,N_13749,N_12413);
or U16269 (N_16269,N_12345,N_15585);
nand U16270 (N_16270,N_12117,N_15224);
or U16271 (N_16271,N_15905,N_12775);
nor U16272 (N_16272,N_13546,N_14933);
and U16273 (N_16273,N_15250,N_15312);
and U16274 (N_16274,N_12260,N_15843);
or U16275 (N_16275,N_13109,N_13186);
and U16276 (N_16276,N_13629,N_13575);
nand U16277 (N_16277,N_14013,N_15291);
xor U16278 (N_16278,N_14764,N_13219);
or U16279 (N_16279,N_12409,N_13614);
nand U16280 (N_16280,N_14002,N_15556);
nand U16281 (N_16281,N_13696,N_14578);
and U16282 (N_16282,N_12445,N_14123);
or U16283 (N_16283,N_14760,N_12832);
and U16284 (N_16284,N_12231,N_14980);
nand U16285 (N_16285,N_15927,N_12559);
nand U16286 (N_16286,N_13281,N_14803);
nor U16287 (N_16287,N_12834,N_12912);
or U16288 (N_16288,N_12120,N_13395);
xor U16289 (N_16289,N_13367,N_14861);
nand U16290 (N_16290,N_14868,N_15813);
or U16291 (N_16291,N_12066,N_15262);
nor U16292 (N_16292,N_14273,N_14838);
nand U16293 (N_16293,N_15965,N_12810);
and U16294 (N_16294,N_14994,N_14059);
and U16295 (N_16295,N_14404,N_15332);
nor U16296 (N_16296,N_14757,N_14378);
nor U16297 (N_16297,N_15545,N_15717);
and U16298 (N_16298,N_13432,N_15096);
and U16299 (N_16299,N_14878,N_13792);
and U16300 (N_16300,N_14143,N_15784);
and U16301 (N_16301,N_12369,N_14248);
nor U16302 (N_16302,N_14787,N_15111);
nor U16303 (N_16303,N_14268,N_15323);
xnor U16304 (N_16304,N_14811,N_13371);
or U16305 (N_16305,N_12263,N_15134);
nor U16306 (N_16306,N_15338,N_14560);
or U16307 (N_16307,N_14132,N_15847);
and U16308 (N_16308,N_14321,N_15812);
nand U16309 (N_16309,N_15402,N_13936);
and U16310 (N_16310,N_12115,N_15265);
or U16311 (N_16311,N_15720,N_13491);
nor U16312 (N_16312,N_14828,N_12275);
nand U16313 (N_16313,N_14529,N_12562);
and U16314 (N_16314,N_13227,N_12644);
nor U16315 (N_16315,N_14526,N_12186);
nand U16316 (N_16316,N_13352,N_12550);
nor U16317 (N_16317,N_13561,N_14609);
nor U16318 (N_16318,N_13809,N_15359);
or U16319 (N_16319,N_13772,N_14436);
nor U16320 (N_16320,N_12342,N_14782);
nand U16321 (N_16321,N_15853,N_15160);
or U16322 (N_16322,N_12107,N_15047);
or U16323 (N_16323,N_12953,N_13274);
or U16324 (N_16324,N_15805,N_14885);
xor U16325 (N_16325,N_15698,N_14416);
or U16326 (N_16326,N_13723,N_12235);
nand U16327 (N_16327,N_14580,N_12317);
nand U16328 (N_16328,N_15067,N_15471);
nor U16329 (N_16329,N_13656,N_14452);
xor U16330 (N_16330,N_12234,N_13440);
and U16331 (N_16331,N_13401,N_12430);
and U16332 (N_16332,N_12267,N_13383);
and U16333 (N_16333,N_13943,N_14915);
or U16334 (N_16334,N_12612,N_14162);
or U16335 (N_16335,N_12800,N_13535);
and U16336 (N_16336,N_12436,N_12620);
nor U16337 (N_16337,N_12497,N_13249);
and U16338 (N_16338,N_14682,N_14050);
or U16339 (N_16339,N_14791,N_14615);
nand U16340 (N_16340,N_15571,N_13140);
nor U16341 (N_16341,N_14610,N_14330);
nand U16342 (N_16342,N_15531,N_15774);
or U16343 (N_16343,N_13078,N_15960);
and U16344 (N_16344,N_12464,N_14105);
nor U16345 (N_16345,N_13539,N_15369);
nand U16346 (N_16346,N_12932,N_14944);
xnor U16347 (N_16347,N_13543,N_13713);
nand U16348 (N_16348,N_13518,N_15697);
and U16349 (N_16349,N_13056,N_12699);
and U16350 (N_16350,N_12214,N_12929);
or U16351 (N_16351,N_14627,N_12815);
nor U16352 (N_16352,N_13256,N_15413);
or U16353 (N_16353,N_13181,N_12793);
nor U16354 (N_16354,N_12385,N_14507);
and U16355 (N_16355,N_14229,N_14139);
nor U16356 (N_16356,N_14075,N_15071);
or U16357 (N_16357,N_13974,N_14969);
and U16358 (N_16358,N_12157,N_13307);
or U16359 (N_16359,N_14765,N_15252);
or U16360 (N_16360,N_12760,N_15983);
xnor U16361 (N_16361,N_13085,N_13977);
and U16362 (N_16362,N_15519,N_15856);
nor U16363 (N_16363,N_15598,N_15013);
nor U16364 (N_16364,N_13847,N_14849);
nand U16365 (N_16365,N_14405,N_12925);
or U16366 (N_16366,N_15898,N_14911);
xor U16367 (N_16367,N_13810,N_15973);
nor U16368 (N_16368,N_15857,N_12482);
and U16369 (N_16369,N_13454,N_13497);
or U16370 (N_16370,N_15771,N_14652);
nand U16371 (N_16371,N_12067,N_15374);
and U16372 (N_16372,N_12370,N_12919);
and U16373 (N_16373,N_13243,N_13951);
nand U16374 (N_16374,N_15615,N_14544);
or U16375 (N_16375,N_14054,N_12148);
and U16376 (N_16376,N_14365,N_15406);
nand U16377 (N_16377,N_12326,N_15057);
and U16378 (N_16378,N_12129,N_15373);
nor U16379 (N_16379,N_14830,N_13517);
nor U16380 (N_16380,N_13466,N_13570);
nand U16381 (N_16381,N_14464,N_14745);
and U16382 (N_16382,N_12062,N_13890);
and U16383 (N_16383,N_13950,N_13648);
nand U16384 (N_16384,N_13342,N_15251);
nand U16385 (N_16385,N_14530,N_13699);
and U16386 (N_16386,N_13859,N_12183);
and U16387 (N_16387,N_12703,N_12866);
nand U16388 (N_16388,N_14348,N_15582);
and U16389 (N_16389,N_12239,N_15919);
or U16390 (N_16390,N_15652,N_13633);
nand U16391 (N_16391,N_14037,N_12744);
nand U16392 (N_16392,N_13787,N_15376);
nor U16393 (N_16393,N_15040,N_14449);
and U16394 (N_16394,N_14130,N_14114);
nand U16395 (N_16395,N_14303,N_12415);
and U16396 (N_16396,N_13316,N_13121);
or U16397 (N_16397,N_13309,N_12616);
or U16398 (N_16398,N_14118,N_14417);
nand U16399 (N_16399,N_15157,N_13143);
or U16400 (N_16400,N_13157,N_15347);
nor U16401 (N_16401,N_13999,N_15817);
xor U16402 (N_16402,N_14515,N_15350);
or U16403 (N_16403,N_12762,N_15525);
nand U16404 (N_16404,N_15802,N_15838);
nand U16405 (N_16405,N_13375,N_13118);
and U16406 (N_16406,N_15073,N_15185);
xnor U16407 (N_16407,N_14136,N_12080);
xnor U16408 (N_16408,N_15387,N_14989);
nor U16409 (N_16409,N_15261,N_14855);
and U16410 (N_16410,N_13133,N_13631);
nand U16411 (N_16411,N_15915,N_12958);
nor U16412 (N_16412,N_14343,N_15661);
and U16413 (N_16413,N_13311,N_15895);
xnor U16414 (N_16414,N_12213,N_12922);
or U16415 (N_16415,N_12025,N_12050);
nand U16416 (N_16416,N_14274,N_13148);
nor U16417 (N_16417,N_13761,N_12259);
nand U16418 (N_16418,N_14207,N_14480);
nand U16419 (N_16419,N_14074,N_15488);
and U16420 (N_16420,N_13417,N_14377);
nor U16421 (N_16421,N_15154,N_13891);
nand U16422 (N_16422,N_14371,N_13675);
nor U16423 (N_16423,N_14055,N_13495);
nor U16424 (N_16424,N_12142,N_13327);
nand U16425 (N_16425,N_15221,N_15816);
nor U16426 (N_16426,N_15302,N_13353);
nand U16427 (N_16427,N_12304,N_13964);
or U16428 (N_16428,N_13889,N_13326);
xor U16429 (N_16429,N_15140,N_14503);
xor U16430 (N_16430,N_13089,N_13294);
nor U16431 (N_16431,N_14511,N_13492);
and U16432 (N_16432,N_15730,N_14997);
xnor U16433 (N_16433,N_14670,N_13875);
and U16434 (N_16434,N_13010,N_14797);
nor U16435 (N_16435,N_12927,N_12774);
nor U16436 (N_16436,N_13529,N_14354);
xnor U16437 (N_16437,N_13452,N_15587);
nand U16438 (N_16438,N_14275,N_13487);
nor U16439 (N_16439,N_14457,N_15886);
or U16440 (N_16440,N_13993,N_12407);
or U16441 (N_16441,N_14807,N_12523);
nor U16442 (N_16442,N_15036,N_14463);
xor U16443 (N_16443,N_12089,N_14673);
nor U16444 (N_16444,N_12624,N_15716);
or U16445 (N_16445,N_14642,N_13734);
xnor U16446 (N_16446,N_12079,N_14697);
xnor U16447 (N_16447,N_15777,N_15521);
nor U16448 (N_16448,N_15509,N_14490);
nor U16449 (N_16449,N_15191,N_13240);
nand U16450 (N_16450,N_13031,N_12747);
and U16451 (N_16451,N_14038,N_12989);
or U16452 (N_16452,N_12736,N_14254);
xnor U16453 (N_16453,N_14032,N_15446);
and U16454 (N_16454,N_13173,N_13261);
nor U16455 (N_16455,N_13978,N_15091);
or U16456 (N_16456,N_14525,N_12167);
or U16457 (N_16457,N_14644,N_15530);
xnor U16458 (N_16458,N_15053,N_12967);
nor U16459 (N_16459,N_12996,N_15095);
xnor U16460 (N_16460,N_13926,N_14049);
and U16461 (N_16461,N_14658,N_14546);
nor U16462 (N_16462,N_15272,N_12966);
nand U16463 (N_16463,N_14993,N_15735);
and U16464 (N_16464,N_15845,N_14800);
and U16465 (N_16465,N_15358,N_12470);
and U16466 (N_16466,N_13151,N_13747);
and U16467 (N_16467,N_15920,N_13861);
nand U16468 (N_16468,N_14168,N_15865);
and U16469 (N_16469,N_12588,N_14373);
or U16470 (N_16470,N_14338,N_13241);
nor U16471 (N_16471,N_14316,N_14899);
and U16472 (N_16472,N_13418,N_15420);
xnor U16473 (N_16473,N_14770,N_13124);
nor U16474 (N_16474,N_12602,N_13664);
or U16475 (N_16475,N_12196,N_13979);
nor U16476 (N_16476,N_12827,N_14900);
nand U16477 (N_16477,N_13929,N_13834);
or U16478 (N_16478,N_14308,N_14538);
nor U16479 (N_16479,N_15984,N_15706);
nand U16480 (N_16480,N_14097,N_14116);
nor U16481 (N_16481,N_13632,N_14641);
or U16482 (N_16482,N_12875,N_13549);
xnor U16483 (N_16483,N_15565,N_14558);
nand U16484 (N_16484,N_13468,N_13339);
nand U16485 (N_16485,N_12558,N_12979);
nor U16486 (N_16486,N_12357,N_14559);
nor U16487 (N_16487,N_14491,N_14829);
and U16488 (N_16488,N_12907,N_14506);
and U16489 (N_16489,N_15620,N_12663);
and U16490 (N_16490,N_15861,N_15193);
nor U16491 (N_16491,N_15676,N_15902);
nor U16492 (N_16492,N_13873,N_12817);
nand U16493 (N_16493,N_14396,N_13945);
nand U16494 (N_16494,N_14845,N_13363);
nor U16495 (N_16495,N_12393,N_14336);
nor U16496 (N_16496,N_14896,N_13838);
or U16497 (N_16497,N_13681,N_12016);
xnor U16498 (N_16498,N_14472,N_15704);
nor U16499 (N_16499,N_13203,N_14071);
and U16500 (N_16500,N_14623,N_14917);
xor U16501 (N_16501,N_14542,N_13502);
and U16502 (N_16502,N_12686,N_13563);
nor U16503 (N_16503,N_13545,N_14774);
and U16504 (N_16504,N_14212,N_13499);
nor U16505 (N_16505,N_14471,N_13060);
and U16506 (N_16506,N_12968,N_12221);
nor U16507 (N_16507,N_14477,N_12719);
or U16508 (N_16508,N_12059,N_15129);
nor U16509 (N_16509,N_12993,N_15694);
nand U16510 (N_16510,N_14951,N_14356);
or U16511 (N_16511,N_13135,N_15766);
or U16512 (N_16512,N_15196,N_12894);
nor U16513 (N_16513,N_14078,N_13226);
nand U16514 (N_16514,N_13510,N_14253);
nor U16515 (N_16515,N_14793,N_12223);
or U16516 (N_16516,N_15156,N_13110);
nand U16517 (N_16517,N_13982,N_14191);
and U16518 (N_16518,N_12401,N_12553);
and U16519 (N_16519,N_13410,N_13178);
nand U16520 (N_16520,N_14149,N_13429);
or U16521 (N_16521,N_15429,N_15510);
xnor U16522 (N_16522,N_12728,N_12483);
nand U16523 (N_16523,N_13465,N_12291);
xor U16524 (N_16524,N_15039,N_15236);
or U16525 (N_16525,N_15343,N_13330);
nand U16526 (N_16526,N_13168,N_12255);
nor U16527 (N_16527,N_15570,N_13369);
xor U16528 (N_16528,N_13323,N_13074);
and U16529 (N_16529,N_12886,N_13163);
nor U16530 (N_16530,N_12920,N_15178);
nand U16531 (N_16531,N_15660,N_13494);
and U16532 (N_16532,N_14466,N_12669);
nand U16533 (N_16533,N_15308,N_12551);
or U16534 (N_16534,N_14945,N_15317);
nor U16535 (N_16535,N_12857,N_12893);
nor U16536 (N_16536,N_13783,N_12382);
nand U16537 (N_16537,N_13564,N_15127);
nor U16538 (N_16538,N_13822,N_12465);
nand U16539 (N_16539,N_14624,N_15658);
and U16540 (N_16540,N_12228,N_13607);
or U16541 (N_16541,N_14533,N_12484);
nor U16542 (N_16542,N_13382,N_15222);
xor U16543 (N_16543,N_13966,N_15592);
and U16544 (N_16544,N_12397,N_12659);
nand U16545 (N_16545,N_12363,N_14926);
or U16546 (N_16546,N_14129,N_15700);
nor U16547 (N_16547,N_14513,N_12341);
xor U16548 (N_16548,N_13896,N_13126);
or U16549 (N_16549,N_14734,N_15481);
and U16550 (N_16550,N_15976,N_12145);
nor U16551 (N_16551,N_14965,N_14984);
and U16552 (N_16552,N_14950,N_15008);
and U16553 (N_16553,N_13892,N_14647);
and U16554 (N_16554,N_12956,N_15056);
and U16555 (N_16555,N_13455,N_13242);
or U16556 (N_16556,N_12452,N_12954);
nand U16557 (N_16557,N_15079,N_15147);
nor U16558 (N_16558,N_13191,N_12930);
nor U16559 (N_16559,N_14048,N_12704);
nor U16560 (N_16560,N_15220,N_13581);
or U16561 (N_16561,N_12031,N_14380);
and U16562 (N_16562,N_15242,N_15901);
nand U16563 (N_16563,N_14996,N_12057);
nor U16564 (N_16564,N_12078,N_13443);
or U16565 (N_16565,N_12751,N_12227);
nor U16566 (N_16566,N_12162,N_13298);
nand U16567 (N_16567,N_12880,N_14454);
nor U16568 (N_16568,N_12014,N_13478);
or U16569 (N_16569,N_15899,N_13623);
or U16570 (N_16570,N_13640,N_15740);
and U16571 (N_16571,N_13356,N_13394);
nor U16572 (N_16572,N_14474,N_13423);
nand U16573 (N_16573,N_13373,N_15664);
nand U16574 (N_16574,N_13880,N_15755);
or U16575 (N_16575,N_15688,N_12220);
nand U16576 (N_16576,N_15331,N_14107);
and U16577 (N_16577,N_12999,N_13660);
or U16578 (N_16578,N_13435,N_14318);
and U16579 (N_16579,N_12546,N_12047);
nand U16580 (N_16580,N_13819,N_14411);
or U16581 (N_16581,N_13208,N_14731);
nand U16582 (N_16582,N_14947,N_14884);
xnor U16583 (N_16583,N_14741,N_14656);
nand U16584 (N_16584,N_15923,N_14661);
nand U16585 (N_16585,N_13961,N_12189);
and U16586 (N_16586,N_13228,N_13855);
or U16587 (N_16587,N_12269,N_15830);
nand U16588 (N_16588,N_12177,N_12096);
or U16589 (N_16589,N_12124,N_15439);
nor U16590 (N_16590,N_15454,N_15793);
and U16591 (N_16591,N_13034,N_14649);
and U16592 (N_16592,N_15741,N_14790);
xor U16593 (N_16593,N_13931,N_14825);
nor U16594 (N_16594,N_15142,N_12941);
or U16595 (N_16595,N_15616,N_12427);
nand U16596 (N_16596,N_13214,N_12159);
nand U16597 (N_16597,N_14470,N_14281);
xnor U16598 (N_16598,N_15554,N_14270);
nor U16599 (N_16599,N_13130,N_13851);
nand U16600 (N_16600,N_12822,N_15245);
nor U16601 (N_16601,N_12224,N_15113);
nand U16602 (N_16602,N_13637,N_12683);
nor U16603 (N_16603,N_13948,N_13084);
nor U16604 (N_16604,N_14759,N_14280);
or U16605 (N_16605,N_15869,N_12392);
nand U16606 (N_16606,N_15753,N_12376);
or U16607 (N_16607,N_13900,N_15050);
xor U16608 (N_16608,N_13515,N_14846);
nand U16609 (N_16609,N_14403,N_12307);
nor U16610 (N_16610,N_14324,N_14601);
nand U16611 (N_16611,N_15285,N_12877);
nand U16612 (N_16612,N_13165,N_14317);
and U16613 (N_16613,N_15781,N_14858);
and U16614 (N_16614,N_12045,N_15477);
or U16615 (N_16615,N_14086,N_12288);
nand U16616 (N_16616,N_12364,N_15846);
nor U16617 (N_16617,N_13604,N_14897);
or U16618 (N_16618,N_14932,N_12974);
and U16619 (N_16619,N_14307,N_14638);
nand U16620 (N_16620,N_15378,N_15908);
xor U16621 (N_16621,N_13531,N_12087);
and U16622 (N_16622,N_14435,N_14505);
and U16623 (N_16623,N_12389,N_13286);
nand U16624 (N_16624,N_15772,N_14028);
and U16625 (N_16625,N_14678,N_13509);
or U16626 (N_16626,N_15460,N_15239);
nor U16627 (N_16627,N_14693,N_15508);
or U16628 (N_16628,N_15596,N_15046);
and U16629 (N_16629,N_14018,N_13123);
xor U16630 (N_16630,N_12349,N_14593);
nand U16631 (N_16631,N_14184,N_14141);
or U16632 (N_16632,N_12766,N_14881);
and U16633 (N_16633,N_15485,N_13036);
xnor U16634 (N_16634,N_13066,N_12708);
nand U16635 (N_16635,N_12237,N_12918);
nor U16636 (N_16636,N_14707,N_15360);
nor U16637 (N_16637,N_15511,N_12495);
and U16638 (N_16638,N_15445,N_12286);
and U16639 (N_16639,N_14943,N_12042);
nand U16640 (N_16640,N_14459,N_15550);
or U16641 (N_16641,N_13731,N_14421);
or U16642 (N_16642,N_12712,N_12211);
and U16643 (N_16643,N_13439,N_13427);
and U16644 (N_16644,N_14931,N_13265);
xor U16645 (N_16645,N_12243,N_12715);
and U16646 (N_16646,N_12845,N_13029);
and U16647 (N_16647,N_13025,N_12273);
xnor U16648 (N_16648,N_13671,N_12240);
xor U16649 (N_16649,N_15579,N_13192);
and U16650 (N_16650,N_15436,N_14519);
or U16651 (N_16651,N_12661,N_14181);
nand U16652 (N_16652,N_12176,N_12887);
nor U16653 (N_16653,N_15672,N_14244);
and U16654 (N_16654,N_13651,N_14026);
nor U16655 (N_16655,N_14903,N_13770);
nor U16656 (N_16656,N_13508,N_13361);
or U16657 (N_16657,N_14991,N_15839);
or U16658 (N_16658,N_13484,N_15893);
and U16659 (N_16659,N_13198,N_13514);
nand U16660 (N_16660,N_14034,N_12476);
and U16661 (N_16661,N_15163,N_12140);
nand U16662 (N_16662,N_14441,N_15289);
or U16663 (N_16663,N_14552,N_15208);
or U16664 (N_16664,N_13801,N_14156);
and U16665 (N_16665,N_14802,N_15754);
and U16666 (N_16666,N_13827,N_15106);
nor U16667 (N_16667,N_15912,N_14548);
and U16668 (N_16668,N_12717,N_13610);
and U16669 (N_16669,N_14810,N_12032);
nor U16670 (N_16670,N_14970,N_15621);
xor U16671 (N_16671,N_15070,N_12552);
xor U16672 (N_16672,N_14655,N_14419);
nand U16673 (N_16673,N_15719,N_14260);
nand U16674 (N_16674,N_12726,N_13639);
xor U16675 (N_16675,N_12467,N_14598);
or U16676 (N_16676,N_13893,N_14434);
or U16677 (N_16677,N_13786,N_13184);
nor U16678 (N_16678,N_12318,N_14909);
nor U16679 (N_16679,N_15061,N_13180);
nor U16680 (N_16680,N_12443,N_14893);
nand U16681 (N_16681,N_14923,N_14001);
nand U16682 (N_16682,N_12309,N_15649);
and U16683 (N_16683,N_14310,N_12068);
nor U16684 (N_16684,N_15546,N_12444);
or U16685 (N_16685,N_12771,N_13842);
nor U16686 (N_16686,N_12992,N_13447);
nor U16687 (N_16687,N_12883,N_15375);
nor U16688 (N_16688,N_14722,N_13212);
nand U16689 (N_16689,N_14877,N_13534);
xnor U16690 (N_16690,N_15851,N_15462);
and U16691 (N_16691,N_15461,N_12680);
and U16692 (N_16692,N_14985,N_13407);
nor U16693 (N_16693,N_15980,N_15703);
nand U16694 (N_16694,N_14277,N_15743);
and U16695 (N_16695,N_12947,N_14219);
xnor U16696 (N_16696,N_14111,N_12438);
nand U16697 (N_16697,N_14391,N_14804);
nor U16698 (N_16698,N_12946,N_13081);
or U16699 (N_16699,N_14847,N_12303);
nand U16700 (N_16700,N_15648,N_13313);
and U16701 (N_16701,N_12981,N_13396);
nand U16702 (N_16702,N_14556,N_15988);
nor U16703 (N_16703,N_15423,N_14495);
and U16704 (N_16704,N_14326,N_12277);
nor U16705 (N_16705,N_15283,N_15255);
and U16706 (N_16706,N_13754,N_15037);
or U16707 (N_16707,N_13397,N_13957);
and U16708 (N_16708,N_13755,N_12936);
nand U16709 (N_16709,N_13213,N_12101);
nor U16710 (N_16710,N_12990,N_13698);
nand U16711 (N_16711,N_13620,N_13355);
nand U16712 (N_16712,N_15522,N_13583);
nor U16713 (N_16713,N_15483,N_13959);
nor U16714 (N_16714,N_15368,N_13366);
nor U16715 (N_16715,N_13843,N_12583);
or U16716 (N_16716,N_15967,N_14869);
or U16717 (N_16717,N_13566,N_13183);
nand U16718 (N_16718,N_15020,N_14189);
nor U16719 (N_16719,N_15430,N_13037);
and U16720 (N_16720,N_12592,N_12995);
and U16721 (N_16721,N_15124,N_15219);
nand U16722 (N_16722,N_12123,N_12481);
nand U16723 (N_16723,N_15932,N_14056);
nand U16724 (N_16724,N_12949,N_12169);
nand U16725 (N_16725,N_15675,N_14986);
or U16726 (N_16726,N_15791,N_12134);
nand U16727 (N_16727,N_13108,N_15609);
xor U16728 (N_16728,N_13189,N_12788);
and U16729 (N_16729,N_13937,N_15780);
and U16730 (N_16730,N_15401,N_12783);
and U16731 (N_16731,N_15034,N_14376);
nor U16732 (N_16732,N_15316,N_15939);
and U16733 (N_16733,N_12556,N_15933);
nor U16734 (N_16734,N_14739,N_12858);
nor U16735 (N_16735,N_15307,N_14127);
and U16736 (N_16736,N_13608,N_12860);
and U16737 (N_16737,N_14728,N_13886);
and U16738 (N_16738,N_13201,N_15187);
nor U16739 (N_16739,N_14590,N_14971);
xor U16740 (N_16740,N_12537,N_15497);
nand U16741 (N_16741,N_13852,N_14748);
nor U16742 (N_16742,N_15778,N_14023);
or U16743 (N_16743,N_12584,N_15547);
nand U16744 (N_16744,N_13406,N_13301);
and U16745 (N_16745,N_15822,N_14701);
nor U16746 (N_16746,N_12619,N_12803);
nor U16747 (N_16747,N_13431,N_15747);
xor U16748 (N_16748,N_14282,N_12358);
and U16749 (N_16749,N_13325,N_15351);
nand U16750 (N_16750,N_15786,N_14462);
nor U16751 (N_16751,N_12563,N_14783);
and U16752 (N_16752,N_14761,N_12836);
and U16753 (N_16753,N_15538,N_14401);
and U16754 (N_16754,N_13477,N_14360);
nor U16755 (N_16755,N_14448,N_13116);
nand U16756 (N_16756,N_15683,N_13763);
nand U16757 (N_16757,N_15345,N_15100);
nor U16758 (N_16758,N_12204,N_15082);
nor U16759 (N_16759,N_15412,N_15090);
or U16760 (N_16760,N_14450,N_15832);
and U16761 (N_16761,N_15680,N_13697);
or U16762 (N_16762,N_12950,N_15733);
or U16763 (N_16763,N_12379,N_13673);
or U16764 (N_16764,N_14565,N_12272);
nand U16765 (N_16765,N_14595,N_13101);
or U16766 (N_16766,N_15557,N_13832);
nand U16767 (N_16767,N_15506,N_14345);
and U16768 (N_16768,N_14455,N_14818);
or U16769 (N_16769,N_14892,N_15300);
and U16770 (N_16770,N_15944,N_12794);
and U16771 (N_16771,N_13296,N_12037);
nand U16772 (N_16772,N_12514,N_14204);
xor U16773 (N_16773,N_12325,N_12852);
nor U16774 (N_16774,N_13972,N_13684);
or U16775 (N_16775,N_12589,N_15418);
or U16776 (N_16776,N_14170,N_12641);
nor U16777 (N_16777,N_12963,N_13653);
or U16778 (N_16778,N_13381,N_14681);
or U16779 (N_16779,N_13717,N_15768);
nor U16780 (N_16780,N_15209,N_12321);
nand U16781 (N_16781,N_15032,N_14630);
xnor U16782 (N_16782,N_15491,N_14864);
or U16783 (N_16783,N_13757,N_12915);
nor U16784 (N_16784,N_15055,N_12988);
and U16785 (N_16785,N_12864,N_13533);
nand U16786 (N_16786,N_14935,N_13041);
nor U16787 (N_16787,N_15770,N_15093);
nor U16788 (N_16788,N_15132,N_12264);
or U16789 (N_16789,N_13912,N_15534);
or U16790 (N_16790,N_15941,N_13704);
or U16791 (N_16791,N_14331,N_13835);
or U16792 (N_16792,N_12733,N_15639);
and U16793 (N_16793,N_13733,N_15329);
nand U16794 (N_16794,N_13259,N_12524);
and U16795 (N_16795,N_14527,N_15015);
nand U16796 (N_16796,N_15959,N_15470);
or U16797 (N_16797,N_12972,N_13252);
nand U16798 (N_16798,N_12039,N_14137);
nand U16799 (N_16799,N_14737,N_12526);
or U16800 (N_16800,N_13746,N_15159);
nand U16801 (N_16801,N_14165,N_15951);
or U16802 (N_16802,N_12088,N_14446);
nand U16803 (N_16803,N_13035,N_14362);
and U16804 (N_16804,N_15364,N_14085);
nor U16805 (N_16805,N_14635,N_12013);
or U16806 (N_16806,N_12871,N_13011);
xnor U16807 (N_16807,N_12640,N_12848);
xor U16808 (N_16808,N_13732,N_15472);
or U16809 (N_16809,N_14574,N_12900);
or U16810 (N_16810,N_14769,N_12878);
and U16811 (N_16811,N_14295,N_14960);
nand U16812 (N_16812,N_14747,N_13700);
nand U16813 (N_16813,N_12490,N_13277);
or U16814 (N_16814,N_12314,N_15367);
or U16815 (N_16815,N_14135,N_15903);
or U16816 (N_16816,N_12511,N_13424);
or U16817 (N_16817,N_14567,N_15396);
nand U16818 (N_16818,N_13414,N_13816);
nor U16819 (N_16819,N_13501,N_14063);
or U16820 (N_16820,N_13134,N_12244);
nand U16821 (N_16821,N_15380,N_13771);
nor U16822 (N_16822,N_14011,N_13350);
and U16823 (N_16823,N_14677,N_15773);
nor U16824 (N_16824,N_15958,N_12833);
nand U16825 (N_16825,N_14397,N_12202);
or U16826 (N_16826,N_12433,N_14174);
nor U16827 (N_16827,N_12531,N_12884);
nor U16828 (N_16828,N_12471,N_13258);
or U16829 (N_16829,N_14857,N_15002);
and U16830 (N_16830,N_12054,N_15819);
or U16831 (N_16831,N_15728,N_14554);
or U16832 (N_16832,N_15335,N_14167);
nor U16833 (N_16833,N_15080,N_15709);
or U16834 (N_16834,N_13197,N_14081);
xnor U16835 (N_16835,N_12030,N_13206);
nand U16836 (N_16836,N_13860,N_14062);
or U16837 (N_16837,N_15820,N_12820);
nor U16838 (N_16838,N_13735,N_14795);
xnor U16839 (N_16839,N_14120,N_14708);
or U16840 (N_16840,N_12867,N_15010);
and U16841 (N_16841,N_15304,N_13471);
or U16842 (N_16842,N_12575,N_13969);
or U16843 (N_16843,N_12121,N_14941);
nand U16844 (N_16844,N_12716,N_12740);
and U16845 (N_16845,N_14286,N_14264);
nor U16846 (N_16846,N_12940,N_13914);
or U16847 (N_16847,N_15931,N_12011);
xnor U16848 (N_16848,N_14066,N_12645);
nor U16849 (N_16849,N_13647,N_12507);
nor U16850 (N_16850,N_12075,N_15862);
and U16851 (N_16851,N_13550,N_14948);
or U16852 (N_16852,N_12454,N_13740);
xor U16853 (N_16853,N_13393,N_12937);
or U16854 (N_16854,N_14271,N_14806);
nand U16855 (N_16855,N_15031,N_12560);
xor U16856 (N_16856,N_15922,N_13042);
nor U16857 (N_16857,N_12714,N_15349);
nor U16858 (N_16858,N_12705,N_12650);
nor U16859 (N_16859,N_15089,N_15890);
xnor U16860 (N_16860,N_12485,N_14146);
and U16861 (N_16861,N_14010,N_14239);
nor U16862 (N_16862,N_14052,N_13998);
and U16863 (N_16863,N_15785,N_14355);
nand U16864 (N_16864,N_14592,N_13224);
nand U16865 (N_16865,N_14400,N_14151);
or U16866 (N_16866,N_13836,N_15757);
and U16867 (N_16867,N_15987,N_12913);
nor U16868 (N_16868,N_14438,N_15017);
nor U16869 (N_16869,N_14694,N_14831);
nand U16870 (N_16870,N_13122,N_13536);
nor U16871 (N_16871,N_13022,N_14946);
nand U16872 (N_16872,N_13941,N_12001);
nor U16873 (N_16873,N_14796,N_14198);
and U16874 (N_16874,N_15821,N_15696);
nor U16875 (N_16875,N_14850,N_14418);
nand U16876 (N_16876,N_14573,N_13305);
or U16877 (N_16877,N_12713,N_12792);
xor U16878 (N_16878,N_15586,N_14880);
xor U16879 (N_16879,N_14660,N_14006);
or U16880 (N_16880,N_12970,N_14007);
nor U16881 (N_16881,N_15033,N_15029);
or U16882 (N_16882,N_12201,N_13512);
nor U16883 (N_16883,N_12897,N_12106);
xor U16884 (N_16884,N_15707,N_12294);
nor U16885 (N_16885,N_13802,N_13024);
or U16886 (N_16886,N_13800,N_13058);
nor U16887 (N_16887,N_12870,N_15288);
nand U16888 (N_16888,N_14596,N_12541);
nand U16889 (N_16889,N_13789,N_12449);
or U16890 (N_16890,N_15383,N_15201);
or U16891 (N_16891,N_13658,N_15882);
nand U16892 (N_16892,N_13160,N_13605);
or U16893 (N_16893,N_13023,N_15850);
or U16894 (N_16894,N_12904,N_15006);
and U16895 (N_16895,N_14208,N_15761);
nand U16896 (N_16896,N_14159,N_12207);
and U16897 (N_16897,N_15787,N_14949);
or U16898 (N_16898,N_14579,N_13582);
or U16899 (N_16899,N_13762,N_14501);
and U16900 (N_16900,N_14017,N_12198);
nor U16901 (N_16901,N_14566,N_12394);
nand U16902 (N_16902,N_14608,N_12676);
and U16903 (N_16903,N_12252,N_13217);
nand U16904 (N_16904,N_14361,N_13341);
xnor U16905 (N_16905,N_15441,N_15228);
nor U16906 (N_16906,N_15357,N_14126);
and U16907 (N_16907,N_13649,N_15650);
nand U16908 (N_16908,N_15841,N_14494);
and U16909 (N_16909,N_15014,N_15438);
nand U16910 (N_16910,N_12590,N_12965);
nor U16911 (N_16911,N_13884,N_15514);
nand U16912 (N_16912,N_13026,N_12926);
nand U16913 (N_16913,N_14249,N_12188);
nand U16914 (N_16914,N_12156,N_14092);
nand U16915 (N_16915,N_14955,N_15469);
or U16916 (N_16916,N_12534,N_14808);
nor U16917 (N_16917,N_13004,N_12765);
nor U16918 (N_16918,N_14504,N_12257);
or U16919 (N_16919,N_14340,N_15235);
and U16920 (N_16920,N_12056,N_14133);
xnor U16921 (N_16921,N_14691,N_12797);
nor U16922 (N_16922,N_12125,N_15078);
or U16923 (N_16923,N_15169,N_14732);
or U16924 (N_16924,N_15732,N_13511);
nor U16925 (N_16925,N_12574,N_14663);
nor U16926 (N_16926,N_15361,N_12128);
nand U16927 (N_16927,N_12007,N_14498);
nand U16928 (N_16928,N_13811,N_15849);
nand U16929 (N_16929,N_12667,N_13668);
or U16930 (N_16930,N_12383,N_14201);
or U16931 (N_16931,N_15164,N_12629);
nand U16932 (N_16932,N_13408,N_15210);
or U16933 (N_16933,N_15101,N_13237);
xor U16934 (N_16934,N_14975,N_14646);
nand U16935 (N_16935,N_12895,N_13476);
nor U16936 (N_16936,N_15385,N_13378);
nor U16937 (N_16937,N_14487,N_12843);
nand U16938 (N_16938,N_15356,N_13175);
nand U16939 (N_16939,N_12085,N_12300);
nor U16940 (N_16940,N_14676,N_13540);
or U16941 (N_16941,N_14221,N_15225);
or U16942 (N_16942,N_14349,N_15314);
xor U16943 (N_16943,N_14532,N_12625);
xor U16944 (N_16944,N_12840,N_14024);
xnor U16945 (N_16945,N_15197,N_15505);
nor U16946 (N_16946,N_14058,N_12677);
nor U16947 (N_16947,N_12666,N_12440);
nor U16948 (N_16948,N_13958,N_14812);
or U16949 (N_16949,N_12809,N_15643);
nand U16950 (N_16950,N_12171,N_15981);
nor U16951 (N_16951,N_15767,N_15909);
nand U16952 (N_16952,N_14599,N_13678);
or U16953 (N_16953,N_12456,N_13567);
and U16954 (N_16954,N_14102,N_13932);
and U16955 (N_16955,N_14414,N_14144);
and U16956 (N_16956,N_13038,N_15206);
nand U16957 (N_16957,N_15961,N_13513);
or U16958 (N_16958,N_12729,N_15894);
xor U16959 (N_16959,N_12984,N_14128);
and U16960 (N_16960,N_13409,N_12416);
or U16961 (N_16961,N_15811,N_12170);
and U16962 (N_16962,N_14974,N_12150);
nand U16963 (N_16963,N_13032,N_14964);
nor U16964 (N_16964,N_14101,N_12172);
and U16965 (N_16965,N_12632,N_13223);
or U16966 (N_16966,N_13726,N_13798);
or U16967 (N_16967,N_12786,N_15623);
nor U16968 (N_16968,N_13939,N_12069);
nand U16969 (N_16969,N_14359,N_12488);
nor U16970 (N_16970,N_13310,N_14616);
xor U16971 (N_16971,N_15306,N_14712);
nand U16972 (N_16972,N_13814,N_14908);
nand U16973 (N_16973,N_13283,N_14669);
nand U16974 (N_16974,N_14104,N_13368);
or U16975 (N_16975,N_13846,N_12814);
nor U16976 (N_16976,N_13030,N_13954);
and U16977 (N_16977,N_15929,N_14192);
nor U16978 (N_16978,N_14591,N_12934);
or U16979 (N_16979,N_13473,N_15043);
and U16980 (N_16980,N_14562,N_14456);
or U16981 (N_16981,N_14484,N_12344);
or U16982 (N_16982,N_13797,N_12350);
nor U16983 (N_16983,N_14461,N_12739);
and U16984 (N_16984,N_13450,N_12784);
and U16985 (N_16985,N_15866,N_12828);
nand U16986 (N_16986,N_12579,N_12182);
nand U16987 (N_16987,N_15705,N_12496);
and U16988 (N_16988,N_13267,N_12906);
and U16989 (N_16989,N_13193,N_14833);
and U16990 (N_16990,N_15617,N_13741);
and U16991 (N_16991,N_12971,N_12960);
nand U16992 (N_16992,N_12469,N_13942);
xnor U16993 (N_16993,N_13479,N_12185);
or U16994 (N_16994,N_12225,N_14041);
xor U16995 (N_16995,N_12343,N_13289);
nor U16996 (N_16996,N_12701,N_12097);
and U16997 (N_16997,N_12447,N_14763);
xor U16998 (N_16998,N_15588,N_12461);
or U16999 (N_16999,N_13990,N_13602);
and U17000 (N_17000,N_13597,N_13844);
or U17001 (N_17001,N_13033,N_13850);
nor U17002 (N_17002,N_12028,N_14205);
or U17003 (N_17003,N_15194,N_12908);
nand U17004 (N_17004,N_15622,N_13854);
or U17005 (N_17005,N_15086,N_13337);
nor U17006 (N_17006,N_12613,N_14364);
nand U17007 (N_17007,N_12381,N_14392);
or U17008 (N_17008,N_15456,N_13686);
and U17009 (N_17009,N_13480,N_12697);
xnor U17010 (N_17010,N_15473,N_13344);
and U17011 (N_17011,N_12872,N_14103);
nor U17012 (N_17012,N_13946,N_13069);
nor U17013 (N_17013,N_14938,N_15182);
nand U17014 (N_17014,N_12103,N_14246);
and U17015 (N_17015,N_14265,N_14981);
and U17016 (N_17016,N_14285,N_15576);
or U17017 (N_17017,N_13621,N_13280);
xor U17018 (N_17018,N_13781,N_15173);
nand U17019 (N_17019,N_15657,N_12478);
and U17020 (N_17020,N_15937,N_13288);
nand U17021 (N_17021,N_14328,N_15212);
or U17022 (N_17022,N_13504,N_13716);
or U17023 (N_17023,N_12282,N_12781);
or U17024 (N_17024,N_15128,N_15161);
xor U17025 (N_17025,N_12746,N_14968);
nor U17026 (N_17026,N_15975,N_13488);
nand U17027 (N_17027,N_15278,N_13112);
nor U17028 (N_17028,N_15346,N_13618);
or U17029 (N_17029,N_12637,N_12043);
xor U17030 (N_17030,N_12340,N_15400);
nor U17031 (N_17031,N_14197,N_14617);
and U17032 (N_17032,N_13565,N_14125);
nor U17033 (N_17033,N_14882,N_14848);
or U17034 (N_17034,N_12595,N_14115);
nor U17035 (N_17035,N_12412,N_15665);
nor U17036 (N_17036,N_14304,N_12805);
or U17037 (N_17037,N_12437,N_14768);
nor U17038 (N_17038,N_12486,N_12600);
or U17039 (N_17039,N_15437,N_15280);
and U17040 (N_17040,N_12290,N_14684);
or U17041 (N_17041,N_13169,N_13433);
and U17042 (N_17042,N_12811,N_15455);
nand U17043 (N_17043,N_13744,N_13400);
nand U17044 (N_17044,N_13694,N_14351);
nand U17045 (N_17045,N_12633,N_15798);
and U17046 (N_17046,N_13839,N_14262);
nand U17047 (N_17047,N_15807,N_12004);
nor U17048 (N_17048,N_12033,N_12618);
or U17049 (N_17049,N_14902,N_12741);
xor U17050 (N_17050,N_15150,N_13019);
nand U17051 (N_17051,N_12854,N_15181);
nor U17052 (N_17052,N_15925,N_15405);
xnor U17053 (N_17053,N_15138,N_13306);
and U17054 (N_17054,N_12391,N_14534);
or U17055 (N_17055,N_15671,N_15443);
nor U17056 (N_17056,N_15354,N_13609);
xnor U17057 (N_17057,N_13021,N_15883);
and U17058 (N_17058,N_14726,N_12682);
and U17059 (N_17059,N_15542,N_14147);
nor U17060 (N_17060,N_15956,N_12305);
xnor U17061 (N_17061,N_12544,N_15607);
nand U17062 (N_17062,N_13449,N_13706);
nor U17063 (N_17063,N_13158,N_13248);
nand U17064 (N_17064,N_14413,N_15726);
or U17065 (N_17065,N_13707,N_13445);
xor U17066 (N_17066,N_14196,N_14325);
nor U17067 (N_17067,N_13667,N_14607);
and U17068 (N_17068,N_14142,N_15416);
and U17069 (N_17069,N_15738,N_15718);
nand U17070 (N_17070,N_12826,N_12608);
nand U17071 (N_17071,N_12276,N_13626);
or U17072 (N_17072,N_14689,N_12212);
nand U17073 (N_17073,N_12405,N_13719);
nand U17074 (N_17074,N_13727,N_13094);
nand U17075 (N_17075,N_12299,N_13606);
nand U17076 (N_17076,N_12432,N_15162);
nor U17077 (N_17077,N_14333,N_12408);
or U17078 (N_17078,N_12779,N_14589);
and U17079 (N_17079,N_15995,N_13773);
nor U17080 (N_17080,N_13587,N_13532);
nand U17081 (N_17081,N_15938,N_12297);
nor U17082 (N_17082,N_15190,N_12181);
and U17083 (N_17083,N_13210,N_15974);
nand U17084 (N_17084,N_13453,N_15814);
and U17085 (N_17085,N_15558,N_14703);
nor U17086 (N_17086,N_13956,N_15240);
nand U17087 (N_17087,N_13918,N_15910);
and U17088 (N_17088,N_13752,N_12015);
nor U17089 (N_17089,N_15673,N_12249);
nand U17090 (N_17090,N_13824,N_15286);
or U17091 (N_17091,N_15467,N_14238);
nor U17092 (N_17092,N_15259,N_14904);
or U17093 (N_17093,N_13156,N_15678);
xor U17094 (N_17094,N_13150,N_15524);
or U17095 (N_17095,N_12772,N_12053);
xor U17096 (N_17096,N_15858,N_13973);
or U17097 (N_17097,N_13938,N_14632);
xor U17098 (N_17098,N_12853,N_12603);
nand U17099 (N_17099,N_14718,N_12646);
and U17100 (N_17100,N_12161,N_15263);
or U17101 (N_17101,N_13144,N_13027);
nor U17102 (N_17102,N_13087,N_12361);
nor U17103 (N_17103,N_13166,N_15337);
and U17104 (N_17104,N_12475,N_15353);
and U17105 (N_17105,N_12734,N_15021);
and U17106 (N_17106,N_13869,N_14131);
or U17107 (N_17107,N_12113,N_13823);
nor U17108 (N_17108,N_12678,N_14322);
nor U17109 (N_17109,N_14014,N_13818);
and U17110 (N_17110,N_15797,N_13092);
nor U17111 (N_17111,N_14805,N_15695);
and U17112 (N_17112,N_14779,N_15392);
nor U17113 (N_17113,N_12597,N_13102);
nand U17114 (N_17114,N_14068,N_15826);
and U17115 (N_17115,N_12422,N_14809);
nor U17116 (N_17116,N_12174,N_15426);
or U17117 (N_17117,N_14651,N_15681);
and U17118 (N_17118,N_15007,N_12468);
nor U17119 (N_17119,N_12525,N_12356);
xnor U17120 (N_17120,N_15644,N_13867);
nand U17121 (N_17121,N_13593,N_12256);
or U17122 (N_17122,N_12065,N_12874);
or U17123 (N_17123,N_12492,N_15192);
nand U17124 (N_17124,N_13235,N_12642);
nand U17125 (N_17125,N_15549,N_13916);
nor U17126 (N_17126,N_12656,N_13595);
or U17127 (N_17127,N_12769,N_15953);
xnor U17128 (N_17128,N_15667,N_14046);
and U17129 (N_17129,N_12419,N_14299);
xor U17130 (N_17130,N_13642,N_14194);
and U17131 (N_17131,N_13930,N_13451);
or U17132 (N_17132,N_14749,N_15434);
and U17133 (N_17133,N_15076,N_12126);
xnor U17134 (N_17134,N_15852,N_15911);
nor U17135 (N_17135,N_15444,N_12076);
nand U17136 (N_17136,N_12916,N_15563);
nor U17137 (N_17137,N_12921,N_12819);
xnor U17138 (N_17138,N_13145,N_12755);
or U17139 (N_17139,N_14065,N_15026);
nand U17140 (N_17140,N_13612,N_15094);
nor U17141 (N_17141,N_15790,N_13728);
and U17142 (N_17142,N_12319,N_13863);
or U17143 (N_17143,N_14276,N_15815);
or U17144 (N_17144,N_15996,N_14705);
nand U17145 (N_17145,N_13619,N_14227);
nand U17146 (N_17146,N_15168,N_14305);
or U17147 (N_17147,N_14236,N_12593);
nor U17148 (N_17148,N_12758,N_13768);
nand U17149 (N_17149,N_15736,N_15363);
and U17150 (N_17150,N_14138,N_13928);
and U17151 (N_17151,N_13229,N_13190);
nand U17152 (N_17152,N_14814,N_14190);
nor U17153 (N_17153,N_14040,N_15205);
nand U17154 (N_17154,N_13596,N_14199);
nand U17155 (N_17155,N_12165,N_12052);
xor U17156 (N_17156,N_12548,N_12084);
nor U17157 (N_17157,N_13592,N_15917);
or U17158 (N_17158,N_13114,N_15410);
xnor U17159 (N_17159,N_14817,N_12945);
nand U17160 (N_17160,N_13117,N_12539);
nor U17161 (N_17161,N_14699,N_14633);
nand U17162 (N_17162,N_14875,N_13692);
and U17163 (N_17163,N_13663,N_12429);
and U17164 (N_17164,N_13568,N_14076);
or U17165 (N_17165,N_12226,N_13063);
xnor U17166 (N_17166,N_14667,N_14645);
and U17167 (N_17167,N_13953,N_15552);
xor U17168 (N_17168,N_14329,N_14871);
and U17169 (N_17169,N_13554,N_14217);
nand U17170 (N_17170,N_12060,N_13008);
nand U17171 (N_17171,N_12105,N_14934);
nor U17172 (N_17172,N_14583,N_12731);
nor U17173 (N_17173,N_13009,N_13147);
or U17174 (N_17174,N_12086,N_14570);
nor U17175 (N_17175,N_14835,N_13250);
nand U17176 (N_17176,N_14730,N_15260);
nand U17177 (N_17177,N_12865,N_13390);
nand U17178 (N_17178,N_13730,N_14776);
and U17179 (N_17179,N_14402,N_13047);
xor U17180 (N_17180,N_14177,N_15764);
or U17181 (N_17181,N_12890,N_15966);
or U17182 (N_17182,N_13001,N_12528);
nor U17183 (N_17183,N_14098,N_13055);
nand U17184 (N_17184,N_13984,N_13645);
nor U17185 (N_17185,N_14613,N_13096);
or U17186 (N_17186,N_15388,N_12210);
nor U17187 (N_17187,N_15794,N_13199);
or U17188 (N_17188,N_14954,N_13333);
or U17189 (N_17189,N_13272,N_15536);
and U17190 (N_17190,N_14821,N_15818);
nand U17191 (N_17191,N_14148,N_15174);
nand U17192 (N_17192,N_13693,N_13780);
or U17193 (N_17193,N_13486,N_13578);
nand U17194 (N_17194,N_13881,N_14634);
nor U17195 (N_17195,N_15044,N_13360);
nor U17196 (N_17196,N_14368,N_15669);
and U17197 (N_17197,N_12127,N_15313);
nor U17198 (N_17198,N_14729,N_15012);
nand U17199 (N_17199,N_15468,N_15195);
nor U17200 (N_17200,N_13251,N_14451);
and U17201 (N_17201,N_14856,N_14547);
and U17202 (N_17202,N_15799,N_14200);
or U17203 (N_17203,N_13268,N_13902);
and U17204 (N_17204,N_13128,N_15763);
nor U17205 (N_17205,N_12693,N_15548);
or U17206 (N_17206,N_12217,N_15608);
or U17207 (N_17207,N_14597,N_13100);
or U17208 (N_17208,N_12153,N_12029);
or U17209 (N_17209,N_13625,N_15062);
or U17210 (N_17210,N_12241,N_15999);
nor U17211 (N_17211,N_13091,N_15299);
and U17212 (N_17212,N_15723,N_15528);
xnor U17213 (N_17213,N_15271,N_12576);
and U17214 (N_17214,N_14256,N_13136);
or U17215 (N_17215,N_14278,N_15739);
or U17216 (N_17216,N_12730,N_14762);
and U17217 (N_17217,N_13919,N_15878);
nand U17218 (N_17218,N_12230,N_12424);
nor U17219 (N_17219,N_15074,N_13925);
or U17220 (N_17220,N_12499,N_14690);
nor U17221 (N_17221,N_15679,N_15918);
nand U17222 (N_17222,N_15276,N_15891);
nor U17223 (N_17223,N_15936,N_14886);
nor U17224 (N_17224,N_12406,N_14936);
or U17225 (N_17225,N_14313,N_12725);
nand U17226 (N_17226,N_13420,N_13661);
xnor U17227 (N_17227,N_14577,N_12061);
nor U17228 (N_17228,N_13054,N_14100);
and U17229 (N_17229,N_12081,N_14925);
and U17230 (N_17230,N_13988,N_14920);
nand U17231 (N_17231,N_14576,N_14088);
nor U17232 (N_17232,N_15533,N_15273);
and U17233 (N_17233,N_12111,N_12862);
and U17234 (N_17234,N_13105,N_12055);
xor U17235 (N_17235,N_12694,N_15411);
and U17236 (N_17236,N_12331,N_14618);
nor U17237 (N_17237,N_14887,N_13182);
and U17238 (N_17238,N_13898,N_15028);
xor U17239 (N_17239,N_14258,N_12529);
nor U17240 (N_17240,N_14582,N_12998);
nand U17241 (N_17241,N_12742,N_12505);
nor U17242 (N_17242,N_15371,N_15875);
and U17243 (N_17243,N_12756,N_15319);
and U17244 (N_17244,N_15584,N_13273);
or U17245 (N_17245,N_12503,N_12058);
xor U17246 (N_17246,N_14202,N_14255);
nand U17247 (N_17247,N_14553,N_13775);
nand U17248 (N_17248,N_14228,N_13095);
or U17249 (N_17249,N_13387,N_12175);
nor U17250 (N_17250,N_14302,N_14341);
or U17251 (N_17251,N_15352,N_12917);
or U17252 (N_17252,N_15188,N_15599);
xnor U17253 (N_17253,N_12521,N_15048);
nand U17254 (N_17254,N_12660,N_13254);
or U17255 (N_17255,N_15342,N_13795);
and U17256 (N_17256,N_14733,N_13917);
or U17257 (N_17257,N_12614,N_12420);
nor U17258 (N_17258,N_14288,N_14213);
and U17259 (N_17259,N_12199,N_14724);
nor U17260 (N_17260,N_14840,N_14374);
nor U17261 (N_17261,N_13120,N_15631);
and U17262 (N_17262,N_13167,N_13403);
and U17263 (N_17263,N_14961,N_12549);
nor U17264 (N_17264,N_12943,N_15148);
or U17265 (N_17265,N_13384,N_15318);
or U17266 (N_17266,N_15527,N_12414);
xnor U17267 (N_17267,N_15264,N_15145);
or U17268 (N_17268,N_12248,N_12035);
or U17269 (N_17269,N_15268,N_14631);
and U17270 (N_17270,N_15427,N_12903);
nor U17271 (N_17271,N_14492,N_12323);
nor U17272 (N_17272,N_12994,N_15305);
and U17273 (N_17273,N_14549,N_13318);
nor U17274 (N_17274,N_12191,N_12038);
or U17275 (N_17275,N_14714,N_14686);
and U17276 (N_17276,N_12441,N_15867);
nand U17277 (N_17277,N_13005,N_12179);
nor U17278 (N_17278,N_12573,N_12987);
nand U17279 (N_17279,N_14022,N_12839);
or U17280 (N_17280,N_14267,N_12585);
nand U17281 (N_17281,N_15107,N_15016);
or U17282 (N_17282,N_15213,N_13635);
or U17283 (N_17283,N_14473,N_12168);
xor U17284 (N_17284,N_12083,N_15290);
or U17285 (N_17285,N_12910,N_13083);
xnor U17286 (N_17286,N_13683,N_13541);
and U17287 (N_17287,N_14517,N_12681);
xnor U17288 (N_17288,N_15137,N_12388);
and U17289 (N_17289,N_15465,N_12498);
nand U17290 (N_17290,N_15518,N_15120);
nor U17291 (N_17291,N_15379,N_12487);
nor U17292 (N_17292,N_14679,N_14242);
nor U17293 (N_17293,N_15611,N_12684);
nor U17294 (N_17294,N_15714,N_13576);
and U17295 (N_17295,N_12951,N_13115);
or U17296 (N_17296,N_13654,N_14297);
nand U17297 (N_17297,N_13246,N_14211);
nand U17298 (N_17298,N_15110,N_12139);
nand U17299 (N_17299,N_13677,N_15482);
nor U17300 (N_17300,N_13590,N_15833);
nand U17301 (N_17301,N_15486,N_15097);
and U17302 (N_17302,N_15765,N_15641);
nand U17303 (N_17303,N_14522,N_13172);
xor U17304 (N_17304,N_12582,N_13573);
and U17305 (N_17305,N_13718,N_15227);
and U17306 (N_17306,N_12236,N_12289);
nor U17307 (N_17307,N_12377,N_15248);
nor U17308 (N_17308,N_13245,N_15092);
or U17309 (N_17309,N_15873,N_13840);
and U17310 (N_17310,N_14347,N_13287);
nor U17311 (N_17311,N_12835,N_12010);
and U17312 (N_17312,N_15602,N_14311);
nor U17313 (N_17313,N_15834,N_14428);
and U17314 (N_17314,N_15633,N_15121);
nor U17315 (N_17315,N_12801,N_15083);
nand U17316 (N_17316,N_12410,N_13137);
nor U17317 (N_17317,N_13460,N_14895);
nand U17318 (N_17318,N_15625,N_12752);
nor U17319 (N_17319,N_12009,N_12112);
nor U17320 (N_17320,N_15712,N_13351);
or U17321 (N_17321,N_13794,N_12754);
or U17322 (N_17322,N_15662,N_13833);
or U17323 (N_17323,N_12335,N_14218);
nor U17324 (N_17324,N_15480,N_14178);
and U17325 (N_17325,N_12823,N_14155);
or U17326 (N_17326,N_15464,N_15390);
nand U17327 (N_17327,N_15119,N_14543);
nor U17328 (N_17328,N_14119,N_13335);
and U17329 (N_17329,N_14709,N_15404);
nand U17330 (N_17330,N_15828,N_12292);
or U17331 (N_17331,N_14706,N_12403);
or U17332 (N_17332,N_13015,N_12671);
nor U17333 (N_17333,N_15407,N_12518);
nand U17334 (N_17334,N_15435,N_15414);
nor U17335 (N_17335,N_14020,N_12311);
and U17336 (N_17336,N_13405,N_15344);
xnor U17337 (N_17337,N_15594,N_13185);
nor U17338 (N_17338,N_13622,N_13413);
nor U17339 (N_17339,N_12116,N_14385);
nand U17340 (N_17340,N_13070,N_14106);
nor U17341 (N_17341,N_13933,N_15684);
xnor U17342 (N_17342,N_15868,N_12577);
and U17343 (N_17343,N_14606,N_15561);
nor U17344 (N_17344,N_12194,N_12711);
nand U17345 (N_17345,N_12596,N_15844);
or U17346 (N_17346,N_14121,N_12973);
nor U17347 (N_17347,N_13177,N_14272);
xor U17348 (N_17348,N_14788,N_15992);
xor U17349 (N_17349,N_15153,N_14386);
nor U17350 (N_17350,N_14912,N_15762);
nand U17351 (N_17351,N_14735,N_13388);
or U17352 (N_17352,N_12516,N_12418);
or U17353 (N_17353,N_14237,N_12959);
nand U17354 (N_17354,N_15417,N_12957);
or U17355 (N_17355,N_14602,N_13584);
nand U17356 (N_17356,N_15311,N_15692);
and U17357 (N_17357,N_12136,N_12662);
nor U17358 (N_17358,N_14425,N_14467);
and U17359 (N_17359,N_13061,N_12635);
and U17360 (N_17360,N_12707,N_12636);
or U17361 (N_17361,N_15949,N_15442);
or U17362 (N_17362,N_12520,N_14540);
or U17363 (N_17363,N_12695,N_15340);
nor U17364 (N_17364,N_12690,N_12359);
or U17365 (N_17365,N_13555,N_13312);
nand U17366 (N_17366,N_13065,N_12914);
nor U17367 (N_17367,N_15151,N_13202);
nand U17368 (N_17368,N_14959,N_12426);
and U17369 (N_17369,N_15229,N_12439);
or U17370 (N_17370,N_14905,N_12026);
nand U17371 (N_17371,N_14502,N_15341);
and U17372 (N_17372,N_15328,N_15393);
nand U17373 (N_17373,N_15827,N_14163);
and U17374 (N_17374,N_12545,N_14619);
or U17375 (N_17375,N_12737,N_15149);
or U17376 (N_17376,N_13523,N_15060);
and U17377 (N_17377,N_15459,N_13291);
or U17378 (N_17378,N_13230,N_13803);
or U17379 (N_17379,N_15760,N_14090);
and U17380 (N_17380,N_12665,N_14370);
and U17381 (N_17381,N_15751,N_15433);
nor U17382 (N_17382,N_12480,N_14666);
and U17383 (N_17383,N_15613,N_15591);
nor U17384 (N_17384,N_14112,N_14216);
and U17385 (N_17385,N_14070,N_14291);
xor U17386 (N_17386,N_14420,N_13714);
or U17387 (N_17387,N_15282,N_14433);
or U17388 (N_17388,N_15699,N_14269);
or U17389 (N_17389,N_13791,N_13125);
and U17390 (N_17390,N_12399,N_12533);
nand U17391 (N_17391,N_15238,N_13444);
and U17392 (N_17392,N_14150,N_13526);
and U17393 (N_17393,N_12578,N_14289);
xnor U17394 (N_17394,N_13068,N_13650);
nor U17395 (N_17395,N_13715,N_13525);
nand U17396 (N_17396,N_14224,N_15499);
or U17397 (N_17397,N_15249,N_14183);
nand U17398 (N_17398,N_12557,N_15860);
nand U17399 (N_17399,N_12527,N_14153);
nor U17400 (N_17400,N_14700,N_12543);
nor U17401 (N_17401,N_12378,N_14876);
or U17402 (N_17402,N_15244,N_12566);
nor U17403 (N_17403,N_15635,N_15825);
nor U17404 (N_17404,N_15653,N_14509);
nor U17405 (N_17405,N_15950,N_13976);
nor U17406 (N_17406,N_12332,N_15450);
and U17407 (N_17407,N_12863,N_15218);
and U17408 (N_17408,N_12435,N_13300);
nor U17409 (N_17409,N_14231,N_15627);
nand U17410 (N_17410,N_12610,N_14079);
xnor U17411 (N_17411,N_13934,N_13314);
xor U17412 (N_17412,N_13527,N_15804);
xnor U17413 (N_17413,N_12077,N_12668);
and U17414 (N_17414,N_12691,N_13905);
nand U17415 (N_17415,N_15457,N_14605);
nand U17416 (N_17416,N_12670,N_15386);
nand U17417 (N_17417,N_14957,N_12622);
or U17418 (N_17418,N_15256,N_13132);
or U17419 (N_17419,N_14781,N_15632);
or U17420 (N_17420,N_12308,N_15626);
nor U17421 (N_17421,N_14746,N_15115);
or U17422 (N_17422,N_15362,N_13336);
nand U17423 (N_17423,N_12082,N_14358);
nor U17424 (N_17424,N_13830,N_15167);
and U17425 (N_17425,N_15066,N_14432);
xnor U17426 (N_17426,N_13428,N_12380);
nor U17427 (N_17427,N_15216,N_12892);
and U17428 (N_17428,N_15258,N_12938);
and U17429 (N_17429,N_13079,N_15494);
nor U17430 (N_17430,N_15687,N_13831);
and U17431 (N_17431,N_12442,N_15068);
or U17432 (N_17432,N_13883,N_13908);
or U17433 (N_17433,N_15564,N_13467);
nor U17434 (N_17434,N_15993,N_14372);
nor U17435 (N_17435,N_13044,N_12192);
nand U17436 (N_17436,N_15756,N_13045);
nor U17437 (N_17437,N_14440,N_12609);
nor U17438 (N_17438,N_14481,N_13412);
nand U17439 (N_17439,N_13599,N_12802);
or U17440 (N_17440,N_13463,N_13469);
and U17441 (N_17441,N_15935,N_13743);
xnor U17442 (N_17442,N_15977,N_14406);
nand U17443 (N_17443,N_14516,N_15108);
and U17444 (N_17444,N_12512,N_14427);
and U17445 (N_17445,N_15366,N_13574);
and U17446 (N_17446,N_13963,N_14301);
and U17447 (N_17447,N_13358,N_15721);
and U17448 (N_17448,N_14369,N_14179);
and U17449 (N_17449,N_12540,N_14832);
nand U17450 (N_17450,N_15466,N_13419);
nand U17451 (N_17451,N_12891,N_12515);
and U17452 (N_17452,N_13829,N_14929);
and U17453 (N_17453,N_14468,N_14683);
xor U17454 (N_17454,N_13558,N_15985);
nor U17455 (N_17455,N_12776,N_14612);
nor U17456 (N_17456,N_15997,N_15702);
xnor U17457 (N_17457,N_13992,N_12627);
and U17458 (N_17458,N_12279,N_15803);
or U17459 (N_17459,N_12018,N_12387);
nand U17460 (N_17460,N_12262,N_15566);
and U17461 (N_17461,N_15395,N_15742);
or U17462 (N_17462,N_15175,N_12232);
or U17463 (N_17463,N_15098,N_15892);
nand U17464 (N_17464,N_15624,N_13644);
or U17465 (N_17465,N_14245,N_13399);
and U17466 (N_17466,N_15166,N_14799);
nor U17467 (N_17467,N_14648,N_14695);
nor U17468 (N_17468,N_12091,N_12606);
nor U17469 (N_17469,N_12685,N_13456);
and U17470 (N_17470,N_12242,N_12876);
or U17471 (N_17471,N_13813,N_12509);
or U17472 (N_17472,N_13858,N_14901);
nor U17473 (N_17473,N_12501,N_15131);
or U17474 (N_17474,N_15943,N_14247);
nor U17475 (N_17475,N_12778,N_15551);
xor U17476 (N_17476,N_14458,N_13983);
nor U17477 (N_17477,N_13205,N_12281);
nor U17478 (N_17478,N_14426,N_14939);
or U17479 (N_17479,N_12138,N_14314);
nor U17480 (N_17480,N_14976,N_15198);
nand U17481 (N_17481,N_13826,N_13785);
nor U17482 (N_17482,N_13871,N_14910);
xor U17483 (N_17483,N_15541,N_14906);
nand U17484 (N_17484,N_15453,N_15448);
nand U17485 (N_17485,N_14073,N_15907);
and U17486 (N_17486,N_12902,N_12978);
or U17487 (N_17487,N_14752,N_12295);
nor U17488 (N_17488,N_15081,N_14335);
nor U17489 (N_17489,N_15575,N_14837);
nor U17490 (N_17490,N_13365,N_14099);
nand U17491 (N_17491,N_14756,N_15501);
or U17492 (N_17492,N_14015,N_13442);
and U17493 (N_17493,N_15284,N_13955);
nor U17494 (N_17494,N_14721,N_12021);
nand U17495 (N_17495,N_13777,N_15946);
and U17496 (N_17496,N_13685,N_14916);
or U17497 (N_17497,N_12365,N_13003);
nor U17498 (N_17498,N_14203,N_13652);
or U17499 (N_17499,N_13437,N_14497);
or U17500 (N_17500,N_12888,N_13076);
xnor U17501 (N_17501,N_15310,N_15295);
nand U17502 (N_17502,N_13877,N_15836);
nor U17503 (N_17503,N_14000,N_13385);
nor U17504 (N_17504,N_14780,N_15397);
and U17505 (N_17505,N_13421,N_15025);
or U17506 (N_17506,N_14173,N_12352);
or U17507 (N_17507,N_14713,N_15330);
and U17508 (N_17508,N_12722,N_14585);
and U17509 (N_17509,N_13552,N_12868);
and U17510 (N_17510,N_13559,N_14715);
nor U17511 (N_17511,N_13320,N_14195);
and U17512 (N_17512,N_15133,N_12639);
nor U17513 (N_17513,N_14094,N_14972);
nor U17514 (N_17514,N_12155,N_15041);
and U17515 (N_17515,N_13874,N_13215);
xnor U17516 (N_17516,N_13944,N_15991);
nor U17517 (N_17517,N_15476,N_12346);
or U17518 (N_17518,N_12386,N_12962);
xor U17519 (N_17519,N_12869,N_13039);
or U17520 (N_17520,N_15864,N_12453);
xnor U17521 (N_17521,N_14483,N_15170);
nor U17522 (N_17522,N_15504,N_14053);
nor U17523 (N_17523,N_13106,N_12975);
nand U17524 (N_17524,N_12658,N_13271);
or U17525 (N_17525,N_15211,N_13343);
xor U17526 (N_17526,N_15969,N_13113);
and U17527 (N_17527,N_15502,N_12611);
and U17528 (N_17528,N_13207,N_14379);
nor U17529 (N_17529,N_12847,N_12702);
nor U17530 (N_17530,N_13638,N_13481);
or U17531 (N_17531,N_12265,N_14140);
nand U17532 (N_17532,N_13986,N_14977);
nand U17533 (N_17533,N_15647,N_13162);
nand U17534 (N_17534,N_15520,N_13779);
and U17535 (N_17535,N_13662,N_12417);
or U17536 (N_17536,N_15574,N_15298);
nor U17537 (N_17537,N_12851,N_12831);
and U17538 (N_17538,N_14344,N_14045);
or U17539 (N_17539,N_14185,N_15130);
nand U17540 (N_17540,N_13742,N_12245);
and U17541 (N_17541,N_14753,N_13496);
or U17542 (N_17542,N_14650,N_14084);
nand U17543 (N_17543,N_12944,N_14992);
and U17544 (N_17544,N_14822,N_15018);
nor U17545 (N_17545,N_14158,N_13043);
nor U17546 (N_17546,N_15382,N_13303);
nand U17547 (N_17547,N_15835,N_14521);
nor U17548 (N_17548,N_12046,N_15848);
and U17549 (N_17549,N_14357,N_12648);
or U17550 (N_17550,N_13338,N_15618);
and U17551 (N_17551,N_14692,N_12829);
nand U17552 (N_17552,N_14096,N_14514);
or U17553 (N_17553,N_14643,N_12757);
nor U17554 (N_17554,N_13923,N_12873);
nand U17555 (N_17555,N_15573,N_12285);
nand U17556 (N_17556,N_13672,N_14252);
xnor U17557 (N_17557,N_13018,N_14412);
nand U17558 (N_17558,N_12152,N_14639);
nand U17559 (N_17559,N_13170,N_12547);
nand U17560 (N_17560,N_12969,N_15854);
or U17561 (N_17561,N_14259,N_14342);
xnor U17562 (N_17562,N_13878,N_14051);
nor U17563 (N_17563,N_14398,N_15715);
nor U17564 (N_17564,N_13888,N_14327);
nand U17565 (N_17565,N_12764,N_12457);
and U17566 (N_17566,N_13103,N_15871);
nand U17567 (N_17567,N_12149,N_13981);
and U17568 (N_17568,N_15779,N_14720);
nor U17569 (N_17569,N_13521,N_12535);
or U17570 (N_17570,N_15087,N_15748);
nor U17571 (N_17571,N_15619,N_14704);
nand U17572 (N_17572,N_13868,N_13528);
nor U17573 (N_17573,N_12473,N_15979);
or U17574 (N_17574,N_14866,N_13082);
and U17575 (N_17575,N_13897,N_15440);
nand U17576 (N_17576,N_13000,N_15913);
nand U17577 (N_17577,N_13935,N_12147);
and U17578 (N_17578,N_13952,N_13149);
xnor U17579 (N_17579,N_13872,N_12838);
xnor U17580 (N_17580,N_12313,N_15889);
and U17581 (N_17581,N_12804,N_14792);
and U17582 (N_17582,N_13322,N_14999);
nand U17583 (N_17583,N_13099,N_15503);
or U17584 (N_17584,N_12787,N_12591);
and U17585 (N_17585,N_12785,N_15496);
nor U17586 (N_17586,N_12692,N_13216);
or U17587 (N_17587,N_13793,N_14531);
and U17588 (N_17588,N_15424,N_12881);
nand U17589 (N_17589,N_14859,N_14767);
nor U17590 (N_17590,N_15200,N_13901);
nor U17591 (N_17591,N_15880,N_15580);
and U17592 (N_17592,N_13516,N_12073);
and U17593 (N_17593,N_13304,N_13585);
and U17594 (N_17594,N_13828,N_15172);
nand U17595 (N_17595,N_15246,N_14030);
nand U17596 (N_17596,N_14422,N_15752);
or U17597 (N_17597,N_14841,N_12931);
or U17598 (N_17598,N_15381,N_13438);
or U17599 (N_17599,N_13815,N_13474);
nand U17600 (N_17600,N_13987,N_14870);
or U17601 (N_17601,N_14588,N_12721);
nand U17602 (N_17602,N_14751,N_12233);
or U17603 (N_17603,N_15415,N_13104);
nor U17604 (N_17604,N_13315,N_13422);
and U17605 (N_17605,N_15266,N_14083);
and U17606 (N_17606,N_12980,N_12187);
or U17607 (N_17607,N_12355,N_15024);
xor U17608 (N_17608,N_14029,N_12727);
or U17609 (N_17609,N_13340,N_13537);
and U17610 (N_17610,N_12337,N_15322);
and U17611 (N_17611,N_12479,N_12796);
and U17612 (N_17612,N_14873,N_14486);
or U17613 (N_17613,N_13703,N_13615);
nand U17614 (N_17614,N_15640,N_14064);
and U17615 (N_17615,N_15171,N_12500);
and U17616 (N_17616,N_14520,N_15921);
or U17617 (N_17617,N_13359,N_14798);
nand U17618 (N_17618,N_15507,N_14918);
and U17619 (N_17619,N_15737,N_14966);
nor U17620 (N_17620,N_14061,N_15144);
or U17621 (N_17621,N_12327,N_15523);
and U17622 (N_17622,N_12090,N_12709);
or U17623 (N_17623,N_13676,N_13572);
nor U17624 (N_17624,N_12158,N_15126);
nand U17625 (N_17625,N_13020,N_13669);
nor U17626 (N_17626,N_13729,N_13721);
nand U17627 (N_17627,N_12184,N_12654);
and U17628 (N_17628,N_14430,N_12976);
xor U17629 (N_17629,N_12673,N_14685);
xnor U17630 (N_17630,N_13498,N_13807);
nor U17631 (N_17631,N_12504,N_15971);
nor U17632 (N_17632,N_12020,N_12206);
nor U17633 (N_17633,N_13234,N_12208);
or U17634 (N_17634,N_15049,N_13270);
xor U17635 (N_17635,N_15004,N_13046);
nand U17636 (N_17636,N_14834,N_14390);
nand U17637 (N_17637,N_12813,N_15237);
and U17638 (N_17638,N_15336,N_14889);
or U17639 (N_17639,N_13275,N_13848);
nand U17640 (N_17640,N_12178,N_12247);
nor U17641 (N_17641,N_14035,N_13222);
nand U17642 (N_17642,N_13129,N_12222);
nor U17643 (N_17643,N_13580,N_13086);
nand U17644 (N_17644,N_15141,N_15123);
xnor U17645 (N_17645,N_14789,N_13257);
or U17646 (N_17646,N_15432,N_12354);
and U17647 (N_17647,N_15515,N_12368);
and U17648 (N_17648,N_14489,N_15746);
xor U17649 (N_17649,N_13906,N_13856);
nor U17650 (N_17650,N_15782,N_15214);
or U17651 (N_17651,N_13737,N_13392);
nor U17652 (N_17652,N_13887,N_12909);
nor U17653 (N_17653,N_15487,N_14429);
nand U17654 (N_17654,N_13209,N_13601);
and U17655 (N_17655,N_14047,N_13402);
and U17656 (N_17656,N_13882,N_14488);
and U17657 (N_17657,N_15792,N_13705);
nor U17658 (N_17658,N_14176,N_12750);
nand U17659 (N_17659,N_12846,N_13370);
and U17660 (N_17660,N_15600,N_14862);
nor U17661 (N_17661,N_13821,N_15685);
and U17662 (N_17662,N_13225,N_15498);
nand U17663 (N_17663,N_14320,N_12246);
and U17664 (N_17664,N_14998,N_13720);
xnor U17665 (N_17665,N_13862,N_13903);
and U17666 (N_17666,N_13980,N_14963);
nor U17667 (N_17667,N_12474,N_15125);
or U17668 (N_17668,N_13997,N_12777);
or U17669 (N_17669,N_13994,N_12782);
xor U17670 (N_17670,N_14851,N_14423);
or U17671 (N_17671,N_12339,N_15333);
nand U17672 (N_17672,N_13975,N_12812);
nor U17673 (N_17673,N_15027,N_15572);
nor U17674 (N_17674,N_15677,N_14122);
nand U17675 (N_17675,N_12141,N_15982);
xor U17676 (N_17676,N_12948,N_13187);
or U17677 (N_17677,N_14874,N_15659);
nand U17678 (N_17678,N_14569,N_14036);
and U17679 (N_17679,N_14571,N_13598);
nand U17680 (N_17680,N_14786,N_14393);
nor U17681 (N_17681,N_12849,N_12070);
or U17682 (N_17682,N_13204,N_14479);
nor U17683 (N_17683,N_13404,N_12672);
nor U17684 (N_17684,N_15722,N_13317);
and U17685 (N_17685,N_15139,N_13064);
or U17686 (N_17686,N_15001,N_12477);
and U17687 (N_17687,N_13334,N_15560);
nor U17688 (N_17688,N_13796,N_13591);
nor U17689 (N_17689,N_14775,N_13806);
nand U17690 (N_17690,N_12330,N_15842);
nand U17691 (N_17691,N_14031,N_13503);
and U17692 (N_17692,N_12100,N_15884);
nor U17693 (N_17693,N_13764,N_15334);
xnor U17694 (N_17694,N_12991,N_14702);
nor U17695 (N_17695,N_13013,N_14772);
or U17696 (N_17696,N_15666,N_12024);
or U17697 (N_17697,N_14785,N_12761);
xnor U17698 (N_17698,N_12022,N_14995);
nor U17699 (N_17699,N_15117,N_12209);
or U17700 (N_17700,N_13179,N_15568);
nor U17701 (N_17701,N_14883,N_14913);
or U17702 (N_17702,N_14057,N_12005);
or U17703 (N_17703,N_13617,N_13285);
nand U17704 (N_17704,N_15634,N_14898);
or U17705 (N_17705,N_14021,N_15731);
nand U17706 (N_17706,N_13075,N_14653);
nand U17707 (N_17707,N_13002,N_14528);
nand U17708 (N_17708,N_13646,N_13119);
xnor U17709 (N_17709,N_14408,N_14220);
or U17710 (N_17710,N_13947,N_12229);
nor U17711 (N_17711,N_13107,N_15968);
or U17712 (N_17712,N_12570,N_14523);
or U17713 (N_17713,N_15303,N_15122);
nor U17714 (N_17714,N_14604,N_13485);
or U17715 (N_17715,N_15578,N_14674);
xor U17716 (N_17716,N_13682,N_12118);
or U17717 (N_17717,N_13098,N_14842);
or U17718 (N_17718,N_13062,N_12807);
nand U17719 (N_17719,N_15365,N_14584);
nor U17720 (N_17720,N_12763,N_14145);
nand U17721 (N_17721,N_12258,N_15934);
and U17722 (N_17722,N_14853,N_13196);
nor U17723 (N_17723,N_14110,N_14575);
nand U17724 (N_17724,N_12513,N_12431);
and U17725 (N_17725,N_13739,N_12251);
nand U17726 (N_17726,N_12218,N_15789);
nor U17727 (N_17727,N_12044,N_14375);
or U17728 (N_17728,N_15152,N_12048);
nand U17729 (N_17729,N_13910,N_12638);
nand U17730 (N_17730,N_14382,N_14561);
and U17731 (N_17731,N_15463,N_12283);
xor U17732 (N_17732,N_13524,N_15243);
or U17733 (N_17733,N_14283,N_14292);
nand U17734 (N_17734,N_14234,N_12748);
nand U17735 (N_17735,N_15888,N_12706);
xnor U17736 (N_17736,N_15321,N_15710);
or U17737 (N_17737,N_12351,N_15749);
nand U17738 (N_17738,N_13362,N_14535);
or U17739 (N_17739,N_12310,N_13665);
or U17740 (N_17740,N_14512,N_14671);
nor U17741 (N_17741,N_12630,N_14290);
and U17742 (N_17742,N_12425,N_12743);
xnor U17743 (N_17743,N_14293,N_15109);
or U17744 (N_17744,N_12253,N_15075);
and U17745 (N_17745,N_14171,N_12859);
and U17746 (N_17746,N_15553,N_15963);
nand U17747 (N_17747,N_12799,N_14659);
or U17748 (N_17748,N_14568,N_13774);
and U17749 (N_17749,N_14894,N_14687);
nor U17750 (N_17750,N_14636,N_13507);
and U17751 (N_17751,N_14537,N_15690);
nor U17752 (N_17752,N_14956,N_13080);
and U17753 (N_17753,N_15051,N_13461);
or U17754 (N_17754,N_12561,N_15489);
nor U17755 (N_17755,N_14824,N_12219);
nor U17756 (N_17756,N_14166,N_15686);
nand U17757 (N_17757,N_12601,N_12532);
or U17758 (N_17758,N_14323,N_14710);
nor U17759 (N_17759,N_13913,N_13146);
and U17760 (N_17760,N_14485,N_12580);
nand U17761 (N_17761,N_13962,N_15301);
and U17762 (N_17762,N_12568,N_13391);
nand U17763 (N_17763,N_13712,N_14654);
or U17764 (N_17764,N_14924,N_14863);
or U17765 (N_17765,N_15881,N_14442);
or U17766 (N_17766,N_14206,N_12428);
or U17767 (N_17767,N_15645,N_12647);
nand U17768 (N_17768,N_14089,N_14482);
nand U17769 (N_17769,N_12855,N_13153);
and U17770 (N_17770,N_14223,N_14942);
xnor U17771 (N_17771,N_15348,N_15583);
and U17772 (N_17772,N_14215,N_12749);
nand U17773 (N_17773,N_13293,N_12586);
and U17774 (N_17774,N_13812,N_15253);
and U17775 (N_17775,N_12448,N_12555);
or U17776 (N_17776,N_12008,N_13920);
and U17777 (N_17777,N_14080,N_13127);
or U17778 (N_17778,N_13766,N_13864);
or U17779 (N_17779,N_13782,N_12110);
xor U17780 (N_17780,N_14740,N_12360);
nand U17781 (N_17781,N_14298,N_13430);
or U17782 (N_17782,N_13347,N_13915);
and U17783 (N_17783,N_12143,N_13389);
nor U17784 (N_17784,N_12395,N_12621);
and U17785 (N_17785,N_15116,N_13611);
or U17786 (N_17786,N_12144,N_15419);
nor U17787 (N_17787,N_12163,N_13176);
nand U17788 (N_17788,N_13603,N_15297);
nor U17789 (N_17789,N_15916,N_14186);
or U17790 (N_17790,N_13895,N_12166);
and U17791 (N_17791,N_15409,N_12649);
nor U17792 (N_17792,N_12049,N_12367);
or U17793 (N_17793,N_12195,N_13263);
nand U17794 (N_17794,N_12718,N_15269);
and U17795 (N_17795,N_12462,N_13904);
nand U17796 (N_17796,N_12675,N_14665);
nor U17797 (N_17797,N_12000,N_13088);
and U17798 (N_17798,N_13970,N_13553);
nand U17799 (N_17799,N_12019,N_12375);
or U17800 (N_17800,N_13586,N_14008);
xor U17801 (N_17801,N_13231,N_15102);
nand U17802 (N_17802,N_13164,N_12374);
and U17803 (N_17803,N_13849,N_13459);
nand U17804 (N_17804,N_13154,N_12051);
xor U17805 (N_17805,N_13415,N_14820);
nand U17806 (N_17806,N_13426,N_14005);
nor U17807 (N_17807,N_12301,N_14240);
or U17808 (N_17808,N_12071,N_12284);
nor U17809 (N_17809,N_15431,N_13244);
nand U17810 (N_17810,N_14839,N_13899);
or U17811 (N_17811,N_13760,N_12607);
nor U17812 (N_17812,N_15165,N_13996);
and U17813 (N_17813,N_15023,N_13482);
nand U17814 (N_17814,N_13967,N_13348);
or U17815 (N_17815,N_15544,N_14827);
xor U17816 (N_17816,N_13279,N_14263);
nor U17817 (N_17817,N_14367,N_12753);
and U17818 (N_17818,N_14339,N_15281);
xor U17819 (N_17819,N_12791,N_12928);
nor U17820 (N_17820,N_13155,N_12093);
and U17821 (N_17821,N_14250,N_14990);
nand U17822 (N_17822,N_15447,N_15543);
or U17823 (N_17823,N_14987,N_14640);
nand U17824 (N_17824,N_12423,N_13071);
xnor U17825 (N_17825,N_13885,N_12094);
nand U17826 (N_17826,N_15484,N_15512);
and U17827 (N_17827,N_15808,N_13751);
xnor U17828 (N_17828,N_14363,N_13808);
xor U17829 (N_17829,N_13321,N_13500);
nand U17830 (N_17830,N_15947,N_12837);
nand U17831 (N_17831,N_12768,N_15948);
xor U17832 (N_17832,N_15275,N_15215);
or U17833 (N_17833,N_13142,N_15207);
nand U17834 (N_17834,N_14952,N_12160);
or U17835 (N_17835,N_14637,N_12338);
or U17836 (N_17836,N_12933,N_13853);
or U17837 (N_17837,N_15970,N_13748);
and U17838 (N_17838,N_15458,N_13756);
nand U17839 (N_17839,N_15567,N_13506);
or U17840 (N_17840,N_13949,N_12825);
and U17841 (N_17841,N_12510,N_15030);
nand U17842 (N_17842,N_12830,N_12334);
or U17843 (N_17843,N_12336,N_12316);
nor U17844 (N_17844,N_13670,N_15135);
nand U17845 (N_17845,N_15745,N_15326);
and U17846 (N_17846,N_12653,N_13616);
xnor U17847 (N_17847,N_12489,N_14117);
or U17848 (N_17848,N_15370,N_14388);
nand U17849 (N_17849,N_15914,N_13657);
nor U17850 (N_17850,N_15339,N_12626);
and U17851 (N_17851,N_13483,N_13857);
nand U17852 (N_17852,N_15231,N_15955);
xnor U17853 (N_17853,N_14226,N_12254);
xor U17854 (N_17854,N_13817,N_13238);
nand U17855 (N_17855,N_12074,N_13040);
nand U17856 (N_17856,N_14243,N_13520);
nand U17857 (N_17857,N_12353,N_15226);
and U17858 (N_17858,N_13161,N_15577);
or U17859 (N_17859,N_12402,N_15879);
or U17860 (N_17860,N_12939,N_15490);
and U17861 (N_17861,N_13097,N_12466);
nor U17862 (N_17862,N_13628,N_14266);
or U17863 (N_17863,N_13057,N_15744);
or U17864 (N_17864,N_12270,N_13159);
or U17865 (N_17865,N_14352,N_14447);
nand U17866 (N_17866,N_13778,N_13688);
nor U17867 (N_17867,N_13505,N_14953);
xnor U17868 (N_17868,N_13448,N_15495);
or U17869 (N_17869,N_15876,N_12554);
and U17870 (N_17870,N_15234,N_13349);
nor U17871 (N_17871,N_13724,N_12773);
or U17872 (N_17872,N_13989,N_14983);
or U17873 (N_17873,N_13446,N_13357);
and U17874 (N_17874,N_13909,N_12197);
or U17875 (N_17875,N_12808,N_14766);
nor U17876 (N_17876,N_12594,N_14060);
nand U17877 (N_17877,N_14409,N_14979);
nor U17878 (N_17878,N_12955,N_12818);
nand U17879 (N_17879,N_13247,N_12901);
and U17880 (N_17880,N_14387,N_14134);
and U17881 (N_17881,N_12135,N_14095);
nand U17882 (N_17882,N_14958,N_13845);
nor U17883 (N_17883,N_15990,N_15247);
nor U17884 (N_17884,N_14611,N_14043);
and U17885 (N_17885,N_14334,N_12268);
and U17886 (N_17886,N_12587,N_15986);
nand U17887 (N_17887,N_15500,N_12542);
nor U17888 (N_17888,N_14621,N_14415);
and U17889 (N_17889,N_13292,N_15775);
nor U17890 (N_17890,N_14879,N_14625);
nor U17891 (N_17891,N_14620,N_13641);
nor U17892 (N_17892,N_13232,N_13971);
nand U17893 (N_17893,N_15425,N_15630);
or U17894 (N_17894,N_12952,N_14306);
nor U17895 (N_17895,N_15701,N_13679);
nand U17896 (N_17896,N_13111,N_14622);
nor U17897 (N_17897,N_15475,N_13870);
nand U17898 (N_17898,N_12372,N_13067);
or U17899 (N_17899,N_14319,N_13016);
xor U17900 (N_17900,N_12770,N_12398);
and U17901 (N_17901,N_15179,N_13139);
and U17902 (N_17902,N_13266,N_13345);
nor U17903 (N_17903,N_15035,N_12133);
and U17904 (N_17904,N_14453,N_14016);
nor U17905 (N_17905,N_15428,N_14819);
and U17906 (N_17906,N_14978,N_14108);
nor U17907 (N_17907,N_14233,N_13090);
or U17908 (N_17908,N_15713,N_13200);
nor U17909 (N_17909,N_12132,N_14536);
nor U17910 (N_17910,N_15800,N_13985);
or U17911 (N_17911,N_15292,N_12137);
nor U17912 (N_17912,N_15202,N_12012);
nor U17913 (N_17913,N_12745,N_15072);
and U17914 (N_17914,N_12446,N_13837);
nor U17915 (N_17915,N_15887,N_14465);
and U17916 (N_17916,N_14930,N_14914);
nor U17917 (N_17917,N_13489,N_13927);
or U17918 (N_17918,N_14813,N_13331);
and U17919 (N_17919,N_15452,N_12861);
nand U17920 (N_17920,N_13302,N_13006);
nor U17921 (N_17921,N_12698,N_13841);
nor U17922 (N_17922,N_13702,N_13753);
and U17923 (N_17923,N_13911,N_15824);
and U17924 (N_17924,N_13907,N_13965);
or U17925 (N_17925,N_15930,N_15233);
nor U17926 (N_17926,N_15146,N_15724);
and U17927 (N_17927,N_14962,N_14394);
nor U17928 (N_17928,N_13470,N_15569);
and U17929 (N_17929,N_15942,N_12146);
nand U17930 (N_17930,N_15670,N_13457);
and U17931 (N_17931,N_12615,N_12790);
nand U17932 (N_17932,N_15637,N_13377);
nor U17933 (N_17933,N_14182,N_12459);
nand U17934 (N_17934,N_13411,N_13436);
and U17935 (N_17935,N_14309,N_14510);
nand U17936 (N_17936,N_14557,N_14077);
nand U17937 (N_17937,N_14353,N_14794);
and U17938 (N_17938,N_15011,N_15957);
and U17939 (N_17939,N_14742,N_12109);
or U17940 (N_17940,N_15590,N_15189);
or U17941 (N_17941,N_13879,N_13233);
xor U17942 (N_17942,N_15421,N_15186);
nor U17943 (N_17943,N_15606,N_15118);
nand U17944 (N_17944,N_12841,N_15823);
xor U17945 (N_17945,N_14209,N_14744);
or U17946 (N_17946,N_15526,N_13051);
nor U17947 (N_17947,N_15199,N_12102);
xnor U17948 (N_17948,N_12502,N_12098);
or U17949 (N_17949,N_15906,N_12923);
xnor U17950 (N_17950,N_12942,N_12696);
and U17951 (N_17951,N_14826,N_12806);
or U17952 (N_17952,N_15964,N_13674);
and U17953 (N_17953,N_12688,N_15595);
nor U17954 (N_17954,N_12605,N_15614);
and U17955 (N_17955,N_12404,N_15203);
nor U17956 (N_17956,N_15693,N_12571);
and U17957 (N_17957,N_13141,N_13542);
nor U17958 (N_17958,N_13547,N_15656);
or U17959 (N_17959,N_12215,N_14087);
nand U17960 (N_17960,N_15597,N_15924);
and U17961 (N_17961,N_15872,N_13991);
and U17962 (N_17962,N_14784,N_14967);
or U17963 (N_17963,N_13493,N_15183);
and U17964 (N_17964,N_12347,N_14287);
nor U17965 (N_17965,N_15230,N_15729);
xnor U17966 (N_17966,N_14500,N_13188);
nand U17967 (N_17967,N_12173,N_12780);
nor U17968 (N_17968,N_12723,N_14773);
xnor U17969 (N_17969,N_13425,N_15689);
and U17970 (N_17970,N_14675,N_15952);
or U17971 (N_17971,N_13007,N_15257);
and U17972 (N_17972,N_12567,N_15327);
nor U17973 (N_17973,N_14300,N_14383);
xnor U17974 (N_17974,N_13260,N_12002);
nor U17975 (N_17975,N_14815,N_15112);
and U17976 (N_17976,N_13924,N_15535);
nand U17977 (N_17977,N_13680,N_14072);
nand U17978 (N_17978,N_14907,N_14389);
or U17979 (N_17979,N_13255,N_12844);
or U17980 (N_17980,N_13600,N_14222);
xor U17981 (N_17981,N_14823,N_12924);
and U17982 (N_17982,N_13052,N_12274);
nand U17983 (N_17983,N_12720,N_14091);
nand U17984 (N_17984,N_14852,N_13376);
nor U17985 (N_17985,N_14443,N_13922);
nand U17986 (N_17986,N_14003,N_12824);
or U17987 (N_17987,N_12315,N_14727);
nor U17988 (N_17988,N_15795,N_12328);
xor U17989 (N_17989,N_15940,N_13072);
or U17990 (N_17990,N_13328,N_15241);
nor U17991 (N_17991,N_12203,N_12278);
nor U17992 (N_17992,N_15628,N_14891);
nor U17993 (N_17993,N_14478,N_14586);
or U17994 (N_17994,N_15593,N_15403);
or U17995 (N_17995,N_13738,N_14042);
and U17996 (N_17996,N_12329,N_15783);
and U17997 (N_17997,N_15646,N_12643);
nand U17998 (N_17998,N_15727,N_13876);
nand U17999 (N_17999,N_12451,N_13131);
or U18000 (N_18000,N_12822,N_14630);
xor U18001 (N_18001,N_15403,N_15913);
nor U18002 (N_18002,N_13939,N_12225);
nand U18003 (N_18003,N_12548,N_14471);
nand U18004 (N_18004,N_14914,N_12601);
xor U18005 (N_18005,N_14305,N_13382);
nor U18006 (N_18006,N_15919,N_12989);
and U18007 (N_18007,N_13535,N_15578);
xnor U18008 (N_18008,N_15347,N_12010);
or U18009 (N_18009,N_14758,N_14278);
or U18010 (N_18010,N_15185,N_13509);
nand U18011 (N_18011,N_13765,N_13584);
and U18012 (N_18012,N_12640,N_12857);
or U18013 (N_18013,N_14794,N_15410);
xnor U18014 (N_18014,N_13848,N_12206);
or U18015 (N_18015,N_15157,N_13339);
and U18016 (N_18016,N_14427,N_12526);
and U18017 (N_18017,N_12555,N_13740);
or U18018 (N_18018,N_15797,N_12973);
and U18019 (N_18019,N_13609,N_15949);
nor U18020 (N_18020,N_15824,N_13927);
and U18021 (N_18021,N_12100,N_15217);
nand U18022 (N_18022,N_12148,N_15036);
nor U18023 (N_18023,N_14997,N_15904);
nand U18024 (N_18024,N_13507,N_14009);
and U18025 (N_18025,N_12522,N_13741);
xor U18026 (N_18026,N_15782,N_14504);
xnor U18027 (N_18027,N_15759,N_14411);
nor U18028 (N_18028,N_15120,N_14959);
xnor U18029 (N_18029,N_12810,N_12766);
or U18030 (N_18030,N_12211,N_14944);
nor U18031 (N_18031,N_14417,N_13275);
nand U18032 (N_18032,N_15799,N_12611);
nor U18033 (N_18033,N_15324,N_13889);
and U18034 (N_18034,N_14112,N_12822);
and U18035 (N_18035,N_12415,N_14033);
and U18036 (N_18036,N_15776,N_15643);
nand U18037 (N_18037,N_13445,N_12008);
and U18038 (N_18038,N_15019,N_13155);
nand U18039 (N_18039,N_12631,N_14555);
and U18040 (N_18040,N_13860,N_15609);
nor U18041 (N_18041,N_14519,N_14075);
nor U18042 (N_18042,N_15094,N_15704);
nor U18043 (N_18043,N_14514,N_14596);
or U18044 (N_18044,N_12525,N_12138);
or U18045 (N_18045,N_14654,N_15795);
nand U18046 (N_18046,N_13340,N_15097);
and U18047 (N_18047,N_13049,N_13877);
xor U18048 (N_18048,N_15494,N_12947);
and U18049 (N_18049,N_15755,N_13565);
nand U18050 (N_18050,N_14050,N_15119);
nand U18051 (N_18051,N_15549,N_14692);
or U18052 (N_18052,N_12042,N_13506);
nor U18053 (N_18053,N_12853,N_15854);
or U18054 (N_18054,N_15803,N_14919);
or U18055 (N_18055,N_15419,N_13746);
or U18056 (N_18056,N_15728,N_15289);
or U18057 (N_18057,N_12108,N_12175);
nor U18058 (N_18058,N_15132,N_15131);
or U18059 (N_18059,N_13340,N_12832);
or U18060 (N_18060,N_13846,N_15145);
xor U18061 (N_18061,N_15054,N_14878);
nor U18062 (N_18062,N_14689,N_13499);
xor U18063 (N_18063,N_15608,N_15194);
nand U18064 (N_18064,N_14604,N_12675);
nor U18065 (N_18065,N_15750,N_15424);
and U18066 (N_18066,N_12595,N_13988);
or U18067 (N_18067,N_15685,N_13276);
nand U18068 (N_18068,N_15961,N_13161);
nor U18069 (N_18069,N_13754,N_15862);
and U18070 (N_18070,N_13301,N_13207);
nor U18071 (N_18071,N_15086,N_12137);
nand U18072 (N_18072,N_14846,N_14973);
nand U18073 (N_18073,N_13121,N_15821);
nor U18074 (N_18074,N_14518,N_13453);
or U18075 (N_18075,N_12560,N_12052);
xor U18076 (N_18076,N_15849,N_13643);
nand U18077 (N_18077,N_15153,N_12574);
nand U18078 (N_18078,N_13047,N_13413);
nor U18079 (N_18079,N_15930,N_12560);
or U18080 (N_18080,N_15736,N_13110);
nor U18081 (N_18081,N_14336,N_14373);
xor U18082 (N_18082,N_13616,N_15538);
nand U18083 (N_18083,N_15377,N_12180);
and U18084 (N_18084,N_14898,N_14454);
nand U18085 (N_18085,N_13490,N_12987);
and U18086 (N_18086,N_12981,N_13213);
and U18087 (N_18087,N_14079,N_15951);
or U18088 (N_18088,N_14499,N_12122);
nor U18089 (N_18089,N_13065,N_12079);
nor U18090 (N_18090,N_15836,N_14303);
nor U18091 (N_18091,N_14458,N_14248);
nand U18092 (N_18092,N_12178,N_12411);
nor U18093 (N_18093,N_13795,N_15637);
nand U18094 (N_18094,N_13119,N_12897);
nor U18095 (N_18095,N_15468,N_13515);
nand U18096 (N_18096,N_15180,N_13956);
nand U18097 (N_18097,N_13449,N_14380);
or U18098 (N_18098,N_13434,N_13184);
and U18099 (N_18099,N_13427,N_12977);
nor U18100 (N_18100,N_13317,N_14858);
nand U18101 (N_18101,N_15429,N_13418);
or U18102 (N_18102,N_13389,N_14632);
nor U18103 (N_18103,N_15646,N_13759);
and U18104 (N_18104,N_13950,N_15143);
nand U18105 (N_18105,N_15957,N_13414);
xnor U18106 (N_18106,N_14837,N_13243);
or U18107 (N_18107,N_15017,N_13332);
and U18108 (N_18108,N_12166,N_15149);
nor U18109 (N_18109,N_15234,N_15843);
nor U18110 (N_18110,N_13090,N_13336);
nand U18111 (N_18111,N_12504,N_12832);
xor U18112 (N_18112,N_13419,N_13682);
and U18113 (N_18113,N_15424,N_13155);
or U18114 (N_18114,N_14962,N_15081);
or U18115 (N_18115,N_13610,N_12251);
and U18116 (N_18116,N_13891,N_12391);
xnor U18117 (N_18117,N_15015,N_15149);
nand U18118 (N_18118,N_15697,N_15982);
nand U18119 (N_18119,N_15853,N_12382);
nor U18120 (N_18120,N_13775,N_14419);
nand U18121 (N_18121,N_14173,N_12594);
nor U18122 (N_18122,N_15506,N_12470);
and U18123 (N_18123,N_12290,N_12726);
nand U18124 (N_18124,N_12649,N_15927);
or U18125 (N_18125,N_13782,N_15128);
or U18126 (N_18126,N_15632,N_15370);
xnor U18127 (N_18127,N_12717,N_14304);
or U18128 (N_18128,N_13678,N_15415);
or U18129 (N_18129,N_12115,N_13095);
or U18130 (N_18130,N_13035,N_14518);
and U18131 (N_18131,N_13857,N_13420);
nor U18132 (N_18132,N_14317,N_14827);
nor U18133 (N_18133,N_14200,N_13872);
nor U18134 (N_18134,N_15967,N_12225);
nand U18135 (N_18135,N_14775,N_14603);
nand U18136 (N_18136,N_13112,N_13535);
nand U18137 (N_18137,N_12188,N_15373);
or U18138 (N_18138,N_15201,N_13996);
or U18139 (N_18139,N_14728,N_12182);
xnor U18140 (N_18140,N_15464,N_12385);
or U18141 (N_18141,N_15348,N_13862);
nand U18142 (N_18142,N_13781,N_12118);
nand U18143 (N_18143,N_14708,N_14724);
xnor U18144 (N_18144,N_15812,N_13898);
nand U18145 (N_18145,N_14504,N_13202);
nor U18146 (N_18146,N_14416,N_14386);
or U18147 (N_18147,N_13397,N_12448);
nor U18148 (N_18148,N_12574,N_12076);
and U18149 (N_18149,N_15833,N_14939);
and U18150 (N_18150,N_13899,N_15426);
or U18151 (N_18151,N_12278,N_14970);
or U18152 (N_18152,N_15634,N_14153);
nand U18153 (N_18153,N_13331,N_12490);
and U18154 (N_18154,N_13931,N_12274);
nor U18155 (N_18155,N_14557,N_14272);
and U18156 (N_18156,N_15831,N_15319);
nor U18157 (N_18157,N_12910,N_14860);
nand U18158 (N_18158,N_14690,N_14401);
nand U18159 (N_18159,N_12416,N_14662);
or U18160 (N_18160,N_14365,N_13637);
nor U18161 (N_18161,N_12961,N_12205);
nand U18162 (N_18162,N_12456,N_15006);
or U18163 (N_18163,N_12728,N_14768);
nand U18164 (N_18164,N_15740,N_15794);
nand U18165 (N_18165,N_13872,N_12860);
or U18166 (N_18166,N_15818,N_12299);
or U18167 (N_18167,N_12205,N_15128);
or U18168 (N_18168,N_13248,N_12212);
nand U18169 (N_18169,N_14517,N_13625);
and U18170 (N_18170,N_15246,N_15659);
nor U18171 (N_18171,N_14001,N_14021);
and U18172 (N_18172,N_12759,N_12355);
nand U18173 (N_18173,N_13661,N_12985);
xnor U18174 (N_18174,N_12139,N_15166);
and U18175 (N_18175,N_14159,N_13647);
nor U18176 (N_18176,N_13181,N_13257);
or U18177 (N_18177,N_12255,N_15609);
nand U18178 (N_18178,N_13808,N_13059);
nand U18179 (N_18179,N_15197,N_15034);
nand U18180 (N_18180,N_14590,N_14895);
or U18181 (N_18181,N_14061,N_12446);
xor U18182 (N_18182,N_14934,N_12781);
and U18183 (N_18183,N_14313,N_12983);
nand U18184 (N_18184,N_13355,N_12135);
nand U18185 (N_18185,N_14484,N_12828);
and U18186 (N_18186,N_15639,N_15591);
or U18187 (N_18187,N_15018,N_14637);
nor U18188 (N_18188,N_13283,N_13970);
nor U18189 (N_18189,N_15626,N_15443);
and U18190 (N_18190,N_14762,N_13668);
nor U18191 (N_18191,N_13858,N_14334);
or U18192 (N_18192,N_15232,N_13206);
and U18193 (N_18193,N_12954,N_13565);
or U18194 (N_18194,N_15476,N_15963);
or U18195 (N_18195,N_15570,N_14772);
nand U18196 (N_18196,N_14089,N_15072);
and U18197 (N_18197,N_13276,N_13521);
nand U18198 (N_18198,N_15862,N_13083);
nor U18199 (N_18199,N_14560,N_14937);
nor U18200 (N_18200,N_14491,N_14714);
nand U18201 (N_18201,N_13539,N_15693);
nand U18202 (N_18202,N_14748,N_14567);
or U18203 (N_18203,N_15322,N_13131);
nand U18204 (N_18204,N_14242,N_12866);
or U18205 (N_18205,N_13261,N_15478);
and U18206 (N_18206,N_14244,N_13767);
and U18207 (N_18207,N_13501,N_12302);
and U18208 (N_18208,N_12071,N_12478);
or U18209 (N_18209,N_12816,N_12790);
nand U18210 (N_18210,N_15074,N_13843);
nor U18211 (N_18211,N_14836,N_15986);
and U18212 (N_18212,N_15724,N_13550);
and U18213 (N_18213,N_15776,N_13603);
nand U18214 (N_18214,N_12758,N_15066);
nand U18215 (N_18215,N_15655,N_14520);
or U18216 (N_18216,N_12155,N_12908);
and U18217 (N_18217,N_12178,N_12772);
nand U18218 (N_18218,N_15027,N_12811);
nor U18219 (N_18219,N_15964,N_12780);
or U18220 (N_18220,N_12300,N_14963);
nand U18221 (N_18221,N_15634,N_14981);
nor U18222 (N_18222,N_12998,N_14366);
and U18223 (N_18223,N_12686,N_14478);
nor U18224 (N_18224,N_13238,N_12856);
nand U18225 (N_18225,N_14235,N_15121);
and U18226 (N_18226,N_12549,N_15354);
nor U18227 (N_18227,N_15815,N_15910);
nor U18228 (N_18228,N_13920,N_15203);
or U18229 (N_18229,N_14479,N_13600);
nand U18230 (N_18230,N_15191,N_12214);
nand U18231 (N_18231,N_14968,N_12393);
or U18232 (N_18232,N_12380,N_13816);
nand U18233 (N_18233,N_12642,N_14389);
nand U18234 (N_18234,N_12118,N_14935);
nand U18235 (N_18235,N_14834,N_12165);
nor U18236 (N_18236,N_13823,N_13293);
and U18237 (N_18237,N_13251,N_12687);
or U18238 (N_18238,N_12749,N_14550);
nand U18239 (N_18239,N_12002,N_15550);
nor U18240 (N_18240,N_14088,N_13521);
or U18241 (N_18241,N_12379,N_12102);
xnor U18242 (N_18242,N_12351,N_12499);
and U18243 (N_18243,N_13432,N_14678);
and U18244 (N_18244,N_14203,N_15076);
nor U18245 (N_18245,N_14200,N_12611);
nor U18246 (N_18246,N_15342,N_12434);
nor U18247 (N_18247,N_15970,N_12752);
nor U18248 (N_18248,N_12704,N_13828);
nand U18249 (N_18249,N_12898,N_12985);
or U18250 (N_18250,N_13468,N_12883);
nand U18251 (N_18251,N_15617,N_15782);
and U18252 (N_18252,N_14736,N_13997);
nor U18253 (N_18253,N_14176,N_15496);
nor U18254 (N_18254,N_13242,N_14140);
nor U18255 (N_18255,N_14167,N_15680);
or U18256 (N_18256,N_12579,N_12666);
or U18257 (N_18257,N_13283,N_12074);
nor U18258 (N_18258,N_13218,N_12716);
and U18259 (N_18259,N_14448,N_14421);
xor U18260 (N_18260,N_12127,N_14420);
and U18261 (N_18261,N_12165,N_15033);
nor U18262 (N_18262,N_14948,N_13685);
or U18263 (N_18263,N_13902,N_12689);
and U18264 (N_18264,N_12093,N_13854);
or U18265 (N_18265,N_14613,N_12544);
nor U18266 (N_18266,N_13324,N_14707);
nor U18267 (N_18267,N_14175,N_12783);
nor U18268 (N_18268,N_12617,N_15661);
nand U18269 (N_18269,N_14990,N_14421);
nand U18270 (N_18270,N_15366,N_13294);
nor U18271 (N_18271,N_14539,N_14495);
and U18272 (N_18272,N_13304,N_13973);
xnor U18273 (N_18273,N_14242,N_15262);
nand U18274 (N_18274,N_13296,N_14774);
nor U18275 (N_18275,N_14489,N_12659);
nor U18276 (N_18276,N_14546,N_14094);
or U18277 (N_18277,N_12101,N_14569);
nor U18278 (N_18278,N_13995,N_15053);
nand U18279 (N_18279,N_13143,N_12598);
xor U18280 (N_18280,N_14090,N_15211);
or U18281 (N_18281,N_13472,N_13093);
nor U18282 (N_18282,N_14879,N_14639);
nand U18283 (N_18283,N_12390,N_12055);
xnor U18284 (N_18284,N_15324,N_14243);
or U18285 (N_18285,N_12549,N_14287);
and U18286 (N_18286,N_14773,N_14838);
nand U18287 (N_18287,N_12615,N_13121);
or U18288 (N_18288,N_15592,N_15046);
and U18289 (N_18289,N_13118,N_14079);
nand U18290 (N_18290,N_15092,N_12482);
nand U18291 (N_18291,N_14140,N_13025);
nand U18292 (N_18292,N_13131,N_15013);
or U18293 (N_18293,N_12184,N_14239);
nand U18294 (N_18294,N_14881,N_14277);
nand U18295 (N_18295,N_13721,N_15543);
and U18296 (N_18296,N_12389,N_13907);
nand U18297 (N_18297,N_12426,N_14292);
nor U18298 (N_18298,N_15072,N_14141);
or U18299 (N_18299,N_12805,N_15883);
or U18300 (N_18300,N_13335,N_12579);
nand U18301 (N_18301,N_12332,N_13038);
or U18302 (N_18302,N_12638,N_14536);
nand U18303 (N_18303,N_15601,N_13381);
nand U18304 (N_18304,N_14718,N_13103);
and U18305 (N_18305,N_13748,N_12934);
xor U18306 (N_18306,N_15434,N_13059);
and U18307 (N_18307,N_14027,N_13246);
nand U18308 (N_18308,N_12038,N_13931);
or U18309 (N_18309,N_12269,N_15643);
xnor U18310 (N_18310,N_13685,N_15963);
nand U18311 (N_18311,N_14196,N_12990);
and U18312 (N_18312,N_13810,N_13468);
and U18313 (N_18313,N_14882,N_13146);
and U18314 (N_18314,N_13440,N_15393);
xor U18315 (N_18315,N_14326,N_15082);
nand U18316 (N_18316,N_13480,N_12973);
and U18317 (N_18317,N_15473,N_14768);
nor U18318 (N_18318,N_15578,N_12482);
and U18319 (N_18319,N_12936,N_13415);
and U18320 (N_18320,N_13195,N_14062);
nand U18321 (N_18321,N_13488,N_15019);
and U18322 (N_18322,N_13130,N_12532);
and U18323 (N_18323,N_12129,N_15560);
nor U18324 (N_18324,N_15503,N_15748);
or U18325 (N_18325,N_15391,N_12557);
or U18326 (N_18326,N_14858,N_14336);
and U18327 (N_18327,N_14190,N_13292);
nor U18328 (N_18328,N_13088,N_13199);
nor U18329 (N_18329,N_13735,N_12046);
nor U18330 (N_18330,N_14300,N_12230);
nand U18331 (N_18331,N_15238,N_15558);
xnor U18332 (N_18332,N_13430,N_12512);
nor U18333 (N_18333,N_13792,N_14994);
xnor U18334 (N_18334,N_12019,N_15450);
xor U18335 (N_18335,N_12692,N_15824);
or U18336 (N_18336,N_12216,N_14906);
nor U18337 (N_18337,N_15533,N_13790);
nand U18338 (N_18338,N_12977,N_14630);
or U18339 (N_18339,N_14111,N_15689);
nand U18340 (N_18340,N_14723,N_14211);
or U18341 (N_18341,N_12578,N_14518);
and U18342 (N_18342,N_14294,N_12845);
nand U18343 (N_18343,N_13749,N_14199);
and U18344 (N_18344,N_14060,N_15909);
and U18345 (N_18345,N_14482,N_13951);
nor U18346 (N_18346,N_13756,N_13367);
or U18347 (N_18347,N_12176,N_12279);
nor U18348 (N_18348,N_13507,N_13716);
and U18349 (N_18349,N_13563,N_12344);
nor U18350 (N_18350,N_12580,N_15884);
xnor U18351 (N_18351,N_13515,N_14101);
or U18352 (N_18352,N_14827,N_12626);
nor U18353 (N_18353,N_14261,N_15028);
or U18354 (N_18354,N_15442,N_14185);
and U18355 (N_18355,N_13607,N_12125);
nor U18356 (N_18356,N_13777,N_14536);
or U18357 (N_18357,N_12092,N_15355);
nand U18358 (N_18358,N_14812,N_15548);
or U18359 (N_18359,N_14529,N_14258);
xor U18360 (N_18360,N_15154,N_14538);
and U18361 (N_18361,N_15932,N_14401);
nand U18362 (N_18362,N_12338,N_13260);
and U18363 (N_18363,N_12667,N_14606);
xor U18364 (N_18364,N_12961,N_13361);
and U18365 (N_18365,N_14782,N_15103);
and U18366 (N_18366,N_14310,N_15997);
xor U18367 (N_18367,N_13146,N_13710);
or U18368 (N_18368,N_12956,N_14642);
nor U18369 (N_18369,N_14624,N_12472);
xor U18370 (N_18370,N_15711,N_15604);
or U18371 (N_18371,N_14182,N_13291);
and U18372 (N_18372,N_13492,N_13442);
and U18373 (N_18373,N_14763,N_14321);
or U18374 (N_18374,N_15127,N_15233);
nand U18375 (N_18375,N_13610,N_12970);
or U18376 (N_18376,N_13005,N_12210);
or U18377 (N_18377,N_13634,N_15939);
and U18378 (N_18378,N_13363,N_14705);
nand U18379 (N_18379,N_12257,N_14003);
nand U18380 (N_18380,N_15623,N_13167);
nor U18381 (N_18381,N_14519,N_13452);
and U18382 (N_18382,N_13983,N_15379);
and U18383 (N_18383,N_13303,N_14231);
or U18384 (N_18384,N_12810,N_14112);
nor U18385 (N_18385,N_15157,N_15231);
xnor U18386 (N_18386,N_15916,N_13559);
or U18387 (N_18387,N_14108,N_15987);
nand U18388 (N_18388,N_15166,N_12605);
nand U18389 (N_18389,N_12108,N_14251);
nor U18390 (N_18390,N_12742,N_14468);
or U18391 (N_18391,N_12891,N_12948);
and U18392 (N_18392,N_15084,N_15197);
xnor U18393 (N_18393,N_14795,N_13329);
and U18394 (N_18394,N_12487,N_15925);
or U18395 (N_18395,N_12082,N_12639);
xor U18396 (N_18396,N_13289,N_12083);
nor U18397 (N_18397,N_15362,N_14511);
or U18398 (N_18398,N_15333,N_15966);
nor U18399 (N_18399,N_15202,N_13711);
xor U18400 (N_18400,N_15626,N_12627);
nor U18401 (N_18401,N_14019,N_15885);
nand U18402 (N_18402,N_12949,N_14852);
xor U18403 (N_18403,N_12247,N_12548);
xnor U18404 (N_18404,N_13075,N_14883);
and U18405 (N_18405,N_12962,N_14630);
and U18406 (N_18406,N_13520,N_15715);
nor U18407 (N_18407,N_12364,N_12965);
and U18408 (N_18408,N_12667,N_12689);
and U18409 (N_18409,N_12413,N_14259);
or U18410 (N_18410,N_14216,N_12186);
nand U18411 (N_18411,N_12203,N_14586);
nor U18412 (N_18412,N_14065,N_12802);
nor U18413 (N_18413,N_15935,N_12815);
and U18414 (N_18414,N_13381,N_12715);
nand U18415 (N_18415,N_13988,N_14738);
nor U18416 (N_18416,N_15157,N_14345);
nand U18417 (N_18417,N_12270,N_12127);
xor U18418 (N_18418,N_12894,N_12361);
nor U18419 (N_18419,N_12881,N_14070);
nand U18420 (N_18420,N_12995,N_13941);
or U18421 (N_18421,N_13755,N_15206);
or U18422 (N_18422,N_12707,N_15666);
and U18423 (N_18423,N_14481,N_14432);
xnor U18424 (N_18424,N_12134,N_12556);
nor U18425 (N_18425,N_13469,N_13802);
and U18426 (N_18426,N_14082,N_15845);
nor U18427 (N_18427,N_13342,N_14947);
and U18428 (N_18428,N_13107,N_15013);
or U18429 (N_18429,N_14984,N_12718);
or U18430 (N_18430,N_12626,N_12176);
nand U18431 (N_18431,N_15823,N_12454);
nand U18432 (N_18432,N_15334,N_15215);
or U18433 (N_18433,N_15206,N_13179);
nand U18434 (N_18434,N_14222,N_14737);
nand U18435 (N_18435,N_13982,N_15806);
and U18436 (N_18436,N_12750,N_13347);
nand U18437 (N_18437,N_13835,N_13596);
or U18438 (N_18438,N_12649,N_14683);
or U18439 (N_18439,N_14497,N_15810);
or U18440 (N_18440,N_15206,N_13524);
or U18441 (N_18441,N_14704,N_14877);
nor U18442 (N_18442,N_12737,N_15880);
nand U18443 (N_18443,N_12202,N_13625);
xnor U18444 (N_18444,N_13911,N_12292);
nor U18445 (N_18445,N_15321,N_12871);
and U18446 (N_18446,N_12577,N_15412);
or U18447 (N_18447,N_14391,N_13211);
nor U18448 (N_18448,N_13190,N_14759);
nor U18449 (N_18449,N_13569,N_13418);
and U18450 (N_18450,N_15521,N_14041);
nand U18451 (N_18451,N_15337,N_15539);
or U18452 (N_18452,N_14490,N_12968);
nand U18453 (N_18453,N_15873,N_14670);
and U18454 (N_18454,N_15438,N_13773);
and U18455 (N_18455,N_15087,N_13220);
nand U18456 (N_18456,N_14422,N_14011);
or U18457 (N_18457,N_12237,N_15837);
nand U18458 (N_18458,N_12075,N_14369);
nor U18459 (N_18459,N_14294,N_14972);
nand U18460 (N_18460,N_12081,N_13582);
or U18461 (N_18461,N_12917,N_12176);
nor U18462 (N_18462,N_14762,N_14575);
or U18463 (N_18463,N_15109,N_15378);
nor U18464 (N_18464,N_14648,N_13335);
nor U18465 (N_18465,N_14377,N_13777);
nand U18466 (N_18466,N_13380,N_13456);
xor U18467 (N_18467,N_12088,N_13446);
and U18468 (N_18468,N_15374,N_14105);
nor U18469 (N_18469,N_12463,N_15234);
or U18470 (N_18470,N_14341,N_13787);
nand U18471 (N_18471,N_14210,N_13583);
or U18472 (N_18472,N_15261,N_14136);
nand U18473 (N_18473,N_15487,N_15846);
or U18474 (N_18474,N_13750,N_15748);
or U18475 (N_18475,N_12798,N_12154);
or U18476 (N_18476,N_15362,N_15699);
nor U18477 (N_18477,N_14029,N_12665);
and U18478 (N_18478,N_12191,N_13753);
nor U18479 (N_18479,N_12350,N_13772);
and U18480 (N_18480,N_14470,N_13926);
and U18481 (N_18481,N_14467,N_13062);
nor U18482 (N_18482,N_13494,N_15361);
or U18483 (N_18483,N_14413,N_15577);
nand U18484 (N_18484,N_13731,N_12262);
xnor U18485 (N_18485,N_15714,N_12622);
nand U18486 (N_18486,N_14048,N_13348);
and U18487 (N_18487,N_14508,N_12525);
or U18488 (N_18488,N_12383,N_13254);
nand U18489 (N_18489,N_14921,N_14753);
or U18490 (N_18490,N_12143,N_15287);
nand U18491 (N_18491,N_15884,N_13569);
and U18492 (N_18492,N_13685,N_13200);
or U18493 (N_18493,N_15413,N_13117);
and U18494 (N_18494,N_14879,N_14482);
and U18495 (N_18495,N_13744,N_13076);
or U18496 (N_18496,N_14980,N_15624);
and U18497 (N_18497,N_15729,N_14056);
and U18498 (N_18498,N_13591,N_13100);
nor U18499 (N_18499,N_14744,N_15626);
nor U18500 (N_18500,N_14694,N_13326);
nand U18501 (N_18501,N_14902,N_14357);
nand U18502 (N_18502,N_15615,N_14967);
nand U18503 (N_18503,N_14681,N_14276);
nor U18504 (N_18504,N_13004,N_15307);
nand U18505 (N_18505,N_15729,N_15127);
or U18506 (N_18506,N_12985,N_12806);
nor U18507 (N_18507,N_13799,N_13460);
nand U18508 (N_18508,N_13853,N_12807);
nand U18509 (N_18509,N_13943,N_15839);
nor U18510 (N_18510,N_13547,N_12411);
nor U18511 (N_18511,N_12917,N_15937);
and U18512 (N_18512,N_14495,N_14386);
xor U18513 (N_18513,N_14347,N_14094);
nor U18514 (N_18514,N_14443,N_14001);
nand U18515 (N_18515,N_14681,N_13953);
or U18516 (N_18516,N_15351,N_14725);
and U18517 (N_18517,N_14576,N_14704);
nand U18518 (N_18518,N_14957,N_15103);
nand U18519 (N_18519,N_13871,N_14602);
and U18520 (N_18520,N_15362,N_15604);
nand U18521 (N_18521,N_12488,N_14766);
nand U18522 (N_18522,N_13854,N_15802);
nand U18523 (N_18523,N_12258,N_14847);
or U18524 (N_18524,N_15509,N_14948);
or U18525 (N_18525,N_15279,N_13702);
or U18526 (N_18526,N_13326,N_12390);
nor U18527 (N_18527,N_12502,N_15333);
or U18528 (N_18528,N_13089,N_15212);
xnor U18529 (N_18529,N_15710,N_12873);
or U18530 (N_18530,N_12004,N_15681);
nand U18531 (N_18531,N_13733,N_15771);
and U18532 (N_18532,N_15972,N_14885);
nor U18533 (N_18533,N_15273,N_13725);
and U18534 (N_18534,N_13522,N_15583);
nor U18535 (N_18535,N_12182,N_15747);
and U18536 (N_18536,N_15580,N_12433);
nand U18537 (N_18537,N_12659,N_13922);
and U18538 (N_18538,N_15910,N_12581);
or U18539 (N_18539,N_15213,N_15949);
or U18540 (N_18540,N_13250,N_14695);
nand U18541 (N_18541,N_15587,N_14660);
and U18542 (N_18542,N_12494,N_15023);
nand U18543 (N_18543,N_14585,N_13940);
and U18544 (N_18544,N_15794,N_15494);
or U18545 (N_18545,N_13172,N_15908);
nor U18546 (N_18546,N_12755,N_12973);
nand U18547 (N_18547,N_12251,N_13966);
or U18548 (N_18548,N_12283,N_13708);
nor U18549 (N_18549,N_13013,N_12179);
or U18550 (N_18550,N_14809,N_12056);
nand U18551 (N_18551,N_12469,N_15476);
or U18552 (N_18552,N_15078,N_15384);
or U18553 (N_18553,N_14108,N_12560);
and U18554 (N_18554,N_12901,N_14281);
or U18555 (N_18555,N_12063,N_14347);
or U18556 (N_18556,N_14486,N_12696);
or U18557 (N_18557,N_14810,N_14182);
xor U18558 (N_18558,N_12880,N_13489);
nor U18559 (N_18559,N_15052,N_15176);
and U18560 (N_18560,N_15119,N_14476);
nand U18561 (N_18561,N_15330,N_13032);
nand U18562 (N_18562,N_13279,N_12210);
nand U18563 (N_18563,N_13269,N_13839);
and U18564 (N_18564,N_13345,N_12864);
nor U18565 (N_18565,N_15919,N_14286);
and U18566 (N_18566,N_14890,N_14040);
and U18567 (N_18567,N_12993,N_14378);
nor U18568 (N_18568,N_12519,N_13176);
nand U18569 (N_18569,N_14201,N_15091);
or U18570 (N_18570,N_15073,N_14067);
nand U18571 (N_18571,N_13067,N_14857);
or U18572 (N_18572,N_13229,N_14090);
xor U18573 (N_18573,N_15898,N_15092);
or U18574 (N_18574,N_12428,N_13923);
nand U18575 (N_18575,N_14928,N_13189);
xnor U18576 (N_18576,N_14758,N_14919);
nor U18577 (N_18577,N_12015,N_12477);
nor U18578 (N_18578,N_15773,N_13008);
and U18579 (N_18579,N_14304,N_12363);
and U18580 (N_18580,N_14830,N_13389);
and U18581 (N_18581,N_14787,N_12217);
or U18582 (N_18582,N_15457,N_13077);
nor U18583 (N_18583,N_12732,N_12466);
or U18584 (N_18584,N_13132,N_12719);
nand U18585 (N_18585,N_15834,N_15003);
and U18586 (N_18586,N_13562,N_13670);
and U18587 (N_18587,N_15523,N_15059);
and U18588 (N_18588,N_12772,N_13463);
nor U18589 (N_18589,N_12120,N_14949);
and U18590 (N_18590,N_12574,N_14899);
nor U18591 (N_18591,N_14068,N_13734);
nand U18592 (N_18592,N_13300,N_12735);
and U18593 (N_18593,N_14600,N_13422);
nor U18594 (N_18594,N_12643,N_12063);
nor U18595 (N_18595,N_13059,N_15084);
xor U18596 (N_18596,N_14574,N_12575);
nand U18597 (N_18597,N_12131,N_14571);
or U18598 (N_18598,N_13968,N_13119);
nand U18599 (N_18599,N_15227,N_14941);
or U18600 (N_18600,N_14202,N_14887);
and U18601 (N_18601,N_14932,N_14808);
or U18602 (N_18602,N_15152,N_14653);
and U18603 (N_18603,N_13272,N_14530);
xnor U18604 (N_18604,N_15724,N_15088);
or U18605 (N_18605,N_15513,N_13675);
and U18606 (N_18606,N_12548,N_12435);
nor U18607 (N_18607,N_14399,N_15922);
and U18608 (N_18608,N_15898,N_13815);
and U18609 (N_18609,N_15438,N_15833);
nor U18610 (N_18610,N_15882,N_12511);
nor U18611 (N_18611,N_14048,N_13270);
nand U18612 (N_18612,N_12498,N_15819);
and U18613 (N_18613,N_13479,N_12411);
xnor U18614 (N_18614,N_13534,N_14002);
or U18615 (N_18615,N_14626,N_13028);
nand U18616 (N_18616,N_14555,N_12785);
and U18617 (N_18617,N_12867,N_13694);
and U18618 (N_18618,N_15890,N_12204);
and U18619 (N_18619,N_14253,N_12950);
and U18620 (N_18620,N_14011,N_12916);
and U18621 (N_18621,N_14549,N_14103);
xor U18622 (N_18622,N_12403,N_13230);
and U18623 (N_18623,N_15111,N_12503);
nor U18624 (N_18624,N_14864,N_15702);
and U18625 (N_18625,N_13160,N_13797);
xor U18626 (N_18626,N_14043,N_14618);
and U18627 (N_18627,N_13987,N_15378);
and U18628 (N_18628,N_14464,N_13124);
and U18629 (N_18629,N_15191,N_13614);
nor U18630 (N_18630,N_15708,N_14134);
nor U18631 (N_18631,N_14047,N_12849);
or U18632 (N_18632,N_14661,N_13408);
nor U18633 (N_18633,N_14318,N_12779);
or U18634 (N_18634,N_14369,N_12726);
nor U18635 (N_18635,N_12376,N_12838);
nor U18636 (N_18636,N_14023,N_15111);
or U18637 (N_18637,N_12760,N_12966);
and U18638 (N_18638,N_14123,N_14417);
and U18639 (N_18639,N_15780,N_13575);
nand U18640 (N_18640,N_12763,N_13752);
nand U18641 (N_18641,N_15297,N_15648);
or U18642 (N_18642,N_12494,N_15155);
nand U18643 (N_18643,N_15662,N_13977);
or U18644 (N_18644,N_15554,N_14111);
or U18645 (N_18645,N_12209,N_15015);
xnor U18646 (N_18646,N_13183,N_15390);
nor U18647 (N_18647,N_14413,N_14937);
nand U18648 (N_18648,N_12731,N_12159);
or U18649 (N_18649,N_13892,N_13264);
and U18650 (N_18650,N_12221,N_12358);
or U18651 (N_18651,N_14792,N_14247);
and U18652 (N_18652,N_14390,N_13226);
nor U18653 (N_18653,N_14431,N_14491);
or U18654 (N_18654,N_13629,N_12819);
and U18655 (N_18655,N_14397,N_12654);
or U18656 (N_18656,N_14115,N_15236);
nor U18657 (N_18657,N_15753,N_13313);
and U18658 (N_18658,N_14435,N_13824);
nand U18659 (N_18659,N_15820,N_15892);
nand U18660 (N_18660,N_15730,N_12354);
xnor U18661 (N_18661,N_13905,N_14086);
or U18662 (N_18662,N_14083,N_15185);
and U18663 (N_18663,N_14882,N_14746);
and U18664 (N_18664,N_13889,N_14892);
or U18665 (N_18665,N_14303,N_13842);
and U18666 (N_18666,N_15688,N_12158);
nor U18667 (N_18667,N_13868,N_12024);
nand U18668 (N_18668,N_13391,N_13238);
or U18669 (N_18669,N_14058,N_13247);
nand U18670 (N_18670,N_13759,N_14178);
or U18671 (N_18671,N_15276,N_13919);
xnor U18672 (N_18672,N_15413,N_13677);
nor U18673 (N_18673,N_15643,N_14135);
and U18674 (N_18674,N_15468,N_12692);
and U18675 (N_18675,N_15480,N_14703);
or U18676 (N_18676,N_12402,N_12878);
nor U18677 (N_18677,N_12047,N_14214);
or U18678 (N_18678,N_13958,N_13461);
and U18679 (N_18679,N_15876,N_12500);
xnor U18680 (N_18680,N_13545,N_14367);
nor U18681 (N_18681,N_13541,N_13875);
and U18682 (N_18682,N_12889,N_12257);
nand U18683 (N_18683,N_14478,N_15275);
nand U18684 (N_18684,N_12165,N_12131);
and U18685 (N_18685,N_12773,N_12307);
xnor U18686 (N_18686,N_14333,N_12744);
or U18687 (N_18687,N_14856,N_15946);
and U18688 (N_18688,N_14535,N_12429);
nor U18689 (N_18689,N_12422,N_15820);
nor U18690 (N_18690,N_14872,N_14557);
or U18691 (N_18691,N_13104,N_13064);
xor U18692 (N_18692,N_15044,N_12396);
nor U18693 (N_18693,N_13227,N_13862);
or U18694 (N_18694,N_13980,N_13779);
nor U18695 (N_18695,N_13625,N_15827);
nand U18696 (N_18696,N_15752,N_13400);
xor U18697 (N_18697,N_15619,N_15336);
nand U18698 (N_18698,N_14822,N_12350);
or U18699 (N_18699,N_12423,N_12340);
xor U18700 (N_18700,N_14771,N_14294);
or U18701 (N_18701,N_14140,N_12661);
nand U18702 (N_18702,N_12737,N_15760);
nand U18703 (N_18703,N_15724,N_12290);
nor U18704 (N_18704,N_15155,N_14394);
or U18705 (N_18705,N_12828,N_15161);
nand U18706 (N_18706,N_14101,N_13230);
xnor U18707 (N_18707,N_12200,N_14047);
nand U18708 (N_18708,N_15137,N_15494);
nor U18709 (N_18709,N_15508,N_15566);
or U18710 (N_18710,N_14367,N_13516);
nand U18711 (N_18711,N_14924,N_14174);
nand U18712 (N_18712,N_12241,N_15962);
and U18713 (N_18713,N_15518,N_13118);
nor U18714 (N_18714,N_12984,N_15338);
or U18715 (N_18715,N_15389,N_14350);
nor U18716 (N_18716,N_12620,N_14520);
nand U18717 (N_18717,N_13688,N_14187);
nor U18718 (N_18718,N_15517,N_14473);
or U18719 (N_18719,N_14573,N_14469);
and U18720 (N_18720,N_13535,N_15356);
xnor U18721 (N_18721,N_12520,N_12740);
nand U18722 (N_18722,N_12127,N_15533);
nor U18723 (N_18723,N_14407,N_12934);
or U18724 (N_18724,N_15853,N_14985);
nand U18725 (N_18725,N_15845,N_14480);
nand U18726 (N_18726,N_14686,N_13267);
and U18727 (N_18727,N_15496,N_12159);
or U18728 (N_18728,N_12341,N_13335);
or U18729 (N_18729,N_15064,N_14234);
nand U18730 (N_18730,N_15411,N_13969);
and U18731 (N_18731,N_14827,N_15674);
nand U18732 (N_18732,N_13033,N_13704);
and U18733 (N_18733,N_15674,N_15600);
nand U18734 (N_18734,N_12284,N_12797);
and U18735 (N_18735,N_13072,N_13605);
or U18736 (N_18736,N_14665,N_13549);
or U18737 (N_18737,N_13849,N_14621);
and U18738 (N_18738,N_13300,N_14061);
or U18739 (N_18739,N_13873,N_14715);
and U18740 (N_18740,N_14453,N_14998);
nor U18741 (N_18741,N_12419,N_12835);
and U18742 (N_18742,N_12061,N_12067);
and U18743 (N_18743,N_12918,N_12514);
or U18744 (N_18744,N_12660,N_12494);
xor U18745 (N_18745,N_14635,N_12146);
nor U18746 (N_18746,N_12662,N_15756);
or U18747 (N_18747,N_15916,N_12149);
nor U18748 (N_18748,N_14161,N_13788);
nand U18749 (N_18749,N_13400,N_15504);
nor U18750 (N_18750,N_13616,N_15433);
or U18751 (N_18751,N_14770,N_13677);
or U18752 (N_18752,N_13487,N_15622);
nand U18753 (N_18753,N_15460,N_12853);
or U18754 (N_18754,N_15082,N_13674);
nand U18755 (N_18755,N_14968,N_15895);
or U18756 (N_18756,N_13362,N_12774);
and U18757 (N_18757,N_14081,N_15365);
or U18758 (N_18758,N_14281,N_14404);
and U18759 (N_18759,N_12147,N_13315);
or U18760 (N_18760,N_15317,N_12166);
or U18761 (N_18761,N_12297,N_12305);
nand U18762 (N_18762,N_12598,N_15194);
nand U18763 (N_18763,N_15056,N_14792);
and U18764 (N_18764,N_14783,N_15817);
xnor U18765 (N_18765,N_12476,N_12630);
nor U18766 (N_18766,N_12000,N_13054);
or U18767 (N_18767,N_15950,N_14140);
or U18768 (N_18768,N_14227,N_14499);
nor U18769 (N_18769,N_15607,N_15846);
and U18770 (N_18770,N_13943,N_12187);
xor U18771 (N_18771,N_12514,N_12304);
or U18772 (N_18772,N_14767,N_15150);
or U18773 (N_18773,N_14466,N_14222);
nor U18774 (N_18774,N_12364,N_15580);
nand U18775 (N_18775,N_15580,N_13847);
and U18776 (N_18776,N_12948,N_15789);
nand U18777 (N_18777,N_12153,N_13453);
nor U18778 (N_18778,N_15533,N_12640);
or U18779 (N_18779,N_14017,N_13716);
or U18780 (N_18780,N_14065,N_15352);
nor U18781 (N_18781,N_14129,N_13296);
and U18782 (N_18782,N_12199,N_13569);
and U18783 (N_18783,N_15167,N_12969);
and U18784 (N_18784,N_12127,N_13519);
or U18785 (N_18785,N_12595,N_14938);
nor U18786 (N_18786,N_13328,N_13191);
and U18787 (N_18787,N_14960,N_14657);
nand U18788 (N_18788,N_14543,N_12975);
nand U18789 (N_18789,N_14685,N_12238);
and U18790 (N_18790,N_12146,N_15282);
nand U18791 (N_18791,N_15468,N_13268);
nand U18792 (N_18792,N_12215,N_13336);
nand U18793 (N_18793,N_12240,N_13185);
or U18794 (N_18794,N_15810,N_15764);
nand U18795 (N_18795,N_14650,N_12062);
nor U18796 (N_18796,N_15748,N_15708);
nand U18797 (N_18797,N_13538,N_12222);
and U18798 (N_18798,N_13341,N_12466);
xnor U18799 (N_18799,N_15166,N_12102);
nor U18800 (N_18800,N_15564,N_15113);
or U18801 (N_18801,N_13861,N_15839);
nor U18802 (N_18802,N_14558,N_15155);
nor U18803 (N_18803,N_13044,N_13097);
nand U18804 (N_18804,N_15236,N_15778);
or U18805 (N_18805,N_13910,N_12637);
and U18806 (N_18806,N_15135,N_12741);
or U18807 (N_18807,N_12011,N_13595);
nand U18808 (N_18808,N_15573,N_15243);
or U18809 (N_18809,N_15774,N_13160);
nand U18810 (N_18810,N_15235,N_14523);
nand U18811 (N_18811,N_12214,N_12564);
or U18812 (N_18812,N_14434,N_14727);
or U18813 (N_18813,N_15118,N_12783);
or U18814 (N_18814,N_14499,N_14091);
or U18815 (N_18815,N_14464,N_13459);
or U18816 (N_18816,N_14812,N_14541);
nand U18817 (N_18817,N_15740,N_13358);
or U18818 (N_18818,N_14317,N_12125);
xor U18819 (N_18819,N_15132,N_15409);
or U18820 (N_18820,N_13491,N_12569);
nor U18821 (N_18821,N_14429,N_13487);
nor U18822 (N_18822,N_13021,N_12818);
and U18823 (N_18823,N_12036,N_15301);
or U18824 (N_18824,N_12396,N_14471);
and U18825 (N_18825,N_12100,N_13570);
and U18826 (N_18826,N_12632,N_15084);
nor U18827 (N_18827,N_15548,N_14411);
nand U18828 (N_18828,N_14986,N_15482);
or U18829 (N_18829,N_15275,N_14469);
xor U18830 (N_18830,N_14818,N_12048);
xnor U18831 (N_18831,N_13135,N_15088);
and U18832 (N_18832,N_14446,N_13052);
or U18833 (N_18833,N_12792,N_12267);
nand U18834 (N_18834,N_13723,N_15058);
and U18835 (N_18835,N_13278,N_14266);
and U18836 (N_18836,N_14083,N_14030);
and U18837 (N_18837,N_12092,N_12377);
xnor U18838 (N_18838,N_15822,N_12719);
nand U18839 (N_18839,N_13600,N_15623);
nor U18840 (N_18840,N_15197,N_12485);
or U18841 (N_18841,N_12921,N_15961);
or U18842 (N_18842,N_15088,N_13165);
nand U18843 (N_18843,N_13822,N_14775);
or U18844 (N_18844,N_13640,N_12145);
xor U18845 (N_18845,N_12983,N_15787);
nor U18846 (N_18846,N_14272,N_15126);
and U18847 (N_18847,N_12018,N_14102);
nor U18848 (N_18848,N_15865,N_15910);
nor U18849 (N_18849,N_13794,N_13228);
or U18850 (N_18850,N_14223,N_14386);
nor U18851 (N_18851,N_13061,N_14132);
and U18852 (N_18852,N_12455,N_15962);
nor U18853 (N_18853,N_13683,N_13492);
nand U18854 (N_18854,N_12209,N_13934);
nor U18855 (N_18855,N_15753,N_15679);
or U18856 (N_18856,N_13339,N_13650);
xnor U18857 (N_18857,N_13977,N_13937);
or U18858 (N_18858,N_12695,N_15019);
xor U18859 (N_18859,N_12476,N_14186);
nand U18860 (N_18860,N_12728,N_13615);
and U18861 (N_18861,N_12219,N_14065);
nor U18862 (N_18862,N_13246,N_15382);
nand U18863 (N_18863,N_12150,N_13456);
nor U18864 (N_18864,N_12038,N_13670);
nor U18865 (N_18865,N_12474,N_14802);
and U18866 (N_18866,N_15864,N_12154);
nor U18867 (N_18867,N_12402,N_13002);
and U18868 (N_18868,N_13612,N_13196);
and U18869 (N_18869,N_13763,N_14240);
nand U18870 (N_18870,N_15403,N_14065);
xor U18871 (N_18871,N_14213,N_15162);
nand U18872 (N_18872,N_15383,N_15227);
nand U18873 (N_18873,N_14182,N_14642);
and U18874 (N_18874,N_15198,N_15913);
nand U18875 (N_18875,N_14578,N_14435);
nor U18876 (N_18876,N_12843,N_13564);
or U18877 (N_18877,N_14288,N_15653);
xnor U18878 (N_18878,N_15731,N_13750);
or U18879 (N_18879,N_15311,N_12308);
and U18880 (N_18880,N_14345,N_12646);
nand U18881 (N_18881,N_14643,N_12401);
and U18882 (N_18882,N_14181,N_15563);
xnor U18883 (N_18883,N_12979,N_13426);
nor U18884 (N_18884,N_14453,N_12248);
nand U18885 (N_18885,N_14542,N_12894);
xor U18886 (N_18886,N_12467,N_14510);
or U18887 (N_18887,N_12756,N_15214);
nor U18888 (N_18888,N_15811,N_12754);
nor U18889 (N_18889,N_14573,N_12891);
xor U18890 (N_18890,N_14608,N_14035);
xor U18891 (N_18891,N_15834,N_12622);
or U18892 (N_18892,N_12607,N_13549);
nor U18893 (N_18893,N_15189,N_14767);
nand U18894 (N_18894,N_12342,N_15592);
or U18895 (N_18895,N_13748,N_14307);
nand U18896 (N_18896,N_14820,N_14878);
nor U18897 (N_18897,N_13550,N_15704);
xnor U18898 (N_18898,N_15232,N_13210);
and U18899 (N_18899,N_15841,N_12594);
xor U18900 (N_18900,N_14016,N_15015);
nor U18901 (N_18901,N_13765,N_15675);
and U18902 (N_18902,N_15252,N_12596);
xor U18903 (N_18903,N_15190,N_12233);
nor U18904 (N_18904,N_12332,N_12203);
nor U18905 (N_18905,N_12754,N_14171);
nand U18906 (N_18906,N_13177,N_13478);
nor U18907 (N_18907,N_14277,N_15871);
and U18908 (N_18908,N_12752,N_14017);
nand U18909 (N_18909,N_15620,N_13087);
or U18910 (N_18910,N_12197,N_12676);
and U18911 (N_18911,N_15231,N_14364);
and U18912 (N_18912,N_15763,N_14828);
nand U18913 (N_18913,N_14087,N_14810);
and U18914 (N_18914,N_15694,N_12332);
nor U18915 (N_18915,N_13478,N_14678);
nand U18916 (N_18916,N_15869,N_15202);
nand U18917 (N_18917,N_13567,N_15471);
or U18918 (N_18918,N_12286,N_13543);
or U18919 (N_18919,N_15098,N_14105);
nor U18920 (N_18920,N_14046,N_12144);
or U18921 (N_18921,N_15036,N_13616);
or U18922 (N_18922,N_15315,N_14427);
xor U18923 (N_18923,N_12596,N_14665);
and U18924 (N_18924,N_13251,N_14558);
and U18925 (N_18925,N_15403,N_15777);
nor U18926 (N_18926,N_12479,N_12909);
nand U18927 (N_18927,N_13341,N_13550);
xnor U18928 (N_18928,N_12250,N_12043);
nor U18929 (N_18929,N_13794,N_12669);
nand U18930 (N_18930,N_14131,N_15366);
nand U18931 (N_18931,N_15458,N_14956);
nor U18932 (N_18932,N_12040,N_14540);
nand U18933 (N_18933,N_13066,N_15510);
nand U18934 (N_18934,N_12257,N_14775);
or U18935 (N_18935,N_14299,N_14124);
and U18936 (N_18936,N_12108,N_15871);
xnor U18937 (N_18937,N_14305,N_13252);
nor U18938 (N_18938,N_15945,N_15219);
and U18939 (N_18939,N_13847,N_14989);
or U18940 (N_18940,N_14105,N_15057);
nor U18941 (N_18941,N_13092,N_14447);
nor U18942 (N_18942,N_13934,N_15833);
nand U18943 (N_18943,N_15508,N_12619);
or U18944 (N_18944,N_15651,N_15180);
or U18945 (N_18945,N_14350,N_15005);
or U18946 (N_18946,N_14179,N_15052);
nand U18947 (N_18947,N_15288,N_12194);
nor U18948 (N_18948,N_14454,N_15666);
xnor U18949 (N_18949,N_14225,N_12605);
and U18950 (N_18950,N_13809,N_15654);
and U18951 (N_18951,N_12586,N_12943);
nor U18952 (N_18952,N_13363,N_13963);
or U18953 (N_18953,N_14056,N_13419);
nor U18954 (N_18954,N_14116,N_15800);
or U18955 (N_18955,N_12479,N_13749);
nor U18956 (N_18956,N_12258,N_14697);
nand U18957 (N_18957,N_14189,N_14789);
or U18958 (N_18958,N_15040,N_15442);
nand U18959 (N_18959,N_15002,N_12040);
nand U18960 (N_18960,N_14628,N_14566);
nand U18961 (N_18961,N_13660,N_15047);
nand U18962 (N_18962,N_12087,N_15937);
or U18963 (N_18963,N_13364,N_12162);
nor U18964 (N_18964,N_15679,N_13461);
xor U18965 (N_18965,N_13912,N_13579);
nand U18966 (N_18966,N_14517,N_14109);
or U18967 (N_18967,N_13986,N_13074);
nor U18968 (N_18968,N_15969,N_13581);
nor U18969 (N_18969,N_14758,N_12978);
nand U18970 (N_18970,N_12531,N_13033);
or U18971 (N_18971,N_14474,N_12325);
and U18972 (N_18972,N_13103,N_14777);
nand U18973 (N_18973,N_13484,N_15952);
nand U18974 (N_18974,N_15565,N_15484);
nor U18975 (N_18975,N_15668,N_14131);
and U18976 (N_18976,N_12592,N_13342);
nand U18977 (N_18977,N_13275,N_12411);
and U18978 (N_18978,N_13360,N_12820);
and U18979 (N_18979,N_13484,N_12232);
nor U18980 (N_18980,N_15966,N_14503);
nand U18981 (N_18981,N_13463,N_13753);
or U18982 (N_18982,N_14862,N_14024);
nor U18983 (N_18983,N_13508,N_13569);
nand U18984 (N_18984,N_13807,N_12610);
or U18985 (N_18985,N_15296,N_15800);
and U18986 (N_18986,N_12714,N_12671);
nand U18987 (N_18987,N_15947,N_13328);
xor U18988 (N_18988,N_13669,N_15588);
nand U18989 (N_18989,N_15067,N_13051);
or U18990 (N_18990,N_15398,N_13505);
or U18991 (N_18991,N_13968,N_15928);
or U18992 (N_18992,N_13883,N_12977);
or U18993 (N_18993,N_13987,N_13440);
xor U18994 (N_18994,N_13051,N_15453);
and U18995 (N_18995,N_13264,N_14201);
nand U18996 (N_18996,N_14105,N_14776);
nand U18997 (N_18997,N_15038,N_14275);
nor U18998 (N_18998,N_14876,N_15310);
nand U18999 (N_18999,N_12999,N_14928);
and U19000 (N_19000,N_12234,N_13133);
and U19001 (N_19001,N_15473,N_14717);
nand U19002 (N_19002,N_14704,N_14002);
nand U19003 (N_19003,N_14663,N_14620);
xor U19004 (N_19004,N_15215,N_15205);
xor U19005 (N_19005,N_14528,N_12858);
or U19006 (N_19006,N_14532,N_13981);
xnor U19007 (N_19007,N_14871,N_13279);
or U19008 (N_19008,N_14710,N_15997);
xnor U19009 (N_19009,N_13746,N_13115);
nor U19010 (N_19010,N_13318,N_12132);
nand U19011 (N_19011,N_13948,N_14744);
nand U19012 (N_19012,N_13269,N_12864);
nand U19013 (N_19013,N_15521,N_15260);
nor U19014 (N_19014,N_14878,N_13587);
and U19015 (N_19015,N_14398,N_15251);
and U19016 (N_19016,N_12504,N_13325);
nor U19017 (N_19017,N_14051,N_15716);
and U19018 (N_19018,N_15726,N_12769);
or U19019 (N_19019,N_15448,N_13022);
xnor U19020 (N_19020,N_12607,N_13218);
and U19021 (N_19021,N_13728,N_14839);
nand U19022 (N_19022,N_12444,N_14851);
or U19023 (N_19023,N_15124,N_13638);
xor U19024 (N_19024,N_15709,N_14468);
or U19025 (N_19025,N_13305,N_12530);
nor U19026 (N_19026,N_15828,N_13862);
and U19027 (N_19027,N_13194,N_13928);
nand U19028 (N_19028,N_15256,N_12520);
nor U19029 (N_19029,N_13421,N_14777);
nand U19030 (N_19030,N_15491,N_12595);
nand U19031 (N_19031,N_15595,N_13654);
and U19032 (N_19032,N_14707,N_14289);
nand U19033 (N_19033,N_13393,N_12834);
and U19034 (N_19034,N_13421,N_14149);
and U19035 (N_19035,N_12452,N_15018);
xnor U19036 (N_19036,N_14645,N_12593);
or U19037 (N_19037,N_12881,N_12788);
and U19038 (N_19038,N_14769,N_15629);
and U19039 (N_19039,N_14702,N_14354);
nand U19040 (N_19040,N_12621,N_15986);
or U19041 (N_19041,N_12500,N_12077);
nand U19042 (N_19042,N_14669,N_13823);
and U19043 (N_19043,N_13507,N_13451);
xnor U19044 (N_19044,N_15462,N_15022);
or U19045 (N_19045,N_13138,N_13509);
or U19046 (N_19046,N_15633,N_15399);
nor U19047 (N_19047,N_15186,N_14177);
nor U19048 (N_19048,N_13164,N_14056);
and U19049 (N_19049,N_14300,N_13304);
nor U19050 (N_19050,N_15838,N_15550);
and U19051 (N_19051,N_12974,N_14827);
nand U19052 (N_19052,N_15770,N_12564);
nor U19053 (N_19053,N_15817,N_15371);
or U19054 (N_19054,N_12075,N_14375);
and U19055 (N_19055,N_12632,N_13649);
or U19056 (N_19056,N_15723,N_14174);
nand U19057 (N_19057,N_15971,N_14855);
or U19058 (N_19058,N_12215,N_15118);
nor U19059 (N_19059,N_12957,N_14264);
and U19060 (N_19060,N_13123,N_15674);
nand U19061 (N_19061,N_13873,N_12457);
xor U19062 (N_19062,N_14527,N_15336);
nand U19063 (N_19063,N_15581,N_14731);
nand U19064 (N_19064,N_12667,N_13004);
nor U19065 (N_19065,N_15556,N_14221);
nand U19066 (N_19066,N_14216,N_15582);
nor U19067 (N_19067,N_14746,N_14830);
xor U19068 (N_19068,N_15288,N_15484);
nor U19069 (N_19069,N_14080,N_13337);
or U19070 (N_19070,N_13020,N_12987);
nand U19071 (N_19071,N_15971,N_15817);
or U19072 (N_19072,N_13828,N_13251);
and U19073 (N_19073,N_12884,N_13111);
xor U19074 (N_19074,N_13293,N_14371);
or U19075 (N_19075,N_15255,N_14293);
and U19076 (N_19076,N_12481,N_12010);
nand U19077 (N_19077,N_14585,N_12889);
nand U19078 (N_19078,N_14347,N_14943);
and U19079 (N_19079,N_13331,N_12587);
nor U19080 (N_19080,N_14831,N_12165);
nand U19081 (N_19081,N_12369,N_15632);
and U19082 (N_19082,N_15618,N_14757);
and U19083 (N_19083,N_12843,N_15373);
or U19084 (N_19084,N_15749,N_13874);
nand U19085 (N_19085,N_12521,N_12669);
and U19086 (N_19086,N_12302,N_14045);
or U19087 (N_19087,N_14192,N_14698);
or U19088 (N_19088,N_13084,N_12395);
and U19089 (N_19089,N_15379,N_14832);
or U19090 (N_19090,N_15986,N_14468);
xor U19091 (N_19091,N_14488,N_12237);
nand U19092 (N_19092,N_12251,N_14734);
nor U19093 (N_19093,N_13967,N_15903);
or U19094 (N_19094,N_13074,N_14073);
or U19095 (N_19095,N_13084,N_13364);
and U19096 (N_19096,N_13255,N_14342);
or U19097 (N_19097,N_14656,N_15776);
xnor U19098 (N_19098,N_12743,N_12363);
nand U19099 (N_19099,N_14177,N_13118);
or U19100 (N_19100,N_12850,N_14256);
or U19101 (N_19101,N_15474,N_12419);
and U19102 (N_19102,N_15967,N_12833);
nor U19103 (N_19103,N_13371,N_15053);
nand U19104 (N_19104,N_14798,N_14625);
and U19105 (N_19105,N_12304,N_14822);
nor U19106 (N_19106,N_12561,N_13213);
nand U19107 (N_19107,N_15888,N_13829);
xnor U19108 (N_19108,N_15720,N_15436);
nor U19109 (N_19109,N_12790,N_13567);
nor U19110 (N_19110,N_13228,N_12601);
nand U19111 (N_19111,N_14004,N_12386);
and U19112 (N_19112,N_15733,N_12808);
and U19113 (N_19113,N_15087,N_15009);
nand U19114 (N_19114,N_14727,N_12161);
and U19115 (N_19115,N_13092,N_14674);
xor U19116 (N_19116,N_13420,N_12535);
nand U19117 (N_19117,N_12630,N_13221);
nor U19118 (N_19118,N_13489,N_13089);
nor U19119 (N_19119,N_15748,N_14677);
and U19120 (N_19120,N_13976,N_13797);
xor U19121 (N_19121,N_12181,N_13340);
and U19122 (N_19122,N_12398,N_14221);
and U19123 (N_19123,N_12551,N_14214);
nor U19124 (N_19124,N_14783,N_15964);
or U19125 (N_19125,N_13623,N_13063);
and U19126 (N_19126,N_13714,N_15815);
or U19127 (N_19127,N_14395,N_15278);
and U19128 (N_19128,N_13500,N_14164);
or U19129 (N_19129,N_15232,N_14556);
and U19130 (N_19130,N_14584,N_14692);
nand U19131 (N_19131,N_15596,N_14932);
xnor U19132 (N_19132,N_12323,N_13336);
and U19133 (N_19133,N_15008,N_12780);
nand U19134 (N_19134,N_15112,N_13695);
nor U19135 (N_19135,N_13238,N_15246);
or U19136 (N_19136,N_14467,N_13468);
and U19137 (N_19137,N_12885,N_15726);
or U19138 (N_19138,N_15264,N_15209);
nor U19139 (N_19139,N_13773,N_13815);
xnor U19140 (N_19140,N_15250,N_15752);
nand U19141 (N_19141,N_15209,N_15936);
or U19142 (N_19142,N_13996,N_15702);
xnor U19143 (N_19143,N_12736,N_14878);
and U19144 (N_19144,N_12720,N_13577);
and U19145 (N_19145,N_12400,N_12810);
and U19146 (N_19146,N_14386,N_15105);
nand U19147 (N_19147,N_14094,N_15805);
and U19148 (N_19148,N_14468,N_13650);
or U19149 (N_19149,N_13582,N_12595);
nand U19150 (N_19150,N_15277,N_14770);
nand U19151 (N_19151,N_15384,N_15780);
or U19152 (N_19152,N_14796,N_15057);
nor U19153 (N_19153,N_15155,N_14277);
or U19154 (N_19154,N_15986,N_14628);
nand U19155 (N_19155,N_13500,N_15673);
and U19156 (N_19156,N_12347,N_13460);
xor U19157 (N_19157,N_14054,N_13084);
and U19158 (N_19158,N_14726,N_14218);
or U19159 (N_19159,N_12068,N_14919);
and U19160 (N_19160,N_14159,N_13855);
and U19161 (N_19161,N_12247,N_15507);
nor U19162 (N_19162,N_12839,N_14341);
nor U19163 (N_19163,N_13104,N_13489);
nor U19164 (N_19164,N_15529,N_15740);
xor U19165 (N_19165,N_15553,N_15619);
and U19166 (N_19166,N_12345,N_15015);
nand U19167 (N_19167,N_13081,N_12050);
nand U19168 (N_19168,N_12194,N_13678);
nor U19169 (N_19169,N_15306,N_12536);
or U19170 (N_19170,N_13468,N_15094);
or U19171 (N_19171,N_14325,N_13484);
nand U19172 (N_19172,N_15867,N_12714);
xor U19173 (N_19173,N_13997,N_14752);
and U19174 (N_19174,N_14622,N_14898);
or U19175 (N_19175,N_14240,N_13064);
nor U19176 (N_19176,N_13292,N_13341);
and U19177 (N_19177,N_15375,N_13888);
and U19178 (N_19178,N_15452,N_15141);
nor U19179 (N_19179,N_15440,N_15926);
nor U19180 (N_19180,N_15109,N_15170);
xnor U19181 (N_19181,N_12719,N_12509);
or U19182 (N_19182,N_15551,N_13732);
and U19183 (N_19183,N_15260,N_15342);
nand U19184 (N_19184,N_15742,N_14667);
nor U19185 (N_19185,N_15262,N_15218);
nand U19186 (N_19186,N_13464,N_12732);
nand U19187 (N_19187,N_15884,N_15186);
nor U19188 (N_19188,N_13887,N_13935);
and U19189 (N_19189,N_15778,N_15831);
nor U19190 (N_19190,N_14513,N_14312);
nand U19191 (N_19191,N_13947,N_14312);
nand U19192 (N_19192,N_15606,N_12311);
nor U19193 (N_19193,N_15368,N_12503);
nor U19194 (N_19194,N_12103,N_12654);
xnor U19195 (N_19195,N_14987,N_14979);
nand U19196 (N_19196,N_15278,N_13320);
and U19197 (N_19197,N_14149,N_12037);
and U19198 (N_19198,N_14035,N_15862);
nand U19199 (N_19199,N_13352,N_14523);
or U19200 (N_19200,N_13300,N_12578);
xor U19201 (N_19201,N_14188,N_12788);
xor U19202 (N_19202,N_15617,N_15563);
nor U19203 (N_19203,N_15055,N_15545);
nand U19204 (N_19204,N_12093,N_15394);
and U19205 (N_19205,N_13803,N_13060);
or U19206 (N_19206,N_14362,N_15482);
xor U19207 (N_19207,N_14462,N_15019);
nor U19208 (N_19208,N_15288,N_12051);
and U19209 (N_19209,N_15274,N_14120);
and U19210 (N_19210,N_14417,N_13033);
or U19211 (N_19211,N_15585,N_13212);
or U19212 (N_19212,N_14344,N_14524);
or U19213 (N_19213,N_13895,N_13632);
nor U19214 (N_19214,N_12119,N_13987);
or U19215 (N_19215,N_12241,N_13959);
or U19216 (N_19216,N_12539,N_14728);
or U19217 (N_19217,N_15828,N_12390);
or U19218 (N_19218,N_13040,N_13871);
or U19219 (N_19219,N_15509,N_14944);
nand U19220 (N_19220,N_14945,N_14647);
nand U19221 (N_19221,N_13866,N_14282);
and U19222 (N_19222,N_13632,N_14992);
nor U19223 (N_19223,N_14592,N_14179);
and U19224 (N_19224,N_15038,N_15706);
or U19225 (N_19225,N_13419,N_14545);
or U19226 (N_19226,N_13068,N_15191);
nor U19227 (N_19227,N_12417,N_13752);
nand U19228 (N_19228,N_12598,N_15329);
nand U19229 (N_19229,N_12535,N_12214);
nand U19230 (N_19230,N_14362,N_12506);
nor U19231 (N_19231,N_13947,N_12334);
nand U19232 (N_19232,N_12429,N_13199);
and U19233 (N_19233,N_12940,N_14974);
or U19234 (N_19234,N_12338,N_15786);
and U19235 (N_19235,N_14811,N_14519);
or U19236 (N_19236,N_14380,N_15709);
and U19237 (N_19237,N_13683,N_14016);
nor U19238 (N_19238,N_13861,N_14512);
or U19239 (N_19239,N_12638,N_12378);
xnor U19240 (N_19240,N_12609,N_13329);
or U19241 (N_19241,N_15674,N_15801);
and U19242 (N_19242,N_15557,N_14471);
nand U19243 (N_19243,N_14188,N_14836);
nand U19244 (N_19244,N_14899,N_15194);
nor U19245 (N_19245,N_12249,N_15085);
and U19246 (N_19246,N_14794,N_15071);
nor U19247 (N_19247,N_12628,N_14854);
or U19248 (N_19248,N_14878,N_13856);
or U19249 (N_19249,N_14982,N_15789);
or U19250 (N_19250,N_12690,N_14823);
or U19251 (N_19251,N_12347,N_14669);
nand U19252 (N_19252,N_14225,N_14310);
and U19253 (N_19253,N_12538,N_14062);
and U19254 (N_19254,N_13721,N_15752);
xnor U19255 (N_19255,N_14633,N_15440);
and U19256 (N_19256,N_14132,N_13808);
or U19257 (N_19257,N_14293,N_13012);
nand U19258 (N_19258,N_14087,N_13063);
nand U19259 (N_19259,N_15452,N_15254);
nor U19260 (N_19260,N_13570,N_14845);
and U19261 (N_19261,N_14022,N_13583);
or U19262 (N_19262,N_15097,N_12411);
nor U19263 (N_19263,N_14138,N_15492);
nand U19264 (N_19264,N_12218,N_12776);
and U19265 (N_19265,N_14250,N_15160);
and U19266 (N_19266,N_15952,N_14982);
or U19267 (N_19267,N_12651,N_14507);
nor U19268 (N_19268,N_13754,N_15795);
nor U19269 (N_19269,N_13774,N_15043);
and U19270 (N_19270,N_12661,N_12373);
xor U19271 (N_19271,N_13543,N_14581);
nand U19272 (N_19272,N_13463,N_15406);
nand U19273 (N_19273,N_13921,N_12334);
and U19274 (N_19274,N_14953,N_12825);
nor U19275 (N_19275,N_14988,N_13136);
or U19276 (N_19276,N_15912,N_15755);
or U19277 (N_19277,N_12689,N_14792);
nand U19278 (N_19278,N_14444,N_15212);
nand U19279 (N_19279,N_13954,N_15735);
nand U19280 (N_19280,N_13385,N_15234);
and U19281 (N_19281,N_12023,N_12339);
xor U19282 (N_19282,N_13007,N_13413);
or U19283 (N_19283,N_12250,N_12579);
nand U19284 (N_19284,N_13933,N_15273);
nand U19285 (N_19285,N_12248,N_14988);
and U19286 (N_19286,N_12579,N_13831);
or U19287 (N_19287,N_12371,N_12832);
nand U19288 (N_19288,N_13348,N_13496);
and U19289 (N_19289,N_12012,N_13437);
and U19290 (N_19290,N_15763,N_12333);
nand U19291 (N_19291,N_13918,N_13554);
or U19292 (N_19292,N_13112,N_15744);
or U19293 (N_19293,N_14766,N_12217);
xnor U19294 (N_19294,N_12731,N_13885);
xnor U19295 (N_19295,N_13799,N_15051);
and U19296 (N_19296,N_14451,N_15059);
or U19297 (N_19297,N_12872,N_14142);
or U19298 (N_19298,N_15193,N_15608);
nand U19299 (N_19299,N_15737,N_12449);
nor U19300 (N_19300,N_15193,N_15061);
or U19301 (N_19301,N_13536,N_13529);
xnor U19302 (N_19302,N_12582,N_14167);
or U19303 (N_19303,N_14960,N_12351);
or U19304 (N_19304,N_15438,N_14974);
and U19305 (N_19305,N_12790,N_12857);
or U19306 (N_19306,N_15208,N_14952);
nor U19307 (N_19307,N_12120,N_14932);
xor U19308 (N_19308,N_12295,N_12529);
nor U19309 (N_19309,N_12410,N_13170);
nand U19310 (N_19310,N_15467,N_14389);
and U19311 (N_19311,N_13281,N_13803);
and U19312 (N_19312,N_12759,N_13701);
and U19313 (N_19313,N_15348,N_15526);
and U19314 (N_19314,N_14060,N_15271);
nand U19315 (N_19315,N_15653,N_15616);
nor U19316 (N_19316,N_13938,N_13884);
nand U19317 (N_19317,N_13050,N_15439);
or U19318 (N_19318,N_15587,N_15488);
or U19319 (N_19319,N_14202,N_13149);
nand U19320 (N_19320,N_12296,N_15513);
nor U19321 (N_19321,N_12163,N_12306);
nand U19322 (N_19322,N_14753,N_14984);
or U19323 (N_19323,N_15747,N_15848);
or U19324 (N_19324,N_14998,N_12797);
xnor U19325 (N_19325,N_14041,N_12284);
and U19326 (N_19326,N_14279,N_14795);
or U19327 (N_19327,N_15534,N_13072);
nor U19328 (N_19328,N_15592,N_14179);
and U19329 (N_19329,N_14834,N_15705);
nand U19330 (N_19330,N_13107,N_13962);
nand U19331 (N_19331,N_13065,N_13363);
nand U19332 (N_19332,N_14991,N_12320);
nand U19333 (N_19333,N_13248,N_14602);
and U19334 (N_19334,N_12830,N_13734);
and U19335 (N_19335,N_12028,N_14924);
xnor U19336 (N_19336,N_12329,N_12336);
nor U19337 (N_19337,N_13168,N_12743);
nand U19338 (N_19338,N_13479,N_15298);
and U19339 (N_19339,N_15193,N_14292);
nor U19340 (N_19340,N_13487,N_12541);
and U19341 (N_19341,N_15715,N_12777);
and U19342 (N_19342,N_13016,N_12111);
nand U19343 (N_19343,N_14749,N_12647);
nor U19344 (N_19344,N_12672,N_12728);
nand U19345 (N_19345,N_13833,N_15257);
and U19346 (N_19346,N_14100,N_14924);
nand U19347 (N_19347,N_15252,N_12664);
nor U19348 (N_19348,N_12659,N_14716);
nor U19349 (N_19349,N_13980,N_12058);
nand U19350 (N_19350,N_14845,N_15265);
nor U19351 (N_19351,N_13111,N_12015);
or U19352 (N_19352,N_13168,N_13503);
nor U19353 (N_19353,N_13646,N_13479);
or U19354 (N_19354,N_15791,N_15617);
xnor U19355 (N_19355,N_12470,N_13174);
nor U19356 (N_19356,N_15379,N_12862);
nand U19357 (N_19357,N_12554,N_12491);
or U19358 (N_19358,N_13140,N_13417);
nand U19359 (N_19359,N_15124,N_13449);
and U19360 (N_19360,N_14014,N_14592);
and U19361 (N_19361,N_12118,N_14007);
nand U19362 (N_19362,N_12828,N_14078);
xnor U19363 (N_19363,N_12118,N_12840);
and U19364 (N_19364,N_14769,N_15913);
nor U19365 (N_19365,N_13578,N_14724);
nand U19366 (N_19366,N_13028,N_12869);
xnor U19367 (N_19367,N_12896,N_13895);
nor U19368 (N_19368,N_14981,N_13290);
xor U19369 (N_19369,N_15232,N_12863);
and U19370 (N_19370,N_14566,N_13040);
or U19371 (N_19371,N_13958,N_15007);
nand U19372 (N_19372,N_13625,N_13538);
and U19373 (N_19373,N_15665,N_13499);
or U19374 (N_19374,N_13134,N_14367);
nand U19375 (N_19375,N_14683,N_12693);
xnor U19376 (N_19376,N_13990,N_12538);
or U19377 (N_19377,N_13702,N_14993);
nand U19378 (N_19378,N_15248,N_15858);
xor U19379 (N_19379,N_15208,N_13464);
xor U19380 (N_19380,N_15609,N_12066);
nor U19381 (N_19381,N_12135,N_13268);
nand U19382 (N_19382,N_13548,N_15501);
or U19383 (N_19383,N_14074,N_13296);
nand U19384 (N_19384,N_12364,N_15343);
or U19385 (N_19385,N_14961,N_12667);
and U19386 (N_19386,N_13608,N_15547);
and U19387 (N_19387,N_15578,N_15505);
nor U19388 (N_19388,N_13549,N_12224);
or U19389 (N_19389,N_15650,N_15426);
nand U19390 (N_19390,N_13713,N_15692);
or U19391 (N_19391,N_15938,N_14722);
and U19392 (N_19392,N_14156,N_12696);
or U19393 (N_19393,N_13022,N_13779);
xor U19394 (N_19394,N_15208,N_15715);
or U19395 (N_19395,N_15889,N_12252);
or U19396 (N_19396,N_13438,N_12858);
nand U19397 (N_19397,N_13293,N_15250);
or U19398 (N_19398,N_15261,N_12927);
nor U19399 (N_19399,N_15680,N_13676);
nor U19400 (N_19400,N_13857,N_12499);
or U19401 (N_19401,N_15987,N_12780);
nand U19402 (N_19402,N_12967,N_15766);
xor U19403 (N_19403,N_12719,N_13023);
nor U19404 (N_19404,N_14904,N_15621);
and U19405 (N_19405,N_13376,N_14826);
nor U19406 (N_19406,N_12020,N_15787);
and U19407 (N_19407,N_13862,N_12113);
and U19408 (N_19408,N_13829,N_13901);
and U19409 (N_19409,N_14101,N_14580);
and U19410 (N_19410,N_13311,N_15566);
nand U19411 (N_19411,N_12947,N_15191);
xnor U19412 (N_19412,N_12198,N_13422);
or U19413 (N_19413,N_14180,N_15067);
and U19414 (N_19414,N_15912,N_13839);
xor U19415 (N_19415,N_15670,N_13093);
nor U19416 (N_19416,N_14331,N_15578);
or U19417 (N_19417,N_14672,N_13197);
and U19418 (N_19418,N_12068,N_12974);
nand U19419 (N_19419,N_15682,N_14447);
or U19420 (N_19420,N_14877,N_15902);
nor U19421 (N_19421,N_15115,N_12575);
nand U19422 (N_19422,N_13281,N_13672);
and U19423 (N_19423,N_12631,N_15667);
nand U19424 (N_19424,N_13044,N_13008);
nand U19425 (N_19425,N_14941,N_13123);
nor U19426 (N_19426,N_15163,N_12327);
nand U19427 (N_19427,N_14109,N_12765);
xnor U19428 (N_19428,N_13047,N_15461);
and U19429 (N_19429,N_14874,N_12004);
nor U19430 (N_19430,N_14427,N_13858);
and U19431 (N_19431,N_14426,N_14344);
or U19432 (N_19432,N_14314,N_13416);
nand U19433 (N_19433,N_12456,N_13687);
nand U19434 (N_19434,N_15268,N_15767);
or U19435 (N_19435,N_13400,N_15553);
and U19436 (N_19436,N_12659,N_15864);
or U19437 (N_19437,N_13991,N_14346);
xor U19438 (N_19438,N_13918,N_14317);
nor U19439 (N_19439,N_13629,N_15223);
and U19440 (N_19440,N_15419,N_15834);
or U19441 (N_19441,N_13196,N_12101);
nand U19442 (N_19442,N_13475,N_14603);
nand U19443 (N_19443,N_15146,N_12080);
and U19444 (N_19444,N_13252,N_14891);
and U19445 (N_19445,N_15524,N_14614);
and U19446 (N_19446,N_12546,N_14672);
nor U19447 (N_19447,N_15192,N_13724);
nand U19448 (N_19448,N_15790,N_14848);
nor U19449 (N_19449,N_15380,N_14903);
nor U19450 (N_19450,N_14370,N_14565);
nand U19451 (N_19451,N_13044,N_15998);
nor U19452 (N_19452,N_15355,N_14929);
and U19453 (N_19453,N_12574,N_12658);
nand U19454 (N_19454,N_13112,N_12767);
or U19455 (N_19455,N_14246,N_15199);
nor U19456 (N_19456,N_14135,N_12254);
or U19457 (N_19457,N_12186,N_13997);
or U19458 (N_19458,N_15423,N_14916);
or U19459 (N_19459,N_13293,N_15244);
nand U19460 (N_19460,N_13470,N_15102);
nor U19461 (N_19461,N_14858,N_14380);
xnor U19462 (N_19462,N_14638,N_13568);
nand U19463 (N_19463,N_13258,N_14259);
and U19464 (N_19464,N_15643,N_13968);
nor U19465 (N_19465,N_14263,N_13220);
and U19466 (N_19466,N_12980,N_14691);
or U19467 (N_19467,N_15439,N_14099);
nand U19468 (N_19468,N_15615,N_12634);
or U19469 (N_19469,N_15895,N_12117);
or U19470 (N_19470,N_14795,N_15018);
xnor U19471 (N_19471,N_12895,N_14078);
nand U19472 (N_19472,N_12866,N_13764);
nor U19473 (N_19473,N_14413,N_14255);
nor U19474 (N_19474,N_15108,N_12720);
or U19475 (N_19475,N_13813,N_12544);
nand U19476 (N_19476,N_12759,N_13926);
and U19477 (N_19477,N_15852,N_15578);
and U19478 (N_19478,N_12704,N_14880);
nand U19479 (N_19479,N_13759,N_13422);
and U19480 (N_19480,N_14594,N_13594);
nor U19481 (N_19481,N_13484,N_13073);
nand U19482 (N_19482,N_12280,N_13955);
and U19483 (N_19483,N_12735,N_14454);
nor U19484 (N_19484,N_13516,N_12377);
nand U19485 (N_19485,N_12165,N_14571);
nand U19486 (N_19486,N_13970,N_15514);
xor U19487 (N_19487,N_13499,N_15315);
nand U19488 (N_19488,N_12113,N_13009);
and U19489 (N_19489,N_13678,N_14333);
nand U19490 (N_19490,N_15027,N_15053);
nand U19491 (N_19491,N_13845,N_15634);
nor U19492 (N_19492,N_13513,N_14114);
nand U19493 (N_19493,N_12553,N_15505);
nand U19494 (N_19494,N_13547,N_12412);
nor U19495 (N_19495,N_12671,N_15661);
nor U19496 (N_19496,N_14299,N_15781);
nand U19497 (N_19497,N_13127,N_12144);
nor U19498 (N_19498,N_15196,N_12200);
or U19499 (N_19499,N_14688,N_12989);
or U19500 (N_19500,N_13505,N_15914);
nand U19501 (N_19501,N_14076,N_15492);
nand U19502 (N_19502,N_15123,N_15388);
or U19503 (N_19503,N_13547,N_12282);
nor U19504 (N_19504,N_15788,N_12845);
nor U19505 (N_19505,N_13915,N_12921);
and U19506 (N_19506,N_14335,N_15600);
nor U19507 (N_19507,N_13453,N_13744);
nand U19508 (N_19508,N_13171,N_14816);
nand U19509 (N_19509,N_14090,N_15192);
or U19510 (N_19510,N_12491,N_12873);
or U19511 (N_19511,N_14127,N_13629);
nand U19512 (N_19512,N_13533,N_13566);
and U19513 (N_19513,N_13804,N_15225);
xor U19514 (N_19514,N_14112,N_12083);
xor U19515 (N_19515,N_14186,N_12899);
or U19516 (N_19516,N_13592,N_12882);
xnor U19517 (N_19517,N_15698,N_15528);
nand U19518 (N_19518,N_14531,N_12819);
nor U19519 (N_19519,N_13632,N_14994);
nor U19520 (N_19520,N_15586,N_13272);
nor U19521 (N_19521,N_15576,N_13596);
and U19522 (N_19522,N_14422,N_13304);
and U19523 (N_19523,N_12966,N_14934);
nand U19524 (N_19524,N_12270,N_14197);
xnor U19525 (N_19525,N_13392,N_14924);
nor U19526 (N_19526,N_13491,N_15860);
nand U19527 (N_19527,N_15747,N_13642);
nand U19528 (N_19528,N_13547,N_12758);
or U19529 (N_19529,N_13974,N_14992);
and U19530 (N_19530,N_15672,N_15295);
and U19531 (N_19531,N_12493,N_14867);
xor U19532 (N_19532,N_14818,N_14077);
or U19533 (N_19533,N_15875,N_15770);
nor U19534 (N_19534,N_14902,N_12185);
and U19535 (N_19535,N_12893,N_14377);
and U19536 (N_19536,N_14970,N_14420);
xor U19537 (N_19537,N_13213,N_13485);
nand U19538 (N_19538,N_13393,N_12293);
nor U19539 (N_19539,N_13327,N_13811);
nand U19540 (N_19540,N_15538,N_15085);
nand U19541 (N_19541,N_15014,N_13458);
nand U19542 (N_19542,N_13411,N_13682);
or U19543 (N_19543,N_14791,N_14328);
nand U19544 (N_19544,N_15625,N_15716);
or U19545 (N_19545,N_14968,N_13216);
and U19546 (N_19546,N_13357,N_13308);
nand U19547 (N_19547,N_13108,N_12975);
nand U19548 (N_19548,N_15406,N_15107);
or U19549 (N_19549,N_14249,N_13389);
or U19550 (N_19550,N_12960,N_13763);
or U19551 (N_19551,N_13781,N_15384);
and U19552 (N_19552,N_12919,N_13070);
nand U19553 (N_19553,N_15909,N_12897);
nor U19554 (N_19554,N_13301,N_15466);
or U19555 (N_19555,N_12834,N_14002);
nand U19556 (N_19556,N_14643,N_13745);
and U19557 (N_19557,N_14243,N_12579);
nand U19558 (N_19558,N_13285,N_12343);
and U19559 (N_19559,N_13246,N_15716);
nor U19560 (N_19560,N_14721,N_14219);
and U19561 (N_19561,N_14246,N_12895);
and U19562 (N_19562,N_14726,N_14348);
or U19563 (N_19563,N_15724,N_15791);
xnor U19564 (N_19564,N_14395,N_14691);
and U19565 (N_19565,N_13321,N_13132);
nand U19566 (N_19566,N_15264,N_14839);
and U19567 (N_19567,N_15106,N_14102);
and U19568 (N_19568,N_12986,N_12461);
nor U19569 (N_19569,N_12897,N_12998);
or U19570 (N_19570,N_15047,N_13461);
nand U19571 (N_19571,N_12534,N_14213);
or U19572 (N_19572,N_15861,N_15735);
or U19573 (N_19573,N_13865,N_15123);
or U19574 (N_19574,N_12604,N_14547);
or U19575 (N_19575,N_15908,N_14715);
nand U19576 (N_19576,N_15912,N_14157);
and U19577 (N_19577,N_14516,N_15401);
nand U19578 (N_19578,N_14430,N_12559);
and U19579 (N_19579,N_15215,N_12054);
nand U19580 (N_19580,N_13999,N_13658);
xnor U19581 (N_19581,N_14301,N_15925);
nor U19582 (N_19582,N_14716,N_15090);
and U19583 (N_19583,N_13528,N_15357);
or U19584 (N_19584,N_13253,N_13696);
or U19585 (N_19585,N_14675,N_14425);
and U19586 (N_19586,N_14480,N_14377);
and U19587 (N_19587,N_14642,N_13707);
nand U19588 (N_19588,N_15072,N_13795);
and U19589 (N_19589,N_14088,N_14583);
nand U19590 (N_19590,N_12262,N_12466);
or U19591 (N_19591,N_13574,N_14997);
and U19592 (N_19592,N_12783,N_13943);
nor U19593 (N_19593,N_13503,N_15715);
nand U19594 (N_19594,N_15586,N_14131);
or U19595 (N_19595,N_12145,N_14915);
nand U19596 (N_19596,N_13898,N_12799);
nor U19597 (N_19597,N_14724,N_14377);
and U19598 (N_19598,N_15733,N_12419);
nand U19599 (N_19599,N_15703,N_12545);
nor U19600 (N_19600,N_13514,N_14402);
nand U19601 (N_19601,N_15780,N_12678);
nand U19602 (N_19602,N_13642,N_13917);
nand U19603 (N_19603,N_12233,N_13030);
nor U19604 (N_19604,N_12133,N_15912);
and U19605 (N_19605,N_14613,N_13839);
or U19606 (N_19606,N_13273,N_12539);
and U19607 (N_19607,N_15845,N_15186);
or U19608 (N_19608,N_15754,N_13054);
nor U19609 (N_19609,N_12684,N_15771);
nand U19610 (N_19610,N_13346,N_15478);
nor U19611 (N_19611,N_13126,N_15900);
nor U19612 (N_19612,N_15340,N_13974);
nand U19613 (N_19613,N_15020,N_14210);
or U19614 (N_19614,N_13225,N_13257);
nor U19615 (N_19615,N_12313,N_13234);
xnor U19616 (N_19616,N_15709,N_13704);
nand U19617 (N_19617,N_12981,N_14013);
and U19618 (N_19618,N_14548,N_15784);
and U19619 (N_19619,N_12965,N_13055);
nand U19620 (N_19620,N_12199,N_15259);
or U19621 (N_19621,N_13889,N_13695);
and U19622 (N_19622,N_13255,N_15743);
or U19623 (N_19623,N_14678,N_12918);
nor U19624 (N_19624,N_15595,N_12406);
and U19625 (N_19625,N_12987,N_15938);
nand U19626 (N_19626,N_12307,N_12530);
and U19627 (N_19627,N_15463,N_15170);
and U19628 (N_19628,N_12229,N_15817);
or U19629 (N_19629,N_14718,N_13185);
and U19630 (N_19630,N_14119,N_15710);
or U19631 (N_19631,N_14235,N_14024);
or U19632 (N_19632,N_13622,N_15750);
nand U19633 (N_19633,N_12057,N_13472);
and U19634 (N_19634,N_14230,N_15445);
or U19635 (N_19635,N_12940,N_12233);
nand U19636 (N_19636,N_14405,N_13770);
and U19637 (N_19637,N_14188,N_13045);
or U19638 (N_19638,N_13303,N_13881);
nor U19639 (N_19639,N_12945,N_15407);
nand U19640 (N_19640,N_13557,N_12108);
or U19641 (N_19641,N_12943,N_14215);
or U19642 (N_19642,N_12924,N_14802);
nor U19643 (N_19643,N_14158,N_15161);
nor U19644 (N_19644,N_13112,N_12566);
and U19645 (N_19645,N_13063,N_14312);
nand U19646 (N_19646,N_14523,N_15361);
nand U19647 (N_19647,N_13167,N_12420);
or U19648 (N_19648,N_15065,N_14098);
and U19649 (N_19649,N_12863,N_12440);
nor U19650 (N_19650,N_14416,N_14571);
or U19651 (N_19651,N_12904,N_14684);
nor U19652 (N_19652,N_14034,N_13057);
nor U19653 (N_19653,N_13386,N_15546);
nor U19654 (N_19654,N_15569,N_13839);
and U19655 (N_19655,N_14631,N_15034);
or U19656 (N_19656,N_13305,N_15174);
nor U19657 (N_19657,N_14641,N_14136);
and U19658 (N_19658,N_13282,N_12036);
and U19659 (N_19659,N_12658,N_13235);
and U19660 (N_19660,N_14803,N_12166);
and U19661 (N_19661,N_13501,N_13201);
nor U19662 (N_19662,N_13421,N_14413);
or U19663 (N_19663,N_15656,N_14954);
nor U19664 (N_19664,N_13337,N_15349);
and U19665 (N_19665,N_12867,N_14982);
and U19666 (N_19666,N_14565,N_12422);
or U19667 (N_19667,N_13435,N_12847);
nand U19668 (N_19668,N_15862,N_15823);
and U19669 (N_19669,N_13018,N_15190);
and U19670 (N_19670,N_12385,N_15655);
xor U19671 (N_19671,N_13526,N_15801);
xnor U19672 (N_19672,N_13083,N_12854);
and U19673 (N_19673,N_13593,N_15715);
or U19674 (N_19674,N_15452,N_12906);
and U19675 (N_19675,N_15863,N_15318);
xnor U19676 (N_19676,N_13676,N_13115);
xnor U19677 (N_19677,N_14244,N_15365);
nor U19678 (N_19678,N_14853,N_14771);
and U19679 (N_19679,N_15052,N_13645);
nor U19680 (N_19680,N_15952,N_13146);
nor U19681 (N_19681,N_14430,N_13801);
nor U19682 (N_19682,N_14418,N_14368);
nand U19683 (N_19683,N_13346,N_13635);
or U19684 (N_19684,N_12120,N_15268);
or U19685 (N_19685,N_12824,N_13656);
nand U19686 (N_19686,N_15282,N_13323);
nor U19687 (N_19687,N_12269,N_14366);
or U19688 (N_19688,N_13685,N_14507);
or U19689 (N_19689,N_15467,N_15798);
or U19690 (N_19690,N_13599,N_15888);
nand U19691 (N_19691,N_13566,N_14133);
and U19692 (N_19692,N_13819,N_12510);
nand U19693 (N_19693,N_15430,N_13972);
and U19694 (N_19694,N_15592,N_13750);
xor U19695 (N_19695,N_13214,N_14731);
nor U19696 (N_19696,N_15456,N_12314);
nand U19697 (N_19697,N_15976,N_12911);
or U19698 (N_19698,N_14943,N_14276);
nor U19699 (N_19699,N_15762,N_14167);
or U19700 (N_19700,N_15366,N_14972);
and U19701 (N_19701,N_15022,N_12075);
nor U19702 (N_19702,N_15832,N_13500);
or U19703 (N_19703,N_15685,N_15335);
nand U19704 (N_19704,N_13110,N_15655);
or U19705 (N_19705,N_14824,N_14766);
nor U19706 (N_19706,N_13829,N_15886);
or U19707 (N_19707,N_13074,N_13473);
nor U19708 (N_19708,N_15291,N_14698);
or U19709 (N_19709,N_14034,N_14111);
or U19710 (N_19710,N_13717,N_13551);
nand U19711 (N_19711,N_13229,N_14359);
xor U19712 (N_19712,N_15934,N_12848);
nor U19713 (N_19713,N_13970,N_12292);
or U19714 (N_19714,N_15575,N_13038);
and U19715 (N_19715,N_14347,N_12993);
nor U19716 (N_19716,N_14266,N_13655);
xor U19717 (N_19717,N_13238,N_13552);
nor U19718 (N_19718,N_12793,N_12701);
or U19719 (N_19719,N_12402,N_12887);
and U19720 (N_19720,N_12887,N_15912);
nand U19721 (N_19721,N_12102,N_14375);
or U19722 (N_19722,N_15055,N_13225);
or U19723 (N_19723,N_13551,N_12808);
xnor U19724 (N_19724,N_12915,N_12930);
and U19725 (N_19725,N_15630,N_12976);
nand U19726 (N_19726,N_15497,N_13498);
or U19727 (N_19727,N_13422,N_15039);
xnor U19728 (N_19728,N_12456,N_14820);
nor U19729 (N_19729,N_14473,N_15730);
and U19730 (N_19730,N_15833,N_14199);
or U19731 (N_19731,N_12978,N_12170);
or U19732 (N_19732,N_13721,N_15183);
nor U19733 (N_19733,N_15577,N_15177);
nand U19734 (N_19734,N_12454,N_12138);
nand U19735 (N_19735,N_14311,N_13423);
or U19736 (N_19736,N_14319,N_13715);
xor U19737 (N_19737,N_12066,N_12456);
and U19738 (N_19738,N_13408,N_13801);
nand U19739 (N_19739,N_15101,N_14305);
nand U19740 (N_19740,N_15684,N_13742);
nand U19741 (N_19741,N_14433,N_14630);
nand U19742 (N_19742,N_15213,N_12791);
and U19743 (N_19743,N_14252,N_13734);
and U19744 (N_19744,N_15233,N_13924);
nor U19745 (N_19745,N_15692,N_15009);
and U19746 (N_19746,N_12395,N_15122);
nand U19747 (N_19747,N_12935,N_15691);
xnor U19748 (N_19748,N_13380,N_14085);
and U19749 (N_19749,N_13808,N_14849);
nor U19750 (N_19750,N_15643,N_12887);
and U19751 (N_19751,N_15220,N_14591);
nand U19752 (N_19752,N_14865,N_13574);
nand U19753 (N_19753,N_14847,N_15877);
and U19754 (N_19754,N_13384,N_13269);
nor U19755 (N_19755,N_13630,N_15906);
or U19756 (N_19756,N_14819,N_15910);
xnor U19757 (N_19757,N_12627,N_15051);
and U19758 (N_19758,N_12556,N_12027);
nor U19759 (N_19759,N_14954,N_13909);
nor U19760 (N_19760,N_12807,N_15633);
or U19761 (N_19761,N_13457,N_15884);
nand U19762 (N_19762,N_15142,N_13211);
nand U19763 (N_19763,N_12919,N_13190);
and U19764 (N_19764,N_15823,N_15054);
or U19765 (N_19765,N_15697,N_12789);
and U19766 (N_19766,N_14725,N_15852);
or U19767 (N_19767,N_13198,N_14416);
and U19768 (N_19768,N_13771,N_12236);
or U19769 (N_19769,N_13521,N_12909);
nor U19770 (N_19770,N_12584,N_15658);
nor U19771 (N_19771,N_12116,N_14352);
nand U19772 (N_19772,N_13898,N_12746);
xor U19773 (N_19773,N_14745,N_13141);
nand U19774 (N_19774,N_15465,N_12282);
nor U19775 (N_19775,N_13268,N_13063);
xnor U19776 (N_19776,N_12605,N_14945);
or U19777 (N_19777,N_15547,N_15758);
or U19778 (N_19778,N_13083,N_14749);
or U19779 (N_19779,N_13437,N_15989);
or U19780 (N_19780,N_15228,N_13843);
nand U19781 (N_19781,N_13099,N_12408);
xnor U19782 (N_19782,N_15524,N_12171);
and U19783 (N_19783,N_14692,N_15154);
nand U19784 (N_19784,N_14749,N_13005);
or U19785 (N_19785,N_14879,N_15461);
or U19786 (N_19786,N_12093,N_13813);
nand U19787 (N_19787,N_12045,N_15890);
nor U19788 (N_19788,N_14759,N_15103);
nand U19789 (N_19789,N_15326,N_13451);
nand U19790 (N_19790,N_15663,N_14017);
nand U19791 (N_19791,N_15430,N_15406);
or U19792 (N_19792,N_12416,N_12796);
nand U19793 (N_19793,N_15088,N_13246);
or U19794 (N_19794,N_15663,N_15521);
and U19795 (N_19795,N_14462,N_15432);
nor U19796 (N_19796,N_13378,N_12450);
nor U19797 (N_19797,N_13925,N_14453);
and U19798 (N_19798,N_15615,N_15389);
and U19799 (N_19799,N_13273,N_12425);
and U19800 (N_19800,N_14338,N_15396);
or U19801 (N_19801,N_13418,N_14983);
nor U19802 (N_19802,N_14406,N_13900);
nand U19803 (N_19803,N_13951,N_15579);
and U19804 (N_19804,N_13664,N_15302);
nand U19805 (N_19805,N_15505,N_12253);
nand U19806 (N_19806,N_15892,N_15039);
or U19807 (N_19807,N_14294,N_15903);
nor U19808 (N_19808,N_14055,N_13679);
and U19809 (N_19809,N_13051,N_13544);
xor U19810 (N_19810,N_12153,N_14173);
or U19811 (N_19811,N_12104,N_13786);
or U19812 (N_19812,N_14038,N_12666);
and U19813 (N_19813,N_13109,N_12130);
nor U19814 (N_19814,N_15659,N_12946);
nand U19815 (N_19815,N_14214,N_13605);
and U19816 (N_19816,N_12422,N_15124);
and U19817 (N_19817,N_15005,N_15022);
nor U19818 (N_19818,N_12362,N_12428);
nand U19819 (N_19819,N_13742,N_14902);
and U19820 (N_19820,N_15809,N_13747);
nor U19821 (N_19821,N_14626,N_12268);
and U19822 (N_19822,N_15474,N_12779);
and U19823 (N_19823,N_12572,N_14204);
xnor U19824 (N_19824,N_12331,N_15537);
or U19825 (N_19825,N_14073,N_13420);
or U19826 (N_19826,N_12778,N_12481);
or U19827 (N_19827,N_14098,N_12074);
or U19828 (N_19828,N_13752,N_15830);
and U19829 (N_19829,N_12753,N_12926);
nor U19830 (N_19830,N_12986,N_13659);
nand U19831 (N_19831,N_13697,N_14971);
and U19832 (N_19832,N_13401,N_14716);
and U19833 (N_19833,N_13486,N_12241);
nor U19834 (N_19834,N_13795,N_13758);
nor U19835 (N_19835,N_14021,N_13469);
or U19836 (N_19836,N_12773,N_13758);
nand U19837 (N_19837,N_12910,N_15496);
nand U19838 (N_19838,N_12788,N_13697);
and U19839 (N_19839,N_14593,N_15093);
or U19840 (N_19840,N_15597,N_13486);
and U19841 (N_19841,N_12313,N_15289);
and U19842 (N_19842,N_15564,N_13376);
nand U19843 (N_19843,N_13496,N_14661);
nand U19844 (N_19844,N_15052,N_15491);
nand U19845 (N_19845,N_12715,N_14818);
and U19846 (N_19846,N_12662,N_12112);
or U19847 (N_19847,N_13954,N_14785);
and U19848 (N_19848,N_13063,N_13743);
xor U19849 (N_19849,N_14775,N_12395);
and U19850 (N_19850,N_12828,N_15367);
and U19851 (N_19851,N_13535,N_15078);
and U19852 (N_19852,N_15506,N_12953);
nor U19853 (N_19853,N_13616,N_14811);
nor U19854 (N_19854,N_12226,N_14123);
or U19855 (N_19855,N_14842,N_14626);
xnor U19856 (N_19856,N_13226,N_13818);
and U19857 (N_19857,N_14289,N_15709);
or U19858 (N_19858,N_14057,N_14845);
nor U19859 (N_19859,N_14154,N_15196);
or U19860 (N_19860,N_13595,N_12107);
or U19861 (N_19861,N_13233,N_12455);
nand U19862 (N_19862,N_12800,N_12631);
nand U19863 (N_19863,N_12097,N_12162);
or U19864 (N_19864,N_12763,N_13032);
or U19865 (N_19865,N_14213,N_14265);
xor U19866 (N_19866,N_14339,N_14269);
nand U19867 (N_19867,N_13134,N_12512);
nor U19868 (N_19868,N_12287,N_15307);
and U19869 (N_19869,N_14311,N_13011);
or U19870 (N_19870,N_14945,N_14607);
or U19871 (N_19871,N_12489,N_14969);
and U19872 (N_19872,N_13024,N_15290);
or U19873 (N_19873,N_15656,N_14774);
nor U19874 (N_19874,N_14235,N_13841);
and U19875 (N_19875,N_13420,N_13739);
nand U19876 (N_19876,N_13294,N_12805);
nand U19877 (N_19877,N_13233,N_15023);
nor U19878 (N_19878,N_12522,N_14332);
xnor U19879 (N_19879,N_12648,N_13905);
and U19880 (N_19880,N_15835,N_12375);
nand U19881 (N_19881,N_13235,N_12641);
xor U19882 (N_19882,N_13926,N_14410);
or U19883 (N_19883,N_13498,N_14884);
xor U19884 (N_19884,N_12420,N_13475);
nand U19885 (N_19885,N_15858,N_12956);
nand U19886 (N_19886,N_13946,N_12611);
and U19887 (N_19887,N_14372,N_15195);
nand U19888 (N_19888,N_15418,N_15505);
and U19889 (N_19889,N_15747,N_13169);
and U19890 (N_19890,N_13813,N_14294);
and U19891 (N_19891,N_13627,N_15374);
xor U19892 (N_19892,N_12523,N_13669);
nand U19893 (N_19893,N_15674,N_15013);
or U19894 (N_19894,N_15882,N_14524);
and U19895 (N_19895,N_14776,N_15025);
nand U19896 (N_19896,N_14542,N_14938);
nor U19897 (N_19897,N_14701,N_13168);
and U19898 (N_19898,N_13768,N_14403);
or U19899 (N_19899,N_14695,N_12777);
nor U19900 (N_19900,N_13037,N_15568);
or U19901 (N_19901,N_14102,N_12315);
and U19902 (N_19902,N_14170,N_12957);
and U19903 (N_19903,N_12496,N_15329);
or U19904 (N_19904,N_13629,N_12938);
xor U19905 (N_19905,N_15741,N_12896);
xnor U19906 (N_19906,N_12637,N_12505);
or U19907 (N_19907,N_13491,N_15800);
xnor U19908 (N_19908,N_14188,N_15118);
and U19909 (N_19909,N_13424,N_13118);
nand U19910 (N_19910,N_14467,N_15101);
nor U19911 (N_19911,N_15110,N_14881);
nand U19912 (N_19912,N_12091,N_15208);
and U19913 (N_19913,N_13918,N_15663);
nor U19914 (N_19914,N_15581,N_13406);
or U19915 (N_19915,N_14031,N_15409);
nand U19916 (N_19916,N_12798,N_13188);
and U19917 (N_19917,N_12247,N_14243);
nand U19918 (N_19918,N_13752,N_14006);
or U19919 (N_19919,N_12846,N_15737);
and U19920 (N_19920,N_13385,N_12794);
nand U19921 (N_19921,N_13842,N_13771);
nand U19922 (N_19922,N_15015,N_12600);
nand U19923 (N_19923,N_14338,N_12204);
nand U19924 (N_19924,N_12844,N_15927);
nand U19925 (N_19925,N_14238,N_15098);
nor U19926 (N_19926,N_14176,N_15253);
nand U19927 (N_19927,N_15595,N_12850);
nand U19928 (N_19928,N_14804,N_13965);
and U19929 (N_19929,N_15551,N_14595);
nor U19930 (N_19930,N_13591,N_13664);
nor U19931 (N_19931,N_15292,N_15493);
nand U19932 (N_19932,N_15811,N_12719);
nand U19933 (N_19933,N_13210,N_13377);
or U19934 (N_19934,N_12889,N_12862);
nand U19935 (N_19935,N_14146,N_15228);
nand U19936 (N_19936,N_13014,N_15847);
nand U19937 (N_19937,N_13350,N_15960);
nor U19938 (N_19938,N_12980,N_14225);
nor U19939 (N_19939,N_13086,N_14005);
nand U19940 (N_19940,N_12853,N_12128);
nand U19941 (N_19941,N_15459,N_14970);
xor U19942 (N_19942,N_15175,N_13685);
and U19943 (N_19943,N_12454,N_14249);
or U19944 (N_19944,N_14208,N_15640);
or U19945 (N_19945,N_15484,N_14841);
and U19946 (N_19946,N_15367,N_12098);
or U19947 (N_19947,N_14288,N_13793);
nand U19948 (N_19948,N_12562,N_12339);
or U19949 (N_19949,N_13127,N_13988);
and U19950 (N_19950,N_14667,N_14783);
or U19951 (N_19951,N_14079,N_13331);
nor U19952 (N_19952,N_14632,N_13992);
or U19953 (N_19953,N_13693,N_14659);
or U19954 (N_19954,N_13075,N_14856);
xnor U19955 (N_19955,N_14943,N_14137);
nand U19956 (N_19956,N_14602,N_13016);
and U19957 (N_19957,N_14150,N_15689);
nor U19958 (N_19958,N_13543,N_15677);
or U19959 (N_19959,N_15003,N_13010);
nor U19960 (N_19960,N_15656,N_12589);
nor U19961 (N_19961,N_13259,N_14927);
xor U19962 (N_19962,N_12383,N_14882);
nor U19963 (N_19963,N_14219,N_14808);
and U19964 (N_19964,N_14135,N_12857);
nor U19965 (N_19965,N_13065,N_15040);
nand U19966 (N_19966,N_12762,N_14720);
xnor U19967 (N_19967,N_15751,N_14445);
and U19968 (N_19968,N_15718,N_15638);
or U19969 (N_19969,N_15800,N_13923);
nand U19970 (N_19970,N_12661,N_15672);
and U19971 (N_19971,N_12798,N_15375);
nor U19972 (N_19972,N_13845,N_14462);
and U19973 (N_19973,N_15093,N_14010);
nand U19974 (N_19974,N_12500,N_13411);
nand U19975 (N_19975,N_12155,N_13814);
nor U19976 (N_19976,N_12779,N_14384);
or U19977 (N_19977,N_13081,N_12859);
or U19978 (N_19978,N_13157,N_15795);
nand U19979 (N_19979,N_15954,N_15776);
and U19980 (N_19980,N_13211,N_12987);
nor U19981 (N_19981,N_13206,N_14408);
or U19982 (N_19982,N_14053,N_13954);
nand U19983 (N_19983,N_15212,N_14998);
and U19984 (N_19984,N_13436,N_13293);
or U19985 (N_19985,N_15838,N_15663);
or U19986 (N_19986,N_14896,N_13768);
nand U19987 (N_19987,N_14912,N_13396);
and U19988 (N_19988,N_12594,N_15077);
and U19989 (N_19989,N_14554,N_15533);
xnor U19990 (N_19990,N_12057,N_15106);
xor U19991 (N_19991,N_13529,N_14849);
and U19992 (N_19992,N_12352,N_15495);
and U19993 (N_19993,N_14042,N_15034);
and U19994 (N_19994,N_15114,N_13709);
nor U19995 (N_19995,N_13000,N_15317);
and U19996 (N_19996,N_14645,N_13576);
xor U19997 (N_19997,N_13750,N_12203);
nor U19998 (N_19998,N_12512,N_13562);
or U19999 (N_19999,N_13076,N_12412);
and UO_0 (O_0,N_16705,N_17158);
and UO_1 (O_1,N_17409,N_18572);
nand UO_2 (O_2,N_16691,N_16876);
nand UO_3 (O_3,N_16805,N_19633);
nand UO_4 (O_4,N_19737,N_17199);
and UO_5 (O_5,N_18850,N_17735);
nand UO_6 (O_6,N_17713,N_17228);
xnor UO_7 (O_7,N_16143,N_18989);
and UO_8 (O_8,N_17476,N_18442);
or UO_9 (O_9,N_17705,N_16409);
and UO_10 (O_10,N_18844,N_17312);
nor UO_11 (O_11,N_16325,N_16600);
or UO_12 (O_12,N_16245,N_16071);
nor UO_13 (O_13,N_17696,N_19078);
nand UO_14 (O_14,N_19261,N_16759);
xnor UO_15 (O_15,N_16666,N_17806);
nand UO_16 (O_16,N_19543,N_17103);
or UO_17 (O_17,N_19129,N_19949);
and UO_18 (O_18,N_19370,N_19808);
or UO_19 (O_19,N_18041,N_17813);
nand UO_20 (O_20,N_16768,N_19158);
nor UO_21 (O_21,N_18072,N_16144);
or UO_22 (O_22,N_16178,N_19740);
or UO_23 (O_23,N_17542,N_17336);
xnor UO_24 (O_24,N_19312,N_16998);
or UO_25 (O_25,N_17453,N_18998);
nor UO_26 (O_26,N_16785,N_19752);
nor UO_27 (O_27,N_16947,N_16561);
or UO_28 (O_28,N_18305,N_19528);
and UO_29 (O_29,N_19564,N_18722);
nand UO_30 (O_30,N_16251,N_16447);
or UO_31 (O_31,N_18524,N_17485);
nand UO_32 (O_32,N_18925,N_16311);
nand UO_33 (O_33,N_17610,N_19332);
xor UO_34 (O_34,N_17971,N_17405);
nor UO_35 (O_35,N_19552,N_19235);
and UO_36 (O_36,N_18943,N_16990);
or UO_37 (O_37,N_18431,N_18045);
and UO_38 (O_38,N_16308,N_16858);
and UO_39 (O_39,N_17845,N_19276);
xnor UO_40 (O_40,N_17297,N_17611);
nand UO_41 (O_41,N_16132,N_16243);
nand UO_42 (O_42,N_16033,N_16031);
nor UO_43 (O_43,N_16389,N_18293);
or UO_44 (O_44,N_17464,N_16174);
xor UO_45 (O_45,N_19239,N_18455);
and UO_46 (O_46,N_19353,N_17354);
nand UO_47 (O_47,N_17757,N_16271);
or UO_48 (O_48,N_17767,N_16266);
or UO_49 (O_49,N_17896,N_17750);
or UO_50 (O_50,N_19594,N_17461);
nor UO_51 (O_51,N_19833,N_18176);
nand UO_52 (O_52,N_17765,N_18854);
and UO_53 (O_53,N_16503,N_17707);
xnor UO_54 (O_54,N_18508,N_16092);
and UO_55 (O_55,N_18742,N_16514);
or UO_56 (O_56,N_17247,N_18997);
nor UO_57 (O_57,N_18818,N_16029);
and UO_58 (O_58,N_19970,N_18785);
or UO_59 (O_59,N_18438,N_19950);
nor UO_60 (O_60,N_19400,N_16761);
or UO_61 (O_61,N_16475,N_19605);
nand UO_62 (O_62,N_19124,N_16813);
xnor UO_63 (O_63,N_17715,N_18758);
nand UO_64 (O_64,N_19601,N_17535);
nand UO_65 (O_65,N_17057,N_18714);
or UO_66 (O_66,N_18685,N_16487);
or UO_67 (O_67,N_16939,N_17974);
nand UO_68 (O_68,N_19100,N_16778);
nor UO_69 (O_69,N_19316,N_16655);
nand UO_70 (O_70,N_18081,N_16852);
nand UO_71 (O_71,N_17601,N_16450);
or UO_72 (O_72,N_19579,N_16110);
and UO_73 (O_73,N_18095,N_18027);
nand UO_74 (O_74,N_19850,N_17788);
nor UO_75 (O_75,N_16402,N_18213);
nor UO_76 (O_76,N_16648,N_16495);
nor UO_77 (O_77,N_17808,N_16142);
nand UO_78 (O_78,N_16793,N_17321);
nand UO_79 (O_79,N_17555,N_19367);
and UO_80 (O_80,N_19548,N_18398);
nand UO_81 (O_81,N_18511,N_18316);
xnor UO_82 (O_82,N_16963,N_17142);
nand UO_83 (O_83,N_18744,N_16378);
nor UO_84 (O_84,N_19018,N_16592);
or UO_85 (O_85,N_19466,N_19984);
or UO_86 (O_86,N_18001,N_17731);
and UO_87 (O_87,N_18986,N_17078);
nand UO_88 (O_88,N_16364,N_16969);
and UO_89 (O_89,N_17474,N_17167);
or UO_90 (O_90,N_18253,N_17112);
nor UO_91 (O_91,N_19913,N_19785);
or UO_92 (O_92,N_19348,N_19423);
nor UO_93 (O_93,N_16150,N_17108);
xor UO_94 (O_94,N_19039,N_16777);
nand UO_95 (O_95,N_17445,N_18167);
nor UO_96 (O_96,N_19569,N_19803);
and UO_97 (O_97,N_19773,N_18912);
or UO_98 (O_98,N_18236,N_18324);
or UO_99 (O_99,N_19067,N_17101);
nand UO_100 (O_100,N_19396,N_19005);
or UO_101 (O_101,N_19098,N_18955);
nor UO_102 (O_102,N_18183,N_16304);
nand UO_103 (O_103,N_17334,N_18050);
or UO_104 (O_104,N_19643,N_19211);
nand UO_105 (O_105,N_19150,N_18494);
nand UO_106 (O_106,N_16638,N_16258);
xor UO_107 (O_107,N_16326,N_16548);
xnor UO_108 (O_108,N_19991,N_19973);
nor UO_109 (O_109,N_17121,N_19728);
or UO_110 (O_110,N_16256,N_17604);
xnor UO_111 (O_111,N_16718,N_16436);
nor UO_112 (O_112,N_18344,N_19198);
nand UO_113 (O_113,N_17457,N_16301);
nor UO_114 (O_114,N_16595,N_17643);
nor UO_115 (O_115,N_17728,N_16373);
and UO_116 (O_116,N_19856,N_19020);
nor UO_117 (O_117,N_18876,N_19186);
and UO_118 (O_118,N_19929,N_18839);
and UO_119 (O_119,N_17599,N_16698);
and UO_120 (O_120,N_19416,N_16264);
or UO_121 (O_121,N_18142,N_19671);
xnor UO_122 (O_122,N_19160,N_16797);
or UO_123 (O_123,N_19016,N_18161);
nor UO_124 (O_124,N_18110,N_19194);
nand UO_125 (O_125,N_17248,N_16242);
nand UO_126 (O_126,N_18583,N_17390);
nor UO_127 (O_127,N_18127,N_18520);
or UO_128 (O_128,N_17651,N_17920);
nor UO_129 (O_129,N_18152,N_16690);
nor UO_130 (O_130,N_18238,N_18426);
nor UO_131 (O_131,N_18547,N_16467);
and UO_132 (O_132,N_17137,N_17937);
nor UO_133 (O_133,N_17202,N_18332);
nor UO_134 (O_134,N_18975,N_18191);
or UO_135 (O_135,N_16111,N_18138);
xor UO_136 (O_136,N_18732,N_18527);
and UO_137 (O_137,N_17968,N_18929);
nand UO_138 (O_138,N_18846,N_16629);
xnor UO_139 (O_139,N_16088,N_16729);
and UO_140 (O_140,N_18469,N_18739);
or UO_141 (O_141,N_16396,N_17590);
and UO_142 (O_142,N_18171,N_17349);
nand UO_143 (O_143,N_18761,N_17055);
and UO_144 (O_144,N_17682,N_18674);
and UO_145 (O_145,N_18342,N_16683);
or UO_146 (O_146,N_19527,N_19575);
nand UO_147 (O_147,N_19406,N_16814);
or UO_148 (O_148,N_19443,N_18004);
nor UO_149 (O_149,N_17416,N_16321);
nor UO_150 (O_150,N_17675,N_19924);
xnor UO_151 (O_151,N_18054,N_18919);
nand UO_152 (O_152,N_18406,N_16250);
or UO_153 (O_153,N_19074,N_16199);
nand UO_154 (O_154,N_16987,N_16585);
and UO_155 (O_155,N_16593,N_17560);
nor UO_156 (O_156,N_17553,N_17825);
and UO_157 (O_157,N_18239,N_16244);
or UO_158 (O_158,N_18057,N_16730);
nand UO_159 (O_159,N_16073,N_17428);
or UO_160 (O_160,N_18498,N_17411);
nor UO_161 (O_161,N_18403,N_19557);
nor UO_162 (O_162,N_17591,N_16306);
or UO_163 (O_163,N_17098,N_18179);
nor UO_164 (O_164,N_16614,N_17570);
nor UO_165 (O_165,N_19111,N_16589);
or UO_166 (O_166,N_18907,N_16290);
nand UO_167 (O_167,N_16933,N_18680);
nor UO_168 (O_168,N_16567,N_19214);
nor UO_169 (O_169,N_18084,N_17410);
nor UO_170 (O_170,N_19137,N_19901);
and UO_171 (O_171,N_19843,N_17885);
nand UO_172 (O_172,N_17626,N_19931);
nor UO_173 (O_173,N_18856,N_19588);
and UO_174 (O_174,N_17949,N_16541);
and UO_175 (O_175,N_18783,N_17091);
nor UO_176 (O_176,N_19884,N_19299);
nor UO_177 (O_177,N_18805,N_19590);
xnor UO_178 (O_178,N_18189,N_19816);
nor UO_179 (O_179,N_16607,N_16889);
or UO_180 (O_180,N_18329,N_19278);
nor UO_181 (O_181,N_17725,N_18617);
or UO_182 (O_182,N_17332,N_19864);
nor UO_183 (O_183,N_19921,N_18078);
nand UO_184 (O_184,N_19897,N_16848);
nor UO_185 (O_185,N_16238,N_17779);
nor UO_186 (O_186,N_17880,N_18800);
or UO_187 (O_187,N_18321,N_16726);
and UO_188 (O_188,N_18297,N_19600);
nand UO_189 (O_189,N_19867,N_19758);
or UO_190 (O_190,N_19483,N_19424);
xnor UO_191 (O_191,N_18291,N_16625);
or UO_192 (O_192,N_16387,N_16932);
nor UO_193 (O_193,N_18088,N_17690);
nor UO_194 (O_194,N_16343,N_17217);
and UO_195 (O_195,N_16505,N_18210);
nor UO_196 (O_196,N_18985,N_19701);
nor UO_197 (O_197,N_17391,N_17567);
nor UO_198 (O_198,N_19486,N_19070);
nor UO_199 (O_199,N_18574,N_17619);
or UO_200 (O_200,N_16123,N_19553);
nor UO_201 (O_201,N_19065,N_17181);
nor UO_202 (O_202,N_18266,N_19749);
nor UO_203 (O_203,N_17344,N_18683);
and UO_204 (O_204,N_18735,N_18120);
and UO_205 (O_205,N_16298,N_19189);
nand UO_206 (O_206,N_19980,N_16803);
nand UO_207 (O_207,N_17618,N_19978);
and UO_208 (O_208,N_19667,N_16757);
and UO_209 (O_209,N_16135,N_19031);
nand UO_210 (O_210,N_18273,N_19322);
or UO_211 (O_211,N_19906,N_17315);
xnor UO_212 (O_212,N_18162,N_16860);
nand UO_213 (O_213,N_17685,N_17339);
and UO_214 (O_214,N_16509,N_18639);
or UO_215 (O_215,N_18383,N_17669);
or UO_216 (O_216,N_19591,N_16623);
and UO_217 (O_217,N_18112,N_19300);
or UO_218 (O_218,N_18651,N_16010);
nand UO_219 (O_219,N_16553,N_18390);
nand UO_220 (O_220,N_16292,N_17270);
nor UO_221 (O_221,N_16671,N_19414);
and UO_222 (O_222,N_19102,N_19355);
nor UO_223 (O_223,N_17094,N_16072);
and UO_224 (O_224,N_19580,N_18654);
or UO_225 (O_225,N_18663,N_19159);
and UO_226 (O_226,N_19644,N_16380);
and UO_227 (O_227,N_16583,N_19654);
nand UO_228 (O_228,N_16480,N_18462);
and UO_229 (O_229,N_19987,N_16740);
xnor UO_230 (O_230,N_17446,N_17901);
nand UO_231 (O_231,N_16197,N_17141);
nor UO_232 (O_232,N_16315,N_18423);
or UO_233 (O_233,N_16949,N_18312);
and UO_234 (O_234,N_19257,N_19148);
nand UO_235 (O_235,N_19217,N_18252);
and UO_236 (O_236,N_19948,N_16191);
nand UO_237 (O_237,N_19138,N_19730);
or UO_238 (O_238,N_17293,N_17117);
nor UO_239 (O_239,N_17206,N_17481);
xor UO_240 (O_240,N_18757,N_18107);
or UO_241 (O_241,N_18275,N_17291);
nor UO_242 (O_242,N_17089,N_17663);
nand UO_243 (O_243,N_17631,N_19969);
nand UO_244 (O_244,N_16171,N_19676);
xor UO_245 (O_245,N_18822,N_16388);
or UO_246 (O_246,N_19000,N_18377);
nand UO_247 (O_247,N_17493,N_17805);
xnor UO_248 (O_248,N_18021,N_16512);
nand UO_249 (O_249,N_17970,N_18678);
nand UO_250 (O_250,N_18348,N_16130);
nand UO_251 (O_251,N_19751,N_17525);
nor UO_252 (O_252,N_18351,N_16981);
and UO_253 (O_253,N_18550,N_16910);
and UO_254 (O_254,N_17285,N_17150);
nor UO_255 (O_255,N_19647,N_19133);
nor UO_256 (O_256,N_18477,N_18737);
xor UO_257 (O_257,N_17085,N_17828);
nand UO_258 (O_258,N_17658,N_19522);
and UO_259 (O_259,N_16064,N_17853);
or UO_260 (O_260,N_18770,N_19887);
xor UO_261 (O_261,N_16067,N_19272);
and UO_262 (O_262,N_18217,N_16265);
nand UO_263 (O_263,N_16145,N_18056);
xnor UO_264 (O_264,N_17488,N_16547);
and UO_265 (O_265,N_17062,N_18791);
nand UO_266 (O_266,N_18365,N_17869);
and UO_267 (O_267,N_19517,N_18094);
nand UO_268 (O_268,N_17956,N_18144);
nand UO_269 (O_269,N_19729,N_17165);
xnor UO_270 (O_270,N_16097,N_18801);
or UO_271 (O_271,N_18388,N_19904);
nand UO_272 (O_272,N_18151,N_19254);
or UO_273 (O_273,N_19456,N_19834);
or UO_274 (O_274,N_16838,N_17277);
xnor UO_275 (O_275,N_19255,N_17382);
and UO_276 (O_276,N_17007,N_16416);
and UO_277 (O_277,N_18020,N_18495);
xnor UO_278 (O_278,N_16140,N_18047);
or UO_279 (O_279,N_19465,N_19338);
nor UO_280 (O_280,N_16479,N_19546);
nand UO_281 (O_281,N_17575,N_17340);
or UO_282 (O_282,N_17614,N_19755);
nor UO_283 (O_283,N_19051,N_16058);
nand UO_284 (O_284,N_16517,N_17634);
nand UO_285 (O_285,N_17215,N_17388);
nor UO_286 (O_286,N_18241,N_16108);
nand UO_287 (O_287,N_18774,N_18671);
nor UO_288 (O_288,N_18540,N_17694);
nand UO_289 (O_289,N_19452,N_16383);
or UO_290 (O_290,N_17807,N_18855);
nand UO_291 (O_291,N_16115,N_16166);
and UO_292 (O_292,N_18080,N_18009);
nand UO_293 (O_293,N_16363,N_16232);
nor UO_294 (O_294,N_17208,N_16113);
xor UO_295 (O_295,N_19464,N_17637);
nor UO_296 (O_296,N_18954,N_16076);
or UO_297 (O_297,N_19380,N_16820);
and UO_298 (O_298,N_19857,N_19110);
nor UO_299 (O_299,N_17514,N_16225);
or UO_300 (O_300,N_18489,N_18734);
or UO_301 (O_301,N_19253,N_19873);
nor UO_302 (O_302,N_19567,N_16531);
nor UO_303 (O_303,N_16751,N_17664);
and UO_304 (O_304,N_17529,N_17162);
nand UO_305 (O_305,N_19865,N_19576);
nand UO_306 (O_306,N_17419,N_19462);
nor UO_307 (O_307,N_18804,N_19637);
nand UO_308 (O_308,N_19373,N_16642);
xor UO_309 (O_309,N_16737,N_18620);
nand UO_310 (O_310,N_19687,N_18870);
nand UO_311 (O_311,N_19054,N_18113);
and UO_312 (O_312,N_17284,N_16627);
nor UO_313 (O_313,N_18689,N_17099);
xor UO_314 (O_314,N_19872,N_17432);
xor UO_315 (O_315,N_18773,N_16369);
and UO_316 (O_316,N_16156,N_16557);
nor UO_317 (O_317,N_18513,N_19478);
nor UO_318 (O_318,N_19045,N_19310);
nand UO_319 (O_319,N_18279,N_16610);
xnor UO_320 (O_320,N_19750,N_17144);
nor UO_321 (O_321,N_19918,N_18308);
xor UO_322 (O_322,N_19115,N_18936);
and UO_323 (O_323,N_17819,N_17522);
nor UO_324 (O_324,N_16339,N_16755);
or UO_325 (O_325,N_18437,N_18750);
or UO_326 (O_326,N_18718,N_16438);
or UO_327 (O_327,N_17179,N_19279);
nor UO_328 (O_328,N_18802,N_17781);
xor UO_329 (O_329,N_17484,N_18432);
nand UO_330 (O_330,N_17246,N_19679);
nand UO_331 (O_331,N_19963,N_17090);
and UO_332 (O_332,N_18402,N_19571);
nor UO_333 (O_333,N_17743,N_17021);
and UO_334 (O_334,N_18143,N_19975);
and UO_335 (O_335,N_19153,N_17931);
nor UO_336 (O_336,N_18254,N_19377);
or UO_337 (O_337,N_18972,N_17596);
nor UO_338 (O_338,N_18204,N_18182);
nor UO_339 (O_339,N_18798,N_19336);
xor UO_340 (O_340,N_18341,N_19706);
or UO_341 (O_341,N_18851,N_17691);
and UO_342 (O_342,N_18769,N_19280);
xnor UO_343 (O_343,N_16764,N_16005);
nor UO_344 (O_344,N_18824,N_18130);
and UO_345 (O_345,N_16714,N_16159);
or UO_346 (O_346,N_19774,N_17362);
nand UO_347 (O_347,N_17519,N_16964);
nor UO_348 (O_348,N_17161,N_17163);
xor UO_349 (O_349,N_17938,N_18705);
and UO_350 (O_350,N_18434,N_18367);
nand UO_351 (O_351,N_18945,N_18139);
or UO_352 (O_352,N_16526,N_16370);
or UO_353 (O_353,N_17223,N_19800);
nor UO_354 (O_354,N_19034,N_17904);
or UO_355 (O_355,N_17407,N_17052);
or UO_356 (O_356,N_18096,N_18759);
or UO_357 (O_357,N_16272,N_16725);
nand UO_358 (O_358,N_18728,N_16771);
and UO_359 (O_359,N_16189,N_17787);
xnor UO_360 (O_360,N_18010,N_18267);
and UO_361 (O_361,N_17071,N_19815);
nor UO_362 (O_362,N_18160,N_19088);
and UO_363 (O_363,N_17566,N_19086);
nor UO_364 (O_364,N_16239,N_19477);
nand UO_365 (O_365,N_17274,N_19632);
nand UO_366 (O_366,N_16448,N_17492);
or UO_367 (O_367,N_19246,N_19069);
and UO_368 (O_368,N_18257,N_16839);
nor UO_369 (O_369,N_19429,N_18303);
nor UO_370 (O_370,N_17443,N_18747);
or UO_371 (O_371,N_16635,N_17255);
nand UO_372 (O_372,N_17660,N_18089);
nand UO_373 (O_373,N_16346,N_17612);
and UO_374 (O_374,N_16749,N_19083);
nand UO_375 (O_375,N_16350,N_18395);
nor UO_376 (O_376,N_16367,N_18396);
nor UO_377 (O_377,N_16566,N_19819);
xor UO_378 (O_378,N_19058,N_18227);
or UO_379 (O_379,N_19568,N_19435);
or UO_380 (O_380,N_17424,N_18011);
nor UO_381 (O_381,N_19014,N_19173);
nand UO_382 (O_382,N_16536,N_18389);
nand UO_383 (O_383,N_16282,N_16390);
or UO_384 (O_384,N_17774,N_19689);
and UO_385 (O_385,N_17871,N_19835);
nand UO_386 (O_386,N_19981,N_17360);
and UO_387 (O_387,N_17554,N_18382);
nor UO_388 (O_388,N_18033,N_16177);
or UO_389 (O_389,N_17908,N_16911);
and UO_390 (O_390,N_16921,N_19983);
nand UO_391 (O_391,N_16167,N_17292);
nand UO_392 (O_392,N_19692,N_18710);
and UO_393 (O_393,N_19945,N_17458);
and UO_394 (O_394,N_18313,N_19555);
nand UO_395 (O_395,N_16283,N_19589);
nand UO_396 (O_396,N_16784,N_19177);
xnor UO_397 (O_397,N_17517,N_18032);
and UO_398 (O_398,N_17977,N_17925);
or UO_399 (O_399,N_17744,N_19718);
nor UO_400 (O_400,N_17483,N_19028);
or UO_401 (O_401,N_18833,N_17160);
or UO_402 (O_402,N_19281,N_19955);
or UO_403 (O_403,N_17238,N_18886);
nor UO_404 (O_404,N_17965,N_17383);
nor UO_405 (O_405,N_16275,N_18368);
and UO_406 (O_406,N_17646,N_17689);
and UO_407 (O_407,N_18884,N_17303);
nor UO_408 (O_408,N_17086,N_18720);
or UO_409 (O_409,N_16670,N_19320);
nand UO_410 (O_410,N_16875,N_18772);
or UO_411 (O_411,N_19275,N_19908);
nor UO_412 (O_412,N_18662,N_17438);
or UO_413 (O_413,N_18156,N_18949);
or UO_414 (O_414,N_16418,N_16894);
and UO_415 (O_415,N_17841,N_18430);
or UO_416 (O_416,N_16327,N_19165);
and UO_417 (O_417,N_19716,N_19216);
nand UO_418 (O_418,N_16429,N_19121);
and UO_419 (O_419,N_17840,N_18128);
nor UO_420 (O_420,N_19611,N_18192);
or UO_421 (O_421,N_19182,N_19109);
or UO_422 (O_422,N_17895,N_19747);
nor UO_423 (O_423,N_18569,N_18199);
nand UO_424 (O_424,N_17550,N_18883);
nor UO_425 (O_425,N_18965,N_19721);
nor UO_426 (O_426,N_18594,N_17692);
nor UO_427 (O_427,N_17040,N_17135);
or UO_428 (O_428,N_18386,N_18061);
or UO_429 (O_429,N_18981,N_18840);
or UO_430 (O_430,N_19116,N_19412);
or UO_431 (O_431,N_17119,N_18480);
nand UO_432 (O_432,N_17156,N_18283);
nand UO_433 (O_433,N_18537,N_16020);
nor UO_434 (O_434,N_19019,N_19037);
nor UO_435 (O_435,N_17231,N_19925);
nor UO_436 (O_436,N_19351,N_19723);
and UO_437 (O_437,N_19314,N_19357);
and UO_438 (O_438,N_19459,N_16011);
or UO_439 (O_439,N_17768,N_18542);
or UO_440 (O_440,N_19744,N_19335);
or UO_441 (O_441,N_17835,N_16731);
and UO_442 (O_442,N_18519,N_18708);
and UO_443 (O_443,N_18463,N_17572);
nand UO_444 (O_444,N_16065,N_18675);
xor UO_445 (O_445,N_19087,N_19940);
and UO_446 (O_446,N_18416,N_16224);
nor UO_447 (O_447,N_17319,N_16125);
and UO_448 (O_448,N_18361,N_18871);
nor UO_449 (O_449,N_16529,N_17770);
or UO_450 (O_450,N_16781,N_19410);
and UO_451 (O_451,N_17565,N_16832);
nand UO_452 (O_452,N_18046,N_16904);
and UO_453 (O_453,N_16796,N_19989);
nand UO_454 (O_454,N_18729,N_19824);
and UO_455 (O_455,N_19610,N_17673);
or UO_456 (O_456,N_16053,N_17102);
nand UO_457 (O_457,N_18169,N_19563);
and UO_458 (O_458,N_17623,N_19577);
nor UO_459 (O_459,N_17183,N_17615);
nor UO_460 (O_460,N_19957,N_19099);
and UO_461 (O_461,N_18278,N_16034);
and UO_462 (O_462,N_19157,N_19089);
or UO_463 (O_463,N_18349,N_16825);
nand UO_464 (O_464,N_17919,N_17644);
or UO_465 (O_465,N_16030,N_19195);
nand UO_466 (O_466,N_16345,N_19467);
nand UO_467 (O_467,N_19842,N_19418);
xnor UO_468 (O_468,N_18845,N_17531);
or UO_469 (O_469,N_19821,N_17916);
or UO_470 (O_470,N_18897,N_19293);
and UO_471 (O_471,N_17816,N_19652);
nor UO_472 (O_472,N_17834,N_19670);
or UO_473 (O_473,N_17393,N_16446);
or UO_474 (O_474,N_17678,N_16334);
nor UO_475 (O_475,N_19140,N_16483);
nand UO_476 (O_476,N_19771,N_16697);
and UO_477 (O_477,N_18019,N_19495);
and UO_478 (O_478,N_19003,N_16849);
xnor UO_479 (O_479,N_19958,N_16277);
and UO_480 (O_480,N_19229,N_16172);
or UO_481 (O_481,N_19776,N_19994);
nand UO_482 (O_482,N_18793,N_19743);
and UO_483 (O_483,N_18911,N_16712);
and UO_484 (O_484,N_19473,N_16128);
and UO_485 (O_485,N_18193,N_17982);
xnor UO_486 (O_486,N_19056,N_18079);
nand UO_487 (O_487,N_18225,N_19068);
nor UO_488 (O_488,N_18541,N_19809);
xnor UO_489 (O_489,N_19917,N_18420);
nor UO_490 (O_490,N_19509,N_17899);
xor UO_491 (O_491,N_18930,N_16294);
nor UO_492 (O_492,N_18566,N_16508);
nand UO_493 (O_493,N_18853,N_18559);
nor UO_494 (O_494,N_19232,N_17969);
nor UO_495 (O_495,N_19782,N_19995);
nor UO_496 (O_496,N_19386,N_16482);
nand UO_497 (O_497,N_17724,N_17939);
and UO_498 (O_498,N_19167,N_19362);
nor UO_499 (O_499,N_17234,N_17837);
or UO_500 (O_500,N_17338,N_18300);
nand UO_501 (O_501,N_16300,N_16219);
nor UO_502 (O_502,N_19053,N_16161);
xor UO_503 (O_503,N_19878,N_19264);
nand UO_504 (O_504,N_18509,N_17510);
xnor UO_505 (O_505,N_16464,N_19787);
and UO_506 (O_506,N_16087,N_16649);
nor UO_507 (O_507,N_18433,N_18022);
xnor UO_508 (O_508,N_17734,N_17929);
nor UO_509 (O_509,N_19330,N_17472);
and UO_510 (O_510,N_17347,N_19391);
nand UO_511 (O_511,N_16916,N_16582);
or UO_512 (O_512,N_19218,N_16750);
and UO_513 (O_513,N_19007,N_17365);
or UO_514 (O_514,N_18755,N_19892);
and UO_515 (O_515,N_19799,N_19027);
nand UO_516 (O_516,N_19085,N_18746);
nand UO_517 (O_517,N_19304,N_17113);
and UO_518 (O_518,N_17741,N_17552);
or UO_519 (O_519,N_16957,N_19715);
nor UO_520 (O_520,N_18314,N_19529);
or UO_521 (O_521,N_19966,N_18366);
nor UO_522 (O_522,N_16180,N_16074);
nor UO_523 (O_523,N_18533,N_17041);
nor UO_524 (O_524,N_17733,N_16270);
nand UO_525 (O_525,N_19566,N_18724);
nor UO_526 (O_526,N_17544,N_18863);
xnor UO_527 (O_527,N_19656,N_18554);
xnor UO_528 (O_528,N_17975,N_17239);
nand UO_529 (O_529,N_16422,N_16414);
nand UO_530 (O_530,N_18150,N_19442);
or UO_531 (O_531,N_17887,N_16375);
or UO_532 (O_532,N_18058,N_16192);
or UO_533 (O_533,N_16485,N_19979);
and UO_534 (O_534,N_16486,N_17043);
and UO_535 (O_535,N_17586,N_19700);
and UO_536 (O_536,N_17537,N_19309);
and UO_537 (O_537,N_18235,N_18082);
nand UO_538 (O_538,N_17191,N_17942);
nand UO_539 (O_539,N_17569,N_19061);
xnor UO_540 (O_540,N_18820,N_16774);
nand UO_541 (O_541,N_17076,N_16558);
nand UO_542 (O_542,N_16310,N_16175);
nand UO_543 (O_543,N_16728,N_19993);
or UO_544 (O_544,N_17872,N_16057);
nor UO_545 (O_545,N_19678,N_16982);
or UO_546 (O_546,N_18548,N_18147);
or UO_547 (O_547,N_19457,N_18399);
nor UO_548 (O_548,N_19447,N_17515);
nor UO_549 (O_549,N_18940,N_17389);
or UO_550 (O_550,N_16496,N_16856);
xnor UO_551 (O_551,N_18613,N_17494);
and UO_552 (O_552,N_16701,N_19584);
nor UO_553 (O_553,N_16559,N_17778);
and UO_554 (O_554,N_17065,N_17301);
nor UO_555 (O_555,N_18704,N_16163);
nand UO_556 (O_556,N_19811,N_16898);
or UO_557 (O_557,N_19493,N_18137);
or UO_558 (O_558,N_17762,N_19853);
nand UO_559 (O_559,N_17385,N_19283);
nand UO_560 (O_560,N_18439,N_17928);
nor UO_561 (O_561,N_16782,N_18226);
xnor UO_562 (O_562,N_19927,N_19448);
or UO_563 (O_563,N_16018,N_16504);
nor UO_564 (O_564,N_16309,N_16657);
or UO_565 (O_565,N_19712,N_19869);
xnor UO_566 (O_566,N_18240,N_16901);
and UO_567 (O_567,N_17317,N_18295);
nand UO_568 (O_568,N_18756,N_17988);
and UO_569 (O_569,N_19844,N_19942);
xor UO_570 (O_570,N_16395,N_18378);
nor UO_571 (O_571,N_18282,N_17376);
xor UO_572 (O_572,N_18319,N_16520);
nand UO_573 (O_573,N_19708,N_17502);
xor UO_574 (O_574,N_18966,N_18221);
nand UO_575 (O_575,N_18565,N_16107);
or UO_576 (O_576,N_17249,N_16056);
nor UO_577 (O_577,N_19727,N_19792);
and UO_578 (O_578,N_18544,N_18302);
or UO_579 (O_579,N_19144,N_17263);
nor UO_580 (O_580,N_18523,N_19612);
nor UO_581 (O_581,N_16591,N_19139);
or UO_582 (O_582,N_16870,N_18375);
nand UO_583 (O_583,N_17775,N_17784);
or UO_584 (O_584,N_17984,N_18914);
nor UO_585 (O_585,N_18825,N_16153);
nor UO_586 (O_586,N_18413,N_18077);
or UO_587 (O_587,N_18201,N_16241);
nand UO_588 (O_588,N_19685,N_19860);
or UO_589 (O_589,N_18355,N_16709);
xnor UO_590 (O_590,N_19358,N_19401);
nor UO_591 (O_591,N_16080,N_16524);
or UO_592 (O_592,N_17288,N_18263);
or UO_593 (O_593,N_19559,N_19832);
xnor UO_594 (O_594,N_16506,N_17536);
nor UO_595 (O_595,N_16736,N_19407);
nand UO_596 (O_596,N_16336,N_16746);
nor UO_597 (O_597,N_17736,N_18899);
xnor UO_598 (O_598,N_17730,N_16465);
and UO_599 (O_599,N_19282,N_19862);
xnor UO_600 (O_600,N_19474,N_18093);
or UO_601 (O_601,N_17079,N_19388);
nand UO_602 (O_602,N_19625,N_18562);
and UO_603 (O_603,N_17469,N_18953);
or UO_604 (O_604,N_19179,N_18973);
nor UO_605 (O_605,N_19428,N_17681);
nand UO_606 (O_606,N_18626,N_16687);
and UO_607 (O_607,N_17633,N_18570);
nand UO_608 (O_608,N_16023,N_19620);
nor UO_609 (O_609,N_18440,N_19907);
nor UO_610 (O_610,N_17527,N_19174);
or UO_611 (O_611,N_19193,N_18376);
nor UO_612 (O_612,N_17210,N_18579);
nor UO_613 (O_613,N_17595,N_16425);
xor UO_614 (O_614,N_19939,N_19769);
nor UO_615 (O_615,N_16223,N_17386);
and UO_616 (O_616,N_17789,N_19036);
nand UO_617 (O_617,N_17014,N_16476);
and UO_618 (O_618,N_16662,N_19480);
xor UO_619 (O_619,N_17006,N_19664);
nor UO_620 (O_620,N_17314,N_18256);
nor UO_621 (O_621,N_17944,N_19104);
nor UO_622 (O_622,N_19935,N_19852);
and UO_623 (O_623,N_19561,N_17214);
or UO_624 (O_624,N_18903,N_16443);
nor UO_625 (O_625,N_17257,N_16316);
or UO_626 (O_626,N_17972,N_19836);
xnor UO_627 (O_627,N_17296,N_16626);
and UO_628 (O_628,N_16684,N_18646);
and UO_629 (O_629,N_19343,N_16442);
nand UO_630 (O_630,N_17034,N_18103);
nand UO_631 (O_631,N_16912,N_18373);
xor UO_632 (O_632,N_19971,N_19651);
xor UO_633 (O_633,N_19032,N_17143);
and UO_634 (O_634,N_16024,N_18306);
or UO_635 (O_635,N_19941,N_19947);
nor UO_636 (O_636,N_19657,N_19191);
or UO_637 (O_637,N_19879,N_17256);
nand UO_638 (O_638,N_19840,N_17350);
nor UO_639 (O_639,N_18379,N_18778);
nand UO_640 (O_640,N_18516,N_19877);
nor UO_641 (O_641,N_19513,N_19622);
nor UO_642 (O_642,N_17683,N_17548);
nand UO_643 (O_643,N_19413,N_18441);
xor UO_644 (O_644,N_17854,N_19900);
or UO_645 (O_645,N_16634,N_17478);
xnor UO_646 (O_646,N_18948,N_16540);
or UO_647 (O_647,N_16606,N_16358);
and UO_648 (O_648,N_17630,N_18357);
and UO_649 (O_649,N_17940,N_19952);
or UO_650 (O_650,N_18534,N_18893);
nand UO_651 (O_651,N_18175,N_17903);
nand UO_652 (O_652,N_19839,N_16609);
or UO_653 (O_653,N_17702,N_19350);
nand UO_654 (O_654,N_16928,N_18100);
and UO_655 (O_655,N_17613,N_17253);
or UO_656 (O_656,N_17024,N_19784);
and UO_657 (O_657,N_16833,N_17077);
nor UO_658 (O_658,N_19004,N_16651);
and UO_659 (O_659,N_17232,N_17668);
and UO_660 (O_660,N_19488,N_18034);
or UO_661 (O_661,N_16493,N_17373);
xnor UO_662 (O_662,N_18106,N_17374);
xnor UO_663 (O_663,N_17576,N_19233);
xor UO_664 (O_664,N_19545,N_18172);
or UO_665 (O_665,N_16590,N_18532);
nor UO_666 (O_666,N_18449,N_18809);
or UO_667 (O_667,N_19172,N_19641);
nor UO_668 (O_668,N_16499,N_16287);
nand UO_669 (O_669,N_18743,N_17136);
nand UO_670 (O_670,N_16988,N_16945);
nor UO_671 (O_671,N_17499,N_16361);
nor UO_672 (O_672,N_19866,N_17574);
and UO_673 (O_673,N_19041,N_19812);
nand UO_674 (O_674,N_19315,N_18748);
or UO_675 (O_675,N_17511,N_18959);
and UO_676 (O_676,N_18391,N_19030);
nor UO_677 (O_677,N_16544,N_19746);
nand UO_678 (O_678,N_17518,N_18325);
or UO_679 (O_679,N_17387,N_16428);
nand UO_680 (O_680,N_16124,N_19756);
or UO_681 (O_681,N_19364,N_18937);
and UO_682 (O_682,N_17738,N_18866);
and UO_683 (O_683,N_17688,N_18924);
xnor UO_684 (O_684,N_19992,N_18075);
and UO_685 (O_685,N_19263,N_17342);
nor UO_686 (O_686,N_19823,N_17561);
xnor UO_687 (O_687,N_19013,N_17271);
and UO_688 (O_688,N_19521,N_17399);
or UO_689 (O_689,N_17002,N_16799);
or UO_690 (O_690,N_19602,N_17960);
xnor UO_691 (O_691,N_16940,N_18353);
or UO_692 (O_692,N_16492,N_16466);
nand UO_693 (O_693,N_18531,N_19734);
or UO_694 (O_694,N_16867,N_18472);
nand UO_695 (O_695,N_17027,N_19722);
xnor UO_696 (O_696,N_16890,N_17073);
and UO_697 (O_697,N_16680,N_16686);
or UO_698 (O_698,N_16203,N_16542);
and UO_699 (O_699,N_17512,N_18676);
or UO_700 (O_700,N_16040,N_19366);
nor UO_701 (O_701,N_16555,N_16263);
and UO_702 (O_702,N_17655,N_18885);
nor UO_703 (O_703,N_18040,N_17441);
nand UO_704 (O_704,N_19226,N_19210);
or UO_705 (O_705,N_17473,N_19302);
or UO_706 (O_706,N_16456,N_18684);
nor UO_707 (O_707,N_16012,N_17990);
nor UO_708 (O_708,N_17295,N_19634);
or UO_709 (O_709,N_17580,N_18573);
or UO_710 (O_710,N_19932,N_19849);
and UO_711 (O_711,N_18887,N_17286);
or UO_712 (O_712,N_17397,N_16394);
nor UO_713 (O_713,N_18512,N_18682);
and UO_714 (O_714,N_16575,N_17201);
and UO_715 (O_715,N_18900,N_18085);
nand UO_716 (O_716,N_18957,N_17653);
and UO_717 (O_717,N_17697,N_18792);
nor UO_718 (O_718,N_19301,N_17357);
and UO_719 (O_719,N_19063,N_19585);
nor UO_720 (O_720,N_16812,N_18504);
nand UO_721 (O_721,N_18634,N_16739);
or UO_722 (O_722,N_16377,N_16953);
nor UO_723 (O_723,N_17280,N_19026);
nand UO_724 (O_724,N_17283,N_16299);
or UO_725 (O_725,N_18589,N_17368);
and UO_726 (O_726,N_17421,N_19273);
and UO_727 (O_727,N_19709,N_16248);
and UO_728 (O_728,N_19277,N_18765);
and UO_729 (O_729,N_19183,N_16909);
nand UO_730 (O_730,N_17505,N_17211);
and UO_731 (O_731,N_17890,N_19245);
or UO_732 (O_732,N_18878,N_18835);
and UO_733 (O_733,N_18690,N_16118);
nor UO_734 (O_734,N_19319,N_19072);
nor UO_735 (O_735,N_19613,N_19841);
nand UO_736 (O_736,N_17915,N_17000);
and UO_737 (O_737,N_17126,N_19489);
xor UO_738 (O_738,N_18115,N_17714);
nor UO_739 (O_739,N_18418,N_17718);
and UO_740 (O_740,N_19896,N_18996);
nor UO_741 (O_741,N_17985,N_19650);
or UO_742 (O_742,N_19234,N_19704);
and UO_743 (O_743,N_19530,N_18700);
or UO_744 (O_744,N_18317,N_17241);
nor UO_745 (O_745,N_18723,N_17993);
nor UO_746 (O_746,N_17420,N_17687);
nor UO_747 (O_747,N_16767,N_19937);
or UO_748 (O_748,N_19471,N_17771);
nor UO_749 (O_749,N_18672,N_18190);
xor UO_750 (O_750,N_19222,N_17495);
xor UO_751 (O_751,N_19363,N_16700);
and UO_752 (O_752,N_17140,N_16179);
or UO_753 (O_753,N_19888,N_17384);
nand UO_754 (O_754,N_19365,N_19269);
xor UO_755 (O_755,N_17918,N_19859);
nand UO_756 (O_756,N_17026,N_16046);
nor UO_757 (O_757,N_17657,N_17860);
nor UO_758 (O_758,N_18237,N_17900);
xnor UO_759 (O_759,N_17111,N_16637);
nand UO_760 (O_760,N_17521,N_18872);
and UO_761 (O_761,N_17498,N_19668);
nand UO_762 (O_762,N_18796,N_18141);
and UO_763 (O_763,N_19847,N_18637);
or UO_764 (O_764,N_16895,N_17196);
nand UO_765 (O_765,N_18841,N_17226);
or UO_766 (O_766,N_16673,N_19376);
nor UO_767 (O_767,N_19691,N_19017);
and UO_768 (O_768,N_18005,N_17997);
nor UO_769 (O_769,N_19573,N_18625);
and UO_770 (O_770,N_17981,N_17562);
and UO_771 (O_771,N_18507,N_19262);
nor UO_772 (O_772,N_18372,N_18067);
nor UO_773 (O_773,N_18727,N_17621);
nand UO_774 (O_774,N_19184,N_16973);
nand UO_775 (O_775,N_16286,N_19415);
nor UO_776 (O_776,N_17017,N_19192);
or UO_777 (O_777,N_18484,N_16624);
xor UO_778 (O_778,N_16679,N_18336);
nor UO_779 (O_779,N_19520,N_16511);
nor UO_780 (O_780,N_16303,N_17361);
or UO_781 (O_781,N_16488,N_18421);
and UO_782 (O_782,N_18777,N_17645);
and UO_783 (O_783,N_19399,N_18281);
nand UO_784 (O_784,N_19379,N_16743);
or UO_785 (O_785,N_18060,N_19627);
or UO_786 (O_786,N_16193,N_18363);
or UO_787 (O_787,N_17168,N_18429);
nand UO_788 (O_788,N_16221,N_16455);
xnor UO_789 (O_789,N_16305,N_19898);
nor UO_790 (O_790,N_19720,N_19492);
or UO_791 (O_791,N_19899,N_19499);
nor UO_792 (O_792,N_19735,N_18970);
nand UO_793 (O_793,N_18788,N_17881);
and UO_794 (O_794,N_18053,N_18539);
or UO_795 (O_795,N_19943,N_16007);
nor UO_796 (O_796,N_19166,N_16724);
nor UO_797 (O_797,N_16228,N_16114);
nand UO_798 (O_798,N_16424,N_17272);
or UO_799 (O_799,N_18956,N_18208);
and UO_800 (O_800,N_17811,N_18298);
nor UO_801 (O_801,N_16693,N_16992);
or UO_802 (O_802,N_17431,N_18042);
nand UO_803 (O_803,N_16371,N_18668);
nand UO_804 (O_804,N_19270,N_19922);
and UO_805 (O_805,N_16855,N_18738);
or UO_806 (O_806,N_16117,N_16723);
or UO_807 (O_807,N_19127,N_17497);
or UO_808 (O_808,N_16176,N_16944);
or UO_809 (O_809,N_17727,N_17375);
nor UO_810 (O_810,N_18581,N_17116);
and UO_811 (O_811,N_16773,N_18934);
and UO_812 (O_812,N_17720,N_19204);
nor UO_813 (O_813,N_16515,N_16411);
nor UO_814 (O_814,N_19398,N_19092);
nor UO_815 (O_815,N_19544,N_17851);
and UO_816 (O_816,N_16577,N_19738);
and UO_817 (O_817,N_19064,N_18561);
nand UO_818 (O_818,N_19617,N_19535);
and UO_819 (O_819,N_16568,N_16605);
xnor UO_820 (O_820,N_19453,N_17149);
nor UO_821 (O_821,N_18601,N_17025);
or UO_822 (O_822,N_17299,N_17850);
or UO_823 (O_823,N_18698,N_18693);
nor UO_824 (O_824,N_18163,N_19096);
nor UO_825 (O_825,N_16891,N_17978);
or UO_826 (O_826,N_16967,N_18496);
or UO_827 (O_827,N_19445,N_16061);
or UO_828 (O_828,N_19858,N_19334);
nand UO_829 (O_829,N_19893,N_17867);
xor UO_830 (O_830,N_16817,N_16042);
nor UO_831 (O_831,N_18043,N_16019);
nor UO_832 (O_832,N_18311,N_17874);
nor UO_833 (O_833,N_18582,N_17568);
xnor UO_834 (O_834,N_17482,N_18923);
and UO_835 (O_835,N_16401,N_18099);
or UO_836 (O_836,N_19540,N_17022);
or UO_837 (O_837,N_17114,N_18401);
or UO_838 (O_838,N_19472,N_16406);
xnor UO_839 (O_839,N_16815,N_19250);
and UO_840 (O_840,N_19550,N_16722);
or UO_841 (O_841,N_19796,N_16162);
nand UO_842 (O_842,N_18214,N_16314);
and UO_843 (O_843,N_16846,N_16762);
nor UO_844 (O_844,N_19287,N_18906);
nand UO_845 (O_845,N_18666,N_16484);
nand UO_846 (O_846,N_19661,N_19132);
or UO_847 (O_847,N_19011,N_19463);
and UO_848 (O_848,N_19810,N_19558);
xor UO_849 (O_849,N_19105,N_19337);
nand UO_850 (O_850,N_16960,N_18926);
nor UO_851 (O_851,N_16386,N_16578);
xnor UO_852 (O_852,N_18415,N_16468);
nor UO_853 (O_853,N_16116,N_19593);
xnor UO_854 (O_854,N_17508,N_18448);
nand UO_855 (O_855,N_17146,N_18338);
nor UO_856 (O_856,N_19506,N_17245);
and UO_857 (O_857,N_17273,N_18272);
nand UO_858 (O_858,N_16332,N_16752);
xnor UO_859 (O_859,N_16716,N_18725);
or UO_860 (O_860,N_16979,N_19251);
nor UO_861 (O_861,N_17617,N_16043);
nor UO_862 (O_862,N_19164,N_19342);
nand UO_863 (O_863,N_16196,N_17772);
nand UO_864 (O_864,N_17487,N_18648);
nor UO_865 (O_865,N_18553,N_16903);
nand UO_866 (O_866,N_17298,N_17109);
or UO_867 (O_867,N_18908,N_19838);
or UO_868 (O_868,N_18116,N_16845);
nand UO_869 (O_869,N_19914,N_17962);
nor UO_870 (O_870,N_19976,N_16268);
nand UO_871 (O_871,N_16643,N_18691);
and UO_872 (O_872,N_19271,N_17470);
and UO_873 (O_873,N_18024,N_19510);
nor UO_874 (O_874,N_17701,N_19403);
nor UO_875 (O_875,N_17019,N_18307);
nand UO_876 (O_876,N_17679,N_18310);
and UO_877 (O_877,N_18114,N_17131);
nor UO_878 (O_878,N_16794,N_18808);
or UO_879 (O_879,N_17946,N_16943);
nand UO_880 (O_880,N_18568,N_18794);
or UO_881 (O_881,N_19055,N_17858);
and UO_882 (O_882,N_16708,N_18751);
nor UO_883 (O_883,N_17500,N_17677);
xnor UO_884 (O_884,N_16384,N_19220);
and UO_885 (O_885,N_19073,N_16611);
nand UO_886 (O_886,N_18468,N_19196);
or UO_887 (O_887,N_17654,N_18265);
nand UO_888 (O_888,N_16208,N_17240);
nand UO_889 (O_889,N_16147,N_17044);
or UO_890 (O_890,N_16550,N_17030);
nand UO_891 (O_891,N_16748,N_17279);
nor UO_892 (O_892,N_18942,N_17909);
nor UO_893 (O_893,N_16404,N_18713);
nand UO_894 (O_894,N_17608,N_18688);
or UO_895 (O_895,N_19662,N_18950);
or UO_896 (O_896,N_17693,N_18428);
or UO_897 (O_897,N_18202,N_16397);
nand UO_898 (O_898,N_17801,N_19498);
and UO_899 (O_899,N_19359,N_16216);
nand UO_900 (O_900,N_19781,N_18460);
nand UO_901 (O_901,N_19188,N_17859);
nor UO_902 (O_902,N_16942,N_17749);
xnor UO_903 (O_903,N_19437,N_18069);
nand UO_904 (O_904,N_18860,N_18787);
or UO_905 (O_905,N_16439,N_16413);
nor UO_906 (O_906,N_16588,N_18600);
xor UO_907 (O_907,N_18502,N_17465);
and UO_908 (O_908,N_17254,N_19103);
and UO_909 (O_909,N_16675,N_17821);
nand UO_910 (O_910,N_19012,N_17056);
or UO_911 (O_911,N_18806,N_16044);
xnor UO_912 (O_912,N_19046,N_18196);
or UO_913 (O_913,N_16792,N_17153);
nor UO_914 (O_914,N_16213,N_18073);
nor UO_915 (O_915,N_17480,N_18644);
or UO_916 (O_916,N_17989,N_18795);
nor UO_917 (O_917,N_16121,N_16417);
and UO_918 (O_918,N_17300,N_16462);
nor UO_919 (O_919,N_18330,N_16278);
nor UO_920 (O_920,N_16886,N_17607);
and UO_921 (O_921,N_19982,N_16276);
and UO_922 (O_922,N_19060,N_18036);
xnor UO_923 (O_923,N_18935,N_17166);
and UO_924 (O_924,N_18521,N_16337);
or UO_925 (O_925,N_16449,N_16654);
xor UO_926 (O_926,N_16780,N_17699);
nand UO_927 (O_927,N_17377,N_17005);
or UO_928 (O_928,N_19518,N_16915);
xor UO_929 (O_929,N_16313,N_18917);
xnor UO_930 (O_930,N_16295,N_18309);
or UO_931 (O_931,N_16719,N_17105);
nor UO_932 (O_932,N_16950,N_19331);
or UO_933 (O_933,N_17324,N_18875);
xnor UO_934 (O_934,N_19082,N_17973);
or UO_935 (O_935,N_16220,N_17406);
nor UO_936 (O_936,N_19122,N_19626);
nand UO_937 (O_937,N_18641,N_16806);
nand UO_938 (O_938,N_19880,N_18643);
and UO_939 (O_939,N_19514,N_17875);
nand UO_940 (O_940,N_18315,N_19960);
nor UO_941 (O_941,N_19107,N_19988);
nand UO_942 (O_942,N_18580,N_19674);
nand UO_943 (O_943,N_17394,N_16929);
nand UO_944 (O_944,N_16365,N_16528);
or UO_945 (O_945,N_17463,N_17058);
or UO_946 (O_946,N_19430,N_18247);
nand UO_947 (O_947,N_19469,N_18538);
and UO_948 (O_948,N_17792,N_16398);
nand UO_949 (O_949,N_16359,N_16170);
xnor UO_950 (O_950,N_16821,N_16628);
and UO_951 (O_951,N_19441,N_18486);
or UO_952 (O_952,N_19936,N_16747);
xor UO_953 (O_953,N_16914,N_18660);
nand UO_954 (O_954,N_16881,N_17980);
xor UO_955 (O_955,N_17766,N_17987);
nor UO_956 (O_956,N_18503,N_16518);
nand UO_957 (O_957,N_16616,N_16050);
or UO_958 (O_958,N_18610,N_16210);
or UO_959 (O_959,N_19190,N_16842);
or UO_960 (O_960,N_18928,N_17400);
or UO_961 (O_961,N_19326,N_19916);
xor UO_962 (O_962,N_16754,N_17012);
or UO_963 (O_963,N_19628,N_18347);
and UO_964 (O_964,N_19845,N_16352);
nor UO_965 (O_965,N_16157,N_19340);
nor UO_966 (O_966,N_16859,N_19775);
nand UO_967 (O_967,N_19381,N_17036);
nor UO_968 (O_968,N_17809,N_19905);
and UO_969 (O_969,N_19427,N_16644);
and UO_970 (O_970,N_16137,N_19768);
and UO_971 (O_971,N_17823,N_17897);
or UO_972 (O_972,N_18301,N_17810);
and UO_973 (O_973,N_16689,N_19372);
and UO_974 (O_974,N_19224,N_16924);
and UO_975 (O_975,N_17087,N_17593);
and UO_976 (O_976,N_18318,N_18412);
and UO_977 (O_977,N_17069,N_18200);
nor UO_978 (O_978,N_17462,N_18016);
nor UO_979 (O_979,N_17171,N_16211);
nor UO_980 (O_980,N_19642,N_18339);
nor UO_981 (O_981,N_17333,N_19536);
xor UO_982 (O_982,N_19586,N_19291);
or UO_983 (O_983,N_16127,N_19742);
and UO_984 (O_984,N_18971,N_17124);
nand UO_985 (O_985,N_17477,N_18995);
nor UO_986 (O_986,N_19693,N_19409);
or UO_987 (O_987,N_16884,N_19990);
xor UO_988 (O_988,N_18381,N_16574);
and UO_989 (O_989,N_18473,N_17746);
or UO_990 (O_990,N_18932,N_19871);
xnor UO_991 (O_991,N_19848,N_18655);
xor UO_992 (O_992,N_17933,N_18028);
nand UO_993 (O_993,N_17258,N_19996);
nand UO_994 (O_994,N_18555,N_19683);
nor UO_995 (O_995,N_17471,N_18506);
xnor UO_996 (O_996,N_17032,N_19460);
and UO_997 (O_997,N_16844,N_16000);
nand UO_998 (O_998,N_17008,N_19790);
nor UO_999 (O_999,N_19870,N_16936);
nand UO_1000 (O_1000,N_16291,N_17155);
and UO_1001 (O_1001,N_17950,N_16009);
or UO_1002 (O_1002,N_17647,N_16534);
nand UO_1003 (O_1003,N_16112,N_18546);
and UO_1004 (O_1004,N_18474,N_18611);
nor UO_1005 (O_1005,N_18345,N_16322);
xnor UO_1006 (O_1006,N_19703,N_16296);
nor UO_1007 (O_1007,N_17686,N_16151);
nor UO_1008 (O_1008,N_18764,N_18014);
nor UO_1009 (O_1009,N_18149,N_16786);
nor UO_1010 (O_1010,N_17589,N_18960);
nand UO_1011 (O_1011,N_17379,N_16457);
and UO_1012 (O_1012,N_17656,N_19475);
nand UO_1013 (O_1013,N_17169,N_17396);
and UO_1014 (O_1014,N_17320,N_16598);
nand UO_1015 (O_1015,N_17182,N_16091);
nor UO_1016 (O_1016,N_19534,N_17995);
and UO_1017 (O_1017,N_19855,N_16993);
and UO_1018 (O_1018,N_19986,N_18627);
nand UO_1019 (O_1019,N_16676,N_16391);
and UO_1020 (O_1020,N_18849,N_18335);
and UO_1021 (O_1021,N_19603,N_18910);
nand UO_1022 (O_1022,N_19292,N_16252);
or UO_1023 (O_1023,N_19814,N_17366);
xor UO_1024 (O_1024,N_17588,N_18834);
or UO_1025 (O_1025,N_19006,N_16869);
and UO_1026 (O_1026,N_16267,N_18994);
nand UO_1027 (O_1027,N_17712,N_17754);
nand UO_1028 (O_1028,N_18178,N_16079);
nor UO_1029 (O_1029,N_18927,N_18446);
nand UO_1030 (O_1030,N_18451,N_18362);
nand UO_1031 (O_1031,N_16016,N_16699);
nand UO_1032 (O_1032,N_16965,N_17412);
or UO_1033 (O_1033,N_18400,N_17145);
and UO_1034 (O_1034,N_17864,N_16459);
and UO_1035 (O_1035,N_17506,N_19289);
nand UO_1036 (O_1036,N_16099,N_16619);
nand UO_1037 (O_1037,N_19249,N_17773);
and UO_1038 (O_1038,N_16647,N_17170);
or UO_1039 (O_1039,N_19237,N_16923);
and UO_1040 (O_1040,N_16766,N_19209);
and UO_1041 (O_1041,N_16758,N_17849);
nand UO_1042 (O_1042,N_16897,N_16338);
or UO_1043 (O_1043,N_16381,N_17976);
nand UO_1044 (O_1044,N_17907,N_18180);
nand UO_1045 (O_1045,N_19934,N_16620);
or UO_1046 (O_1046,N_19659,N_19236);
nand UO_1047 (O_1047,N_18068,N_19432);
nand UO_1048 (O_1048,N_17661,N_17451);
and UO_1049 (O_1049,N_17763,N_17004);
xor UO_1050 (O_1050,N_16955,N_19450);
nand UO_1051 (O_1051,N_17259,N_17952);
or UO_1052 (O_1052,N_16917,N_19079);
xnor UO_1053 (O_1053,N_16204,N_17911);
nor UO_1054 (O_1054,N_19484,N_19436);
nand UO_1055 (O_1055,N_19181,N_17275);
xnor UO_1056 (O_1056,N_17587,N_18304);
nor UO_1057 (O_1057,N_16317,N_17097);
or UO_1058 (O_1058,N_19770,N_16255);
or UO_1059 (O_1059,N_19533,N_18695);
nor UO_1060 (O_1060,N_16983,N_17695);
nand UO_1061 (O_1061,N_18784,N_18422);
and UO_1062 (O_1062,N_19347,N_19919);
and UO_1063 (O_1063,N_19677,N_19223);
nor UO_1064 (O_1064,N_19047,N_19417);
nand UO_1065 (O_1065,N_17371,N_18612);
or UO_1066 (O_1066,N_17491,N_16002);
or UO_1067 (O_1067,N_18686,N_18915);
nand UO_1068 (O_1068,N_17882,N_19205);
xor UO_1069 (O_1069,N_19247,N_17752);
and UO_1070 (O_1070,N_19024,N_18677);
and UO_1071 (O_1071,N_16810,N_17489);
nand UO_1072 (O_1072,N_17533,N_17598);
nand UO_1073 (O_1073,N_16068,N_17577);
nand UO_1074 (O_1074,N_16274,N_16995);
or UO_1075 (O_1075,N_18155,N_19886);
nor UO_1076 (O_1076,N_16372,N_16653);
and UO_1077 (O_1077,N_17174,N_16640);
and UO_1078 (O_1078,N_19077,N_16941);
and UO_1079 (O_1079,N_17546,N_16866);
or UO_1080 (O_1080,N_16837,N_16584);
and UO_1081 (O_1081,N_17289,N_17680);
or UO_1082 (O_1082,N_18487,N_16084);
nand UO_1083 (O_1083,N_19961,N_18223);
nor UO_1084 (O_1084,N_18650,N_19387);
or UO_1085 (O_1085,N_17430,N_18188);
or UO_1086 (O_1086,N_16878,N_16580);
and UO_1087 (O_1087,N_16622,N_18716);
nand UO_1088 (O_1088,N_16996,N_18198);
and UO_1089 (O_1089,N_18712,N_19883);
xor UO_1090 (O_1090,N_16190,N_19168);
nand UO_1091 (O_1091,N_17028,N_18615);
nor UO_1092 (O_1092,N_17045,N_16082);
nand UO_1093 (O_1093,N_16340,N_19126);
nand UO_1094 (O_1094,N_18522,N_16594);
nor UO_1095 (O_1095,N_18133,N_16184);
or UO_1096 (O_1096,N_16356,N_18640);
and UO_1097 (O_1097,N_18425,N_17068);
and UO_1098 (O_1098,N_18007,N_16769);
nand UO_1099 (O_1099,N_18605,N_19675);
nand UO_1100 (O_1100,N_19515,N_16745);
or UO_1101 (O_1101,N_16054,N_17839);
nand UO_1102 (O_1102,N_19208,N_17230);
or UO_1103 (O_1103,N_16727,N_19541);
or UO_1104 (O_1104,N_18164,N_19946);
and UO_1105 (O_1105,N_19731,N_16400);
nor UO_1106 (O_1106,N_19374,N_17551);
and UO_1107 (O_1107,N_19876,N_19136);
or UO_1108 (O_1108,N_19500,N_19178);
and UO_1109 (O_1109,N_18481,N_19361);
nor UO_1110 (O_1110,N_19383,N_17084);
or UO_1111 (O_1111,N_17838,N_18323);
and UO_1112 (O_1112,N_18258,N_17719);
nand UO_1113 (O_1113,N_17648,N_18135);
and UO_1114 (O_1114,N_16507,N_18635);
xor UO_1115 (O_1115,N_19539,N_17635);
nand UO_1116 (O_1116,N_19596,N_18117);
or UO_1117 (O_1117,N_19649,N_17983);
nor UO_1118 (O_1118,N_18260,N_16141);
xor UO_1119 (O_1119,N_19713,N_19938);
nor UO_1120 (O_1120,N_18008,N_17082);
and UO_1121 (O_1121,N_16312,N_19015);
and UO_1122 (O_1122,N_19653,N_18055);
and UO_1123 (O_1123,N_17092,N_16596);
and UO_1124 (O_1124,N_17636,N_19959);
and UO_1125 (O_1125,N_18059,N_17829);
nand UO_1126 (O_1126,N_18857,N_18947);
nor UO_1127 (O_1127,N_16865,N_16770);
nor UO_1128 (O_1128,N_17629,N_19248);
and UO_1129 (O_1129,N_18371,N_19125);
or UO_1130 (O_1130,N_17865,N_19889);
and UO_1131 (O_1131,N_19228,N_18987);
or UO_1132 (O_1132,N_19152,N_16354);
xor UO_1133 (O_1133,N_16695,N_19725);
nand UO_1134 (O_1134,N_18408,N_18719);
and UO_1135 (O_1135,N_17070,N_16452);
or UO_1136 (O_1136,N_18901,N_17652);
nor UO_1137 (O_1137,N_16280,N_17709);
nor UO_1138 (O_1138,N_19071,N_18717);
or UO_1139 (O_1139,N_17876,N_19805);
and UO_1140 (O_1140,N_18065,N_16863);
and UO_1141 (O_1141,N_17556,N_18545);
and UO_1142 (O_1142,N_19360,N_18427);
and UO_1143 (O_1143,N_16677,N_17541);
nand UO_1144 (O_1144,N_16519,N_17437);
nand UO_1145 (O_1145,N_19669,N_19296);
and UO_1146 (O_1146,N_19408,N_16986);
nor UO_1147 (O_1147,N_17600,N_17642);
xor UO_1148 (O_1148,N_16658,N_17822);
nor UO_1149 (O_1149,N_17549,N_16521);
nor UO_1150 (O_1150,N_16146,N_16974);
or UO_1151 (O_1151,N_19438,N_16430);
xnor UO_1152 (O_1152,N_17095,N_17776);
nor UO_1153 (O_1153,N_16905,N_16545);
nor UO_1154 (O_1154,N_18549,N_19997);
and UO_1155 (O_1155,N_16302,N_19106);
or UO_1156 (O_1156,N_17742,N_18664);
nor UO_1157 (O_1157,N_18558,N_18920);
xnor UO_1158 (O_1158,N_18224,N_18817);
nand UO_1159 (O_1159,N_19672,N_16471);
or UO_1160 (O_1160,N_18328,N_17721);
and UO_1161 (O_1161,N_17242,N_16217);
nor UO_1162 (O_1162,N_19043,N_18505);
or UO_1163 (O_1163,N_17737,N_18921);
xnor UO_1164 (O_1164,N_18333,N_19630);
nor UO_1165 (O_1165,N_17516,N_17582);
and UO_1166 (O_1166,N_17039,N_18157);
and UO_1167 (O_1167,N_17133,N_17698);
nor UO_1168 (O_1168,N_17138,N_19663);
or UO_1169 (O_1169,N_19385,N_19213);
nand UO_1170 (O_1170,N_19806,N_16892);
nand UO_1171 (O_1171,N_19243,N_17640);
nand UO_1172 (O_1172,N_19496,N_17381);
nand UO_1173 (O_1173,N_19490,N_16261);
nor UO_1174 (O_1174,N_18243,N_17120);
nand UO_1175 (O_1175,N_18246,N_18370);
nor UO_1176 (O_1176,N_16014,N_17526);
xnor UO_1177 (O_1177,N_17127,N_17831);
and UO_1178 (O_1178,N_17826,N_19614);
nor UO_1179 (O_1179,N_18290,N_18444);
nor UO_1180 (O_1180,N_16738,N_16652);
nor UO_1181 (O_1181,N_17716,N_19426);
nand UO_1182 (O_1182,N_17459,N_16333);
nand UO_1183 (O_1183,N_16906,N_19972);
or UO_1184 (O_1184,N_17031,N_18002);
and UO_1185 (O_1185,N_16804,N_17912);
and UO_1186 (O_1186,N_16100,N_19505);
and UO_1187 (O_1187,N_17748,N_18624);
and UO_1188 (O_1188,N_18753,N_18405);
or UO_1189 (O_1189,N_19763,N_18411);
nand UO_1190 (O_1190,N_16927,N_17096);
and UO_1191 (O_1191,N_17751,N_16229);
nor UO_1192 (O_1192,N_19686,N_17799);
nand UO_1193 (O_1193,N_17224,N_19631);
or UO_1194 (O_1194,N_16227,N_16379);
nor UO_1195 (O_1195,N_18064,N_17797);
xor UO_1196 (O_1196,N_18780,N_17236);
and UO_1197 (O_1197,N_16347,N_19284);
or UO_1198 (O_1198,N_17759,N_18013);
nor UO_1199 (O_1199,N_17268,N_16956);
nand UO_1200 (O_1200,N_18242,N_18993);
and UO_1201 (O_1201,N_19052,N_18350);
nor UO_1202 (O_1202,N_19451,N_19108);
or UO_1203 (O_1203,N_16807,N_18961);
and UO_1204 (O_1204,N_18810,N_16222);
or UO_1205 (O_1205,N_19974,N_19549);
nand UO_1206 (O_1206,N_19042,N_18173);
xnor UO_1207 (O_1207,N_17180,N_19411);
nor UO_1208 (O_1208,N_19507,N_18815);
and UO_1209 (O_1209,N_16047,N_16478);
nor UO_1210 (O_1210,N_19230,N_16075);
xor UO_1211 (O_1211,N_18590,N_16882);
or UO_1212 (O_1212,N_18126,N_19817);
nor UO_1213 (O_1213,N_16385,N_19519);
and UO_1214 (O_1214,N_19434,N_17507);
and UO_1215 (O_1215,N_18864,N_17352);
nand UO_1216 (O_1216,N_19325,N_16154);
and UO_1217 (O_1217,N_18593,N_17935);
and UO_1218 (O_1218,N_19801,N_17846);
xor UO_1219 (O_1219,N_17786,N_19753);
nor UO_1220 (O_1220,N_19818,N_17581);
nor UO_1221 (O_1221,N_19757,N_19764);
nand UO_1222 (O_1222,N_18285,N_18749);
and UO_1223 (O_1223,N_19732,N_19739);
or UO_1224 (O_1224,N_19206,N_17212);
and UO_1225 (O_1225,N_19333,N_19062);
nor UO_1226 (O_1226,N_17513,N_19556);
nand UO_1227 (O_1227,N_18097,N_19719);
nand UO_1228 (O_1228,N_18584,N_18944);
or UO_1229 (O_1229,N_19798,N_17700);
xnor UO_1230 (O_1230,N_16601,N_17364);
or UO_1231 (O_1231,N_16681,N_16461);
nand UO_1232 (O_1232,N_18340,N_17417);
xor UO_1233 (O_1233,N_19592,N_18888);
nand UO_1234 (O_1234,N_17281,N_18352);
and UO_1235 (O_1235,N_19163,N_17018);
nor UO_1236 (O_1236,N_19468,N_19009);
and UO_1237 (O_1237,N_16202,N_16603);
xnor UO_1238 (O_1238,N_16120,N_18969);
nor UO_1239 (O_1239,N_19694,N_17827);
nand UO_1240 (O_1240,N_17963,N_18632);
and UO_1241 (O_1241,N_18575,N_19033);
nor UO_1242 (O_1242,N_19479,N_18048);
and UO_1243 (O_1243,N_19697,N_17460);
and UO_1244 (O_1244,N_16212,N_16741);
and UO_1245 (O_1245,N_16823,N_17178);
nand UO_1246 (O_1246,N_18443,N_17540);
or UO_1247 (O_1247,N_18184,N_18858);
and UO_1248 (O_1248,N_18026,N_18485);
or UO_1249 (O_1249,N_16613,N_17605);
and UO_1250 (O_1250,N_17110,N_16775);
nor UO_1251 (O_1251,N_17123,N_16899);
or UO_1252 (O_1252,N_18086,N_16063);
nand UO_1253 (O_1253,N_16661,N_17403);
nand UO_1254 (O_1254,N_19578,N_17866);
and UO_1255 (O_1255,N_19440,N_18380);
nor UO_1256 (O_1256,N_19560,N_19175);
nand UO_1257 (O_1257,N_19795,N_17624);
and UO_1258 (O_1258,N_16538,N_18445);
nor UO_1259 (O_1259,N_16645,N_18364);
nor UO_1260 (O_1260,N_16039,N_17666);
xor UO_1261 (O_1261,N_19497,N_16937);
nand UO_1262 (O_1262,N_18951,N_18862);
or UO_1263 (O_1263,N_19645,N_19851);
xnor UO_1264 (O_1264,N_18299,N_16581);
nor UO_1265 (O_1265,N_17147,N_16744);
nor UO_1266 (O_1266,N_17722,N_17957);
and UO_1267 (O_1267,N_18230,N_19964);
nor UO_1268 (O_1268,N_17917,N_18557);
or UO_1269 (O_1269,N_18331,N_17824);
nor UO_1270 (O_1270,N_17426,N_17922);
or UO_1271 (O_1271,N_18123,N_16329);
nand UO_1272 (O_1272,N_18606,N_19537);
nand UO_1273 (O_1273,N_16403,N_19212);
and UO_1274 (O_1274,N_19682,N_17926);
or UO_1275 (O_1275,N_19482,N_19390);
nand UO_1276 (O_1276,N_16554,N_19512);
and UO_1277 (O_1277,N_17966,N_18346);
nor UO_1278 (O_1278,N_18394,N_16523);
or UO_1279 (O_1279,N_17609,N_19025);
nor UO_1280 (O_1280,N_17311,N_18608);
nand UO_1281 (O_1281,N_17233,N_18816);
or UO_1282 (O_1282,N_17729,N_18812);
and UO_1283 (O_1283,N_17216,N_16587);
xnor UO_1284 (O_1284,N_16095,N_19286);
or UO_1285 (O_1285,N_17603,N_19926);
and UO_1286 (O_1286,N_16931,N_16349);
nor UO_1287 (O_1287,N_19710,N_17676);
nor UO_1288 (O_1288,N_18799,N_16822);
or UO_1289 (O_1289,N_17456,N_17325);
nor UO_1290 (O_1290,N_19185,N_16032);
nor UO_1291 (O_1291,N_16861,N_18083);
nand UO_1292 (O_1292,N_18262,N_16198);
and UO_1293 (O_1293,N_18832,N_19207);
nor UO_1294 (O_1294,N_18977,N_18706);
nor UO_1295 (O_1295,N_19008,N_17539);
nand UO_1296 (O_1296,N_18933,N_19711);
nand UO_1297 (O_1297,N_19802,N_17927);
or UO_1298 (O_1298,N_18209,N_19215);
xnor UO_1299 (O_1299,N_17584,N_18476);
or UO_1300 (O_1300,N_16826,N_17106);
or UO_1301 (O_1301,N_18771,N_17132);
nand UO_1302 (O_1302,N_16036,N_16841);
nand UO_1303 (O_1303,N_17139,N_19684);
and UO_1304 (O_1304,N_17639,N_17758);
or UO_1305 (O_1305,N_19405,N_16318);
nand UO_1306 (O_1306,N_16078,N_19581);
or UO_1307 (O_1307,N_17450,N_16948);
xnor UO_1308 (O_1308,N_18633,N_16249);
or UO_1309 (O_1309,N_18327,N_18879);
nor UO_1310 (O_1310,N_16169,N_18483);
and UO_1311 (O_1311,N_16234,N_18018);
nand UO_1312 (O_1312,N_18424,N_17921);
nor UO_1313 (O_1313,N_16410,N_17020);
and UO_1314 (O_1314,N_19023,N_18670);
and UO_1315 (O_1315,N_16579,N_17415);
or UO_1316 (O_1316,N_16500,N_16883);
nor UO_1317 (O_1317,N_19736,N_19766);
or UO_1318 (O_1318,N_18699,N_16665);
nand UO_1319 (O_1319,N_19882,N_17010);
or UO_1320 (O_1320,N_19531,N_17104);
or UO_1321 (O_1321,N_16022,N_17532);
xnor UO_1322 (O_1322,N_17442,N_17072);
nand UO_1323 (O_1323,N_17861,N_19621);
xor UO_1324 (O_1324,N_18898,N_16195);
and UO_1325 (O_1325,N_17190,N_19238);
xnor UO_1326 (O_1326,N_18457,N_17862);
xor UO_1327 (O_1327,N_16980,N_16004);
and UO_1328 (O_1328,N_16173,N_17905);
and UO_1329 (O_1329,N_17003,N_16214);
nor UO_1330 (O_1330,N_16659,N_19135);
or UO_1331 (O_1331,N_17064,N_16368);
nor UO_1332 (O_1332,N_17870,N_18991);
or UO_1333 (O_1333,N_16836,N_18592);
nor UO_1334 (O_1334,N_19894,N_17898);
and UO_1335 (O_1335,N_18464,N_16279);
or UO_1336 (O_1336,N_18248,N_18092);
xnor UO_1337 (O_1337,N_18665,N_16035);
and UO_1338 (O_1338,N_17830,N_17961);
nand UO_1339 (O_1339,N_16281,N_17848);
or UO_1340 (O_1340,N_19227,N_17836);
xor UO_1341 (O_1341,N_17795,N_17408);
nand UO_1342 (O_1342,N_17327,N_17528);
nor UO_1343 (O_1343,N_16618,N_18153);
xor UO_1344 (O_1344,N_18873,N_18552);
nand UO_1345 (O_1345,N_18721,N_16972);
or UO_1346 (O_1346,N_18467,N_16472);
and UO_1347 (O_1347,N_16498,N_19666);
nand UO_1348 (O_1348,N_19985,N_16419);
nor UO_1349 (O_1349,N_16535,N_18090);
or UO_1350 (O_1350,N_16185,N_19562);
xnor UO_1351 (O_1351,N_16328,N_18649);
or UO_1352 (O_1352,N_18101,N_18894);
or UO_1353 (O_1353,N_16783,N_19131);
or UO_1354 (O_1354,N_17037,N_16563);
and UO_1355 (O_1355,N_17534,N_17359);
or UO_1356 (O_1356,N_19874,N_19180);
xnor UO_1357 (O_1357,N_18414,N_17454);
and UO_1358 (O_1358,N_17439,N_16348);
and UO_1359 (O_1359,N_19352,N_19084);
and UO_1360 (O_1360,N_17671,N_19487);
nand UO_1361 (O_1361,N_19080,N_16262);
nor UO_1362 (O_1362,N_18195,N_18233);
nor UO_1363 (O_1363,N_19665,N_19142);
nor UO_1364 (O_1364,N_19890,N_16490);
nand UO_1365 (O_1365,N_16160,N_17802);
nor UO_1366 (O_1366,N_19511,N_18636);
or UO_1367 (O_1367,N_19252,N_17951);
nand UO_1368 (O_1368,N_17011,N_17622);
nand UO_1369 (O_1369,N_18322,N_16900);
nor UO_1370 (O_1370,N_18436,N_17794);
or UO_1371 (O_1371,N_19371,N_17798);
xor UO_1372 (O_1372,N_18530,N_16572);
nor UO_1373 (O_1373,N_18326,N_17418);
xnor UO_1374 (O_1374,N_17447,N_16608);
xor UO_1375 (O_1375,N_19639,N_18697);
or UO_1376 (O_1376,N_18596,N_18261);
nand UO_1377 (O_1377,N_16230,N_16632);
or UO_1378 (O_1378,N_16441,N_17302);
nand UO_1379 (O_1379,N_16152,N_17125);
nand UO_1380 (O_1380,N_18563,N_19444);
xnor UO_1381 (O_1381,N_17638,N_18964);
or UO_1382 (O_1382,N_17307,N_17016);
or UO_1383 (O_1383,N_16351,N_17194);
or UO_1384 (O_1384,N_18478,N_18913);
or UO_1385 (O_1385,N_16907,N_18104);
or UO_1386 (O_1386,N_19820,N_19861);
or UO_1387 (O_1387,N_17176,N_19696);
nand UO_1388 (O_1388,N_16667,N_18492);
or UO_1389 (O_1389,N_17341,N_16285);
or UO_1390 (O_1390,N_17934,N_16235);
or UO_1391 (O_1391,N_19305,N_17747);
nand UO_1392 (O_1392,N_16126,N_16489);
nor UO_1393 (O_1393,N_18218,N_17198);
and UO_1394 (O_1394,N_17665,N_17192);
nor UO_1395 (O_1395,N_18207,N_17913);
nor UO_1396 (O_1396,N_16233,N_17331);
nand UO_1397 (O_1397,N_16850,N_16664);
nor UO_1398 (O_1398,N_16122,N_16970);
xor UO_1399 (O_1399,N_18535,N_17038);
nor UO_1400 (O_1400,N_18621,N_19470);
and UO_1401 (O_1401,N_17061,N_18603);
and UO_1402 (O_1402,N_17186,N_16756);
xnor UO_1403 (O_1403,N_16494,N_16656);
nand UO_1404 (O_1404,N_19274,N_18616);
nor UO_1405 (O_1405,N_18166,N_16357);
nor UO_1406 (O_1406,N_16879,N_16918);
nand UO_1407 (O_1407,N_18891,N_19094);
xor UO_1408 (O_1408,N_18337,N_19570);
and UO_1409 (O_1409,N_19895,N_18296);
nor UO_1410 (O_1410,N_19699,N_19389);
or UO_1411 (O_1411,N_17225,N_18454);
nor UO_1412 (O_1412,N_17100,N_19928);
xor UO_1413 (O_1413,N_19854,N_17029);
nor UO_1414 (O_1414,N_19998,N_17048);
nor UO_1415 (O_1415,N_19266,N_19788);
nand UO_1416 (O_1416,N_19329,N_17433);
and UO_1417 (O_1417,N_17817,N_19419);
nand UO_1418 (O_1418,N_18479,N_17583);
and UO_1419 (O_1419,N_18752,N_16549);
nand UO_1420 (O_1420,N_17509,N_17130);
and UO_1421 (O_1421,N_17063,N_16297);
and UO_1422 (O_1422,N_16062,N_17081);
nor UO_1423 (O_1423,N_18842,N_19112);
or UO_1424 (O_1424,N_19965,N_16320);
nor UO_1425 (O_1425,N_16434,N_17213);
nand UO_1426 (O_1426,N_16164,N_17856);
and UO_1427 (O_1427,N_16307,N_17053);
nand UO_1428 (O_1428,N_17783,N_16854);
or UO_1429 (O_1429,N_16013,N_19454);
nor UO_1430 (O_1430,N_19313,N_19141);
nor UO_1431 (O_1431,N_19655,N_18289);
nand UO_1432 (O_1432,N_17842,N_17684);
or UO_1433 (O_1433,N_18861,N_16081);
nand UO_1434 (O_1434,N_18393,N_17543);
xor UO_1435 (O_1435,N_18211,N_19146);
and UO_1436 (O_1436,N_16393,N_17290);
nand UO_1437 (O_1437,N_17923,N_17222);
nor UO_1438 (O_1438,N_19930,N_17316);
xnor UO_1439 (O_1439,N_17367,N_16707);
nand UO_1440 (O_1440,N_19231,N_18588);
xor UO_1441 (O_1441,N_16951,N_16711);
and UO_1442 (O_1442,N_19902,N_19702);
nor UO_1443 (O_1443,N_18631,N_19977);
or UO_1444 (O_1444,N_19298,N_16006);
nand UO_1445 (O_1445,N_16038,N_18782);
nand UO_1446 (O_1446,N_17164,N_18938);
or UO_1447 (O_1447,N_17979,N_18629);
xor UO_1448 (O_1448,N_17229,N_17093);
nand UO_1449 (O_1449,N_17994,N_16543);
and UO_1450 (O_1450,N_19640,N_17346);
or UO_1451 (O_1451,N_18614,N_19199);
nand UO_1452 (O_1452,N_17358,N_17001);
xor UO_1453 (O_1453,N_19658,N_19503);
nand UO_1454 (O_1454,N_18909,N_18168);
or UO_1455 (O_1455,N_17083,N_18999);
nor UO_1456 (O_1456,N_17054,N_16811);
nand UO_1457 (O_1457,N_17667,N_17524);
xnor UO_1458 (O_1458,N_17329,N_16330);
or UO_1459 (O_1459,N_16857,N_16090);
and UO_1460 (O_1460,N_19404,N_18896);
nand UO_1461 (O_1461,N_16562,N_19393);
nand UO_1462 (O_1462,N_18874,N_18659);
and UO_1463 (O_1463,N_16760,N_16999);
nor UO_1464 (O_1464,N_16293,N_17832);
nor UO_1465 (O_1465,N_17475,N_19145);
and UO_1466 (O_1466,N_18963,N_16788);
xor UO_1467 (O_1467,N_18354,N_19828);
nand UO_1468 (O_1468,N_16715,N_18186);
and UO_1469 (O_1469,N_19597,N_18837);
nand UO_1470 (O_1470,N_17269,N_19794);
nand UO_1471 (O_1471,N_16066,N_16129);
xnor UO_1472 (O_1472,N_16678,N_16586);
nand UO_1473 (O_1473,N_17468,N_19609);
and UO_1474 (O_1474,N_17276,N_16597);
or UO_1475 (O_1475,N_16059,N_17578);
and UO_1476 (O_1476,N_18661,N_18652);
and UO_1477 (O_1477,N_16959,N_16209);
nor UO_1478 (O_1478,N_17959,N_18733);
xnor UO_1479 (O_1479,N_16997,N_16926);
and UO_1480 (O_1480,N_16978,N_19369);
and UO_1481 (O_1481,N_18984,N_17237);
nand UO_1482 (O_1482,N_17501,N_18459);
nor UO_1483 (O_1483,N_18049,N_19779);
xnor UO_1484 (O_1484,N_16015,N_18630);
nand UO_1485 (O_1485,N_19944,N_16829);
or UO_1486 (O_1486,N_18889,N_19123);
nand UO_1487 (O_1487,N_16808,N_18458);
and UO_1488 (O_1488,N_18826,N_17855);
nor UO_1489 (O_1489,N_16742,N_18407);
nor UO_1490 (O_1490,N_17844,N_17353);
nand UO_1491 (O_1491,N_18905,N_17425);
and UO_1492 (O_1492,N_16639,N_18419);
and UO_1493 (O_1493,N_19368,N_18692);
and UO_1494 (O_1494,N_16257,N_19968);
and UO_1495 (O_1495,N_17820,N_16809);
and UO_1496 (O_1496,N_16800,N_16136);
or UO_1497 (O_1497,N_18578,N_19203);
nor UO_1498 (O_1498,N_18006,N_19599);
or UO_1499 (O_1499,N_17452,N_16181);
nor UO_1500 (O_1500,N_16226,N_17243);
xor UO_1501 (O_1501,N_19885,N_18268);
nor UO_1502 (O_1502,N_16843,N_16240);
and UO_1503 (O_1503,N_19265,N_17843);
nor UO_1504 (O_1504,N_19169,N_19219);
nand UO_1505 (O_1505,N_19303,N_19384);
nor UO_1506 (O_1506,N_19911,N_18767);
nor UO_1507 (O_1507,N_17118,N_18577);
xor UO_1508 (O_1508,N_17227,N_18982);
and UO_1509 (O_1509,N_18843,N_19648);
nand UO_1510 (O_1510,N_19048,N_16872);
xnor UO_1511 (O_1511,N_16985,N_17047);
and UO_1512 (O_1512,N_16440,N_16525);
xnor UO_1513 (O_1513,N_19826,N_16564);
and UO_1514 (O_1514,N_18023,N_18471);
nor UO_1515 (O_1515,N_19202,N_19827);
and UO_1516 (O_1516,N_16470,N_17888);
and UO_1517 (O_1517,N_16003,N_19646);
and UO_1518 (O_1518,N_19242,N_17265);
or UO_1519 (O_1519,N_17308,N_19076);
or UO_1520 (O_1520,N_18417,N_17122);
nand UO_1521 (O_1521,N_16896,N_16148);
or UO_1522 (O_1522,N_17013,N_18493);
or UO_1523 (O_1523,N_18181,N_18244);
or UO_1524 (O_1524,N_16341,N_17740);
nor UO_1525 (O_1525,N_19294,N_19962);
xnor UO_1526 (O_1526,N_18125,N_18711);
xor UO_1527 (O_1527,N_17427,N_18726);
and UO_1528 (O_1528,N_18435,N_19502);
xnor UO_1529 (O_1529,N_16668,N_16218);
nand UO_1530 (O_1530,N_18528,N_17597);
and UO_1531 (O_1531,N_17486,N_17625);
xor UO_1532 (O_1532,N_19176,N_19345);
nand UO_1533 (O_1533,N_16546,N_17088);
or UO_1534 (O_1534,N_18931,N_18859);
nor UO_1535 (O_1535,N_18754,N_16433);
and UO_1536 (O_1536,N_17287,N_18453);
nor UO_1537 (O_1537,N_18037,N_18488);
and UO_1538 (O_1538,N_19119,N_17504);
and UO_1539 (O_1539,N_18515,N_17563);
nand UO_1540 (O_1540,N_17185,N_19606);
nand UO_1541 (O_1541,N_17947,N_16893);
nor UO_1542 (O_1542,N_16362,N_19397);
nor UO_1543 (O_1543,N_16435,N_17627);
nor UO_1544 (O_1544,N_19690,N_17782);
and UO_1545 (O_1545,N_18194,N_16802);
xor UO_1546 (O_1546,N_17318,N_18707);
nand UO_1547 (O_1547,N_17345,N_19688);
or UO_1548 (O_1548,N_18294,N_17440);
nand UO_1549 (O_1549,N_17218,N_16052);
or UO_1550 (O_1550,N_16934,N_16421);
or UO_1551 (O_1551,N_18622,N_18087);
or UO_1552 (O_1552,N_16862,N_19375);
nor UO_1553 (O_1553,N_17833,N_16831);
nor UO_1554 (O_1554,N_16787,N_19780);
or UO_1555 (O_1555,N_17739,N_19542);
nor UO_1556 (O_1556,N_17251,N_17209);
xnor UO_1557 (O_1557,N_16086,N_18990);
or UO_1558 (O_1558,N_19829,N_18490);
and UO_1559 (O_1559,N_19956,N_17200);
nand UO_1560 (O_1560,N_17602,N_18786);
and UO_1561 (O_1561,N_18595,N_18384);
nand UO_1562 (O_1562,N_16961,N_17594);
or UO_1563 (O_1563,N_16288,N_16432);
or UO_1564 (O_1564,N_17306,N_19745);
nor UO_1565 (O_1565,N_17128,N_18586);
xnor UO_1566 (O_1566,N_18715,N_19636);
nand UO_1567 (O_1567,N_18983,N_18450);
or UO_1568 (O_1568,N_17889,N_18827);
nor UO_1569 (O_1569,N_16617,N_18251);
nand UO_1570 (O_1570,N_19420,N_17559);
nor UO_1571 (O_1571,N_17717,N_17330);
nor UO_1572 (O_1572,N_19604,N_17955);
and UO_1573 (O_1573,N_18234,N_16920);
nor UO_1574 (O_1574,N_17708,N_17761);
and UO_1575 (O_1575,N_16105,N_19525);
nor UO_1576 (O_1576,N_18556,N_19726);
or UO_1577 (O_1577,N_16453,N_19097);
xnor UO_1578 (O_1578,N_18452,N_16408);
nor UO_1579 (O_1579,N_16201,N_19091);
and UO_1580 (O_1580,N_19130,N_18029);
or UO_1581 (O_1581,N_17703,N_16284);
or UO_1582 (O_1582,N_19002,N_18497);
or UO_1583 (O_1583,N_17706,N_17764);
nand UO_1584 (O_1584,N_16289,N_16532);
and UO_1585 (O_1585,N_19793,N_16106);
or UO_1586 (O_1586,N_17992,N_18789);
and UO_1587 (O_1587,N_17606,N_19339);
and UO_1588 (O_1588,N_16646,N_18158);
and UO_1589 (O_1589,N_16798,N_18410);
or UO_1590 (O_1590,N_17193,N_18232);
and UO_1591 (O_1591,N_17964,N_16458);
nor UO_1592 (O_1592,N_17134,N_18219);
or UO_1593 (O_1593,N_16102,N_19891);
or UO_1594 (O_1594,N_17564,N_16828);
nor UO_1595 (O_1595,N_16925,N_16426);
nor UO_1596 (O_1596,N_19778,N_19147);
nand UO_1597 (O_1597,N_19421,N_16669);
nand UO_1598 (O_1598,N_18882,N_18134);
nand UO_1599 (O_1599,N_16237,N_16631);
or UO_1600 (O_1600,N_16694,N_19767);
and UO_1601 (O_1601,N_17235,N_18228);
nor UO_1602 (O_1602,N_17777,N_16026);
or UO_1603 (O_1603,N_18358,N_19491);
nor UO_1604 (O_1604,N_16602,N_19923);
or UO_1605 (O_1605,N_16497,N_18819);
or UO_1606 (O_1606,N_16335,N_16094);
or UO_1607 (O_1607,N_17893,N_16104);
or UO_1608 (O_1608,N_17868,N_18526);
nand UO_1609 (O_1609,N_16269,N_17363);
xor UO_1610 (O_1610,N_19308,N_16834);
or UO_1611 (O_1611,N_19118,N_19001);
nor UO_1612 (O_1612,N_19765,N_18781);
nand UO_1613 (O_1613,N_17035,N_17278);
nand UO_1614 (O_1614,N_17892,N_16431);
nor UO_1615 (O_1615,N_16323,N_19910);
or UO_1616 (O_1616,N_17310,N_16060);
nand UO_1617 (O_1617,N_19574,N_17910);
nor UO_1618 (O_1618,N_19619,N_17954);
nor UO_1619 (O_1619,N_17879,N_16188);
nand UO_1620 (O_1620,N_16824,N_19075);
and UO_1621 (O_1621,N_19439,N_17670);
xnor UO_1622 (O_1622,N_16672,N_18499);
or UO_1623 (O_1623,N_17266,N_19040);
and UO_1624 (O_1624,N_17066,N_18571);
nand UO_1625 (O_1625,N_16469,N_17902);
nand UO_1626 (O_1626,N_18334,N_16405);
nor UO_1627 (O_1627,N_19394,N_16660);
nor UO_1628 (O_1628,N_18916,N_18847);
nand UO_1629 (O_1629,N_17847,N_17343);
nor UO_1630 (O_1630,N_16477,N_17304);
or UO_1631 (O_1631,N_16025,N_18475);
and UO_1632 (O_1632,N_18797,N_17943);
and UO_1633 (O_1633,N_16454,N_16420);
nor UO_1634 (O_1634,N_17818,N_17337);
nand UO_1635 (O_1635,N_17579,N_18591);
or UO_1636 (O_1636,N_17414,N_19572);
nor UO_1637 (O_1637,N_17175,N_19458);
or UO_1638 (O_1638,N_17571,N_17998);
and UO_1639 (O_1639,N_18881,N_19029);
nand UO_1640 (O_1640,N_17250,N_18039);
nand UO_1641 (O_1641,N_19681,N_18736);
or UO_1642 (O_1642,N_16685,N_16253);
and UO_1643 (O_1643,N_16236,N_18992);
or UO_1644 (O_1644,N_19290,N_17796);
and UO_1645 (O_1645,N_17267,N_17785);
nor UO_1646 (O_1646,N_16717,N_16819);
xor UO_1647 (O_1647,N_16008,N_18052);
and UO_1648 (O_1648,N_19761,N_17435);
xor UO_1649 (O_1649,N_16077,N_17009);
nor UO_1650 (O_1650,N_19134,N_16789);
nor UO_1651 (O_1651,N_18976,N_16551);
nor UO_1652 (O_1652,N_19501,N_16138);
and UO_1653 (O_1653,N_16412,N_19772);
nor UO_1654 (O_1654,N_19344,N_19951);
xor UO_1655 (O_1655,N_19244,N_19461);
nor UO_1656 (O_1656,N_16273,N_16165);
or UO_1657 (O_1657,N_19881,N_18003);
nor UO_1658 (O_1658,N_19341,N_16474);
xnor UO_1659 (O_1659,N_17941,N_16734);
or UO_1660 (O_1660,N_19909,N_18374);
or UO_1661 (O_1661,N_18409,N_16324);
and UO_1662 (O_1662,N_19526,N_19128);
nand UO_1663 (O_1663,N_16355,N_18501);
nor UO_1664 (O_1664,N_17753,N_16427);
nand UO_1665 (O_1665,N_17046,N_17914);
nor UO_1666 (O_1666,N_17074,N_18146);
and UO_1667 (O_1667,N_17755,N_19318);
nor UO_1668 (O_1668,N_16704,N_19698);
nor UO_1669 (O_1669,N_17075,N_18212);
nand UO_1670 (O_1670,N_18250,N_18731);
nand UO_1671 (O_1671,N_16570,N_16706);
and UO_1672 (O_1672,N_16415,N_18177);
nand UO_1673 (O_1673,N_17015,N_19789);
nor UO_1674 (O_1674,N_19508,N_18482);
nand UO_1675 (O_1675,N_18129,N_19485);
nand UO_1676 (O_1676,N_18159,N_19954);
xnor UO_1677 (O_1677,N_16342,N_17732);
and UO_1678 (O_1678,N_19022,N_17672);
xor UO_1679 (O_1679,N_16207,N_19117);
and UO_1680 (O_1680,N_17184,N_16984);
and UO_1681 (O_1681,N_17050,N_17172);
nand UO_1682 (O_1682,N_17726,N_18587);
or UO_1683 (O_1683,N_18941,N_16183);
nand UO_1684 (O_1684,N_16360,N_19035);
nor UO_1685 (O_1685,N_17423,N_17348);
nor UO_1686 (O_1686,N_16382,N_17033);
and UO_1687 (O_1687,N_19481,N_19113);
and UO_1688 (O_1688,N_17195,N_17967);
or UO_1689 (O_1689,N_17891,N_17313);
xnor UO_1690 (O_1690,N_16946,N_16827);
nand UO_1691 (O_1691,N_18647,N_16615);
xor UO_1692 (O_1692,N_16200,N_19095);
or UO_1693 (O_1693,N_18918,N_19200);
xnor UO_1694 (O_1694,N_18807,N_17999);
nand UO_1695 (O_1695,N_16344,N_18124);
xor UO_1696 (O_1696,N_17355,N_18249);
xnor UO_1697 (O_1697,N_16522,N_18287);
nor UO_1698 (O_1698,N_19021,N_17205);
or UO_1699 (O_1699,N_18709,N_18821);
and UO_1700 (O_1700,N_16260,N_18276);
or UO_1701 (O_1701,N_17628,N_17769);
and UO_1702 (O_1702,N_16913,N_17906);
and UO_1703 (O_1703,N_18880,N_18132);
or UO_1704 (O_1704,N_17545,N_16502);
nand UO_1705 (O_1705,N_16366,N_19933);
nor UO_1706 (O_1706,N_16791,N_16975);
and UO_1707 (O_1707,N_18904,N_18154);
and UO_1708 (O_1708,N_19288,N_17791);
and UO_1709 (O_1709,N_17372,N_16763);
nand UO_1710 (O_1710,N_16922,N_18946);
or UO_1711 (O_1711,N_19151,N_16853);
and UO_1712 (O_1712,N_16692,N_18988);
nand UO_1713 (O_1713,N_18645,N_18245);
or UO_1714 (O_1714,N_16194,N_16510);
xnor UO_1715 (O_1715,N_16885,N_19660);
or UO_1716 (O_1716,N_18958,N_19629);
nor UO_1717 (O_1717,N_16445,N_18514);
nand UO_1718 (O_1718,N_18597,N_17051);
xor UO_1719 (O_1719,N_19422,N_19638);
nor UO_1720 (O_1720,N_18197,N_17080);
or UO_1721 (O_1721,N_19259,N_16187);
nor UO_1722 (O_1722,N_18392,N_18604);
nor UO_1723 (O_1723,N_18838,N_18284);
nand UO_1724 (O_1724,N_18470,N_17812);
or UO_1725 (O_1725,N_18598,N_17404);
xnor UO_1726 (O_1726,N_17220,N_17886);
nand UO_1727 (O_1727,N_18939,N_16041);
or UO_1728 (O_1728,N_19038,N_17159);
xnor UO_1729 (O_1729,N_17067,N_16873);
xnor UO_1730 (O_1730,N_18741,N_18038);
nor UO_1731 (O_1731,N_18848,N_16491);
nand UO_1732 (O_1732,N_19090,N_16633);
nand UO_1733 (O_1733,N_18576,N_18567);
nor UO_1734 (O_1734,N_17042,N_17592);
or UO_1735 (O_1735,N_16818,N_16565);
xnor UO_1736 (O_1736,N_19221,N_17650);
or UO_1737 (O_1737,N_18760,N_16139);
xor UO_1738 (O_1738,N_16713,N_19010);
or UO_1739 (O_1739,N_18830,N_18609);
and UO_1740 (O_1740,N_18140,N_17953);
nand UO_1741 (O_1741,N_18015,N_16473);
and UO_1742 (O_1742,N_17380,N_19155);
or UO_1743 (O_1743,N_19258,N_17530);
nor UO_1744 (O_1744,N_19392,N_17401);
xnor UO_1745 (O_1745,N_19695,N_16847);
and UO_1746 (O_1746,N_18702,N_16902);
and UO_1747 (O_1747,N_17328,N_17189);
and UO_1748 (O_1748,N_19635,N_16049);
and UO_1749 (O_1749,N_18051,N_19433);
nand UO_1750 (O_1750,N_18585,N_19783);
xor UO_1751 (O_1751,N_18070,N_19831);
or UO_1752 (O_1752,N_18776,N_17745);
or UO_1753 (O_1753,N_17309,N_17878);
and UO_1754 (O_1754,N_16119,N_16051);
and UO_1755 (O_1755,N_16772,N_18074);
nor UO_1756 (O_1756,N_19953,N_16186);
or UO_1757 (O_1757,N_16463,N_17264);
or UO_1758 (O_1758,N_16888,N_17711);
nor UO_1759 (O_1759,N_17503,N_17804);
xnor UO_1760 (O_1760,N_17197,N_19717);
or UO_1761 (O_1761,N_19777,N_17262);
nand UO_1762 (O_1762,N_18274,N_19149);
nor UO_1763 (O_1763,N_19624,N_16103);
nor UO_1764 (O_1764,N_18280,N_19762);
nor UO_1765 (O_1765,N_18967,N_19547);
nand UO_1766 (O_1766,N_16437,N_19523);
and UO_1767 (O_1767,N_18877,N_18813);
and UO_1768 (O_1768,N_16392,N_17157);
and UO_1769 (O_1769,N_19049,N_16017);
nor UO_1770 (O_1770,N_19327,N_18867);
nand UO_1771 (O_1771,N_16938,N_16795);
nand UO_1772 (O_1772,N_17322,N_19066);
and UO_1773 (O_1773,N_16460,N_16037);
nand UO_1774 (O_1774,N_18701,N_16319);
nand UO_1775 (O_1775,N_18385,N_19583);
and UO_1776 (O_1776,N_18619,N_19346);
nor UO_1777 (O_1777,N_19297,N_18320);
nor UO_1778 (O_1778,N_19786,N_17060);
or UO_1779 (O_1779,N_18170,N_19328);
and UO_1780 (O_1780,N_18145,N_18745);
xor UO_1781 (O_1781,N_16513,N_16968);
or UO_1782 (O_1782,N_19797,N_18952);
nor UO_1783 (O_1783,N_17413,N_19044);
or UO_1784 (O_1784,N_16527,N_16246);
or UO_1785 (O_1785,N_16976,N_17649);
and UO_1786 (O_1786,N_18062,N_19349);
nand UO_1787 (O_1787,N_19197,N_18397);
nand UO_1788 (O_1788,N_16149,N_16735);
or UO_1789 (O_1789,N_17444,N_18404);
and UO_1790 (O_1790,N_19093,N_18525);
nand UO_1791 (O_1791,N_17107,N_16994);
xnor UO_1792 (O_1792,N_17674,N_16573);
or UO_1793 (O_1793,N_19081,N_16537);
and UO_1794 (O_1794,N_18387,N_18174);
nand UO_1795 (O_1795,N_18679,N_19114);
or UO_1796 (O_1796,N_19920,N_17177);
or UO_1797 (O_1797,N_19162,N_19846);
or UO_1798 (O_1798,N_19705,N_16732);
xnor UO_1799 (O_1799,N_17207,N_16871);
xor UO_1800 (O_1800,N_18669,N_16481);
nor UO_1801 (O_1801,N_18359,N_18491);
nor UO_1802 (O_1802,N_18119,N_17188);
or UO_1803 (O_1803,N_16612,N_19225);
nor UO_1804 (O_1804,N_18206,N_18369);
and UO_1805 (O_1805,N_18030,N_18076);
nor UO_1806 (O_1806,N_19618,N_18779);
nand UO_1807 (O_1807,N_19754,N_17351);
nand UO_1808 (O_1808,N_16131,N_17659);
nor UO_1809 (O_1809,N_18811,N_16501);
nand UO_1810 (O_1810,N_19307,N_18979);
or UO_1811 (O_1811,N_18259,N_16753);
or UO_1812 (O_1812,N_16399,N_17790);
nor UO_1813 (O_1813,N_18628,N_18288);
nand UO_1814 (O_1814,N_16930,N_16215);
and UO_1815 (O_1815,N_17370,N_16089);
xor UO_1816 (O_1816,N_18730,N_18216);
or UO_1817 (O_1817,N_17884,N_17780);
xnor UO_1818 (O_1818,N_16259,N_18102);
or UO_1819 (O_1819,N_19912,N_16830);
nor UO_1820 (O_1820,N_19565,N_17305);
nand UO_1821 (O_1821,N_18768,N_16908);
nor UO_1822 (O_1822,N_16636,N_16604);
nor UO_1823 (O_1823,N_16864,N_16556);
xnor UO_1824 (O_1824,N_19354,N_18185);
and UO_1825 (O_1825,N_19582,N_16331);
nand UO_1826 (O_1826,N_17873,N_17187);
nor UO_1827 (O_1827,N_18187,N_19268);
or UO_1828 (O_1828,N_16205,N_18836);
or UO_1829 (O_1829,N_18536,N_17704);
or UO_1830 (O_1830,N_18852,N_18466);
and UO_1831 (O_1831,N_18109,N_17115);
or UO_1832 (O_1832,N_19903,N_18869);
or UO_1833 (O_1833,N_19161,N_19356);
nor UO_1834 (O_1834,N_16733,N_18136);
nand UO_1835 (O_1835,N_18974,N_18343);
nand UO_1836 (O_1836,N_19476,N_16096);
nand UO_1837 (O_1837,N_16028,N_18618);
or UO_1838 (O_1838,N_18694,N_16374);
or UO_1839 (O_1839,N_16720,N_16407);
nand UO_1840 (O_1840,N_19395,N_17620);
nand UO_1841 (O_1841,N_17479,N_19154);
and UO_1842 (O_1842,N_19321,N_16134);
and UO_1843 (O_1843,N_19260,N_16133);
nor UO_1844 (O_1844,N_18978,N_18902);
nor UO_1845 (O_1845,N_18277,N_18560);
or UO_1846 (O_1846,N_18360,N_16801);
nand UO_1847 (O_1847,N_18510,N_16840);
or UO_1848 (O_1848,N_16835,N_18071);
nand UO_1849 (O_1849,N_17585,N_19748);
or UO_1850 (O_1850,N_16069,N_17958);
nand UO_1851 (O_1851,N_17378,N_16696);
or UO_1852 (O_1852,N_17392,N_19915);
nand UO_1853 (O_1853,N_19554,N_16560);
and UO_1854 (O_1854,N_16576,N_18696);
nor UO_1855 (O_1855,N_16779,N_18638);
nand UO_1856 (O_1856,N_16971,N_16206);
nor UO_1857 (O_1857,N_18681,N_18500);
and UO_1858 (O_1858,N_17936,N_17996);
and UO_1859 (O_1859,N_16663,N_17323);
nand UO_1860 (O_1860,N_17129,N_19724);
xnor UO_1861 (O_1861,N_19295,N_16048);
nor UO_1862 (O_1862,N_17538,N_17883);
xor UO_1863 (O_1863,N_18111,N_17260);
nand UO_1864 (O_1864,N_18968,N_19306);
and UO_1865 (O_1865,N_19201,N_16530);
xor UO_1866 (O_1866,N_18657,N_17173);
or UO_1867 (O_1867,N_17467,N_19171);
nor UO_1868 (O_1868,N_17402,N_18829);
or UO_1869 (O_1869,N_18017,N_18203);
or UO_1870 (O_1870,N_18461,N_16101);
or UO_1871 (O_1871,N_17369,N_17282);
or UO_1872 (O_1872,N_17422,N_19494);
nor UO_1873 (O_1873,N_16569,N_16790);
nor UO_1874 (O_1874,N_18035,N_17523);
nor UO_1875 (O_1875,N_18763,N_16630);
nor UO_1876 (O_1876,N_19830,N_16045);
nand UO_1877 (O_1877,N_18667,N_17852);
nor UO_1878 (O_1878,N_19598,N_16880);
and UO_1879 (O_1879,N_17662,N_18962);
xor UO_1880 (O_1880,N_17049,N_19311);
nand UO_1881 (O_1881,N_16868,N_19504);
and UO_1882 (O_1882,N_16353,N_18642);
nand UO_1883 (O_1883,N_18066,N_18890);
or UO_1884 (O_1884,N_16001,N_18790);
or UO_1885 (O_1885,N_17151,N_18517);
and UO_1886 (O_1886,N_19714,N_19804);
nor UO_1887 (O_1887,N_17803,N_19551);
or UO_1888 (O_1888,N_16703,N_18264);
nor UO_1889 (O_1889,N_18465,N_18868);
and UO_1890 (O_1890,N_17059,N_17924);
nor UO_1891 (O_1891,N_17814,N_17632);
nand UO_1892 (O_1892,N_18831,N_19680);
and UO_1893 (O_1893,N_19707,N_19324);
nand UO_1894 (O_1894,N_18231,N_17244);
and UO_1895 (O_1895,N_18131,N_16954);
or UO_1896 (O_1896,N_17335,N_19323);
and UO_1897 (O_1897,N_17490,N_16887);
nor UO_1898 (O_1898,N_19059,N_18922);
or UO_1899 (O_1899,N_17466,N_18000);
or UO_1900 (O_1900,N_19101,N_19760);
nor UO_1901 (O_1901,N_17945,N_19759);
nor UO_1902 (O_1902,N_17154,N_16874);
xnor UO_1903 (O_1903,N_19449,N_19156);
nand UO_1904 (O_1904,N_17203,N_17496);
or UO_1905 (O_1905,N_18148,N_16674);
xnor UO_1906 (O_1906,N_18980,N_16977);
nor UO_1907 (O_1907,N_19825,N_19240);
nor UO_1908 (O_1908,N_16021,N_18270);
xor UO_1909 (O_1909,N_19863,N_19431);
and UO_1910 (O_1910,N_19382,N_17815);
nand UO_1911 (O_1911,N_17148,N_18220);
and UO_1912 (O_1912,N_16776,N_18025);
and UO_1913 (O_1913,N_19607,N_17434);
and UO_1914 (O_1914,N_17398,N_19402);
nand UO_1915 (O_1915,N_16158,N_19267);
or UO_1916 (O_1916,N_19608,N_18892);
nor UO_1917 (O_1917,N_16070,N_17326);
or UO_1918 (O_1918,N_17894,N_16027);
and UO_1919 (O_1919,N_16682,N_18687);
nor UO_1920 (O_1920,N_18456,N_17356);
or UO_1921 (O_1921,N_18356,N_19516);
and UO_1922 (O_1922,N_16571,N_19587);
nand UO_1923 (O_1923,N_16231,N_16247);
and UO_1924 (O_1924,N_18222,N_18518);
nor UO_1925 (O_1925,N_18118,N_16952);
or UO_1926 (O_1926,N_18762,N_17641);
nor UO_1927 (O_1927,N_18599,N_16702);
or UO_1928 (O_1928,N_16919,N_16958);
nand UO_1929 (O_1929,N_16989,N_17723);
nand UO_1930 (O_1930,N_19868,N_18255);
nand UO_1931 (O_1931,N_16533,N_16641);
or UO_1932 (O_1932,N_18098,N_17800);
or UO_1933 (O_1933,N_18623,N_18814);
nor UO_1934 (O_1934,N_17710,N_18205);
nand UO_1935 (O_1935,N_19538,N_17793);
nand UO_1936 (O_1936,N_17857,N_17449);
nor UO_1937 (O_1937,N_16877,N_17204);
nor UO_1938 (O_1938,N_18673,N_17932);
nand UO_1939 (O_1939,N_16539,N_17261);
and UO_1940 (O_1940,N_18105,N_18803);
xor UO_1941 (O_1941,N_16650,N_19378);
nor UO_1942 (O_1942,N_18658,N_17760);
or UO_1943 (O_1943,N_18607,N_18215);
nand UO_1944 (O_1944,N_18229,N_18653);
nand UO_1945 (O_1945,N_18108,N_18895);
nand UO_1946 (O_1946,N_17616,N_16621);
nor UO_1947 (O_1947,N_19615,N_18703);
or UO_1948 (O_1948,N_18740,N_19595);
and UO_1949 (O_1949,N_18271,N_18543);
nand UO_1950 (O_1950,N_19822,N_19813);
nor UO_1951 (O_1951,N_18775,N_19967);
and UO_1952 (O_1952,N_18551,N_18766);
nand UO_1953 (O_1953,N_17930,N_19673);
nor UO_1954 (O_1954,N_18447,N_16109);
xnor UO_1955 (O_1955,N_18656,N_19733);
nand UO_1956 (O_1956,N_18269,N_19837);
nor UO_1957 (O_1957,N_16055,N_16451);
or UO_1958 (O_1958,N_16444,N_19120);
nor UO_1959 (O_1959,N_19616,N_19317);
nor UO_1960 (O_1960,N_17448,N_16765);
or UO_1961 (O_1961,N_16710,N_18602);
nor UO_1962 (O_1962,N_18012,N_17395);
nand UO_1963 (O_1963,N_17221,N_16085);
nand UO_1964 (O_1964,N_17294,N_17455);
and UO_1965 (O_1965,N_19057,N_16083);
nor UO_1966 (O_1966,N_18044,N_17547);
xnor UO_1967 (O_1967,N_17756,N_16376);
nand UO_1968 (O_1968,N_17436,N_16599);
nor UO_1969 (O_1969,N_17219,N_16935);
nor UO_1970 (O_1970,N_17573,N_17986);
or UO_1971 (O_1971,N_16966,N_19455);
and UO_1972 (O_1972,N_18031,N_17558);
and UO_1973 (O_1973,N_19623,N_17023);
nand UO_1974 (O_1974,N_18122,N_19170);
or UO_1975 (O_1975,N_17252,N_18165);
nor UO_1976 (O_1976,N_17429,N_17877);
or UO_1977 (O_1977,N_19875,N_16991);
or UO_1978 (O_1978,N_18564,N_16816);
nor UO_1979 (O_1979,N_16552,N_19446);
nor UO_1980 (O_1980,N_16688,N_18529);
or UO_1981 (O_1981,N_16516,N_19050);
xor UO_1982 (O_1982,N_16168,N_16721);
nor UO_1983 (O_1983,N_18828,N_16423);
nor UO_1984 (O_1984,N_19807,N_19425);
xnor UO_1985 (O_1985,N_18091,N_18286);
nor UO_1986 (O_1986,N_17948,N_17991);
and UO_1987 (O_1987,N_16182,N_19999);
or UO_1988 (O_1988,N_18121,N_19256);
and UO_1989 (O_1989,N_16254,N_16962);
and UO_1990 (O_1990,N_19285,N_17520);
nand UO_1991 (O_1991,N_17152,N_19241);
nor UO_1992 (O_1992,N_16155,N_19741);
or UO_1993 (O_1993,N_18865,N_17557);
and UO_1994 (O_1994,N_19143,N_19524);
nand UO_1995 (O_1995,N_19187,N_17863);
or UO_1996 (O_1996,N_18063,N_18292);
xnor UO_1997 (O_1997,N_16093,N_19791);
and UO_1998 (O_1998,N_19532,N_18823);
and UO_1999 (O_1999,N_16098,N_16851);
or UO_2000 (O_2000,N_16358,N_19132);
nor UO_2001 (O_2001,N_16576,N_19651);
xnor UO_2002 (O_2002,N_19186,N_17002);
and UO_2003 (O_2003,N_19421,N_16613);
nand UO_2004 (O_2004,N_18104,N_16287);
or UO_2005 (O_2005,N_19753,N_16062);
and UO_2006 (O_2006,N_19198,N_19933);
and UO_2007 (O_2007,N_17564,N_17037);
or UO_2008 (O_2008,N_16188,N_18095);
nand UO_2009 (O_2009,N_16660,N_16739);
xnor UO_2010 (O_2010,N_16232,N_18164);
and UO_2011 (O_2011,N_18748,N_16012);
and UO_2012 (O_2012,N_16405,N_19444);
nor UO_2013 (O_2013,N_19736,N_19419);
and UO_2014 (O_2014,N_19674,N_17459);
or UO_2015 (O_2015,N_19303,N_16631);
nor UO_2016 (O_2016,N_18713,N_17928);
nand UO_2017 (O_2017,N_16065,N_19338);
nand UO_2018 (O_2018,N_17005,N_17609);
xnor UO_2019 (O_2019,N_19747,N_17512);
xor UO_2020 (O_2020,N_19523,N_16968);
xnor UO_2021 (O_2021,N_18391,N_18151);
nor UO_2022 (O_2022,N_18984,N_17845);
and UO_2023 (O_2023,N_19781,N_18869);
nand UO_2024 (O_2024,N_17025,N_18853);
nor UO_2025 (O_2025,N_18632,N_19219);
or UO_2026 (O_2026,N_18760,N_18407);
and UO_2027 (O_2027,N_16961,N_16923);
xnor UO_2028 (O_2028,N_18571,N_16923);
and UO_2029 (O_2029,N_19965,N_19569);
nand UO_2030 (O_2030,N_16559,N_17661);
and UO_2031 (O_2031,N_16873,N_16901);
xor UO_2032 (O_2032,N_16069,N_19136);
nand UO_2033 (O_2033,N_18259,N_16152);
and UO_2034 (O_2034,N_16563,N_18242);
and UO_2035 (O_2035,N_18237,N_19434);
nand UO_2036 (O_2036,N_16031,N_18153);
or UO_2037 (O_2037,N_18486,N_16871);
and UO_2038 (O_2038,N_19021,N_16644);
and UO_2039 (O_2039,N_18481,N_19920);
or UO_2040 (O_2040,N_19934,N_17028);
nand UO_2041 (O_2041,N_18000,N_17002);
and UO_2042 (O_2042,N_18540,N_19819);
nand UO_2043 (O_2043,N_19292,N_16967);
xnor UO_2044 (O_2044,N_16359,N_19989);
nor UO_2045 (O_2045,N_17260,N_18168);
or UO_2046 (O_2046,N_17589,N_18174);
nor UO_2047 (O_2047,N_17129,N_16410);
nand UO_2048 (O_2048,N_17387,N_17865);
nor UO_2049 (O_2049,N_17091,N_18882);
nor UO_2050 (O_2050,N_16324,N_18650);
xor UO_2051 (O_2051,N_16722,N_18839);
or UO_2052 (O_2052,N_17173,N_19396);
and UO_2053 (O_2053,N_17453,N_16323);
nor UO_2054 (O_2054,N_17715,N_16639);
nor UO_2055 (O_2055,N_19685,N_17402);
xor UO_2056 (O_2056,N_17643,N_18123);
nor UO_2057 (O_2057,N_18915,N_18706);
xnor UO_2058 (O_2058,N_19872,N_16132);
or UO_2059 (O_2059,N_16314,N_16903);
nand UO_2060 (O_2060,N_17935,N_19210);
nor UO_2061 (O_2061,N_17641,N_19407);
nor UO_2062 (O_2062,N_18864,N_17453);
or UO_2063 (O_2063,N_17117,N_17076);
nor UO_2064 (O_2064,N_18771,N_19922);
or UO_2065 (O_2065,N_17575,N_17532);
and UO_2066 (O_2066,N_18285,N_18077);
and UO_2067 (O_2067,N_19866,N_17119);
and UO_2068 (O_2068,N_18654,N_17410);
or UO_2069 (O_2069,N_17715,N_18845);
and UO_2070 (O_2070,N_18825,N_17932);
or UO_2071 (O_2071,N_19020,N_17399);
and UO_2072 (O_2072,N_18187,N_17505);
or UO_2073 (O_2073,N_18201,N_16233);
nand UO_2074 (O_2074,N_19819,N_17636);
nand UO_2075 (O_2075,N_16286,N_18557);
and UO_2076 (O_2076,N_16065,N_16986);
and UO_2077 (O_2077,N_17049,N_19874);
nand UO_2078 (O_2078,N_16644,N_16347);
xor UO_2079 (O_2079,N_17656,N_18882);
nor UO_2080 (O_2080,N_18943,N_18761);
and UO_2081 (O_2081,N_19047,N_18713);
or UO_2082 (O_2082,N_18513,N_16778);
or UO_2083 (O_2083,N_17596,N_16194);
nor UO_2084 (O_2084,N_16182,N_19016);
nor UO_2085 (O_2085,N_18956,N_16023);
and UO_2086 (O_2086,N_17520,N_16671);
or UO_2087 (O_2087,N_16295,N_18386);
nand UO_2088 (O_2088,N_16211,N_16673);
or UO_2089 (O_2089,N_17586,N_17222);
nor UO_2090 (O_2090,N_16155,N_17315);
and UO_2091 (O_2091,N_18696,N_16997);
and UO_2092 (O_2092,N_17885,N_16563);
nor UO_2093 (O_2093,N_18502,N_17827);
nand UO_2094 (O_2094,N_16981,N_16904);
nor UO_2095 (O_2095,N_16090,N_18979);
and UO_2096 (O_2096,N_16866,N_16448);
and UO_2097 (O_2097,N_19144,N_19870);
nor UO_2098 (O_2098,N_16636,N_19209);
nor UO_2099 (O_2099,N_17803,N_18811);
and UO_2100 (O_2100,N_17368,N_17546);
or UO_2101 (O_2101,N_17286,N_19500);
nor UO_2102 (O_2102,N_17588,N_18963);
and UO_2103 (O_2103,N_19699,N_18823);
nand UO_2104 (O_2104,N_19862,N_17552);
and UO_2105 (O_2105,N_18194,N_18843);
nand UO_2106 (O_2106,N_18519,N_18131);
and UO_2107 (O_2107,N_18995,N_16567);
or UO_2108 (O_2108,N_19705,N_19872);
or UO_2109 (O_2109,N_19828,N_17709);
and UO_2110 (O_2110,N_19742,N_19052);
nor UO_2111 (O_2111,N_17932,N_19568);
or UO_2112 (O_2112,N_19996,N_16902);
nor UO_2113 (O_2113,N_16491,N_16366);
nand UO_2114 (O_2114,N_18739,N_16575);
and UO_2115 (O_2115,N_17157,N_17775);
nand UO_2116 (O_2116,N_16341,N_17631);
or UO_2117 (O_2117,N_18536,N_17272);
or UO_2118 (O_2118,N_19626,N_18216);
nor UO_2119 (O_2119,N_17932,N_16603);
or UO_2120 (O_2120,N_18665,N_16890);
and UO_2121 (O_2121,N_18620,N_17585);
xor UO_2122 (O_2122,N_18088,N_19279);
or UO_2123 (O_2123,N_16705,N_19960);
nand UO_2124 (O_2124,N_19889,N_16343);
or UO_2125 (O_2125,N_17700,N_16585);
and UO_2126 (O_2126,N_18808,N_17779);
nor UO_2127 (O_2127,N_19948,N_19344);
and UO_2128 (O_2128,N_17605,N_18213);
or UO_2129 (O_2129,N_16992,N_17850);
nand UO_2130 (O_2130,N_17050,N_19993);
or UO_2131 (O_2131,N_17364,N_19975);
and UO_2132 (O_2132,N_16354,N_19935);
and UO_2133 (O_2133,N_18286,N_18083);
nand UO_2134 (O_2134,N_17701,N_18408);
and UO_2135 (O_2135,N_18331,N_17346);
and UO_2136 (O_2136,N_17572,N_17594);
xnor UO_2137 (O_2137,N_16861,N_16065);
or UO_2138 (O_2138,N_17243,N_19459);
nand UO_2139 (O_2139,N_16986,N_18791);
or UO_2140 (O_2140,N_18058,N_19656);
nor UO_2141 (O_2141,N_16294,N_16455);
nand UO_2142 (O_2142,N_19188,N_16644);
or UO_2143 (O_2143,N_17466,N_16896);
and UO_2144 (O_2144,N_19903,N_16089);
nand UO_2145 (O_2145,N_18395,N_19316);
nand UO_2146 (O_2146,N_18119,N_16054);
or UO_2147 (O_2147,N_16331,N_17592);
and UO_2148 (O_2148,N_17977,N_17051);
or UO_2149 (O_2149,N_18781,N_18210);
or UO_2150 (O_2150,N_18423,N_19916);
nor UO_2151 (O_2151,N_19884,N_19105);
and UO_2152 (O_2152,N_16967,N_16106);
and UO_2153 (O_2153,N_19092,N_18170);
nand UO_2154 (O_2154,N_17170,N_17059);
and UO_2155 (O_2155,N_16657,N_17396);
nor UO_2156 (O_2156,N_16941,N_16728);
and UO_2157 (O_2157,N_17616,N_16600);
xor UO_2158 (O_2158,N_16863,N_17667);
nor UO_2159 (O_2159,N_17860,N_17788);
or UO_2160 (O_2160,N_16602,N_16776);
xor UO_2161 (O_2161,N_18793,N_17733);
and UO_2162 (O_2162,N_17049,N_17148);
and UO_2163 (O_2163,N_17009,N_18709);
or UO_2164 (O_2164,N_17801,N_18579);
and UO_2165 (O_2165,N_19266,N_17081);
xor UO_2166 (O_2166,N_19339,N_17159);
or UO_2167 (O_2167,N_16008,N_19107);
and UO_2168 (O_2168,N_17208,N_19196);
and UO_2169 (O_2169,N_17890,N_19873);
xor UO_2170 (O_2170,N_18192,N_18085);
nor UO_2171 (O_2171,N_17657,N_16139);
or UO_2172 (O_2172,N_18582,N_16370);
nand UO_2173 (O_2173,N_16447,N_19809);
or UO_2174 (O_2174,N_16577,N_19989);
or UO_2175 (O_2175,N_19665,N_18688);
nor UO_2176 (O_2176,N_16438,N_16678);
and UO_2177 (O_2177,N_16316,N_17741);
nand UO_2178 (O_2178,N_19700,N_18305);
nor UO_2179 (O_2179,N_19006,N_19430);
nand UO_2180 (O_2180,N_18656,N_18107);
xnor UO_2181 (O_2181,N_19338,N_19839);
or UO_2182 (O_2182,N_16369,N_18425);
xor UO_2183 (O_2183,N_17384,N_19349);
or UO_2184 (O_2184,N_18036,N_16148);
nor UO_2185 (O_2185,N_16962,N_18358);
nor UO_2186 (O_2186,N_19298,N_19725);
or UO_2187 (O_2187,N_19831,N_17667);
and UO_2188 (O_2188,N_19041,N_16568);
and UO_2189 (O_2189,N_19902,N_16094);
and UO_2190 (O_2190,N_18945,N_17105);
or UO_2191 (O_2191,N_17046,N_18573);
xnor UO_2192 (O_2192,N_19591,N_17705);
and UO_2193 (O_2193,N_17183,N_17216);
or UO_2194 (O_2194,N_18474,N_17229);
xnor UO_2195 (O_2195,N_18687,N_16368);
and UO_2196 (O_2196,N_19339,N_17823);
and UO_2197 (O_2197,N_18779,N_16238);
and UO_2198 (O_2198,N_19076,N_17095);
nor UO_2199 (O_2199,N_19056,N_19285);
or UO_2200 (O_2200,N_18714,N_16517);
and UO_2201 (O_2201,N_16586,N_16812);
and UO_2202 (O_2202,N_18447,N_19316);
or UO_2203 (O_2203,N_17024,N_17595);
nand UO_2204 (O_2204,N_19045,N_19565);
nor UO_2205 (O_2205,N_17514,N_17769);
nor UO_2206 (O_2206,N_17344,N_19364);
nand UO_2207 (O_2207,N_17576,N_19054);
and UO_2208 (O_2208,N_19327,N_18765);
nand UO_2209 (O_2209,N_17164,N_18694);
or UO_2210 (O_2210,N_17966,N_17432);
or UO_2211 (O_2211,N_19997,N_19323);
nand UO_2212 (O_2212,N_18070,N_18173);
nand UO_2213 (O_2213,N_17235,N_17402);
or UO_2214 (O_2214,N_17578,N_18680);
nor UO_2215 (O_2215,N_17621,N_16372);
or UO_2216 (O_2216,N_19955,N_18032);
or UO_2217 (O_2217,N_16679,N_18641);
and UO_2218 (O_2218,N_18700,N_16286);
or UO_2219 (O_2219,N_17059,N_19510);
or UO_2220 (O_2220,N_17360,N_19462);
nand UO_2221 (O_2221,N_18467,N_16764);
or UO_2222 (O_2222,N_16818,N_17279);
and UO_2223 (O_2223,N_19529,N_18426);
nand UO_2224 (O_2224,N_19975,N_16777);
nor UO_2225 (O_2225,N_19465,N_19044);
nand UO_2226 (O_2226,N_19269,N_16749);
nand UO_2227 (O_2227,N_19630,N_19357);
xnor UO_2228 (O_2228,N_18360,N_17890);
xor UO_2229 (O_2229,N_16472,N_19005);
nor UO_2230 (O_2230,N_19657,N_18336);
xnor UO_2231 (O_2231,N_17923,N_19153);
or UO_2232 (O_2232,N_16816,N_19263);
nand UO_2233 (O_2233,N_19728,N_19270);
nor UO_2234 (O_2234,N_17598,N_19878);
nand UO_2235 (O_2235,N_18188,N_19265);
and UO_2236 (O_2236,N_18881,N_18989);
nor UO_2237 (O_2237,N_19732,N_17038);
and UO_2238 (O_2238,N_18529,N_16731);
xor UO_2239 (O_2239,N_19871,N_17280);
or UO_2240 (O_2240,N_16657,N_16524);
nor UO_2241 (O_2241,N_18430,N_18335);
and UO_2242 (O_2242,N_17930,N_17013);
and UO_2243 (O_2243,N_16514,N_18145);
nor UO_2244 (O_2244,N_18582,N_17008);
nand UO_2245 (O_2245,N_18372,N_17529);
or UO_2246 (O_2246,N_18386,N_16135);
or UO_2247 (O_2247,N_19737,N_16468);
and UO_2248 (O_2248,N_17705,N_19414);
nor UO_2249 (O_2249,N_16179,N_17264);
nand UO_2250 (O_2250,N_17487,N_18866);
and UO_2251 (O_2251,N_18001,N_19351);
and UO_2252 (O_2252,N_18011,N_19637);
nand UO_2253 (O_2253,N_16291,N_17265);
and UO_2254 (O_2254,N_16743,N_19858);
nand UO_2255 (O_2255,N_16462,N_18552);
nor UO_2256 (O_2256,N_16032,N_19592);
nor UO_2257 (O_2257,N_16348,N_16029);
nand UO_2258 (O_2258,N_19937,N_19204);
and UO_2259 (O_2259,N_17113,N_17528);
or UO_2260 (O_2260,N_16034,N_18103);
xor UO_2261 (O_2261,N_18383,N_18235);
or UO_2262 (O_2262,N_16942,N_16265);
or UO_2263 (O_2263,N_18794,N_17914);
or UO_2264 (O_2264,N_16930,N_16505);
nor UO_2265 (O_2265,N_17509,N_17024);
or UO_2266 (O_2266,N_19749,N_19508);
nand UO_2267 (O_2267,N_19780,N_17596);
nand UO_2268 (O_2268,N_17689,N_16773);
or UO_2269 (O_2269,N_17853,N_17447);
xor UO_2270 (O_2270,N_16056,N_19998);
or UO_2271 (O_2271,N_19621,N_19637);
and UO_2272 (O_2272,N_16016,N_19636);
nor UO_2273 (O_2273,N_19265,N_16131);
and UO_2274 (O_2274,N_16256,N_18287);
and UO_2275 (O_2275,N_17356,N_18501);
or UO_2276 (O_2276,N_16433,N_17518);
xor UO_2277 (O_2277,N_17994,N_16555);
nor UO_2278 (O_2278,N_16007,N_16849);
or UO_2279 (O_2279,N_16378,N_19869);
or UO_2280 (O_2280,N_19745,N_18026);
nor UO_2281 (O_2281,N_18511,N_16916);
nor UO_2282 (O_2282,N_17349,N_17965);
and UO_2283 (O_2283,N_18735,N_19396);
and UO_2284 (O_2284,N_19913,N_17872);
or UO_2285 (O_2285,N_18882,N_18423);
or UO_2286 (O_2286,N_17717,N_16811);
nand UO_2287 (O_2287,N_19116,N_16059);
or UO_2288 (O_2288,N_16000,N_16643);
nand UO_2289 (O_2289,N_17846,N_17936);
xnor UO_2290 (O_2290,N_18352,N_16985);
or UO_2291 (O_2291,N_19162,N_16819);
or UO_2292 (O_2292,N_17403,N_19303);
and UO_2293 (O_2293,N_17065,N_17763);
nor UO_2294 (O_2294,N_19454,N_18786);
nor UO_2295 (O_2295,N_18448,N_16680);
nor UO_2296 (O_2296,N_19383,N_18027);
nor UO_2297 (O_2297,N_16515,N_17561);
and UO_2298 (O_2298,N_19595,N_17862);
and UO_2299 (O_2299,N_16663,N_17758);
nor UO_2300 (O_2300,N_17213,N_16765);
nor UO_2301 (O_2301,N_16089,N_17119);
or UO_2302 (O_2302,N_16170,N_16548);
and UO_2303 (O_2303,N_19343,N_19309);
nor UO_2304 (O_2304,N_17704,N_17747);
nor UO_2305 (O_2305,N_16459,N_17735);
or UO_2306 (O_2306,N_18694,N_18191);
nor UO_2307 (O_2307,N_16694,N_18103);
and UO_2308 (O_2308,N_16480,N_18576);
and UO_2309 (O_2309,N_17322,N_17142);
and UO_2310 (O_2310,N_19860,N_18144);
and UO_2311 (O_2311,N_18726,N_17949);
nor UO_2312 (O_2312,N_19112,N_19541);
and UO_2313 (O_2313,N_17674,N_19237);
and UO_2314 (O_2314,N_19054,N_16340);
xnor UO_2315 (O_2315,N_19524,N_19802);
or UO_2316 (O_2316,N_19274,N_19427);
or UO_2317 (O_2317,N_19036,N_18816);
nor UO_2318 (O_2318,N_19878,N_16135);
or UO_2319 (O_2319,N_17044,N_16667);
nor UO_2320 (O_2320,N_17244,N_18473);
nand UO_2321 (O_2321,N_17618,N_16378);
nor UO_2322 (O_2322,N_19112,N_17758);
and UO_2323 (O_2323,N_18306,N_18642);
and UO_2324 (O_2324,N_18160,N_16101);
xnor UO_2325 (O_2325,N_18625,N_16721);
or UO_2326 (O_2326,N_19267,N_17269);
and UO_2327 (O_2327,N_18356,N_17870);
and UO_2328 (O_2328,N_16078,N_17857);
nor UO_2329 (O_2329,N_17442,N_17467);
or UO_2330 (O_2330,N_17279,N_19032);
nor UO_2331 (O_2331,N_19275,N_16860);
or UO_2332 (O_2332,N_16265,N_16638);
or UO_2333 (O_2333,N_19344,N_17453);
nand UO_2334 (O_2334,N_18959,N_16159);
or UO_2335 (O_2335,N_18551,N_18453);
nor UO_2336 (O_2336,N_17042,N_17703);
and UO_2337 (O_2337,N_19166,N_18223);
nor UO_2338 (O_2338,N_17904,N_19332);
and UO_2339 (O_2339,N_19842,N_17431);
xnor UO_2340 (O_2340,N_17110,N_18847);
and UO_2341 (O_2341,N_17108,N_18661);
xor UO_2342 (O_2342,N_18686,N_19428);
nor UO_2343 (O_2343,N_16794,N_18272);
or UO_2344 (O_2344,N_19579,N_19922);
nor UO_2345 (O_2345,N_19287,N_16969);
nor UO_2346 (O_2346,N_17400,N_18549);
nor UO_2347 (O_2347,N_18663,N_17334);
and UO_2348 (O_2348,N_17770,N_16476);
nand UO_2349 (O_2349,N_19393,N_18155);
or UO_2350 (O_2350,N_18546,N_17344);
and UO_2351 (O_2351,N_18510,N_19591);
xnor UO_2352 (O_2352,N_18143,N_16487);
and UO_2353 (O_2353,N_18259,N_19393);
and UO_2354 (O_2354,N_17821,N_19066);
nor UO_2355 (O_2355,N_19273,N_16021);
or UO_2356 (O_2356,N_16454,N_16423);
or UO_2357 (O_2357,N_16910,N_17599);
nor UO_2358 (O_2358,N_18254,N_19669);
nand UO_2359 (O_2359,N_17782,N_19806);
or UO_2360 (O_2360,N_19193,N_18996);
or UO_2361 (O_2361,N_16385,N_17779);
and UO_2362 (O_2362,N_19917,N_16618);
xnor UO_2363 (O_2363,N_19067,N_18424);
xor UO_2364 (O_2364,N_17735,N_18966);
and UO_2365 (O_2365,N_17200,N_18183);
nor UO_2366 (O_2366,N_18568,N_17539);
nor UO_2367 (O_2367,N_18384,N_19099);
nor UO_2368 (O_2368,N_17057,N_17897);
or UO_2369 (O_2369,N_17837,N_16535);
and UO_2370 (O_2370,N_19739,N_16767);
nor UO_2371 (O_2371,N_17746,N_19850);
and UO_2372 (O_2372,N_19081,N_17712);
and UO_2373 (O_2373,N_17743,N_16277);
and UO_2374 (O_2374,N_16725,N_16078);
nand UO_2375 (O_2375,N_19023,N_17406);
and UO_2376 (O_2376,N_18954,N_18069);
and UO_2377 (O_2377,N_17901,N_16387);
nor UO_2378 (O_2378,N_18129,N_19978);
xnor UO_2379 (O_2379,N_18333,N_16341);
or UO_2380 (O_2380,N_18059,N_18464);
nand UO_2381 (O_2381,N_18136,N_17472);
or UO_2382 (O_2382,N_17940,N_18631);
nand UO_2383 (O_2383,N_16423,N_17562);
nor UO_2384 (O_2384,N_17227,N_18385);
and UO_2385 (O_2385,N_17550,N_18641);
nand UO_2386 (O_2386,N_18238,N_19684);
or UO_2387 (O_2387,N_18003,N_17297);
and UO_2388 (O_2388,N_18744,N_17462);
nand UO_2389 (O_2389,N_19272,N_16925);
nand UO_2390 (O_2390,N_17376,N_19161);
or UO_2391 (O_2391,N_18730,N_17640);
nor UO_2392 (O_2392,N_17958,N_18378);
nand UO_2393 (O_2393,N_17641,N_18988);
nor UO_2394 (O_2394,N_19647,N_18206);
nor UO_2395 (O_2395,N_17008,N_19061);
or UO_2396 (O_2396,N_16472,N_17346);
xnor UO_2397 (O_2397,N_19950,N_18556);
and UO_2398 (O_2398,N_18629,N_17070);
nand UO_2399 (O_2399,N_16766,N_19850);
or UO_2400 (O_2400,N_19295,N_19151);
nand UO_2401 (O_2401,N_16082,N_17281);
or UO_2402 (O_2402,N_18073,N_16097);
and UO_2403 (O_2403,N_19014,N_19390);
nand UO_2404 (O_2404,N_19478,N_18489);
and UO_2405 (O_2405,N_16486,N_19819);
xor UO_2406 (O_2406,N_17689,N_19584);
or UO_2407 (O_2407,N_18137,N_19311);
xor UO_2408 (O_2408,N_16162,N_16588);
nor UO_2409 (O_2409,N_17476,N_19975);
and UO_2410 (O_2410,N_18113,N_19774);
or UO_2411 (O_2411,N_19117,N_17450);
nand UO_2412 (O_2412,N_17103,N_19659);
or UO_2413 (O_2413,N_17554,N_19123);
or UO_2414 (O_2414,N_17733,N_19320);
nor UO_2415 (O_2415,N_16751,N_18396);
or UO_2416 (O_2416,N_18893,N_16320);
or UO_2417 (O_2417,N_19140,N_18773);
nor UO_2418 (O_2418,N_19763,N_17155);
nand UO_2419 (O_2419,N_19439,N_16011);
xnor UO_2420 (O_2420,N_17497,N_18722);
xnor UO_2421 (O_2421,N_19269,N_16140);
or UO_2422 (O_2422,N_18111,N_17808);
xor UO_2423 (O_2423,N_17947,N_19378);
nand UO_2424 (O_2424,N_17370,N_16214);
or UO_2425 (O_2425,N_18234,N_18010);
nor UO_2426 (O_2426,N_17914,N_16936);
nand UO_2427 (O_2427,N_17736,N_18930);
nand UO_2428 (O_2428,N_19320,N_17466);
nor UO_2429 (O_2429,N_18354,N_16886);
xnor UO_2430 (O_2430,N_16547,N_17432);
or UO_2431 (O_2431,N_18410,N_19308);
nor UO_2432 (O_2432,N_19999,N_16055);
and UO_2433 (O_2433,N_17406,N_19370);
nand UO_2434 (O_2434,N_18305,N_16078);
and UO_2435 (O_2435,N_18661,N_16825);
or UO_2436 (O_2436,N_17844,N_16835);
or UO_2437 (O_2437,N_18755,N_18231);
nor UO_2438 (O_2438,N_17962,N_18696);
nand UO_2439 (O_2439,N_18736,N_17684);
nor UO_2440 (O_2440,N_17889,N_16722);
or UO_2441 (O_2441,N_19268,N_18414);
nor UO_2442 (O_2442,N_17572,N_18979);
and UO_2443 (O_2443,N_19252,N_17837);
or UO_2444 (O_2444,N_16771,N_16130);
or UO_2445 (O_2445,N_16022,N_16001);
or UO_2446 (O_2446,N_19114,N_17041);
and UO_2447 (O_2447,N_18705,N_19299);
nand UO_2448 (O_2448,N_17340,N_18169);
or UO_2449 (O_2449,N_18511,N_16242);
nor UO_2450 (O_2450,N_16306,N_17260);
xnor UO_2451 (O_2451,N_17328,N_18787);
nand UO_2452 (O_2452,N_17327,N_17482);
nand UO_2453 (O_2453,N_19647,N_18203);
and UO_2454 (O_2454,N_19732,N_17795);
and UO_2455 (O_2455,N_19433,N_18807);
and UO_2456 (O_2456,N_17925,N_16955);
nand UO_2457 (O_2457,N_19045,N_17637);
or UO_2458 (O_2458,N_19410,N_19425);
and UO_2459 (O_2459,N_18305,N_16936);
nand UO_2460 (O_2460,N_18747,N_18989);
xnor UO_2461 (O_2461,N_19185,N_19241);
or UO_2462 (O_2462,N_18867,N_17351);
nand UO_2463 (O_2463,N_19067,N_19432);
nand UO_2464 (O_2464,N_17683,N_19406);
or UO_2465 (O_2465,N_16457,N_18292);
nand UO_2466 (O_2466,N_17255,N_19816);
and UO_2467 (O_2467,N_17445,N_16931);
xnor UO_2468 (O_2468,N_16693,N_16976);
xor UO_2469 (O_2469,N_18842,N_18181);
nand UO_2470 (O_2470,N_16498,N_18510);
nand UO_2471 (O_2471,N_19923,N_19067);
xor UO_2472 (O_2472,N_17738,N_16927);
nand UO_2473 (O_2473,N_19418,N_19654);
xnor UO_2474 (O_2474,N_16486,N_18155);
nor UO_2475 (O_2475,N_16363,N_16734);
or UO_2476 (O_2476,N_18768,N_16830);
nor UO_2477 (O_2477,N_18973,N_19663);
and UO_2478 (O_2478,N_19806,N_19059);
or UO_2479 (O_2479,N_19997,N_16731);
nand UO_2480 (O_2480,N_19604,N_19561);
xnor UO_2481 (O_2481,N_19495,N_18975);
and UO_2482 (O_2482,N_18998,N_16995);
and UO_2483 (O_2483,N_16728,N_19681);
nand UO_2484 (O_2484,N_17214,N_18215);
nand UO_2485 (O_2485,N_16204,N_19384);
nand UO_2486 (O_2486,N_17407,N_17160);
nand UO_2487 (O_2487,N_17015,N_18135);
nand UO_2488 (O_2488,N_17954,N_17086);
xor UO_2489 (O_2489,N_19744,N_17094);
and UO_2490 (O_2490,N_16053,N_18941);
and UO_2491 (O_2491,N_18500,N_16554);
and UO_2492 (O_2492,N_19421,N_16566);
nand UO_2493 (O_2493,N_17781,N_18538);
or UO_2494 (O_2494,N_16472,N_16167);
nor UO_2495 (O_2495,N_16470,N_16344);
nand UO_2496 (O_2496,N_19877,N_16741);
nand UO_2497 (O_2497,N_19098,N_19161);
xor UO_2498 (O_2498,N_18488,N_16607);
nand UO_2499 (O_2499,N_19799,N_16858);
endmodule