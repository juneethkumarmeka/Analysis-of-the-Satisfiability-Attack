module basic_500_3000_500_4_levels_2xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_5,In_38);
nor U1 (N_1,In_178,In_44);
xor U2 (N_2,In_268,In_191);
nand U3 (N_3,In_395,In_243);
or U4 (N_4,In_215,In_394);
nand U5 (N_5,In_27,In_55);
or U6 (N_6,In_238,In_190);
nor U7 (N_7,In_35,In_116);
nand U8 (N_8,In_150,In_401);
nand U9 (N_9,In_365,In_0);
nand U10 (N_10,In_407,In_318);
nor U11 (N_11,In_67,In_281);
and U12 (N_12,In_240,In_18);
nor U13 (N_13,In_165,In_46);
and U14 (N_14,In_313,In_154);
nand U15 (N_15,In_287,In_471);
and U16 (N_16,In_284,In_270);
and U17 (N_17,In_175,In_170);
nor U18 (N_18,In_301,In_378);
or U19 (N_19,In_349,In_264);
nor U20 (N_20,In_206,In_379);
and U21 (N_21,In_292,In_193);
or U22 (N_22,In_263,In_4);
and U23 (N_23,In_332,In_380);
or U24 (N_24,In_414,In_455);
nor U25 (N_25,In_48,In_452);
nand U26 (N_26,In_107,In_129);
nor U27 (N_27,In_406,In_295);
or U28 (N_28,In_152,In_119);
nand U29 (N_29,In_135,In_197);
nor U30 (N_30,In_381,In_446);
nor U31 (N_31,In_346,In_312);
or U32 (N_32,In_290,In_438);
or U33 (N_33,In_338,In_239);
nor U34 (N_34,In_54,In_192);
nand U35 (N_35,In_299,In_445);
nor U36 (N_36,In_498,In_147);
or U37 (N_37,In_84,In_242);
nor U38 (N_38,In_371,In_288);
nor U39 (N_39,In_164,In_128);
and U40 (N_40,In_294,In_337);
nor U41 (N_41,In_134,In_50);
or U42 (N_42,In_443,In_375);
nor U43 (N_43,In_405,In_462);
nand U44 (N_44,In_361,In_343);
or U45 (N_45,In_77,In_335);
and U46 (N_46,In_391,In_427);
or U47 (N_47,In_228,In_141);
nand U48 (N_48,In_199,In_248);
nor U49 (N_49,In_465,In_389);
or U50 (N_50,In_61,In_326);
nor U51 (N_51,In_384,In_354);
nor U52 (N_52,In_212,In_103);
xnor U53 (N_53,In_467,In_201);
nand U54 (N_54,In_473,In_475);
and U55 (N_55,In_196,In_433);
or U56 (N_56,In_220,In_278);
and U57 (N_57,In_227,In_366);
nand U58 (N_58,In_101,In_367);
or U59 (N_59,In_83,In_132);
and U60 (N_60,In_202,In_72);
nand U61 (N_61,In_120,In_280);
nand U62 (N_62,In_321,In_320);
nand U63 (N_63,In_183,In_194);
and U64 (N_64,In_355,In_73);
and U65 (N_65,In_151,In_344);
and U66 (N_66,In_252,In_89);
nor U67 (N_67,In_167,In_114);
nor U68 (N_68,In_159,In_26);
nor U69 (N_69,In_370,In_417);
and U70 (N_70,In_289,In_250);
and U71 (N_71,In_231,In_125);
nor U72 (N_72,In_226,In_444);
or U73 (N_73,In_13,In_496);
nor U74 (N_74,In_81,In_387);
nor U75 (N_75,In_492,In_99);
and U76 (N_76,In_442,In_87);
nand U77 (N_77,In_112,In_385);
or U78 (N_78,In_277,In_260);
nand U79 (N_79,In_23,In_434);
and U80 (N_80,In_230,In_65);
and U81 (N_81,In_482,In_136);
nand U82 (N_82,In_138,In_42);
nor U83 (N_83,In_432,In_398);
nand U84 (N_84,In_483,In_341);
or U85 (N_85,In_169,In_168);
or U86 (N_86,In_91,In_106);
nor U87 (N_87,In_499,In_68);
nor U88 (N_88,In_291,In_78);
or U89 (N_89,In_70,In_340);
and U90 (N_90,In_353,In_10);
or U91 (N_91,In_461,In_262);
nand U92 (N_92,In_342,In_241);
or U93 (N_93,In_454,In_331);
nor U94 (N_94,In_397,In_113);
nor U95 (N_95,In_45,In_56);
nand U96 (N_96,In_31,In_362);
nor U97 (N_97,In_53,In_180);
nor U98 (N_98,In_286,In_182);
nor U99 (N_99,In_143,In_396);
and U100 (N_100,In_484,In_328);
nand U101 (N_101,In_276,In_425);
nand U102 (N_102,In_124,In_75);
or U103 (N_103,In_118,In_450);
or U104 (N_104,In_181,In_439);
or U105 (N_105,In_259,In_24);
and U106 (N_106,In_121,In_356);
or U107 (N_107,In_255,In_184);
nor U108 (N_108,In_93,In_3);
or U109 (N_109,In_11,In_464);
nand U110 (N_110,In_373,In_36);
and U111 (N_111,In_218,In_400);
and U112 (N_112,In_51,In_198);
or U113 (N_113,In_495,In_244);
nor U114 (N_114,In_58,In_90);
nor U115 (N_115,In_265,In_123);
or U116 (N_116,In_74,In_98);
nand U117 (N_117,In_383,In_494);
nand U118 (N_118,In_470,In_488);
nor U119 (N_119,In_177,In_40);
or U120 (N_120,In_350,In_279);
or U121 (N_121,In_127,In_79);
nand U122 (N_122,In_322,In_57);
or U123 (N_123,In_217,In_115);
nor U124 (N_124,In_66,In_360);
nand U125 (N_125,In_359,In_108);
or U126 (N_126,In_305,In_310);
and U127 (N_127,In_413,In_109);
and U128 (N_128,In_453,In_148);
and U129 (N_129,In_448,In_261);
nand U130 (N_130,In_298,In_430);
or U131 (N_131,In_176,In_12);
or U132 (N_132,In_21,In_145);
and U133 (N_133,In_80,In_166);
nor U134 (N_134,In_497,In_411);
nand U135 (N_135,In_8,In_86);
nand U136 (N_136,In_348,In_97);
and U137 (N_137,In_418,In_219);
or U138 (N_138,In_468,In_296);
or U139 (N_139,In_306,In_352);
nor U140 (N_140,In_333,In_102);
or U141 (N_141,In_369,In_173);
or U142 (N_142,In_133,In_232);
nor U143 (N_143,In_222,In_372);
or U144 (N_144,In_363,In_161);
nor U145 (N_145,In_476,In_315);
nand U146 (N_146,In_386,In_474);
nor U147 (N_147,In_424,In_308);
nor U148 (N_148,In_142,In_330);
and U149 (N_149,In_449,In_304);
and U150 (N_150,In_25,In_358);
and U151 (N_151,In_325,In_157);
and U152 (N_152,In_428,In_236);
or U153 (N_153,In_435,In_481);
nor U154 (N_154,In_456,In_282);
and U155 (N_155,In_478,In_156);
and U156 (N_156,In_104,In_221);
nor U157 (N_157,In_63,In_186);
xor U158 (N_158,In_303,In_82);
nor U159 (N_159,In_345,In_19);
nand U160 (N_160,In_162,In_160);
nand U161 (N_161,In_216,In_420);
or U162 (N_162,In_28,In_200);
nand U163 (N_163,In_419,In_211);
nand U164 (N_164,In_188,In_149);
or U165 (N_165,In_34,In_253);
nor U166 (N_166,In_88,In_293);
nor U167 (N_167,In_334,In_69);
nand U168 (N_168,In_33,In_213);
xnor U169 (N_169,In_457,In_30);
xnor U170 (N_170,In_22,In_451);
nand U171 (N_171,In_437,In_59);
or U172 (N_172,In_426,In_210);
nor U173 (N_173,In_285,In_440);
nand U174 (N_174,In_17,In_122);
nand U175 (N_175,In_377,In_324);
nand U176 (N_176,In_62,In_158);
and U177 (N_177,In_126,In_466);
and U178 (N_178,In_302,In_195);
nor U179 (N_179,In_96,In_117);
and U180 (N_180,In_267,In_441);
nor U181 (N_181,In_409,In_105);
or U182 (N_182,In_410,In_472);
or U183 (N_183,In_272,In_404);
nor U184 (N_184,In_273,In_469);
nor U185 (N_185,In_347,In_274);
nor U186 (N_186,In_137,In_94);
and U187 (N_187,In_64,In_20);
or U188 (N_188,In_275,In_95);
and U189 (N_189,In_208,In_459);
or U190 (N_190,In_447,In_487);
xnor U191 (N_191,In_237,In_214);
or U192 (N_192,In_390,In_283);
nor U193 (N_193,In_485,In_32);
nand U194 (N_194,In_76,In_323);
nand U195 (N_195,In_39,In_174);
or U196 (N_196,In_131,In_402);
xnor U197 (N_197,In_144,In_209);
nand U198 (N_198,In_60,In_7);
and U199 (N_199,In_223,In_235);
and U200 (N_200,In_140,In_171);
and U201 (N_201,In_431,In_258);
or U202 (N_202,In_153,In_14);
nand U203 (N_203,In_52,In_155);
nand U204 (N_204,In_480,In_43);
and U205 (N_205,In_9,In_463);
and U206 (N_206,In_388,In_203);
xnor U207 (N_207,In_336,In_392);
and U208 (N_208,In_204,In_491);
or U209 (N_209,In_269,In_234);
and U210 (N_210,In_139,In_316);
and U211 (N_211,In_225,In_319);
nor U212 (N_212,In_412,In_300);
and U213 (N_213,In_172,In_16);
xor U214 (N_214,In_339,In_374);
nand U215 (N_215,In_247,In_15);
nand U216 (N_216,In_179,In_364);
and U217 (N_217,In_329,In_256);
nor U218 (N_218,In_49,In_246);
nor U219 (N_219,In_85,In_408);
and U220 (N_220,In_205,In_403);
and U221 (N_221,In_111,In_271);
and U222 (N_222,In_41,In_429);
nor U223 (N_223,In_245,In_146);
nand U224 (N_224,In_399,In_229);
nand U225 (N_225,In_490,In_479);
and U226 (N_226,In_314,In_29);
nor U227 (N_227,In_207,In_233);
nand U228 (N_228,In_393,In_100);
and U229 (N_229,In_460,In_130);
nand U230 (N_230,In_421,In_416);
nand U231 (N_231,In_185,In_309);
nand U232 (N_232,In_317,In_351);
and U233 (N_233,In_307,In_187);
and U234 (N_234,In_254,In_415);
or U235 (N_235,In_6,In_2);
and U236 (N_236,In_311,In_189);
nand U237 (N_237,In_224,In_297);
and U238 (N_238,In_436,In_327);
or U239 (N_239,In_37,In_257);
nand U240 (N_240,In_71,In_251);
nand U241 (N_241,In_163,In_368);
and U242 (N_242,In_493,In_376);
and U243 (N_243,In_1,In_357);
nand U244 (N_244,In_47,In_110);
nand U245 (N_245,In_486,In_458);
nand U246 (N_246,In_422,In_477);
or U247 (N_247,In_489,In_423);
or U248 (N_248,In_249,In_266);
nor U249 (N_249,In_382,In_92);
nand U250 (N_250,In_66,In_72);
or U251 (N_251,In_140,In_238);
and U252 (N_252,In_397,In_414);
or U253 (N_253,In_405,In_458);
and U254 (N_254,In_166,In_266);
or U255 (N_255,In_273,In_282);
nor U256 (N_256,In_376,In_240);
nor U257 (N_257,In_177,In_80);
nor U258 (N_258,In_188,In_343);
and U259 (N_259,In_430,In_445);
or U260 (N_260,In_368,In_52);
or U261 (N_261,In_75,In_421);
and U262 (N_262,In_69,In_317);
nand U263 (N_263,In_490,In_459);
xor U264 (N_264,In_477,In_173);
nand U265 (N_265,In_303,In_231);
and U266 (N_266,In_325,In_71);
and U267 (N_267,In_181,In_447);
xor U268 (N_268,In_317,In_145);
and U269 (N_269,In_463,In_33);
nand U270 (N_270,In_151,In_361);
or U271 (N_271,In_43,In_136);
and U272 (N_272,In_28,In_497);
nand U273 (N_273,In_76,In_66);
nand U274 (N_274,In_420,In_12);
nor U275 (N_275,In_434,In_261);
nor U276 (N_276,In_453,In_420);
nor U277 (N_277,In_439,In_496);
nand U278 (N_278,In_124,In_313);
nor U279 (N_279,In_78,In_223);
and U280 (N_280,In_120,In_104);
nor U281 (N_281,In_80,In_185);
nor U282 (N_282,In_285,In_484);
or U283 (N_283,In_270,In_198);
nor U284 (N_284,In_40,In_468);
nor U285 (N_285,In_149,In_381);
or U286 (N_286,In_115,In_358);
or U287 (N_287,In_436,In_340);
xnor U288 (N_288,In_27,In_76);
or U289 (N_289,In_64,In_306);
and U290 (N_290,In_445,In_340);
nor U291 (N_291,In_439,In_321);
nand U292 (N_292,In_297,In_82);
nor U293 (N_293,In_390,In_107);
nand U294 (N_294,In_352,In_108);
and U295 (N_295,In_45,In_28);
and U296 (N_296,In_364,In_330);
and U297 (N_297,In_130,In_150);
or U298 (N_298,In_114,In_190);
nor U299 (N_299,In_452,In_173);
and U300 (N_300,In_270,In_137);
or U301 (N_301,In_238,In_356);
nor U302 (N_302,In_416,In_401);
or U303 (N_303,In_252,In_296);
or U304 (N_304,In_118,In_287);
nand U305 (N_305,In_442,In_40);
or U306 (N_306,In_140,In_235);
or U307 (N_307,In_257,In_118);
nor U308 (N_308,In_400,In_405);
and U309 (N_309,In_317,In_78);
nor U310 (N_310,In_485,In_270);
or U311 (N_311,In_403,In_412);
nand U312 (N_312,In_145,In_382);
and U313 (N_313,In_267,In_472);
nor U314 (N_314,In_204,In_380);
nor U315 (N_315,In_238,In_33);
and U316 (N_316,In_7,In_385);
and U317 (N_317,In_245,In_53);
nand U318 (N_318,In_240,In_257);
or U319 (N_319,In_319,In_265);
xnor U320 (N_320,In_397,In_48);
or U321 (N_321,In_423,In_201);
nor U322 (N_322,In_182,In_252);
or U323 (N_323,In_239,In_400);
nor U324 (N_324,In_253,In_233);
nor U325 (N_325,In_371,In_67);
nor U326 (N_326,In_0,In_358);
and U327 (N_327,In_202,In_467);
nand U328 (N_328,In_64,In_459);
nor U329 (N_329,In_228,In_109);
nor U330 (N_330,In_359,In_149);
nand U331 (N_331,In_496,In_481);
nor U332 (N_332,In_76,In_361);
nand U333 (N_333,In_454,In_491);
nand U334 (N_334,In_316,In_15);
nand U335 (N_335,In_66,In_114);
nand U336 (N_336,In_328,In_73);
or U337 (N_337,In_331,In_432);
nand U338 (N_338,In_171,In_419);
and U339 (N_339,In_396,In_254);
or U340 (N_340,In_205,In_203);
and U341 (N_341,In_443,In_460);
or U342 (N_342,In_143,In_216);
nand U343 (N_343,In_478,In_225);
nor U344 (N_344,In_384,In_80);
or U345 (N_345,In_415,In_63);
nand U346 (N_346,In_69,In_423);
or U347 (N_347,In_10,In_105);
and U348 (N_348,In_239,In_11);
nand U349 (N_349,In_13,In_25);
nand U350 (N_350,In_28,In_491);
nor U351 (N_351,In_347,In_70);
nor U352 (N_352,In_81,In_243);
nand U353 (N_353,In_474,In_15);
and U354 (N_354,In_353,In_290);
nand U355 (N_355,In_47,In_247);
or U356 (N_356,In_212,In_210);
and U357 (N_357,In_303,In_432);
and U358 (N_358,In_43,In_425);
or U359 (N_359,In_433,In_430);
nand U360 (N_360,In_267,In_430);
or U361 (N_361,In_390,In_387);
nor U362 (N_362,In_216,In_14);
nand U363 (N_363,In_379,In_298);
or U364 (N_364,In_333,In_240);
and U365 (N_365,In_111,In_58);
nand U366 (N_366,In_421,In_257);
or U367 (N_367,In_428,In_385);
and U368 (N_368,In_123,In_460);
nor U369 (N_369,In_110,In_418);
nand U370 (N_370,In_114,In_352);
or U371 (N_371,In_131,In_224);
nor U372 (N_372,In_261,In_58);
and U373 (N_373,In_242,In_440);
nand U374 (N_374,In_280,In_236);
and U375 (N_375,In_277,In_218);
and U376 (N_376,In_126,In_349);
and U377 (N_377,In_375,In_478);
or U378 (N_378,In_330,In_234);
and U379 (N_379,In_419,In_333);
nand U380 (N_380,In_453,In_316);
nor U381 (N_381,In_324,In_29);
and U382 (N_382,In_106,In_231);
and U383 (N_383,In_457,In_105);
or U384 (N_384,In_28,In_213);
and U385 (N_385,In_22,In_273);
and U386 (N_386,In_105,In_406);
and U387 (N_387,In_106,In_311);
nand U388 (N_388,In_478,In_393);
nor U389 (N_389,In_449,In_477);
nand U390 (N_390,In_492,In_335);
nand U391 (N_391,In_89,In_358);
nand U392 (N_392,In_260,In_345);
and U393 (N_393,In_57,In_119);
and U394 (N_394,In_165,In_241);
or U395 (N_395,In_225,In_182);
nand U396 (N_396,In_3,In_438);
nand U397 (N_397,In_126,In_481);
nand U398 (N_398,In_371,In_476);
and U399 (N_399,In_63,In_243);
nor U400 (N_400,In_268,In_95);
and U401 (N_401,In_420,In_304);
nor U402 (N_402,In_95,In_36);
or U403 (N_403,In_131,In_338);
and U404 (N_404,In_195,In_83);
nor U405 (N_405,In_348,In_423);
nand U406 (N_406,In_260,In_58);
and U407 (N_407,In_441,In_161);
nand U408 (N_408,In_302,In_20);
nand U409 (N_409,In_97,In_324);
and U410 (N_410,In_471,In_111);
nand U411 (N_411,In_71,In_272);
and U412 (N_412,In_463,In_295);
nand U413 (N_413,In_483,In_111);
xor U414 (N_414,In_248,In_371);
nor U415 (N_415,In_269,In_370);
and U416 (N_416,In_495,In_18);
and U417 (N_417,In_59,In_65);
or U418 (N_418,In_224,In_218);
or U419 (N_419,In_244,In_499);
or U420 (N_420,In_306,In_343);
nor U421 (N_421,In_387,In_360);
or U422 (N_422,In_69,In_389);
nor U423 (N_423,In_375,In_228);
xnor U424 (N_424,In_226,In_425);
and U425 (N_425,In_296,In_22);
and U426 (N_426,In_166,In_475);
or U427 (N_427,In_156,In_268);
and U428 (N_428,In_101,In_163);
or U429 (N_429,In_194,In_122);
or U430 (N_430,In_208,In_374);
nor U431 (N_431,In_162,In_154);
or U432 (N_432,In_216,In_329);
nand U433 (N_433,In_413,In_122);
and U434 (N_434,In_59,In_388);
nor U435 (N_435,In_489,In_156);
and U436 (N_436,In_417,In_439);
nor U437 (N_437,In_320,In_295);
nor U438 (N_438,In_139,In_244);
and U439 (N_439,In_379,In_122);
and U440 (N_440,In_163,In_470);
nand U441 (N_441,In_103,In_316);
nor U442 (N_442,In_34,In_333);
nor U443 (N_443,In_245,In_33);
nor U444 (N_444,In_65,In_274);
or U445 (N_445,In_138,In_284);
nand U446 (N_446,In_127,In_392);
nor U447 (N_447,In_145,In_207);
and U448 (N_448,In_108,In_294);
or U449 (N_449,In_382,In_77);
nor U450 (N_450,In_52,In_390);
and U451 (N_451,In_340,In_342);
nand U452 (N_452,In_297,In_295);
or U453 (N_453,In_116,In_295);
or U454 (N_454,In_340,In_229);
and U455 (N_455,In_265,In_466);
nor U456 (N_456,In_247,In_377);
and U457 (N_457,In_216,In_125);
or U458 (N_458,In_312,In_406);
nand U459 (N_459,In_67,In_43);
and U460 (N_460,In_338,In_130);
nand U461 (N_461,In_362,In_369);
nand U462 (N_462,In_155,In_341);
nor U463 (N_463,In_37,In_61);
or U464 (N_464,In_406,In_493);
nand U465 (N_465,In_328,In_72);
nor U466 (N_466,In_362,In_2);
or U467 (N_467,In_424,In_261);
nand U468 (N_468,In_153,In_384);
and U469 (N_469,In_393,In_48);
and U470 (N_470,In_416,In_154);
or U471 (N_471,In_482,In_45);
or U472 (N_472,In_98,In_342);
and U473 (N_473,In_75,In_16);
nor U474 (N_474,In_231,In_315);
nor U475 (N_475,In_31,In_365);
or U476 (N_476,In_179,In_422);
nor U477 (N_477,In_120,In_85);
nor U478 (N_478,In_479,In_377);
nor U479 (N_479,In_70,In_127);
nand U480 (N_480,In_94,In_26);
nand U481 (N_481,In_155,In_157);
nor U482 (N_482,In_93,In_0);
and U483 (N_483,In_41,In_452);
nor U484 (N_484,In_145,In_98);
nand U485 (N_485,In_244,In_175);
or U486 (N_486,In_28,In_131);
and U487 (N_487,In_234,In_298);
or U488 (N_488,In_449,In_51);
nor U489 (N_489,In_282,In_422);
and U490 (N_490,In_168,In_126);
nand U491 (N_491,In_384,In_206);
or U492 (N_492,In_375,In_12);
nor U493 (N_493,In_78,In_172);
xor U494 (N_494,In_103,In_344);
or U495 (N_495,In_351,In_391);
nor U496 (N_496,In_300,In_458);
nor U497 (N_497,In_469,In_125);
nand U498 (N_498,In_236,In_184);
and U499 (N_499,In_261,In_404);
or U500 (N_500,In_135,In_183);
nor U501 (N_501,In_384,In_295);
or U502 (N_502,In_401,In_371);
nand U503 (N_503,In_32,In_369);
or U504 (N_504,In_241,In_264);
and U505 (N_505,In_494,In_15);
or U506 (N_506,In_107,In_378);
nand U507 (N_507,In_177,In_342);
and U508 (N_508,In_449,In_239);
nand U509 (N_509,In_232,In_187);
or U510 (N_510,In_285,In_130);
and U511 (N_511,In_302,In_154);
nand U512 (N_512,In_405,In_224);
nor U513 (N_513,In_47,In_425);
nand U514 (N_514,In_148,In_101);
nand U515 (N_515,In_181,In_343);
nand U516 (N_516,In_191,In_238);
or U517 (N_517,In_15,In_289);
nand U518 (N_518,In_38,In_442);
nor U519 (N_519,In_348,In_133);
or U520 (N_520,In_447,In_439);
nor U521 (N_521,In_397,In_168);
and U522 (N_522,In_154,In_454);
and U523 (N_523,In_195,In_13);
nor U524 (N_524,In_103,In_296);
nor U525 (N_525,In_464,In_121);
or U526 (N_526,In_387,In_398);
and U527 (N_527,In_174,In_126);
and U528 (N_528,In_461,In_445);
and U529 (N_529,In_259,In_464);
and U530 (N_530,In_380,In_41);
nand U531 (N_531,In_383,In_142);
and U532 (N_532,In_358,In_62);
nor U533 (N_533,In_472,In_448);
nor U534 (N_534,In_44,In_43);
nor U535 (N_535,In_283,In_448);
or U536 (N_536,In_299,In_110);
nor U537 (N_537,In_390,In_340);
or U538 (N_538,In_472,In_414);
and U539 (N_539,In_238,In_125);
nor U540 (N_540,In_399,In_134);
nand U541 (N_541,In_0,In_408);
and U542 (N_542,In_55,In_22);
nand U543 (N_543,In_19,In_494);
nand U544 (N_544,In_261,In_117);
nor U545 (N_545,In_61,In_266);
nor U546 (N_546,In_276,In_135);
nor U547 (N_547,In_193,In_463);
nand U548 (N_548,In_428,In_52);
nor U549 (N_549,In_228,In_66);
nor U550 (N_550,In_443,In_368);
or U551 (N_551,In_305,In_142);
nand U552 (N_552,In_119,In_106);
nor U553 (N_553,In_121,In_6);
nor U554 (N_554,In_424,In_450);
nand U555 (N_555,In_418,In_28);
or U556 (N_556,In_3,In_313);
nor U557 (N_557,In_151,In_258);
or U558 (N_558,In_227,In_76);
nor U559 (N_559,In_332,In_411);
or U560 (N_560,In_102,In_134);
and U561 (N_561,In_295,In_379);
or U562 (N_562,In_94,In_404);
or U563 (N_563,In_56,In_147);
nor U564 (N_564,In_285,In_302);
and U565 (N_565,In_493,In_47);
nand U566 (N_566,In_266,In_244);
xnor U567 (N_567,In_375,In_252);
nand U568 (N_568,In_249,In_287);
nor U569 (N_569,In_24,In_3);
nor U570 (N_570,In_342,In_322);
or U571 (N_571,In_286,In_451);
xor U572 (N_572,In_373,In_239);
nor U573 (N_573,In_181,In_14);
nand U574 (N_574,In_376,In_424);
nand U575 (N_575,In_126,In_152);
nor U576 (N_576,In_414,In_423);
nor U577 (N_577,In_180,In_186);
or U578 (N_578,In_316,In_69);
or U579 (N_579,In_385,In_41);
nor U580 (N_580,In_96,In_493);
nand U581 (N_581,In_94,In_355);
nor U582 (N_582,In_489,In_150);
and U583 (N_583,In_344,In_474);
nor U584 (N_584,In_147,In_51);
or U585 (N_585,In_335,In_419);
nor U586 (N_586,In_481,In_134);
and U587 (N_587,In_451,In_267);
nor U588 (N_588,In_491,In_174);
xnor U589 (N_589,In_309,In_56);
nand U590 (N_590,In_228,In_7);
nor U591 (N_591,In_24,In_93);
or U592 (N_592,In_415,In_88);
nand U593 (N_593,In_202,In_452);
nand U594 (N_594,In_295,In_402);
nand U595 (N_595,In_200,In_290);
and U596 (N_596,In_130,In_18);
nor U597 (N_597,In_216,In_240);
or U598 (N_598,In_374,In_286);
nand U599 (N_599,In_85,In_111);
and U600 (N_600,In_161,In_179);
nor U601 (N_601,In_199,In_441);
or U602 (N_602,In_162,In_487);
nand U603 (N_603,In_402,In_359);
and U604 (N_604,In_448,In_63);
nand U605 (N_605,In_320,In_104);
nand U606 (N_606,In_109,In_89);
nand U607 (N_607,In_250,In_141);
and U608 (N_608,In_280,In_468);
and U609 (N_609,In_310,In_410);
or U610 (N_610,In_293,In_64);
and U611 (N_611,In_412,In_356);
nand U612 (N_612,In_417,In_466);
nand U613 (N_613,In_458,In_263);
and U614 (N_614,In_78,In_128);
and U615 (N_615,In_14,In_402);
nand U616 (N_616,In_145,In_331);
nand U617 (N_617,In_332,In_410);
nand U618 (N_618,In_92,In_13);
or U619 (N_619,In_118,In_71);
and U620 (N_620,In_306,In_245);
nand U621 (N_621,In_461,In_475);
and U622 (N_622,In_482,In_389);
and U623 (N_623,In_155,In_443);
nand U624 (N_624,In_303,In_221);
nor U625 (N_625,In_369,In_65);
nor U626 (N_626,In_428,In_137);
xor U627 (N_627,In_119,In_18);
nor U628 (N_628,In_78,In_67);
nand U629 (N_629,In_36,In_303);
or U630 (N_630,In_369,In_129);
or U631 (N_631,In_363,In_374);
or U632 (N_632,In_379,In_372);
nand U633 (N_633,In_183,In_472);
or U634 (N_634,In_354,In_345);
nand U635 (N_635,In_199,In_477);
nor U636 (N_636,In_334,In_275);
nand U637 (N_637,In_357,In_113);
and U638 (N_638,In_419,In_125);
and U639 (N_639,In_162,In_64);
nand U640 (N_640,In_355,In_317);
nand U641 (N_641,In_458,In_138);
or U642 (N_642,In_287,In_448);
nor U643 (N_643,In_161,In_17);
and U644 (N_644,In_397,In_428);
nor U645 (N_645,In_272,In_330);
or U646 (N_646,In_380,In_212);
and U647 (N_647,In_286,In_168);
nand U648 (N_648,In_126,In_452);
nor U649 (N_649,In_117,In_204);
and U650 (N_650,In_134,In_105);
or U651 (N_651,In_402,In_37);
and U652 (N_652,In_441,In_45);
nand U653 (N_653,In_29,In_148);
nor U654 (N_654,In_476,In_273);
nand U655 (N_655,In_5,In_429);
or U656 (N_656,In_404,In_378);
nand U657 (N_657,In_77,In_310);
nand U658 (N_658,In_468,In_264);
nor U659 (N_659,In_200,In_7);
and U660 (N_660,In_440,In_27);
or U661 (N_661,In_430,In_135);
nor U662 (N_662,In_356,In_267);
or U663 (N_663,In_280,In_432);
nand U664 (N_664,In_255,In_391);
nor U665 (N_665,In_133,In_245);
nand U666 (N_666,In_412,In_256);
or U667 (N_667,In_179,In_240);
or U668 (N_668,In_332,In_221);
or U669 (N_669,In_204,In_266);
and U670 (N_670,In_74,In_183);
or U671 (N_671,In_100,In_346);
and U672 (N_672,In_169,In_13);
or U673 (N_673,In_331,In_173);
nand U674 (N_674,In_210,In_435);
and U675 (N_675,In_212,In_23);
nand U676 (N_676,In_312,In_439);
or U677 (N_677,In_4,In_359);
nor U678 (N_678,In_40,In_250);
nand U679 (N_679,In_168,In_406);
and U680 (N_680,In_148,In_414);
nand U681 (N_681,In_328,In_18);
nor U682 (N_682,In_351,In_300);
nand U683 (N_683,In_93,In_284);
nor U684 (N_684,In_207,In_206);
and U685 (N_685,In_148,In_323);
or U686 (N_686,In_447,In_79);
xor U687 (N_687,In_6,In_295);
nand U688 (N_688,In_151,In_306);
or U689 (N_689,In_57,In_425);
or U690 (N_690,In_47,In_133);
nand U691 (N_691,In_486,In_330);
nand U692 (N_692,In_220,In_374);
or U693 (N_693,In_433,In_203);
and U694 (N_694,In_414,In_21);
or U695 (N_695,In_296,In_42);
nand U696 (N_696,In_137,In_287);
or U697 (N_697,In_497,In_118);
nor U698 (N_698,In_1,In_282);
nor U699 (N_699,In_409,In_209);
nor U700 (N_700,In_347,In_480);
nor U701 (N_701,In_118,In_135);
nand U702 (N_702,In_464,In_169);
and U703 (N_703,In_192,In_158);
and U704 (N_704,In_9,In_213);
and U705 (N_705,In_448,In_393);
or U706 (N_706,In_238,In_44);
nand U707 (N_707,In_13,In_93);
nor U708 (N_708,In_27,In_60);
nand U709 (N_709,In_67,In_56);
and U710 (N_710,In_79,In_133);
nor U711 (N_711,In_256,In_157);
or U712 (N_712,In_83,In_158);
nand U713 (N_713,In_130,In_69);
nor U714 (N_714,In_225,In_308);
and U715 (N_715,In_435,In_226);
nand U716 (N_716,In_66,In_128);
nor U717 (N_717,In_311,In_308);
and U718 (N_718,In_283,In_395);
nand U719 (N_719,In_201,In_253);
and U720 (N_720,In_120,In_92);
or U721 (N_721,In_399,In_223);
nor U722 (N_722,In_162,In_422);
nor U723 (N_723,In_318,In_295);
nand U724 (N_724,In_240,In_24);
and U725 (N_725,In_353,In_21);
nor U726 (N_726,In_0,In_498);
nor U727 (N_727,In_200,In_425);
or U728 (N_728,In_10,In_152);
and U729 (N_729,In_150,In_432);
and U730 (N_730,In_143,In_259);
nand U731 (N_731,In_338,In_105);
nor U732 (N_732,In_164,In_271);
and U733 (N_733,In_79,In_333);
nor U734 (N_734,In_34,In_184);
or U735 (N_735,In_280,In_374);
nor U736 (N_736,In_311,In_154);
nor U737 (N_737,In_394,In_429);
nand U738 (N_738,In_141,In_394);
or U739 (N_739,In_294,In_380);
or U740 (N_740,In_354,In_298);
and U741 (N_741,In_167,In_123);
or U742 (N_742,In_206,In_132);
and U743 (N_743,In_463,In_180);
nand U744 (N_744,In_409,In_234);
nor U745 (N_745,In_87,In_204);
and U746 (N_746,In_314,In_130);
nand U747 (N_747,In_475,In_484);
and U748 (N_748,In_235,In_263);
nand U749 (N_749,In_184,In_168);
nand U750 (N_750,N_346,N_131);
xnor U751 (N_751,N_392,N_628);
nand U752 (N_752,N_583,N_66);
or U753 (N_753,N_182,N_744);
and U754 (N_754,N_63,N_247);
nor U755 (N_755,N_322,N_132);
or U756 (N_756,N_613,N_353);
nor U757 (N_757,N_422,N_690);
nor U758 (N_758,N_205,N_499);
nor U759 (N_759,N_437,N_229);
or U760 (N_760,N_442,N_526);
or U761 (N_761,N_407,N_98);
or U762 (N_762,N_308,N_696);
and U763 (N_763,N_553,N_279);
nand U764 (N_764,N_725,N_710);
nand U765 (N_765,N_298,N_697);
or U766 (N_766,N_103,N_577);
nand U767 (N_767,N_562,N_644);
nand U768 (N_768,N_221,N_27);
and U769 (N_769,N_579,N_109);
or U770 (N_770,N_162,N_77);
or U771 (N_771,N_248,N_505);
nand U772 (N_772,N_328,N_657);
nand U773 (N_773,N_151,N_508);
nor U774 (N_774,N_715,N_303);
or U775 (N_775,N_480,N_128);
and U776 (N_776,N_184,N_159);
or U777 (N_777,N_438,N_133);
and U778 (N_778,N_101,N_211);
or U779 (N_779,N_317,N_224);
and U780 (N_780,N_114,N_246);
nand U781 (N_781,N_209,N_739);
and U782 (N_782,N_724,N_196);
or U783 (N_783,N_73,N_576);
nand U784 (N_784,N_30,N_389);
nor U785 (N_785,N_462,N_412);
nor U786 (N_786,N_471,N_306);
or U787 (N_787,N_15,N_496);
xnor U788 (N_788,N_378,N_520);
nor U789 (N_789,N_222,N_423);
nand U790 (N_790,N_380,N_141);
nor U791 (N_791,N_347,N_646);
nor U792 (N_792,N_268,N_108);
nor U793 (N_793,N_460,N_507);
and U794 (N_794,N_403,N_519);
or U795 (N_795,N_321,N_71);
or U796 (N_796,N_603,N_421);
nand U797 (N_797,N_194,N_21);
nand U798 (N_798,N_326,N_714);
or U799 (N_799,N_623,N_273);
and U800 (N_800,N_381,N_700);
and U801 (N_801,N_351,N_129);
nor U802 (N_802,N_521,N_658);
nand U803 (N_803,N_656,N_459);
nand U804 (N_804,N_388,N_664);
nor U805 (N_805,N_626,N_284);
and U806 (N_806,N_722,N_427);
and U807 (N_807,N_467,N_271);
nand U808 (N_808,N_568,N_594);
nand U809 (N_809,N_359,N_22);
nand U810 (N_810,N_622,N_58);
nor U811 (N_811,N_361,N_534);
nand U812 (N_812,N_340,N_174);
or U813 (N_813,N_34,N_226);
and U814 (N_814,N_208,N_160);
nor U815 (N_815,N_400,N_153);
nor U816 (N_816,N_681,N_466);
nand U817 (N_817,N_698,N_627);
and U818 (N_818,N_572,N_530);
nor U819 (N_819,N_201,N_425);
or U820 (N_820,N_147,N_483);
nand U821 (N_821,N_26,N_563);
and U822 (N_822,N_629,N_90);
and U823 (N_823,N_197,N_587);
or U824 (N_824,N_500,N_255);
xor U825 (N_825,N_189,N_416);
nor U826 (N_826,N_327,N_625);
nand U827 (N_827,N_558,N_431);
xor U828 (N_828,N_81,N_447);
nor U829 (N_829,N_83,N_238);
and U830 (N_830,N_741,N_14);
nor U831 (N_831,N_379,N_213);
and U832 (N_832,N_580,N_72);
nor U833 (N_833,N_158,N_297);
nand U834 (N_834,N_310,N_239);
nor U835 (N_835,N_4,N_355);
nor U836 (N_836,N_60,N_706);
and U837 (N_837,N_64,N_228);
or U838 (N_838,N_316,N_143);
or U839 (N_839,N_343,N_193);
or U840 (N_840,N_53,N_104);
and U841 (N_841,N_111,N_481);
nand U842 (N_842,N_608,N_149);
or U843 (N_843,N_0,N_542);
and U844 (N_844,N_288,N_296);
nand U845 (N_845,N_533,N_417);
or U846 (N_846,N_641,N_91);
or U847 (N_847,N_446,N_348);
or U848 (N_848,N_44,N_142);
or U849 (N_849,N_490,N_282);
nor U850 (N_850,N_396,N_509);
or U851 (N_851,N_589,N_736);
and U852 (N_852,N_430,N_274);
or U853 (N_853,N_721,N_391);
nand U854 (N_854,N_694,N_666);
and U855 (N_855,N_107,N_212);
or U856 (N_856,N_119,N_102);
or U857 (N_857,N_541,N_59);
nand U858 (N_858,N_537,N_514);
and U859 (N_859,N_311,N_262);
nor U860 (N_860,N_707,N_640);
or U861 (N_861,N_332,N_597);
xnor U862 (N_862,N_299,N_426);
nor U863 (N_863,N_614,N_390);
or U864 (N_864,N_555,N_305);
nand U865 (N_865,N_254,N_415);
xor U866 (N_866,N_80,N_188);
or U867 (N_867,N_538,N_32);
and U868 (N_868,N_344,N_635);
nor U869 (N_869,N_257,N_264);
nor U870 (N_870,N_662,N_146);
and U871 (N_871,N_670,N_200);
and U872 (N_872,N_410,N_419);
and U873 (N_873,N_424,N_740);
or U874 (N_874,N_470,N_660);
or U875 (N_875,N_55,N_548);
nand U876 (N_876,N_74,N_746);
or U877 (N_877,N_561,N_515);
or U878 (N_878,N_632,N_293);
and U879 (N_879,N_588,N_38);
or U880 (N_880,N_445,N_675);
nand U881 (N_881,N_144,N_56);
and U882 (N_882,N_99,N_653);
and U883 (N_883,N_186,N_337);
or U884 (N_884,N_281,N_312);
or U885 (N_885,N_270,N_105);
or U886 (N_886,N_525,N_749);
nor U887 (N_887,N_37,N_365);
nand U888 (N_888,N_287,N_461);
or U889 (N_889,N_550,N_349);
nand U890 (N_890,N_643,N_573);
and U891 (N_891,N_180,N_605);
and U892 (N_892,N_259,N_527);
nor U893 (N_893,N_713,N_16);
and U894 (N_894,N_733,N_176);
nor U895 (N_895,N_23,N_214);
nor U896 (N_896,N_649,N_127);
and U897 (N_897,N_371,N_253);
and U898 (N_898,N_155,N_2);
or U899 (N_899,N_290,N_518);
or U900 (N_900,N_258,N_479);
nand U901 (N_901,N_5,N_168);
nand U902 (N_902,N_263,N_225);
and U903 (N_903,N_528,N_374);
or U904 (N_904,N_171,N_592);
nand U905 (N_905,N_708,N_249);
and U906 (N_906,N_36,N_596);
nor U907 (N_907,N_604,N_448);
nor U908 (N_908,N_130,N_731);
and U909 (N_909,N_712,N_165);
and U910 (N_910,N_41,N_336);
nor U911 (N_911,N_89,N_190);
or U912 (N_912,N_630,N_484);
nor U913 (N_913,N_590,N_680);
and U914 (N_914,N_511,N_54);
nor U915 (N_915,N_338,N_601);
nand U916 (N_916,N_362,N_70);
nand U917 (N_917,N_325,N_642);
xor U918 (N_918,N_11,N_637);
or U919 (N_919,N_172,N_323);
nand U920 (N_920,N_384,N_702);
and U921 (N_921,N_12,N_455);
and U922 (N_922,N_345,N_547);
and U923 (N_923,N_18,N_354);
nor U924 (N_924,N_185,N_1);
or U925 (N_925,N_84,N_156);
and U926 (N_926,N_535,N_230);
nand U927 (N_927,N_616,N_251);
xnor U928 (N_928,N_95,N_450);
nand U929 (N_929,N_19,N_112);
nand U930 (N_930,N_350,N_401);
nor U931 (N_931,N_676,N_621);
or U932 (N_932,N_652,N_494);
nor U933 (N_933,N_339,N_543);
nand U934 (N_934,N_598,N_244);
nor U935 (N_935,N_639,N_20);
nand U936 (N_936,N_567,N_24);
or U937 (N_937,N_96,N_217);
and U938 (N_938,N_469,N_210);
nand U939 (N_939,N_352,N_25);
or U940 (N_940,N_309,N_117);
nor U941 (N_941,N_385,N_517);
and U942 (N_942,N_689,N_647);
and U943 (N_943,N_748,N_687);
and U944 (N_944,N_62,N_408);
nor U945 (N_945,N_223,N_28);
or U946 (N_946,N_357,N_31);
nor U947 (N_947,N_115,N_522);
nand U948 (N_948,N_650,N_192);
nand U949 (N_949,N_586,N_655);
nand U950 (N_950,N_68,N_49);
or U951 (N_951,N_178,N_314);
or U952 (N_952,N_584,N_397);
or U953 (N_953,N_283,N_50);
nand U954 (N_954,N_559,N_585);
and U955 (N_955,N_612,N_599);
nand U956 (N_956,N_454,N_506);
nand U957 (N_957,N_595,N_57);
nand U958 (N_958,N_728,N_665);
nand U959 (N_959,N_154,N_368);
nor U960 (N_960,N_175,N_79);
nor U961 (N_961,N_705,N_669);
nand U962 (N_962,N_219,N_651);
nor U963 (N_963,N_566,N_560);
nand U964 (N_964,N_711,N_33);
xnor U965 (N_965,N_110,N_181);
or U966 (N_966,N_512,N_449);
nand U967 (N_967,N_377,N_668);
nor U968 (N_968,N_418,N_444);
nand U969 (N_969,N_206,N_315);
nand U970 (N_970,N_491,N_93);
and U971 (N_971,N_234,N_545);
or U972 (N_972,N_198,N_574);
nor U973 (N_973,N_717,N_285);
nor U974 (N_974,N_157,N_456);
nand U975 (N_975,N_593,N_659);
nand U976 (N_976,N_497,N_243);
nand U977 (N_977,N_709,N_732);
nand U978 (N_978,N_126,N_406);
nor U979 (N_979,N_360,N_363);
and U980 (N_980,N_477,N_75);
nand U981 (N_981,N_683,N_204);
and U982 (N_982,N_672,N_493);
or U983 (N_983,N_654,N_578);
nor U984 (N_984,N_17,N_123);
nand U985 (N_985,N_602,N_276);
xor U986 (N_986,N_420,N_743);
and U987 (N_987,N_39,N_367);
nand U988 (N_988,N_536,N_277);
nand U989 (N_989,N_47,N_723);
nand U990 (N_990,N_398,N_638);
nor U991 (N_991,N_125,N_730);
nand U992 (N_992,N_386,N_393);
nor U993 (N_993,N_402,N_51);
or U994 (N_994,N_726,N_674);
nor U995 (N_995,N_358,N_240);
nor U996 (N_996,N_693,N_742);
nand U997 (N_997,N_729,N_435);
nor U998 (N_998,N_13,N_439);
and U999 (N_999,N_195,N_611);
nor U1000 (N_1000,N_301,N_502);
or U1001 (N_1001,N_256,N_472);
nand U1002 (N_1002,N_624,N_161);
nor U1003 (N_1003,N_556,N_453);
or U1004 (N_1004,N_241,N_679);
nor U1005 (N_1005,N_387,N_292);
nor U1006 (N_1006,N_82,N_250);
nor U1007 (N_1007,N_510,N_600);
nand U1008 (N_1008,N_554,N_695);
nor U1009 (N_1009,N_463,N_571);
and U1010 (N_1010,N_342,N_320);
and U1011 (N_1011,N_570,N_546);
or U1012 (N_1012,N_235,N_451);
and U1013 (N_1013,N_474,N_458);
or U1014 (N_1014,N_313,N_747);
and U1015 (N_1015,N_513,N_489);
nor U1016 (N_1016,N_9,N_475);
nor U1017 (N_1017,N_35,N_3);
nor U1018 (N_1018,N_183,N_607);
nand U1019 (N_1019,N_356,N_61);
and U1020 (N_1020,N_395,N_699);
and U1021 (N_1021,N_164,N_330);
nand U1022 (N_1022,N_366,N_242);
nand U1023 (N_1023,N_267,N_120);
and U1024 (N_1024,N_544,N_187);
nand U1025 (N_1025,N_122,N_615);
nor U1026 (N_1026,N_436,N_409);
nor U1027 (N_1027,N_7,N_482);
nor U1028 (N_1028,N_324,N_488);
and U1029 (N_1029,N_487,N_734);
nand U1030 (N_1030,N_43,N_701);
nand U1031 (N_1031,N_45,N_452);
nand U1032 (N_1032,N_434,N_684);
nand U1033 (N_1033,N_331,N_231);
and U1034 (N_1034,N_485,N_202);
and U1035 (N_1035,N_100,N_719);
and U1036 (N_1036,N_617,N_302);
or U1037 (N_1037,N_745,N_688);
nand U1038 (N_1038,N_272,N_220);
nand U1039 (N_1039,N_404,N_682);
nor U1040 (N_1040,N_40,N_76);
and U1041 (N_1041,N_245,N_432);
or U1042 (N_1042,N_118,N_227);
nor U1043 (N_1043,N_163,N_85);
nor U1044 (N_1044,N_692,N_501);
nor U1045 (N_1045,N_166,N_370);
nand U1046 (N_1046,N_703,N_464);
and U1047 (N_1047,N_620,N_121);
nor U1048 (N_1048,N_631,N_531);
or U1049 (N_1049,N_179,N_138);
nor U1050 (N_1050,N_411,N_405);
or U1051 (N_1051,N_372,N_106);
and U1052 (N_1052,N_465,N_215);
nor U1053 (N_1053,N_291,N_275);
and U1054 (N_1054,N_232,N_648);
nand U1055 (N_1055,N_116,N_591);
or U1056 (N_1056,N_318,N_335);
nor U1057 (N_1057,N_294,N_504);
nand U1058 (N_1058,N_428,N_307);
nor U1059 (N_1059,N_609,N_457);
or U1060 (N_1060,N_295,N_286);
or U1061 (N_1061,N_261,N_619);
nand U1062 (N_1062,N_492,N_382);
or U1063 (N_1063,N_29,N_685);
and U1064 (N_1064,N_8,N_678);
or U1065 (N_1065,N_486,N_532);
and U1066 (N_1066,N_341,N_565);
or U1067 (N_1067,N_236,N_581);
nor U1068 (N_1068,N_167,N_667);
nor U1069 (N_1069,N_124,N_375);
or U1070 (N_1070,N_139,N_280);
or U1071 (N_1071,N_704,N_414);
nor U1072 (N_1072,N_52,N_495);
nand U1073 (N_1073,N_237,N_191);
nor U1074 (N_1074,N_720,N_319);
nor U1075 (N_1075,N_671,N_373);
nand U1076 (N_1076,N_476,N_333);
or U1077 (N_1077,N_473,N_92);
and U1078 (N_1078,N_46,N_300);
and U1079 (N_1079,N_718,N_42);
or U1080 (N_1080,N_218,N_569);
nor U1081 (N_1081,N_441,N_216);
and U1082 (N_1082,N_478,N_65);
or U1083 (N_1083,N_140,N_737);
nand U1084 (N_1084,N_364,N_413);
or U1085 (N_1085,N_252,N_67);
or U1086 (N_1086,N_97,N_94);
nor U1087 (N_1087,N_661,N_429);
or U1088 (N_1088,N_78,N_334);
and U1089 (N_1089,N_6,N_673);
or U1090 (N_1090,N_524,N_289);
nor U1091 (N_1091,N_686,N_260);
and U1092 (N_1092,N_134,N_443);
nor U1093 (N_1093,N_691,N_735);
and U1094 (N_1094,N_369,N_169);
nor U1095 (N_1095,N_113,N_634);
nand U1096 (N_1096,N_173,N_177);
nand U1097 (N_1097,N_87,N_633);
xor U1098 (N_1098,N_266,N_48);
nand U1099 (N_1099,N_440,N_606);
nor U1100 (N_1100,N_636,N_552);
and U1101 (N_1101,N_551,N_663);
nand U1102 (N_1102,N_137,N_738);
and U1103 (N_1103,N_540,N_265);
nor U1104 (N_1104,N_549,N_557);
or U1105 (N_1105,N_399,N_278);
nor U1106 (N_1106,N_575,N_618);
nor U1107 (N_1107,N_207,N_145);
and U1108 (N_1108,N_170,N_468);
nor U1109 (N_1109,N_329,N_383);
nor U1110 (N_1110,N_529,N_10);
nor U1111 (N_1111,N_610,N_376);
and U1112 (N_1112,N_516,N_150);
nand U1113 (N_1113,N_539,N_152);
and U1114 (N_1114,N_304,N_269);
and U1115 (N_1115,N_199,N_564);
nand U1116 (N_1116,N_233,N_677);
and U1117 (N_1117,N_394,N_86);
nand U1118 (N_1118,N_523,N_645);
nand U1119 (N_1119,N_69,N_727);
and U1120 (N_1120,N_203,N_433);
or U1121 (N_1121,N_135,N_498);
nor U1122 (N_1122,N_136,N_148);
nand U1123 (N_1123,N_88,N_582);
nor U1124 (N_1124,N_503,N_716);
or U1125 (N_1125,N_319,N_178);
nand U1126 (N_1126,N_513,N_534);
and U1127 (N_1127,N_18,N_669);
nor U1128 (N_1128,N_555,N_641);
nand U1129 (N_1129,N_636,N_363);
or U1130 (N_1130,N_592,N_152);
or U1131 (N_1131,N_487,N_52);
nor U1132 (N_1132,N_327,N_420);
nor U1133 (N_1133,N_609,N_474);
nand U1134 (N_1134,N_680,N_50);
nand U1135 (N_1135,N_330,N_38);
and U1136 (N_1136,N_305,N_494);
and U1137 (N_1137,N_594,N_142);
nor U1138 (N_1138,N_131,N_50);
or U1139 (N_1139,N_669,N_63);
nand U1140 (N_1140,N_424,N_674);
and U1141 (N_1141,N_557,N_9);
and U1142 (N_1142,N_18,N_204);
nand U1143 (N_1143,N_685,N_674);
or U1144 (N_1144,N_76,N_470);
nand U1145 (N_1145,N_665,N_690);
or U1146 (N_1146,N_256,N_345);
nor U1147 (N_1147,N_748,N_279);
xnor U1148 (N_1148,N_739,N_384);
and U1149 (N_1149,N_663,N_76);
or U1150 (N_1150,N_708,N_729);
and U1151 (N_1151,N_168,N_271);
or U1152 (N_1152,N_115,N_298);
nand U1153 (N_1153,N_680,N_424);
and U1154 (N_1154,N_135,N_446);
nand U1155 (N_1155,N_510,N_341);
xor U1156 (N_1156,N_486,N_624);
or U1157 (N_1157,N_686,N_180);
or U1158 (N_1158,N_118,N_3);
and U1159 (N_1159,N_557,N_384);
nor U1160 (N_1160,N_278,N_725);
nor U1161 (N_1161,N_505,N_250);
nor U1162 (N_1162,N_639,N_421);
nor U1163 (N_1163,N_420,N_511);
and U1164 (N_1164,N_585,N_451);
or U1165 (N_1165,N_69,N_463);
and U1166 (N_1166,N_150,N_305);
nor U1167 (N_1167,N_523,N_349);
nand U1168 (N_1168,N_20,N_40);
and U1169 (N_1169,N_277,N_34);
and U1170 (N_1170,N_663,N_521);
or U1171 (N_1171,N_91,N_437);
or U1172 (N_1172,N_105,N_641);
nor U1173 (N_1173,N_338,N_340);
nand U1174 (N_1174,N_308,N_152);
nand U1175 (N_1175,N_242,N_727);
or U1176 (N_1176,N_391,N_701);
and U1177 (N_1177,N_593,N_112);
nor U1178 (N_1178,N_352,N_416);
nor U1179 (N_1179,N_486,N_185);
and U1180 (N_1180,N_619,N_383);
or U1181 (N_1181,N_215,N_574);
and U1182 (N_1182,N_162,N_628);
nand U1183 (N_1183,N_331,N_77);
nor U1184 (N_1184,N_502,N_241);
and U1185 (N_1185,N_10,N_206);
or U1186 (N_1186,N_164,N_45);
or U1187 (N_1187,N_483,N_650);
nand U1188 (N_1188,N_440,N_531);
nand U1189 (N_1189,N_87,N_21);
nor U1190 (N_1190,N_90,N_743);
nor U1191 (N_1191,N_728,N_51);
nand U1192 (N_1192,N_683,N_9);
or U1193 (N_1193,N_19,N_79);
nand U1194 (N_1194,N_647,N_584);
nor U1195 (N_1195,N_698,N_657);
nand U1196 (N_1196,N_178,N_4);
and U1197 (N_1197,N_736,N_203);
nand U1198 (N_1198,N_585,N_356);
nand U1199 (N_1199,N_590,N_41);
nor U1200 (N_1200,N_541,N_397);
and U1201 (N_1201,N_670,N_388);
nand U1202 (N_1202,N_287,N_688);
and U1203 (N_1203,N_543,N_343);
or U1204 (N_1204,N_1,N_426);
or U1205 (N_1205,N_68,N_576);
or U1206 (N_1206,N_291,N_433);
or U1207 (N_1207,N_24,N_7);
or U1208 (N_1208,N_686,N_141);
or U1209 (N_1209,N_436,N_178);
nand U1210 (N_1210,N_679,N_8);
and U1211 (N_1211,N_213,N_65);
or U1212 (N_1212,N_524,N_123);
nor U1213 (N_1213,N_391,N_191);
nor U1214 (N_1214,N_259,N_331);
or U1215 (N_1215,N_684,N_563);
and U1216 (N_1216,N_441,N_338);
nand U1217 (N_1217,N_87,N_444);
or U1218 (N_1218,N_271,N_587);
and U1219 (N_1219,N_341,N_298);
nor U1220 (N_1220,N_317,N_110);
and U1221 (N_1221,N_252,N_687);
nor U1222 (N_1222,N_692,N_82);
nand U1223 (N_1223,N_566,N_71);
nand U1224 (N_1224,N_725,N_685);
or U1225 (N_1225,N_425,N_583);
and U1226 (N_1226,N_589,N_652);
nand U1227 (N_1227,N_192,N_98);
and U1228 (N_1228,N_533,N_440);
or U1229 (N_1229,N_111,N_161);
and U1230 (N_1230,N_467,N_486);
or U1231 (N_1231,N_397,N_120);
nand U1232 (N_1232,N_664,N_133);
and U1233 (N_1233,N_702,N_579);
and U1234 (N_1234,N_511,N_694);
or U1235 (N_1235,N_737,N_696);
nor U1236 (N_1236,N_4,N_388);
nor U1237 (N_1237,N_692,N_216);
nand U1238 (N_1238,N_43,N_431);
or U1239 (N_1239,N_362,N_3);
or U1240 (N_1240,N_636,N_642);
nand U1241 (N_1241,N_421,N_265);
nand U1242 (N_1242,N_577,N_165);
and U1243 (N_1243,N_346,N_340);
or U1244 (N_1244,N_175,N_204);
or U1245 (N_1245,N_148,N_620);
nand U1246 (N_1246,N_197,N_596);
or U1247 (N_1247,N_98,N_126);
or U1248 (N_1248,N_461,N_435);
or U1249 (N_1249,N_749,N_372);
or U1250 (N_1250,N_258,N_328);
or U1251 (N_1251,N_209,N_729);
and U1252 (N_1252,N_285,N_594);
or U1253 (N_1253,N_81,N_343);
nand U1254 (N_1254,N_730,N_164);
and U1255 (N_1255,N_483,N_38);
nand U1256 (N_1256,N_321,N_553);
nand U1257 (N_1257,N_747,N_184);
nor U1258 (N_1258,N_256,N_728);
nor U1259 (N_1259,N_707,N_2);
or U1260 (N_1260,N_4,N_36);
nor U1261 (N_1261,N_351,N_176);
xor U1262 (N_1262,N_483,N_692);
or U1263 (N_1263,N_63,N_663);
nor U1264 (N_1264,N_555,N_520);
and U1265 (N_1265,N_445,N_184);
or U1266 (N_1266,N_632,N_525);
nand U1267 (N_1267,N_128,N_20);
xor U1268 (N_1268,N_478,N_22);
nand U1269 (N_1269,N_415,N_12);
nand U1270 (N_1270,N_427,N_9);
nand U1271 (N_1271,N_360,N_144);
nor U1272 (N_1272,N_654,N_619);
and U1273 (N_1273,N_278,N_167);
or U1274 (N_1274,N_201,N_462);
nor U1275 (N_1275,N_144,N_740);
nand U1276 (N_1276,N_188,N_198);
nand U1277 (N_1277,N_155,N_576);
nor U1278 (N_1278,N_614,N_659);
nor U1279 (N_1279,N_258,N_290);
or U1280 (N_1280,N_256,N_557);
or U1281 (N_1281,N_262,N_618);
and U1282 (N_1282,N_717,N_467);
nor U1283 (N_1283,N_241,N_674);
and U1284 (N_1284,N_216,N_495);
nor U1285 (N_1285,N_705,N_501);
or U1286 (N_1286,N_267,N_722);
and U1287 (N_1287,N_129,N_7);
nor U1288 (N_1288,N_135,N_288);
nand U1289 (N_1289,N_447,N_74);
xor U1290 (N_1290,N_608,N_152);
nand U1291 (N_1291,N_207,N_645);
nor U1292 (N_1292,N_696,N_472);
nor U1293 (N_1293,N_347,N_282);
nor U1294 (N_1294,N_369,N_738);
nor U1295 (N_1295,N_523,N_231);
and U1296 (N_1296,N_589,N_638);
and U1297 (N_1297,N_90,N_372);
xor U1298 (N_1298,N_503,N_35);
and U1299 (N_1299,N_45,N_635);
nand U1300 (N_1300,N_547,N_383);
or U1301 (N_1301,N_110,N_91);
nand U1302 (N_1302,N_128,N_262);
xor U1303 (N_1303,N_665,N_635);
nand U1304 (N_1304,N_217,N_276);
and U1305 (N_1305,N_672,N_179);
or U1306 (N_1306,N_519,N_648);
and U1307 (N_1307,N_22,N_677);
or U1308 (N_1308,N_558,N_669);
nand U1309 (N_1309,N_723,N_370);
nand U1310 (N_1310,N_622,N_445);
or U1311 (N_1311,N_434,N_635);
nand U1312 (N_1312,N_197,N_666);
or U1313 (N_1313,N_407,N_110);
or U1314 (N_1314,N_680,N_461);
nand U1315 (N_1315,N_397,N_484);
nand U1316 (N_1316,N_745,N_284);
nand U1317 (N_1317,N_132,N_593);
nor U1318 (N_1318,N_262,N_506);
nand U1319 (N_1319,N_65,N_136);
and U1320 (N_1320,N_719,N_84);
and U1321 (N_1321,N_725,N_503);
nand U1322 (N_1322,N_171,N_666);
or U1323 (N_1323,N_607,N_670);
nand U1324 (N_1324,N_379,N_399);
nand U1325 (N_1325,N_552,N_733);
or U1326 (N_1326,N_561,N_343);
and U1327 (N_1327,N_588,N_15);
and U1328 (N_1328,N_609,N_132);
xnor U1329 (N_1329,N_670,N_225);
nor U1330 (N_1330,N_479,N_307);
and U1331 (N_1331,N_42,N_164);
and U1332 (N_1332,N_599,N_406);
and U1333 (N_1333,N_731,N_624);
or U1334 (N_1334,N_358,N_300);
xor U1335 (N_1335,N_382,N_363);
nand U1336 (N_1336,N_685,N_446);
nand U1337 (N_1337,N_366,N_216);
and U1338 (N_1338,N_195,N_337);
nand U1339 (N_1339,N_375,N_537);
nor U1340 (N_1340,N_69,N_228);
or U1341 (N_1341,N_535,N_719);
xor U1342 (N_1342,N_643,N_229);
or U1343 (N_1343,N_351,N_334);
nor U1344 (N_1344,N_106,N_5);
nor U1345 (N_1345,N_212,N_611);
or U1346 (N_1346,N_649,N_740);
and U1347 (N_1347,N_739,N_396);
nand U1348 (N_1348,N_76,N_534);
or U1349 (N_1349,N_164,N_294);
and U1350 (N_1350,N_410,N_37);
nand U1351 (N_1351,N_738,N_221);
nand U1352 (N_1352,N_249,N_91);
nand U1353 (N_1353,N_547,N_688);
and U1354 (N_1354,N_590,N_128);
nor U1355 (N_1355,N_326,N_235);
or U1356 (N_1356,N_361,N_629);
xnor U1357 (N_1357,N_224,N_540);
and U1358 (N_1358,N_410,N_507);
and U1359 (N_1359,N_396,N_219);
nor U1360 (N_1360,N_646,N_14);
and U1361 (N_1361,N_30,N_376);
nor U1362 (N_1362,N_351,N_135);
nor U1363 (N_1363,N_332,N_735);
nand U1364 (N_1364,N_95,N_482);
nor U1365 (N_1365,N_696,N_84);
or U1366 (N_1366,N_274,N_648);
and U1367 (N_1367,N_418,N_691);
or U1368 (N_1368,N_708,N_41);
nor U1369 (N_1369,N_138,N_522);
nand U1370 (N_1370,N_122,N_653);
or U1371 (N_1371,N_447,N_191);
or U1372 (N_1372,N_652,N_339);
and U1373 (N_1373,N_722,N_308);
and U1374 (N_1374,N_84,N_431);
nor U1375 (N_1375,N_631,N_437);
nor U1376 (N_1376,N_163,N_276);
and U1377 (N_1377,N_371,N_2);
nand U1378 (N_1378,N_144,N_248);
or U1379 (N_1379,N_489,N_134);
nand U1380 (N_1380,N_577,N_643);
and U1381 (N_1381,N_180,N_169);
and U1382 (N_1382,N_68,N_564);
nand U1383 (N_1383,N_652,N_349);
and U1384 (N_1384,N_22,N_162);
and U1385 (N_1385,N_568,N_253);
and U1386 (N_1386,N_578,N_729);
nor U1387 (N_1387,N_143,N_490);
or U1388 (N_1388,N_722,N_452);
nor U1389 (N_1389,N_82,N_99);
or U1390 (N_1390,N_744,N_468);
nor U1391 (N_1391,N_274,N_450);
nor U1392 (N_1392,N_329,N_216);
nand U1393 (N_1393,N_700,N_338);
or U1394 (N_1394,N_52,N_287);
or U1395 (N_1395,N_515,N_413);
nor U1396 (N_1396,N_602,N_339);
nor U1397 (N_1397,N_172,N_166);
and U1398 (N_1398,N_395,N_35);
or U1399 (N_1399,N_128,N_109);
and U1400 (N_1400,N_675,N_707);
and U1401 (N_1401,N_444,N_139);
nand U1402 (N_1402,N_594,N_262);
nor U1403 (N_1403,N_300,N_160);
nor U1404 (N_1404,N_533,N_14);
and U1405 (N_1405,N_523,N_499);
nor U1406 (N_1406,N_172,N_109);
nor U1407 (N_1407,N_508,N_434);
nand U1408 (N_1408,N_638,N_54);
nor U1409 (N_1409,N_287,N_41);
and U1410 (N_1410,N_197,N_276);
nand U1411 (N_1411,N_307,N_180);
or U1412 (N_1412,N_571,N_383);
nor U1413 (N_1413,N_238,N_511);
nor U1414 (N_1414,N_193,N_7);
or U1415 (N_1415,N_331,N_215);
nand U1416 (N_1416,N_469,N_596);
nand U1417 (N_1417,N_645,N_276);
nor U1418 (N_1418,N_661,N_603);
nand U1419 (N_1419,N_463,N_320);
nand U1420 (N_1420,N_112,N_512);
nand U1421 (N_1421,N_466,N_127);
nand U1422 (N_1422,N_392,N_275);
or U1423 (N_1423,N_121,N_655);
nor U1424 (N_1424,N_655,N_25);
nor U1425 (N_1425,N_374,N_702);
nor U1426 (N_1426,N_717,N_448);
or U1427 (N_1427,N_90,N_451);
and U1428 (N_1428,N_278,N_687);
nand U1429 (N_1429,N_271,N_235);
nand U1430 (N_1430,N_190,N_196);
nand U1431 (N_1431,N_415,N_163);
nor U1432 (N_1432,N_370,N_126);
nor U1433 (N_1433,N_746,N_303);
nand U1434 (N_1434,N_29,N_708);
xnor U1435 (N_1435,N_57,N_414);
and U1436 (N_1436,N_62,N_423);
nor U1437 (N_1437,N_160,N_395);
nand U1438 (N_1438,N_211,N_350);
and U1439 (N_1439,N_295,N_506);
and U1440 (N_1440,N_689,N_411);
and U1441 (N_1441,N_462,N_393);
nor U1442 (N_1442,N_518,N_651);
and U1443 (N_1443,N_569,N_82);
nand U1444 (N_1444,N_179,N_257);
or U1445 (N_1445,N_253,N_579);
nor U1446 (N_1446,N_256,N_666);
nand U1447 (N_1447,N_369,N_218);
or U1448 (N_1448,N_463,N_468);
and U1449 (N_1449,N_366,N_520);
and U1450 (N_1450,N_535,N_317);
and U1451 (N_1451,N_576,N_430);
nand U1452 (N_1452,N_223,N_547);
or U1453 (N_1453,N_441,N_247);
and U1454 (N_1454,N_391,N_212);
and U1455 (N_1455,N_59,N_239);
nand U1456 (N_1456,N_641,N_741);
and U1457 (N_1457,N_376,N_586);
nand U1458 (N_1458,N_632,N_560);
xnor U1459 (N_1459,N_600,N_347);
and U1460 (N_1460,N_520,N_632);
and U1461 (N_1461,N_693,N_212);
nor U1462 (N_1462,N_170,N_112);
nor U1463 (N_1463,N_688,N_136);
and U1464 (N_1464,N_600,N_214);
or U1465 (N_1465,N_617,N_692);
nor U1466 (N_1466,N_471,N_589);
or U1467 (N_1467,N_375,N_268);
and U1468 (N_1468,N_4,N_554);
nand U1469 (N_1469,N_184,N_154);
nor U1470 (N_1470,N_280,N_688);
nor U1471 (N_1471,N_566,N_692);
nand U1472 (N_1472,N_220,N_255);
nand U1473 (N_1473,N_706,N_216);
and U1474 (N_1474,N_498,N_84);
nor U1475 (N_1475,N_601,N_381);
nand U1476 (N_1476,N_460,N_161);
or U1477 (N_1477,N_699,N_642);
nor U1478 (N_1478,N_389,N_21);
nand U1479 (N_1479,N_45,N_224);
nor U1480 (N_1480,N_296,N_371);
nor U1481 (N_1481,N_222,N_526);
and U1482 (N_1482,N_581,N_610);
or U1483 (N_1483,N_632,N_582);
nand U1484 (N_1484,N_62,N_106);
or U1485 (N_1485,N_558,N_684);
and U1486 (N_1486,N_7,N_696);
nor U1487 (N_1487,N_466,N_11);
nand U1488 (N_1488,N_556,N_171);
nand U1489 (N_1489,N_81,N_201);
or U1490 (N_1490,N_732,N_493);
nand U1491 (N_1491,N_749,N_568);
nand U1492 (N_1492,N_666,N_0);
and U1493 (N_1493,N_709,N_115);
nor U1494 (N_1494,N_384,N_234);
nand U1495 (N_1495,N_337,N_77);
and U1496 (N_1496,N_678,N_124);
or U1497 (N_1497,N_261,N_505);
nor U1498 (N_1498,N_38,N_549);
nand U1499 (N_1499,N_243,N_295);
and U1500 (N_1500,N_757,N_1322);
or U1501 (N_1501,N_765,N_793);
or U1502 (N_1502,N_957,N_760);
nor U1503 (N_1503,N_785,N_798);
or U1504 (N_1504,N_1102,N_1338);
and U1505 (N_1505,N_1137,N_890);
or U1506 (N_1506,N_1491,N_886);
and U1507 (N_1507,N_1301,N_1429);
or U1508 (N_1508,N_1187,N_1100);
nand U1509 (N_1509,N_1479,N_1198);
or U1510 (N_1510,N_998,N_1378);
nand U1511 (N_1511,N_900,N_1110);
nand U1512 (N_1512,N_1190,N_1360);
nor U1513 (N_1513,N_1080,N_1094);
nor U1514 (N_1514,N_825,N_887);
or U1515 (N_1515,N_1475,N_806);
and U1516 (N_1516,N_1457,N_1087);
nor U1517 (N_1517,N_849,N_939);
xnor U1518 (N_1518,N_1139,N_1085);
and U1519 (N_1519,N_927,N_1395);
nand U1520 (N_1520,N_770,N_1040);
or U1521 (N_1521,N_788,N_1052);
and U1522 (N_1522,N_842,N_1202);
or U1523 (N_1523,N_923,N_846);
or U1524 (N_1524,N_1363,N_1297);
nor U1525 (N_1525,N_1465,N_895);
nor U1526 (N_1526,N_1261,N_873);
and U1527 (N_1527,N_1304,N_979);
and U1528 (N_1528,N_1096,N_1462);
and U1529 (N_1529,N_876,N_1369);
nor U1530 (N_1530,N_1163,N_1485);
nor U1531 (N_1531,N_1207,N_1061);
nand U1532 (N_1532,N_1263,N_1490);
nand U1533 (N_1533,N_1018,N_801);
or U1534 (N_1534,N_1302,N_1318);
nor U1535 (N_1535,N_1006,N_1436);
xor U1536 (N_1536,N_855,N_1313);
and U1537 (N_1537,N_950,N_764);
or U1538 (N_1538,N_1141,N_1404);
nand U1539 (N_1539,N_1142,N_1168);
or U1540 (N_1540,N_815,N_1218);
or U1541 (N_1541,N_936,N_1420);
and U1542 (N_1542,N_1192,N_1216);
or U1543 (N_1543,N_1194,N_1160);
nor U1544 (N_1544,N_1219,N_1407);
or U1545 (N_1545,N_1396,N_1265);
nand U1546 (N_1546,N_1138,N_1430);
or U1547 (N_1547,N_903,N_1268);
or U1548 (N_1548,N_1405,N_1489);
and U1549 (N_1549,N_1306,N_1358);
and U1550 (N_1550,N_924,N_1081);
nor U1551 (N_1551,N_915,N_1346);
xnor U1552 (N_1552,N_1258,N_1185);
nor U1553 (N_1553,N_1175,N_754);
nor U1554 (N_1554,N_1010,N_1364);
nor U1555 (N_1555,N_1337,N_1329);
and U1556 (N_1556,N_879,N_1482);
xor U1557 (N_1557,N_852,N_1051);
or U1558 (N_1558,N_1298,N_916);
and U1559 (N_1559,N_906,N_938);
nor U1560 (N_1560,N_1264,N_1325);
or U1561 (N_1561,N_1031,N_816);
nand U1562 (N_1562,N_1345,N_1312);
and U1563 (N_1563,N_860,N_1365);
or U1564 (N_1564,N_791,N_1162);
and U1565 (N_1565,N_1048,N_1356);
and U1566 (N_1566,N_1097,N_1158);
and U1567 (N_1567,N_902,N_1106);
nand U1568 (N_1568,N_1382,N_780);
nand U1569 (N_1569,N_1497,N_1022);
nor U1570 (N_1570,N_1201,N_913);
or U1571 (N_1571,N_1154,N_1336);
nand U1572 (N_1572,N_1353,N_1488);
nor U1573 (N_1573,N_1444,N_1251);
or U1574 (N_1574,N_1438,N_1361);
or U1575 (N_1575,N_756,N_1038);
and U1576 (N_1576,N_982,N_953);
nand U1577 (N_1577,N_1045,N_1245);
or U1578 (N_1578,N_1419,N_1088);
or U1579 (N_1579,N_776,N_1406);
xor U1580 (N_1580,N_1240,N_1370);
nor U1581 (N_1581,N_1493,N_1053);
nand U1582 (N_1582,N_922,N_966);
nand U1583 (N_1583,N_897,N_755);
nor U1584 (N_1584,N_1324,N_819);
and U1585 (N_1585,N_1288,N_919);
nand U1586 (N_1586,N_858,N_1256);
or U1587 (N_1587,N_1095,N_1310);
nand U1588 (N_1588,N_1205,N_1411);
nor U1589 (N_1589,N_1077,N_1208);
nor U1590 (N_1590,N_1422,N_1450);
and U1591 (N_1591,N_975,N_993);
or U1592 (N_1592,N_821,N_1432);
and U1593 (N_1593,N_1357,N_1026);
nor U1594 (N_1594,N_1209,N_1127);
nand U1595 (N_1595,N_1233,N_1123);
nand U1596 (N_1596,N_1033,N_848);
nand U1597 (N_1597,N_1147,N_1066);
nor U1598 (N_1598,N_1107,N_910);
nand U1599 (N_1599,N_1311,N_1266);
and U1600 (N_1600,N_1200,N_983);
nand U1601 (N_1601,N_847,N_1355);
or U1602 (N_1602,N_1428,N_1433);
and U1603 (N_1603,N_838,N_805);
nand U1604 (N_1604,N_1440,N_1291);
and U1605 (N_1605,N_1449,N_961);
and U1606 (N_1606,N_926,N_991);
nand U1607 (N_1607,N_1156,N_1276);
and U1608 (N_1608,N_1165,N_996);
or U1609 (N_1609,N_809,N_934);
nor U1610 (N_1610,N_1002,N_1435);
nand U1611 (N_1611,N_1280,N_834);
and U1612 (N_1612,N_912,N_1159);
or U1613 (N_1613,N_1410,N_954);
or U1614 (N_1614,N_1328,N_1173);
nand U1615 (N_1615,N_1034,N_1003);
or U1616 (N_1616,N_1460,N_972);
nor U1617 (N_1617,N_952,N_1471);
and U1618 (N_1618,N_1001,N_1092);
nand U1619 (N_1619,N_1134,N_1055);
and U1620 (N_1620,N_908,N_813);
nor U1621 (N_1621,N_1029,N_1012);
nand U1622 (N_1622,N_1290,N_971);
nand U1623 (N_1623,N_1009,N_1443);
or U1624 (N_1624,N_937,N_837);
or U1625 (N_1625,N_1494,N_1456);
and U1626 (N_1626,N_1400,N_1191);
nand U1627 (N_1627,N_1184,N_851);
and U1628 (N_1628,N_1255,N_856);
nand U1629 (N_1629,N_874,N_1466);
nand U1630 (N_1630,N_1445,N_1149);
or U1631 (N_1631,N_835,N_1319);
nand U1632 (N_1632,N_968,N_1119);
nand U1633 (N_1633,N_1238,N_1180);
or U1634 (N_1634,N_1343,N_750);
or U1635 (N_1635,N_1469,N_1109);
nand U1636 (N_1636,N_1124,N_1082);
and U1637 (N_1637,N_1118,N_1412);
nor U1638 (N_1638,N_1354,N_1246);
nand U1639 (N_1639,N_973,N_826);
nor U1640 (N_1640,N_1321,N_985);
xor U1641 (N_1641,N_896,N_877);
or U1642 (N_1642,N_767,N_1197);
nand U1643 (N_1643,N_1499,N_1453);
and U1644 (N_1644,N_1305,N_1316);
and U1645 (N_1645,N_911,N_1376);
and U1646 (N_1646,N_1212,N_1043);
nand U1647 (N_1647,N_828,N_1065);
nor U1648 (N_1648,N_1387,N_830);
and U1649 (N_1649,N_1332,N_931);
and U1650 (N_1650,N_1252,N_967);
nor U1651 (N_1651,N_1495,N_1386);
nor U1652 (N_1652,N_841,N_1307);
nand U1653 (N_1653,N_1086,N_889);
or U1654 (N_1654,N_1063,N_1274);
or U1655 (N_1655,N_1069,N_1078);
or U1656 (N_1656,N_1232,N_1132);
nor U1657 (N_1657,N_1249,N_1446);
xor U1658 (N_1658,N_1373,N_1007);
and U1659 (N_1659,N_1186,N_1015);
nor U1660 (N_1660,N_789,N_905);
nand U1661 (N_1661,N_1047,N_1220);
nor U1662 (N_1662,N_786,N_1064);
nor U1663 (N_1663,N_758,N_892);
and U1664 (N_1664,N_1108,N_868);
and U1665 (N_1665,N_945,N_1380);
nor U1666 (N_1666,N_1222,N_907);
nand U1667 (N_1667,N_1211,N_1388);
and U1668 (N_1668,N_1027,N_1231);
nor U1669 (N_1669,N_883,N_784);
or U1670 (N_1670,N_1042,N_1021);
and U1671 (N_1671,N_1215,N_1442);
or U1672 (N_1672,N_1224,N_1103);
nor U1673 (N_1673,N_751,N_917);
nand U1674 (N_1674,N_824,N_1320);
and U1675 (N_1675,N_942,N_984);
nand U1676 (N_1676,N_1121,N_1285);
or U1677 (N_1677,N_810,N_1056);
nand U1678 (N_1678,N_1384,N_1303);
or U1679 (N_1679,N_843,N_762);
nor U1680 (N_1680,N_965,N_1035);
nor U1681 (N_1681,N_1114,N_988);
nand U1682 (N_1682,N_761,N_955);
or U1683 (N_1683,N_1403,N_1133);
nand U1684 (N_1684,N_1176,N_795);
nand U1685 (N_1685,N_1111,N_866);
and U1686 (N_1686,N_947,N_850);
nor U1687 (N_1687,N_1071,N_1199);
and U1688 (N_1688,N_1352,N_769);
and U1689 (N_1689,N_999,N_1293);
nand U1690 (N_1690,N_1178,N_1225);
nor U1691 (N_1691,N_1214,N_794);
and U1692 (N_1692,N_959,N_1230);
and U1693 (N_1693,N_1447,N_1183);
nor U1694 (N_1694,N_827,N_1130);
or U1695 (N_1695,N_1389,N_1401);
or U1696 (N_1696,N_1213,N_1496);
or U1697 (N_1697,N_1284,N_1234);
nor U1698 (N_1698,N_1135,N_1339);
nor U1699 (N_1699,N_1177,N_1236);
and U1700 (N_1700,N_1451,N_1260);
nor U1701 (N_1701,N_1070,N_1253);
nand U1702 (N_1702,N_882,N_1166);
nand U1703 (N_1703,N_1367,N_759);
or U1704 (N_1704,N_1351,N_1275);
nor U1705 (N_1705,N_1289,N_1068);
and U1706 (N_1706,N_1333,N_1282);
nand U1707 (N_1707,N_814,N_1459);
or U1708 (N_1708,N_875,N_901);
or U1709 (N_1709,N_1072,N_822);
or U1710 (N_1710,N_1146,N_1145);
nor U1711 (N_1711,N_914,N_1241);
or U1712 (N_1712,N_1448,N_980);
and U1713 (N_1713,N_1417,N_1148);
or U1714 (N_1714,N_1366,N_832);
and U1715 (N_1715,N_1383,N_1458);
nor U1716 (N_1716,N_777,N_1091);
and U1717 (N_1717,N_1487,N_925);
or U1718 (N_1718,N_1331,N_783);
nand U1719 (N_1719,N_1076,N_948);
or U1720 (N_1720,N_1464,N_1182);
or U1721 (N_1721,N_1425,N_1084);
nor U1722 (N_1722,N_1083,N_1299);
or U1723 (N_1723,N_1414,N_811);
nand U1724 (N_1724,N_1480,N_1437);
nor U1725 (N_1725,N_1334,N_1402);
and U1726 (N_1726,N_1287,N_808);
and U1727 (N_1727,N_1409,N_1242);
nand U1728 (N_1728,N_768,N_943);
and U1729 (N_1729,N_958,N_909);
nand U1730 (N_1730,N_1171,N_1195);
and U1731 (N_1731,N_899,N_1079);
nand U1732 (N_1732,N_986,N_1424);
or U1733 (N_1733,N_1292,N_976);
and U1734 (N_1734,N_1413,N_1120);
nor U1735 (N_1735,N_992,N_1140);
nor U1736 (N_1736,N_1004,N_820);
nand U1737 (N_1737,N_987,N_1016);
and U1738 (N_1738,N_978,N_1172);
or U1739 (N_1739,N_779,N_1294);
nand U1740 (N_1740,N_1341,N_1326);
nor U1741 (N_1741,N_823,N_1005);
or U1742 (N_1742,N_1269,N_1093);
nor U1743 (N_1743,N_1032,N_960);
nand U1744 (N_1744,N_949,N_1481);
nand U1745 (N_1745,N_1206,N_1327);
nand U1746 (N_1746,N_904,N_1024);
or U1747 (N_1747,N_1267,N_1073);
nor U1748 (N_1748,N_773,N_1335);
nor U1749 (N_1749,N_962,N_1028);
and U1750 (N_1750,N_1210,N_1181);
xnor U1751 (N_1751,N_1421,N_970);
nand U1752 (N_1752,N_1478,N_833);
nor U1753 (N_1753,N_1270,N_1074);
and U1754 (N_1754,N_1008,N_990);
or U1755 (N_1755,N_1483,N_891);
nand U1756 (N_1756,N_1467,N_1362);
nand U1757 (N_1757,N_752,N_1330);
and U1758 (N_1758,N_885,N_796);
or U1759 (N_1759,N_1309,N_1011);
nor U1760 (N_1760,N_1323,N_1125);
and U1761 (N_1761,N_862,N_981);
nor U1762 (N_1762,N_1427,N_1461);
and U1763 (N_1763,N_766,N_1039);
or U1764 (N_1764,N_1271,N_1030);
nor U1765 (N_1765,N_1023,N_1342);
nor U1766 (N_1766,N_864,N_1227);
nand U1767 (N_1767,N_1434,N_1473);
nor U1768 (N_1768,N_804,N_929);
nand U1769 (N_1769,N_1189,N_1057);
and U1770 (N_1770,N_1101,N_1000);
nor U1771 (N_1771,N_865,N_944);
and U1772 (N_1772,N_836,N_994);
nand U1773 (N_1773,N_1398,N_799);
or U1774 (N_1774,N_1243,N_1228);
or U1775 (N_1775,N_1196,N_863);
or U1776 (N_1776,N_1277,N_829);
or U1777 (N_1777,N_1375,N_1239);
or U1778 (N_1778,N_1164,N_1037);
nand U1779 (N_1779,N_956,N_782);
nand U1780 (N_1780,N_1454,N_1143);
or U1781 (N_1781,N_869,N_1050);
nand U1782 (N_1782,N_1116,N_921);
xor U1783 (N_1783,N_1468,N_878);
nor U1784 (N_1784,N_1060,N_964);
nand U1785 (N_1785,N_1167,N_1408);
nor U1786 (N_1786,N_1278,N_1283);
xor U1787 (N_1787,N_1151,N_1019);
nand U1788 (N_1788,N_1392,N_1144);
nand U1789 (N_1789,N_1439,N_840);
nand U1790 (N_1790,N_1296,N_802);
nand U1791 (N_1791,N_974,N_918);
nor U1792 (N_1792,N_1498,N_1344);
or U1793 (N_1793,N_1372,N_1455);
or U1794 (N_1794,N_1046,N_1098);
nand U1795 (N_1795,N_1157,N_1477);
nand U1796 (N_1796,N_1020,N_818);
nor U1797 (N_1797,N_1090,N_1416);
nand U1798 (N_1798,N_1262,N_867);
or U1799 (N_1799,N_1415,N_1394);
and U1800 (N_1800,N_807,N_1169);
nand U1801 (N_1801,N_845,N_790);
or U1802 (N_1802,N_1013,N_920);
nor U1803 (N_1803,N_1131,N_1247);
or U1804 (N_1804,N_817,N_1221);
nor U1805 (N_1805,N_1126,N_1426);
or U1806 (N_1806,N_1188,N_1431);
and U1807 (N_1807,N_1463,N_1397);
nor U1808 (N_1808,N_1272,N_1244);
or U1809 (N_1809,N_1281,N_932);
or U1810 (N_1810,N_1203,N_894);
nor U1811 (N_1811,N_1152,N_1044);
nor U1812 (N_1812,N_951,N_1472);
and U1813 (N_1813,N_1025,N_1254);
and U1814 (N_1814,N_941,N_1286);
or U1815 (N_1815,N_1054,N_1014);
nand U1816 (N_1816,N_933,N_1223);
nor U1817 (N_1817,N_1229,N_1170);
and U1818 (N_1818,N_1340,N_774);
nand U1819 (N_1819,N_1374,N_1391);
nand U1820 (N_1820,N_963,N_854);
nand U1821 (N_1821,N_1476,N_1381);
and U1822 (N_1822,N_1153,N_1058);
and U1823 (N_1823,N_1259,N_1105);
nand U1824 (N_1824,N_871,N_1390);
nor U1825 (N_1825,N_839,N_1150);
nand U1826 (N_1826,N_1204,N_803);
nand U1827 (N_1827,N_1347,N_1250);
or U1828 (N_1828,N_1036,N_893);
and U1829 (N_1829,N_1129,N_1122);
nand U1830 (N_1830,N_1041,N_1295);
or U1831 (N_1831,N_1075,N_1368);
or U1832 (N_1832,N_1452,N_1226);
nor U1833 (N_1833,N_1441,N_1486);
or U1834 (N_1834,N_861,N_888);
or U1835 (N_1835,N_1349,N_1235);
nor U1836 (N_1836,N_792,N_772);
and U1837 (N_1837,N_969,N_797);
xor U1838 (N_1838,N_1308,N_1161);
nand U1839 (N_1839,N_1371,N_1492);
nand U1840 (N_1840,N_1273,N_753);
or U1841 (N_1841,N_1359,N_1067);
nor U1842 (N_1842,N_881,N_995);
nand U1843 (N_1843,N_1049,N_1350);
nand U1844 (N_1844,N_946,N_853);
nor U1845 (N_1845,N_831,N_898);
and U1846 (N_1846,N_781,N_1279);
nand U1847 (N_1847,N_1136,N_1117);
and U1848 (N_1848,N_1315,N_930);
or U1849 (N_1849,N_1174,N_997);
nor U1850 (N_1850,N_884,N_1237);
or U1851 (N_1851,N_1317,N_1484);
or U1852 (N_1852,N_1393,N_1257);
or U1853 (N_1853,N_812,N_763);
and U1854 (N_1854,N_1099,N_800);
or U1855 (N_1855,N_1385,N_1470);
nor U1856 (N_1856,N_1474,N_1248);
nor U1857 (N_1857,N_1104,N_977);
or U1858 (N_1858,N_1217,N_1115);
or U1859 (N_1859,N_880,N_1423);
or U1860 (N_1860,N_1314,N_1300);
nor U1861 (N_1861,N_859,N_928);
nor U1862 (N_1862,N_1179,N_872);
or U1863 (N_1863,N_1089,N_787);
or U1864 (N_1864,N_1113,N_1193);
or U1865 (N_1865,N_844,N_1348);
xnor U1866 (N_1866,N_1155,N_857);
and U1867 (N_1867,N_778,N_1377);
and U1868 (N_1868,N_1418,N_1112);
nor U1869 (N_1869,N_1379,N_771);
nand U1870 (N_1870,N_1128,N_1062);
or U1871 (N_1871,N_870,N_940);
nor U1872 (N_1872,N_935,N_989);
nand U1873 (N_1873,N_1017,N_775);
and U1874 (N_1874,N_1399,N_1059);
nor U1875 (N_1875,N_775,N_1365);
and U1876 (N_1876,N_1293,N_1485);
nand U1877 (N_1877,N_1339,N_1215);
and U1878 (N_1878,N_1488,N_987);
nor U1879 (N_1879,N_1003,N_1017);
and U1880 (N_1880,N_1442,N_1223);
nor U1881 (N_1881,N_1111,N_1037);
or U1882 (N_1882,N_983,N_1499);
or U1883 (N_1883,N_859,N_965);
nand U1884 (N_1884,N_1157,N_947);
nor U1885 (N_1885,N_981,N_1293);
nor U1886 (N_1886,N_821,N_1100);
and U1887 (N_1887,N_779,N_943);
and U1888 (N_1888,N_795,N_1222);
nor U1889 (N_1889,N_1401,N_1361);
nand U1890 (N_1890,N_1121,N_1145);
nand U1891 (N_1891,N_1456,N_1485);
or U1892 (N_1892,N_807,N_1228);
and U1893 (N_1893,N_1238,N_756);
or U1894 (N_1894,N_1282,N_1065);
and U1895 (N_1895,N_1060,N_1223);
and U1896 (N_1896,N_1201,N_1173);
nand U1897 (N_1897,N_1315,N_811);
nor U1898 (N_1898,N_1035,N_1218);
nor U1899 (N_1899,N_1299,N_862);
or U1900 (N_1900,N_1150,N_768);
nor U1901 (N_1901,N_1142,N_1117);
nor U1902 (N_1902,N_802,N_1416);
or U1903 (N_1903,N_1402,N_1066);
nor U1904 (N_1904,N_1082,N_1461);
and U1905 (N_1905,N_1471,N_953);
nor U1906 (N_1906,N_1003,N_1128);
nor U1907 (N_1907,N_819,N_1276);
and U1908 (N_1908,N_1043,N_966);
nor U1909 (N_1909,N_1387,N_1080);
nor U1910 (N_1910,N_1065,N_1183);
and U1911 (N_1911,N_1436,N_1325);
and U1912 (N_1912,N_849,N_1128);
or U1913 (N_1913,N_903,N_884);
nor U1914 (N_1914,N_1143,N_868);
xor U1915 (N_1915,N_846,N_1231);
nor U1916 (N_1916,N_767,N_1162);
or U1917 (N_1917,N_1258,N_939);
nor U1918 (N_1918,N_1250,N_1133);
or U1919 (N_1919,N_1064,N_1218);
or U1920 (N_1920,N_785,N_1224);
and U1921 (N_1921,N_1484,N_1139);
or U1922 (N_1922,N_1111,N_1078);
nor U1923 (N_1923,N_1455,N_908);
or U1924 (N_1924,N_998,N_1309);
nor U1925 (N_1925,N_1108,N_1313);
or U1926 (N_1926,N_1447,N_1244);
nand U1927 (N_1927,N_1479,N_1420);
nor U1928 (N_1928,N_854,N_755);
nor U1929 (N_1929,N_1136,N_903);
xor U1930 (N_1930,N_1141,N_1092);
nor U1931 (N_1931,N_1059,N_1293);
and U1932 (N_1932,N_931,N_1446);
nor U1933 (N_1933,N_1417,N_1068);
nand U1934 (N_1934,N_1448,N_1353);
and U1935 (N_1935,N_993,N_864);
nor U1936 (N_1936,N_960,N_1426);
and U1937 (N_1937,N_1445,N_1215);
nor U1938 (N_1938,N_1086,N_897);
nor U1939 (N_1939,N_1394,N_1053);
nand U1940 (N_1940,N_1415,N_1312);
or U1941 (N_1941,N_1240,N_1467);
or U1942 (N_1942,N_1445,N_865);
or U1943 (N_1943,N_1095,N_1432);
and U1944 (N_1944,N_1298,N_884);
or U1945 (N_1945,N_852,N_1120);
nand U1946 (N_1946,N_1014,N_1435);
nand U1947 (N_1947,N_914,N_1362);
nor U1948 (N_1948,N_1257,N_812);
nand U1949 (N_1949,N_1428,N_1143);
nor U1950 (N_1950,N_1334,N_1341);
nor U1951 (N_1951,N_1145,N_851);
or U1952 (N_1952,N_1250,N_831);
or U1953 (N_1953,N_1010,N_1293);
nand U1954 (N_1954,N_1170,N_1240);
or U1955 (N_1955,N_1355,N_1226);
nor U1956 (N_1956,N_1375,N_1150);
nor U1957 (N_1957,N_847,N_1097);
nor U1958 (N_1958,N_1278,N_1435);
and U1959 (N_1959,N_821,N_868);
or U1960 (N_1960,N_1445,N_945);
or U1961 (N_1961,N_773,N_1018);
or U1962 (N_1962,N_1208,N_1313);
nand U1963 (N_1963,N_1102,N_1460);
nor U1964 (N_1964,N_1234,N_1429);
and U1965 (N_1965,N_1068,N_1155);
nor U1966 (N_1966,N_975,N_793);
or U1967 (N_1967,N_940,N_1421);
or U1968 (N_1968,N_1234,N_1164);
and U1969 (N_1969,N_1322,N_1097);
xor U1970 (N_1970,N_846,N_1032);
nand U1971 (N_1971,N_1432,N_1051);
nor U1972 (N_1972,N_793,N_1405);
nor U1973 (N_1973,N_948,N_1408);
or U1974 (N_1974,N_878,N_961);
nand U1975 (N_1975,N_1035,N_1438);
nand U1976 (N_1976,N_1093,N_1404);
and U1977 (N_1977,N_848,N_932);
nor U1978 (N_1978,N_1008,N_926);
and U1979 (N_1979,N_1083,N_1404);
nand U1980 (N_1980,N_917,N_1061);
nand U1981 (N_1981,N_1403,N_1117);
nor U1982 (N_1982,N_1135,N_943);
or U1983 (N_1983,N_905,N_1374);
or U1984 (N_1984,N_1346,N_1211);
or U1985 (N_1985,N_782,N_1355);
nor U1986 (N_1986,N_1127,N_1027);
and U1987 (N_1987,N_1147,N_886);
nor U1988 (N_1988,N_1012,N_1150);
and U1989 (N_1989,N_1459,N_1295);
nor U1990 (N_1990,N_1156,N_870);
nand U1991 (N_1991,N_1400,N_900);
or U1992 (N_1992,N_944,N_976);
nand U1993 (N_1993,N_1073,N_1206);
nand U1994 (N_1994,N_1109,N_1074);
and U1995 (N_1995,N_813,N_1262);
nor U1996 (N_1996,N_1118,N_907);
nand U1997 (N_1997,N_751,N_1319);
nand U1998 (N_1998,N_1288,N_757);
or U1999 (N_1999,N_1220,N_1363);
nor U2000 (N_2000,N_1250,N_1359);
nand U2001 (N_2001,N_1362,N_1113);
nor U2002 (N_2002,N_817,N_1089);
nand U2003 (N_2003,N_1094,N_1058);
and U2004 (N_2004,N_1079,N_1154);
and U2005 (N_2005,N_930,N_1062);
or U2006 (N_2006,N_1050,N_1035);
or U2007 (N_2007,N_874,N_754);
xnor U2008 (N_2008,N_845,N_1315);
nand U2009 (N_2009,N_1345,N_1223);
nand U2010 (N_2010,N_967,N_972);
or U2011 (N_2011,N_994,N_1156);
nor U2012 (N_2012,N_1277,N_1326);
or U2013 (N_2013,N_1024,N_785);
nor U2014 (N_2014,N_1177,N_1460);
nor U2015 (N_2015,N_1334,N_1220);
nor U2016 (N_2016,N_1135,N_934);
or U2017 (N_2017,N_1324,N_1317);
and U2018 (N_2018,N_1491,N_750);
or U2019 (N_2019,N_1043,N_892);
and U2020 (N_2020,N_1358,N_1459);
nand U2021 (N_2021,N_1303,N_959);
and U2022 (N_2022,N_1179,N_1106);
nor U2023 (N_2023,N_1234,N_828);
nand U2024 (N_2024,N_764,N_931);
and U2025 (N_2025,N_1139,N_793);
and U2026 (N_2026,N_1203,N_1372);
nand U2027 (N_2027,N_835,N_1437);
nand U2028 (N_2028,N_1382,N_1342);
nand U2029 (N_2029,N_1401,N_1123);
nand U2030 (N_2030,N_987,N_959);
or U2031 (N_2031,N_1367,N_1365);
nand U2032 (N_2032,N_952,N_1095);
xnor U2033 (N_2033,N_1242,N_1218);
and U2034 (N_2034,N_948,N_1237);
nor U2035 (N_2035,N_1072,N_1142);
and U2036 (N_2036,N_1045,N_917);
and U2037 (N_2037,N_1479,N_775);
xnor U2038 (N_2038,N_1433,N_820);
and U2039 (N_2039,N_965,N_1468);
and U2040 (N_2040,N_1446,N_1258);
nor U2041 (N_2041,N_980,N_1169);
nor U2042 (N_2042,N_882,N_1126);
nand U2043 (N_2043,N_774,N_787);
xor U2044 (N_2044,N_764,N_1037);
and U2045 (N_2045,N_1256,N_1401);
xnor U2046 (N_2046,N_1287,N_1229);
nor U2047 (N_2047,N_1174,N_1201);
or U2048 (N_2048,N_1105,N_1035);
or U2049 (N_2049,N_800,N_909);
nor U2050 (N_2050,N_1367,N_816);
or U2051 (N_2051,N_1146,N_1188);
nor U2052 (N_2052,N_1084,N_1261);
and U2053 (N_2053,N_1422,N_774);
nor U2054 (N_2054,N_1441,N_1225);
xnor U2055 (N_2055,N_1201,N_833);
nand U2056 (N_2056,N_1394,N_761);
xnor U2057 (N_2057,N_758,N_995);
nor U2058 (N_2058,N_939,N_1076);
nand U2059 (N_2059,N_1451,N_845);
or U2060 (N_2060,N_1307,N_1039);
nand U2061 (N_2061,N_968,N_957);
nor U2062 (N_2062,N_1337,N_1066);
and U2063 (N_2063,N_1427,N_1098);
nand U2064 (N_2064,N_798,N_1432);
and U2065 (N_2065,N_1343,N_1199);
nand U2066 (N_2066,N_1226,N_761);
nor U2067 (N_2067,N_907,N_872);
and U2068 (N_2068,N_1035,N_1032);
nor U2069 (N_2069,N_962,N_819);
nor U2070 (N_2070,N_1353,N_941);
nand U2071 (N_2071,N_1277,N_1075);
nand U2072 (N_2072,N_1070,N_956);
nand U2073 (N_2073,N_1195,N_779);
nor U2074 (N_2074,N_788,N_801);
nand U2075 (N_2075,N_896,N_1084);
nand U2076 (N_2076,N_1160,N_1077);
xor U2077 (N_2077,N_1180,N_805);
nand U2078 (N_2078,N_1140,N_1303);
or U2079 (N_2079,N_847,N_1119);
nor U2080 (N_2080,N_1133,N_1015);
nor U2081 (N_2081,N_1015,N_1339);
nor U2082 (N_2082,N_854,N_1281);
or U2083 (N_2083,N_1145,N_1232);
nor U2084 (N_2084,N_1473,N_1236);
or U2085 (N_2085,N_1288,N_1471);
xnor U2086 (N_2086,N_1369,N_966);
or U2087 (N_2087,N_1345,N_865);
nand U2088 (N_2088,N_1428,N_921);
and U2089 (N_2089,N_1175,N_1205);
and U2090 (N_2090,N_1242,N_1435);
or U2091 (N_2091,N_1105,N_1069);
and U2092 (N_2092,N_1180,N_1132);
or U2093 (N_2093,N_1486,N_1398);
nor U2094 (N_2094,N_774,N_1445);
nor U2095 (N_2095,N_1342,N_1153);
nor U2096 (N_2096,N_1448,N_1432);
or U2097 (N_2097,N_1363,N_1089);
or U2098 (N_2098,N_947,N_1404);
nand U2099 (N_2099,N_1341,N_1080);
and U2100 (N_2100,N_1257,N_841);
nand U2101 (N_2101,N_1402,N_770);
and U2102 (N_2102,N_1131,N_1068);
nor U2103 (N_2103,N_1091,N_1113);
nand U2104 (N_2104,N_1247,N_1166);
and U2105 (N_2105,N_860,N_966);
and U2106 (N_2106,N_1454,N_1135);
nand U2107 (N_2107,N_1030,N_837);
xor U2108 (N_2108,N_851,N_1431);
or U2109 (N_2109,N_990,N_1115);
nand U2110 (N_2110,N_1302,N_751);
nor U2111 (N_2111,N_1387,N_1494);
or U2112 (N_2112,N_779,N_822);
nor U2113 (N_2113,N_1128,N_946);
nand U2114 (N_2114,N_999,N_1391);
or U2115 (N_2115,N_1336,N_1283);
and U2116 (N_2116,N_1247,N_896);
nand U2117 (N_2117,N_1224,N_1317);
and U2118 (N_2118,N_1408,N_1182);
or U2119 (N_2119,N_1224,N_769);
nand U2120 (N_2120,N_1328,N_1160);
or U2121 (N_2121,N_1354,N_939);
nand U2122 (N_2122,N_988,N_1216);
or U2123 (N_2123,N_1046,N_1190);
xnor U2124 (N_2124,N_1003,N_1135);
or U2125 (N_2125,N_1317,N_916);
nor U2126 (N_2126,N_932,N_1006);
or U2127 (N_2127,N_1040,N_873);
nor U2128 (N_2128,N_880,N_1202);
nor U2129 (N_2129,N_849,N_1390);
nor U2130 (N_2130,N_1485,N_1125);
or U2131 (N_2131,N_1314,N_779);
and U2132 (N_2132,N_779,N_1158);
or U2133 (N_2133,N_929,N_1271);
nand U2134 (N_2134,N_1188,N_1435);
nor U2135 (N_2135,N_875,N_867);
or U2136 (N_2136,N_1187,N_1177);
or U2137 (N_2137,N_906,N_1126);
nand U2138 (N_2138,N_846,N_1435);
or U2139 (N_2139,N_1223,N_777);
xor U2140 (N_2140,N_1019,N_938);
nand U2141 (N_2141,N_1324,N_779);
nor U2142 (N_2142,N_1126,N_822);
or U2143 (N_2143,N_1143,N_1037);
nor U2144 (N_2144,N_1322,N_1497);
and U2145 (N_2145,N_1481,N_1348);
nor U2146 (N_2146,N_1320,N_1316);
nand U2147 (N_2147,N_1443,N_1257);
nor U2148 (N_2148,N_1029,N_1467);
and U2149 (N_2149,N_1209,N_1280);
nand U2150 (N_2150,N_787,N_1227);
or U2151 (N_2151,N_904,N_1046);
nand U2152 (N_2152,N_1382,N_1307);
or U2153 (N_2153,N_1103,N_1298);
or U2154 (N_2154,N_1023,N_972);
or U2155 (N_2155,N_1180,N_1172);
nor U2156 (N_2156,N_932,N_1228);
nor U2157 (N_2157,N_1167,N_1448);
nand U2158 (N_2158,N_1250,N_1346);
nand U2159 (N_2159,N_1325,N_1066);
nor U2160 (N_2160,N_1155,N_784);
and U2161 (N_2161,N_956,N_966);
or U2162 (N_2162,N_1460,N_1431);
nand U2163 (N_2163,N_1038,N_806);
xor U2164 (N_2164,N_1373,N_1092);
nor U2165 (N_2165,N_818,N_1156);
nand U2166 (N_2166,N_1231,N_1439);
nor U2167 (N_2167,N_1078,N_896);
nor U2168 (N_2168,N_1395,N_1442);
nor U2169 (N_2169,N_1210,N_948);
or U2170 (N_2170,N_901,N_1357);
and U2171 (N_2171,N_1031,N_1474);
and U2172 (N_2172,N_1471,N_1032);
nor U2173 (N_2173,N_1255,N_1178);
nand U2174 (N_2174,N_756,N_1488);
and U2175 (N_2175,N_1087,N_1047);
nor U2176 (N_2176,N_869,N_1205);
and U2177 (N_2177,N_1475,N_829);
nor U2178 (N_2178,N_858,N_1428);
or U2179 (N_2179,N_804,N_1046);
and U2180 (N_2180,N_1414,N_936);
xnor U2181 (N_2181,N_1448,N_1370);
nand U2182 (N_2182,N_1295,N_1139);
or U2183 (N_2183,N_1242,N_941);
and U2184 (N_2184,N_1223,N_1190);
nand U2185 (N_2185,N_1138,N_1289);
xor U2186 (N_2186,N_1388,N_1163);
or U2187 (N_2187,N_1066,N_848);
nand U2188 (N_2188,N_1062,N_1197);
nor U2189 (N_2189,N_1046,N_802);
nor U2190 (N_2190,N_1194,N_1264);
and U2191 (N_2191,N_1391,N_1354);
and U2192 (N_2192,N_934,N_816);
or U2193 (N_2193,N_923,N_1113);
or U2194 (N_2194,N_1017,N_1131);
nand U2195 (N_2195,N_1047,N_1330);
nor U2196 (N_2196,N_982,N_903);
and U2197 (N_2197,N_1124,N_893);
or U2198 (N_2198,N_1117,N_894);
and U2199 (N_2199,N_1075,N_1461);
nor U2200 (N_2200,N_854,N_1363);
nand U2201 (N_2201,N_893,N_946);
and U2202 (N_2202,N_1087,N_1060);
and U2203 (N_2203,N_947,N_788);
or U2204 (N_2204,N_945,N_1113);
nor U2205 (N_2205,N_1427,N_1409);
or U2206 (N_2206,N_1431,N_1358);
nor U2207 (N_2207,N_855,N_1160);
nand U2208 (N_2208,N_928,N_1145);
nand U2209 (N_2209,N_1389,N_1211);
nand U2210 (N_2210,N_916,N_1229);
nor U2211 (N_2211,N_768,N_1238);
xor U2212 (N_2212,N_842,N_1415);
and U2213 (N_2213,N_1453,N_931);
or U2214 (N_2214,N_826,N_1124);
xor U2215 (N_2215,N_918,N_1264);
and U2216 (N_2216,N_1021,N_874);
nor U2217 (N_2217,N_1156,N_1031);
or U2218 (N_2218,N_1047,N_1052);
nand U2219 (N_2219,N_928,N_766);
and U2220 (N_2220,N_1394,N_1422);
or U2221 (N_2221,N_1012,N_1324);
and U2222 (N_2222,N_976,N_1330);
nor U2223 (N_2223,N_1152,N_1102);
or U2224 (N_2224,N_1276,N_1419);
nor U2225 (N_2225,N_1133,N_810);
nor U2226 (N_2226,N_1352,N_1191);
and U2227 (N_2227,N_893,N_982);
or U2228 (N_2228,N_932,N_1285);
nor U2229 (N_2229,N_1135,N_1343);
or U2230 (N_2230,N_1281,N_1394);
nand U2231 (N_2231,N_804,N_1356);
nor U2232 (N_2232,N_1032,N_1444);
or U2233 (N_2233,N_875,N_849);
nand U2234 (N_2234,N_829,N_1087);
nor U2235 (N_2235,N_1106,N_779);
and U2236 (N_2236,N_1158,N_1403);
nor U2237 (N_2237,N_754,N_1106);
or U2238 (N_2238,N_1013,N_828);
or U2239 (N_2239,N_882,N_927);
and U2240 (N_2240,N_1445,N_803);
or U2241 (N_2241,N_1175,N_1105);
and U2242 (N_2242,N_1450,N_884);
nand U2243 (N_2243,N_841,N_1142);
nand U2244 (N_2244,N_1137,N_933);
and U2245 (N_2245,N_1179,N_1046);
xnor U2246 (N_2246,N_1362,N_1274);
nand U2247 (N_2247,N_1417,N_1290);
and U2248 (N_2248,N_1296,N_778);
and U2249 (N_2249,N_1439,N_1044);
nand U2250 (N_2250,N_2101,N_1535);
or U2251 (N_2251,N_1997,N_1959);
xnor U2252 (N_2252,N_1669,N_1576);
nand U2253 (N_2253,N_1981,N_1696);
nand U2254 (N_2254,N_1604,N_1904);
or U2255 (N_2255,N_1601,N_2161);
nand U2256 (N_2256,N_2205,N_2151);
or U2257 (N_2257,N_1549,N_1731);
or U2258 (N_2258,N_1763,N_1870);
nand U2259 (N_2259,N_1898,N_1721);
nor U2260 (N_2260,N_2087,N_1500);
and U2261 (N_2261,N_1820,N_1761);
nand U2262 (N_2262,N_1903,N_1891);
nand U2263 (N_2263,N_2040,N_2050);
nand U2264 (N_2264,N_1631,N_2170);
or U2265 (N_2265,N_2222,N_1725);
nand U2266 (N_2266,N_1936,N_1862);
nor U2267 (N_2267,N_1680,N_1988);
nor U2268 (N_2268,N_1619,N_1778);
nand U2269 (N_2269,N_1732,N_1503);
nor U2270 (N_2270,N_1706,N_1611);
nand U2271 (N_2271,N_1733,N_1938);
or U2272 (N_2272,N_1691,N_1925);
and U2273 (N_2273,N_2042,N_2013);
or U2274 (N_2274,N_1743,N_2107);
and U2275 (N_2275,N_1530,N_1976);
and U2276 (N_2276,N_2143,N_1547);
or U2277 (N_2277,N_2194,N_1784);
and U2278 (N_2278,N_1849,N_1569);
and U2279 (N_2279,N_1753,N_1768);
or U2280 (N_2280,N_1799,N_2160);
nand U2281 (N_2281,N_1990,N_1756);
and U2282 (N_2282,N_1739,N_2103);
or U2283 (N_2283,N_1823,N_1970);
nor U2284 (N_2284,N_1765,N_2247);
nand U2285 (N_2285,N_2022,N_2196);
and U2286 (N_2286,N_2169,N_1962);
nor U2287 (N_2287,N_1865,N_2185);
or U2288 (N_2288,N_2071,N_2159);
nor U2289 (N_2289,N_1996,N_1740);
nand U2290 (N_2290,N_1634,N_1512);
and U2291 (N_2291,N_1840,N_2031);
nor U2292 (N_2292,N_1558,N_1557);
or U2293 (N_2293,N_2081,N_1617);
nor U2294 (N_2294,N_2093,N_1502);
nand U2295 (N_2295,N_2051,N_1718);
nor U2296 (N_2296,N_1638,N_2238);
nand U2297 (N_2297,N_1562,N_1827);
or U2298 (N_2298,N_1519,N_2116);
and U2299 (N_2299,N_1808,N_2084);
and U2300 (N_2300,N_1801,N_1987);
nor U2301 (N_2301,N_2211,N_2122);
nand U2302 (N_2302,N_1626,N_2124);
and U2303 (N_2303,N_1847,N_1821);
nor U2304 (N_2304,N_1881,N_2063);
nor U2305 (N_2305,N_1615,N_2055);
or U2306 (N_2306,N_2078,N_1846);
nor U2307 (N_2307,N_2057,N_2006);
nand U2308 (N_2308,N_1693,N_1662);
nor U2309 (N_2309,N_1672,N_1501);
and U2310 (N_2310,N_1586,N_2008);
or U2311 (N_2311,N_1689,N_2121);
or U2312 (N_2312,N_2241,N_1596);
nand U2313 (N_2313,N_2167,N_1864);
nand U2314 (N_2314,N_2073,N_1647);
nor U2315 (N_2315,N_1878,N_1629);
and U2316 (N_2316,N_1888,N_1606);
or U2317 (N_2317,N_2060,N_1979);
nor U2318 (N_2318,N_1782,N_1687);
nor U2319 (N_2319,N_2033,N_1661);
and U2320 (N_2320,N_1949,N_2190);
and U2321 (N_2321,N_1532,N_1614);
nand U2322 (N_2322,N_2157,N_1873);
and U2323 (N_2323,N_1723,N_1651);
nor U2324 (N_2324,N_2045,N_2164);
nand U2325 (N_2325,N_1975,N_1991);
nor U2326 (N_2326,N_1663,N_2133);
or U2327 (N_2327,N_1704,N_1828);
nand U2328 (N_2328,N_1800,N_1710);
and U2329 (N_2329,N_1831,N_1525);
nor U2330 (N_2330,N_2027,N_1678);
xnor U2331 (N_2331,N_2016,N_1514);
nand U2332 (N_2332,N_1599,N_1946);
or U2333 (N_2333,N_1931,N_1565);
or U2334 (N_2334,N_1955,N_2220);
or U2335 (N_2335,N_1914,N_1553);
nor U2336 (N_2336,N_1934,N_1509);
and U2337 (N_2337,N_2110,N_1977);
and U2338 (N_2338,N_2023,N_1790);
and U2339 (N_2339,N_1958,N_1793);
and U2340 (N_2340,N_1655,N_1924);
or U2341 (N_2341,N_1961,N_1792);
nor U2342 (N_2342,N_1589,N_2011);
nor U2343 (N_2343,N_2208,N_2155);
or U2344 (N_2344,N_1795,N_2004);
nor U2345 (N_2345,N_2195,N_1625);
or U2346 (N_2346,N_2009,N_1602);
nand U2347 (N_2347,N_1843,N_1892);
nand U2348 (N_2348,N_2127,N_2059);
xnor U2349 (N_2349,N_1741,N_2002);
nor U2350 (N_2350,N_1600,N_2158);
nand U2351 (N_2351,N_1728,N_1912);
and U2352 (N_2352,N_1755,N_2210);
or U2353 (N_2353,N_2131,N_1513);
nor U2354 (N_2354,N_1620,N_1966);
nor U2355 (N_2355,N_2092,N_2123);
nand U2356 (N_2356,N_2219,N_1818);
nand U2357 (N_2357,N_1886,N_2153);
nor U2358 (N_2358,N_2005,N_1715);
xor U2359 (N_2359,N_1835,N_2145);
nor U2360 (N_2360,N_2213,N_2174);
or U2361 (N_2361,N_2139,N_1572);
nor U2362 (N_2362,N_1695,N_2245);
and U2363 (N_2363,N_2079,N_1730);
nand U2364 (N_2364,N_1563,N_2216);
or U2365 (N_2365,N_2089,N_2019);
and U2366 (N_2366,N_1571,N_2049);
nor U2367 (N_2367,N_2191,N_1758);
nand U2368 (N_2368,N_1650,N_2147);
or U2369 (N_2369,N_1694,N_2198);
or U2370 (N_2370,N_2162,N_2119);
nor U2371 (N_2371,N_2214,N_1842);
or U2372 (N_2372,N_1720,N_1552);
and U2373 (N_2373,N_1568,N_1561);
nor U2374 (N_2374,N_1692,N_1508);
nand U2375 (N_2375,N_2086,N_2020);
nor U2376 (N_2376,N_1964,N_2248);
and U2377 (N_2377,N_2118,N_2041);
nor U2378 (N_2378,N_1608,N_1637);
nor U2379 (N_2379,N_1890,N_1524);
and U2380 (N_2380,N_2066,N_1957);
and U2381 (N_2381,N_1587,N_2172);
nor U2382 (N_2382,N_1909,N_1633);
nor U2383 (N_2383,N_2077,N_2070);
and U2384 (N_2384,N_2212,N_1829);
nand U2385 (N_2385,N_2244,N_1861);
nor U2386 (N_2386,N_1699,N_1989);
or U2387 (N_2387,N_1935,N_1839);
nand U2388 (N_2388,N_1775,N_2035);
nand U2389 (N_2389,N_1697,N_1592);
or U2390 (N_2390,N_2193,N_2156);
nand U2391 (N_2391,N_1985,N_1983);
and U2392 (N_2392,N_1984,N_2171);
nor U2393 (N_2393,N_1883,N_1844);
or U2394 (N_2394,N_1830,N_1866);
and U2395 (N_2395,N_1684,N_1666);
or U2396 (N_2396,N_1762,N_2154);
nor U2397 (N_2397,N_2228,N_1591);
and U2398 (N_2398,N_1777,N_2173);
or U2399 (N_2399,N_1559,N_2148);
nand U2400 (N_2400,N_1548,N_2025);
nor U2401 (N_2401,N_2186,N_2236);
and U2402 (N_2402,N_1875,N_2100);
nand U2403 (N_2403,N_2017,N_1664);
nor U2404 (N_2404,N_1887,N_2014);
nor U2405 (N_2405,N_2012,N_1927);
nor U2406 (N_2406,N_1911,N_1856);
and U2407 (N_2407,N_1670,N_1560);
and U2408 (N_2408,N_2115,N_1556);
or U2409 (N_2409,N_1877,N_1813);
nand U2410 (N_2410,N_2065,N_1879);
or U2411 (N_2411,N_1885,N_1564);
nor U2412 (N_2412,N_2053,N_2090);
xnor U2413 (N_2413,N_2234,N_2015);
nor U2414 (N_2414,N_1716,N_1566);
nand U2415 (N_2415,N_1677,N_1915);
nand U2416 (N_2416,N_1635,N_1658);
nand U2417 (N_2417,N_1744,N_1896);
nor U2418 (N_2418,N_1965,N_1956);
and U2419 (N_2419,N_2140,N_1567);
nor U2420 (N_2420,N_1579,N_1627);
nor U2421 (N_2421,N_2074,N_1807);
nor U2422 (N_2422,N_1855,N_1766);
and U2423 (N_2423,N_1834,N_1838);
and U2424 (N_2424,N_2163,N_1610);
nand U2425 (N_2425,N_2226,N_2237);
or U2426 (N_2426,N_2243,N_1948);
nand U2427 (N_2427,N_1544,N_2111);
nand U2428 (N_2428,N_1906,N_1688);
nand U2429 (N_2429,N_2180,N_2109);
nand U2430 (N_2430,N_1652,N_2037);
and U2431 (N_2431,N_1641,N_2128);
nand U2432 (N_2432,N_1644,N_1708);
nor U2433 (N_2433,N_2126,N_2030);
and U2434 (N_2434,N_1752,N_1700);
nand U2435 (N_2435,N_1971,N_1803);
nand U2436 (N_2436,N_2141,N_1690);
nand U2437 (N_2437,N_2150,N_2200);
or U2438 (N_2438,N_1986,N_2221);
nor U2439 (N_2439,N_1901,N_1825);
and U2440 (N_2440,N_2189,N_1645);
nand U2441 (N_2441,N_2104,N_1918);
or U2442 (N_2442,N_1998,N_1642);
or U2443 (N_2443,N_1817,N_1590);
nor U2444 (N_2444,N_1701,N_1806);
nand U2445 (N_2445,N_1794,N_1654);
nand U2446 (N_2446,N_1570,N_1908);
nor U2447 (N_2447,N_2204,N_2038);
and U2448 (N_2448,N_1506,N_2209);
and U2449 (N_2449,N_1769,N_2099);
and U2450 (N_2450,N_1812,N_1802);
or U2451 (N_2451,N_1791,N_1523);
xnor U2452 (N_2452,N_1832,N_1526);
nor U2453 (N_2453,N_1616,N_1969);
and U2454 (N_2454,N_2114,N_1554);
or U2455 (N_2455,N_1555,N_2007);
nand U2456 (N_2456,N_1518,N_1967);
nand U2457 (N_2457,N_1538,N_1707);
nor U2458 (N_2458,N_1796,N_2018);
and U2459 (N_2459,N_1999,N_1528);
nand U2460 (N_2460,N_1505,N_2149);
nand U2461 (N_2461,N_1593,N_1711);
nand U2462 (N_2462,N_1895,N_1869);
and U2463 (N_2463,N_2215,N_2029);
and U2464 (N_2464,N_2058,N_2240);
or U2465 (N_2465,N_1729,N_2064);
and U2466 (N_2466,N_2021,N_1673);
or U2467 (N_2467,N_1923,N_1994);
or U2468 (N_2468,N_1871,N_1907);
or U2469 (N_2469,N_2024,N_1876);
or U2470 (N_2470,N_1722,N_2094);
nor U2471 (N_2471,N_1679,N_1863);
nand U2472 (N_2472,N_2003,N_1880);
and U2473 (N_2473,N_2091,N_1852);
xor U2474 (N_2474,N_2225,N_1698);
or U2475 (N_2475,N_1899,N_1954);
nor U2476 (N_2476,N_1780,N_1712);
and U2477 (N_2477,N_2113,N_1841);
and U2478 (N_2478,N_1609,N_2054);
and U2479 (N_2479,N_1632,N_1760);
or U2480 (N_2480,N_1546,N_1787);
nor U2481 (N_2481,N_1724,N_1926);
and U2482 (N_2482,N_1582,N_1960);
and U2483 (N_2483,N_1939,N_1575);
and U2484 (N_2484,N_1776,N_1685);
nor U2485 (N_2485,N_1816,N_1797);
xor U2486 (N_2486,N_2235,N_1759);
nor U2487 (N_2487,N_1972,N_1771);
nand U2488 (N_2488,N_1941,N_1848);
nor U2489 (N_2489,N_1742,N_2181);
nor U2490 (N_2490,N_2207,N_2152);
nand U2491 (N_2491,N_2043,N_1646);
nand U2492 (N_2492,N_2052,N_1750);
nand U2493 (N_2493,N_1919,N_1814);
nor U2494 (N_2494,N_2138,N_1653);
nand U2495 (N_2495,N_2095,N_2230);
and U2496 (N_2496,N_2082,N_1618);
and U2497 (N_2497,N_1713,N_2075);
and U2498 (N_2498,N_1902,N_1580);
or U2499 (N_2499,N_2223,N_1588);
and U2500 (N_2500,N_2056,N_1913);
nand U2501 (N_2501,N_2108,N_2176);
nand U2502 (N_2502,N_2217,N_1534);
or U2503 (N_2503,N_1836,N_1943);
and U2504 (N_2504,N_1850,N_1703);
and U2505 (N_2505,N_1992,N_1515);
or U2506 (N_2506,N_1815,N_2129);
nand U2507 (N_2507,N_1674,N_1630);
nor U2508 (N_2508,N_2085,N_1920);
nor U2509 (N_2509,N_2047,N_1751);
and U2510 (N_2510,N_1545,N_1540);
and U2511 (N_2511,N_1953,N_2125);
and U2512 (N_2512,N_2231,N_1621);
nor U2513 (N_2513,N_1809,N_2246);
nand U2514 (N_2514,N_1573,N_1860);
nand U2515 (N_2515,N_1681,N_1810);
nand U2516 (N_2516,N_2130,N_1734);
and U2517 (N_2517,N_1507,N_2242);
and U2518 (N_2518,N_1717,N_1665);
nor U2519 (N_2519,N_1636,N_1749);
nand U2520 (N_2520,N_1910,N_2097);
nor U2521 (N_2521,N_1702,N_1735);
or U2522 (N_2522,N_2000,N_1772);
and U2523 (N_2523,N_1811,N_1932);
or U2524 (N_2524,N_1851,N_1668);
nand U2525 (N_2525,N_2080,N_1682);
nand U2526 (N_2526,N_2096,N_2135);
or U2527 (N_2527,N_1671,N_1624);
nor U2528 (N_2528,N_2178,N_1510);
and U2529 (N_2529,N_2046,N_1940);
and U2530 (N_2530,N_1623,N_1822);
nor U2531 (N_2531,N_1785,N_1622);
or U2532 (N_2532,N_1950,N_2187);
and U2533 (N_2533,N_1612,N_2203);
xor U2534 (N_2534,N_1947,N_1736);
and U2535 (N_2535,N_1952,N_1853);
nor U2536 (N_2536,N_2137,N_1516);
nand U2537 (N_2537,N_1779,N_1585);
nand U2538 (N_2538,N_2083,N_1656);
nand U2539 (N_2539,N_1660,N_2183);
and U2540 (N_2540,N_1854,N_2061);
nor U2541 (N_2541,N_2227,N_1824);
nor U2542 (N_2542,N_1933,N_1597);
nand U2543 (N_2543,N_1922,N_1773);
nand U2544 (N_2544,N_2146,N_1584);
nand U2545 (N_2545,N_1714,N_1942);
xnor U2546 (N_2546,N_1826,N_1737);
nand U2547 (N_2547,N_2098,N_1648);
nand U2548 (N_2548,N_2034,N_1894);
or U2549 (N_2549,N_1709,N_1537);
nand U2550 (N_2550,N_1858,N_1639);
nand U2551 (N_2551,N_1905,N_1921);
and U2552 (N_2552,N_1640,N_1819);
or U2553 (N_2553,N_1884,N_2067);
xnor U2554 (N_2554,N_2175,N_1900);
nand U2555 (N_2555,N_1551,N_2218);
nor U2556 (N_2556,N_1521,N_2102);
xor U2557 (N_2557,N_1745,N_2120);
nor U2558 (N_2558,N_1951,N_2069);
nor U2559 (N_2559,N_2179,N_1872);
nor U2560 (N_2560,N_2184,N_1993);
and U2561 (N_2561,N_1789,N_1764);
and U2562 (N_2562,N_1874,N_1542);
nand U2563 (N_2563,N_1963,N_1719);
nor U2564 (N_2564,N_1788,N_1536);
or U2565 (N_2565,N_1837,N_1613);
nor U2566 (N_2566,N_1945,N_2032);
or U2567 (N_2567,N_1605,N_1804);
nor U2568 (N_2568,N_2062,N_2199);
nor U2569 (N_2569,N_1973,N_1726);
nor U2570 (N_2570,N_1930,N_1686);
or U2571 (N_2571,N_1774,N_2026);
or U2572 (N_2572,N_1511,N_2239);
xor U2573 (N_2573,N_2182,N_1767);
nand U2574 (N_2574,N_1867,N_1916);
and U2575 (N_2575,N_1781,N_1643);
or U2576 (N_2576,N_1603,N_2166);
xnor U2577 (N_2577,N_2142,N_2168);
nor U2578 (N_2578,N_1882,N_2202);
nand U2579 (N_2579,N_1757,N_2001);
or U2580 (N_2580,N_1995,N_1676);
nand U2581 (N_2581,N_1531,N_1980);
and U2582 (N_2582,N_1857,N_2132);
nand U2583 (N_2583,N_2249,N_1628);
and U2584 (N_2584,N_2224,N_1595);
or U2585 (N_2585,N_1859,N_1578);
nand U2586 (N_2586,N_2105,N_1937);
nand U2587 (N_2587,N_1978,N_1770);
nand U2588 (N_2588,N_1929,N_1868);
or U2589 (N_2589,N_1527,N_1517);
or U2590 (N_2590,N_1727,N_1607);
nand U2591 (N_2591,N_1968,N_2165);
or U2592 (N_2592,N_2136,N_2028);
nor U2593 (N_2593,N_1659,N_1543);
or U2594 (N_2594,N_1539,N_1705);
xor U2595 (N_2595,N_1798,N_1583);
nor U2596 (N_2596,N_2039,N_1522);
nand U2597 (N_2597,N_2072,N_2233);
and U2598 (N_2598,N_2088,N_2229);
nand U2599 (N_2599,N_1541,N_2232);
xor U2600 (N_2600,N_2068,N_1805);
and U2601 (N_2601,N_2188,N_1683);
nand U2602 (N_2602,N_1533,N_2192);
or U2603 (N_2603,N_1667,N_2112);
and U2604 (N_2604,N_1657,N_1649);
and U2605 (N_2605,N_2117,N_1889);
nor U2606 (N_2606,N_1581,N_1833);
and U2607 (N_2607,N_2197,N_1928);
nand U2608 (N_2608,N_1574,N_1893);
and U2609 (N_2609,N_1944,N_1754);
nor U2610 (N_2610,N_1550,N_2201);
and U2611 (N_2611,N_2134,N_1783);
and U2612 (N_2612,N_1577,N_1738);
nand U2613 (N_2613,N_1974,N_2206);
and U2614 (N_2614,N_1598,N_1520);
nor U2615 (N_2615,N_1748,N_2106);
nand U2616 (N_2616,N_1529,N_2010);
nand U2617 (N_2617,N_1982,N_2144);
nand U2618 (N_2618,N_1675,N_1504);
or U2619 (N_2619,N_2076,N_2036);
or U2620 (N_2620,N_2048,N_1786);
nor U2621 (N_2621,N_1845,N_1897);
nand U2622 (N_2622,N_1746,N_1917);
nor U2623 (N_2623,N_2044,N_2177);
and U2624 (N_2624,N_1594,N_1747);
nor U2625 (N_2625,N_1590,N_1942);
and U2626 (N_2626,N_1515,N_1781);
nand U2627 (N_2627,N_2072,N_1649);
or U2628 (N_2628,N_1509,N_2063);
nand U2629 (N_2629,N_2110,N_2048);
nor U2630 (N_2630,N_1902,N_1719);
nand U2631 (N_2631,N_1544,N_1711);
nor U2632 (N_2632,N_1625,N_2050);
nor U2633 (N_2633,N_2030,N_1691);
nand U2634 (N_2634,N_1543,N_1883);
nand U2635 (N_2635,N_2078,N_1734);
nor U2636 (N_2636,N_1947,N_2212);
nand U2637 (N_2637,N_2025,N_1695);
or U2638 (N_2638,N_1769,N_2033);
and U2639 (N_2639,N_1803,N_2042);
or U2640 (N_2640,N_1885,N_1589);
nand U2641 (N_2641,N_1704,N_2119);
nor U2642 (N_2642,N_2119,N_1898);
nor U2643 (N_2643,N_2134,N_1950);
or U2644 (N_2644,N_1930,N_1831);
nand U2645 (N_2645,N_1576,N_2141);
nor U2646 (N_2646,N_1876,N_1750);
nor U2647 (N_2647,N_1676,N_2227);
and U2648 (N_2648,N_2099,N_1702);
and U2649 (N_2649,N_1970,N_1620);
nor U2650 (N_2650,N_2249,N_1531);
nand U2651 (N_2651,N_1552,N_1897);
nor U2652 (N_2652,N_2245,N_1713);
and U2653 (N_2653,N_2208,N_1931);
or U2654 (N_2654,N_2223,N_1967);
xor U2655 (N_2655,N_1830,N_2013);
and U2656 (N_2656,N_1782,N_1746);
and U2657 (N_2657,N_1948,N_1624);
or U2658 (N_2658,N_1907,N_2122);
nor U2659 (N_2659,N_1502,N_2235);
nand U2660 (N_2660,N_2130,N_1684);
or U2661 (N_2661,N_1736,N_1782);
nor U2662 (N_2662,N_2219,N_1741);
nand U2663 (N_2663,N_1967,N_2235);
or U2664 (N_2664,N_2067,N_1926);
and U2665 (N_2665,N_1657,N_1620);
and U2666 (N_2666,N_2052,N_1921);
and U2667 (N_2667,N_1974,N_1558);
nor U2668 (N_2668,N_1973,N_1553);
and U2669 (N_2669,N_2235,N_2139);
nand U2670 (N_2670,N_2158,N_1855);
nor U2671 (N_2671,N_1588,N_2217);
and U2672 (N_2672,N_1891,N_1900);
nand U2673 (N_2673,N_1962,N_2073);
nor U2674 (N_2674,N_1578,N_1602);
or U2675 (N_2675,N_1867,N_2069);
nand U2676 (N_2676,N_1594,N_1753);
nor U2677 (N_2677,N_1618,N_1986);
nor U2678 (N_2678,N_1945,N_1818);
and U2679 (N_2679,N_1577,N_1735);
or U2680 (N_2680,N_2127,N_1910);
or U2681 (N_2681,N_1730,N_1609);
nor U2682 (N_2682,N_2018,N_2093);
xnor U2683 (N_2683,N_1931,N_2145);
or U2684 (N_2684,N_1899,N_1840);
nor U2685 (N_2685,N_2106,N_1507);
nand U2686 (N_2686,N_2082,N_1950);
nand U2687 (N_2687,N_2164,N_1802);
nor U2688 (N_2688,N_1849,N_2090);
nor U2689 (N_2689,N_1978,N_2047);
nand U2690 (N_2690,N_1928,N_2048);
nor U2691 (N_2691,N_1762,N_2126);
nand U2692 (N_2692,N_1510,N_1604);
xnor U2693 (N_2693,N_1979,N_1539);
nand U2694 (N_2694,N_1602,N_2020);
nor U2695 (N_2695,N_1710,N_1752);
nor U2696 (N_2696,N_2024,N_1751);
nor U2697 (N_2697,N_1992,N_2044);
nand U2698 (N_2698,N_1673,N_1902);
nand U2699 (N_2699,N_1981,N_1581);
and U2700 (N_2700,N_1806,N_1599);
nor U2701 (N_2701,N_2010,N_1751);
nor U2702 (N_2702,N_1922,N_1714);
nand U2703 (N_2703,N_2174,N_2179);
or U2704 (N_2704,N_1993,N_2075);
and U2705 (N_2705,N_1563,N_1590);
nand U2706 (N_2706,N_2239,N_1639);
or U2707 (N_2707,N_1634,N_1735);
and U2708 (N_2708,N_2003,N_1742);
nor U2709 (N_2709,N_2085,N_1913);
and U2710 (N_2710,N_1667,N_2187);
or U2711 (N_2711,N_1501,N_1854);
nor U2712 (N_2712,N_2085,N_1576);
or U2713 (N_2713,N_1530,N_1947);
or U2714 (N_2714,N_1617,N_2168);
or U2715 (N_2715,N_2145,N_2043);
nand U2716 (N_2716,N_1843,N_2123);
and U2717 (N_2717,N_2033,N_1607);
nand U2718 (N_2718,N_1739,N_1782);
and U2719 (N_2719,N_2160,N_2249);
and U2720 (N_2720,N_1757,N_2089);
nand U2721 (N_2721,N_2216,N_1667);
nand U2722 (N_2722,N_1611,N_1828);
nor U2723 (N_2723,N_2232,N_1950);
and U2724 (N_2724,N_1966,N_1756);
or U2725 (N_2725,N_1890,N_1879);
or U2726 (N_2726,N_2138,N_1522);
and U2727 (N_2727,N_2010,N_1571);
and U2728 (N_2728,N_1596,N_1946);
nand U2729 (N_2729,N_1834,N_1980);
nand U2730 (N_2730,N_1758,N_2064);
or U2731 (N_2731,N_1666,N_2237);
nor U2732 (N_2732,N_1795,N_1965);
or U2733 (N_2733,N_1934,N_2227);
or U2734 (N_2734,N_1533,N_1610);
nand U2735 (N_2735,N_1949,N_2120);
nor U2736 (N_2736,N_1992,N_2210);
and U2737 (N_2737,N_1954,N_2212);
or U2738 (N_2738,N_2103,N_1804);
nor U2739 (N_2739,N_1738,N_2069);
nor U2740 (N_2740,N_1543,N_1665);
and U2741 (N_2741,N_1519,N_1953);
or U2742 (N_2742,N_1757,N_2069);
or U2743 (N_2743,N_1775,N_2243);
nand U2744 (N_2744,N_1884,N_1771);
and U2745 (N_2745,N_2187,N_2156);
nor U2746 (N_2746,N_2158,N_1536);
nor U2747 (N_2747,N_1878,N_1843);
nor U2748 (N_2748,N_1965,N_2189);
nor U2749 (N_2749,N_1873,N_1856);
or U2750 (N_2750,N_1868,N_2180);
or U2751 (N_2751,N_2164,N_1954);
and U2752 (N_2752,N_1517,N_1852);
nor U2753 (N_2753,N_2201,N_1720);
nand U2754 (N_2754,N_1689,N_1830);
or U2755 (N_2755,N_2113,N_1858);
or U2756 (N_2756,N_1593,N_1511);
nand U2757 (N_2757,N_1846,N_1666);
or U2758 (N_2758,N_2046,N_2010);
nand U2759 (N_2759,N_1994,N_1647);
nand U2760 (N_2760,N_1781,N_2061);
nand U2761 (N_2761,N_2187,N_1783);
and U2762 (N_2762,N_1767,N_1900);
xnor U2763 (N_2763,N_1590,N_1764);
and U2764 (N_2764,N_2073,N_1848);
nor U2765 (N_2765,N_1564,N_2225);
or U2766 (N_2766,N_1914,N_1595);
nor U2767 (N_2767,N_2081,N_1840);
nand U2768 (N_2768,N_2159,N_1569);
and U2769 (N_2769,N_2166,N_1612);
and U2770 (N_2770,N_1758,N_1692);
or U2771 (N_2771,N_1956,N_2085);
nand U2772 (N_2772,N_1609,N_2033);
nand U2773 (N_2773,N_2108,N_1708);
nor U2774 (N_2774,N_1880,N_1574);
nor U2775 (N_2775,N_1598,N_2016);
nor U2776 (N_2776,N_1813,N_2049);
or U2777 (N_2777,N_1762,N_1685);
or U2778 (N_2778,N_1750,N_1787);
nor U2779 (N_2779,N_2181,N_1677);
nand U2780 (N_2780,N_1522,N_1555);
nor U2781 (N_2781,N_1999,N_1876);
nand U2782 (N_2782,N_2191,N_1764);
xor U2783 (N_2783,N_1803,N_1942);
and U2784 (N_2784,N_1614,N_1829);
and U2785 (N_2785,N_1894,N_1824);
or U2786 (N_2786,N_1913,N_1662);
or U2787 (N_2787,N_1882,N_2014);
nand U2788 (N_2788,N_1975,N_1812);
nor U2789 (N_2789,N_2150,N_2038);
nor U2790 (N_2790,N_1570,N_1799);
and U2791 (N_2791,N_1880,N_1714);
nor U2792 (N_2792,N_2092,N_1665);
and U2793 (N_2793,N_2108,N_1677);
or U2794 (N_2794,N_2051,N_2151);
or U2795 (N_2795,N_1676,N_2176);
or U2796 (N_2796,N_2120,N_1991);
or U2797 (N_2797,N_1630,N_2112);
nand U2798 (N_2798,N_1597,N_1707);
nor U2799 (N_2799,N_2015,N_1771);
nor U2800 (N_2800,N_2220,N_1514);
and U2801 (N_2801,N_1853,N_1524);
and U2802 (N_2802,N_1862,N_2054);
nor U2803 (N_2803,N_1884,N_2181);
nand U2804 (N_2804,N_1654,N_1865);
and U2805 (N_2805,N_2221,N_1705);
nor U2806 (N_2806,N_1673,N_1620);
xor U2807 (N_2807,N_1972,N_1823);
xor U2808 (N_2808,N_2171,N_1834);
and U2809 (N_2809,N_1850,N_1848);
nor U2810 (N_2810,N_1573,N_1852);
or U2811 (N_2811,N_1553,N_2042);
and U2812 (N_2812,N_1710,N_1965);
and U2813 (N_2813,N_1553,N_1600);
or U2814 (N_2814,N_2101,N_2065);
and U2815 (N_2815,N_1778,N_1597);
nor U2816 (N_2816,N_1509,N_2135);
nor U2817 (N_2817,N_1765,N_1625);
nor U2818 (N_2818,N_1599,N_1778);
and U2819 (N_2819,N_1692,N_1984);
and U2820 (N_2820,N_1915,N_1663);
xor U2821 (N_2821,N_1614,N_1563);
nand U2822 (N_2822,N_2070,N_1695);
nand U2823 (N_2823,N_1707,N_1983);
nor U2824 (N_2824,N_1951,N_1937);
nor U2825 (N_2825,N_2000,N_2105);
nor U2826 (N_2826,N_1512,N_1763);
nor U2827 (N_2827,N_1641,N_2227);
nor U2828 (N_2828,N_1638,N_2058);
nand U2829 (N_2829,N_1755,N_1621);
or U2830 (N_2830,N_2070,N_1940);
and U2831 (N_2831,N_2099,N_1759);
or U2832 (N_2832,N_1560,N_1686);
nand U2833 (N_2833,N_2225,N_2145);
or U2834 (N_2834,N_1548,N_2248);
and U2835 (N_2835,N_1669,N_2123);
and U2836 (N_2836,N_2190,N_1584);
nor U2837 (N_2837,N_1765,N_1694);
and U2838 (N_2838,N_2105,N_1922);
and U2839 (N_2839,N_1988,N_1736);
nor U2840 (N_2840,N_2069,N_1621);
nand U2841 (N_2841,N_1712,N_1830);
nor U2842 (N_2842,N_1663,N_1875);
nand U2843 (N_2843,N_1800,N_1569);
nor U2844 (N_2844,N_1509,N_2069);
nand U2845 (N_2845,N_1906,N_2195);
xor U2846 (N_2846,N_2094,N_1949);
or U2847 (N_2847,N_1822,N_1849);
nor U2848 (N_2848,N_2083,N_1743);
or U2849 (N_2849,N_1684,N_1890);
nor U2850 (N_2850,N_2207,N_1510);
or U2851 (N_2851,N_1891,N_2018);
and U2852 (N_2852,N_1992,N_2081);
and U2853 (N_2853,N_1632,N_2156);
nand U2854 (N_2854,N_2247,N_1629);
nor U2855 (N_2855,N_1938,N_1926);
nand U2856 (N_2856,N_1744,N_1793);
nand U2857 (N_2857,N_1557,N_1795);
and U2858 (N_2858,N_1846,N_1850);
nor U2859 (N_2859,N_1795,N_1976);
and U2860 (N_2860,N_1735,N_2102);
and U2861 (N_2861,N_2137,N_1830);
and U2862 (N_2862,N_1851,N_2027);
nand U2863 (N_2863,N_2088,N_2167);
xnor U2864 (N_2864,N_1513,N_1806);
nand U2865 (N_2865,N_1919,N_1855);
or U2866 (N_2866,N_1803,N_1557);
or U2867 (N_2867,N_2112,N_1877);
or U2868 (N_2868,N_1509,N_1908);
or U2869 (N_2869,N_1876,N_2004);
and U2870 (N_2870,N_1545,N_1561);
nand U2871 (N_2871,N_1508,N_2007);
nand U2872 (N_2872,N_1698,N_1875);
nand U2873 (N_2873,N_1545,N_2055);
nor U2874 (N_2874,N_1903,N_2118);
nor U2875 (N_2875,N_1858,N_1637);
nor U2876 (N_2876,N_1506,N_1632);
or U2877 (N_2877,N_1703,N_1904);
and U2878 (N_2878,N_2010,N_2231);
nand U2879 (N_2879,N_1536,N_2202);
nor U2880 (N_2880,N_1637,N_1800);
or U2881 (N_2881,N_1661,N_1579);
nor U2882 (N_2882,N_1729,N_1582);
nor U2883 (N_2883,N_1508,N_1731);
xnor U2884 (N_2884,N_2081,N_2032);
nor U2885 (N_2885,N_2115,N_1500);
nand U2886 (N_2886,N_1880,N_1836);
nand U2887 (N_2887,N_2230,N_1828);
or U2888 (N_2888,N_2083,N_2071);
nor U2889 (N_2889,N_2039,N_1984);
or U2890 (N_2890,N_1941,N_2195);
and U2891 (N_2891,N_1819,N_1598);
and U2892 (N_2892,N_1745,N_2124);
nand U2893 (N_2893,N_1786,N_1767);
nor U2894 (N_2894,N_2214,N_1699);
or U2895 (N_2895,N_2134,N_1721);
and U2896 (N_2896,N_1592,N_1740);
nand U2897 (N_2897,N_1504,N_1952);
nor U2898 (N_2898,N_1722,N_1879);
and U2899 (N_2899,N_2045,N_1785);
or U2900 (N_2900,N_1892,N_2122);
or U2901 (N_2901,N_1858,N_1565);
or U2902 (N_2902,N_1896,N_1581);
and U2903 (N_2903,N_2153,N_1647);
and U2904 (N_2904,N_2114,N_1916);
or U2905 (N_2905,N_1524,N_1739);
or U2906 (N_2906,N_1559,N_2147);
and U2907 (N_2907,N_1651,N_1510);
nand U2908 (N_2908,N_1821,N_2130);
and U2909 (N_2909,N_1741,N_1532);
and U2910 (N_2910,N_2229,N_1824);
nor U2911 (N_2911,N_1606,N_1784);
nor U2912 (N_2912,N_1933,N_2249);
nand U2913 (N_2913,N_2235,N_1768);
nor U2914 (N_2914,N_1888,N_1573);
nand U2915 (N_2915,N_1548,N_1688);
or U2916 (N_2916,N_1798,N_1823);
and U2917 (N_2917,N_1947,N_1860);
and U2918 (N_2918,N_2075,N_1791);
nand U2919 (N_2919,N_1707,N_2067);
nor U2920 (N_2920,N_1892,N_2009);
nor U2921 (N_2921,N_1731,N_1695);
and U2922 (N_2922,N_1980,N_1529);
xor U2923 (N_2923,N_2150,N_2106);
nand U2924 (N_2924,N_2001,N_2000);
nor U2925 (N_2925,N_1645,N_2027);
and U2926 (N_2926,N_1950,N_2165);
nor U2927 (N_2927,N_1587,N_2149);
nand U2928 (N_2928,N_1665,N_1628);
or U2929 (N_2929,N_1582,N_1878);
or U2930 (N_2930,N_2087,N_1740);
and U2931 (N_2931,N_1710,N_1735);
nor U2932 (N_2932,N_1717,N_1553);
and U2933 (N_2933,N_2131,N_2178);
and U2934 (N_2934,N_2239,N_1716);
or U2935 (N_2935,N_1785,N_2213);
or U2936 (N_2936,N_2125,N_1924);
or U2937 (N_2937,N_1833,N_2099);
or U2938 (N_2938,N_2121,N_2237);
nor U2939 (N_2939,N_1806,N_2027);
or U2940 (N_2940,N_1829,N_1923);
or U2941 (N_2941,N_2145,N_1679);
or U2942 (N_2942,N_1726,N_1975);
nor U2943 (N_2943,N_2067,N_1881);
nand U2944 (N_2944,N_1694,N_1657);
nor U2945 (N_2945,N_2128,N_1659);
or U2946 (N_2946,N_1789,N_2156);
or U2947 (N_2947,N_2045,N_1632);
nand U2948 (N_2948,N_1865,N_1555);
and U2949 (N_2949,N_2139,N_2075);
or U2950 (N_2950,N_1505,N_1825);
nor U2951 (N_2951,N_1854,N_2237);
nand U2952 (N_2952,N_1635,N_1649);
nor U2953 (N_2953,N_2112,N_1532);
nor U2954 (N_2954,N_1750,N_1719);
nand U2955 (N_2955,N_1738,N_1879);
nor U2956 (N_2956,N_1982,N_1766);
nand U2957 (N_2957,N_1832,N_1510);
or U2958 (N_2958,N_2057,N_2088);
or U2959 (N_2959,N_1981,N_1575);
or U2960 (N_2960,N_1638,N_1970);
nor U2961 (N_2961,N_1894,N_2059);
nand U2962 (N_2962,N_2096,N_1597);
and U2963 (N_2963,N_1752,N_1996);
or U2964 (N_2964,N_2224,N_1835);
nor U2965 (N_2965,N_2121,N_1771);
nor U2966 (N_2966,N_1990,N_1804);
nor U2967 (N_2967,N_1969,N_1622);
and U2968 (N_2968,N_2089,N_1799);
nand U2969 (N_2969,N_1850,N_1943);
nand U2970 (N_2970,N_1552,N_2141);
xnor U2971 (N_2971,N_1721,N_1830);
or U2972 (N_2972,N_1926,N_1899);
and U2973 (N_2973,N_1858,N_1544);
xor U2974 (N_2974,N_2235,N_1810);
nand U2975 (N_2975,N_1670,N_2241);
or U2976 (N_2976,N_1947,N_1617);
or U2977 (N_2977,N_2133,N_2114);
and U2978 (N_2978,N_1784,N_1866);
or U2979 (N_2979,N_1694,N_1714);
and U2980 (N_2980,N_1723,N_2133);
nor U2981 (N_2981,N_1774,N_1553);
nand U2982 (N_2982,N_1718,N_1740);
or U2983 (N_2983,N_1632,N_1728);
or U2984 (N_2984,N_2153,N_1968);
nand U2985 (N_2985,N_1869,N_2038);
nor U2986 (N_2986,N_2063,N_2150);
or U2987 (N_2987,N_1601,N_2244);
or U2988 (N_2988,N_1501,N_1518);
and U2989 (N_2989,N_2008,N_2157);
nand U2990 (N_2990,N_1613,N_2233);
nor U2991 (N_2991,N_1956,N_2200);
nand U2992 (N_2992,N_2231,N_1912);
nand U2993 (N_2993,N_2026,N_1720);
and U2994 (N_2994,N_1542,N_1990);
nand U2995 (N_2995,N_1561,N_1728);
and U2996 (N_2996,N_2219,N_2142);
or U2997 (N_2997,N_2051,N_1927);
or U2998 (N_2998,N_2072,N_1572);
and U2999 (N_2999,N_2012,N_1711);
nand UO_0 (O_0,N_2982,N_2770);
or UO_1 (O_1,N_2603,N_2955);
and UO_2 (O_2,N_2963,N_2341);
or UO_3 (O_3,N_2752,N_2609);
or UO_4 (O_4,N_2654,N_2939);
or UO_5 (O_5,N_2507,N_2504);
or UO_6 (O_6,N_2840,N_2488);
nor UO_7 (O_7,N_2505,N_2586);
or UO_8 (O_8,N_2605,N_2427);
and UO_9 (O_9,N_2989,N_2338);
or UO_10 (O_10,N_2816,N_2523);
or UO_11 (O_11,N_2506,N_2792);
and UO_12 (O_12,N_2995,N_2283);
nor UO_13 (O_13,N_2592,N_2635);
nor UO_14 (O_14,N_2743,N_2289);
nand UO_15 (O_15,N_2465,N_2735);
and UO_16 (O_16,N_2621,N_2458);
nand UO_17 (O_17,N_2492,N_2571);
nor UO_18 (O_18,N_2869,N_2539);
nand UO_19 (O_19,N_2565,N_2443);
nor UO_20 (O_20,N_2904,N_2815);
xor UO_21 (O_21,N_2489,N_2469);
and UO_22 (O_22,N_2763,N_2852);
or UO_23 (O_23,N_2751,N_2940);
and UO_24 (O_24,N_2864,N_2513);
nand UO_25 (O_25,N_2994,N_2818);
and UO_26 (O_26,N_2876,N_2351);
and UO_27 (O_27,N_2472,N_2951);
nor UO_28 (O_28,N_2528,N_2857);
or UO_29 (O_29,N_2447,N_2633);
or UO_30 (O_30,N_2516,N_2533);
nor UO_31 (O_31,N_2634,N_2430);
nor UO_32 (O_32,N_2777,N_2629);
or UO_33 (O_33,N_2898,N_2789);
nand UO_34 (O_34,N_2705,N_2267);
nand UO_35 (O_35,N_2658,N_2845);
nor UO_36 (O_36,N_2623,N_2286);
and UO_37 (O_37,N_2525,N_2415);
or UO_38 (O_38,N_2487,N_2464);
nor UO_39 (O_39,N_2992,N_2302);
or UO_40 (O_40,N_2374,N_2457);
nand UO_41 (O_41,N_2713,N_2295);
nor UO_42 (O_42,N_2391,N_2961);
xor UO_43 (O_43,N_2663,N_2952);
or UO_44 (O_44,N_2970,N_2502);
or UO_45 (O_45,N_2759,N_2461);
or UO_46 (O_46,N_2574,N_2440);
and UO_47 (O_47,N_2954,N_2964);
nor UO_48 (O_48,N_2354,N_2870);
and UO_49 (O_49,N_2710,N_2331);
nor UO_50 (O_50,N_2493,N_2846);
and UO_51 (O_51,N_2686,N_2819);
nor UO_52 (O_52,N_2606,N_2591);
and UO_53 (O_53,N_2510,N_2874);
nor UO_54 (O_54,N_2801,N_2608);
nand UO_55 (O_55,N_2316,N_2611);
or UO_56 (O_56,N_2687,N_2875);
nor UO_57 (O_57,N_2991,N_2948);
nor UO_58 (O_58,N_2726,N_2290);
or UO_59 (O_59,N_2426,N_2938);
nor UO_60 (O_60,N_2403,N_2908);
nand UO_61 (O_61,N_2647,N_2556);
or UO_62 (O_62,N_2917,N_2388);
and UO_63 (O_63,N_2828,N_2709);
or UO_64 (O_64,N_2402,N_2424);
nand UO_65 (O_65,N_2337,N_2536);
nor UO_66 (O_66,N_2805,N_2596);
nand UO_67 (O_67,N_2262,N_2776);
and UO_68 (O_68,N_2432,N_2787);
nor UO_69 (O_69,N_2600,N_2930);
or UO_70 (O_70,N_2561,N_2958);
or UO_71 (O_71,N_2442,N_2669);
or UO_72 (O_72,N_2750,N_2682);
nor UO_73 (O_73,N_2274,N_2993);
nand UO_74 (O_74,N_2401,N_2913);
nand UO_75 (O_75,N_2837,N_2292);
and UO_76 (O_76,N_2667,N_2406);
or UO_77 (O_77,N_2478,N_2378);
and UO_78 (O_78,N_2671,N_2614);
or UO_79 (O_79,N_2355,N_2367);
and UO_80 (O_80,N_2903,N_2646);
nor UO_81 (O_81,N_2383,N_2340);
nand UO_82 (O_82,N_2325,N_2741);
or UO_83 (O_83,N_2546,N_2485);
nor UO_84 (O_84,N_2333,N_2888);
nand UO_85 (O_85,N_2632,N_2990);
or UO_86 (O_86,N_2980,N_2307);
nand UO_87 (O_87,N_2740,N_2330);
nand UO_88 (O_88,N_2799,N_2589);
or UO_89 (O_89,N_2254,N_2416);
nor UO_90 (O_90,N_2923,N_2508);
and UO_91 (O_91,N_2534,N_2916);
or UO_92 (O_92,N_2643,N_2620);
and UO_93 (O_93,N_2277,N_2684);
nand UO_94 (O_94,N_2676,N_2257);
and UO_95 (O_95,N_2618,N_2924);
nand UO_96 (O_96,N_2637,N_2454);
or UO_97 (O_97,N_2661,N_2593);
and UO_98 (O_98,N_2664,N_2827);
nand UO_99 (O_99,N_2610,N_2317);
nor UO_100 (O_100,N_2548,N_2907);
and UO_101 (O_101,N_2582,N_2865);
and UO_102 (O_102,N_2419,N_2467);
nand UO_103 (O_103,N_2395,N_2365);
nand UO_104 (O_104,N_2971,N_2882);
and UO_105 (O_105,N_2662,N_2891);
nand UO_106 (O_106,N_2261,N_2694);
nand UO_107 (O_107,N_2681,N_2880);
or UO_108 (O_108,N_2832,N_2371);
or UO_109 (O_109,N_2739,N_2973);
xor UO_110 (O_110,N_2878,N_2619);
nor UO_111 (O_111,N_2791,N_2328);
or UO_112 (O_112,N_2967,N_2968);
and UO_113 (O_113,N_2937,N_2369);
or UO_114 (O_114,N_2657,N_2588);
or UO_115 (O_115,N_2300,N_2518);
nor UO_116 (O_116,N_2280,N_2400);
and UO_117 (O_117,N_2576,N_2358);
and UO_118 (O_118,N_2851,N_2714);
and UO_119 (O_119,N_2324,N_2537);
nor UO_120 (O_120,N_2474,N_2644);
nand UO_121 (O_121,N_2305,N_2639);
nand UO_122 (O_122,N_2883,N_2260);
or UO_123 (O_123,N_2481,N_2833);
or UO_124 (O_124,N_2298,N_2947);
and UO_125 (O_125,N_2725,N_2503);
nand UO_126 (O_126,N_2754,N_2717);
nand UO_127 (O_127,N_2414,N_2384);
or UO_128 (O_128,N_2612,N_2793);
or UO_129 (O_129,N_2407,N_2455);
nor UO_130 (O_130,N_2284,N_2526);
nand UO_131 (O_131,N_2742,N_2381);
or UO_132 (O_132,N_2860,N_2486);
nor UO_133 (O_133,N_2479,N_2699);
nand UO_134 (O_134,N_2519,N_2567);
nor UO_135 (O_135,N_2800,N_2933);
and UO_136 (O_136,N_2602,N_2368);
nand UO_137 (O_137,N_2312,N_2781);
or UO_138 (O_138,N_2696,N_2413);
and UO_139 (O_139,N_2497,N_2547);
nor UO_140 (O_140,N_2420,N_2275);
nand UO_141 (O_141,N_2842,N_2597);
nor UO_142 (O_142,N_2692,N_2718);
nand UO_143 (O_143,N_2988,N_2417);
nor UO_144 (O_144,N_2737,N_2631);
and UO_145 (O_145,N_2303,N_2691);
nand UO_146 (O_146,N_2861,N_2444);
or UO_147 (O_147,N_2890,N_2270);
and UO_148 (O_148,N_2564,N_2640);
and UO_149 (O_149,N_2881,N_2969);
or UO_150 (O_150,N_2674,N_2838);
nor UO_151 (O_151,N_2931,N_2960);
or UO_152 (O_152,N_2987,N_2797);
and UO_153 (O_153,N_2382,N_2445);
nor UO_154 (O_154,N_2934,N_2767);
nand UO_155 (O_155,N_2893,N_2665);
nor UO_156 (O_156,N_2310,N_2728);
or UO_157 (O_157,N_2380,N_2531);
or UO_158 (O_158,N_2912,N_2841);
and UO_159 (O_159,N_2269,N_2577);
nand UO_160 (O_160,N_2884,N_2746);
nand UO_161 (O_161,N_2517,N_2941);
xnor UO_162 (O_162,N_2348,N_2810);
and UO_163 (O_163,N_2701,N_2825);
or UO_164 (O_164,N_2950,N_2282);
or UO_165 (O_165,N_2482,N_2702);
xor UO_166 (O_166,N_2352,N_2688);
or UO_167 (O_167,N_2649,N_2583);
and UO_168 (O_168,N_2595,N_2343);
xor UO_169 (O_169,N_2500,N_2285);
nor UO_170 (O_170,N_2919,N_2788);
or UO_171 (O_171,N_2820,N_2377);
nor UO_172 (O_172,N_2423,N_2693);
and UO_173 (O_173,N_2731,N_2753);
nor UO_174 (O_174,N_2981,N_2509);
or UO_175 (O_175,N_2360,N_2345);
nand UO_176 (O_176,N_2524,N_2834);
nand UO_177 (O_177,N_2765,N_2585);
or UO_178 (O_178,N_2451,N_2768);
or UO_179 (O_179,N_2764,N_2578);
nand UO_180 (O_180,N_2659,N_2920);
nor UO_181 (O_181,N_2638,N_2690);
xor UO_182 (O_182,N_2601,N_2978);
xor UO_183 (O_183,N_2297,N_2703);
nand UO_184 (O_184,N_2342,N_2738);
or UO_185 (O_185,N_2334,N_2326);
and UO_186 (O_186,N_2678,N_2498);
nand UO_187 (O_187,N_2306,N_2977);
and UO_188 (O_188,N_2652,N_2986);
or UO_189 (O_189,N_2673,N_2495);
or UO_190 (O_190,N_2397,N_2813);
or UO_191 (O_191,N_2796,N_2868);
or UO_192 (O_192,N_2555,N_2824);
nor UO_193 (O_193,N_2854,N_2480);
nand UO_194 (O_194,N_2641,N_2715);
or UO_195 (O_195,N_2441,N_2910);
and UO_196 (O_196,N_2779,N_2604);
nor UO_197 (O_197,N_2685,N_2922);
nor UO_198 (O_198,N_2786,N_2594);
nand UO_199 (O_199,N_2812,N_2945);
or UO_200 (O_200,N_2719,N_2272);
and UO_201 (O_201,N_2772,N_2376);
and UO_202 (O_202,N_2821,N_2258);
and UO_203 (O_203,N_2872,N_2587);
xnor UO_204 (O_204,N_2732,N_2449);
or UO_205 (O_205,N_2895,N_2894);
nor UO_206 (O_206,N_2859,N_2918);
and UO_207 (O_207,N_2829,N_2625);
or UO_208 (O_208,N_2642,N_2748);
or UO_209 (O_209,N_2323,N_2672);
nand UO_210 (O_210,N_2871,N_2346);
nor UO_211 (O_211,N_2396,N_2901);
and UO_212 (O_212,N_2545,N_2900);
nor UO_213 (O_213,N_2501,N_2744);
nor UO_214 (O_214,N_2613,N_2550);
and UO_215 (O_215,N_2428,N_2256);
nor UO_216 (O_216,N_2867,N_2944);
or UO_217 (O_217,N_2389,N_2483);
nand UO_218 (O_218,N_2724,N_2873);
or UO_219 (O_219,N_2551,N_2999);
nor UO_220 (O_220,N_2532,N_2911);
and UO_221 (O_221,N_2965,N_2757);
and UO_222 (O_222,N_2538,N_2496);
or UO_223 (O_223,N_2668,N_2327);
nor UO_224 (O_224,N_2301,N_2251);
or UO_225 (O_225,N_2450,N_2373);
or UO_226 (O_226,N_2392,N_2892);
or UO_227 (O_227,N_2855,N_2656);
nor UO_228 (O_228,N_2798,N_2405);
nor UO_229 (O_229,N_2268,N_2733);
and UO_230 (O_230,N_2263,N_2749);
and UO_231 (O_231,N_2804,N_2790);
and UO_232 (O_232,N_2766,N_2926);
nor UO_233 (O_233,N_2802,N_2356);
nand UO_234 (O_234,N_2385,N_2466);
and UO_235 (O_235,N_2535,N_2499);
nand UO_236 (O_236,N_2784,N_2344);
nor UO_237 (O_237,N_2452,N_2409);
and UO_238 (O_238,N_2296,N_2288);
or UO_239 (O_239,N_2708,N_2858);
nand UO_240 (O_240,N_2683,N_2549);
and UO_241 (O_241,N_2729,N_2830);
nand UO_242 (O_242,N_2253,N_2785);
nand UO_243 (O_243,N_2736,N_2885);
and UO_244 (O_244,N_2808,N_2946);
and UO_245 (O_245,N_2250,N_2760);
or UO_246 (O_246,N_2627,N_2886);
and UO_247 (O_247,N_2529,N_2372);
nand UO_248 (O_248,N_2569,N_2972);
nor UO_249 (O_249,N_2817,N_2712);
and UO_250 (O_250,N_2491,N_2771);
and UO_251 (O_251,N_2252,N_2782);
nor UO_252 (O_252,N_2552,N_2366);
or UO_253 (O_253,N_2848,N_2541);
nor UO_254 (O_254,N_2581,N_2942);
and UO_255 (O_255,N_2936,N_2411);
and UO_256 (O_256,N_2957,N_2722);
and UO_257 (O_257,N_2336,N_2320);
nor UO_258 (O_258,N_2679,N_2943);
and UO_259 (O_259,N_2425,N_2278);
nand UO_260 (O_260,N_2666,N_2677);
nand UO_261 (O_261,N_2716,N_2421);
nand UO_262 (O_262,N_2580,N_2573);
or UO_263 (O_263,N_2932,N_2698);
or UO_264 (O_264,N_2675,N_2459);
xnor UO_265 (O_265,N_2935,N_2559);
and UO_266 (O_266,N_2359,N_2522);
and UO_267 (O_267,N_2949,N_2446);
and UO_268 (O_268,N_2953,N_2349);
or UO_269 (O_269,N_2599,N_2543);
nand UO_270 (O_270,N_2778,N_2839);
and UO_271 (O_271,N_2959,N_2921);
or UO_272 (O_272,N_2814,N_2755);
and UO_273 (O_273,N_2616,N_2515);
or UO_274 (O_274,N_2475,N_2689);
nor UO_275 (O_275,N_2615,N_2844);
nand UO_276 (O_276,N_2648,N_2866);
and UO_277 (O_277,N_2266,N_2730);
nor UO_278 (O_278,N_2562,N_2607);
and UO_279 (O_279,N_2379,N_2774);
nor UO_280 (O_280,N_2811,N_2394);
and UO_281 (O_281,N_2847,N_2975);
or UO_282 (O_282,N_2264,N_2463);
nor UO_283 (O_283,N_2470,N_2645);
or UO_284 (O_284,N_2575,N_2807);
and UO_285 (O_285,N_2780,N_2490);
nand UO_286 (O_286,N_2436,N_2512);
and UO_287 (O_287,N_2370,N_2437);
nand UO_288 (O_288,N_2271,N_2795);
or UO_289 (O_289,N_2849,N_2477);
or UO_290 (O_290,N_2695,N_2905);
and UO_291 (O_291,N_2293,N_2471);
nor UO_292 (O_292,N_2311,N_2255);
or UO_293 (O_293,N_2769,N_2889);
or UO_294 (O_294,N_2319,N_2927);
nand UO_295 (O_295,N_2563,N_2393);
and UO_296 (O_296,N_2476,N_2353);
nand UO_297 (O_297,N_2363,N_2626);
or UO_298 (O_298,N_2542,N_2362);
and UO_299 (O_299,N_2704,N_2418);
nor UO_300 (O_300,N_2322,N_2598);
and UO_301 (O_301,N_2364,N_2899);
nand UO_302 (O_302,N_2514,N_2783);
nand UO_303 (O_303,N_2711,N_2747);
nand UO_304 (O_304,N_2456,N_2985);
or UO_305 (O_305,N_2398,N_2462);
nand UO_306 (O_306,N_2265,N_2494);
xor UO_307 (O_307,N_2756,N_2622);
and UO_308 (O_308,N_2318,N_2335);
nand UO_309 (O_309,N_2836,N_2636);
nor UO_310 (O_310,N_2521,N_2439);
and UO_311 (O_311,N_2617,N_2655);
nor UO_312 (O_312,N_2761,N_2339);
nand UO_313 (O_313,N_2387,N_2434);
and UO_314 (O_314,N_2294,N_2758);
and UO_315 (O_315,N_2929,N_2332);
xnor UO_316 (O_316,N_2315,N_2408);
or UO_317 (O_317,N_2721,N_2628);
nor UO_318 (O_318,N_2299,N_2279);
nand UO_319 (O_319,N_2473,N_2734);
or UO_320 (O_320,N_2308,N_2956);
or UO_321 (O_321,N_2511,N_2321);
nor UO_322 (O_322,N_2570,N_2794);
nand UO_323 (O_323,N_2557,N_2979);
nor UO_324 (O_324,N_2877,N_2706);
nand UO_325 (O_325,N_2314,N_2412);
nor UO_326 (O_326,N_2762,N_2544);
nand UO_327 (O_327,N_2996,N_2700);
nor UO_328 (O_328,N_2448,N_2435);
and UO_329 (O_329,N_2727,N_2520);
and UO_330 (O_330,N_2404,N_2826);
or UO_331 (O_331,N_2723,N_2558);
or UO_332 (O_332,N_2773,N_2896);
nor UO_333 (O_333,N_2572,N_2484);
or UO_334 (O_334,N_2745,N_2630);
or UO_335 (O_335,N_2914,N_2579);
and UO_336 (O_336,N_2361,N_2806);
xor UO_337 (O_337,N_2902,N_2273);
and UO_338 (O_338,N_2823,N_2928);
xnor UO_339 (O_339,N_2997,N_2998);
or UO_340 (O_340,N_2803,N_2925);
or UO_341 (O_341,N_2350,N_2976);
nand UO_342 (O_342,N_2707,N_2915);
nor UO_343 (O_343,N_2566,N_2680);
nor UO_344 (O_344,N_2410,N_2863);
or UO_345 (O_345,N_2304,N_2309);
and UO_346 (O_346,N_2879,N_2527);
nand UO_347 (O_347,N_2697,N_2720);
and UO_348 (O_348,N_2453,N_2468);
nand UO_349 (O_349,N_2399,N_2966);
nand UO_350 (O_350,N_2974,N_2438);
or UO_351 (O_351,N_2433,N_2390);
nor UO_352 (O_352,N_2422,N_2897);
and UO_353 (O_353,N_2862,N_2983);
nand UO_354 (O_354,N_2809,N_2431);
or UO_355 (O_355,N_2313,N_2853);
and UO_356 (O_356,N_2670,N_2530);
or UO_357 (O_357,N_2375,N_2560);
xnor UO_358 (O_358,N_2584,N_2835);
or UO_359 (O_359,N_2660,N_2650);
nor UO_360 (O_360,N_2287,N_2906);
or UO_361 (O_361,N_2850,N_2259);
nor UO_362 (O_362,N_2386,N_2540);
and UO_363 (O_363,N_2554,N_2429);
nand UO_364 (O_364,N_2347,N_2887);
and UO_365 (O_365,N_2553,N_2568);
nor UO_366 (O_366,N_2843,N_2357);
and UO_367 (O_367,N_2653,N_2856);
nand UO_368 (O_368,N_2291,N_2984);
nor UO_369 (O_369,N_2775,N_2831);
nor UO_370 (O_370,N_2590,N_2822);
or UO_371 (O_371,N_2651,N_2281);
and UO_372 (O_372,N_2624,N_2460);
nand UO_373 (O_373,N_2909,N_2329);
and UO_374 (O_374,N_2276,N_2962);
nand UO_375 (O_375,N_2287,N_2261);
nor UO_376 (O_376,N_2706,N_2502);
or UO_377 (O_377,N_2266,N_2389);
nor UO_378 (O_378,N_2604,N_2757);
and UO_379 (O_379,N_2844,N_2992);
nand UO_380 (O_380,N_2342,N_2909);
or UO_381 (O_381,N_2990,N_2543);
nand UO_382 (O_382,N_2911,N_2985);
nand UO_383 (O_383,N_2462,N_2297);
and UO_384 (O_384,N_2528,N_2285);
nand UO_385 (O_385,N_2481,N_2351);
nand UO_386 (O_386,N_2271,N_2496);
nor UO_387 (O_387,N_2341,N_2902);
nand UO_388 (O_388,N_2354,N_2641);
nand UO_389 (O_389,N_2786,N_2563);
or UO_390 (O_390,N_2564,N_2444);
nor UO_391 (O_391,N_2393,N_2257);
nand UO_392 (O_392,N_2806,N_2771);
or UO_393 (O_393,N_2381,N_2562);
or UO_394 (O_394,N_2902,N_2424);
and UO_395 (O_395,N_2269,N_2834);
nor UO_396 (O_396,N_2400,N_2299);
and UO_397 (O_397,N_2800,N_2812);
nand UO_398 (O_398,N_2740,N_2358);
nand UO_399 (O_399,N_2489,N_2294);
and UO_400 (O_400,N_2338,N_2784);
or UO_401 (O_401,N_2927,N_2476);
xor UO_402 (O_402,N_2269,N_2786);
and UO_403 (O_403,N_2749,N_2489);
nor UO_404 (O_404,N_2265,N_2576);
nor UO_405 (O_405,N_2710,N_2814);
nor UO_406 (O_406,N_2881,N_2253);
nand UO_407 (O_407,N_2468,N_2636);
nor UO_408 (O_408,N_2289,N_2617);
nor UO_409 (O_409,N_2310,N_2288);
nand UO_410 (O_410,N_2888,N_2877);
xnor UO_411 (O_411,N_2970,N_2921);
nand UO_412 (O_412,N_2620,N_2505);
nor UO_413 (O_413,N_2991,N_2799);
and UO_414 (O_414,N_2512,N_2305);
nor UO_415 (O_415,N_2740,N_2431);
or UO_416 (O_416,N_2374,N_2506);
nand UO_417 (O_417,N_2833,N_2875);
and UO_418 (O_418,N_2697,N_2748);
nand UO_419 (O_419,N_2460,N_2981);
nor UO_420 (O_420,N_2848,N_2349);
nor UO_421 (O_421,N_2480,N_2706);
nand UO_422 (O_422,N_2475,N_2297);
and UO_423 (O_423,N_2877,N_2373);
nor UO_424 (O_424,N_2974,N_2583);
nor UO_425 (O_425,N_2891,N_2387);
nor UO_426 (O_426,N_2359,N_2892);
nand UO_427 (O_427,N_2538,N_2485);
nor UO_428 (O_428,N_2927,N_2864);
nand UO_429 (O_429,N_2763,N_2855);
nor UO_430 (O_430,N_2576,N_2399);
and UO_431 (O_431,N_2827,N_2869);
and UO_432 (O_432,N_2514,N_2292);
nand UO_433 (O_433,N_2967,N_2417);
nand UO_434 (O_434,N_2297,N_2353);
nand UO_435 (O_435,N_2694,N_2838);
nor UO_436 (O_436,N_2661,N_2848);
nand UO_437 (O_437,N_2485,N_2954);
or UO_438 (O_438,N_2378,N_2895);
or UO_439 (O_439,N_2495,N_2651);
and UO_440 (O_440,N_2848,N_2472);
and UO_441 (O_441,N_2648,N_2879);
nand UO_442 (O_442,N_2253,N_2392);
nand UO_443 (O_443,N_2853,N_2927);
or UO_444 (O_444,N_2519,N_2508);
nor UO_445 (O_445,N_2891,N_2695);
and UO_446 (O_446,N_2808,N_2378);
nand UO_447 (O_447,N_2422,N_2898);
or UO_448 (O_448,N_2556,N_2850);
nand UO_449 (O_449,N_2764,N_2503);
and UO_450 (O_450,N_2968,N_2307);
and UO_451 (O_451,N_2698,N_2934);
or UO_452 (O_452,N_2309,N_2810);
nand UO_453 (O_453,N_2854,N_2846);
nand UO_454 (O_454,N_2296,N_2828);
nor UO_455 (O_455,N_2474,N_2894);
xor UO_456 (O_456,N_2762,N_2512);
nor UO_457 (O_457,N_2583,N_2421);
nor UO_458 (O_458,N_2518,N_2498);
nand UO_459 (O_459,N_2520,N_2662);
nor UO_460 (O_460,N_2558,N_2533);
and UO_461 (O_461,N_2586,N_2906);
and UO_462 (O_462,N_2598,N_2359);
nor UO_463 (O_463,N_2512,N_2917);
nor UO_464 (O_464,N_2830,N_2423);
or UO_465 (O_465,N_2655,N_2770);
or UO_466 (O_466,N_2530,N_2416);
nand UO_467 (O_467,N_2568,N_2408);
or UO_468 (O_468,N_2915,N_2686);
nor UO_469 (O_469,N_2860,N_2660);
nor UO_470 (O_470,N_2804,N_2277);
nor UO_471 (O_471,N_2312,N_2795);
nand UO_472 (O_472,N_2563,N_2797);
xor UO_473 (O_473,N_2342,N_2505);
nand UO_474 (O_474,N_2830,N_2782);
nor UO_475 (O_475,N_2696,N_2750);
nor UO_476 (O_476,N_2716,N_2324);
nor UO_477 (O_477,N_2968,N_2806);
nand UO_478 (O_478,N_2861,N_2293);
nand UO_479 (O_479,N_2839,N_2752);
or UO_480 (O_480,N_2410,N_2376);
xor UO_481 (O_481,N_2719,N_2511);
nor UO_482 (O_482,N_2647,N_2918);
or UO_483 (O_483,N_2440,N_2439);
nand UO_484 (O_484,N_2598,N_2580);
nand UO_485 (O_485,N_2832,N_2334);
and UO_486 (O_486,N_2959,N_2936);
nand UO_487 (O_487,N_2679,N_2732);
and UO_488 (O_488,N_2283,N_2498);
or UO_489 (O_489,N_2637,N_2933);
nand UO_490 (O_490,N_2736,N_2797);
nand UO_491 (O_491,N_2267,N_2457);
nor UO_492 (O_492,N_2259,N_2486);
nand UO_493 (O_493,N_2469,N_2617);
or UO_494 (O_494,N_2887,N_2552);
nor UO_495 (O_495,N_2559,N_2751);
or UO_496 (O_496,N_2609,N_2939);
and UO_497 (O_497,N_2653,N_2513);
and UO_498 (O_498,N_2480,N_2297);
nand UO_499 (O_499,N_2597,N_2991);
endmodule