module basic_750_5000_1000_10_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_36,In_522);
and U1 (N_1,In_681,In_596);
or U2 (N_2,In_109,In_157);
and U3 (N_3,In_316,In_641);
nor U4 (N_4,In_319,In_636);
nor U5 (N_5,In_541,In_373);
and U6 (N_6,In_435,In_103);
nand U7 (N_7,In_720,In_533);
nor U8 (N_8,In_63,In_51);
and U9 (N_9,In_348,In_259);
nand U10 (N_10,In_45,In_651);
or U11 (N_11,In_405,In_657);
nand U12 (N_12,In_526,In_660);
or U13 (N_13,In_472,In_217);
and U14 (N_14,In_5,In_444);
or U15 (N_15,In_739,In_179);
and U16 (N_16,In_420,In_666);
or U17 (N_17,In_297,In_135);
nand U18 (N_18,In_79,In_618);
and U19 (N_19,In_177,In_647);
and U20 (N_20,In_126,In_2);
and U21 (N_21,In_637,In_452);
nand U22 (N_22,In_461,In_223);
xnor U23 (N_23,In_449,In_245);
nand U24 (N_24,In_576,In_352);
or U25 (N_25,In_570,In_107);
nand U26 (N_26,In_494,In_735);
nor U27 (N_27,In_184,In_4);
nand U28 (N_28,In_571,In_729);
or U29 (N_29,In_410,In_482);
nor U30 (N_30,In_395,In_221);
or U31 (N_31,In_355,In_476);
xnor U32 (N_32,In_285,In_158);
nor U33 (N_33,In_178,In_23);
and U34 (N_34,In_505,In_699);
nand U35 (N_35,In_68,In_585);
nand U36 (N_36,In_451,In_549);
and U37 (N_37,In_548,In_349);
or U38 (N_38,In_457,In_628);
or U39 (N_39,In_293,In_35);
nand U40 (N_40,In_580,In_170);
or U41 (N_41,In_278,In_668);
xor U42 (N_42,In_281,In_421);
and U43 (N_43,In_474,In_193);
nand U44 (N_44,In_380,In_210);
and U45 (N_45,In_587,In_554);
or U46 (N_46,In_543,In_586);
and U47 (N_47,In_624,In_33);
or U48 (N_48,In_347,In_434);
or U49 (N_49,In_528,In_602);
nor U50 (N_50,In_694,In_363);
or U51 (N_51,In_84,In_140);
and U52 (N_52,In_683,In_26);
nor U53 (N_53,In_325,In_268);
nand U54 (N_54,In_492,In_60);
nor U55 (N_55,In_385,In_558);
nand U56 (N_56,In_414,In_493);
and U57 (N_57,In_569,In_390);
and U58 (N_58,In_161,In_18);
and U59 (N_59,In_194,In_11);
nor U60 (N_60,In_697,In_58);
and U61 (N_61,In_251,In_630);
or U62 (N_62,In_53,In_215);
or U63 (N_63,In_669,In_430);
nand U64 (N_64,In_345,In_656);
or U65 (N_65,In_582,In_273);
or U66 (N_66,In_534,In_253);
or U67 (N_67,In_300,In_160);
nand U68 (N_68,In_340,In_743);
xnor U69 (N_69,In_392,In_25);
nand U70 (N_70,In_200,In_484);
nor U71 (N_71,In_315,In_320);
nor U72 (N_72,In_662,In_118);
xnor U73 (N_73,In_439,In_736);
or U74 (N_74,In_64,In_578);
or U75 (N_75,In_201,In_552);
and U76 (N_76,In_696,In_21);
or U77 (N_77,In_102,In_460);
and U78 (N_78,In_137,In_607);
and U79 (N_79,In_69,In_272);
nor U80 (N_80,In_220,In_232);
or U81 (N_81,In_535,In_145);
nand U82 (N_82,In_588,In_356);
and U83 (N_83,In_593,In_331);
nand U84 (N_84,In_466,In_31);
nor U85 (N_85,In_364,In_263);
and U86 (N_86,In_341,In_547);
or U87 (N_87,In_250,In_719);
nor U88 (N_88,In_61,In_346);
or U89 (N_89,In_305,In_41);
nand U90 (N_90,In_591,In_659);
or U91 (N_91,In_143,In_407);
nand U92 (N_92,In_458,In_121);
and U93 (N_93,In_302,In_727);
nand U94 (N_94,In_610,In_747);
nor U95 (N_95,In_133,In_469);
nor U96 (N_96,In_86,In_181);
nor U97 (N_97,In_446,In_168);
nand U98 (N_98,In_74,In_332);
or U99 (N_99,In_129,In_56);
or U100 (N_100,In_115,In_370);
or U101 (N_101,In_164,In_698);
nor U102 (N_102,In_382,In_709);
or U103 (N_103,In_289,In_116);
nor U104 (N_104,In_83,In_208);
or U105 (N_105,In_677,In_402);
nand U106 (N_106,In_214,In_500);
nor U107 (N_107,In_67,In_545);
or U108 (N_108,In_227,In_626);
or U109 (N_109,In_687,In_519);
or U110 (N_110,In_594,In_165);
and U111 (N_111,In_640,In_287);
and U112 (N_112,In_550,In_692);
nor U113 (N_113,In_447,In_358);
nor U114 (N_114,In_511,In_504);
and U115 (N_115,In_676,In_89);
nor U116 (N_116,In_236,In_240);
or U117 (N_117,In_573,In_324);
nand U118 (N_118,In_520,In_509);
nand U119 (N_119,In_92,In_524);
or U120 (N_120,In_128,In_483);
or U121 (N_121,In_303,In_506);
nand U122 (N_122,In_312,In_49);
nor U123 (N_123,In_599,In_714);
nand U124 (N_124,In_746,In_213);
and U125 (N_125,In_94,In_478);
nor U126 (N_126,In_517,In_703);
and U127 (N_127,In_650,In_243);
nor U128 (N_128,In_646,In_288);
and U129 (N_129,In_112,In_639);
nand U130 (N_130,In_96,In_124);
and U131 (N_131,In_485,In_706);
or U132 (N_132,In_516,In_199);
or U133 (N_133,In_387,In_108);
nand U134 (N_134,In_191,In_368);
nand U135 (N_135,In_396,In_12);
and U136 (N_136,In_713,In_189);
xnor U137 (N_137,In_415,In_555);
nor U138 (N_138,In_633,In_66);
and U139 (N_139,In_411,In_498);
nor U140 (N_140,In_427,In_1);
nor U141 (N_141,In_665,In_50);
and U142 (N_142,In_52,In_322);
nor U143 (N_143,In_514,In_216);
and U144 (N_144,In_538,In_423);
nor U145 (N_145,In_621,In_675);
or U146 (N_146,In_725,In_737);
or U147 (N_147,In_47,In_575);
or U148 (N_148,In_684,In_235);
nand U149 (N_149,In_65,In_441);
nand U150 (N_150,In_156,In_601);
nor U151 (N_151,In_562,In_613);
or U152 (N_152,In_330,In_615);
and U153 (N_153,In_44,In_529);
or U154 (N_154,In_173,In_314);
and U155 (N_155,In_323,In_450);
nand U156 (N_156,In_432,In_691);
nand U157 (N_157,In_30,In_301);
nand U158 (N_158,In_603,In_304);
and U159 (N_159,In_391,In_686);
and U160 (N_160,In_142,In_672);
and U161 (N_161,In_360,In_530);
nor U162 (N_162,In_404,In_748);
or U163 (N_163,In_75,In_667);
and U164 (N_164,In_98,In_611);
or U165 (N_165,In_123,In_371);
nor U166 (N_166,In_635,In_551);
or U167 (N_167,In_682,In_311);
nand U168 (N_168,In_393,In_95);
and U169 (N_169,In_604,In_581);
and U170 (N_170,In_367,In_234);
or U171 (N_171,In_480,In_211);
nor U172 (N_172,In_172,In_704);
nor U173 (N_173,In_564,In_117);
nor U174 (N_174,In_507,In_634);
nand U175 (N_175,In_486,In_379);
and U176 (N_176,In_231,In_206);
nand U177 (N_177,In_166,In_671);
or U178 (N_178,In_261,In_241);
nor U179 (N_179,In_34,In_680);
nor U180 (N_180,In_632,In_260);
nor U181 (N_181,In_623,In_462);
and U182 (N_182,In_544,In_617);
nand U183 (N_183,In_648,In_495);
nand U184 (N_184,In_563,In_336);
nor U185 (N_185,In_744,In_375);
nand U186 (N_186,In_233,In_612);
and U187 (N_187,In_359,In_350);
or U188 (N_188,In_417,In_280);
nand U189 (N_189,In_328,In_521);
nor U190 (N_190,In_14,In_284);
nand U191 (N_191,In_337,In_433);
nand U192 (N_192,In_275,In_489);
nor U193 (N_193,In_605,In_207);
nand U194 (N_194,In_196,In_182);
and U195 (N_195,In_335,In_32);
nor U196 (N_196,In_372,In_119);
nor U197 (N_197,In_282,In_749);
or U198 (N_198,In_690,In_497);
or U199 (N_199,In_475,In_459);
or U200 (N_200,In_503,In_388);
nand U201 (N_201,In_631,In_146);
nand U202 (N_202,In_664,In_515);
or U203 (N_203,In_333,In_219);
nand U204 (N_204,In_180,In_147);
nand U205 (N_205,In_292,In_369);
nand U206 (N_206,In_740,In_127);
or U207 (N_207,In_176,In_153);
nor U208 (N_208,In_3,In_353);
nand U209 (N_209,In_20,In_225);
or U210 (N_210,In_111,In_154);
and U211 (N_211,In_643,In_155);
nor U212 (N_212,In_249,In_386);
or U213 (N_213,In_408,In_440);
nand U214 (N_214,In_203,In_228);
nand U215 (N_215,In_310,In_443);
or U216 (N_216,In_546,In_523);
nand U217 (N_217,In_334,In_57);
and U218 (N_218,In_244,In_274);
and U219 (N_219,In_366,In_579);
or U220 (N_220,In_429,In_508);
nor U221 (N_221,In_357,In_431);
xnor U222 (N_222,In_708,In_139);
or U223 (N_223,In_652,In_726);
nor U224 (N_224,In_299,In_183);
nor U225 (N_225,In_378,In_38);
nand U226 (N_226,In_125,In_717);
nor U227 (N_227,In_572,In_710);
or U228 (N_228,In_695,In_198);
and U229 (N_229,In_342,In_384);
and U230 (N_230,In_295,In_711);
and U231 (N_231,In_583,In_252);
or U232 (N_232,In_269,In_678);
nand U233 (N_233,In_365,In_670);
and U234 (N_234,In_590,In_553);
nor U235 (N_235,In_187,In_374);
nor U236 (N_236,In_383,In_638);
nand U237 (N_237,In_255,In_470);
or U238 (N_238,In_693,In_413);
and U239 (N_239,In_267,In_307);
and U240 (N_240,In_501,In_190);
nor U241 (N_241,In_625,In_700);
and U242 (N_242,In_531,In_454);
nor U243 (N_243,In_130,In_418);
and U244 (N_244,In_8,In_653);
and U245 (N_245,In_39,In_649);
nand U246 (N_246,In_271,In_453);
and U247 (N_247,In_192,In_463);
or U248 (N_248,In_565,In_162);
and U249 (N_249,In_242,In_202);
or U250 (N_250,In_105,In_707);
xnor U251 (N_251,In_724,In_502);
nand U252 (N_252,In_270,In_138);
nand U253 (N_253,In_85,In_560);
or U254 (N_254,In_655,In_151);
nor U255 (N_255,In_209,In_19);
nor U256 (N_256,In_150,In_689);
nor U257 (N_257,In_702,In_291);
and U258 (N_258,In_467,In_81);
or U259 (N_259,In_141,In_398);
nand U260 (N_260,In_256,In_149);
and U261 (N_261,In_425,In_688);
nand U262 (N_262,In_701,In_91);
nand U263 (N_263,In_309,In_163);
nor U264 (N_264,In_473,In_577);
nand U265 (N_265,In_110,In_557);
or U266 (N_266,In_597,In_186);
nand U267 (N_267,In_442,In_169);
or U268 (N_268,In_80,In_204);
or U269 (N_269,In_377,In_229);
nor U270 (N_270,In_481,In_403);
and U271 (N_271,In_589,In_394);
nand U272 (N_272,In_445,In_77);
nor U273 (N_273,In_264,In_600);
nor U274 (N_274,In_479,In_15);
and U275 (N_275,In_721,In_620);
nand U276 (N_276,In_471,In_513);
nand U277 (N_277,In_286,In_663);
nor U278 (N_278,In_16,In_327);
nand U279 (N_279,In_422,In_246);
nand U280 (N_280,In_732,In_661);
nand U281 (N_281,In_400,In_438);
nor U282 (N_282,In_627,In_71);
or U283 (N_283,In_428,In_595);
nor U284 (N_284,In_344,In_424);
nor U285 (N_285,In_37,In_188);
or U286 (N_286,In_131,In_247);
nand U287 (N_287,In_10,In_351);
or U288 (N_288,In_90,In_237);
and U289 (N_289,In_134,In_88);
and U290 (N_290,In_313,In_0);
nor U291 (N_291,In_100,In_113);
or U292 (N_292,In_298,In_70);
and U293 (N_293,In_464,In_195);
nor U294 (N_294,In_510,In_468);
nor U295 (N_295,In_512,In_27);
nand U296 (N_296,In_745,In_362);
nor U297 (N_297,In_629,In_87);
nor U298 (N_298,In_321,In_658);
and U299 (N_299,In_17,In_24);
nand U300 (N_300,In_22,In_722);
nor U301 (N_301,In_226,In_419);
or U302 (N_302,In_222,In_496);
nand U303 (N_303,In_437,In_290);
nor U304 (N_304,In_265,In_448);
and U305 (N_305,In_326,In_416);
and U306 (N_306,In_426,In_487);
nand U307 (N_307,In_401,In_93);
and U308 (N_308,In_584,In_13);
or U309 (N_309,In_120,In_258);
or U310 (N_310,In_55,In_152);
or U311 (N_311,In_532,In_317);
or U312 (N_312,In_306,In_318);
nor U313 (N_313,In_642,In_574);
and U314 (N_314,In_540,In_536);
nor U315 (N_315,In_59,In_716);
or U316 (N_316,In_72,In_525);
nand U317 (N_317,In_712,In_338);
and U318 (N_318,In_224,In_136);
or U319 (N_319,In_568,In_205);
nor U320 (N_320,In_742,In_499);
nor U321 (N_321,In_389,In_619);
nand U322 (N_322,In_114,In_361);
and U323 (N_323,In_456,In_539);
nand U324 (N_324,In_718,In_144);
nand U325 (N_325,In_644,In_248);
or U326 (N_326,In_616,In_238);
nor U327 (N_327,In_43,In_376);
nand U328 (N_328,In_608,In_465);
nand U329 (N_329,In_556,In_354);
and U330 (N_330,In_9,In_609);
nor U331 (N_331,In_673,In_174);
nor U332 (N_332,In_46,In_406);
xnor U333 (N_333,In_339,In_159);
nand U334 (N_334,In_622,In_308);
nor U335 (N_335,In_685,In_7);
or U336 (N_336,In_490,In_542);
nor U337 (N_337,In_132,In_488);
nand U338 (N_338,In_715,In_76);
and U339 (N_339,In_29,In_679);
nand U340 (N_340,In_537,In_399);
and U341 (N_341,In_436,In_294);
and U342 (N_342,In_566,In_705);
or U343 (N_343,In_381,In_296);
nor U344 (N_344,In_477,In_343);
or U345 (N_345,In_42,In_171);
and U346 (N_346,In_527,In_175);
or U347 (N_347,In_674,In_266);
and U348 (N_348,In_97,In_101);
or U349 (N_349,In_276,In_730);
or U350 (N_350,In_409,In_723);
nor U351 (N_351,In_212,In_277);
nor U352 (N_352,In_329,In_598);
nand U353 (N_353,In_122,In_733);
and U354 (N_354,In_731,In_254);
nor U355 (N_355,In_561,In_728);
nand U356 (N_356,In_73,In_412);
or U357 (N_357,In_54,In_257);
and U358 (N_358,In_279,In_62);
and U359 (N_359,In_734,In_28);
or U360 (N_360,In_230,In_78);
or U361 (N_361,In_99,In_106);
and U362 (N_362,In_48,In_455);
xor U363 (N_363,In_645,In_606);
and U364 (N_364,In_397,In_592);
nand U365 (N_365,In_218,In_654);
or U366 (N_366,In_239,In_40);
nand U367 (N_367,In_148,In_185);
or U368 (N_368,In_197,In_518);
or U369 (N_369,In_741,In_738);
or U370 (N_370,In_6,In_104);
or U371 (N_371,In_167,In_283);
nand U372 (N_372,In_262,In_567);
or U373 (N_373,In_614,In_491);
or U374 (N_374,In_559,In_82);
nor U375 (N_375,In_120,In_74);
and U376 (N_376,In_587,In_114);
nor U377 (N_377,In_564,In_14);
and U378 (N_378,In_300,In_151);
nor U379 (N_379,In_739,In_121);
nand U380 (N_380,In_140,In_273);
nor U381 (N_381,In_738,In_250);
nand U382 (N_382,In_57,In_367);
nor U383 (N_383,In_681,In_556);
nor U384 (N_384,In_384,In_691);
and U385 (N_385,In_156,In_92);
and U386 (N_386,In_101,In_410);
nand U387 (N_387,In_565,In_462);
and U388 (N_388,In_395,In_123);
xor U389 (N_389,In_541,In_557);
nor U390 (N_390,In_660,In_718);
or U391 (N_391,In_667,In_406);
nand U392 (N_392,In_523,In_328);
and U393 (N_393,In_408,In_352);
nor U394 (N_394,In_267,In_284);
nand U395 (N_395,In_309,In_274);
nand U396 (N_396,In_133,In_475);
or U397 (N_397,In_26,In_695);
nand U398 (N_398,In_230,In_107);
or U399 (N_399,In_335,In_239);
and U400 (N_400,In_29,In_389);
or U401 (N_401,In_238,In_555);
nand U402 (N_402,In_460,In_624);
nor U403 (N_403,In_485,In_145);
and U404 (N_404,In_560,In_272);
nand U405 (N_405,In_550,In_691);
nand U406 (N_406,In_142,In_548);
and U407 (N_407,In_95,In_6);
or U408 (N_408,In_676,In_35);
nor U409 (N_409,In_611,In_631);
nor U410 (N_410,In_369,In_574);
and U411 (N_411,In_532,In_480);
or U412 (N_412,In_506,In_160);
and U413 (N_413,In_433,In_216);
or U414 (N_414,In_495,In_432);
and U415 (N_415,In_449,In_109);
nand U416 (N_416,In_39,In_5);
nand U417 (N_417,In_95,In_610);
nor U418 (N_418,In_269,In_533);
and U419 (N_419,In_581,In_180);
and U420 (N_420,In_428,In_258);
and U421 (N_421,In_622,In_365);
nand U422 (N_422,In_619,In_410);
or U423 (N_423,In_426,In_231);
and U424 (N_424,In_130,In_557);
and U425 (N_425,In_672,In_301);
nor U426 (N_426,In_214,In_725);
nor U427 (N_427,In_425,In_29);
or U428 (N_428,In_269,In_345);
and U429 (N_429,In_302,In_181);
nand U430 (N_430,In_66,In_536);
or U431 (N_431,In_291,In_33);
or U432 (N_432,In_640,In_358);
nor U433 (N_433,In_193,In_19);
nand U434 (N_434,In_300,In_548);
and U435 (N_435,In_69,In_625);
nor U436 (N_436,In_573,In_199);
and U437 (N_437,In_275,In_534);
and U438 (N_438,In_573,In_323);
or U439 (N_439,In_367,In_55);
or U440 (N_440,In_645,In_578);
and U441 (N_441,In_349,In_88);
nor U442 (N_442,In_732,In_598);
and U443 (N_443,In_682,In_140);
nor U444 (N_444,In_483,In_207);
nor U445 (N_445,In_29,In_320);
nor U446 (N_446,In_670,In_547);
nor U447 (N_447,In_569,In_670);
xnor U448 (N_448,In_114,In_289);
or U449 (N_449,In_189,In_238);
or U450 (N_450,In_210,In_738);
or U451 (N_451,In_439,In_194);
xor U452 (N_452,In_492,In_318);
and U453 (N_453,In_5,In_518);
or U454 (N_454,In_164,In_682);
nor U455 (N_455,In_475,In_310);
nor U456 (N_456,In_308,In_286);
nor U457 (N_457,In_173,In_502);
or U458 (N_458,In_87,In_110);
nand U459 (N_459,In_120,In_297);
nand U460 (N_460,In_604,In_260);
nand U461 (N_461,In_211,In_447);
nor U462 (N_462,In_731,In_314);
and U463 (N_463,In_563,In_510);
nand U464 (N_464,In_395,In_136);
or U465 (N_465,In_290,In_738);
or U466 (N_466,In_31,In_244);
and U467 (N_467,In_351,In_154);
and U468 (N_468,In_722,In_353);
nor U469 (N_469,In_374,In_518);
nor U470 (N_470,In_564,In_472);
and U471 (N_471,In_520,In_358);
nand U472 (N_472,In_714,In_460);
nand U473 (N_473,In_730,In_473);
nand U474 (N_474,In_396,In_554);
or U475 (N_475,In_407,In_563);
nand U476 (N_476,In_165,In_602);
nand U477 (N_477,In_114,In_323);
nor U478 (N_478,In_470,In_460);
nor U479 (N_479,In_155,In_292);
and U480 (N_480,In_234,In_404);
nand U481 (N_481,In_695,In_529);
or U482 (N_482,In_746,In_388);
nor U483 (N_483,In_143,In_697);
or U484 (N_484,In_724,In_608);
or U485 (N_485,In_469,In_253);
or U486 (N_486,In_93,In_720);
nand U487 (N_487,In_416,In_317);
or U488 (N_488,In_622,In_354);
nor U489 (N_489,In_499,In_689);
or U490 (N_490,In_250,In_473);
or U491 (N_491,In_298,In_357);
and U492 (N_492,In_160,In_420);
or U493 (N_493,In_611,In_379);
or U494 (N_494,In_427,In_167);
and U495 (N_495,In_481,In_24);
nand U496 (N_496,In_3,In_80);
or U497 (N_497,In_144,In_681);
and U498 (N_498,In_209,In_242);
xnor U499 (N_499,In_107,In_55);
xor U500 (N_500,N_283,N_177);
nand U501 (N_501,N_434,N_199);
nor U502 (N_502,N_13,N_27);
or U503 (N_503,N_285,N_247);
nand U504 (N_504,N_31,N_408);
nand U505 (N_505,N_427,N_61);
and U506 (N_506,N_221,N_160);
or U507 (N_507,N_87,N_116);
or U508 (N_508,N_43,N_293);
nor U509 (N_509,N_89,N_451);
or U510 (N_510,N_146,N_329);
nor U511 (N_511,N_461,N_278);
nor U512 (N_512,N_447,N_294);
or U513 (N_513,N_345,N_231);
and U514 (N_514,N_20,N_196);
or U515 (N_515,N_53,N_50);
or U516 (N_516,N_430,N_432);
nor U517 (N_517,N_284,N_218);
or U518 (N_518,N_289,N_21);
nor U519 (N_519,N_230,N_173);
nand U520 (N_520,N_378,N_307);
or U521 (N_521,N_471,N_356);
nor U522 (N_522,N_26,N_236);
or U523 (N_523,N_172,N_438);
nand U524 (N_524,N_141,N_426);
and U525 (N_525,N_475,N_321);
or U526 (N_526,N_128,N_277);
nor U527 (N_527,N_286,N_16);
or U528 (N_528,N_342,N_224);
or U529 (N_529,N_275,N_263);
nor U530 (N_530,N_202,N_117);
and U531 (N_531,N_454,N_120);
nand U532 (N_532,N_25,N_291);
nand U533 (N_533,N_373,N_193);
or U534 (N_534,N_166,N_32);
nand U535 (N_535,N_241,N_181);
xnor U536 (N_536,N_17,N_445);
nor U537 (N_537,N_317,N_153);
and U538 (N_538,N_330,N_467);
nand U539 (N_539,N_155,N_338);
and U540 (N_540,N_387,N_499);
nand U541 (N_541,N_94,N_298);
nand U542 (N_542,N_246,N_41);
nand U543 (N_543,N_110,N_431);
and U544 (N_544,N_418,N_44);
and U545 (N_545,N_93,N_389);
xor U546 (N_546,N_287,N_424);
and U547 (N_547,N_425,N_316);
nand U548 (N_548,N_464,N_79);
nand U549 (N_549,N_487,N_92);
nor U550 (N_550,N_481,N_310);
nand U551 (N_551,N_111,N_207);
or U552 (N_552,N_295,N_114);
nand U553 (N_553,N_201,N_56);
nor U554 (N_554,N_337,N_349);
nand U555 (N_555,N_96,N_282);
nand U556 (N_556,N_159,N_30);
nand U557 (N_557,N_194,N_86);
nor U558 (N_558,N_200,N_409);
and U559 (N_559,N_136,N_491);
and U560 (N_560,N_394,N_103);
nor U561 (N_561,N_149,N_419);
nand U562 (N_562,N_211,N_290);
or U563 (N_563,N_353,N_229);
nand U564 (N_564,N_217,N_164);
nor U565 (N_565,N_142,N_182);
nand U566 (N_566,N_122,N_152);
or U567 (N_567,N_492,N_348);
xor U568 (N_568,N_299,N_335);
and U569 (N_569,N_390,N_302);
nand U570 (N_570,N_130,N_102);
and U571 (N_571,N_242,N_145);
nor U572 (N_572,N_137,N_305);
nor U573 (N_573,N_77,N_188);
nor U574 (N_574,N_95,N_465);
and U575 (N_575,N_429,N_386);
nand U576 (N_576,N_380,N_139);
and U577 (N_577,N_273,N_352);
nand U578 (N_578,N_165,N_51);
nor U579 (N_579,N_148,N_197);
nand U580 (N_580,N_466,N_473);
nand U581 (N_581,N_113,N_483);
nand U582 (N_582,N_112,N_456);
and U583 (N_583,N_272,N_163);
or U584 (N_584,N_151,N_187);
or U585 (N_585,N_311,N_253);
nor U586 (N_586,N_174,N_453);
or U587 (N_587,N_192,N_365);
nand U588 (N_588,N_267,N_0);
nand U589 (N_589,N_458,N_281);
or U590 (N_590,N_367,N_479);
or U591 (N_591,N_180,N_393);
nand U592 (N_592,N_4,N_333);
or U593 (N_593,N_439,N_78);
nand U594 (N_594,N_39,N_476);
or U595 (N_595,N_470,N_379);
nand U596 (N_596,N_279,N_7);
nand U597 (N_597,N_171,N_227);
nand U598 (N_598,N_248,N_369);
nand U599 (N_599,N_400,N_140);
or U600 (N_600,N_54,N_340);
and U601 (N_601,N_433,N_167);
and U602 (N_602,N_143,N_260);
nor U603 (N_603,N_416,N_144);
nand U604 (N_604,N_161,N_269);
and U605 (N_605,N_407,N_257);
nand U606 (N_606,N_175,N_449);
and U607 (N_607,N_405,N_119);
or U608 (N_608,N_147,N_63);
and U609 (N_609,N_360,N_64);
nor U610 (N_610,N_15,N_88);
nand U611 (N_611,N_233,N_3);
nand U612 (N_612,N_57,N_325);
and U613 (N_613,N_239,N_462);
or U614 (N_614,N_245,N_437);
nor U615 (N_615,N_14,N_127);
and U616 (N_616,N_420,N_238);
nor U617 (N_617,N_318,N_326);
or U618 (N_618,N_399,N_251);
and U619 (N_619,N_309,N_176);
nor U620 (N_620,N_355,N_489);
nor U621 (N_621,N_10,N_359);
xnor U622 (N_622,N_395,N_480);
nand U623 (N_623,N_252,N_327);
nand U624 (N_624,N_34,N_324);
and U625 (N_625,N_341,N_381);
nor U626 (N_626,N_372,N_108);
or U627 (N_627,N_109,N_169);
nor U628 (N_628,N_19,N_448);
and U629 (N_629,N_126,N_339);
nor U630 (N_630,N_125,N_216);
nand U631 (N_631,N_186,N_457);
or U632 (N_632,N_235,N_361);
nor U633 (N_633,N_121,N_459);
or U634 (N_634,N_132,N_304);
nor U635 (N_635,N_314,N_158);
nor U636 (N_636,N_268,N_226);
and U637 (N_637,N_262,N_370);
or U638 (N_638,N_336,N_375);
or U639 (N_639,N_313,N_244);
or U640 (N_640,N_203,N_351);
nor U641 (N_641,N_477,N_406);
nor U642 (N_642,N_123,N_40);
nor U643 (N_643,N_71,N_206);
nand U644 (N_644,N_168,N_98);
or U645 (N_645,N_357,N_358);
nor U646 (N_646,N_133,N_38);
nand U647 (N_647,N_261,N_495);
or U648 (N_648,N_240,N_300);
nand U649 (N_649,N_37,N_366);
and U650 (N_650,N_412,N_150);
nand U651 (N_651,N_320,N_368);
nand U652 (N_652,N_414,N_255);
and U653 (N_653,N_446,N_450);
and U654 (N_654,N_403,N_65);
nand U655 (N_655,N_234,N_100);
nor U656 (N_656,N_69,N_1);
or U657 (N_657,N_463,N_97);
and U658 (N_658,N_440,N_76);
or U659 (N_659,N_410,N_208);
and U660 (N_660,N_67,N_484);
nor U661 (N_661,N_225,N_296);
nand U662 (N_662,N_343,N_488);
and U663 (N_663,N_129,N_398);
nand U664 (N_664,N_280,N_156);
and U665 (N_665,N_232,N_328);
or U666 (N_666,N_415,N_11);
or U667 (N_667,N_347,N_68);
nand U668 (N_668,N_460,N_5);
and U669 (N_669,N_350,N_250);
and U670 (N_670,N_266,N_179);
nor U671 (N_671,N_22,N_362);
nand U672 (N_672,N_170,N_472);
nand U673 (N_673,N_18,N_292);
and U674 (N_674,N_254,N_388);
or U675 (N_675,N_131,N_383);
and U676 (N_676,N_376,N_198);
and U677 (N_677,N_178,N_308);
and U678 (N_678,N_82,N_402);
or U679 (N_679,N_259,N_223);
or U680 (N_680,N_29,N_212);
and U681 (N_681,N_443,N_482);
xor U682 (N_682,N_490,N_469);
and U683 (N_683,N_452,N_70);
and U684 (N_684,N_478,N_58);
and U685 (N_685,N_72,N_84);
nand U686 (N_686,N_334,N_363);
nor U687 (N_687,N_497,N_104);
nor U688 (N_688,N_9,N_306);
nand U689 (N_689,N_256,N_138);
nand U690 (N_690,N_377,N_391);
or U691 (N_691,N_49,N_190);
nor U692 (N_692,N_297,N_485);
or U693 (N_693,N_28,N_6);
and U694 (N_694,N_24,N_271);
nand U695 (N_695,N_185,N_411);
and U696 (N_696,N_189,N_237);
nor U697 (N_697,N_105,N_134);
nor U698 (N_698,N_220,N_66);
nor U699 (N_699,N_396,N_118);
nand U700 (N_700,N_83,N_213);
and U701 (N_701,N_428,N_344);
nand U702 (N_702,N_493,N_374);
nor U703 (N_703,N_417,N_401);
and U704 (N_704,N_195,N_397);
nand U705 (N_705,N_46,N_115);
nand U706 (N_706,N_332,N_73);
or U707 (N_707,N_59,N_486);
or U708 (N_708,N_91,N_214);
or U709 (N_709,N_364,N_274);
and U710 (N_710,N_288,N_81);
nor U711 (N_711,N_47,N_496);
nor U712 (N_712,N_382,N_184);
nor U713 (N_713,N_312,N_8);
or U714 (N_714,N_441,N_45);
nor U715 (N_715,N_423,N_205);
and U716 (N_716,N_107,N_42);
xnor U717 (N_717,N_209,N_270);
nand U718 (N_718,N_183,N_162);
and U719 (N_719,N_422,N_35);
nand U720 (N_720,N_191,N_468);
nand U721 (N_721,N_258,N_36);
or U722 (N_722,N_99,N_85);
or U723 (N_723,N_62,N_33);
and U724 (N_724,N_55,N_319);
nor U725 (N_725,N_265,N_210);
nand U726 (N_726,N_74,N_384);
nor U727 (N_727,N_301,N_228);
nand U728 (N_728,N_474,N_80);
nand U729 (N_729,N_222,N_276);
or U730 (N_730,N_90,N_264);
nand U731 (N_731,N_494,N_346);
and U732 (N_732,N_135,N_2);
nand U733 (N_733,N_421,N_442);
and U734 (N_734,N_75,N_215);
or U735 (N_735,N_106,N_249);
and U736 (N_736,N_204,N_371);
or U737 (N_737,N_455,N_124);
nor U738 (N_738,N_303,N_498);
and U739 (N_739,N_444,N_243);
and U740 (N_740,N_392,N_436);
nand U741 (N_741,N_12,N_101);
or U742 (N_742,N_354,N_331);
nand U743 (N_743,N_404,N_154);
or U744 (N_744,N_385,N_219);
nor U745 (N_745,N_23,N_322);
or U746 (N_746,N_52,N_435);
and U747 (N_747,N_157,N_60);
nand U748 (N_748,N_413,N_315);
nand U749 (N_749,N_323,N_48);
nand U750 (N_750,N_200,N_4);
or U751 (N_751,N_233,N_421);
and U752 (N_752,N_285,N_40);
or U753 (N_753,N_486,N_334);
nor U754 (N_754,N_458,N_6);
and U755 (N_755,N_361,N_392);
or U756 (N_756,N_33,N_52);
or U757 (N_757,N_316,N_163);
nor U758 (N_758,N_156,N_284);
nor U759 (N_759,N_313,N_129);
and U760 (N_760,N_225,N_83);
nand U761 (N_761,N_438,N_226);
or U762 (N_762,N_160,N_297);
nor U763 (N_763,N_418,N_188);
nor U764 (N_764,N_171,N_48);
nor U765 (N_765,N_465,N_491);
or U766 (N_766,N_47,N_282);
or U767 (N_767,N_203,N_118);
nor U768 (N_768,N_70,N_340);
nor U769 (N_769,N_287,N_11);
or U770 (N_770,N_280,N_457);
nor U771 (N_771,N_268,N_9);
nor U772 (N_772,N_226,N_193);
nor U773 (N_773,N_316,N_52);
or U774 (N_774,N_17,N_431);
nand U775 (N_775,N_419,N_377);
nand U776 (N_776,N_57,N_470);
nor U777 (N_777,N_248,N_401);
nor U778 (N_778,N_157,N_44);
nand U779 (N_779,N_45,N_450);
nor U780 (N_780,N_272,N_45);
nand U781 (N_781,N_175,N_97);
nand U782 (N_782,N_141,N_475);
and U783 (N_783,N_213,N_389);
or U784 (N_784,N_84,N_93);
nor U785 (N_785,N_434,N_454);
or U786 (N_786,N_493,N_385);
nor U787 (N_787,N_479,N_127);
nand U788 (N_788,N_422,N_116);
nor U789 (N_789,N_491,N_191);
and U790 (N_790,N_96,N_459);
or U791 (N_791,N_422,N_211);
and U792 (N_792,N_343,N_16);
nor U793 (N_793,N_250,N_442);
nand U794 (N_794,N_494,N_398);
or U795 (N_795,N_152,N_176);
nor U796 (N_796,N_156,N_315);
or U797 (N_797,N_485,N_190);
nor U798 (N_798,N_484,N_252);
nor U799 (N_799,N_450,N_250);
nor U800 (N_800,N_266,N_84);
and U801 (N_801,N_276,N_383);
and U802 (N_802,N_190,N_69);
and U803 (N_803,N_322,N_273);
nor U804 (N_804,N_408,N_271);
nand U805 (N_805,N_495,N_446);
nand U806 (N_806,N_144,N_433);
nand U807 (N_807,N_254,N_173);
and U808 (N_808,N_122,N_113);
nand U809 (N_809,N_259,N_459);
nor U810 (N_810,N_371,N_462);
or U811 (N_811,N_249,N_346);
nand U812 (N_812,N_217,N_262);
nor U813 (N_813,N_484,N_442);
and U814 (N_814,N_485,N_434);
or U815 (N_815,N_192,N_324);
and U816 (N_816,N_413,N_70);
and U817 (N_817,N_274,N_232);
or U818 (N_818,N_63,N_76);
nor U819 (N_819,N_469,N_259);
and U820 (N_820,N_157,N_398);
nand U821 (N_821,N_283,N_452);
nand U822 (N_822,N_479,N_340);
or U823 (N_823,N_225,N_99);
and U824 (N_824,N_262,N_219);
or U825 (N_825,N_153,N_145);
and U826 (N_826,N_97,N_462);
xnor U827 (N_827,N_346,N_403);
nor U828 (N_828,N_386,N_486);
and U829 (N_829,N_118,N_418);
nand U830 (N_830,N_438,N_84);
and U831 (N_831,N_174,N_49);
and U832 (N_832,N_138,N_450);
xnor U833 (N_833,N_287,N_169);
or U834 (N_834,N_124,N_356);
nor U835 (N_835,N_106,N_237);
or U836 (N_836,N_422,N_426);
nor U837 (N_837,N_30,N_486);
nand U838 (N_838,N_385,N_392);
or U839 (N_839,N_443,N_40);
and U840 (N_840,N_466,N_434);
and U841 (N_841,N_355,N_276);
nand U842 (N_842,N_333,N_363);
or U843 (N_843,N_122,N_314);
nor U844 (N_844,N_146,N_401);
and U845 (N_845,N_393,N_166);
or U846 (N_846,N_269,N_81);
or U847 (N_847,N_193,N_258);
nand U848 (N_848,N_450,N_344);
nand U849 (N_849,N_298,N_320);
and U850 (N_850,N_381,N_492);
nand U851 (N_851,N_212,N_138);
and U852 (N_852,N_377,N_125);
nand U853 (N_853,N_231,N_43);
nor U854 (N_854,N_16,N_403);
nand U855 (N_855,N_431,N_429);
nor U856 (N_856,N_31,N_336);
and U857 (N_857,N_199,N_325);
nor U858 (N_858,N_116,N_400);
xor U859 (N_859,N_416,N_427);
and U860 (N_860,N_324,N_482);
or U861 (N_861,N_394,N_240);
nand U862 (N_862,N_11,N_304);
nor U863 (N_863,N_215,N_375);
or U864 (N_864,N_306,N_210);
and U865 (N_865,N_239,N_34);
or U866 (N_866,N_391,N_94);
and U867 (N_867,N_269,N_211);
nand U868 (N_868,N_191,N_46);
nand U869 (N_869,N_293,N_0);
or U870 (N_870,N_62,N_152);
or U871 (N_871,N_65,N_104);
and U872 (N_872,N_382,N_226);
or U873 (N_873,N_406,N_358);
nand U874 (N_874,N_260,N_34);
nand U875 (N_875,N_62,N_413);
or U876 (N_876,N_375,N_424);
nor U877 (N_877,N_410,N_475);
xnor U878 (N_878,N_437,N_480);
nor U879 (N_879,N_251,N_382);
nand U880 (N_880,N_35,N_36);
nand U881 (N_881,N_303,N_327);
or U882 (N_882,N_424,N_166);
and U883 (N_883,N_35,N_460);
nor U884 (N_884,N_115,N_28);
nand U885 (N_885,N_490,N_135);
or U886 (N_886,N_12,N_384);
or U887 (N_887,N_80,N_455);
nor U888 (N_888,N_157,N_54);
and U889 (N_889,N_376,N_492);
or U890 (N_890,N_488,N_492);
or U891 (N_891,N_323,N_137);
nor U892 (N_892,N_316,N_295);
nor U893 (N_893,N_409,N_13);
xnor U894 (N_894,N_332,N_461);
nor U895 (N_895,N_287,N_4);
nand U896 (N_896,N_397,N_345);
nor U897 (N_897,N_153,N_477);
and U898 (N_898,N_231,N_254);
and U899 (N_899,N_91,N_38);
nand U900 (N_900,N_282,N_432);
nand U901 (N_901,N_156,N_185);
nand U902 (N_902,N_124,N_472);
nand U903 (N_903,N_174,N_284);
xor U904 (N_904,N_279,N_185);
and U905 (N_905,N_494,N_129);
and U906 (N_906,N_135,N_111);
or U907 (N_907,N_309,N_246);
or U908 (N_908,N_71,N_353);
nor U909 (N_909,N_156,N_18);
nand U910 (N_910,N_210,N_452);
nor U911 (N_911,N_338,N_334);
nand U912 (N_912,N_337,N_273);
and U913 (N_913,N_120,N_395);
or U914 (N_914,N_322,N_308);
nor U915 (N_915,N_489,N_365);
or U916 (N_916,N_89,N_98);
nand U917 (N_917,N_111,N_455);
or U918 (N_918,N_66,N_210);
and U919 (N_919,N_189,N_144);
or U920 (N_920,N_172,N_272);
nand U921 (N_921,N_157,N_337);
and U922 (N_922,N_243,N_91);
nand U923 (N_923,N_331,N_33);
nand U924 (N_924,N_255,N_3);
nand U925 (N_925,N_112,N_271);
and U926 (N_926,N_262,N_93);
and U927 (N_927,N_211,N_267);
or U928 (N_928,N_471,N_406);
or U929 (N_929,N_165,N_220);
or U930 (N_930,N_356,N_268);
nand U931 (N_931,N_146,N_46);
nor U932 (N_932,N_3,N_390);
or U933 (N_933,N_451,N_433);
nor U934 (N_934,N_447,N_305);
nor U935 (N_935,N_173,N_136);
nand U936 (N_936,N_231,N_476);
nand U937 (N_937,N_91,N_205);
or U938 (N_938,N_420,N_415);
nor U939 (N_939,N_229,N_188);
nor U940 (N_940,N_447,N_345);
nand U941 (N_941,N_496,N_251);
and U942 (N_942,N_88,N_152);
and U943 (N_943,N_411,N_312);
and U944 (N_944,N_492,N_304);
or U945 (N_945,N_230,N_158);
or U946 (N_946,N_140,N_428);
and U947 (N_947,N_271,N_258);
and U948 (N_948,N_413,N_433);
and U949 (N_949,N_98,N_472);
nor U950 (N_950,N_325,N_441);
and U951 (N_951,N_72,N_92);
or U952 (N_952,N_40,N_130);
nor U953 (N_953,N_185,N_349);
nand U954 (N_954,N_275,N_127);
nor U955 (N_955,N_79,N_269);
nor U956 (N_956,N_394,N_492);
and U957 (N_957,N_279,N_411);
nand U958 (N_958,N_108,N_161);
and U959 (N_959,N_488,N_61);
nand U960 (N_960,N_145,N_76);
and U961 (N_961,N_231,N_81);
nand U962 (N_962,N_117,N_56);
nand U963 (N_963,N_337,N_313);
nand U964 (N_964,N_318,N_2);
nand U965 (N_965,N_225,N_151);
nor U966 (N_966,N_348,N_300);
or U967 (N_967,N_334,N_359);
nand U968 (N_968,N_2,N_240);
and U969 (N_969,N_182,N_85);
and U970 (N_970,N_58,N_89);
and U971 (N_971,N_453,N_399);
nand U972 (N_972,N_481,N_85);
nand U973 (N_973,N_429,N_175);
nor U974 (N_974,N_160,N_189);
nor U975 (N_975,N_111,N_125);
and U976 (N_976,N_376,N_207);
nor U977 (N_977,N_124,N_170);
or U978 (N_978,N_135,N_229);
nand U979 (N_979,N_257,N_289);
and U980 (N_980,N_353,N_93);
or U981 (N_981,N_163,N_48);
and U982 (N_982,N_278,N_231);
and U983 (N_983,N_269,N_205);
and U984 (N_984,N_305,N_207);
nor U985 (N_985,N_70,N_120);
and U986 (N_986,N_89,N_119);
and U987 (N_987,N_357,N_294);
nand U988 (N_988,N_304,N_60);
and U989 (N_989,N_125,N_435);
nor U990 (N_990,N_44,N_249);
and U991 (N_991,N_197,N_99);
nand U992 (N_992,N_448,N_114);
nand U993 (N_993,N_398,N_380);
and U994 (N_994,N_133,N_394);
nand U995 (N_995,N_276,N_175);
or U996 (N_996,N_70,N_272);
or U997 (N_997,N_254,N_392);
xor U998 (N_998,N_240,N_347);
nand U999 (N_999,N_114,N_80);
nor U1000 (N_1000,N_880,N_820);
nor U1001 (N_1001,N_641,N_972);
nand U1002 (N_1002,N_976,N_857);
nand U1003 (N_1003,N_510,N_682);
nand U1004 (N_1004,N_518,N_526);
nand U1005 (N_1005,N_954,N_996);
or U1006 (N_1006,N_602,N_728);
or U1007 (N_1007,N_715,N_568);
nand U1008 (N_1008,N_765,N_712);
or U1009 (N_1009,N_872,N_590);
nand U1010 (N_1010,N_891,N_726);
nand U1011 (N_1011,N_612,N_595);
or U1012 (N_1012,N_981,N_901);
or U1013 (N_1013,N_893,N_779);
or U1014 (N_1014,N_713,N_608);
nor U1015 (N_1015,N_607,N_994);
or U1016 (N_1016,N_500,N_960);
nor U1017 (N_1017,N_830,N_883);
nor U1018 (N_1018,N_642,N_801);
nor U1019 (N_1019,N_906,N_787);
nor U1020 (N_1020,N_863,N_523);
nand U1021 (N_1021,N_747,N_889);
nand U1022 (N_1022,N_767,N_599);
or U1023 (N_1023,N_720,N_622);
nand U1024 (N_1024,N_977,N_986);
and U1025 (N_1025,N_967,N_625);
nand U1026 (N_1026,N_667,N_824);
nor U1027 (N_1027,N_845,N_885);
and U1028 (N_1028,N_604,N_714);
or U1029 (N_1029,N_818,N_882);
nor U1030 (N_1030,N_907,N_837);
and U1031 (N_1031,N_511,N_690);
and U1032 (N_1032,N_925,N_598);
and U1033 (N_1033,N_609,N_653);
or U1034 (N_1034,N_633,N_825);
nand U1035 (N_1035,N_640,N_763);
or U1036 (N_1036,N_528,N_742);
nor U1037 (N_1037,N_658,N_855);
nand U1038 (N_1038,N_538,N_797);
or U1039 (N_1039,N_563,N_521);
nand U1040 (N_1040,N_539,N_634);
and U1041 (N_1041,N_921,N_851);
nand U1042 (N_1042,N_852,N_811);
and U1043 (N_1043,N_744,N_927);
and U1044 (N_1044,N_639,N_803);
nor U1045 (N_1045,N_535,N_947);
nand U1046 (N_1046,N_847,N_616);
and U1047 (N_1047,N_950,N_694);
nand U1048 (N_1048,N_512,N_984);
nand U1049 (N_1049,N_541,N_740);
nor U1050 (N_1050,N_532,N_971);
and U1051 (N_1051,N_989,N_507);
nand U1052 (N_1052,N_773,N_887);
or U1053 (N_1053,N_681,N_566);
nor U1054 (N_1054,N_661,N_585);
nand U1055 (N_1055,N_513,N_644);
and U1056 (N_1056,N_540,N_549);
or U1057 (N_1057,N_696,N_544);
nand U1058 (N_1058,N_832,N_762);
nor U1059 (N_1059,N_809,N_716);
nand U1060 (N_1060,N_669,N_955);
nor U1061 (N_1061,N_517,N_973);
nor U1062 (N_1062,N_582,N_503);
and U1063 (N_1063,N_591,N_868);
and U1064 (N_1064,N_579,N_686);
and U1065 (N_1065,N_968,N_522);
nand U1066 (N_1066,N_623,N_516);
nor U1067 (N_1067,N_569,N_772);
or U1068 (N_1068,N_679,N_647);
and U1069 (N_1069,N_804,N_597);
and U1070 (N_1070,N_923,N_958);
or U1071 (N_1071,N_583,N_525);
or U1072 (N_1072,N_853,N_703);
nand U1073 (N_1073,N_865,N_869);
nand U1074 (N_1074,N_659,N_683);
nand U1075 (N_1075,N_542,N_561);
and U1076 (N_1076,N_769,N_547);
or U1077 (N_1077,N_939,N_905);
nor U1078 (N_1078,N_732,N_789);
or U1079 (N_1079,N_570,N_932);
and U1080 (N_1080,N_723,N_735);
nor U1081 (N_1081,N_731,N_506);
nand U1082 (N_1082,N_663,N_819);
nor U1083 (N_1083,N_738,N_613);
or U1084 (N_1084,N_838,N_618);
and U1085 (N_1085,N_788,N_778);
or U1086 (N_1086,N_688,N_861);
nand U1087 (N_1087,N_888,N_897);
or U1088 (N_1088,N_594,N_520);
or U1089 (N_1089,N_991,N_700);
nand U1090 (N_1090,N_993,N_926);
nand U1091 (N_1091,N_965,N_892);
and U1092 (N_1092,N_980,N_783);
and U1093 (N_1093,N_979,N_707);
nor U1094 (N_1094,N_527,N_550);
or U1095 (N_1095,N_890,N_760);
nor U1096 (N_1096,N_571,N_557);
or U1097 (N_1097,N_961,N_910);
and U1098 (N_1098,N_756,N_974);
nand U1099 (N_1099,N_737,N_812);
nand U1100 (N_1100,N_533,N_697);
nand U1101 (N_1101,N_759,N_722);
and U1102 (N_1102,N_578,N_922);
and U1103 (N_1103,N_822,N_813);
nand U1104 (N_1104,N_565,N_920);
nor U1105 (N_1105,N_963,N_805);
and U1106 (N_1106,N_970,N_514);
or U1107 (N_1107,N_687,N_877);
and U1108 (N_1108,N_724,N_791);
or U1109 (N_1109,N_727,N_648);
nand U1110 (N_1110,N_560,N_978);
or U1111 (N_1111,N_864,N_781);
and U1112 (N_1112,N_743,N_919);
nand U1113 (N_1113,N_501,N_628);
or U1114 (N_1114,N_534,N_733);
or U1115 (N_1115,N_992,N_775);
nand U1116 (N_1116,N_878,N_556);
or U1117 (N_1117,N_985,N_632);
nand U1118 (N_1118,N_933,N_748);
and U1119 (N_1119,N_706,N_867);
and U1120 (N_1120,N_580,N_531);
and U1121 (N_1121,N_677,N_530);
and U1122 (N_1122,N_678,N_646);
or U1123 (N_1123,N_903,N_546);
nor U1124 (N_1124,N_576,N_745);
and U1125 (N_1125,N_842,N_975);
nor U1126 (N_1126,N_827,N_701);
and U1127 (N_1127,N_573,N_596);
nor U1128 (N_1128,N_929,N_638);
or U1129 (N_1129,N_603,N_586);
nor U1130 (N_1130,N_940,N_806);
nand U1131 (N_1131,N_581,N_934);
nor U1132 (N_1132,N_784,N_785);
nand U1133 (N_1133,N_953,N_899);
or U1134 (N_1134,N_928,N_741);
nand U1135 (N_1135,N_873,N_721);
or U1136 (N_1136,N_957,N_699);
or U1137 (N_1137,N_758,N_635);
nor U1138 (N_1138,N_504,N_786);
and U1139 (N_1139,N_637,N_666);
or U1140 (N_1140,N_990,N_914);
and U1141 (N_1141,N_946,N_774);
nand U1142 (N_1142,N_524,N_770);
nor U1143 (N_1143,N_999,N_614);
and U1144 (N_1144,N_983,N_800);
or U1145 (N_1145,N_761,N_631);
and U1146 (N_1146,N_698,N_515);
nand U1147 (N_1147,N_601,N_898);
or U1148 (N_1148,N_719,N_502);
and U1149 (N_1149,N_691,N_705);
nor U1150 (N_1150,N_636,N_815);
nor U1151 (N_1151,N_757,N_917);
nand U1152 (N_1152,N_900,N_537);
or U1153 (N_1153,N_849,N_508);
nand U1154 (N_1154,N_876,N_587);
nand U1155 (N_1155,N_611,N_567);
nand U1156 (N_1156,N_749,N_650);
or U1157 (N_1157,N_850,N_997);
or U1158 (N_1158,N_718,N_693);
nand U1159 (N_1159,N_657,N_854);
nor U1160 (N_1160,N_895,N_816);
or U1161 (N_1161,N_710,N_952);
nor U1162 (N_1162,N_930,N_894);
nor U1163 (N_1163,N_998,N_552);
nor U1164 (N_1164,N_828,N_966);
and U1165 (N_1165,N_562,N_655);
nand U1166 (N_1166,N_665,N_871);
and U1167 (N_1167,N_776,N_643);
or U1168 (N_1168,N_771,N_629);
nand U1169 (N_1169,N_676,N_944);
and U1170 (N_1170,N_904,N_840);
and U1171 (N_1171,N_675,N_909);
nor U1172 (N_1172,N_754,N_729);
or U1173 (N_1173,N_833,N_555);
and U1174 (N_1174,N_935,N_680);
nor U1175 (N_1175,N_915,N_505);
nand U1176 (N_1176,N_795,N_575);
and U1177 (N_1177,N_793,N_746);
or U1178 (N_1178,N_617,N_689);
and U1179 (N_1179,N_600,N_685);
and U1180 (N_1180,N_777,N_630);
nand U1181 (N_1181,N_931,N_750);
or U1182 (N_1182,N_886,N_870);
nand U1183 (N_1183,N_821,N_624);
and U1184 (N_1184,N_964,N_823);
nand U1185 (N_1185,N_752,N_709);
and U1186 (N_1186,N_662,N_529);
nand U1187 (N_1187,N_558,N_913);
and U1188 (N_1188,N_936,N_551);
or U1189 (N_1189,N_792,N_652);
nor U1190 (N_1190,N_918,N_671);
and U1191 (N_1191,N_645,N_908);
and U1192 (N_1192,N_615,N_817);
and U1193 (N_1193,N_572,N_620);
and U1194 (N_1194,N_577,N_668);
and U1195 (N_1195,N_654,N_768);
and U1196 (N_1196,N_834,N_796);
nor U1197 (N_1197,N_559,N_937);
or U1198 (N_1198,N_651,N_969);
xor U1199 (N_1199,N_841,N_962);
nor U1200 (N_1200,N_672,N_945);
or U1201 (N_1201,N_798,N_995);
nor U1202 (N_1202,N_881,N_826);
and U1203 (N_1203,N_584,N_588);
or U1204 (N_1204,N_988,N_619);
and U1205 (N_1205,N_951,N_938);
nand U1206 (N_1206,N_941,N_725);
nor U1207 (N_1207,N_554,N_564);
nand U1208 (N_1208,N_702,N_649);
nand U1209 (N_1209,N_858,N_553);
nor U1210 (N_1210,N_626,N_835);
nand U1211 (N_1211,N_670,N_943);
nand U1212 (N_1212,N_660,N_692);
nand U1213 (N_1213,N_782,N_807);
nand U1214 (N_1214,N_751,N_704);
nor U1215 (N_1215,N_610,N_808);
xnor U1216 (N_1216,N_896,N_708);
and U1217 (N_1217,N_879,N_831);
or U1218 (N_1218,N_780,N_695);
nor U1219 (N_1219,N_949,N_860);
or U1220 (N_1220,N_673,N_589);
nand U1221 (N_1221,N_734,N_790);
or U1222 (N_1222,N_736,N_924);
nand U1223 (N_1223,N_574,N_753);
and U1224 (N_1224,N_545,N_843);
nor U1225 (N_1225,N_509,N_536);
nand U1226 (N_1226,N_605,N_814);
or U1227 (N_1227,N_846,N_839);
nand U1228 (N_1228,N_766,N_987);
or U1229 (N_1229,N_902,N_875);
nor U1230 (N_1230,N_848,N_656);
or U1231 (N_1231,N_711,N_911);
nand U1232 (N_1232,N_956,N_664);
nand U1233 (N_1233,N_866,N_717);
or U1234 (N_1234,N_859,N_593);
nor U1235 (N_1235,N_856,N_916);
nand U1236 (N_1236,N_862,N_884);
and U1237 (N_1237,N_959,N_739);
nor U1238 (N_1238,N_674,N_519);
nor U1239 (N_1239,N_592,N_794);
and U1240 (N_1240,N_755,N_810);
or U1241 (N_1241,N_829,N_543);
nor U1242 (N_1242,N_802,N_844);
nor U1243 (N_1243,N_621,N_684);
and U1244 (N_1244,N_836,N_874);
nor U1245 (N_1245,N_942,N_912);
or U1246 (N_1246,N_799,N_606);
and U1247 (N_1247,N_730,N_764);
nand U1248 (N_1248,N_548,N_982);
and U1249 (N_1249,N_627,N_948);
nand U1250 (N_1250,N_621,N_562);
and U1251 (N_1251,N_594,N_787);
or U1252 (N_1252,N_815,N_791);
nor U1253 (N_1253,N_519,N_769);
nand U1254 (N_1254,N_802,N_925);
and U1255 (N_1255,N_805,N_621);
or U1256 (N_1256,N_973,N_597);
or U1257 (N_1257,N_935,N_750);
nand U1258 (N_1258,N_568,N_619);
nor U1259 (N_1259,N_876,N_588);
nand U1260 (N_1260,N_580,N_813);
nor U1261 (N_1261,N_938,N_988);
nand U1262 (N_1262,N_695,N_645);
or U1263 (N_1263,N_721,N_558);
nor U1264 (N_1264,N_761,N_897);
nand U1265 (N_1265,N_633,N_502);
nand U1266 (N_1266,N_739,N_682);
nand U1267 (N_1267,N_908,N_782);
nor U1268 (N_1268,N_608,N_611);
nand U1269 (N_1269,N_664,N_757);
and U1270 (N_1270,N_605,N_912);
or U1271 (N_1271,N_779,N_572);
nand U1272 (N_1272,N_917,N_653);
nand U1273 (N_1273,N_934,N_644);
or U1274 (N_1274,N_672,N_669);
nor U1275 (N_1275,N_564,N_728);
nand U1276 (N_1276,N_640,N_607);
nand U1277 (N_1277,N_531,N_579);
or U1278 (N_1278,N_568,N_834);
nand U1279 (N_1279,N_708,N_950);
nand U1280 (N_1280,N_574,N_620);
nor U1281 (N_1281,N_978,N_781);
or U1282 (N_1282,N_671,N_848);
and U1283 (N_1283,N_847,N_934);
and U1284 (N_1284,N_735,N_530);
nor U1285 (N_1285,N_876,N_659);
or U1286 (N_1286,N_698,N_843);
nand U1287 (N_1287,N_603,N_661);
nand U1288 (N_1288,N_973,N_847);
nor U1289 (N_1289,N_939,N_527);
nor U1290 (N_1290,N_987,N_867);
and U1291 (N_1291,N_717,N_648);
or U1292 (N_1292,N_751,N_679);
nand U1293 (N_1293,N_513,N_640);
or U1294 (N_1294,N_827,N_810);
or U1295 (N_1295,N_784,N_993);
nand U1296 (N_1296,N_660,N_920);
or U1297 (N_1297,N_838,N_761);
nor U1298 (N_1298,N_833,N_535);
and U1299 (N_1299,N_695,N_801);
nand U1300 (N_1300,N_696,N_736);
nor U1301 (N_1301,N_616,N_832);
nand U1302 (N_1302,N_673,N_849);
or U1303 (N_1303,N_694,N_604);
nand U1304 (N_1304,N_695,N_520);
and U1305 (N_1305,N_746,N_757);
nor U1306 (N_1306,N_639,N_868);
nor U1307 (N_1307,N_756,N_871);
and U1308 (N_1308,N_750,N_679);
and U1309 (N_1309,N_905,N_645);
nand U1310 (N_1310,N_824,N_772);
nand U1311 (N_1311,N_893,N_502);
or U1312 (N_1312,N_837,N_631);
or U1313 (N_1313,N_807,N_629);
or U1314 (N_1314,N_773,N_904);
or U1315 (N_1315,N_921,N_654);
nor U1316 (N_1316,N_594,N_770);
or U1317 (N_1317,N_729,N_590);
and U1318 (N_1318,N_843,N_920);
nand U1319 (N_1319,N_975,N_574);
nor U1320 (N_1320,N_917,N_763);
nor U1321 (N_1321,N_576,N_992);
and U1322 (N_1322,N_617,N_978);
nand U1323 (N_1323,N_540,N_655);
nor U1324 (N_1324,N_639,N_795);
or U1325 (N_1325,N_934,N_627);
or U1326 (N_1326,N_750,N_609);
nand U1327 (N_1327,N_922,N_729);
nor U1328 (N_1328,N_650,N_628);
or U1329 (N_1329,N_945,N_897);
and U1330 (N_1330,N_873,N_936);
or U1331 (N_1331,N_840,N_590);
nand U1332 (N_1332,N_768,N_731);
and U1333 (N_1333,N_741,N_539);
or U1334 (N_1334,N_954,N_849);
nor U1335 (N_1335,N_611,N_905);
and U1336 (N_1336,N_779,N_914);
nand U1337 (N_1337,N_879,N_814);
nor U1338 (N_1338,N_682,N_530);
and U1339 (N_1339,N_685,N_648);
nand U1340 (N_1340,N_678,N_670);
and U1341 (N_1341,N_517,N_762);
nand U1342 (N_1342,N_542,N_832);
and U1343 (N_1343,N_526,N_589);
and U1344 (N_1344,N_754,N_566);
nor U1345 (N_1345,N_576,N_666);
or U1346 (N_1346,N_703,N_923);
nand U1347 (N_1347,N_663,N_842);
nand U1348 (N_1348,N_627,N_536);
or U1349 (N_1349,N_936,N_684);
or U1350 (N_1350,N_544,N_767);
and U1351 (N_1351,N_790,N_869);
nand U1352 (N_1352,N_682,N_586);
nand U1353 (N_1353,N_733,N_820);
nor U1354 (N_1354,N_707,N_665);
or U1355 (N_1355,N_861,N_655);
and U1356 (N_1356,N_785,N_717);
and U1357 (N_1357,N_709,N_927);
or U1358 (N_1358,N_905,N_598);
and U1359 (N_1359,N_950,N_618);
and U1360 (N_1360,N_589,N_977);
xor U1361 (N_1361,N_853,N_623);
and U1362 (N_1362,N_755,N_862);
or U1363 (N_1363,N_541,N_875);
and U1364 (N_1364,N_794,N_567);
nor U1365 (N_1365,N_917,N_527);
or U1366 (N_1366,N_682,N_524);
or U1367 (N_1367,N_831,N_545);
nor U1368 (N_1368,N_806,N_988);
nor U1369 (N_1369,N_775,N_510);
nand U1370 (N_1370,N_900,N_820);
or U1371 (N_1371,N_799,N_804);
or U1372 (N_1372,N_518,N_552);
nor U1373 (N_1373,N_534,N_644);
nand U1374 (N_1374,N_934,N_864);
or U1375 (N_1375,N_818,N_560);
nor U1376 (N_1376,N_541,N_865);
nor U1377 (N_1377,N_884,N_697);
and U1378 (N_1378,N_712,N_615);
and U1379 (N_1379,N_657,N_903);
and U1380 (N_1380,N_739,N_595);
nor U1381 (N_1381,N_721,N_662);
xnor U1382 (N_1382,N_903,N_919);
and U1383 (N_1383,N_722,N_902);
and U1384 (N_1384,N_821,N_909);
nand U1385 (N_1385,N_734,N_961);
nor U1386 (N_1386,N_504,N_740);
and U1387 (N_1387,N_753,N_737);
nor U1388 (N_1388,N_505,N_866);
nand U1389 (N_1389,N_625,N_950);
and U1390 (N_1390,N_599,N_715);
nand U1391 (N_1391,N_925,N_856);
and U1392 (N_1392,N_664,N_876);
or U1393 (N_1393,N_589,N_710);
nor U1394 (N_1394,N_737,N_511);
and U1395 (N_1395,N_702,N_876);
nor U1396 (N_1396,N_876,N_771);
nor U1397 (N_1397,N_803,N_888);
nor U1398 (N_1398,N_676,N_572);
or U1399 (N_1399,N_529,N_971);
nand U1400 (N_1400,N_636,N_803);
and U1401 (N_1401,N_645,N_812);
or U1402 (N_1402,N_955,N_855);
and U1403 (N_1403,N_975,N_705);
or U1404 (N_1404,N_739,N_768);
nor U1405 (N_1405,N_701,N_826);
or U1406 (N_1406,N_704,N_606);
or U1407 (N_1407,N_552,N_660);
nor U1408 (N_1408,N_930,N_893);
nand U1409 (N_1409,N_669,N_881);
nor U1410 (N_1410,N_540,N_531);
or U1411 (N_1411,N_711,N_761);
nand U1412 (N_1412,N_681,N_952);
and U1413 (N_1413,N_839,N_660);
and U1414 (N_1414,N_806,N_504);
nand U1415 (N_1415,N_660,N_697);
nor U1416 (N_1416,N_615,N_944);
nand U1417 (N_1417,N_586,N_612);
nor U1418 (N_1418,N_714,N_966);
nand U1419 (N_1419,N_923,N_570);
nor U1420 (N_1420,N_962,N_808);
or U1421 (N_1421,N_930,N_973);
nand U1422 (N_1422,N_557,N_597);
nor U1423 (N_1423,N_823,N_977);
and U1424 (N_1424,N_668,N_660);
and U1425 (N_1425,N_755,N_608);
nand U1426 (N_1426,N_661,N_842);
nor U1427 (N_1427,N_831,N_764);
nand U1428 (N_1428,N_887,N_830);
or U1429 (N_1429,N_610,N_837);
nor U1430 (N_1430,N_983,N_998);
nor U1431 (N_1431,N_548,N_980);
nand U1432 (N_1432,N_959,N_518);
or U1433 (N_1433,N_865,N_900);
nand U1434 (N_1434,N_572,N_726);
or U1435 (N_1435,N_760,N_712);
nand U1436 (N_1436,N_879,N_687);
and U1437 (N_1437,N_706,N_805);
nand U1438 (N_1438,N_869,N_675);
nor U1439 (N_1439,N_571,N_609);
nor U1440 (N_1440,N_765,N_930);
or U1441 (N_1441,N_729,N_897);
or U1442 (N_1442,N_996,N_892);
and U1443 (N_1443,N_891,N_803);
or U1444 (N_1444,N_857,N_577);
and U1445 (N_1445,N_506,N_581);
nand U1446 (N_1446,N_845,N_597);
and U1447 (N_1447,N_710,N_512);
nor U1448 (N_1448,N_882,N_736);
nor U1449 (N_1449,N_799,N_530);
nand U1450 (N_1450,N_865,N_836);
and U1451 (N_1451,N_936,N_901);
or U1452 (N_1452,N_522,N_735);
nand U1453 (N_1453,N_602,N_525);
nor U1454 (N_1454,N_673,N_506);
nand U1455 (N_1455,N_834,N_913);
nand U1456 (N_1456,N_734,N_624);
nor U1457 (N_1457,N_524,N_512);
nor U1458 (N_1458,N_513,N_855);
nor U1459 (N_1459,N_563,N_612);
nor U1460 (N_1460,N_740,N_954);
or U1461 (N_1461,N_563,N_876);
or U1462 (N_1462,N_998,N_630);
nor U1463 (N_1463,N_769,N_823);
nand U1464 (N_1464,N_772,N_938);
nor U1465 (N_1465,N_573,N_855);
or U1466 (N_1466,N_949,N_755);
and U1467 (N_1467,N_842,N_556);
nand U1468 (N_1468,N_753,N_971);
nand U1469 (N_1469,N_663,N_705);
or U1470 (N_1470,N_530,N_709);
nand U1471 (N_1471,N_612,N_946);
or U1472 (N_1472,N_745,N_927);
nand U1473 (N_1473,N_836,N_687);
nand U1474 (N_1474,N_763,N_696);
or U1475 (N_1475,N_706,N_584);
and U1476 (N_1476,N_672,N_695);
and U1477 (N_1477,N_661,N_981);
or U1478 (N_1478,N_742,N_939);
and U1479 (N_1479,N_517,N_710);
or U1480 (N_1480,N_965,N_614);
nand U1481 (N_1481,N_938,N_937);
or U1482 (N_1482,N_901,N_676);
or U1483 (N_1483,N_815,N_699);
or U1484 (N_1484,N_660,N_685);
nor U1485 (N_1485,N_686,N_949);
nand U1486 (N_1486,N_972,N_831);
or U1487 (N_1487,N_976,N_596);
and U1488 (N_1488,N_696,N_522);
nand U1489 (N_1489,N_738,N_843);
or U1490 (N_1490,N_781,N_951);
and U1491 (N_1491,N_702,N_720);
or U1492 (N_1492,N_888,N_712);
or U1493 (N_1493,N_586,N_538);
or U1494 (N_1494,N_827,N_764);
nand U1495 (N_1495,N_689,N_524);
or U1496 (N_1496,N_983,N_766);
nand U1497 (N_1497,N_748,N_734);
nor U1498 (N_1498,N_944,N_598);
nor U1499 (N_1499,N_768,N_638);
and U1500 (N_1500,N_1051,N_1055);
xor U1501 (N_1501,N_1220,N_1425);
nand U1502 (N_1502,N_1086,N_1208);
and U1503 (N_1503,N_1497,N_1126);
nand U1504 (N_1504,N_1291,N_1057);
nor U1505 (N_1505,N_1012,N_1016);
and U1506 (N_1506,N_1118,N_1495);
or U1507 (N_1507,N_1364,N_1329);
and U1508 (N_1508,N_1427,N_1370);
xnor U1509 (N_1509,N_1308,N_1139);
nand U1510 (N_1510,N_1150,N_1195);
nor U1511 (N_1511,N_1479,N_1352);
or U1512 (N_1512,N_1242,N_1353);
nand U1513 (N_1513,N_1009,N_1280);
nor U1514 (N_1514,N_1095,N_1162);
nor U1515 (N_1515,N_1363,N_1455);
nor U1516 (N_1516,N_1447,N_1035);
nand U1517 (N_1517,N_1018,N_1359);
or U1518 (N_1518,N_1458,N_1010);
and U1519 (N_1519,N_1309,N_1122);
and U1520 (N_1520,N_1380,N_1134);
nand U1521 (N_1521,N_1070,N_1428);
and U1522 (N_1522,N_1196,N_1266);
nor U1523 (N_1523,N_1171,N_1250);
or U1524 (N_1524,N_1194,N_1333);
or U1525 (N_1525,N_1264,N_1410);
and U1526 (N_1526,N_1330,N_1430);
or U1527 (N_1527,N_1384,N_1047);
nand U1528 (N_1528,N_1401,N_1338);
nand U1529 (N_1529,N_1043,N_1227);
and U1530 (N_1530,N_1015,N_1053);
nor U1531 (N_1531,N_1349,N_1324);
nor U1532 (N_1532,N_1046,N_1112);
and U1533 (N_1533,N_1409,N_1239);
nand U1534 (N_1534,N_1233,N_1222);
nand U1535 (N_1535,N_1300,N_1451);
nand U1536 (N_1536,N_1038,N_1391);
or U1537 (N_1537,N_1360,N_1056);
and U1538 (N_1538,N_1271,N_1140);
nor U1539 (N_1539,N_1002,N_1007);
nand U1540 (N_1540,N_1178,N_1302);
and U1541 (N_1541,N_1022,N_1375);
nand U1542 (N_1542,N_1444,N_1031);
nand U1543 (N_1543,N_1092,N_1422);
and U1544 (N_1544,N_1268,N_1245);
nand U1545 (N_1545,N_1200,N_1164);
and U1546 (N_1546,N_1151,N_1386);
nand U1547 (N_1547,N_1439,N_1045);
or U1548 (N_1548,N_1412,N_1243);
nand U1549 (N_1549,N_1340,N_1026);
nand U1550 (N_1550,N_1481,N_1199);
nor U1551 (N_1551,N_1120,N_1485);
nor U1552 (N_1552,N_1131,N_1322);
nor U1553 (N_1553,N_1278,N_1442);
nor U1554 (N_1554,N_1163,N_1411);
and U1555 (N_1555,N_1385,N_1350);
or U1556 (N_1556,N_1211,N_1377);
nor U1557 (N_1557,N_1389,N_1307);
and U1558 (N_1558,N_1068,N_1011);
and U1559 (N_1559,N_1480,N_1437);
nor U1560 (N_1560,N_1235,N_1170);
or U1561 (N_1561,N_1282,N_1101);
nor U1562 (N_1562,N_1473,N_1418);
nor U1563 (N_1563,N_1339,N_1251);
or U1564 (N_1564,N_1323,N_1269);
nor U1565 (N_1565,N_1314,N_1464);
nand U1566 (N_1566,N_1079,N_1064);
nor U1567 (N_1567,N_1023,N_1260);
nand U1568 (N_1568,N_1219,N_1029);
nand U1569 (N_1569,N_1127,N_1017);
nor U1570 (N_1570,N_1348,N_1311);
nor U1571 (N_1571,N_1335,N_1225);
or U1572 (N_1572,N_1438,N_1144);
nor U1573 (N_1573,N_1261,N_1417);
nand U1574 (N_1574,N_1265,N_1137);
nand U1575 (N_1575,N_1248,N_1492);
and U1576 (N_1576,N_1310,N_1491);
nand U1577 (N_1577,N_1147,N_1087);
and U1578 (N_1578,N_1077,N_1298);
nor U1579 (N_1579,N_1080,N_1406);
nand U1580 (N_1580,N_1423,N_1072);
nor U1581 (N_1581,N_1099,N_1097);
and U1582 (N_1582,N_1237,N_1180);
and U1583 (N_1583,N_1441,N_1136);
or U1584 (N_1584,N_1123,N_1149);
nand U1585 (N_1585,N_1109,N_1416);
nor U1586 (N_1586,N_1284,N_1419);
and U1587 (N_1587,N_1050,N_1244);
or U1588 (N_1588,N_1175,N_1334);
and U1589 (N_1589,N_1078,N_1138);
nand U1590 (N_1590,N_1341,N_1347);
or U1591 (N_1591,N_1117,N_1273);
nor U1592 (N_1592,N_1223,N_1482);
or U1593 (N_1593,N_1212,N_1082);
nand U1594 (N_1594,N_1270,N_1254);
or U1595 (N_1595,N_1289,N_1484);
nand U1596 (N_1596,N_1318,N_1294);
and U1597 (N_1597,N_1295,N_1033);
or U1598 (N_1598,N_1403,N_1125);
and U1599 (N_1599,N_1081,N_1189);
and U1600 (N_1600,N_1332,N_1257);
and U1601 (N_1601,N_1141,N_1096);
and U1602 (N_1602,N_1305,N_1454);
nor U1603 (N_1603,N_1108,N_1106);
nand U1604 (N_1604,N_1342,N_1283);
and U1605 (N_1605,N_1019,N_1207);
and U1606 (N_1606,N_1008,N_1148);
nand U1607 (N_1607,N_1069,N_1119);
nor U1608 (N_1608,N_1299,N_1059);
xnor U1609 (N_1609,N_1037,N_1191);
or U1610 (N_1610,N_1111,N_1337);
and U1611 (N_1611,N_1316,N_1240);
xor U1612 (N_1612,N_1368,N_1303);
nor U1613 (N_1613,N_1467,N_1496);
or U1614 (N_1614,N_1286,N_1474);
or U1615 (N_1615,N_1071,N_1061);
nand U1616 (N_1616,N_1321,N_1249);
nor U1617 (N_1617,N_1312,N_1256);
nor U1618 (N_1618,N_1020,N_1159);
nand U1619 (N_1619,N_1469,N_1446);
nor U1620 (N_1620,N_1434,N_1471);
or U1621 (N_1621,N_1102,N_1408);
nor U1622 (N_1622,N_1371,N_1355);
nand U1623 (N_1623,N_1396,N_1490);
nand U1624 (N_1624,N_1301,N_1392);
nand U1625 (N_1625,N_1030,N_1293);
xnor U1626 (N_1626,N_1165,N_1487);
or U1627 (N_1627,N_1493,N_1004);
or U1628 (N_1628,N_1381,N_1133);
and U1629 (N_1629,N_1076,N_1470);
or U1630 (N_1630,N_1445,N_1452);
or U1631 (N_1631,N_1486,N_1440);
nand U1632 (N_1632,N_1263,N_1367);
nor U1633 (N_1633,N_1168,N_1477);
or U1634 (N_1634,N_1346,N_1083);
nand U1635 (N_1635,N_1098,N_1229);
nand U1636 (N_1636,N_1190,N_1267);
nand U1637 (N_1637,N_1325,N_1369);
nor U1638 (N_1638,N_1317,N_1104);
nor U1639 (N_1639,N_1252,N_1093);
or U1640 (N_1640,N_1028,N_1177);
xnor U1641 (N_1641,N_1166,N_1049);
nand U1642 (N_1642,N_1431,N_1400);
or U1643 (N_1643,N_1376,N_1304);
nor U1644 (N_1644,N_1063,N_1054);
nand U1645 (N_1645,N_1357,N_1090);
or U1646 (N_1646,N_1358,N_1404);
or U1647 (N_1647,N_1209,N_1272);
nor U1648 (N_1648,N_1172,N_1152);
nor U1649 (N_1649,N_1382,N_1459);
and U1650 (N_1650,N_1456,N_1005);
nand U1651 (N_1651,N_1281,N_1494);
nand U1652 (N_1652,N_1036,N_1421);
or U1653 (N_1653,N_1218,N_1021);
nand U1654 (N_1654,N_1292,N_1453);
and U1655 (N_1655,N_1203,N_1183);
and U1656 (N_1656,N_1041,N_1088);
and U1657 (N_1657,N_1279,N_1184);
nand U1658 (N_1658,N_1187,N_1230);
nand U1659 (N_1659,N_1429,N_1013);
nand U1660 (N_1660,N_1356,N_1206);
nor U1661 (N_1661,N_1062,N_1145);
nand U1662 (N_1662,N_1024,N_1488);
and U1663 (N_1663,N_1277,N_1146);
or U1664 (N_1664,N_1085,N_1449);
nand U1665 (N_1665,N_1114,N_1142);
and U1666 (N_1666,N_1226,N_1132);
nand U1667 (N_1667,N_1498,N_1001);
or U1668 (N_1668,N_1306,N_1383);
and U1669 (N_1669,N_1420,N_1228);
nor U1670 (N_1670,N_1124,N_1135);
and U1671 (N_1671,N_1048,N_1204);
or U1672 (N_1672,N_1014,N_1489);
and U1673 (N_1673,N_1378,N_1231);
nor U1674 (N_1674,N_1326,N_1331);
and U1675 (N_1675,N_1372,N_1320);
xor U1676 (N_1676,N_1398,N_1236);
nor U1677 (N_1677,N_1052,N_1067);
nand U1678 (N_1678,N_1472,N_1394);
xor U1679 (N_1679,N_1433,N_1192);
or U1680 (N_1680,N_1032,N_1457);
and U1681 (N_1681,N_1399,N_1275);
or U1682 (N_1682,N_1259,N_1432);
and U1683 (N_1683,N_1193,N_1328);
or U1684 (N_1684,N_1084,N_1110);
and U1685 (N_1685,N_1169,N_1130);
nor U1686 (N_1686,N_1197,N_1006);
or U1687 (N_1687,N_1468,N_1094);
and U1688 (N_1688,N_1361,N_1216);
and U1689 (N_1689,N_1176,N_1224);
and U1690 (N_1690,N_1129,N_1414);
and U1691 (N_1691,N_1091,N_1465);
and U1692 (N_1692,N_1379,N_1089);
and U1693 (N_1693,N_1167,N_1365);
or U1694 (N_1694,N_1246,N_1201);
and U1695 (N_1695,N_1158,N_1424);
nand U1696 (N_1696,N_1460,N_1040);
nand U1697 (N_1697,N_1215,N_1074);
nor U1698 (N_1698,N_1436,N_1255);
or U1699 (N_1699,N_1060,N_1362);
nor U1700 (N_1700,N_1287,N_1039);
nand U1701 (N_1701,N_1156,N_1044);
nor U1702 (N_1702,N_1405,N_1327);
and U1703 (N_1703,N_1402,N_1027);
or U1704 (N_1704,N_1395,N_1160);
nor U1705 (N_1705,N_1448,N_1407);
nand U1706 (N_1706,N_1499,N_1182);
nor U1707 (N_1707,N_1366,N_1107);
nor U1708 (N_1708,N_1185,N_1354);
or U1709 (N_1709,N_1413,N_1116);
or U1710 (N_1710,N_1290,N_1387);
nor U1711 (N_1711,N_1258,N_1397);
or U1712 (N_1712,N_1345,N_1393);
nor U1713 (N_1713,N_1221,N_1475);
nor U1714 (N_1714,N_1313,N_1435);
or U1715 (N_1715,N_1463,N_1154);
or U1716 (N_1716,N_1415,N_1241);
nor U1717 (N_1717,N_1262,N_1000);
or U1718 (N_1718,N_1234,N_1483);
and U1719 (N_1719,N_1297,N_1157);
or U1720 (N_1720,N_1274,N_1161);
and U1721 (N_1721,N_1247,N_1285);
or U1722 (N_1722,N_1153,N_1476);
nor U1723 (N_1723,N_1034,N_1103);
nor U1724 (N_1724,N_1205,N_1121);
nor U1725 (N_1725,N_1374,N_1066);
or U1726 (N_1726,N_1443,N_1343);
nand U1727 (N_1727,N_1188,N_1042);
nor U1728 (N_1728,N_1288,N_1025);
and U1729 (N_1729,N_1276,N_1373);
or U1730 (N_1730,N_1073,N_1214);
nand U1731 (N_1731,N_1003,N_1058);
nand U1732 (N_1732,N_1065,N_1319);
or U1733 (N_1733,N_1115,N_1336);
or U1734 (N_1734,N_1213,N_1113);
and U1735 (N_1735,N_1155,N_1296);
and U1736 (N_1736,N_1186,N_1461);
or U1737 (N_1737,N_1179,N_1388);
nor U1738 (N_1738,N_1478,N_1128);
nor U1739 (N_1739,N_1253,N_1232);
nand U1740 (N_1740,N_1105,N_1174);
and U1741 (N_1741,N_1466,N_1344);
and U1742 (N_1742,N_1426,N_1210);
nor U1743 (N_1743,N_1198,N_1075);
nand U1744 (N_1744,N_1173,N_1351);
or U1745 (N_1745,N_1390,N_1315);
and U1746 (N_1746,N_1462,N_1181);
and U1747 (N_1747,N_1450,N_1143);
nor U1748 (N_1748,N_1217,N_1100);
or U1749 (N_1749,N_1238,N_1202);
nand U1750 (N_1750,N_1440,N_1352);
nor U1751 (N_1751,N_1008,N_1215);
or U1752 (N_1752,N_1337,N_1216);
nand U1753 (N_1753,N_1254,N_1114);
or U1754 (N_1754,N_1474,N_1031);
nand U1755 (N_1755,N_1346,N_1485);
nand U1756 (N_1756,N_1073,N_1477);
nor U1757 (N_1757,N_1299,N_1032);
nor U1758 (N_1758,N_1317,N_1265);
or U1759 (N_1759,N_1395,N_1167);
or U1760 (N_1760,N_1227,N_1473);
nand U1761 (N_1761,N_1483,N_1452);
and U1762 (N_1762,N_1059,N_1315);
and U1763 (N_1763,N_1273,N_1282);
nor U1764 (N_1764,N_1341,N_1063);
nor U1765 (N_1765,N_1061,N_1350);
and U1766 (N_1766,N_1102,N_1283);
and U1767 (N_1767,N_1150,N_1194);
and U1768 (N_1768,N_1277,N_1385);
nand U1769 (N_1769,N_1162,N_1295);
nand U1770 (N_1770,N_1356,N_1411);
or U1771 (N_1771,N_1181,N_1307);
nor U1772 (N_1772,N_1431,N_1057);
nand U1773 (N_1773,N_1454,N_1428);
nor U1774 (N_1774,N_1128,N_1473);
or U1775 (N_1775,N_1300,N_1426);
nand U1776 (N_1776,N_1399,N_1005);
nor U1777 (N_1777,N_1422,N_1006);
nand U1778 (N_1778,N_1463,N_1231);
or U1779 (N_1779,N_1469,N_1084);
and U1780 (N_1780,N_1427,N_1300);
xor U1781 (N_1781,N_1076,N_1100);
nand U1782 (N_1782,N_1153,N_1254);
nor U1783 (N_1783,N_1150,N_1297);
nand U1784 (N_1784,N_1380,N_1291);
nand U1785 (N_1785,N_1016,N_1013);
and U1786 (N_1786,N_1010,N_1154);
xnor U1787 (N_1787,N_1195,N_1447);
nor U1788 (N_1788,N_1099,N_1349);
or U1789 (N_1789,N_1272,N_1491);
and U1790 (N_1790,N_1440,N_1058);
nand U1791 (N_1791,N_1163,N_1104);
nor U1792 (N_1792,N_1441,N_1366);
or U1793 (N_1793,N_1149,N_1261);
or U1794 (N_1794,N_1494,N_1436);
or U1795 (N_1795,N_1332,N_1137);
nor U1796 (N_1796,N_1371,N_1383);
nor U1797 (N_1797,N_1293,N_1344);
and U1798 (N_1798,N_1224,N_1198);
or U1799 (N_1799,N_1215,N_1050);
or U1800 (N_1800,N_1489,N_1448);
and U1801 (N_1801,N_1446,N_1407);
nor U1802 (N_1802,N_1034,N_1242);
and U1803 (N_1803,N_1248,N_1130);
nand U1804 (N_1804,N_1300,N_1394);
nor U1805 (N_1805,N_1131,N_1258);
and U1806 (N_1806,N_1266,N_1473);
nor U1807 (N_1807,N_1414,N_1307);
and U1808 (N_1808,N_1015,N_1242);
nor U1809 (N_1809,N_1338,N_1228);
nor U1810 (N_1810,N_1324,N_1030);
and U1811 (N_1811,N_1451,N_1225);
nor U1812 (N_1812,N_1495,N_1328);
nor U1813 (N_1813,N_1461,N_1476);
nor U1814 (N_1814,N_1083,N_1162);
or U1815 (N_1815,N_1057,N_1197);
and U1816 (N_1816,N_1475,N_1268);
nand U1817 (N_1817,N_1095,N_1008);
nand U1818 (N_1818,N_1220,N_1093);
nand U1819 (N_1819,N_1240,N_1161);
nand U1820 (N_1820,N_1192,N_1424);
nand U1821 (N_1821,N_1433,N_1272);
and U1822 (N_1822,N_1479,N_1279);
or U1823 (N_1823,N_1246,N_1285);
nor U1824 (N_1824,N_1213,N_1337);
nand U1825 (N_1825,N_1241,N_1350);
and U1826 (N_1826,N_1432,N_1115);
nand U1827 (N_1827,N_1201,N_1258);
nand U1828 (N_1828,N_1108,N_1237);
or U1829 (N_1829,N_1428,N_1349);
or U1830 (N_1830,N_1034,N_1314);
and U1831 (N_1831,N_1425,N_1326);
and U1832 (N_1832,N_1385,N_1092);
and U1833 (N_1833,N_1099,N_1183);
nand U1834 (N_1834,N_1113,N_1073);
and U1835 (N_1835,N_1109,N_1304);
or U1836 (N_1836,N_1332,N_1388);
nor U1837 (N_1837,N_1239,N_1240);
or U1838 (N_1838,N_1008,N_1290);
or U1839 (N_1839,N_1306,N_1415);
xor U1840 (N_1840,N_1222,N_1358);
nand U1841 (N_1841,N_1404,N_1326);
nor U1842 (N_1842,N_1018,N_1070);
nand U1843 (N_1843,N_1416,N_1107);
and U1844 (N_1844,N_1407,N_1485);
or U1845 (N_1845,N_1212,N_1327);
nand U1846 (N_1846,N_1344,N_1324);
and U1847 (N_1847,N_1467,N_1348);
or U1848 (N_1848,N_1053,N_1183);
and U1849 (N_1849,N_1374,N_1372);
and U1850 (N_1850,N_1435,N_1009);
and U1851 (N_1851,N_1175,N_1225);
nand U1852 (N_1852,N_1315,N_1464);
or U1853 (N_1853,N_1232,N_1085);
and U1854 (N_1854,N_1275,N_1159);
or U1855 (N_1855,N_1184,N_1395);
or U1856 (N_1856,N_1344,N_1218);
nand U1857 (N_1857,N_1104,N_1185);
nand U1858 (N_1858,N_1139,N_1146);
nand U1859 (N_1859,N_1320,N_1161);
nor U1860 (N_1860,N_1133,N_1418);
and U1861 (N_1861,N_1413,N_1355);
nor U1862 (N_1862,N_1081,N_1330);
and U1863 (N_1863,N_1020,N_1321);
nor U1864 (N_1864,N_1177,N_1157);
and U1865 (N_1865,N_1420,N_1359);
or U1866 (N_1866,N_1370,N_1029);
or U1867 (N_1867,N_1334,N_1365);
nand U1868 (N_1868,N_1101,N_1203);
and U1869 (N_1869,N_1457,N_1290);
or U1870 (N_1870,N_1164,N_1289);
or U1871 (N_1871,N_1017,N_1116);
nor U1872 (N_1872,N_1176,N_1470);
or U1873 (N_1873,N_1383,N_1364);
and U1874 (N_1874,N_1108,N_1292);
or U1875 (N_1875,N_1249,N_1460);
and U1876 (N_1876,N_1392,N_1486);
nor U1877 (N_1877,N_1200,N_1322);
or U1878 (N_1878,N_1264,N_1340);
nand U1879 (N_1879,N_1306,N_1311);
nand U1880 (N_1880,N_1268,N_1021);
and U1881 (N_1881,N_1323,N_1217);
and U1882 (N_1882,N_1428,N_1081);
nand U1883 (N_1883,N_1356,N_1092);
and U1884 (N_1884,N_1273,N_1084);
nor U1885 (N_1885,N_1372,N_1107);
nor U1886 (N_1886,N_1035,N_1176);
or U1887 (N_1887,N_1189,N_1070);
and U1888 (N_1888,N_1420,N_1047);
or U1889 (N_1889,N_1334,N_1499);
or U1890 (N_1890,N_1055,N_1086);
nor U1891 (N_1891,N_1087,N_1153);
or U1892 (N_1892,N_1486,N_1255);
nand U1893 (N_1893,N_1215,N_1245);
or U1894 (N_1894,N_1088,N_1442);
nor U1895 (N_1895,N_1357,N_1031);
or U1896 (N_1896,N_1390,N_1287);
or U1897 (N_1897,N_1400,N_1175);
nand U1898 (N_1898,N_1300,N_1032);
or U1899 (N_1899,N_1054,N_1139);
and U1900 (N_1900,N_1038,N_1468);
and U1901 (N_1901,N_1290,N_1302);
or U1902 (N_1902,N_1158,N_1278);
nand U1903 (N_1903,N_1049,N_1352);
nand U1904 (N_1904,N_1175,N_1267);
or U1905 (N_1905,N_1476,N_1497);
nand U1906 (N_1906,N_1035,N_1175);
nand U1907 (N_1907,N_1203,N_1181);
nor U1908 (N_1908,N_1257,N_1194);
nor U1909 (N_1909,N_1393,N_1379);
or U1910 (N_1910,N_1093,N_1074);
or U1911 (N_1911,N_1081,N_1455);
nor U1912 (N_1912,N_1330,N_1168);
or U1913 (N_1913,N_1116,N_1169);
nand U1914 (N_1914,N_1296,N_1398);
or U1915 (N_1915,N_1467,N_1002);
or U1916 (N_1916,N_1467,N_1318);
nor U1917 (N_1917,N_1383,N_1282);
nor U1918 (N_1918,N_1434,N_1482);
and U1919 (N_1919,N_1091,N_1102);
nand U1920 (N_1920,N_1464,N_1229);
nand U1921 (N_1921,N_1431,N_1409);
nand U1922 (N_1922,N_1217,N_1252);
nand U1923 (N_1923,N_1421,N_1302);
nor U1924 (N_1924,N_1376,N_1087);
or U1925 (N_1925,N_1444,N_1110);
and U1926 (N_1926,N_1206,N_1398);
or U1927 (N_1927,N_1083,N_1039);
and U1928 (N_1928,N_1447,N_1352);
and U1929 (N_1929,N_1314,N_1343);
or U1930 (N_1930,N_1025,N_1325);
and U1931 (N_1931,N_1495,N_1138);
nor U1932 (N_1932,N_1348,N_1274);
and U1933 (N_1933,N_1411,N_1328);
nand U1934 (N_1934,N_1194,N_1328);
nand U1935 (N_1935,N_1151,N_1404);
nand U1936 (N_1936,N_1007,N_1426);
nor U1937 (N_1937,N_1062,N_1472);
nand U1938 (N_1938,N_1308,N_1339);
nand U1939 (N_1939,N_1486,N_1030);
and U1940 (N_1940,N_1084,N_1220);
xor U1941 (N_1941,N_1057,N_1065);
and U1942 (N_1942,N_1156,N_1233);
and U1943 (N_1943,N_1137,N_1050);
nor U1944 (N_1944,N_1326,N_1214);
nor U1945 (N_1945,N_1298,N_1453);
or U1946 (N_1946,N_1088,N_1406);
or U1947 (N_1947,N_1313,N_1245);
nor U1948 (N_1948,N_1115,N_1010);
and U1949 (N_1949,N_1277,N_1462);
nand U1950 (N_1950,N_1469,N_1074);
or U1951 (N_1951,N_1099,N_1325);
and U1952 (N_1952,N_1392,N_1047);
or U1953 (N_1953,N_1292,N_1192);
nor U1954 (N_1954,N_1323,N_1105);
or U1955 (N_1955,N_1149,N_1026);
or U1956 (N_1956,N_1376,N_1481);
and U1957 (N_1957,N_1295,N_1385);
nor U1958 (N_1958,N_1383,N_1319);
or U1959 (N_1959,N_1321,N_1017);
and U1960 (N_1960,N_1467,N_1051);
nor U1961 (N_1961,N_1158,N_1408);
or U1962 (N_1962,N_1078,N_1402);
and U1963 (N_1963,N_1355,N_1303);
and U1964 (N_1964,N_1240,N_1293);
nand U1965 (N_1965,N_1388,N_1341);
nand U1966 (N_1966,N_1085,N_1305);
and U1967 (N_1967,N_1084,N_1280);
or U1968 (N_1968,N_1266,N_1060);
nor U1969 (N_1969,N_1265,N_1100);
nor U1970 (N_1970,N_1408,N_1075);
or U1971 (N_1971,N_1401,N_1383);
and U1972 (N_1972,N_1289,N_1273);
and U1973 (N_1973,N_1014,N_1005);
nor U1974 (N_1974,N_1272,N_1481);
nor U1975 (N_1975,N_1089,N_1021);
nand U1976 (N_1976,N_1314,N_1229);
nand U1977 (N_1977,N_1258,N_1495);
xor U1978 (N_1978,N_1077,N_1010);
or U1979 (N_1979,N_1390,N_1129);
nor U1980 (N_1980,N_1475,N_1027);
nand U1981 (N_1981,N_1066,N_1290);
nor U1982 (N_1982,N_1031,N_1117);
nand U1983 (N_1983,N_1212,N_1488);
and U1984 (N_1984,N_1324,N_1495);
nor U1985 (N_1985,N_1484,N_1025);
or U1986 (N_1986,N_1051,N_1057);
nor U1987 (N_1987,N_1149,N_1058);
nand U1988 (N_1988,N_1465,N_1127);
nor U1989 (N_1989,N_1176,N_1225);
nor U1990 (N_1990,N_1095,N_1318);
and U1991 (N_1991,N_1233,N_1437);
or U1992 (N_1992,N_1191,N_1459);
and U1993 (N_1993,N_1343,N_1072);
or U1994 (N_1994,N_1194,N_1002);
nand U1995 (N_1995,N_1424,N_1300);
nor U1996 (N_1996,N_1166,N_1087);
nand U1997 (N_1997,N_1088,N_1133);
or U1998 (N_1998,N_1099,N_1107);
and U1999 (N_1999,N_1485,N_1317);
or U2000 (N_2000,N_1851,N_1954);
nor U2001 (N_2001,N_1769,N_1876);
nor U2002 (N_2002,N_1818,N_1744);
or U2003 (N_2003,N_1790,N_1674);
or U2004 (N_2004,N_1524,N_1515);
and U2005 (N_2005,N_1574,N_1732);
and U2006 (N_2006,N_1779,N_1770);
or U2007 (N_2007,N_1671,N_1588);
and U2008 (N_2008,N_1705,N_1889);
or U2009 (N_2009,N_1727,N_1942);
nand U2010 (N_2010,N_1991,N_1605);
nand U2011 (N_2011,N_1535,N_1739);
and U2012 (N_2012,N_1645,N_1714);
and U2013 (N_2013,N_1716,N_1718);
and U2014 (N_2014,N_1618,N_1927);
or U2015 (N_2015,N_1850,N_1835);
nand U2016 (N_2016,N_1661,N_1890);
nand U2017 (N_2017,N_1960,N_1776);
nor U2018 (N_2018,N_1978,N_1831);
nor U2019 (N_2019,N_1723,N_1931);
and U2020 (N_2020,N_1803,N_1703);
and U2021 (N_2021,N_1655,N_1575);
and U2022 (N_2022,N_1623,N_1611);
or U2023 (N_2023,N_1741,N_1901);
and U2024 (N_2024,N_1914,N_1865);
nand U2025 (N_2025,N_1516,N_1654);
nand U2026 (N_2026,N_1713,N_1911);
nand U2027 (N_2027,N_1875,N_1893);
and U2028 (N_2028,N_1657,N_1502);
nand U2029 (N_2029,N_1992,N_1707);
or U2030 (N_2030,N_1936,N_1582);
or U2031 (N_2031,N_1529,N_1563);
nor U2032 (N_2032,N_1952,N_1912);
nand U2033 (N_2033,N_1692,N_1728);
nand U2034 (N_2034,N_1640,N_1847);
or U2035 (N_2035,N_1855,N_1988);
nand U2036 (N_2036,N_1682,N_1974);
nand U2037 (N_2037,N_1903,N_1780);
nor U2038 (N_2038,N_1888,N_1816);
and U2039 (N_2039,N_1787,N_1798);
and U2040 (N_2040,N_1965,N_1709);
nor U2041 (N_2041,N_1804,N_1530);
nor U2042 (N_2042,N_1971,N_1885);
nand U2043 (N_2043,N_1592,N_1793);
and U2044 (N_2044,N_1698,N_1670);
and U2045 (N_2045,N_1843,N_1948);
and U2046 (N_2046,N_1724,N_1648);
nand U2047 (N_2047,N_1570,N_1700);
nand U2048 (N_2048,N_1533,N_1603);
and U2049 (N_2049,N_1937,N_1797);
and U2050 (N_2050,N_1925,N_1800);
or U2051 (N_2051,N_1870,N_1677);
nor U2052 (N_2052,N_1848,N_1753);
or U2053 (N_2053,N_1869,N_1560);
nor U2054 (N_2054,N_1627,N_1567);
nor U2055 (N_2055,N_1915,N_1896);
nand U2056 (N_2056,N_1726,N_1695);
and U2057 (N_2057,N_1636,N_1839);
or U2058 (N_2058,N_1752,N_1676);
nor U2059 (N_2059,N_1913,N_1823);
and U2060 (N_2060,N_1842,N_1759);
nor U2061 (N_2061,N_1836,N_1544);
nor U2062 (N_2062,N_1833,N_1970);
and U2063 (N_2063,N_1616,N_1782);
nand U2064 (N_2064,N_1922,N_1987);
nand U2065 (N_2065,N_1550,N_1928);
nor U2066 (N_2066,N_1788,N_1539);
xor U2067 (N_2067,N_1774,N_1761);
nor U2068 (N_2068,N_1555,N_1975);
or U2069 (N_2069,N_1747,N_1950);
nand U2070 (N_2070,N_1758,N_1825);
nand U2071 (N_2071,N_1969,N_1838);
nor U2072 (N_2072,N_1610,N_1880);
or U2073 (N_2073,N_1527,N_1680);
nor U2074 (N_2074,N_1762,N_1900);
and U2075 (N_2075,N_1600,N_1773);
nor U2076 (N_2076,N_1522,N_1660);
or U2077 (N_2077,N_1943,N_1557);
nor U2078 (N_2078,N_1540,N_1568);
nand U2079 (N_2079,N_1523,N_1679);
nor U2080 (N_2080,N_1853,N_1725);
nand U2081 (N_2081,N_1849,N_1852);
nand U2082 (N_2082,N_1829,N_1972);
or U2083 (N_2083,N_1733,N_1646);
and U2084 (N_2084,N_1926,N_1589);
nand U2085 (N_2085,N_1534,N_1772);
nor U2086 (N_2086,N_1897,N_1822);
and U2087 (N_2087,N_1641,N_1510);
nor U2088 (N_2088,N_1854,N_1564);
and U2089 (N_2089,N_1608,N_1979);
or U2090 (N_2090,N_1968,N_1626);
nand U2091 (N_2091,N_1520,N_1580);
nor U2092 (N_2092,N_1953,N_1697);
or U2093 (N_2093,N_1509,N_1919);
and U2094 (N_2094,N_1945,N_1678);
and U2095 (N_2095,N_1559,N_1612);
or U2096 (N_2096,N_1808,N_1624);
or U2097 (N_2097,N_1781,N_1528);
and U2098 (N_2098,N_1899,N_1558);
and U2099 (N_2099,N_1710,N_1916);
nand U2100 (N_2100,N_1814,N_1989);
nor U2101 (N_2101,N_1628,N_1811);
nand U2102 (N_2102,N_1826,N_1751);
nor U2103 (N_2103,N_1562,N_1956);
or U2104 (N_2104,N_1754,N_1879);
and U2105 (N_2105,N_1859,N_1569);
nor U2106 (N_2106,N_1663,N_1910);
or U2107 (N_2107,N_1827,N_1976);
nor U2108 (N_2108,N_1791,N_1507);
xor U2109 (N_2109,N_1668,N_1685);
and U2110 (N_2110,N_1662,N_1946);
or U2111 (N_2111,N_1635,N_1598);
or U2112 (N_2112,N_1750,N_1617);
xor U2113 (N_2113,N_1514,N_1553);
or U2114 (N_2114,N_1696,N_1688);
and U2115 (N_2115,N_1545,N_1934);
nand U2116 (N_2116,N_1656,N_1649);
nor U2117 (N_2117,N_1659,N_1664);
and U2118 (N_2118,N_1891,N_1596);
nand U2119 (N_2119,N_1643,N_1792);
nand U2120 (N_2120,N_1591,N_1977);
or U2121 (N_2121,N_1959,N_1884);
or U2122 (N_2122,N_1898,N_1546);
nor U2123 (N_2123,N_1867,N_1681);
and U2124 (N_2124,N_1666,N_1665);
and U2125 (N_2125,N_1990,N_1862);
nand U2126 (N_2126,N_1737,N_1824);
nand U2127 (N_2127,N_1777,N_1548);
or U2128 (N_2128,N_1887,N_1932);
and U2129 (N_2129,N_1771,N_1929);
nor U2130 (N_2130,N_1506,N_1706);
or U2131 (N_2131,N_1871,N_1973);
and U2132 (N_2132,N_1689,N_1684);
nor U2133 (N_2133,N_1998,N_1923);
and U2134 (N_2134,N_1547,N_1629);
nor U2135 (N_2135,N_1740,N_1607);
nand U2136 (N_2136,N_1730,N_1573);
and U2137 (N_2137,N_1504,N_1519);
or U2138 (N_2138,N_1729,N_1766);
or U2139 (N_2139,N_1642,N_1961);
nand U2140 (N_2140,N_1585,N_1609);
nor U2141 (N_2141,N_1593,N_1860);
nand U2142 (N_2142,N_1693,N_1634);
or U2143 (N_2143,N_1828,N_1743);
and U2144 (N_2144,N_1955,N_1552);
and U2145 (N_2145,N_1651,N_1639);
nand U2146 (N_2146,N_1720,N_1844);
or U2147 (N_2147,N_1561,N_1525);
or U2148 (N_2148,N_1815,N_1531);
nand U2149 (N_2149,N_1819,N_1667);
nor U2150 (N_2150,N_1537,N_1503);
nand U2151 (N_2151,N_1586,N_1918);
and U2152 (N_2152,N_1583,N_1691);
and U2153 (N_2153,N_1981,N_1906);
xnor U2154 (N_2154,N_1637,N_1584);
nor U2155 (N_2155,N_1807,N_1813);
or U2156 (N_2156,N_1638,N_1877);
nand U2157 (N_2157,N_1817,N_1551);
nor U2158 (N_2158,N_1734,N_1783);
and U2159 (N_2159,N_1746,N_1809);
nand U2160 (N_2160,N_1653,N_1511);
nor U2161 (N_2161,N_1505,N_1763);
and U2162 (N_2162,N_1701,N_1576);
nor U2163 (N_2163,N_1631,N_1597);
or U2164 (N_2164,N_1858,N_1602);
nor U2165 (N_2165,N_1837,N_1935);
nor U2166 (N_2166,N_1578,N_1905);
nor U2167 (N_2167,N_1694,N_1538);
nor U2168 (N_2168,N_1983,N_1996);
xor U2169 (N_2169,N_1810,N_1500);
or U2170 (N_2170,N_1687,N_1909);
or U2171 (N_2171,N_1874,N_1601);
and U2172 (N_2172,N_1778,N_1768);
nor U2173 (N_2173,N_1699,N_1513);
nor U2174 (N_2174,N_1556,N_1868);
and U2175 (N_2175,N_1508,N_1658);
or U2176 (N_2176,N_1702,N_1647);
nor U2177 (N_2177,N_1526,N_1886);
and U2178 (N_2178,N_1795,N_1683);
nor U2179 (N_2179,N_1532,N_1963);
nand U2180 (N_2180,N_1721,N_1882);
and U2181 (N_2181,N_1904,N_1731);
nor U2182 (N_2182,N_1669,N_1690);
nor U2183 (N_2183,N_1518,N_1907);
nand U2184 (N_2184,N_1805,N_1748);
and U2185 (N_2185,N_1957,N_1930);
nand U2186 (N_2186,N_1984,N_1599);
nor U2187 (N_2187,N_1986,N_1962);
nand U2188 (N_2188,N_1577,N_1652);
and U2189 (N_2189,N_1866,N_1821);
or U2190 (N_2190,N_1917,N_1846);
or U2191 (N_2191,N_1757,N_1933);
and U2192 (N_2192,N_1673,N_1856);
and U2193 (N_2193,N_1711,N_1796);
or U2194 (N_2194,N_1632,N_1622);
nor U2195 (N_2195,N_1802,N_1881);
or U2196 (N_2196,N_1675,N_1801);
nand U2197 (N_2197,N_1613,N_1764);
or U2198 (N_2198,N_1999,N_1620);
and U2199 (N_2199,N_1841,N_1921);
and U2200 (N_2200,N_1621,N_1615);
nand U2201 (N_2201,N_1994,N_1785);
nand U2202 (N_2202,N_1735,N_1872);
or U2203 (N_2203,N_1966,N_1566);
nor U2204 (N_2204,N_1895,N_1997);
nand U2205 (N_2205,N_1672,N_1630);
or U2206 (N_2206,N_1587,N_1717);
and U2207 (N_2207,N_1834,N_1549);
or U2208 (N_2208,N_1924,N_1995);
and U2209 (N_2209,N_1517,N_1967);
nand U2210 (N_2210,N_1775,N_1765);
nor U2211 (N_2211,N_1938,N_1985);
and U2212 (N_2212,N_1501,N_1820);
nand U2213 (N_2213,N_1614,N_1864);
nor U2214 (N_2214,N_1722,N_1760);
or U2215 (N_2215,N_1543,N_1861);
or U2216 (N_2216,N_1873,N_1736);
nand U2217 (N_2217,N_1715,N_1949);
or U2218 (N_2218,N_1940,N_1939);
or U2219 (N_2219,N_1812,N_1845);
nor U2220 (N_2220,N_1908,N_1840);
or U2221 (N_2221,N_1951,N_1920);
nand U2222 (N_2222,N_1784,N_1958);
and U2223 (N_2223,N_1619,N_1536);
and U2224 (N_2224,N_1786,N_1892);
or U2225 (N_2225,N_1595,N_1644);
or U2226 (N_2226,N_1604,N_1806);
or U2227 (N_2227,N_1944,N_1878);
and U2228 (N_2228,N_1572,N_1708);
or U2229 (N_2229,N_1742,N_1571);
nor U2230 (N_2230,N_1633,N_1964);
nand U2231 (N_2231,N_1755,N_1980);
nand U2232 (N_2232,N_1554,N_1894);
nand U2233 (N_2233,N_1883,N_1650);
or U2234 (N_2234,N_1794,N_1745);
nand U2235 (N_2235,N_1594,N_1993);
or U2236 (N_2236,N_1521,N_1581);
nor U2237 (N_2237,N_1982,N_1902);
nand U2238 (N_2238,N_1947,N_1606);
nor U2239 (N_2239,N_1863,N_1799);
nand U2240 (N_2240,N_1542,N_1541);
and U2241 (N_2241,N_1767,N_1712);
and U2242 (N_2242,N_1686,N_1832);
and U2243 (N_2243,N_1565,N_1756);
or U2244 (N_2244,N_1941,N_1625);
or U2245 (N_2245,N_1579,N_1590);
or U2246 (N_2246,N_1789,N_1738);
or U2247 (N_2247,N_1830,N_1857);
nand U2248 (N_2248,N_1749,N_1719);
and U2249 (N_2249,N_1512,N_1704);
nor U2250 (N_2250,N_1637,N_1852);
nand U2251 (N_2251,N_1811,N_1865);
nand U2252 (N_2252,N_1940,N_1567);
xnor U2253 (N_2253,N_1553,N_1882);
nor U2254 (N_2254,N_1551,N_1621);
and U2255 (N_2255,N_1513,N_1841);
or U2256 (N_2256,N_1991,N_1752);
and U2257 (N_2257,N_1740,N_1510);
nor U2258 (N_2258,N_1929,N_1930);
nor U2259 (N_2259,N_1844,N_1858);
nor U2260 (N_2260,N_1678,N_1772);
and U2261 (N_2261,N_1839,N_1964);
or U2262 (N_2262,N_1638,N_1721);
nor U2263 (N_2263,N_1911,N_1636);
nand U2264 (N_2264,N_1868,N_1589);
nor U2265 (N_2265,N_1588,N_1837);
xor U2266 (N_2266,N_1573,N_1589);
nor U2267 (N_2267,N_1878,N_1686);
nand U2268 (N_2268,N_1831,N_1994);
nand U2269 (N_2269,N_1832,N_1830);
nand U2270 (N_2270,N_1725,N_1519);
nand U2271 (N_2271,N_1902,N_1702);
nor U2272 (N_2272,N_1661,N_1692);
or U2273 (N_2273,N_1754,N_1992);
and U2274 (N_2274,N_1850,N_1675);
and U2275 (N_2275,N_1639,N_1930);
and U2276 (N_2276,N_1891,N_1711);
nand U2277 (N_2277,N_1536,N_1960);
nand U2278 (N_2278,N_1932,N_1675);
nand U2279 (N_2279,N_1950,N_1963);
and U2280 (N_2280,N_1651,N_1979);
nor U2281 (N_2281,N_1576,N_1792);
and U2282 (N_2282,N_1787,N_1732);
nand U2283 (N_2283,N_1761,N_1655);
nand U2284 (N_2284,N_1700,N_1725);
and U2285 (N_2285,N_1873,N_1613);
and U2286 (N_2286,N_1666,N_1866);
xnor U2287 (N_2287,N_1901,N_1623);
or U2288 (N_2288,N_1655,N_1589);
and U2289 (N_2289,N_1855,N_1737);
nand U2290 (N_2290,N_1574,N_1892);
nand U2291 (N_2291,N_1566,N_1907);
nand U2292 (N_2292,N_1720,N_1886);
and U2293 (N_2293,N_1793,N_1913);
nand U2294 (N_2294,N_1664,N_1808);
nand U2295 (N_2295,N_1652,N_1842);
and U2296 (N_2296,N_1650,N_1683);
nor U2297 (N_2297,N_1834,N_1512);
or U2298 (N_2298,N_1585,N_1893);
and U2299 (N_2299,N_1755,N_1575);
nand U2300 (N_2300,N_1544,N_1921);
and U2301 (N_2301,N_1569,N_1717);
or U2302 (N_2302,N_1800,N_1938);
nor U2303 (N_2303,N_1647,N_1988);
nand U2304 (N_2304,N_1628,N_1839);
nand U2305 (N_2305,N_1733,N_1572);
nor U2306 (N_2306,N_1927,N_1724);
nand U2307 (N_2307,N_1559,N_1745);
nor U2308 (N_2308,N_1882,N_1787);
nor U2309 (N_2309,N_1588,N_1917);
nor U2310 (N_2310,N_1893,N_1713);
or U2311 (N_2311,N_1975,N_1554);
nor U2312 (N_2312,N_1658,N_1503);
nor U2313 (N_2313,N_1598,N_1928);
or U2314 (N_2314,N_1667,N_1827);
and U2315 (N_2315,N_1504,N_1949);
and U2316 (N_2316,N_1564,N_1943);
nand U2317 (N_2317,N_1694,N_1773);
and U2318 (N_2318,N_1646,N_1607);
nand U2319 (N_2319,N_1971,N_1974);
and U2320 (N_2320,N_1504,N_1800);
nor U2321 (N_2321,N_1725,N_1520);
xnor U2322 (N_2322,N_1764,N_1954);
and U2323 (N_2323,N_1925,N_1866);
and U2324 (N_2324,N_1513,N_1521);
nor U2325 (N_2325,N_1907,N_1527);
nand U2326 (N_2326,N_1901,N_1579);
and U2327 (N_2327,N_1539,N_1918);
nor U2328 (N_2328,N_1514,N_1761);
or U2329 (N_2329,N_1533,N_1656);
and U2330 (N_2330,N_1568,N_1599);
nand U2331 (N_2331,N_1996,N_1760);
xor U2332 (N_2332,N_1949,N_1823);
nor U2333 (N_2333,N_1880,N_1833);
xor U2334 (N_2334,N_1713,N_1816);
nor U2335 (N_2335,N_1748,N_1974);
nand U2336 (N_2336,N_1805,N_1634);
nor U2337 (N_2337,N_1708,N_1914);
or U2338 (N_2338,N_1512,N_1522);
and U2339 (N_2339,N_1683,N_1547);
and U2340 (N_2340,N_1987,N_1817);
nor U2341 (N_2341,N_1660,N_1622);
and U2342 (N_2342,N_1841,N_1563);
and U2343 (N_2343,N_1902,N_1749);
or U2344 (N_2344,N_1601,N_1871);
and U2345 (N_2345,N_1507,N_1882);
and U2346 (N_2346,N_1855,N_1986);
or U2347 (N_2347,N_1905,N_1811);
or U2348 (N_2348,N_1794,N_1767);
nor U2349 (N_2349,N_1885,N_1557);
and U2350 (N_2350,N_1966,N_1856);
nand U2351 (N_2351,N_1573,N_1822);
or U2352 (N_2352,N_1983,N_1688);
and U2353 (N_2353,N_1722,N_1792);
and U2354 (N_2354,N_1764,N_1526);
nand U2355 (N_2355,N_1684,N_1997);
and U2356 (N_2356,N_1579,N_1638);
or U2357 (N_2357,N_1798,N_1936);
or U2358 (N_2358,N_1946,N_1777);
or U2359 (N_2359,N_1768,N_1782);
and U2360 (N_2360,N_1733,N_1511);
nor U2361 (N_2361,N_1544,N_1504);
nor U2362 (N_2362,N_1639,N_1678);
nand U2363 (N_2363,N_1505,N_1917);
and U2364 (N_2364,N_1955,N_1644);
nand U2365 (N_2365,N_1773,N_1761);
or U2366 (N_2366,N_1849,N_1624);
and U2367 (N_2367,N_1552,N_1724);
and U2368 (N_2368,N_1980,N_1953);
or U2369 (N_2369,N_1625,N_1934);
or U2370 (N_2370,N_1791,N_1547);
nor U2371 (N_2371,N_1777,N_1663);
nand U2372 (N_2372,N_1881,N_1885);
or U2373 (N_2373,N_1511,N_1806);
nand U2374 (N_2374,N_1543,N_1889);
or U2375 (N_2375,N_1822,N_1985);
or U2376 (N_2376,N_1849,N_1839);
and U2377 (N_2377,N_1830,N_1913);
or U2378 (N_2378,N_1946,N_1781);
or U2379 (N_2379,N_1963,N_1795);
nand U2380 (N_2380,N_1851,N_1988);
nor U2381 (N_2381,N_1828,N_1558);
nand U2382 (N_2382,N_1977,N_1559);
and U2383 (N_2383,N_1932,N_1954);
or U2384 (N_2384,N_1805,N_1771);
or U2385 (N_2385,N_1746,N_1771);
nor U2386 (N_2386,N_1787,N_1842);
or U2387 (N_2387,N_1682,N_1810);
and U2388 (N_2388,N_1507,N_1896);
and U2389 (N_2389,N_1809,N_1982);
or U2390 (N_2390,N_1773,N_1987);
nor U2391 (N_2391,N_1898,N_1755);
nor U2392 (N_2392,N_1589,N_1984);
or U2393 (N_2393,N_1976,N_1564);
nor U2394 (N_2394,N_1608,N_1835);
nor U2395 (N_2395,N_1912,N_1868);
nor U2396 (N_2396,N_1516,N_1897);
nand U2397 (N_2397,N_1715,N_1809);
and U2398 (N_2398,N_1618,N_1797);
nand U2399 (N_2399,N_1963,N_1526);
nor U2400 (N_2400,N_1829,N_1712);
nor U2401 (N_2401,N_1971,N_1778);
nand U2402 (N_2402,N_1750,N_1586);
or U2403 (N_2403,N_1810,N_1506);
and U2404 (N_2404,N_1628,N_1608);
nand U2405 (N_2405,N_1598,N_1946);
nor U2406 (N_2406,N_1841,N_1767);
or U2407 (N_2407,N_1758,N_1701);
or U2408 (N_2408,N_1703,N_1597);
nand U2409 (N_2409,N_1747,N_1938);
nand U2410 (N_2410,N_1637,N_1591);
nand U2411 (N_2411,N_1723,N_1794);
and U2412 (N_2412,N_1960,N_1670);
nor U2413 (N_2413,N_1527,N_1858);
and U2414 (N_2414,N_1523,N_1754);
and U2415 (N_2415,N_1740,N_1614);
and U2416 (N_2416,N_1917,N_1899);
nand U2417 (N_2417,N_1768,N_1890);
nand U2418 (N_2418,N_1615,N_1521);
and U2419 (N_2419,N_1947,N_1788);
and U2420 (N_2420,N_1811,N_1627);
or U2421 (N_2421,N_1956,N_1547);
nor U2422 (N_2422,N_1689,N_1728);
and U2423 (N_2423,N_1979,N_1764);
nand U2424 (N_2424,N_1816,N_1629);
or U2425 (N_2425,N_1777,N_1637);
or U2426 (N_2426,N_1938,N_1674);
nor U2427 (N_2427,N_1559,N_1577);
nand U2428 (N_2428,N_1873,N_1518);
nand U2429 (N_2429,N_1628,N_1558);
and U2430 (N_2430,N_1922,N_1838);
nand U2431 (N_2431,N_1769,N_1921);
or U2432 (N_2432,N_1532,N_1516);
nand U2433 (N_2433,N_1873,N_1807);
nand U2434 (N_2434,N_1528,N_1538);
and U2435 (N_2435,N_1787,N_1623);
nor U2436 (N_2436,N_1853,N_1536);
nand U2437 (N_2437,N_1618,N_1560);
or U2438 (N_2438,N_1669,N_1834);
or U2439 (N_2439,N_1686,N_1643);
and U2440 (N_2440,N_1727,N_1658);
nor U2441 (N_2441,N_1898,N_1525);
and U2442 (N_2442,N_1503,N_1693);
nor U2443 (N_2443,N_1970,N_1922);
or U2444 (N_2444,N_1543,N_1841);
and U2445 (N_2445,N_1605,N_1723);
or U2446 (N_2446,N_1614,N_1881);
and U2447 (N_2447,N_1956,N_1976);
and U2448 (N_2448,N_1505,N_1818);
and U2449 (N_2449,N_1523,N_1904);
nor U2450 (N_2450,N_1847,N_1777);
nand U2451 (N_2451,N_1655,N_1986);
or U2452 (N_2452,N_1788,N_1567);
nor U2453 (N_2453,N_1655,N_1605);
and U2454 (N_2454,N_1909,N_1587);
or U2455 (N_2455,N_1638,N_1923);
nor U2456 (N_2456,N_1509,N_1820);
or U2457 (N_2457,N_1696,N_1868);
or U2458 (N_2458,N_1998,N_1769);
nor U2459 (N_2459,N_1826,N_1950);
or U2460 (N_2460,N_1599,N_1971);
and U2461 (N_2461,N_1676,N_1533);
and U2462 (N_2462,N_1545,N_1548);
or U2463 (N_2463,N_1741,N_1740);
and U2464 (N_2464,N_1903,N_1630);
nor U2465 (N_2465,N_1832,N_1675);
nand U2466 (N_2466,N_1581,N_1738);
and U2467 (N_2467,N_1888,N_1511);
nor U2468 (N_2468,N_1849,N_1633);
and U2469 (N_2469,N_1996,N_1697);
nand U2470 (N_2470,N_1826,N_1883);
and U2471 (N_2471,N_1876,N_1714);
and U2472 (N_2472,N_1893,N_1768);
and U2473 (N_2473,N_1692,N_1946);
and U2474 (N_2474,N_1562,N_1683);
or U2475 (N_2475,N_1942,N_1698);
nand U2476 (N_2476,N_1590,N_1714);
or U2477 (N_2477,N_1996,N_1822);
nor U2478 (N_2478,N_1715,N_1831);
or U2479 (N_2479,N_1958,N_1892);
and U2480 (N_2480,N_1621,N_1584);
nor U2481 (N_2481,N_1620,N_1660);
and U2482 (N_2482,N_1741,N_1753);
nor U2483 (N_2483,N_1914,N_1986);
and U2484 (N_2484,N_1850,N_1824);
or U2485 (N_2485,N_1825,N_1783);
or U2486 (N_2486,N_1600,N_1968);
or U2487 (N_2487,N_1695,N_1969);
nor U2488 (N_2488,N_1976,N_1871);
nor U2489 (N_2489,N_1769,N_1658);
nand U2490 (N_2490,N_1961,N_1999);
nor U2491 (N_2491,N_1879,N_1540);
or U2492 (N_2492,N_1638,N_1646);
nor U2493 (N_2493,N_1975,N_1781);
nor U2494 (N_2494,N_1799,N_1990);
or U2495 (N_2495,N_1857,N_1597);
nor U2496 (N_2496,N_1663,N_1873);
and U2497 (N_2497,N_1526,N_1645);
nor U2498 (N_2498,N_1762,N_1656);
nand U2499 (N_2499,N_1951,N_1637);
nor U2500 (N_2500,N_2357,N_2304);
or U2501 (N_2501,N_2072,N_2036);
or U2502 (N_2502,N_2281,N_2391);
and U2503 (N_2503,N_2053,N_2117);
and U2504 (N_2504,N_2340,N_2412);
and U2505 (N_2505,N_2026,N_2074);
and U2506 (N_2506,N_2187,N_2458);
or U2507 (N_2507,N_2297,N_2170);
nand U2508 (N_2508,N_2077,N_2082);
nand U2509 (N_2509,N_2146,N_2103);
and U2510 (N_2510,N_2477,N_2324);
and U2511 (N_2511,N_2333,N_2048);
nor U2512 (N_2512,N_2464,N_2471);
nor U2513 (N_2513,N_2499,N_2075);
nor U2514 (N_2514,N_2439,N_2445);
and U2515 (N_2515,N_2057,N_2001);
and U2516 (N_2516,N_2293,N_2022);
nor U2517 (N_2517,N_2067,N_2438);
nand U2518 (N_2518,N_2420,N_2396);
and U2519 (N_2519,N_2023,N_2237);
nor U2520 (N_2520,N_2392,N_2215);
nor U2521 (N_2521,N_2459,N_2316);
xnor U2522 (N_2522,N_2260,N_2225);
nand U2523 (N_2523,N_2218,N_2119);
or U2524 (N_2524,N_2470,N_2084);
nand U2525 (N_2525,N_2346,N_2494);
nand U2526 (N_2526,N_2247,N_2351);
or U2527 (N_2527,N_2287,N_2227);
nand U2528 (N_2528,N_2448,N_2130);
or U2529 (N_2529,N_2488,N_2358);
nand U2530 (N_2530,N_2276,N_2212);
nor U2531 (N_2531,N_2106,N_2088);
nor U2532 (N_2532,N_2201,N_2175);
or U2533 (N_2533,N_2167,N_2482);
and U2534 (N_2534,N_2123,N_2475);
and U2535 (N_2535,N_2219,N_2262);
or U2536 (N_2536,N_2043,N_2427);
nor U2537 (N_2537,N_2044,N_2289);
nor U2538 (N_2538,N_2416,N_2213);
nor U2539 (N_2539,N_2014,N_2382);
nand U2540 (N_2540,N_2268,N_2151);
nor U2541 (N_2541,N_2331,N_2006);
nor U2542 (N_2542,N_2010,N_2047);
or U2543 (N_2543,N_2131,N_2385);
and U2544 (N_2544,N_2223,N_2334);
and U2545 (N_2545,N_2198,N_2312);
and U2546 (N_2546,N_2430,N_2078);
or U2547 (N_2547,N_2426,N_2216);
nand U2548 (N_2548,N_2296,N_2256);
and U2549 (N_2549,N_2232,N_2042);
and U2550 (N_2550,N_2073,N_2040);
nor U2551 (N_2551,N_2102,N_2097);
nand U2552 (N_2552,N_2128,N_2265);
and U2553 (N_2553,N_2401,N_2343);
nor U2554 (N_2554,N_2361,N_2313);
and U2555 (N_2555,N_2407,N_2479);
and U2556 (N_2556,N_2381,N_2461);
nor U2557 (N_2557,N_2061,N_2178);
nand U2558 (N_2558,N_2059,N_2244);
nor U2559 (N_2559,N_2372,N_2404);
and U2560 (N_2560,N_2148,N_2166);
or U2561 (N_2561,N_2055,N_2094);
nand U2562 (N_2562,N_2422,N_2089);
nand U2563 (N_2563,N_2165,N_2172);
nor U2564 (N_2564,N_2229,N_2342);
nor U2565 (N_2565,N_2034,N_2311);
nor U2566 (N_2566,N_2046,N_2140);
and U2567 (N_2567,N_2104,N_2373);
nor U2568 (N_2568,N_2176,N_2350);
or U2569 (N_2569,N_2386,N_2124);
or U2570 (N_2570,N_2052,N_2085);
nor U2571 (N_2571,N_2231,N_2419);
and U2572 (N_2572,N_2455,N_2363);
nand U2573 (N_2573,N_2467,N_2193);
or U2574 (N_2574,N_2086,N_2491);
and U2575 (N_2575,N_2217,N_2177);
or U2576 (N_2576,N_2326,N_2028);
nand U2577 (N_2577,N_2428,N_2068);
nor U2578 (N_2578,N_2473,N_2498);
or U2579 (N_2579,N_2259,N_2397);
and U2580 (N_2580,N_2323,N_2279);
or U2581 (N_2581,N_2406,N_2414);
and U2582 (N_2582,N_2384,N_2192);
or U2583 (N_2583,N_2242,N_2465);
nand U2584 (N_2584,N_2100,N_2241);
nand U2585 (N_2585,N_2087,N_2222);
nor U2586 (N_2586,N_2054,N_2236);
nand U2587 (N_2587,N_2025,N_2015);
or U2588 (N_2588,N_2024,N_2147);
xnor U2589 (N_2589,N_2474,N_2338);
xor U2590 (N_2590,N_2332,N_2325);
xor U2591 (N_2591,N_2122,N_2487);
or U2592 (N_2592,N_2433,N_2092);
and U2593 (N_2593,N_2181,N_2317);
nor U2594 (N_2594,N_2429,N_2234);
and U2595 (N_2595,N_2337,N_2377);
nor U2596 (N_2596,N_2090,N_2286);
and U2597 (N_2597,N_2248,N_2450);
nor U2598 (N_2598,N_2139,N_2163);
and U2599 (N_2599,N_2288,N_2127);
or U2600 (N_2600,N_2240,N_2011);
nor U2601 (N_2601,N_2310,N_2275);
or U2602 (N_2602,N_2019,N_2121);
and U2603 (N_2603,N_2496,N_2255);
nor U2604 (N_2604,N_2060,N_2126);
or U2605 (N_2605,N_2210,N_2113);
nor U2606 (N_2606,N_2129,N_2457);
nor U2607 (N_2607,N_2370,N_2033);
or U2608 (N_2608,N_2280,N_2105);
nand U2609 (N_2609,N_2356,N_2327);
nand U2610 (N_2610,N_2294,N_2056);
nor U2611 (N_2611,N_2169,N_2417);
nor U2612 (N_2612,N_2190,N_2452);
and U2613 (N_2613,N_2095,N_2435);
nor U2614 (N_2614,N_2418,N_2463);
or U2615 (N_2615,N_2291,N_2149);
nor U2616 (N_2616,N_2132,N_2460);
nor U2617 (N_2617,N_2205,N_2008);
nor U2618 (N_2618,N_2328,N_2305);
and U2619 (N_2619,N_2045,N_2096);
nor U2620 (N_2620,N_2141,N_2079);
and U2621 (N_2621,N_2408,N_2115);
nand U2622 (N_2622,N_2437,N_2250);
nand U2623 (N_2623,N_2069,N_2409);
xor U2624 (N_2624,N_2017,N_2360);
nand U2625 (N_2625,N_2292,N_2191);
nand U2626 (N_2626,N_2387,N_2451);
or U2627 (N_2627,N_2413,N_2233);
and U2628 (N_2628,N_2206,N_2120);
nand U2629 (N_2629,N_2160,N_2239);
nand U2630 (N_2630,N_2497,N_2395);
nor U2631 (N_2631,N_2335,N_2012);
or U2632 (N_2632,N_2037,N_2180);
or U2633 (N_2633,N_2264,N_2137);
nor U2634 (N_2634,N_2303,N_2065);
and U2635 (N_2635,N_2393,N_2299);
and U2636 (N_2636,N_2134,N_2493);
nor U2637 (N_2637,N_2142,N_2155);
nor U2638 (N_2638,N_2005,N_2195);
or U2639 (N_2639,N_2168,N_2194);
and U2640 (N_2640,N_2329,N_2442);
or U2641 (N_2641,N_2355,N_2004);
nor U2642 (N_2642,N_2150,N_2020);
or U2643 (N_2643,N_2318,N_2110);
xor U2644 (N_2644,N_2041,N_2002);
or U2645 (N_2645,N_2203,N_2462);
nor U2646 (N_2646,N_2380,N_2300);
or U2647 (N_2647,N_2032,N_2083);
or U2648 (N_2648,N_2364,N_2295);
nand U2649 (N_2649,N_2179,N_2099);
or U2650 (N_2650,N_2144,N_2258);
or U2651 (N_2651,N_2484,N_2207);
nor U2652 (N_2652,N_2249,N_2270);
nand U2653 (N_2653,N_2447,N_2376);
and U2654 (N_2654,N_2449,N_2421);
and U2655 (N_2655,N_2245,N_2423);
nor U2656 (N_2656,N_2388,N_2378);
and U2657 (N_2657,N_2221,N_2341);
nor U2658 (N_2658,N_2348,N_2336);
or U2659 (N_2659,N_2183,N_2320);
and U2660 (N_2660,N_2220,N_2080);
and U2661 (N_2661,N_2490,N_2368);
nor U2662 (N_2662,N_2064,N_2347);
or U2663 (N_2663,N_2436,N_2306);
and U2664 (N_2664,N_2186,N_2267);
or U2665 (N_2665,N_2302,N_2039);
nand U2666 (N_2666,N_2495,N_2456);
and U2667 (N_2667,N_2062,N_2230);
nand U2668 (N_2668,N_2301,N_2290);
nand U2669 (N_2669,N_2399,N_2481);
and U2670 (N_2670,N_2352,N_2261);
or U2671 (N_2671,N_2107,N_2277);
nand U2672 (N_2672,N_2415,N_2283);
or U2673 (N_2673,N_2112,N_2367);
nand U2674 (N_2674,N_2189,N_2050);
nand U2675 (N_2675,N_2405,N_2272);
or U2676 (N_2676,N_2307,N_2029);
and U2677 (N_2677,N_2111,N_2274);
nor U2678 (N_2678,N_2164,N_2101);
or U2679 (N_2679,N_2365,N_2228);
and U2680 (N_2680,N_2454,N_2108);
nand U2681 (N_2681,N_2251,N_2486);
nor U2682 (N_2682,N_2308,N_2093);
and U2683 (N_2683,N_2330,N_2021);
nand U2684 (N_2684,N_2441,N_2444);
nor U2685 (N_2685,N_2153,N_2161);
nand U2686 (N_2686,N_2271,N_2066);
nor U2687 (N_2687,N_2133,N_2489);
nor U2688 (N_2688,N_2383,N_2480);
or U2689 (N_2689,N_2389,N_2469);
nand U2690 (N_2690,N_2202,N_2063);
and U2691 (N_2691,N_2252,N_2253);
and U2692 (N_2692,N_2362,N_2070);
and U2693 (N_2693,N_2478,N_2214);
nand U2694 (N_2694,N_2114,N_2483);
nor U2695 (N_2695,N_2158,N_2403);
or U2696 (N_2696,N_2109,N_2098);
and U2697 (N_2697,N_2254,N_2321);
and U2698 (N_2698,N_2266,N_2453);
or U2699 (N_2699,N_2319,N_2200);
nor U2700 (N_2700,N_2468,N_2273);
and U2701 (N_2701,N_2199,N_2013);
or U2702 (N_2702,N_2349,N_2138);
nand U2703 (N_2703,N_2027,N_2263);
or U2704 (N_2704,N_2411,N_2071);
and U2705 (N_2705,N_2058,N_2196);
nor U2706 (N_2706,N_2322,N_2173);
and U2707 (N_2707,N_2353,N_2038);
or U2708 (N_2708,N_2211,N_2434);
or U2709 (N_2709,N_2007,N_2440);
or U2710 (N_2710,N_2284,N_2235);
nor U2711 (N_2711,N_2081,N_2091);
and U2712 (N_2712,N_2182,N_2339);
or U2713 (N_2713,N_2354,N_2345);
nand U2714 (N_2714,N_2400,N_2366);
nand U2715 (N_2715,N_2224,N_2174);
nor U2716 (N_2716,N_2118,N_2485);
nand U2717 (N_2717,N_2076,N_2156);
nor U2718 (N_2718,N_2162,N_2315);
and U2719 (N_2719,N_2136,N_2238);
nor U2720 (N_2720,N_2432,N_2371);
nand U2721 (N_2721,N_2185,N_2125);
or U2722 (N_2722,N_2425,N_2446);
or U2723 (N_2723,N_2269,N_2000);
nor U2724 (N_2724,N_2209,N_2009);
or U2725 (N_2725,N_2152,N_2143);
or U2726 (N_2726,N_2476,N_2197);
nand U2727 (N_2727,N_2243,N_2154);
and U2728 (N_2728,N_2379,N_2204);
and U2729 (N_2729,N_2116,N_2157);
nand U2730 (N_2730,N_2018,N_2359);
nand U2731 (N_2731,N_2035,N_2375);
and U2732 (N_2732,N_2282,N_2184);
nand U2733 (N_2733,N_2171,N_2051);
or U2734 (N_2734,N_2208,N_2145);
or U2735 (N_2735,N_2031,N_2402);
or U2736 (N_2736,N_2003,N_2369);
and U2737 (N_2737,N_2285,N_2472);
or U2738 (N_2738,N_2410,N_2188);
nand U2739 (N_2739,N_2298,N_2246);
and U2740 (N_2740,N_2398,N_2394);
nand U2741 (N_2741,N_2257,N_2466);
and U2742 (N_2742,N_2492,N_2226);
and U2743 (N_2743,N_2159,N_2016);
and U2744 (N_2744,N_2278,N_2314);
and U2745 (N_2745,N_2424,N_2344);
and U2746 (N_2746,N_2309,N_2030);
nor U2747 (N_2747,N_2431,N_2390);
nor U2748 (N_2748,N_2049,N_2443);
nand U2749 (N_2749,N_2374,N_2135);
or U2750 (N_2750,N_2405,N_2302);
and U2751 (N_2751,N_2298,N_2305);
nor U2752 (N_2752,N_2428,N_2211);
and U2753 (N_2753,N_2282,N_2022);
nor U2754 (N_2754,N_2164,N_2017);
or U2755 (N_2755,N_2481,N_2110);
nand U2756 (N_2756,N_2002,N_2095);
nor U2757 (N_2757,N_2119,N_2313);
nand U2758 (N_2758,N_2155,N_2169);
and U2759 (N_2759,N_2287,N_2331);
nor U2760 (N_2760,N_2260,N_2097);
or U2761 (N_2761,N_2433,N_2087);
or U2762 (N_2762,N_2331,N_2278);
nand U2763 (N_2763,N_2082,N_2147);
nor U2764 (N_2764,N_2491,N_2378);
nand U2765 (N_2765,N_2225,N_2197);
nand U2766 (N_2766,N_2213,N_2488);
nor U2767 (N_2767,N_2112,N_2375);
xnor U2768 (N_2768,N_2257,N_2175);
nor U2769 (N_2769,N_2045,N_2093);
or U2770 (N_2770,N_2208,N_2418);
or U2771 (N_2771,N_2039,N_2400);
nand U2772 (N_2772,N_2182,N_2038);
and U2773 (N_2773,N_2343,N_2236);
and U2774 (N_2774,N_2000,N_2186);
and U2775 (N_2775,N_2015,N_2315);
nor U2776 (N_2776,N_2056,N_2415);
or U2777 (N_2777,N_2164,N_2130);
nand U2778 (N_2778,N_2048,N_2042);
nand U2779 (N_2779,N_2225,N_2282);
nor U2780 (N_2780,N_2326,N_2128);
or U2781 (N_2781,N_2276,N_2493);
and U2782 (N_2782,N_2233,N_2254);
nand U2783 (N_2783,N_2293,N_2370);
nor U2784 (N_2784,N_2298,N_2363);
and U2785 (N_2785,N_2142,N_2011);
nand U2786 (N_2786,N_2465,N_2442);
nand U2787 (N_2787,N_2139,N_2332);
nand U2788 (N_2788,N_2048,N_2278);
nor U2789 (N_2789,N_2000,N_2104);
and U2790 (N_2790,N_2271,N_2498);
or U2791 (N_2791,N_2154,N_2261);
nand U2792 (N_2792,N_2196,N_2145);
or U2793 (N_2793,N_2120,N_2158);
and U2794 (N_2794,N_2012,N_2039);
or U2795 (N_2795,N_2438,N_2012);
nor U2796 (N_2796,N_2460,N_2424);
nand U2797 (N_2797,N_2052,N_2350);
nor U2798 (N_2798,N_2202,N_2194);
or U2799 (N_2799,N_2392,N_2066);
and U2800 (N_2800,N_2484,N_2274);
nand U2801 (N_2801,N_2019,N_2310);
or U2802 (N_2802,N_2469,N_2382);
and U2803 (N_2803,N_2236,N_2018);
and U2804 (N_2804,N_2368,N_2459);
nand U2805 (N_2805,N_2373,N_2314);
nor U2806 (N_2806,N_2008,N_2053);
xnor U2807 (N_2807,N_2386,N_2068);
or U2808 (N_2808,N_2480,N_2065);
or U2809 (N_2809,N_2042,N_2073);
and U2810 (N_2810,N_2336,N_2118);
and U2811 (N_2811,N_2095,N_2139);
nand U2812 (N_2812,N_2241,N_2395);
or U2813 (N_2813,N_2321,N_2381);
nor U2814 (N_2814,N_2056,N_2060);
nand U2815 (N_2815,N_2386,N_2127);
or U2816 (N_2816,N_2263,N_2069);
nor U2817 (N_2817,N_2360,N_2356);
nand U2818 (N_2818,N_2275,N_2473);
and U2819 (N_2819,N_2471,N_2011);
or U2820 (N_2820,N_2343,N_2135);
nor U2821 (N_2821,N_2040,N_2113);
and U2822 (N_2822,N_2340,N_2255);
nor U2823 (N_2823,N_2471,N_2103);
or U2824 (N_2824,N_2390,N_2241);
nand U2825 (N_2825,N_2446,N_2272);
nor U2826 (N_2826,N_2319,N_2209);
nor U2827 (N_2827,N_2088,N_2162);
or U2828 (N_2828,N_2481,N_2409);
and U2829 (N_2829,N_2141,N_2155);
nor U2830 (N_2830,N_2406,N_2162);
and U2831 (N_2831,N_2143,N_2083);
nor U2832 (N_2832,N_2144,N_2266);
or U2833 (N_2833,N_2310,N_2346);
and U2834 (N_2834,N_2018,N_2174);
and U2835 (N_2835,N_2021,N_2273);
and U2836 (N_2836,N_2359,N_2232);
nand U2837 (N_2837,N_2433,N_2346);
nor U2838 (N_2838,N_2358,N_2477);
or U2839 (N_2839,N_2462,N_2199);
nor U2840 (N_2840,N_2031,N_2276);
nand U2841 (N_2841,N_2270,N_2221);
and U2842 (N_2842,N_2426,N_2344);
or U2843 (N_2843,N_2275,N_2351);
nand U2844 (N_2844,N_2381,N_2100);
nor U2845 (N_2845,N_2083,N_2240);
nor U2846 (N_2846,N_2417,N_2059);
nand U2847 (N_2847,N_2343,N_2092);
and U2848 (N_2848,N_2244,N_2100);
and U2849 (N_2849,N_2365,N_2046);
nor U2850 (N_2850,N_2343,N_2263);
and U2851 (N_2851,N_2454,N_2066);
nand U2852 (N_2852,N_2309,N_2266);
nor U2853 (N_2853,N_2460,N_2018);
nand U2854 (N_2854,N_2100,N_2354);
and U2855 (N_2855,N_2318,N_2157);
nor U2856 (N_2856,N_2112,N_2077);
or U2857 (N_2857,N_2134,N_2314);
nand U2858 (N_2858,N_2422,N_2109);
or U2859 (N_2859,N_2195,N_2164);
nand U2860 (N_2860,N_2138,N_2331);
nor U2861 (N_2861,N_2426,N_2383);
or U2862 (N_2862,N_2094,N_2243);
nand U2863 (N_2863,N_2253,N_2369);
or U2864 (N_2864,N_2107,N_2214);
xnor U2865 (N_2865,N_2161,N_2309);
nand U2866 (N_2866,N_2101,N_2068);
xnor U2867 (N_2867,N_2010,N_2098);
nand U2868 (N_2868,N_2050,N_2324);
nor U2869 (N_2869,N_2084,N_2062);
and U2870 (N_2870,N_2290,N_2373);
or U2871 (N_2871,N_2187,N_2246);
nor U2872 (N_2872,N_2207,N_2440);
nand U2873 (N_2873,N_2257,N_2436);
nand U2874 (N_2874,N_2115,N_2421);
nand U2875 (N_2875,N_2191,N_2300);
and U2876 (N_2876,N_2344,N_2321);
and U2877 (N_2877,N_2499,N_2406);
nand U2878 (N_2878,N_2362,N_2294);
nor U2879 (N_2879,N_2124,N_2281);
and U2880 (N_2880,N_2183,N_2233);
or U2881 (N_2881,N_2056,N_2004);
nand U2882 (N_2882,N_2288,N_2400);
nand U2883 (N_2883,N_2313,N_2011);
nand U2884 (N_2884,N_2034,N_2426);
or U2885 (N_2885,N_2461,N_2392);
nor U2886 (N_2886,N_2447,N_2333);
nand U2887 (N_2887,N_2394,N_2355);
and U2888 (N_2888,N_2478,N_2459);
nand U2889 (N_2889,N_2171,N_2227);
or U2890 (N_2890,N_2055,N_2386);
nor U2891 (N_2891,N_2023,N_2296);
nand U2892 (N_2892,N_2059,N_2168);
nand U2893 (N_2893,N_2181,N_2280);
and U2894 (N_2894,N_2437,N_2148);
nand U2895 (N_2895,N_2445,N_2038);
nand U2896 (N_2896,N_2015,N_2468);
and U2897 (N_2897,N_2233,N_2165);
and U2898 (N_2898,N_2314,N_2081);
or U2899 (N_2899,N_2202,N_2016);
nor U2900 (N_2900,N_2286,N_2089);
nand U2901 (N_2901,N_2086,N_2435);
nand U2902 (N_2902,N_2360,N_2197);
and U2903 (N_2903,N_2499,N_2032);
nand U2904 (N_2904,N_2431,N_2334);
xor U2905 (N_2905,N_2483,N_2084);
xor U2906 (N_2906,N_2380,N_2098);
nor U2907 (N_2907,N_2398,N_2043);
and U2908 (N_2908,N_2033,N_2170);
and U2909 (N_2909,N_2354,N_2168);
nor U2910 (N_2910,N_2355,N_2381);
nor U2911 (N_2911,N_2220,N_2067);
nor U2912 (N_2912,N_2380,N_2148);
or U2913 (N_2913,N_2082,N_2408);
nor U2914 (N_2914,N_2104,N_2316);
nand U2915 (N_2915,N_2386,N_2322);
nand U2916 (N_2916,N_2463,N_2445);
or U2917 (N_2917,N_2460,N_2280);
nand U2918 (N_2918,N_2269,N_2402);
and U2919 (N_2919,N_2187,N_2062);
nor U2920 (N_2920,N_2475,N_2109);
and U2921 (N_2921,N_2087,N_2324);
and U2922 (N_2922,N_2025,N_2246);
nor U2923 (N_2923,N_2029,N_2233);
nand U2924 (N_2924,N_2217,N_2036);
and U2925 (N_2925,N_2308,N_2118);
nand U2926 (N_2926,N_2029,N_2259);
nand U2927 (N_2927,N_2403,N_2255);
and U2928 (N_2928,N_2103,N_2229);
nand U2929 (N_2929,N_2021,N_2391);
or U2930 (N_2930,N_2291,N_2359);
nor U2931 (N_2931,N_2377,N_2036);
and U2932 (N_2932,N_2328,N_2213);
or U2933 (N_2933,N_2363,N_2459);
nand U2934 (N_2934,N_2356,N_2487);
or U2935 (N_2935,N_2383,N_2301);
or U2936 (N_2936,N_2248,N_2228);
nand U2937 (N_2937,N_2260,N_2470);
nand U2938 (N_2938,N_2101,N_2096);
nand U2939 (N_2939,N_2257,N_2479);
and U2940 (N_2940,N_2272,N_2132);
nor U2941 (N_2941,N_2294,N_2365);
and U2942 (N_2942,N_2340,N_2383);
nand U2943 (N_2943,N_2140,N_2148);
nand U2944 (N_2944,N_2472,N_2398);
nor U2945 (N_2945,N_2158,N_2065);
or U2946 (N_2946,N_2394,N_2056);
or U2947 (N_2947,N_2263,N_2021);
or U2948 (N_2948,N_2189,N_2479);
nor U2949 (N_2949,N_2083,N_2131);
and U2950 (N_2950,N_2114,N_2047);
nand U2951 (N_2951,N_2485,N_2228);
and U2952 (N_2952,N_2483,N_2290);
and U2953 (N_2953,N_2442,N_2077);
nor U2954 (N_2954,N_2248,N_2100);
or U2955 (N_2955,N_2049,N_2342);
nor U2956 (N_2956,N_2015,N_2289);
and U2957 (N_2957,N_2168,N_2340);
nand U2958 (N_2958,N_2283,N_2289);
nand U2959 (N_2959,N_2250,N_2267);
or U2960 (N_2960,N_2336,N_2177);
nor U2961 (N_2961,N_2336,N_2491);
nand U2962 (N_2962,N_2227,N_2404);
nor U2963 (N_2963,N_2481,N_2176);
nor U2964 (N_2964,N_2262,N_2243);
or U2965 (N_2965,N_2324,N_2146);
or U2966 (N_2966,N_2420,N_2145);
nand U2967 (N_2967,N_2224,N_2023);
and U2968 (N_2968,N_2326,N_2237);
or U2969 (N_2969,N_2068,N_2413);
nor U2970 (N_2970,N_2439,N_2384);
nand U2971 (N_2971,N_2395,N_2318);
or U2972 (N_2972,N_2107,N_2406);
nor U2973 (N_2973,N_2259,N_2024);
or U2974 (N_2974,N_2247,N_2461);
or U2975 (N_2975,N_2404,N_2439);
nand U2976 (N_2976,N_2097,N_2306);
and U2977 (N_2977,N_2157,N_2357);
nor U2978 (N_2978,N_2009,N_2019);
and U2979 (N_2979,N_2154,N_2457);
or U2980 (N_2980,N_2490,N_2019);
and U2981 (N_2981,N_2465,N_2405);
or U2982 (N_2982,N_2185,N_2090);
nor U2983 (N_2983,N_2361,N_2315);
or U2984 (N_2984,N_2407,N_2317);
or U2985 (N_2985,N_2347,N_2239);
and U2986 (N_2986,N_2413,N_2076);
nand U2987 (N_2987,N_2266,N_2499);
and U2988 (N_2988,N_2052,N_2157);
nand U2989 (N_2989,N_2491,N_2196);
or U2990 (N_2990,N_2132,N_2493);
or U2991 (N_2991,N_2244,N_2161);
and U2992 (N_2992,N_2073,N_2229);
and U2993 (N_2993,N_2446,N_2352);
or U2994 (N_2994,N_2135,N_2290);
nand U2995 (N_2995,N_2131,N_2216);
nand U2996 (N_2996,N_2258,N_2055);
or U2997 (N_2997,N_2221,N_2098);
or U2998 (N_2998,N_2414,N_2195);
nand U2999 (N_2999,N_2393,N_2270);
nand U3000 (N_3000,N_2565,N_2822);
and U3001 (N_3001,N_2848,N_2793);
and U3002 (N_3002,N_2997,N_2801);
nand U3003 (N_3003,N_2641,N_2949);
nor U3004 (N_3004,N_2752,N_2869);
and U3005 (N_3005,N_2998,N_2714);
and U3006 (N_3006,N_2543,N_2847);
and U3007 (N_3007,N_2651,N_2754);
nor U3008 (N_3008,N_2784,N_2776);
nor U3009 (N_3009,N_2757,N_2534);
nor U3010 (N_3010,N_2571,N_2771);
and U3011 (N_3011,N_2620,N_2772);
and U3012 (N_3012,N_2704,N_2599);
and U3013 (N_3013,N_2823,N_2512);
nor U3014 (N_3014,N_2928,N_2549);
nor U3015 (N_3015,N_2900,N_2531);
nand U3016 (N_3016,N_2934,N_2764);
or U3017 (N_3017,N_2581,N_2744);
nor U3018 (N_3018,N_2552,N_2702);
and U3019 (N_3019,N_2777,N_2708);
or U3020 (N_3020,N_2551,N_2547);
and U3021 (N_3021,N_2758,N_2877);
nor U3022 (N_3022,N_2642,N_2890);
and U3023 (N_3023,N_2671,N_2950);
or U3024 (N_3024,N_2954,N_2863);
and U3025 (N_3025,N_2600,N_2661);
or U3026 (N_3026,N_2929,N_2682);
or U3027 (N_3027,N_2861,N_2835);
nor U3028 (N_3028,N_2878,N_2886);
nor U3029 (N_3029,N_2666,N_2767);
nor U3030 (N_3030,N_2616,N_2507);
nor U3031 (N_3031,N_2819,N_2518);
and U3032 (N_3032,N_2660,N_2537);
nand U3033 (N_3033,N_2969,N_2530);
nand U3034 (N_3034,N_2649,N_2559);
nor U3035 (N_3035,N_2967,N_2840);
and U3036 (N_3036,N_2773,N_2629);
and U3037 (N_3037,N_2883,N_2726);
and U3038 (N_3038,N_2546,N_2927);
or U3039 (N_3039,N_2670,N_2946);
or U3040 (N_3040,N_2536,N_2668);
nand U3041 (N_3041,N_2609,N_2992);
and U3042 (N_3042,N_2747,N_2582);
nor U3043 (N_3043,N_2817,N_2523);
nor U3044 (N_3044,N_2831,N_2836);
nor U3045 (N_3045,N_2681,N_2911);
and U3046 (N_3046,N_2880,N_2741);
nor U3047 (N_3047,N_2694,N_2889);
nand U3048 (N_3048,N_2514,N_2919);
or U3049 (N_3049,N_2669,N_2575);
and U3050 (N_3050,N_2795,N_2680);
and U3051 (N_3051,N_2931,N_2685);
and U3052 (N_3052,N_2984,N_2623);
nand U3053 (N_3053,N_2983,N_2516);
nand U3054 (N_3054,N_2809,N_2569);
nand U3055 (N_3055,N_2750,N_2820);
nand U3056 (N_3056,N_2522,N_2985);
nor U3057 (N_3057,N_2715,N_2743);
or U3058 (N_3058,N_2903,N_2686);
or U3059 (N_3059,N_2664,N_2994);
and U3060 (N_3060,N_2789,N_2775);
and U3061 (N_3061,N_2925,N_2755);
nand U3062 (N_3062,N_2828,N_2563);
nand U3063 (N_3063,N_2683,N_2566);
and U3064 (N_3064,N_2924,N_2792);
nand U3065 (N_3065,N_2893,N_2947);
or U3066 (N_3066,N_2562,N_2875);
and U3067 (N_3067,N_2633,N_2802);
and U3068 (N_3068,N_2503,N_2794);
nand U3069 (N_3069,N_2699,N_2850);
nand U3070 (N_3070,N_2937,N_2916);
or U3071 (N_3071,N_2738,N_2711);
nor U3072 (N_3072,N_2885,N_2787);
nand U3073 (N_3073,N_2524,N_2874);
nor U3074 (N_3074,N_2851,N_2548);
nand U3075 (N_3075,N_2695,N_2896);
and U3076 (N_3076,N_2904,N_2596);
and U3077 (N_3077,N_2662,N_2996);
or U3078 (N_3078,N_2979,N_2965);
or U3079 (N_3079,N_2865,N_2712);
nand U3080 (N_3080,N_2605,N_2827);
nand U3081 (N_3081,N_2585,N_2864);
nand U3082 (N_3082,N_2707,N_2756);
nor U3083 (N_3083,N_2923,N_2815);
or U3084 (N_3084,N_2703,N_2824);
nor U3085 (N_3085,N_2811,N_2867);
nor U3086 (N_3086,N_2652,N_2688);
nor U3087 (N_3087,N_2615,N_2719);
and U3088 (N_3088,N_2674,N_2844);
and U3089 (N_3089,N_2834,N_2990);
and U3090 (N_3090,N_2779,N_2991);
and U3091 (N_3091,N_2648,N_2879);
nor U3092 (N_3092,N_2959,N_2635);
nor U3093 (N_3093,N_2604,N_2574);
or U3094 (N_3094,N_2630,N_2568);
nor U3095 (N_3095,N_2625,N_2943);
or U3096 (N_3096,N_2607,N_2636);
nor U3097 (N_3097,N_2706,N_2951);
or U3098 (N_3098,N_2942,N_2519);
or U3099 (N_3099,N_2818,N_2614);
or U3100 (N_3100,N_2945,N_2515);
or U3101 (N_3101,N_2717,N_2800);
or U3102 (N_3102,N_2888,N_2533);
nand U3103 (N_3103,N_2583,N_2940);
and U3104 (N_3104,N_2645,N_2876);
nor U3105 (N_3105,N_2973,N_2899);
nand U3106 (N_3106,N_2692,N_2689);
nor U3107 (N_3107,N_2980,N_2906);
and U3108 (N_3108,N_2866,N_2696);
nor U3109 (N_3109,N_2611,N_2731);
or U3110 (N_3110,N_2729,N_2560);
nand U3111 (N_3111,N_2999,N_2912);
or U3112 (N_3112,N_2976,N_2956);
nor U3113 (N_3113,N_2721,N_2561);
and U3114 (N_3114,N_2868,N_2843);
and U3115 (N_3115,N_2860,N_2753);
and U3116 (N_3116,N_2626,N_2957);
nand U3117 (N_3117,N_2962,N_2908);
nand U3118 (N_3118,N_2513,N_2915);
xor U3119 (N_3119,N_2790,N_2952);
or U3120 (N_3120,N_2541,N_2799);
nor U3121 (N_3121,N_2770,N_2926);
nor U3122 (N_3122,N_2610,N_2986);
or U3123 (N_3123,N_2971,N_2505);
and U3124 (N_3124,N_2544,N_2780);
nand U3125 (N_3125,N_2909,N_2580);
or U3126 (N_3126,N_2601,N_2921);
and U3127 (N_3127,N_2791,N_2778);
or U3128 (N_3128,N_2589,N_2948);
and U3129 (N_3129,N_2989,N_2760);
nor U3130 (N_3130,N_2595,N_2593);
nor U3131 (N_3131,N_2987,N_2691);
or U3132 (N_3132,N_2830,N_2873);
nand U3133 (N_3133,N_2677,N_2558);
nand U3134 (N_3134,N_2759,N_2638);
or U3135 (N_3135,N_2936,N_2578);
or U3136 (N_3136,N_2881,N_2665);
or U3137 (N_3137,N_2631,N_2597);
or U3138 (N_3138,N_2734,N_2720);
nand U3139 (N_3139,N_2826,N_2841);
nand U3140 (N_3140,N_2639,N_2862);
nor U3141 (N_3141,N_2853,N_2540);
nor U3142 (N_3142,N_2837,N_2930);
and U3143 (N_3143,N_2700,N_2748);
nand U3144 (N_3144,N_2829,N_2806);
and U3145 (N_3145,N_2693,N_2598);
nand U3146 (N_3146,N_2849,N_2722);
nand U3147 (N_3147,N_2511,N_2803);
or U3148 (N_3148,N_2872,N_2846);
nand U3149 (N_3149,N_2632,N_2527);
and U3150 (N_3150,N_2643,N_2687);
nor U3151 (N_3151,N_2590,N_2564);
or U3152 (N_3152,N_2594,N_2870);
nor U3153 (N_3153,N_2892,N_2856);
or U3154 (N_3154,N_2619,N_2766);
nor U3155 (N_3155,N_2958,N_2894);
and U3156 (N_3156,N_2628,N_2812);
and U3157 (N_3157,N_2988,N_2902);
and U3158 (N_3158,N_2647,N_2679);
nor U3159 (N_3159,N_2917,N_2898);
nand U3160 (N_3160,N_2586,N_2550);
nor U3161 (N_3161,N_2728,N_2602);
nor U3162 (N_3162,N_2640,N_2520);
and U3163 (N_3163,N_2814,N_2672);
or U3164 (N_3164,N_2521,N_2701);
nand U3165 (N_3165,N_2705,N_2763);
nor U3166 (N_3166,N_2781,N_2933);
nand U3167 (N_3167,N_2939,N_2858);
or U3168 (N_3168,N_2821,N_2656);
nand U3169 (N_3169,N_2972,N_2637);
nor U3170 (N_3170,N_2981,N_2745);
or U3171 (N_3171,N_2723,N_2974);
nand U3172 (N_3172,N_2798,N_2941);
xor U3173 (N_3173,N_2532,N_2622);
or U3174 (N_3174,N_2740,N_2657);
nand U3175 (N_3175,N_2554,N_2910);
or U3176 (N_3176,N_2650,N_2749);
and U3177 (N_3177,N_2684,N_2960);
nand U3178 (N_3178,N_2724,N_2716);
and U3179 (N_3179,N_2774,N_2556);
and U3180 (N_3180,N_2739,N_2993);
and U3181 (N_3181,N_2634,N_2832);
or U3182 (N_3182,N_2810,N_2577);
or U3183 (N_3183,N_2592,N_2653);
or U3184 (N_3184,N_2667,N_2966);
or U3185 (N_3185,N_2735,N_2587);
or U3186 (N_3186,N_2833,N_2504);
nand U3187 (N_3187,N_2528,N_2797);
or U3188 (N_3188,N_2567,N_2783);
nor U3189 (N_3189,N_2839,N_2761);
and U3190 (N_3190,N_2553,N_2570);
nand U3191 (N_3191,N_2808,N_2730);
and U3192 (N_3192,N_2742,N_2857);
or U3193 (N_3193,N_2539,N_2606);
and U3194 (N_3194,N_2975,N_2573);
nand U3195 (N_3195,N_2901,N_2842);
nand U3196 (N_3196,N_2955,N_2502);
and U3197 (N_3197,N_2804,N_2572);
xor U3198 (N_3198,N_2961,N_2644);
nand U3199 (N_3199,N_2506,N_2621);
or U3200 (N_3200,N_2782,N_2646);
nand U3201 (N_3201,N_2768,N_2659);
nand U3202 (N_3202,N_2796,N_2588);
nand U3203 (N_3203,N_2555,N_2557);
nor U3204 (N_3204,N_2525,N_2995);
and U3205 (N_3205,N_2690,N_2938);
nor U3206 (N_3206,N_2963,N_2746);
or U3207 (N_3207,N_2663,N_2913);
nand U3208 (N_3208,N_2612,N_2895);
and U3209 (N_3209,N_2538,N_2732);
or U3210 (N_3210,N_2788,N_2769);
or U3211 (N_3211,N_2968,N_2500);
nor U3212 (N_3212,N_2654,N_2807);
and U3213 (N_3213,N_2545,N_2918);
nor U3214 (N_3214,N_2579,N_2517);
and U3215 (N_3215,N_2964,N_2737);
or U3216 (N_3216,N_2655,N_2709);
and U3217 (N_3217,N_2508,N_2982);
nand U3218 (N_3218,N_2675,N_2953);
nor U3219 (N_3219,N_2627,N_2618);
nand U3220 (N_3220,N_2658,N_2914);
nor U3221 (N_3221,N_2977,N_2584);
nor U3222 (N_3222,N_2617,N_2576);
nand U3223 (N_3223,N_2535,N_2920);
nand U3224 (N_3224,N_2624,N_2932);
or U3225 (N_3225,N_2907,N_2786);
or U3226 (N_3226,N_2736,N_2825);
or U3227 (N_3227,N_2813,N_2762);
nand U3228 (N_3228,N_2854,N_2608);
and U3229 (N_3229,N_2922,N_2526);
nor U3230 (N_3230,N_2698,N_2852);
nor U3231 (N_3231,N_2978,N_2887);
and U3232 (N_3232,N_2529,N_2805);
and U3233 (N_3233,N_2751,N_2501);
and U3234 (N_3234,N_2871,N_2713);
nor U3235 (N_3235,N_2816,N_2542);
nand U3236 (N_3236,N_2678,N_2855);
or U3237 (N_3237,N_2725,N_2676);
or U3238 (N_3238,N_2733,N_2510);
or U3239 (N_3239,N_2884,N_2591);
and U3240 (N_3240,N_2897,N_2944);
nor U3241 (N_3241,N_2882,N_2838);
or U3242 (N_3242,N_2613,N_2935);
or U3243 (N_3243,N_2970,N_2710);
or U3244 (N_3244,N_2509,N_2765);
and U3245 (N_3245,N_2603,N_2785);
and U3246 (N_3246,N_2891,N_2718);
or U3247 (N_3247,N_2859,N_2845);
or U3248 (N_3248,N_2697,N_2905);
and U3249 (N_3249,N_2673,N_2727);
or U3250 (N_3250,N_2835,N_2518);
and U3251 (N_3251,N_2847,N_2674);
nand U3252 (N_3252,N_2721,N_2710);
nor U3253 (N_3253,N_2859,N_2664);
or U3254 (N_3254,N_2863,N_2838);
nand U3255 (N_3255,N_2920,N_2562);
nor U3256 (N_3256,N_2940,N_2732);
and U3257 (N_3257,N_2603,N_2823);
or U3258 (N_3258,N_2538,N_2524);
nand U3259 (N_3259,N_2502,N_2543);
or U3260 (N_3260,N_2662,N_2670);
nand U3261 (N_3261,N_2690,N_2860);
nand U3262 (N_3262,N_2557,N_2903);
and U3263 (N_3263,N_2582,N_2763);
and U3264 (N_3264,N_2516,N_2972);
or U3265 (N_3265,N_2642,N_2507);
nor U3266 (N_3266,N_2900,N_2621);
or U3267 (N_3267,N_2681,N_2710);
nor U3268 (N_3268,N_2670,N_2895);
and U3269 (N_3269,N_2945,N_2976);
nand U3270 (N_3270,N_2756,N_2680);
or U3271 (N_3271,N_2591,N_2628);
and U3272 (N_3272,N_2918,N_2576);
and U3273 (N_3273,N_2647,N_2546);
nand U3274 (N_3274,N_2670,N_2921);
or U3275 (N_3275,N_2565,N_2986);
and U3276 (N_3276,N_2660,N_2812);
nor U3277 (N_3277,N_2742,N_2899);
nor U3278 (N_3278,N_2582,N_2899);
or U3279 (N_3279,N_2823,N_2629);
nand U3280 (N_3280,N_2777,N_2624);
or U3281 (N_3281,N_2824,N_2541);
or U3282 (N_3282,N_2759,N_2670);
nand U3283 (N_3283,N_2868,N_2707);
nand U3284 (N_3284,N_2672,N_2658);
nor U3285 (N_3285,N_2631,N_2876);
nor U3286 (N_3286,N_2561,N_2667);
nor U3287 (N_3287,N_2586,N_2886);
and U3288 (N_3288,N_2539,N_2615);
nand U3289 (N_3289,N_2639,N_2577);
nand U3290 (N_3290,N_2837,N_2941);
nand U3291 (N_3291,N_2961,N_2723);
nor U3292 (N_3292,N_2582,N_2524);
and U3293 (N_3293,N_2569,N_2678);
nand U3294 (N_3294,N_2919,N_2778);
and U3295 (N_3295,N_2609,N_2529);
or U3296 (N_3296,N_2922,N_2882);
nand U3297 (N_3297,N_2538,N_2548);
nand U3298 (N_3298,N_2730,N_2791);
nand U3299 (N_3299,N_2858,N_2575);
or U3300 (N_3300,N_2875,N_2689);
and U3301 (N_3301,N_2669,N_2870);
or U3302 (N_3302,N_2948,N_2539);
nand U3303 (N_3303,N_2621,N_2977);
or U3304 (N_3304,N_2828,N_2904);
nand U3305 (N_3305,N_2673,N_2958);
and U3306 (N_3306,N_2697,N_2542);
and U3307 (N_3307,N_2795,N_2698);
nor U3308 (N_3308,N_2916,N_2641);
and U3309 (N_3309,N_2626,N_2834);
or U3310 (N_3310,N_2763,N_2677);
and U3311 (N_3311,N_2832,N_2825);
and U3312 (N_3312,N_2757,N_2705);
nand U3313 (N_3313,N_2644,N_2656);
nand U3314 (N_3314,N_2903,N_2912);
and U3315 (N_3315,N_2949,N_2596);
and U3316 (N_3316,N_2699,N_2530);
nand U3317 (N_3317,N_2551,N_2535);
nor U3318 (N_3318,N_2900,N_2664);
nor U3319 (N_3319,N_2793,N_2531);
or U3320 (N_3320,N_2942,N_2987);
or U3321 (N_3321,N_2591,N_2906);
nand U3322 (N_3322,N_2575,N_2741);
or U3323 (N_3323,N_2759,N_2956);
nand U3324 (N_3324,N_2921,N_2786);
nor U3325 (N_3325,N_2577,N_2951);
nand U3326 (N_3326,N_2925,N_2934);
or U3327 (N_3327,N_2914,N_2848);
nand U3328 (N_3328,N_2999,N_2904);
and U3329 (N_3329,N_2969,N_2667);
nor U3330 (N_3330,N_2996,N_2677);
nor U3331 (N_3331,N_2761,N_2501);
nor U3332 (N_3332,N_2801,N_2651);
nand U3333 (N_3333,N_2670,N_2630);
nor U3334 (N_3334,N_2549,N_2503);
nand U3335 (N_3335,N_2625,N_2591);
and U3336 (N_3336,N_2611,N_2633);
nor U3337 (N_3337,N_2711,N_2998);
nor U3338 (N_3338,N_2575,N_2690);
or U3339 (N_3339,N_2915,N_2623);
nor U3340 (N_3340,N_2830,N_2528);
xnor U3341 (N_3341,N_2510,N_2962);
and U3342 (N_3342,N_2829,N_2547);
nor U3343 (N_3343,N_2592,N_2726);
nand U3344 (N_3344,N_2905,N_2989);
and U3345 (N_3345,N_2542,N_2503);
nor U3346 (N_3346,N_2710,N_2991);
or U3347 (N_3347,N_2902,N_2911);
and U3348 (N_3348,N_2607,N_2849);
and U3349 (N_3349,N_2817,N_2987);
nand U3350 (N_3350,N_2728,N_2510);
or U3351 (N_3351,N_2972,N_2633);
or U3352 (N_3352,N_2708,N_2929);
xnor U3353 (N_3353,N_2535,N_2897);
or U3354 (N_3354,N_2779,N_2572);
or U3355 (N_3355,N_2738,N_2708);
nand U3356 (N_3356,N_2543,N_2842);
nand U3357 (N_3357,N_2789,N_2894);
nor U3358 (N_3358,N_2698,N_2610);
and U3359 (N_3359,N_2934,N_2967);
and U3360 (N_3360,N_2503,N_2524);
or U3361 (N_3361,N_2612,N_2595);
nand U3362 (N_3362,N_2504,N_2885);
and U3363 (N_3363,N_2600,N_2561);
nor U3364 (N_3364,N_2654,N_2615);
and U3365 (N_3365,N_2653,N_2558);
or U3366 (N_3366,N_2976,N_2963);
or U3367 (N_3367,N_2537,N_2505);
nand U3368 (N_3368,N_2573,N_2827);
nor U3369 (N_3369,N_2673,N_2614);
or U3370 (N_3370,N_2646,N_2955);
nand U3371 (N_3371,N_2923,N_2530);
nand U3372 (N_3372,N_2711,N_2557);
nor U3373 (N_3373,N_2856,N_2502);
nor U3374 (N_3374,N_2579,N_2936);
and U3375 (N_3375,N_2757,N_2799);
nand U3376 (N_3376,N_2796,N_2528);
or U3377 (N_3377,N_2886,N_2604);
nand U3378 (N_3378,N_2824,N_2981);
nor U3379 (N_3379,N_2975,N_2604);
or U3380 (N_3380,N_2928,N_2530);
and U3381 (N_3381,N_2831,N_2969);
nor U3382 (N_3382,N_2537,N_2796);
or U3383 (N_3383,N_2571,N_2818);
nor U3384 (N_3384,N_2970,N_2560);
or U3385 (N_3385,N_2893,N_2747);
nand U3386 (N_3386,N_2652,N_2769);
nor U3387 (N_3387,N_2929,N_2525);
xor U3388 (N_3388,N_2947,N_2900);
and U3389 (N_3389,N_2894,N_2606);
or U3390 (N_3390,N_2874,N_2656);
or U3391 (N_3391,N_2872,N_2985);
nand U3392 (N_3392,N_2989,N_2829);
nand U3393 (N_3393,N_2813,N_2611);
nor U3394 (N_3394,N_2578,N_2653);
or U3395 (N_3395,N_2924,N_2655);
nor U3396 (N_3396,N_2840,N_2725);
and U3397 (N_3397,N_2909,N_2995);
or U3398 (N_3398,N_2651,N_2634);
nor U3399 (N_3399,N_2865,N_2898);
and U3400 (N_3400,N_2984,N_2678);
nand U3401 (N_3401,N_2988,N_2901);
nand U3402 (N_3402,N_2877,N_2544);
nor U3403 (N_3403,N_2741,N_2500);
or U3404 (N_3404,N_2957,N_2504);
nand U3405 (N_3405,N_2701,N_2980);
and U3406 (N_3406,N_2710,N_2694);
or U3407 (N_3407,N_2998,N_2670);
nand U3408 (N_3408,N_2639,N_2987);
nand U3409 (N_3409,N_2715,N_2961);
nand U3410 (N_3410,N_2774,N_2686);
nor U3411 (N_3411,N_2846,N_2738);
and U3412 (N_3412,N_2708,N_2931);
nor U3413 (N_3413,N_2975,N_2890);
and U3414 (N_3414,N_2502,N_2829);
nand U3415 (N_3415,N_2638,N_2657);
or U3416 (N_3416,N_2562,N_2571);
or U3417 (N_3417,N_2591,N_2989);
or U3418 (N_3418,N_2989,N_2575);
or U3419 (N_3419,N_2719,N_2864);
nor U3420 (N_3420,N_2708,N_2758);
or U3421 (N_3421,N_2962,N_2855);
nor U3422 (N_3422,N_2556,N_2997);
nand U3423 (N_3423,N_2850,N_2914);
nand U3424 (N_3424,N_2698,N_2600);
nor U3425 (N_3425,N_2500,N_2523);
nor U3426 (N_3426,N_2859,N_2853);
or U3427 (N_3427,N_2814,N_2559);
nand U3428 (N_3428,N_2838,N_2547);
nor U3429 (N_3429,N_2994,N_2746);
and U3430 (N_3430,N_2825,N_2987);
or U3431 (N_3431,N_2951,N_2910);
nor U3432 (N_3432,N_2988,N_2885);
or U3433 (N_3433,N_2703,N_2549);
xnor U3434 (N_3434,N_2895,N_2796);
and U3435 (N_3435,N_2747,N_2923);
and U3436 (N_3436,N_2741,N_2528);
or U3437 (N_3437,N_2800,N_2899);
nor U3438 (N_3438,N_2888,N_2995);
or U3439 (N_3439,N_2536,N_2740);
nand U3440 (N_3440,N_2545,N_2702);
nor U3441 (N_3441,N_2803,N_2625);
nor U3442 (N_3442,N_2921,N_2704);
nor U3443 (N_3443,N_2632,N_2953);
xnor U3444 (N_3444,N_2651,N_2794);
and U3445 (N_3445,N_2732,N_2848);
nand U3446 (N_3446,N_2892,N_2664);
and U3447 (N_3447,N_2895,N_2603);
nor U3448 (N_3448,N_2755,N_2986);
or U3449 (N_3449,N_2569,N_2954);
nor U3450 (N_3450,N_2981,N_2632);
nand U3451 (N_3451,N_2941,N_2824);
and U3452 (N_3452,N_2620,N_2629);
and U3453 (N_3453,N_2776,N_2988);
and U3454 (N_3454,N_2747,N_2782);
or U3455 (N_3455,N_2513,N_2722);
or U3456 (N_3456,N_2680,N_2834);
and U3457 (N_3457,N_2912,N_2694);
nor U3458 (N_3458,N_2851,N_2657);
xnor U3459 (N_3459,N_2786,N_2811);
or U3460 (N_3460,N_2535,N_2799);
and U3461 (N_3461,N_2879,N_2623);
nand U3462 (N_3462,N_2897,N_2966);
or U3463 (N_3463,N_2963,N_2862);
nand U3464 (N_3464,N_2641,N_2825);
nor U3465 (N_3465,N_2594,N_2781);
or U3466 (N_3466,N_2518,N_2566);
nor U3467 (N_3467,N_2713,N_2674);
nand U3468 (N_3468,N_2810,N_2514);
nand U3469 (N_3469,N_2859,N_2982);
or U3470 (N_3470,N_2585,N_2704);
nor U3471 (N_3471,N_2756,N_2923);
and U3472 (N_3472,N_2899,N_2902);
and U3473 (N_3473,N_2718,N_2678);
nand U3474 (N_3474,N_2922,N_2543);
or U3475 (N_3475,N_2651,N_2927);
nor U3476 (N_3476,N_2598,N_2828);
or U3477 (N_3477,N_2606,N_2647);
nor U3478 (N_3478,N_2500,N_2750);
nor U3479 (N_3479,N_2906,N_2773);
nor U3480 (N_3480,N_2845,N_2717);
and U3481 (N_3481,N_2864,N_2894);
or U3482 (N_3482,N_2566,N_2997);
nand U3483 (N_3483,N_2762,N_2531);
nand U3484 (N_3484,N_2794,N_2903);
nor U3485 (N_3485,N_2917,N_2788);
or U3486 (N_3486,N_2829,N_2857);
nor U3487 (N_3487,N_2890,N_2710);
nand U3488 (N_3488,N_2684,N_2889);
nor U3489 (N_3489,N_2530,N_2526);
or U3490 (N_3490,N_2842,N_2540);
and U3491 (N_3491,N_2855,N_2957);
or U3492 (N_3492,N_2907,N_2709);
nor U3493 (N_3493,N_2505,N_2519);
and U3494 (N_3494,N_2858,N_2584);
nand U3495 (N_3495,N_2970,N_2917);
and U3496 (N_3496,N_2632,N_2682);
nand U3497 (N_3497,N_2916,N_2613);
nor U3498 (N_3498,N_2780,N_2931);
or U3499 (N_3499,N_2533,N_2775);
or U3500 (N_3500,N_3166,N_3139);
or U3501 (N_3501,N_3091,N_3231);
and U3502 (N_3502,N_3301,N_3040);
and U3503 (N_3503,N_3090,N_3425);
or U3504 (N_3504,N_3333,N_3329);
nor U3505 (N_3505,N_3381,N_3335);
nor U3506 (N_3506,N_3495,N_3473);
nor U3507 (N_3507,N_3097,N_3174);
and U3508 (N_3508,N_3374,N_3042);
nand U3509 (N_3509,N_3271,N_3444);
nand U3510 (N_3510,N_3272,N_3110);
nor U3511 (N_3511,N_3406,N_3454);
nand U3512 (N_3512,N_3312,N_3399);
or U3513 (N_3513,N_3325,N_3084);
nand U3514 (N_3514,N_3480,N_3075);
and U3515 (N_3515,N_3402,N_3340);
nand U3516 (N_3516,N_3129,N_3175);
nor U3517 (N_3517,N_3192,N_3177);
or U3518 (N_3518,N_3429,N_3101);
or U3519 (N_3519,N_3135,N_3268);
nand U3520 (N_3520,N_3323,N_3251);
nand U3521 (N_3521,N_3001,N_3147);
and U3522 (N_3522,N_3295,N_3159);
or U3523 (N_3523,N_3274,N_3093);
nand U3524 (N_3524,N_3146,N_3344);
and U3525 (N_3525,N_3490,N_3409);
or U3526 (N_3526,N_3049,N_3071);
nand U3527 (N_3527,N_3311,N_3064);
or U3528 (N_3528,N_3065,N_3125);
nor U3529 (N_3529,N_3099,N_3492);
nor U3530 (N_3530,N_3358,N_3478);
nand U3531 (N_3531,N_3063,N_3489);
nand U3532 (N_3532,N_3127,N_3278);
nor U3533 (N_3533,N_3208,N_3359);
nand U3534 (N_3534,N_3427,N_3293);
or U3535 (N_3535,N_3371,N_3181);
nor U3536 (N_3536,N_3004,N_3463);
xor U3537 (N_3537,N_3169,N_3431);
nor U3538 (N_3538,N_3401,N_3426);
nor U3539 (N_3539,N_3069,N_3390);
and U3540 (N_3540,N_3440,N_3031);
nand U3541 (N_3541,N_3483,N_3441);
or U3542 (N_3542,N_3186,N_3217);
nor U3543 (N_3543,N_3349,N_3354);
and U3544 (N_3544,N_3206,N_3260);
nor U3545 (N_3545,N_3043,N_3417);
nand U3546 (N_3546,N_3336,N_3182);
nand U3547 (N_3547,N_3420,N_3254);
nor U3548 (N_3548,N_3389,N_3000);
nand U3549 (N_3549,N_3197,N_3232);
and U3550 (N_3550,N_3392,N_3403);
and U3551 (N_3551,N_3317,N_3455);
or U3552 (N_3552,N_3434,N_3488);
or U3553 (N_3553,N_3338,N_3202);
or U3554 (N_3554,N_3077,N_3289);
nand U3555 (N_3555,N_3201,N_3112);
nand U3556 (N_3556,N_3252,N_3122);
or U3557 (N_3557,N_3079,N_3423);
and U3558 (N_3558,N_3219,N_3015);
and U3559 (N_3559,N_3060,N_3382);
or U3560 (N_3560,N_3088,N_3210);
nand U3561 (N_3561,N_3350,N_3414);
nor U3562 (N_3562,N_3376,N_3179);
nor U3563 (N_3563,N_3298,N_3357);
nor U3564 (N_3564,N_3080,N_3366);
and U3565 (N_3565,N_3378,N_3249);
and U3566 (N_3566,N_3485,N_3386);
or U3567 (N_3567,N_3356,N_3313);
nand U3568 (N_3568,N_3498,N_3477);
nor U3569 (N_3569,N_3465,N_3324);
and U3570 (N_3570,N_3328,N_3221);
nand U3571 (N_3571,N_3050,N_3243);
nor U3572 (N_3572,N_3062,N_3220);
nand U3573 (N_3573,N_3009,N_3308);
and U3574 (N_3574,N_3235,N_3012);
nor U3575 (N_3575,N_3353,N_3411);
nor U3576 (N_3576,N_3450,N_3037);
nor U3577 (N_3577,N_3173,N_3172);
xnor U3578 (N_3578,N_3261,N_3257);
and U3579 (N_3579,N_3048,N_3472);
and U3580 (N_3580,N_3437,N_3011);
nand U3581 (N_3581,N_3280,N_3092);
nand U3582 (N_3582,N_3034,N_3168);
nand U3583 (N_3583,N_3057,N_3113);
nand U3584 (N_3584,N_3150,N_3292);
or U3585 (N_3585,N_3275,N_3132);
nand U3586 (N_3586,N_3443,N_3006);
and U3587 (N_3587,N_3111,N_3029);
and U3588 (N_3588,N_3459,N_3284);
or U3589 (N_3589,N_3343,N_3041);
or U3590 (N_3590,N_3234,N_3487);
nor U3591 (N_3591,N_3085,N_3046);
nor U3592 (N_3592,N_3475,N_3223);
or U3593 (N_3593,N_3351,N_3380);
or U3594 (N_3594,N_3119,N_3279);
or U3595 (N_3595,N_3167,N_3030);
nor U3596 (N_3596,N_3105,N_3397);
and U3597 (N_3597,N_3385,N_3355);
or U3598 (N_3598,N_3365,N_3089);
nor U3599 (N_3599,N_3209,N_3320);
and U3600 (N_3600,N_3137,N_3290);
and U3601 (N_3601,N_3321,N_3496);
nor U3602 (N_3602,N_3407,N_3019);
and U3603 (N_3603,N_3327,N_3130);
or U3604 (N_3604,N_3400,N_3073);
and U3605 (N_3605,N_3294,N_3368);
nand U3606 (N_3606,N_3044,N_3299);
nor U3607 (N_3607,N_3416,N_3066);
or U3608 (N_3608,N_3203,N_3120);
nand U3609 (N_3609,N_3213,N_3273);
or U3610 (N_3610,N_3449,N_3211);
and U3611 (N_3611,N_3096,N_3204);
nor U3612 (N_3612,N_3134,N_3384);
and U3613 (N_3613,N_3466,N_3003);
or U3614 (N_3614,N_3393,N_3373);
and U3615 (N_3615,N_3348,N_3002);
nand U3616 (N_3616,N_3297,N_3339);
or U3617 (N_3617,N_3047,N_3151);
nor U3618 (N_3618,N_3315,N_3145);
nor U3619 (N_3619,N_3157,N_3133);
and U3620 (N_3620,N_3266,N_3229);
or U3621 (N_3621,N_3238,N_3195);
nor U3622 (N_3622,N_3383,N_3020);
nor U3623 (N_3623,N_3226,N_3141);
nand U3624 (N_3624,N_3458,N_3187);
nand U3625 (N_3625,N_3233,N_3439);
or U3626 (N_3626,N_3218,N_3387);
nor U3627 (N_3627,N_3124,N_3253);
and U3628 (N_3628,N_3337,N_3237);
and U3629 (N_3629,N_3452,N_3413);
or U3630 (N_3630,N_3138,N_3276);
and U3631 (N_3631,N_3013,N_3446);
and U3632 (N_3632,N_3142,N_3281);
and U3633 (N_3633,N_3239,N_3205);
nand U3634 (N_3634,N_3076,N_3410);
or U3635 (N_3635,N_3114,N_3148);
nand U3636 (N_3636,N_3360,N_3149);
and U3637 (N_3637,N_3106,N_3021);
or U3638 (N_3638,N_3072,N_3038);
nor U3639 (N_3639,N_3283,N_3155);
nor U3640 (N_3640,N_3070,N_3265);
nand U3641 (N_3641,N_3161,N_3396);
or U3642 (N_3642,N_3144,N_3225);
nand U3643 (N_3643,N_3282,N_3014);
and U3644 (N_3644,N_3123,N_3055);
and U3645 (N_3645,N_3039,N_3467);
nand U3646 (N_3646,N_3388,N_3346);
or U3647 (N_3647,N_3497,N_3375);
or U3648 (N_3648,N_3164,N_3200);
nor U3649 (N_3649,N_3163,N_3178);
and U3650 (N_3650,N_3116,N_3479);
and U3651 (N_3651,N_3451,N_3468);
nand U3652 (N_3652,N_3422,N_3362);
nand U3653 (N_3653,N_3018,N_3305);
and U3654 (N_3654,N_3140,N_3198);
or U3655 (N_3655,N_3236,N_3121);
and U3656 (N_3656,N_3227,N_3156);
nor U3657 (N_3657,N_3319,N_3436);
nand U3658 (N_3658,N_3094,N_3264);
and U3659 (N_3659,N_3433,N_3215);
or U3660 (N_3660,N_3484,N_3304);
or U3661 (N_3661,N_3185,N_3023);
and U3662 (N_3662,N_3470,N_3082);
and U3663 (N_3663,N_3419,N_3445);
xnor U3664 (N_3664,N_3051,N_3010);
nor U3665 (N_3665,N_3098,N_3054);
nor U3666 (N_3666,N_3053,N_3224);
or U3667 (N_3667,N_3035,N_3394);
or U3668 (N_3668,N_3245,N_3191);
nor U3669 (N_3669,N_3460,N_3270);
nand U3670 (N_3670,N_3430,N_3363);
nor U3671 (N_3671,N_3342,N_3024);
nand U3672 (N_3672,N_3448,N_3412);
nand U3673 (N_3673,N_3153,N_3256);
nor U3674 (N_3674,N_3391,N_3183);
nand U3675 (N_3675,N_3016,N_3118);
or U3676 (N_3676,N_3058,N_3395);
and U3677 (N_3677,N_3322,N_3408);
or U3678 (N_3678,N_3045,N_3469);
nand U3679 (N_3679,N_3115,N_3193);
nand U3680 (N_3680,N_3190,N_3405);
nor U3681 (N_3681,N_3296,N_3222);
or U3682 (N_3682,N_3104,N_3212);
nand U3683 (N_3683,N_3108,N_3165);
and U3684 (N_3684,N_3421,N_3246);
and U3685 (N_3685,N_3109,N_3216);
nor U3686 (N_3686,N_3081,N_3491);
nand U3687 (N_3687,N_3364,N_3083);
nor U3688 (N_3688,N_3314,N_3036);
or U3689 (N_3689,N_3309,N_3310);
nand U3690 (N_3690,N_3248,N_3143);
nor U3691 (N_3691,N_3228,N_3361);
nor U3692 (N_3692,N_3158,N_3418);
nand U3693 (N_3693,N_3347,N_3078);
nor U3694 (N_3694,N_3432,N_3318);
and U3695 (N_3695,N_3474,N_3005);
nand U3696 (N_3696,N_3263,N_3379);
nand U3697 (N_3697,N_3247,N_3059);
and U3698 (N_3698,N_3244,N_3171);
nor U3699 (N_3699,N_3269,N_3230);
or U3700 (N_3700,N_3259,N_3188);
nor U3701 (N_3701,N_3415,N_3100);
and U3702 (N_3702,N_3160,N_3462);
nor U3703 (N_3703,N_3447,N_3131);
nor U3704 (N_3704,N_3067,N_3464);
nor U3705 (N_3705,N_3331,N_3370);
or U3706 (N_3706,N_3471,N_3189);
nand U3707 (N_3707,N_3499,N_3345);
nand U3708 (N_3708,N_3250,N_3287);
nand U3709 (N_3709,N_3061,N_3486);
nor U3710 (N_3710,N_3107,N_3369);
nand U3711 (N_3711,N_3438,N_3482);
nand U3712 (N_3712,N_3493,N_3334);
and U3713 (N_3713,N_3330,N_3095);
or U3714 (N_3714,N_3288,N_3286);
nand U3715 (N_3715,N_3476,N_3128);
nor U3716 (N_3716,N_3306,N_3367);
nand U3717 (N_3717,N_3372,N_3307);
nand U3718 (N_3718,N_3240,N_3291);
nand U3719 (N_3719,N_3398,N_3102);
nand U3720 (N_3720,N_3494,N_3087);
nor U3721 (N_3721,N_3267,N_3007);
nor U3722 (N_3722,N_3285,N_3316);
nor U3723 (N_3723,N_3442,N_3241);
or U3724 (N_3724,N_3207,N_3074);
and U3725 (N_3725,N_3136,N_3377);
nand U3726 (N_3726,N_3277,N_3025);
nor U3727 (N_3727,N_3303,N_3068);
xnor U3728 (N_3728,N_3184,N_3056);
and U3729 (N_3729,N_3326,N_3435);
and U3730 (N_3730,N_3017,N_3332);
and U3731 (N_3731,N_3199,N_3126);
nor U3732 (N_3732,N_3176,N_3152);
or U3733 (N_3733,N_3457,N_3196);
and U3734 (N_3734,N_3026,N_3022);
nand U3735 (N_3735,N_3180,N_3352);
or U3736 (N_3736,N_3428,N_3033);
and U3737 (N_3737,N_3424,N_3117);
and U3738 (N_3738,N_3404,N_3052);
or U3739 (N_3739,N_3194,N_3028);
nor U3740 (N_3740,N_3086,N_3008);
nand U3741 (N_3741,N_3027,N_3341);
or U3742 (N_3742,N_3103,N_3302);
nand U3743 (N_3743,N_3456,N_3162);
nand U3744 (N_3744,N_3170,N_3461);
or U3745 (N_3745,N_3300,N_3032);
nor U3746 (N_3746,N_3242,N_3154);
nor U3747 (N_3747,N_3255,N_3262);
nand U3748 (N_3748,N_3481,N_3258);
or U3749 (N_3749,N_3453,N_3214);
nor U3750 (N_3750,N_3463,N_3065);
nand U3751 (N_3751,N_3435,N_3255);
nor U3752 (N_3752,N_3178,N_3030);
nand U3753 (N_3753,N_3358,N_3232);
xor U3754 (N_3754,N_3137,N_3426);
and U3755 (N_3755,N_3058,N_3328);
nand U3756 (N_3756,N_3419,N_3228);
and U3757 (N_3757,N_3012,N_3055);
or U3758 (N_3758,N_3400,N_3325);
nor U3759 (N_3759,N_3307,N_3004);
and U3760 (N_3760,N_3331,N_3463);
nand U3761 (N_3761,N_3128,N_3086);
and U3762 (N_3762,N_3141,N_3038);
nor U3763 (N_3763,N_3163,N_3291);
and U3764 (N_3764,N_3398,N_3259);
or U3765 (N_3765,N_3082,N_3104);
nor U3766 (N_3766,N_3490,N_3114);
or U3767 (N_3767,N_3157,N_3174);
and U3768 (N_3768,N_3304,N_3211);
or U3769 (N_3769,N_3444,N_3329);
or U3770 (N_3770,N_3024,N_3156);
nor U3771 (N_3771,N_3492,N_3159);
or U3772 (N_3772,N_3057,N_3339);
nand U3773 (N_3773,N_3334,N_3481);
or U3774 (N_3774,N_3229,N_3085);
nand U3775 (N_3775,N_3406,N_3286);
nor U3776 (N_3776,N_3153,N_3098);
or U3777 (N_3777,N_3402,N_3062);
or U3778 (N_3778,N_3325,N_3360);
nand U3779 (N_3779,N_3386,N_3269);
nor U3780 (N_3780,N_3455,N_3287);
and U3781 (N_3781,N_3281,N_3061);
or U3782 (N_3782,N_3265,N_3071);
nor U3783 (N_3783,N_3033,N_3485);
and U3784 (N_3784,N_3367,N_3377);
and U3785 (N_3785,N_3312,N_3313);
nand U3786 (N_3786,N_3324,N_3155);
nand U3787 (N_3787,N_3314,N_3312);
and U3788 (N_3788,N_3346,N_3292);
nor U3789 (N_3789,N_3410,N_3478);
nand U3790 (N_3790,N_3033,N_3363);
nor U3791 (N_3791,N_3225,N_3258);
xnor U3792 (N_3792,N_3383,N_3452);
nor U3793 (N_3793,N_3157,N_3451);
and U3794 (N_3794,N_3349,N_3201);
or U3795 (N_3795,N_3265,N_3201);
nand U3796 (N_3796,N_3395,N_3012);
and U3797 (N_3797,N_3353,N_3323);
nand U3798 (N_3798,N_3277,N_3295);
nand U3799 (N_3799,N_3411,N_3248);
nor U3800 (N_3800,N_3290,N_3261);
nor U3801 (N_3801,N_3077,N_3255);
xor U3802 (N_3802,N_3152,N_3386);
and U3803 (N_3803,N_3323,N_3173);
nor U3804 (N_3804,N_3294,N_3198);
or U3805 (N_3805,N_3282,N_3098);
nor U3806 (N_3806,N_3261,N_3459);
nor U3807 (N_3807,N_3284,N_3458);
nand U3808 (N_3808,N_3370,N_3116);
xor U3809 (N_3809,N_3421,N_3402);
nor U3810 (N_3810,N_3297,N_3131);
or U3811 (N_3811,N_3024,N_3218);
nand U3812 (N_3812,N_3344,N_3100);
or U3813 (N_3813,N_3134,N_3152);
xnor U3814 (N_3814,N_3238,N_3020);
nor U3815 (N_3815,N_3408,N_3172);
nor U3816 (N_3816,N_3404,N_3429);
or U3817 (N_3817,N_3312,N_3276);
nand U3818 (N_3818,N_3199,N_3429);
or U3819 (N_3819,N_3083,N_3493);
nor U3820 (N_3820,N_3358,N_3219);
nand U3821 (N_3821,N_3097,N_3044);
nor U3822 (N_3822,N_3375,N_3365);
and U3823 (N_3823,N_3227,N_3481);
and U3824 (N_3824,N_3415,N_3243);
or U3825 (N_3825,N_3192,N_3200);
nand U3826 (N_3826,N_3372,N_3087);
nand U3827 (N_3827,N_3180,N_3479);
nor U3828 (N_3828,N_3152,N_3304);
nand U3829 (N_3829,N_3320,N_3213);
nor U3830 (N_3830,N_3063,N_3321);
or U3831 (N_3831,N_3018,N_3000);
or U3832 (N_3832,N_3115,N_3008);
nor U3833 (N_3833,N_3443,N_3374);
and U3834 (N_3834,N_3238,N_3082);
nand U3835 (N_3835,N_3469,N_3117);
nor U3836 (N_3836,N_3371,N_3137);
and U3837 (N_3837,N_3451,N_3226);
or U3838 (N_3838,N_3487,N_3111);
nand U3839 (N_3839,N_3182,N_3304);
nor U3840 (N_3840,N_3224,N_3229);
nand U3841 (N_3841,N_3276,N_3373);
and U3842 (N_3842,N_3270,N_3135);
or U3843 (N_3843,N_3027,N_3311);
nor U3844 (N_3844,N_3464,N_3220);
or U3845 (N_3845,N_3428,N_3380);
or U3846 (N_3846,N_3429,N_3469);
and U3847 (N_3847,N_3158,N_3263);
or U3848 (N_3848,N_3012,N_3052);
or U3849 (N_3849,N_3230,N_3407);
or U3850 (N_3850,N_3172,N_3060);
and U3851 (N_3851,N_3330,N_3042);
nand U3852 (N_3852,N_3236,N_3370);
nand U3853 (N_3853,N_3471,N_3075);
nand U3854 (N_3854,N_3360,N_3102);
and U3855 (N_3855,N_3422,N_3069);
or U3856 (N_3856,N_3058,N_3164);
xor U3857 (N_3857,N_3442,N_3255);
and U3858 (N_3858,N_3394,N_3334);
and U3859 (N_3859,N_3379,N_3294);
or U3860 (N_3860,N_3149,N_3335);
and U3861 (N_3861,N_3001,N_3454);
and U3862 (N_3862,N_3145,N_3156);
or U3863 (N_3863,N_3451,N_3065);
xor U3864 (N_3864,N_3302,N_3284);
or U3865 (N_3865,N_3058,N_3126);
and U3866 (N_3866,N_3166,N_3021);
and U3867 (N_3867,N_3087,N_3180);
nand U3868 (N_3868,N_3238,N_3212);
or U3869 (N_3869,N_3129,N_3241);
and U3870 (N_3870,N_3174,N_3354);
or U3871 (N_3871,N_3260,N_3324);
nor U3872 (N_3872,N_3266,N_3414);
and U3873 (N_3873,N_3260,N_3099);
nor U3874 (N_3874,N_3027,N_3344);
or U3875 (N_3875,N_3122,N_3469);
nor U3876 (N_3876,N_3284,N_3004);
or U3877 (N_3877,N_3253,N_3264);
nor U3878 (N_3878,N_3263,N_3002);
nor U3879 (N_3879,N_3184,N_3253);
nor U3880 (N_3880,N_3481,N_3418);
and U3881 (N_3881,N_3065,N_3460);
nor U3882 (N_3882,N_3147,N_3145);
nand U3883 (N_3883,N_3476,N_3269);
nand U3884 (N_3884,N_3453,N_3304);
or U3885 (N_3885,N_3094,N_3054);
or U3886 (N_3886,N_3035,N_3072);
nor U3887 (N_3887,N_3351,N_3153);
nand U3888 (N_3888,N_3190,N_3324);
nor U3889 (N_3889,N_3054,N_3495);
nand U3890 (N_3890,N_3469,N_3448);
nand U3891 (N_3891,N_3353,N_3217);
or U3892 (N_3892,N_3180,N_3455);
xor U3893 (N_3893,N_3055,N_3096);
or U3894 (N_3894,N_3003,N_3461);
or U3895 (N_3895,N_3336,N_3239);
and U3896 (N_3896,N_3393,N_3488);
or U3897 (N_3897,N_3346,N_3443);
and U3898 (N_3898,N_3417,N_3468);
or U3899 (N_3899,N_3200,N_3480);
and U3900 (N_3900,N_3488,N_3030);
nand U3901 (N_3901,N_3231,N_3490);
nand U3902 (N_3902,N_3007,N_3134);
or U3903 (N_3903,N_3250,N_3355);
nor U3904 (N_3904,N_3387,N_3258);
or U3905 (N_3905,N_3181,N_3099);
or U3906 (N_3906,N_3115,N_3052);
nor U3907 (N_3907,N_3289,N_3497);
nand U3908 (N_3908,N_3132,N_3192);
or U3909 (N_3909,N_3056,N_3087);
or U3910 (N_3910,N_3179,N_3156);
nand U3911 (N_3911,N_3229,N_3363);
nand U3912 (N_3912,N_3279,N_3368);
and U3913 (N_3913,N_3000,N_3177);
nand U3914 (N_3914,N_3400,N_3124);
and U3915 (N_3915,N_3151,N_3053);
and U3916 (N_3916,N_3373,N_3090);
or U3917 (N_3917,N_3117,N_3344);
or U3918 (N_3918,N_3326,N_3123);
and U3919 (N_3919,N_3376,N_3459);
nor U3920 (N_3920,N_3328,N_3461);
or U3921 (N_3921,N_3264,N_3412);
or U3922 (N_3922,N_3172,N_3207);
or U3923 (N_3923,N_3271,N_3345);
or U3924 (N_3924,N_3008,N_3077);
nor U3925 (N_3925,N_3131,N_3104);
nand U3926 (N_3926,N_3003,N_3087);
and U3927 (N_3927,N_3132,N_3120);
and U3928 (N_3928,N_3240,N_3242);
nor U3929 (N_3929,N_3184,N_3214);
nand U3930 (N_3930,N_3261,N_3298);
nor U3931 (N_3931,N_3141,N_3377);
nand U3932 (N_3932,N_3018,N_3232);
nor U3933 (N_3933,N_3338,N_3224);
nor U3934 (N_3934,N_3098,N_3205);
nand U3935 (N_3935,N_3473,N_3064);
nor U3936 (N_3936,N_3096,N_3030);
nor U3937 (N_3937,N_3496,N_3375);
or U3938 (N_3938,N_3103,N_3071);
and U3939 (N_3939,N_3470,N_3191);
or U3940 (N_3940,N_3353,N_3310);
nor U3941 (N_3941,N_3256,N_3400);
nor U3942 (N_3942,N_3008,N_3308);
and U3943 (N_3943,N_3019,N_3020);
or U3944 (N_3944,N_3265,N_3170);
nor U3945 (N_3945,N_3174,N_3262);
nor U3946 (N_3946,N_3165,N_3231);
nor U3947 (N_3947,N_3147,N_3156);
and U3948 (N_3948,N_3314,N_3014);
nor U3949 (N_3949,N_3234,N_3063);
nor U3950 (N_3950,N_3257,N_3271);
and U3951 (N_3951,N_3028,N_3133);
xnor U3952 (N_3952,N_3017,N_3275);
nand U3953 (N_3953,N_3348,N_3322);
or U3954 (N_3954,N_3200,N_3404);
or U3955 (N_3955,N_3296,N_3290);
nand U3956 (N_3956,N_3251,N_3188);
nand U3957 (N_3957,N_3225,N_3301);
nand U3958 (N_3958,N_3093,N_3068);
nand U3959 (N_3959,N_3250,N_3232);
nor U3960 (N_3960,N_3212,N_3412);
nor U3961 (N_3961,N_3354,N_3407);
nor U3962 (N_3962,N_3345,N_3161);
nor U3963 (N_3963,N_3050,N_3177);
nand U3964 (N_3964,N_3349,N_3339);
or U3965 (N_3965,N_3294,N_3439);
nor U3966 (N_3966,N_3373,N_3362);
nor U3967 (N_3967,N_3496,N_3350);
nor U3968 (N_3968,N_3131,N_3259);
or U3969 (N_3969,N_3300,N_3239);
nor U3970 (N_3970,N_3267,N_3459);
and U3971 (N_3971,N_3165,N_3136);
and U3972 (N_3972,N_3320,N_3216);
nand U3973 (N_3973,N_3345,N_3147);
nand U3974 (N_3974,N_3049,N_3110);
nand U3975 (N_3975,N_3450,N_3462);
or U3976 (N_3976,N_3150,N_3251);
and U3977 (N_3977,N_3300,N_3084);
nand U3978 (N_3978,N_3094,N_3319);
or U3979 (N_3979,N_3410,N_3361);
nand U3980 (N_3980,N_3354,N_3234);
nor U3981 (N_3981,N_3461,N_3088);
and U3982 (N_3982,N_3496,N_3440);
and U3983 (N_3983,N_3452,N_3446);
or U3984 (N_3984,N_3014,N_3220);
and U3985 (N_3985,N_3403,N_3101);
nand U3986 (N_3986,N_3337,N_3430);
and U3987 (N_3987,N_3428,N_3107);
or U3988 (N_3988,N_3127,N_3288);
nor U3989 (N_3989,N_3358,N_3443);
or U3990 (N_3990,N_3287,N_3178);
nand U3991 (N_3991,N_3291,N_3142);
nand U3992 (N_3992,N_3044,N_3294);
and U3993 (N_3993,N_3247,N_3478);
and U3994 (N_3994,N_3314,N_3359);
nand U3995 (N_3995,N_3208,N_3164);
nor U3996 (N_3996,N_3324,N_3345);
or U3997 (N_3997,N_3196,N_3267);
and U3998 (N_3998,N_3401,N_3208);
nor U3999 (N_3999,N_3044,N_3420);
and U4000 (N_4000,N_3712,N_3797);
and U4001 (N_4001,N_3808,N_3983);
nand U4002 (N_4002,N_3515,N_3771);
and U4003 (N_4003,N_3953,N_3555);
or U4004 (N_4004,N_3973,N_3919);
nor U4005 (N_4005,N_3740,N_3556);
nor U4006 (N_4006,N_3876,N_3718);
or U4007 (N_4007,N_3947,N_3882);
and U4008 (N_4008,N_3747,N_3906);
nand U4009 (N_4009,N_3840,N_3870);
xnor U4010 (N_4010,N_3538,N_3957);
nand U4011 (N_4011,N_3575,N_3867);
nand U4012 (N_4012,N_3801,N_3783);
or U4013 (N_4013,N_3736,N_3595);
and U4014 (N_4014,N_3674,N_3915);
nor U4015 (N_4015,N_3985,N_3651);
nand U4016 (N_4016,N_3652,N_3803);
nand U4017 (N_4017,N_3774,N_3707);
or U4018 (N_4018,N_3883,N_3905);
nand U4019 (N_4019,N_3628,N_3881);
nor U4020 (N_4020,N_3773,N_3787);
or U4021 (N_4021,N_3616,N_3892);
nand U4022 (N_4022,N_3834,N_3946);
nor U4023 (N_4023,N_3578,N_3725);
or U4024 (N_4024,N_3574,N_3990);
nor U4025 (N_4025,N_3654,N_3609);
nor U4026 (N_4026,N_3518,N_3667);
xnor U4027 (N_4027,N_3942,N_3621);
or U4028 (N_4028,N_3878,N_3900);
nand U4029 (N_4029,N_3875,N_3861);
or U4030 (N_4030,N_3891,N_3806);
or U4031 (N_4031,N_3544,N_3733);
nand U4032 (N_4032,N_3799,N_3888);
nor U4033 (N_4033,N_3825,N_3910);
nand U4034 (N_4034,N_3590,N_3577);
nand U4035 (N_4035,N_3970,N_3701);
nor U4036 (N_4036,N_3813,N_3828);
nand U4037 (N_4037,N_3788,N_3535);
nor U4038 (N_4038,N_3602,N_3648);
or U4039 (N_4039,N_3835,N_3673);
and U4040 (N_4040,N_3645,N_3686);
or U4041 (N_4041,N_3899,N_3841);
nand U4042 (N_4042,N_3593,N_3692);
nand U4043 (N_4043,N_3669,N_3713);
and U4044 (N_4044,N_3962,N_3785);
and U4045 (N_4045,N_3711,N_3751);
and U4046 (N_4046,N_3666,N_3534);
nor U4047 (N_4047,N_3683,N_3829);
nand U4048 (N_4048,N_3898,N_3695);
nor U4049 (N_4049,N_3596,N_3597);
nor U4050 (N_4050,N_3814,N_3745);
nand U4051 (N_4051,N_3557,N_3720);
nand U4052 (N_4052,N_3591,N_3930);
nor U4053 (N_4053,N_3606,N_3886);
nor U4054 (N_4054,N_3866,N_3650);
nor U4055 (N_4055,N_3982,N_3506);
or U4056 (N_4056,N_3517,N_3735);
and U4057 (N_4057,N_3913,N_3831);
or U4058 (N_4058,N_3678,N_3991);
and U4059 (N_4059,N_3761,N_3843);
or U4060 (N_4060,N_3681,N_3559);
or U4061 (N_4061,N_3933,N_3805);
nand U4062 (N_4062,N_3880,N_3585);
or U4063 (N_4063,N_3699,N_3945);
or U4064 (N_4064,N_3856,N_3827);
nand U4065 (N_4065,N_3611,N_3586);
nor U4066 (N_4066,N_3721,N_3550);
or U4067 (N_4067,N_3939,N_3649);
and U4068 (N_4068,N_3570,N_3558);
and U4069 (N_4069,N_3975,N_3704);
nand U4070 (N_4070,N_3904,N_3664);
nand U4071 (N_4071,N_3594,N_3708);
nand U4072 (N_4072,N_3858,N_3530);
and U4073 (N_4073,N_3863,N_3765);
and U4074 (N_4074,N_3792,N_3714);
nor U4075 (N_4075,N_3989,N_3917);
and U4076 (N_4076,N_3887,N_3869);
nor U4077 (N_4077,N_3541,N_3694);
and U4078 (N_4078,N_3573,N_3912);
xnor U4079 (N_4079,N_3826,N_3968);
nand U4080 (N_4080,N_3823,N_3855);
or U4081 (N_4081,N_3563,N_3793);
nor U4082 (N_4082,N_3641,N_3763);
nand U4083 (N_4083,N_3642,N_3539);
nor U4084 (N_4084,N_3857,N_3552);
nand U4085 (N_4085,N_3696,N_3723);
nand U4086 (N_4086,N_3737,N_3698);
nand U4087 (N_4087,N_3846,N_3889);
or U4088 (N_4088,N_3922,N_3923);
and U4089 (N_4089,N_3798,N_3647);
or U4090 (N_4090,N_3623,N_3807);
or U4091 (N_4091,N_3706,N_3680);
or U4092 (N_4092,N_3739,N_3503);
or U4093 (N_4093,N_3677,N_3688);
and U4094 (N_4094,N_3546,N_3507);
nor U4095 (N_4095,N_3832,N_3702);
nor U4096 (N_4096,N_3582,N_3971);
nand U4097 (N_4097,N_3786,N_3717);
and U4098 (N_4098,N_3921,N_3655);
and U4099 (N_4099,N_3819,N_3779);
nor U4100 (N_4100,N_3873,N_3693);
and U4101 (N_4101,N_3670,N_3784);
nor U4102 (N_4102,N_3837,N_3938);
nor U4103 (N_4103,N_3551,N_3789);
and U4104 (N_4104,N_3909,N_3662);
nor U4105 (N_4105,N_3948,N_3896);
nand U4106 (N_4106,N_3543,N_3509);
or U4107 (N_4107,N_3589,N_3604);
and U4108 (N_4108,N_3549,N_3511);
and U4109 (N_4109,N_3741,N_3768);
nand U4110 (N_4110,N_3571,N_3620);
or U4111 (N_4111,N_3859,N_3790);
or U4112 (N_4112,N_3979,N_3918);
or U4113 (N_4113,N_3842,N_3569);
nor U4114 (N_4114,N_3622,N_3995);
nor U4115 (N_4115,N_3612,N_3732);
nand U4116 (N_4116,N_3877,N_3929);
or U4117 (N_4117,N_3729,N_3854);
nand U4118 (N_4118,N_3935,N_3734);
nand U4119 (N_4119,N_3653,N_3997);
nand U4120 (N_4120,N_3916,N_3850);
nor U4121 (N_4121,N_3728,N_3775);
nor U4122 (N_4122,N_3944,N_3766);
or U4123 (N_4123,N_3637,N_3848);
nand U4124 (N_4124,N_3522,N_3715);
nor U4125 (N_4125,N_3636,N_3618);
and U4126 (N_4126,N_3791,N_3658);
and U4127 (N_4127,N_3830,N_3601);
nand U4128 (N_4128,N_3526,N_3525);
nand U4129 (N_4129,N_3802,N_3816);
nand U4130 (N_4130,N_3851,N_3505);
and U4131 (N_4131,N_3613,N_3746);
xor U4132 (N_4132,N_3749,N_3588);
nand U4133 (N_4133,N_3685,N_3626);
nor U4134 (N_4134,N_3548,N_3752);
nor U4135 (N_4135,N_3937,N_3849);
and U4136 (N_4136,N_3748,N_3800);
nor U4137 (N_4137,N_3776,N_3926);
and U4138 (N_4138,N_3527,N_3815);
or U4139 (N_4139,N_3572,N_3845);
and U4140 (N_4140,N_3615,N_3890);
nand U4141 (N_4141,N_3540,N_3634);
nor U4142 (N_4142,N_3629,N_3513);
nand U4143 (N_4143,N_3777,N_3853);
nor U4144 (N_4144,N_3821,N_3961);
and U4145 (N_4145,N_3665,N_3812);
and U4146 (N_4146,N_3941,N_3836);
nand U4147 (N_4147,N_3874,N_3980);
or U4148 (N_4148,N_3724,N_3782);
or U4149 (N_4149,N_3565,N_3536);
and U4150 (N_4150,N_3547,N_3762);
and U4151 (N_4151,N_3865,N_3592);
or U4152 (N_4152,N_3633,N_3607);
or U4153 (N_4153,N_3758,N_3719);
nand U4154 (N_4154,N_3566,N_3950);
nand U4155 (N_4155,N_3581,N_3660);
and U4156 (N_4156,N_3967,N_3966);
or U4157 (N_4157,N_3969,N_3999);
or U4158 (N_4158,N_3964,N_3954);
and U4159 (N_4159,N_3772,N_3794);
or U4160 (N_4160,N_3756,N_3675);
or U4161 (N_4161,N_3579,N_3931);
nor U4162 (N_4162,N_3676,N_3608);
nand U4163 (N_4163,N_3753,N_3996);
nand U4164 (N_4164,N_3727,N_3523);
and U4165 (N_4165,N_3600,N_3568);
and U4166 (N_4166,N_3646,N_3895);
and U4167 (N_4167,N_3818,N_3940);
xor U4168 (N_4168,N_3885,N_3998);
or U4169 (N_4169,N_3852,N_3603);
nor U4170 (N_4170,N_3994,N_3679);
nand U4171 (N_4171,N_3532,N_3908);
nor U4172 (N_4172,N_3809,N_3981);
or U4173 (N_4173,N_3778,N_3897);
and U4174 (N_4174,N_3533,N_3770);
or U4175 (N_4175,N_3584,N_3959);
nand U4176 (N_4176,N_3838,N_3730);
nor U4177 (N_4177,N_3760,N_3528);
or U4178 (N_4178,N_3599,N_3907);
and U4179 (N_4179,N_3690,N_3951);
nand U4180 (N_4180,N_3554,N_3716);
and U4181 (N_4181,N_3963,N_3709);
nand U4182 (N_4182,N_3614,N_3847);
nand U4183 (N_4183,N_3965,N_3781);
nor U4184 (N_4184,N_3598,N_3700);
nor U4185 (N_4185,N_3750,N_3619);
nor U4186 (N_4186,N_3769,N_3562);
and U4187 (N_4187,N_3580,N_3710);
nand U4188 (N_4188,N_3510,N_3722);
or U4189 (N_4189,N_3583,N_3864);
nor U4190 (N_4190,N_3820,N_3920);
and U4191 (N_4191,N_3630,N_3817);
nor U4192 (N_4192,N_3810,N_3643);
or U4193 (N_4193,N_3605,N_3757);
and U4194 (N_4194,N_3932,N_3902);
nand U4195 (N_4195,N_3871,N_3671);
and U4196 (N_4196,N_3986,N_3697);
nor U4197 (N_4197,N_3524,N_3610);
nor U4198 (N_4198,N_3537,N_3520);
nor U4199 (N_4199,N_3691,N_3764);
nor U4200 (N_4200,N_3656,N_3925);
and U4201 (N_4201,N_3519,N_3624);
nand U4202 (N_4202,N_3682,N_3639);
and U4203 (N_4203,N_3504,N_3978);
nand U4204 (N_4204,N_3903,N_3934);
and U4205 (N_4205,N_3684,N_3928);
nand U4206 (N_4206,N_3631,N_3663);
and U4207 (N_4207,N_3521,N_3657);
nand U4208 (N_4208,N_3743,N_3635);
and U4209 (N_4209,N_3516,N_3755);
nor U4210 (N_4210,N_3754,N_3705);
or U4211 (N_4211,N_3508,N_3949);
and U4212 (N_4212,N_3644,N_3839);
and U4213 (N_4213,N_3956,N_3884);
nor U4214 (N_4214,N_3512,N_3576);
nor U4215 (N_4215,N_3668,N_3943);
and U4216 (N_4216,N_3759,N_3955);
nor U4217 (N_4217,N_3640,N_3984);
and U4218 (N_4218,N_3738,N_3560);
or U4219 (N_4219,N_3804,N_3868);
and U4220 (N_4220,N_3974,N_3844);
and U4221 (N_4221,N_3514,N_3879);
nand U4222 (N_4222,N_3587,N_3977);
or U4223 (N_4223,N_3795,N_3993);
or U4224 (N_4224,N_3703,N_3914);
nor U4225 (N_4225,N_3726,N_3529);
and U4226 (N_4226,N_3564,N_3893);
nor U4227 (N_4227,N_3862,N_3780);
nand U4228 (N_4228,N_3860,N_3744);
nand U4229 (N_4229,N_3824,N_3811);
or U4230 (N_4230,N_3687,N_3567);
nand U4231 (N_4231,N_3988,N_3972);
or U4232 (N_4232,N_3500,N_3638);
and U4233 (N_4233,N_3632,N_3911);
or U4234 (N_4234,N_3661,N_3822);
or U4235 (N_4235,N_3672,N_3924);
or U4236 (N_4236,N_3742,N_3976);
nand U4237 (N_4237,N_3561,N_3952);
or U4238 (N_4238,N_3894,N_3659);
and U4239 (N_4239,N_3987,N_3796);
nor U4240 (N_4240,N_3960,N_3936);
and U4241 (N_4241,N_3531,N_3767);
and U4242 (N_4242,N_3625,N_3833);
nor U4243 (N_4243,N_3545,N_3731);
and U4244 (N_4244,N_3501,N_3958);
nor U4245 (N_4245,N_3872,N_3542);
nand U4246 (N_4246,N_3901,N_3502);
nand U4247 (N_4247,N_3617,N_3627);
or U4248 (N_4248,N_3992,N_3553);
and U4249 (N_4249,N_3927,N_3689);
and U4250 (N_4250,N_3685,N_3828);
nand U4251 (N_4251,N_3749,N_3762);
or U4252 (N_4252,N_3707,N_3542);
or U4253 (N_4253,N_3502,N_3586);
and U4254 (N_4254,N_3706,N_3634);
or U4255 (N_4255,N_3793,N_3756);
nand U4256 (N_4256,N_3918,N_3924);
nand U4257 (N_4257,N_3604,N_3628);
or U4258 (N_4258,N_3928,N_3614);
or U4259 (N_4259,N_3618,N_3852);
or U4260 (N_4260,N_3598,N_3651);
nor U4261 (N_4261,N_3721,N_3680);
nand U4262 (N_4262,N_3679,N_3732);
nor U4263 (N_4263,N_3570,N_3776);
nand U4264 (N_4264,N_3903,N_3505);
nor U4265 (N_4265,N_3568,N_3880);
and U4266 (N_4266,N_3982,N_3581);
or U4267 (N_4267,N_3516,N_3638);
nand U4268 (N_4268,N_3968,N_3949);
nand U4269 (N_4269,N_3935,N_3502);
nand U4270 (N_4270,N_3604,N_3682);
or U4271 (N_4271,N_3977,N_3884);
or U4272 (N_4272,N_3771,N_3678);
or U4273 (N_4273,N_3869,N_3980);
and U4274 (N_4274,N_3952,N_3623);
and U4275 (N_4275,N_3720,N_3970);
nor U4276 (N_4276,N_3597,N_3753);
nor U4277 (N_4277,N_3544,N_3992);
or U4278 (N_4278,N_3843,N_3619);
and U4279 (N_4279,N_3513,N_3883);
nand U4280 (N_4280,N_3843,N_3778);
nand U4281 (N_4281,N_3829,N_3940);
or U4282 (N_4282,N_3553,N_3501);
or U4283 (N_4283,N_3654,N_3620);
nor U4284 (N_4284,N_3964,N_3550);
nand U4285 (N_4285,N_3726,N_3933);
nor U4286 (N_4286,N_3962,N_3842);
or U4287 (N_4287,N_3617,N_3670);
nand U4288 (N_4288,N_3568,N_3534);
and U4289 (N_4289,N_3765,N_3544);
nand U4290 (N_4290,N_3545,N_3709);
nor U4291 (N_4291,N_3826,N_3792);
nand U4292 (N_4292,N_3916,N_3692);
or U4293 (N_4293,N_3921,N_3710);
or U4294 (N_4294,N_3794,N_3602);
nor U4295 (N_4295,N_3888,N_3786);
nor U4296 (N_4296,N_3957,N_3540);
or U4297 (N_4297,N_3795,N_3990);
nor U4298 (N_4298,N_3561,N_3985);
and U4299 (N_4299,N_3893,N_3960);
nand U4300 (N_4300,N_3512,N_3618);
nand U4301 (N_4301,N_3857,N_3916);
nand U4302 (N_4302,N_3904,N_3539);
nand U4303 (N_4303,N_3515,N_3529);
and U4304 (N_4304,N_3694,N_3528);
and U4305 (N_4305,N_3644,N_3668);
and U4306 (N_4306,N_3627,N_3890);
nor U4307 (N_4307,N_3980,N_3811);
and U4308 (N_4308,N_3502,N_3993);
nor U4309 (N_4309,N_3955,N_3819);
nand U4310 (N_4310,N_3890,N_3600);
or U4311 (N_4311,N_3839,N_3869);
and U4312 (N_4312,N_3940,N_3796);
nand U4313 (N_4313,N_3754,N_3520);
or U4314 (N_4314,N_3669,N_3857);
and U4315 (N_4315,N_3527,N_3971);
nand U4316 (N_4316,N_3660,N_3900);
nand U4317 (N_4317,N_3639,N_3835);
nand U4318 (N_4318,N_3635,N_3549);
nand U4319 (N_4319,N_3659,N_3504);
nor U4320 (N_4320,N_3963,N_3674);
and U4321 (N_4321,N_3740,N_3524);
or U4322 (N_4322,N_3508,N_3770);
nor U4323 (N_4323,N_3912,N_3886);
or U4324 (N_4324,N_3746,N_3707);
and U4325 (N_4325,N_3937,N_3858);
nor U4326 (N_4326,N_3636,N_3758);
nand U4327 (N_4327,N_3886,N_3823);
nor U4328 (N_4328,N_3821,N_3970);
nand U4329 (N_4329,N_3704,N_3880);
and U4330 (N_4330,N_3720,N_3570);
or U4331 (N_4331,N_3772,N_3637);
nor U4332 (N_4332,N_3617,N_3943);
and U4333 (N_4333,N_3760,N_3534);
nor U4334 (N_4334,N_3639,N_3974);
or U4335 (N_4335,N_3882,N_3595);
nand U4336 (N_4336,N_3846,N_3670);
and U4337 (N_4337,N_3528,N_3787);
or U4338 (N_4338,N_3522,N_3560);
nor U4339 (N_4339,N_3811,N_3731);
nor U4340 (N_4340,N_3557,N_3585);
and U4341 (N_4341,N_3993,N_3535);
nand U4342 (N_4342,N_3514,N_3611);
or U4343 (N_4343,N_3916,N_3510);
nand U4344 (N_4344,N_3672,N_3791);
and U4345 (N_4345,N_3956,N_3799);
nand U4346 (N_4346,N_3950,N_3949);
and U4347 (N_4347,N_3507,N_3676);
or U4348 (N_4348,N_3776,N_3697);
and U4349 (N_4349,N_3607,N_3805);
or U4350 (N_4350,N_3542,N_3887);
nand U4351 (N_4351,N_3554,N_3694);
nand U4352 (N_4352,N_3971,N_3667);
nand U4353 (N_4353,N_3816,N_3559);
or U4354 (N_4354,N_3959,N_3662);
nand U4355 (N_4355,N_3954,N_3940);
or U4356 (N_4356,N_3614,N_3885);
or U4357 (N_4357,N_3985,N_3557);
or U4358 (N_4358,N_3988,N_3798);
and U4359 (N_4359,N_3578,N_3548);
nor U4360 (N_4360,N_3852,N_3621);
and U4361 (N_4361,N_3692,N_3697);
or U4362 (N_4362,N_3784,N_3626);
or U4363 (N_4363,N_3844,N_3560);
nor U4364 (N_4364,N_3878,N_3841);
and U4365 (N_4365,N_3886,N_3821);
and U4366 (N_4366,N_3941,N_3916);
and U4367 (N_4367,N_3807,N_3954);
nor U4368 (N_4368,N_3627,N_3805);
and U4369 (N_4369,N_3831,N_3692);
or U4370 (N_4370,N_3950,N_3807);
nand U4371 (N_4371,N_3544,N_3993);
or U4372 (N_4372,N_3892,N_3963);
and U4373 (N_4373,N_3567,N_3580);
nor U4374 (N_4374,N_3792,N_3824);
and U4375 (N_4375,N_3977,N_3803);
or U4376 (N_4376,N_3860,N_3768);
nand U4377 (N_4377,N_3549,N_3545);
and U4378 (N_4378,N_3672,N_3751);
and U4379 (N_4379,N_3526,N_3716);
and U4380 (N_4380,N_3683,N_3764);
and U4381 (N_4381,N_3572,N_3649);
or U4382 (N_4382,N_3779,N_3589);
nor U4383 (N_4383,N_3678,N_3625);
nand U4384 (N_4384,N_3598,N_3538);
nand U4385 (N_4385,N_3927,N_3726);
nor U4386 (N_4386,N_3658,N_3967);
and U4387 (N_4387,N_3912,N_3706);
nand U4388 (N_4388,N_3831,N_3842);
nand U4389 (N_4389,N_3571,N_3595);
nor U4390 (N_4390,N_3971,N_3520);
or U4391 (N_4391,N_3884,N_3907);
and U4392 (N_4392,N_3671,N_3512);
nand U4393 (N_4393,N_3581,N_3594);
nand U4394 (N_4394,N_3879,N_3976);
or U4395 (N_4395,N_3848,N_3750);
or U4396 (N_4396,N_3686,N_3731);
and U4397 (N_4397,N_3922,N_3736);
or U4398 (N_4398,N_3875,N_3907);
and U4399 (N_4399,N_3937,N_3888);
and U4400 (N_4400,N_3528,N_3860);
and U4401 (N_4401,N_3681,N_3957);
nor U4402 (N_4402,N_3757,N_3715);
nand U4403 (N_4403,N_3675,N_3822);
and U4404 (N_4404,N_3935,N_3852);
nand U4405 (N_4405,N_3614,N_3683);
or U4406 (N_4406,N_3658,N_3632);
nor U4407 (N_4407,N_3714,N_3633);
and U4408 (N_4408,N_3678,N_3999);
nor U4409 (N_4409,N_3834,N_3527);
nand U4410 (N_4410,N_3746,N_3691);
or U4411 (N_4411,N_3546,N_3629);
nand U4412 (N_4412,N_3666,N_3769);
nand U4413 (N_4413,N_3866,N_3770);
nand U4414 (N_4414,N_3655,N_3793);
or U4415 (N_4415,N_3873,N_3684);
nor U4416 (N_4416,N_3755,N_3622);
nor U4417 (N_4417,N_3507,N_3754);
nor U4418 (N_4418,N_3730,N_3660);
nand U4419 (N_4419,N_3911,N_3985);
nand U4420 (N_4420,N_3594,N_3732);
and U4421 (N_4421,N_3545,N_3955);
nand U4422 (N_4422,N_3867,N_3916);
nand U4423 (N_4423,N_3908,N_3921);
nor U4424 (N_4424,N_3720,N_3657);
and U4425 (N_4425,N_3954,N_3971);
and U4426 (N_4426,N_3720,N_3988);
and U4427 (N_4427,N_3878,N_3992);
nand U4428 (N_4428,N_3542,N_3993);
nor U4429 (N_4429,N_3741,N_3690);
nor U4430 (N_4430,N_3665,N_3532);
or U4431 (N_4431,N_3748,N_3973);
or U4432 (N_4432,N_3570,N_3835);
or U4433 (N_4433,N_3834,N_3758);
and U4434 (N_4434,N_3861,N_3901);
xor U4435 (N_4435,N_3993,N_3504);
nand U4436 (N_4436,N_3929,N_3536);
nand U4437 (N_4437,N_3952,N_3666);
nand U4438 (N_4438,N_3992,N_3798);
and U4439 (N_4439,N_3656,N_3619);
and U4440 (N_4440,N_3787,N_3955);
and U4441 (N_4441,N_3874,N_3773);
nor U4442 (N_4442,N_3726,N_3653);
nand U4443 (N_4443,N_3643,N_3569);
nor U4444 (N_4444,N_3830,N_3927);
nor U4445 (N_4445,N_3740,N_3586);
nand U4446 (N_4446,N_3977,N_3877);
nand U4447 (N_4447,N_3613,N_3627);
nand U4448 (N_4448,N_3563,N_3552);
nand U4449 (N_4449,N_3761,N_3576);
nand U4450 (N_4450,N_3553,N_3779);
and U4451 (N_4451,N_3730,N_3579);
xor U4452 (N_4452,N_3843,N_3821);
or U4453 (N_4453,N_3824,N_3852);
nor U4454 (N_4454,N_3677,N_3554);
or U4455 (N_4455,N_3867,N_3502);
nor U4456 (N_4456,N_3720,N_3813);
nor U4457 (N_4457,N_3972,N_3744);
nor U4458 (N_4458,N_3985,N_3714);
and U4459 (N_4459,N_3750,N_3902);
nand U4460 (N_4460,N_3630,N_3762);
and U4461 (N_4461,N_3986,N_3875);
nand U4462 (N_4462,N_3673,N_3932);
or U4463 (N_4463,N_3935,N_3987);
nand U4464 (N_4464,N_3647,N_3702);
nand U4465 (N_4465,N_3551,N_3905);
or U4466 (N_4466,N_3873,N_3822);
or U4467 (N_4467,N_3964,N_3909);
or U4468 (N_4468,N_3980,N_3783);
nand U4469 (N_4469,N_3682,N_3894);
nor U4470 (N_4470,N_3978,N_3591);
nor U4471 (N_4471,N_3610,N_3602);
nor U4472 (N_4472,N_3729,N_3920);
nand U4473 (N_4473,N_3689,N_3840);
xor U4474 (N_4474,N_3784,N_3816);
and U4475 (N_4475,N_3975,N_3962);
nand U4476 (N_4476,N_3910,N_3879);
nand U4477 (N_4477,N_3535,N_3934);
nand U4478 (N_4478,N_3658,N_3914);
and U4479 (N_4479,N_3636,N_3962);
nand U4480 (N_4480,N_3569,N_3636);
and U4481 (N_4481,N_3928,N_3777);
and U4482 (N_4482,N_3831,N_3982);
nor U4483 (N_4483,N_3893,N_3782);
or U4484 (N_4484,N_3723,N_3998);
nor U4485 (N_4485,N_3709,N_3772);
nor U4486 (N_4486,N_3665,N_3874);
nor U4487 (N_4487,N_3591,N_3903);
and U4488 (N_4488,N_3567,N_3805);
nand U4489 (N_4489,N_3995,N_3635);
nor U4490 (N_4490,N_3924,N_3895);
and U4491 (N_4491,N_3759,N_3546);
nor U4492 (N_4492,N_3514,N_3756);
nand U4493 (N_4493,N_3625,N_3528);
nand U4494 (N_4494,N_3835,N_3567);
and U4495 (N_4495,N_3988,N_3630);
or U4496 (N_4496,N_3732,N_3812);
or U4497 (N_4497,N_3972,N_3908);
or U4498 (N_4498,N_3980,N_3818);
or U4499 (N_4499,N_3536,N_3764);
nand U4500 (N_4500,N_4372,N_4197);
nor U4501 (N_4501,N_4199,N_4410);
or U4502 (N_4502,N_4336,N_4185);
and U4503 (N_4503,N_4125,N_4433);
nor U4504 (N_4504,N_4061,N_4444);
and U4505 (N_4505,N_4368,N_4473);
and U4506 (N_4506,N_4041,N_4068);
nor U4507 (N_4507,N_4218,N_4394);
nand U4508 (N_4508,N_4173,N_4355);
and U4509 (N_4509,N_4175,N_4145);
and U4510 (N_4510,N_4172,N_4347);
or U4511 (N_4511,N_4134,N_4021);
and U4512 (N_4512,N_4201,N_4076);
nor U4513 (N_4513,N_4111,N_4075);
nor U4514 (N_4514,N_4128,N_4087);
or U4515 (N_4515,N_4077,N_4055);
and U4516 (N_4516,N_4441,N_4256);
nand U4517 (N_4517,N_4406,N_4169);
nor U4518 (N_4518,N_4296,N_4388);
nor U4519 (N_4519,N_4133,N_4019);
nor U4520 (N_4520,N_4074,N_4351);
nand U4521 (N_4521,N_4320,N_4225);
or U4522 (N_4522,N_4426,N_4117);
nor U4523 (N_4523,N_4017,N_4308);
nor U4524 (N_4524,N_4483,N_4335);
or U4525 (N_4525,N_4311,N_4271);
and U4526 (N_4526,N_4385,N_4151);
and U4527 (N_4527,N_4063,N_4094);
or U4528 (N_4528,N_4285,N_4364);
and U4529 (N_4529,N_4162,N_4438);
nor U4530 (N_4530,N_4013,N_4284);
or U4531 (N_4531,N_4227,N_4062);
xor U4532 (N_4532,N_4010,N_4114);
nand U4533 (N_4533,N_4044,N_4238);
nand U4534 (N_4534,N_4290,N_4281);
or U4535 (N_4535,N_4093,N_4069);
nor U4536 (N_4536,N_4480,N_4437);
and U4537 (N_4537,N_4136,N_4179);
nand U4538 (N_4538,N_4052,N_4485);
nand U4539 (N_4539,N_4393,N_4082);
and U4540 (N_4540,N_4064,N_4100);
and U4541 (N_4541,N_4186,N_4229);
nand U4542 (N_4542,N_4342,N_4253);
nor U4543 (N_4543,N_4261,N_4011);
or U4544 (N_4544,N_4423,N_4424);
and U4545 (N_4545,N_4101,N_4325);
nor U4546 (N_4546,N_4371,N_4083);
or U4547 (N_4547,N_4081,N_4251);
nor U4548 (N_4548,N_4012,N_4152);
and U4549 (N_4549,N_4163,N_4331);
or U4550 (N_4550,N_4001,N_4155);
or U4551 (N_4551,N_4436,N_4139);
nand U4552 (N_4552,N_4360,N_4099);
and U4553 (N_4553,N_4432,N_4260);
or U4554 (N_4554,N_4192,N_4334);
nor U4555 (N_4555,N_4465,N_4318);
nand U4556 (N_4556,N_4124,N_4126);
xnor U4557 (N_4557,N_4211,N_4143);
and U4558 (N_4558,N_4291,N_4498);
and U4559 (N_4559,N_4269,N_4427);
nor U4560 (N_4560,N_4065,N_4234);
nand U4561 (N_4561,N_4359,N_4499);
nand U4562 (N_4562,N_4080,N_4088);
or U4563 (N_4563,N_4109,N_4428);
nand U4564 (N_4564,N_4149,N_4419);
and U4565 (N_4565,N_4484,N_4166);
nand U4566 (N_4566,N_4452,N_4210);
and U4567 (N_4567,N_4369,N_4167);
or U4568 (N_4568,N_4206,N_4490);
or U4569 (N_4569,N_4466,N_4130);
nor U4570 (N_4570,N_4110,N_4407);
nand U4571 (N_4571,N_4492,N_4303);
and U4572 (N_4572,N_4242,N_4416);
nor U4573 (N_4573,N_4333,N_4220);
nand U4574 (N_4574,N_4144,N_4178);
or U4575 (N_4575,N_4434,N_4189);
nor U4576 (N_4576,N_4453,N_4383);
nand U4577 (N_4577,N_4298,N_4215);
nand U4578 (N_4578,N_4262,N_4137);
or U4579 (N_4579,N_4038,N_4319);
or U4580 (N_4580,N_4268,N_4121);
nand U4581 (N_4581,N_4307,N_4309);
and U4582 (N_4582,N_4020,N_4397);
or U4583 (N_4583,N_4447,N_4265);
nand U4584 (N_4584,N_4373,N_4187);
nand U4585 (N_4585,N_4207,N_4129);
and U4586 (N_4586,N_4243,N_4079);
or U4587 (N_4587,N_4244,N_4487);
or U4588 (N_4588,N_4366,N_4212);
or U4589 (N_4589,N_4477,N_4050);
or U4590 (N_4590,N_4398,N_4156);
nand U4591 (N_4591,N_4195,N_4247);
or U4592 (N_4592,N_4387,N_4037);
nand U4593 (N_4593,N_4395,N_4203);
nand U4594 (N_4594,N_4131,N_4098);
nor U4595 (N_4595,N_4140,N_4489);
nand U4596 (N_4596,N_4445,N_4159);
nor U4597 (N_4597,N_4002,N_4056);
nand U4598 (N_4598,N_4448,N_4354);
nand U4599 (N_4599,N_4376,N_4408);
nand U4600 (N_4600,N_4022,N_4026);
nand U4601 (N_4601,N_4409,N_4214);
nor U4602 (N_4602,N_4259,N_4328);
nand U4603 (N_4603,N_4246,N_4174);
nor U4604 (N_4604,N_4341,N_4415);
and U4605 (N_4605,N_4405,N_4297);
or U4606 (N_4606,N_4032,N_4435);
nor U4607 (N_4607,N_4177,N_4182);
and U4608 (N_4608,N_4183,N_4067);
nand U4609 (N_4609,N_4420,N_4361);
nor U4610 (N_4610,N_4078,N_4375);
nand U4611 (N_4611,N_4188,N_4289);
nor U4612 (N_4612,N_4232,N_4226);
nand U4613 (N_4613,N_4392,N_4219);
and U4614 (N_4614,N_4272,N_4476);
or U4615 (N_4615,N_4474,N_4497);
and U4616 (N_4616,N_4164,N_4250);
or U4617 (N_4617,N_4115,N_4066);
nor U4618 (N_4618,N_4107,N_4141);
nand U4619 (N_4619,N_4348,N_4165);
and U4620 (N_4620,N_4413,N_4494);
and U4621 (N_4621,N_4469,N_4472);
and U4622 (N_4622,N_4464,N_4058);
or U4623 (N_4623,N_4148,N_4005);
and U4624 (N_4624,N_4326,N_4471);
or U4625 (N_4625,N_4449,N_4299);
or U4626 (N_4626,N_4118,N_4157);
and U4627 (N_4627,N_4198,N_4495);
and U4628 (N_4628,N_4459,N_4209);
nor U4629 (N_4629,N_4488,N_4430);
or U4630 (N_4630,N_4000,N_4034);
and U4631 (N_4631,N_4181,N_4104);
and U4632 (N_4632,N_4193,N_4412);
and U4633 (N_4633,N_4027,N_4016);
or U4634 (N_4634,N_4146,N_4239);
nand U4635 (N_4635,N_4241,N_4377);
nand U4636 (N_4636,N_4270,N_4030);
or U4637 (N_4637,N_4301,N_4329);
and U4638 (N_4638,N_4105,N_4053);
and U4639 (N_4639,N_4302,N_4237);
nand U4640 (N_4640,N_4451,N_4086);
and U4641 (N_4641,N_4120,N_4276);
nor U4642 (N_4642,N_4403,N_4048);
nand U4643 (N_4643,N_4184,N_4442);
nor U4644 (N_4644,N_4305,N_4221);
nor U4645 (N_4645,N_4379,N_4462);
or U4646 (N_4646,N_4386,N_4382);
nand U4647 (N_4647,N_4003,N_4194);
nor U4648 (N_4648,N_4332,N_4071);
or U4649 (N_4649,N_4353,N_4035);
nor U4650 (N_4650,N_4029,N_4092);
nand U4651 (N_4651,N_4421,N_4292);
and U4652 (N_4652,N_4344,N_4028);
nand U4653 (N_4653,N_4127,N_4363);
and U4654 (N_4654,N_4417,N_4240);
and U4655 (N_4655,N_4161,N_4378);
and U4656 (N_4656,N_4425,N_4370);
and U4657 (N_4657,N_4180,N_4039);
or U4658 (N_4658,N_4322,N_4043);
nor U4659 (N_4659,N_4401,N_4264);
or U4660 (N_4660,N_4231,N_4455);
nand U4661 (N_4661,N_4317,N_4147);
nand U4662 (N_4662,N_4249,N_4036);
nor U4663 (N_4663,N_4486,N_4280);
or U4664 (N_4664,N_4481,N_4399);
or U4665 (N_4665,N_4414,N_4084);
or U4666 (N_4666,N_4170,N_4018);
nor U4667 (N_4667,N_4306,N_4461);
nor U4668 (N_4668,N_4337,N_4190);
nand U4669 (N_4669,N_4112,N_4095);
nor U4670 (N_4670,N_4293,N_4321);
or U4671 (N_4671,N_4400,N_4478);
nor U4672 (N_4672,N_4278,N_4257);
or U4673 (N_4673,N_4191,N_4283);
nand U4674 (N_4674,N_4482,N_4491);
nand U4675 (N_4675,N_4224,N_4235);
nor U4676 (N_4676,N_4213,N_4286);
and U4677 (N_4677,N_4357,N_4365);
or U4678 (N_4678,N_4258,N_4205);
nand U4679 (N_4679,N_4277,N_4345);
nor U4680 (N_4680,N_4389,N_4454);
nand U4681 (N_4681,N_4295,N_4054);
nand U4682 (N_4682,N_4255,N_4208);
and U4683 (N_4683,N_4440,N_4315);
nor U4684 (N_4684,N_4443,N_4228);
nand U4685 (N_4685,N_4463,N_4008);
nor U4686 (N_4686,N_4288,N_4047);
and U4687 (N_4687,N_4103,N_4142);
nor U4688 (N_4688,N_4254,N_4340);
nor U4689 (N_4689,N_4304,N_4468);
and U4690 (N_4690,N_4113,N_4279);
nand U4691 (N_4691,N_4362,N_4085);
nand U4692 (N_4692,N_4070,N_4316);
nor U4693 (N_4693,N_4200,N_4116);
and U4694 (N_4694,N_4402,N_4349);
nand U4695 (N_4695,N_4358,N_4324);
nand U4696 (N_4696,N_4346,N_4217);
and U4697 (N_4697,N_4135,N_4352);
nand U4698 (N_4698,N_4356,N_4367);
nand U4699 (N_4699,N_4404,N_4230);
nor U4700 (N_4700,N_4411,N_4381);
and U4701 (N_4701,N_4106,N_4216);
nor U4702 (N_4702,N_4470,N_4431);
or U4703 (N_4703,N_4014,N_4446);
nand U4704 (N_4704,N_4153,N_4097);
and U4705 (N_4705,N_4310,N_4493);
nor U4706 (N_4706,N_4202,N_4294);
nor U4707 (N_4707,N_4275,N_4158);
nand U4708 (N_4708,N_4273,N_4467);
nor U4709 (N_4709,N_4040,N_4327);
xor U4710 (N_4710,N_4073,N_4150);
and U4711 (N_4711,N_4176,N_4096);
nor U4712 (N_4712,N_4015,N_4313);
and U4713 (N_4713,N_4223,N_4004);
and U4714 (N_4714,N_4132,N_4456);
nand U4715 (N_4715,N_4475,N_4204);
nor U4716 (N_4716,N_4245,N_4154);
nand U4717 (N_4717,N_4343,N_4090);
nor U4718 (N_4718,N_4496,N_4060);
or U4719 (N_4719,N_4282,N_4042);
nor U4720 (N_4720,N_4051,N_4045);
and U4721 (N_4721,N_4222,N_4263);
and U4722 (N_4722,N_4009,N_4312);
or U4723 (N_4723,N_4439,N_4160);
and U4724 (N_4724,N_4422,N_4089);
nand U4725 (N_4725,N_4450,N_4057);
nor U4726 (N_4726,N_4300,N_4391);
nor U4727 (N_4727,N_4091,N_4007);
nor U4728 (N_4728,N_4460,N_4390);
nand U4729 (N_4729,N_4023,N_4330);
nand U4730 (N_4730,N_4396,N_4123);
or U4731 (N_4731,N_4102,N_4233);
nor U4732 (N_4732,N_4236,N_4266);
and U4733 (N_4733,N_4457,N_4418);
nor U4734 (N_4734,N_4138,N_4049);
or U4735 (N_4735,N_4033,N_4024);
nand U4736 (N_4736,N_4380,N_4031);
nand U4737 (N_4737,N_4025,N_4314);
nand U4738 (N_4738,N_4274,N_4479);
nand U4739 (N_4739,N_4323,N_4171);
nor U4740 (N_4740,N_4196,N_4338);
or U4741 (N_4741,N_4429,N_4122);
xnor U4742 (N_4742,N_4384,N_4339);
and U4743 (N_4743,N_4119,N_4374);
nor U4744 (N_4744,N_4350,N_4252);
and U4745 (N_4745,N_4248,N_4046);
nand U4746 (N_4746,N_4458,N_4108);
nor U4747 (N_4747,N_4287,N_4072);
or U4748 (N_4748,N_4059,N_4006);
or U4749 (N_4749,N_4267,N_4168);
or U4750 (N_4750,N_4423,N_4466);
nor U4751 (N_4751,N_4109,N_4328);
nor U4752 (N_4752,N_4368,N_4367);
nor U4753 (N_4753,N_4101,N_4465);
nor U4754 (N_4754,N_4290,N_4058);
or U4755 (N_4755,N_4236,N_4156);
and U4756 (N_4756,N_4161,N_4436);
and U4757 (N_4757,N_4078,N_4491);
nand U4758 (N_4758,N_4260,N_4074);
nor U4759 (N_4759,N_4204,N_4187);
or U4760 (N_4760,N_4388,N_4346);
and U4761 (N_4761,N_4286,N_4351);
nor U4762 (N_4762,N_4071,N_4079);
and U4763 (N_4763,N_4382,N_4332);
and U4764 (N_4764,N_4200,N_4378);
and U4765 (N_4765,N_4346,N_4120);
or U4766 (N_4766,N_4006,N_4223);
or U4767 (N_4767,N_4181,N_4332);
nor U4768 (N_4768,N_4267,N_4230);
or U4769 (N_4769,N_4118,N_4068);
or U4770 (N_4770,N_4168,N_4422);
nand U4771 (N_4771,N_4416,N_4431);
nand U4772 (N_4772,N_4396,N_4434);
or U4773 (N_4773,N_4044,N_4492);
and U4774 (N_4774,N_4133,N_4120);
or U4775 (N_4775,N_4185,N_4453);
nor U4776 (N_4776,N_4435,N_4292);
and U4777 (N_4777,N_4476,N_4303);
or U4778 (N_4778,N_4088,N_4422);
nand U4779 (N_4779,N_4158,N_4392);
nor U4780 (N_4780,N_4227,N_4282);
or U4781 (N_4781,N_4290,N_4480);
or U4782 (N_4782,N_4421,N_4340);
nor U4783 (N_4783,N_4126,N_4465);
nor U4784 (N_4784,N_4088,N_4433);
nand U4785 (N_4785,N_4075,N_4156);
or U4786 (N_4786,N_4266,N_4155);
and U4787 (N_4787,N_4236,N_4040);
nand U4788 (N_4788,N_4110,N_4263);
nand U4789 (N_4789,N_4327,N_4387);
nand U4790 (N_4790,N_4127,N_4457);
or U4791 (N_4791,N_4414,N_4491);
or U4792 (N_4792,N_4253,N_4098);
and U4793 (N_4793,N_4364,N_4363);
nor U4794 (N_4794,N_4108,N_4224);
and U4795 (N_4795,N_4245,N_4450);
nand U4796 (N_4796,N_4002,N_4202);
nor U4797 (N_4797,N_4023,N_4392);
or U4798 (N_4798,N_4255,N_4155);
nand U4799 (N_4799,N_4447,N_4286);
or U4800 (N_4800,N_4398,N_4403);
or U4801 (N_4801,N_4274,N_4328);
and U4802 (N_4802,N_4286,N_4352);
nor U4803 (N_4803,N_4269,N_4348);
and U4804 (N_4804,N_4484,N_4381);
or U4805 (N_4805,N_4286,N_4295);
and U4806 (N_4806,N_4014,N_4271);
and U4807 (N_4807,N_4263,N_4224);
and U4808 (N_4808,N_4396,N_4284);
nand U4809 (N_4809,N_4017,N_4439);
or U4810 (N_4810,N_4221,N_4395);
or U4811 (N_4811,N_4094,N_4152);
and U4812 (N_4812,N_4228,N_4264);
nor U4813 (N_4813,N_4023,N_4429);
nand U4814 (N_4814,N_4258,N_4369);
nor U4815 (N_4815,N_4239,N_4384);
xnor U4816 (N_4816,N_4298,N_4278);
or U4817 (N_4817,N_4235,N_4380);
nand U4818 (N_4818,N_4231,N_4070);
or U4819 (N_4819,N_4234,N_4143);
or U4820 (N_4820,N_4161,N_4098);
and U4821 (N_4821,N_4161,N_4078);
nor U4822 (N_4822,N_4410,N_4419);
nand U4823 (N_4823,N_4267,N_4203);
nand U4824 (N_4824,N_4308,N_4204);
nand U4825 (N_4825,N_4372,N_4395);
xnor U4826 (N_4826,N_4096,N_4032);
nand U4827 (N_4827,N_4444,N_4419);
or U4828 (N_4828,N_4484,N_4304);
nand U4829 (N_4829,N_4219,N_4347);
and U4830 (N_4830,N_4433,N_4084);
xor U4831 (N_4831,N_4344,N_4376);
or U4832 (N_4832,N_4182,N_4025);
nor U4833 (N_4833,N_4036,N_4171);
xor U4834 (N_4834,N_4058,N_4187);
and U4835 (N_4835,N_4017,N_4104);
or U4836 (N_4836,N_4276,N_4305);
nor U4837 (N_4837,N_4018,N_4096);
and U4838 (N_4838,N_4130,N_4047);
and U4839 (N_4839,N_4029,N_4208);
nor U4840 (N_4840,N_4222,N_4126);
nor U4841 (N_4841,N_4256,N_4047);
nand U4842 (N_4842,N_4283,N_4093);
nand U4843 (N_4843,N_4277,N_4413);
and U4844 (N_4844,N_4424,N_4200);
or U4845 (N_4845,N_4277,N_4416);
nand U4846 (N_4846,N_4184,N_4128);
and U4847 (N_4847,N_4417,N_4141);
nor U4848 (N_4848,N_4318,N_4395);
or U4849 (N_4849,N_4303,N_4299);
and U4850 (N_4850,N_4371,N_4286);
nand U4851 (N_4851,N_4206,N_4437);
or U4852 (N_4852,N_4073,N_4238);
nand U4853 (N_4853,N_4200,N_4296);
and U4854 (N_4854,N_4371,N_4096);
or U4855 (N_4855,N_4129,N_4264);
nor U4856 (N_4856,N_4126,N_4112);
and U4857 (N_4857,N_4284,N_4434);
nor U4858 (N_4858,N_4089,N_4335);
nand U4859 (N_4859,N_4233,N_4443);
and U4860 (N_4860,N_4065,N_4184);
nor U4861 (N_4861,N_4241,N_4347);
xnor U4862 (N_4862,N_4265,N_4336);
nand U4863 (N_4863,N_4200,N_4351);
nand U4864 (N_4864,N_4493,N_4404);
or U4865 (N_4865,N_4309,N_4259);
or U4866 (N_4866,N_4014,N_4147);
and U4867 (N_4867,N_4078,N_4228);
nand U4868 (N_4868,N_4185,N_4165);
nor U4869 (N_4869,N_4489,N_4109);
and U4870 (N_4870,N_4166,N_4245);
nand U4871 (N_4871,N_4057,N_4202);
nand U4872 (N_4872,N_4080,N_4336);
nand U4873 (N_4873,N_4307,N_4494);
or U4874 (N_4874,N_4151,N_4373);
and U4875 (N_4875,N_4358,N_4024);
nor U4876 (N_4876,N_4279,N_4152);
nand U4877 (N_4877,N_4334,N_4415);
nor U4878 (N_4878,N_4150,N_4311);
nor U4879 (N_4879,N_4222,N_4297);
or U4880 (N_4880,N_4209,N_4477);
nand U4881 (N_4881,N_4218,N_4091);
and U4882 (N_4882,N_4165,N_4484);
or U4883 (N_4883,N_4378,N_4463);
nand U4884 (N_4884,N_4004,N_4114);
or U4885 (N_4885,N_4299,N_4086);
and U4886 (N_4886,N_4104,N_4216);
nand U4887 (N_4887,N_4345,N_4097);
nor U4888 (N_4888,N_4411,N_4252);
xnor U4889 (N_4889,N_4345,N_4438);
or U4890 (N_4890,N_4230,N_4166);
nor U4891 (N_4891,N_4129,N_4137);
nor U4892 (N_4892,N_4311,N_4252);
or U4893 (N_4893,N_4410,N_4333);
nor U4894 (N_4894,N_4387,N_4305);
and U4895 (N_4895,N_4203,N_4254);
nor U4896 (N_4896,N_4454,N_4125);
nor U4897 (N_4897,N_4427,N_4412);
nand U4898 (N_4898,N_4398,N_4053);
nand U4899 (N_4899,N_4304,N_4461);
and U4900 (N_4900,N_4091,N_4289);
or U4901 (N_4901,N_4018,N_4215);
or U4902 (N_4902,N_4218,N_4138);
and U4903 (N_4903,N_4136,N_4440);
and U4904 (N_4904,N_4468,N_4494);
nand U4905 (N_4905,N_4035,N_4146);
or U4906 (N_4906,N_4295,N_4310);
and U4907 (N_4907,N_4198,N_4166);
nor U4908 (N_4908,N_4362,N_4188);
or U4909 (N_4909,N_4331,N_4004);
nor U4910 (N_4910,N_4066,N_4032);
nand U4911 (N_4911,N_4157,N_4097);
and U4912 (N_4912,N_4460,N_4093);
nor U4913 (N_4913,N_4074,N_4266);
nand U4914 (N_4914,N_4019,N_4338);
and U4915 (N_4915,N_4487,N_4079);
nor U4916 (N_4916,N_4313,N_4323);
nor U4917 (N_4917,N_4075,N_4113);
or U4918 (N_4918,N_4370,N_4114);
or U4919 (N_4919,N_4099,N_4105);
nand U4920 (N_4920,N_4104,N_4149);
and U4921 (N_4921,N_4411,N_4023);
nor U4922 (N_4922,N_4428,N_4260);
nand U4923 (N_4923,N_4307,N_4240);
nor U4924 (N_4924,N_4493,N_4473);
nor U4925 (N_4925,N_4158,N_4053);
and U4926 (N_4926,N_4146,N_4333);
nand U4927 (N_4927,N_4224,N_4128);
nor U4928 (N_4928,N_4462,N_4027);
nor U4929 (N_4929,N_4449,N_4189);
nor U4930 (N_4930,N_4460,N_4467);
or U4931 (N_4931,N_4084,N_4040);
nor U4932 (N_4932,N_4405,N_4282);
nand U4933 (N_4933,N_4199,N_4108);
and U4934 (N_4934,N_4131,N_4041);
nor U4935 (N_4935,N_4195,N_4304);
nand U4936 (N_4936,N_4021,N_4430);
and U4937 (N_4937,N_4072,N_4394);
and U4938 (N_4938,N_4255,N_4311);
nand U4939 (N_4939,N_4240,N_4165);
nor U4940 (N_4940,N_4208,N_4109);
and U4941 (N_4941,N_4496,N_4204);
xnor U4942 (N_4942,N_4362,N_4305);
nor U4943 (N_4943,N_4254,N_4213);
nor U4944 (N_4944,N_4388,N_4325);
or U4945 (N_4945,N_4051,N_4028);
nand U4946 (N_4946,N_4023,N_4278);
nand U4947 (N_4947,N_4106,N_4170);
and U4948 (N_4948,N_4250,N_4119);
or U4949 (N_4949,N_4000,N_4251);
nand U4950 (N_4950,N_4251,N_4474);
and U4951 (N_4951,N_4204,N_4216);
and U4952 (N_4952,N_4410,N_4273);
nand U4953 (N_4953,N_4418,N_4349);
nor U4954 (N_4954,N_4326,N_4321);
and U4955 (N_4955,N_4343,N_4289);
or U4956 (N_4956,N_4204,N_4194);
nor U4957 (N_4957,N_4412,N_4302);
or U4958 (N_4958,N_4037,N_4280);
or U4959 (N_4959,N_4122,N_4017);
nor U4960 (N_4960,N_4282,N_4092);
and U4961 (N_4961,N_4458,N_4190);
or U4962 (N_4962,N_4238,N_4352);
nor U4963 (N_4963,N_4027,N_4047);
nor U4964 (N_4964,N_4480,N_4070);
nand U4965 (N_4965,N_4410,N_4318);
or U4966 (N_4966,N_4371,N_4084);
and U4967 (N_4967,N_4148,N_4357);
nor U4968 (N_4968,N_4179,N_4129);
or U4969 (N_4969,N_4329,N_4441);
or U4970 (N_4970,N_4045,N_4067);
nand U4971 (N_4971,N_4386,N_4029);
and U4972 (N_4972,N_4247,N_4234);
and U4973 (N_4973,N_4463,N_4140);
or U4974 (N_4974,N_4100,N_4337);
nand U4975 (N_4975,N_4027,N_4088);
nor U4976 (N_4976,N_4267,N_4301);
nand U4977 (N_4977,N_4366,N_4231);
nor U4978 (N_4978,N_4255,N_4210);
and U4979 (N_4979,N_4269,N_4342);
or U4980 (N_4980,N_4272,N_4499);
nor U4981 (N_4981,N_4192,N_4204);
nor U4982 (N_4982,N_4489,N_4075);
or U4983 (N_4983,N_4379,N_4357);
xnor U4984 (N_4984,N_4366,N_4312);
or U4985 (N_4985,N_4329,N_4036);
nand U4986 (N_4986,N_4328,N_4178);
nor U4987 (N_4987,N_4141,N_4418);
xor U4988 (N_4988,N_4044,N_4456);
nor U4989 (N_4989,N_4098,N_4494);
and U4990 (N_4990,N_4329,N_4296);
nand U4991 (N_4991,N_4098,N_4018);
nor U4992 (N_4992,N_4311,N_4181);
and U4993 (N_4993,N_4101,N_4343);
nand U4994 (N_4994,N_4264,N_4349);
or U4995 (N_4995,N_4248,N_4464);
nor U4996 (N_4996,N_4326,N_4174);
nand U4997 (N_4997,N_4492,N_4413);
and U4998 (N_4998,N_4260,N_4108);
and U4999 (N_4999,N_4261,N_4450);
and UO_0 (O_0,N_4633,N_4868);
nor UO_1 (O_1,N_4695,N_4942);
and UO_2 (O_2,N_4573,N_4660);
and UO_3 (O_3,N_4750,N_4933);
and UO_4 (O_4,N_4534,N_4953);
nand UO_5 (O_5,N_4693,N_4661);
nor UO_6 (O_6,N_4865,N_4882);
and UO_7 (O_7,N_4807,N_4637);
or UO_8 (O_8,N_4909,N_4675);
nor UO_9 (O_9,N_4884,N_4718);
or UO_10 (O_10,N_4649,N_4851);
nor UO_11 (O_11,N_4740,N_4617);
and UO_12 (O_12,N_4793,N_4559);
and UO_13 (O_13,N_4503,N_4611);
or UO_14 (O_14,N_4671,N_4749);
and UO_15 (O_15,N_4915,N_4704);
and UO_16 (O_16,N_4574,N_4841);
and UO_17 (O_17,N_4571,N_4701);
nor UO_18 (O_18,N_4791,N_4698);
and UO_19 (O_19,N_4855,N_4581);
nor UO_20 (O_20,N_4713,N_4993);
nand UO_21 (O_21,N_4619,N_4829);
nand UO_22 (O_22,N_4715,N_4759);
nand UO_23 (O_23,N_4557,N_4594);
nand UO_24 (O_24,N_4522,N_4625);
or UO_25 (O_25,N_4858,N_4586);
or UO_26 (O_26,N_4642,N_4958);
nand UO_27 (O_27,N_4732,N_4847);
nand UO_28 (O_28,N_4856,N_4945);
nand UO_29 (O_29,N_4610,N_4859);
nor UO_30 (O_30,N_4912,N_4919);
nor UO_31 (O_31,N_4816,N_4543);
or UO_32 (O_32,N_4954,N_4735);
and UO_33 (O_33,N_4795,N_4570);
and UO_34 (O_34,N_4881,N_4502);
or UO_35 (O_35,N_4639,N_4947);
nor UO_36 (O_36,N_4579,N_4827);
and UO_37 (O_37,N_4746,N_4836);
nor UO_38 (O_38,N_4777,N_4929);
or UO_39 (O_39,N_4553,N_4584);
nor UO_40 (O_40,N_4600,N_4688);
nor UO_41 (O_41,N_4897,N_4667);
nand UO_42 (O_42,N_4591,N_4950);
or UO_43 (O_43,N_4849,N_4900);
xor UO_44 (O_44,N_4870,N_4500);
or UO_45 (O_45,N_4853,N_4575);
nor UO_46 (O_46,N_4934,N_4566);
or UO_47 (O_47,N_4788,N_4833);
nand UO_48 (O_48,N_4668,N_4694);
xor UO_49 (O_49,N_4558,N_4869);
nand UO_50 (O_50,N_4938,N_4814);
nand UO_51 (O_51,N_4769,N_4602);
and UO_52 (O_52,N_4561,N_4647);
nand UO_53 (O_53,N_4648,N_4696);
and UO_54 (O_54,N_4968,N_4967);
nor UO_55 (O_55,N_4927,N_4507);
nand UO_56 (O_56,N_4519,N_4564);
nand UO_57 (O_57,N_4901,N_4775);
xor UO_58 (O_58,N_4813,N_4614);
nor UO_59 (O_59,N_4681,N_4665);
nor UO_60 (O_60,N_4944,N_4504);
nor UO_61 (O_61,N_4547,N_4666);
nand UO_62 (O_62,N_4823,N_4781);
nor UO_63 (O_63,N_4632,N_4555);
nor UO_64 (O_64,N_4726,N_4508);
xnor UO_65 (O_65,N_4772,N_4689);
and UO_66 (O_66,N_4634,N_4678);
or UO_67 (O_67,N_4982,N_4505);
or UO_68 (O_68,N_4866,N_4804);
nand UO_69 (O_69,N_4615,N_4976);
and UO_70 (O_70,N_4805,N_4748);
or UO_71 (O_71,N_4578,N_4757);
and UO_72 (O_72,N_4545,N_4518);
or UO_73 (O_73,N_4994,N_4810);
and UO_74 (O_74,N_4902,N_4623);
and UO_75 (O_75,N_4990,N_4532);
nor UO_76 (O_76,N_4593,N_4825);
nand UO_77 (O_77,N_4501,N_4939);
and UO_78 (O_78,N_4685,N_4935);
and UO_79 (O_79,N_4515,N_4984);
nand UO_80 (O_80,N_4562,N_4910);
nor UO_81 (O_81,N_4690,N_4747);
nand UO_82 (O_82,N_4554,N_4756);
nand UO_83 (O_83,N_4716,N_4708);
nand UO_84 (O_84,N_4659,N_4729);
and UO_85 (O_85,N_4991,N_4609);
nor UO_86 (O_86,N_4714,N_4636);
nand UO_87 (O_87,N_4758,N_4817);
nand UO_88 (O_88,N_4932,N_4686);
or UO_89 (O_89,N_4819,N_4645);
nand UO_90 (O_90,N_4673,N_4871);
and UO_91 (O_91,N_4974,N_4514);
or UO_92 (O_92,N_4630,N_4717);
or UO_93 (O_93,N_4620,N_4966);
nand UO_94 (O_94,N_4955,N_4525);
nor UO_95 (O_95,N_4771,N_4782);
nand UO_96 (O_96,N_4996,N_4551);
nor UO_97 (O_97,N_4962,N_4539);
nor UO_98 (O_98,N_4583,N_4899);
and UO_99 (O_99,N_4744,N_4755);
nor UO_100 (O_100,N_4510,N_4887);
or UO_101 (O_101,N_4808,N_4761);
nand UO_102 (O_102,N_4702,N_4700);
and UO_103 (O_103,N_4576,N_4784);
and UO_104 (O_104,N_4905,N_4618);
nand UO_105 (O_105,N_4896,N_4520);
or UO_106 (O_106,N_4957,N_4831);
nor UO_107 (O_107,N_4533,N_4995);
nor UO_108 (O_108,N_4926,N_4707);
nand UO_109 (O_109,N_4780,N_4509);
and UO_110 (O_110,N_4542,N_4628);
nand UO_111 (O_111,N_4592,N_4923);
and UO_112 (O_112,N_4567,N_4683);
and UO_113 (O_113,N_4658,N_4589);
or UO_114 (O_114,N_4809,N_4980);
nor UO_115 (O_115,N_4890,N_4692);
nor UO_116 (O_116,N_4960,N_4821);
and UO_117 (O_117,N_4601,N_4986);
nor UO_118 (O_118,N_4604,N_4722);
and UO_119 (O_119,N_4754,N_4674);
nor UO_120 (O_120,N_4940,N_4530);
or UO_121 (O_121,N_4842,N_4641);
and UO_122 (O_122,N_4977,N_4834);
or UO_123 (O_123,N_4599,N_4796);
nor UO_124 (O_124,N_4513,N_4626);
or UO_125 (O_125,N_4965,N_4768);
nor UO_126 (O_126,N_4656,N_4818);
nor UO_127 (O_127,N_4911,N_4999);
nand UO_128 (O_128,N_4652,N_4751);
nor UO_129 (O_129,N_4850,N_4907);
or UO_130 (O_130,N_4998,N_4811);
nand UO_131 (O_131,N_4767,N_4638);
or UO_132 (O_132,N_4789,N_4597);
nand UO_133 (O_133,N_4846,N_4948);
nand UO_134 (O_134,N_4569,N_4843);
or UO_135 (O_135,N_4725,N_4981);
nor UO_136 (O_136,N_4800,N_4529);
nor UO_137 (O_137,N_4541,N_4627);
and UO_138 (O_138,N_4875,N_4524);
or UO_139 (O_139,N_4941,N_4580);
nand UO_140 (O_140,N_4724,N_4745);
or UO_141 (O_141,N_4760,N_4640);
and UO_142 (O_142,N_4663,N_4815);
xnor UO_143 (O_143,N_4864,N_4587);
or UO_144 (O_144,N_4550,N_4526);
and UO_145 (O_145,N_4709,N_4839);
nand UO_146 (O_146,N_4613,N_4528);
and UO_147 (O_147,N_4883,N_4824);
nor UO_148 (O_148,N_4585,N_4785);
or UO_149 (O_149,N_4979,N_4635);
nor UO_150 (O_150,N_4798,N_4914);
or UO_151 (O_151,N_4738,N_4787);
nor UO_152 (O_152,N_4603,N_4874);
nand UO_153 (O_153,N_4572,N_4535);
nor UO_154 (O_154,N_4721,N_4873);
and UO_155 (O_155,N_4857,N_4605);
nand UO_156 (O_156,N_4790,N_4538);
and UO_157 (O_157,N_4672,N_4770);
or UO_158 (O_158,N_4906,N_4959);
nor UO_159 (O_159,N_4920,N_4854);
nand UO_160 (O_160,N_4983,N_4973);
or UO_161 (O_161,N_4844,N_4670);
nor UO_162 (O_162,N_4560,N_4891);
nand UO_163 (O_163,N_4898,N_4917);
nor UO_164 (O_164,N_4679,N_4943);
and UO_165 (O_165,N_4728,N_4631);
nor UO_166 (O_166,N_4931,N_4852);
xnor UO_167 (O_167,N_4963,N_4680);
nand UO_168 (O_168,N_4616,N_4886);
nor UO_169 (O_169,N_4687,N_4621);
and UO_170 (O_170,N_4826,N_4964);
or UO_171 (O_171,N_4880,N_4622);
nor UO_172 (O_172,N_4877,N_4565);
nor UO_173 (O_173,N_4650,N_4992);
nor UO_174 (O_174,N_4512,N_4664);
or UO_175 (O_175,N_4516,N_4588);
nor UO_176 (O_176,N_4764,N_4765);
or UO_177 (O_177,N_4822,N_4792);
nor UO_178 (O_178,N_4606,N_4946);
and UO_179 (O_179,N_4506,N_4766);
xnor UO_180 (O_180,N_4969,N_4916);
nand UO_181 (O_181,N_4568,N_4997);
or UO_182 (O_182,N_4577,N_4861);
and UO_183 (O_183,N_4918,N_4802);
nand UO_184 (O_184,N_4596,N_4952);
or UO_185 (O_185,N_4607,N_4972);
nor UO_186 (O_186,N_4903,N_4803);
or UO_187 (O_187,N_4753,N_4951);
nor UO_188 (O_188,N_4863,N_4786);
nand UO_189 (O_189,N_4908,N_4985);
and UO_190 (O_190,N_4876,N_4527);
and UO_191 (O_191,N_4676,N_4723);
and UO_192 (O_192,N_4949,N_4904);
nor UO_193 (O_193,N_4970,N_4537);
nand UO_194 (O_194,N_4889,N_4736);
or UO_195 (O_195,N_4894,N_4536);
nand UO_196 (O_196,N_4895,N_4867);
or UO_197 (O_197,N_4521,N_4752);
nor UO_198 (O_198,N_4921,N_4598);
or UO_199 (O_199,N_4860,N_4651);
xor UO_200 (O_200,N_4608,N_4511);
or UO_201 (O_201,N_4779,N_4892);
nand UO_202 (O_202,N_4662,N_4727);
nor UO_203 (O_203,N_4544,N_4936);
or UO_204 (O_204,N_4989,N_4540);
or UO_205 (O_205,N_4832,N_4654);
nor UO_206 (O_206,N_4978,N_4739);
nor UO_207 (O_207,N_4697,N_4848);
and UO_208 (O_208,N_4595,N_4612);
or UO_209 (O_209,N_4878,N_4523);
and UO_210 (O_210,N_4743,N_4806);
nand UO_211 (O_211,N_4922,N_4799);
nand UO_212 (O_212,N_4763,N_4961);
nand UO_213 (O_213,N_4655,N_4776);
or UO_214 (O_214,N_4699,N_4705);
nor UO_215 (O_215,N_4517,N_4924);
nor UO_216 (O_216,N_4644,N_4837);
nand UO_217 (O_217,N_4590,N_4975);
and UO_218 (O_218,N_4987,N_4773);
and UO_219 (O_219,N_4937,N_4731);
nand UO_220 (O_220,N_4872,N_4734);
or UO_221 (O_221,N_4531,N_4712);
and UO_222 (O_222,N_4719,N_4893);
and UO_223 (O_223,N_4925,N_4838);
or UO_224 (O_224,N_4552,N_4742);
nor UO_225 (O_225,N_4885,N_4971);
nor UO_226 (O_226,N_4956,N_4624);
or UO_227 (O_227,N_4930,N_4774);
and UO_228 (O_228,N_4711,N_4684);
and UO_229 (O_229,N_4862,N_4794);
or UO_230 (O_230,N_4546,N_4646);
nor UO_231 (O_231,N_4828,N_4548);
and UO_232 (O_232,N_4720,N_4778);
nor UO_233 (O_233,N_4653,N_4888);
and UO_234 (O_234,N_4988,N_4783);
or UO_235 (O_235,N_4741,N_4710);
nand UO_236 (O_236,N_4913,N_4703);
nor UO_237 (O_237,N_4812,N_4691);
or UO_238 (O_238,N_4643,N_4730);
nor UO_239 (O_239,N_4835,N_4556);
nand UO_240 (O_240,N_4928,N_4629);
nor UO_241 (O_241,N_4549,N_4879);
nor UO_242 (O_242,N_4682,N_4733);
and UO_243 (O_243,N_4830,N_4797);
nor UO_244 (O_244,N_4669,N_4677);
and UO_245 (O_245,N_4706,N_4737);
nor UO_246 (O_246,N_4762,N_4840);
nor UO_247 (O_247,N_4820,N_4801);
nand UO_248 (O_248,N_4657,N_4845);
or UO_249 (O_249,N_4563,N_4582);
or UO_250 (O_250,N_4582,N_4864);
and UO_251 (O_251,N_4722,N_4978);
nand UO_252 (O_252,N_4775,N_4958);
nand UO_253 (O_253,N_4755,N_4724);
nor UO_254 (O_254,N_4735,N_4803);
and UO_255 (O_255,N_4571,N_4523);
and UO_256 (O_256,N_4619,N_4689);
and UO_257 (O_257,N_4727,N_4621);
nand UO_258 (O_258,N_4749,N_4728);
and UO_259 (O_259,N_4739,N_4846);
and UO_260 (O_260,N_4925,N_4563);
or UO_261 (O_261,N_4805,N_4954);
and UO_262 (O_262,N_4547,N_4786);
and UO_263 (O_263,N_4705,N_4694);
nand UO_264 (O_264,N_4721,N_4675);
or UO_265 (O_265,N_4951,N_4974);
xnor UO_266 (O_266,N_4544,N_4683);
nand UO_267 (O_267,N_4883,N_4540);
or UO_268 (O_268,N_4671,N_4982);
and UO_269 (O_269,N_4967,N_4784);
or UO_270 (O_270,N_4809,N_4855);
nand UO_271 (O_271,N_4998,N_4762);
and UO_272 (O_272,N_4556,N_4862);
nor UO_273 (O_273,N_4778,N_4685);
and UO_274 (O_274,N_4505,N_4868);
nor UO_275 (O_275,N_4516,N_4773);
nand UO_276 (O_276,N_4732,N_4694);
nand UO_277 (O_277,N_4700,N_4630);
nor UO_278 (O_278,N_4654,N_4509);
nand UO_279 (O_279,N_4559,N_4813);
or UO_280 (O_280,N_4814,N_4525);
nor UO_281 (O_281,N_4633,N_4528);
nor UO_282 (O_282,N_4534,N_4582);
and UO_283 (O_283,N_4746,N_4955);
or UO_284 (O_284,N_4806,N_4527);
nor UO_285 (O_285,N_4568,N_4989);
xor UO_286 (O_286,N_4562,N_4823);
and UO_287 (O_287,N_4977,N_4686);
and UO_288 (O_288,N_4701,N_4949);
nand UO_289 (O_289,N_4640,N_4928);
and UO_290 (O_290,N_4865,N_4709);
nor UO_291 (O_291,N_4606,N_4679);
and UO_292 (O_292,N_4639,N_4608);
nand UO_293 (O_293,N_4707,N_4777);
xnor UO_294 (O_294,N_4960,N_4866);
and UO_295 (O_295,N_4943,N_4986);
or UO_296 (O_296,N_4649,N_4645);
and UO_297 (O_297,N_4905,N_4685);
and UO_298 (O_298,N_4581,N_4879);
nand UO_299 (O_299,N_4967,N_4921);
and UO_300 (O_300,N_4697,N_4723);
nor UO_301 (O_301,N_4661,N_4777);
nand UO_302 (O_302,N_4665,N_4973);
and UO_303 (O_303,N_4619,N_4983);
or UO_304 (O_304,N_4943,N_4841);
and UO_305 (O_305,N_4759,N_4972);
and UO_306 (O_306,N_4681,N_4909);
nor UO_307 (O_307,N_4886,N_4521);
nand UO_308 (O_308,N_4967,N_4945);
or UO_309 (O_309,N_4613,N_4770);
and UO_310 (O_310,N_4574,N_4803);
or UO_311 (O_311,N_4778,N_4838);
nor UO_312 (O_312,N_4963,N_4946);
or UO_313 (O_313,N_4600,N_4978);
or UO_314 (O_314,N_4692,N_4794);
nand UO_315 (O_315,N_4531,N_4823);
and UO_316 (O_316,N_4583,N_4819);
and UO_317 (O_317,N_4972,N_4638);
or UO_318 (O_318,N_4874,N_4760);
nor UO_319 (O_319,N_4504,N_4520);
or UO_320 (O_320,N_4843,N_4667);
or UO_321 (O_321,N_4920,N_4712);
or UO_322 (O_322,N_4825,N_4543);
nand UO_323 (O_323,N_4818,N_4752);
and UO_324 (O_324,N_4662,N_4691);
and UO_325 (O_325,N_4746,N_4613);
nor UO_326 (O_326,N_4754,N_4601);
and UO_327 (O_327,N_4817,N_4982);
nand UO_328 (O_328,N_4606,N_4865);
nor UO_329 (O_329,N_4602,N_4724);
nor UO_330 (O_330,N_4534,N_4644);
nor UO_331 (O_331,N_4579,N_4523);
or UO_332 (O_332,N_4992,N_4613);
nor UO_333 (O_333,N_4864,N_4859);
or UO_334 (O_334,N_4542,N_4761);
or UO_335 (O_335,N_4926,N_4805);
nor UO_336 (O_336,N_4557,N_4694);
or UO_337 (O_337,N_4508,N_4874);
nand UO_338 (O_338,N_4659,N_4676);
nor UO_339 (O_339,N_4997,N_4827);
or UO_340 (O_340,N_4909,N_4657);
or UO_341 (O_341,N_4960,N_4764);
or UO_342 (O_342,N_4810,N_4721);
nand UO_343 (O_343,N_4570,N_4524);
and UO_344 (O_344,N_4528,N_4904);
and UO_345 (O_345,N_4920,N_4771);
xor UO_346 (O_346,N_4940,N_4723);
or UO_347 (O_347,N_4766,N_4557);
or UO_348 (O_348,N_4731,N_4594);
nor UO_349 (O_349,N_4911,N_4939);
nand UO_350 (O_350,N_4864,N_4735);
nor UO_351 (O_351,N_4770,N_4954);
and UO_352 (O_352,N_4922,N_4611);
nand UO_353 (O_353,N_4762,N_4804);
and UO_354 (O_354,N_4753,N_4570);
nand UO_355 (O_355,N_4774,N_4653);
and UO_356 (O_356,N_4706,N_4651);
nor UO_357 (O_357,N_4652,N_4665);
nor UO_358 (O_358,N_4747,N_4621);
or UO_359 (O_359,N_4727,N_4533);
and UO_360 (O_360,N_4838,N_4535);
xnor UO_361 (O_361,N_4577,N_4909);
nor UO_362 (O_362,N_4883,N_4610);
nand UO_363 (O_363,N_4624,N_4872);
nor UO_364 (O_364,N_4586,N_4975);
or UO_365 (O_365,N_4694,N_4576);
nor UO_366 (O_366,N_4719,N_4723);
nand UO_367 (O_367,N_4600,N_4566);
nand UO_368 (O_368,N_4923,N_4944);
nand UO_369 (O_369,N_4724,N_4608);
or UO_370 (O_370,N_4532,N_4744);
nor UO_371 (O_371,N_4785,N_4939);
nor UO_372 (O_372,N_4814,N_4769);
and UO_373 (O_373,N_4616,N_4709);
nand UO_374 (O_374,N_4983,N_4738);
nor UO_375 (O_375,N_4525,N_4835);
nor UO_376 (O_376,N_4562,N_4839);
nor UO_377 (O_377,N_4573,N_4929);
and UO_378 (O_378,N_4670,N_4953);
nand UO_379 (O_379,N_4883,N_4865);
and UO_380 (O_380,N_4901,N_4822);
nand UO_381 (O_381,N_4938,N_4877);
and UO_382 (O_382,N_4740,N_4813);
and UO_383 (O_383,N_4979,N_4934);
or UO_384 (O_384,N_4841,N_4752);
or UO_385 (O_385,N_4799,N_4894);
or UO_386 (O_386,N_4708,N_4600);
nand UO_387 (O_387,N_4676,N_4539);
nor UO_388 (O_388,N_4858,N_4853);
or UO_389 (O_389,N_4728,N_4648);
and UO_390 (O_390,N_4769,N_4723);
and UO_391 (O_391,N_4912,N_4648);
and UO_392 (O_392,N_4505,N_4561);
nor UO_393 (O_393,N_4886,N_4636);
nor UO_394 (O_394,N_4999,N_4937);
or UO_395 (O_395,N_4754,N_4637);
or UO_396 (O_396,N_4938,N_4830);
and UO_397 (O_397,N_4619,N_4546);
or UO_398 (O_398,N_4589,N_4619);
nand UO_399 (O_399,N_4708,N_4776);
or UO_400 (O_400,N_4639,N_4641);
nand UO_401 (O_401,N_4738,N_4679);
nand UO_402 (O_402,N_4606,N_4611);
xor UO_403 (O_403,N_4924,N_4721);
and UO_404 (O_404,N_4735,N_4897);
and UO_405 (O_405,N_4609,N_4864);
nor UO_406 (O_406,N_4725,N_4694);
and UO_407 (O_407,N_4653,N_4990);
nand UO_408 (O_408,N_4939,N_4520);
nor UO_409 (O_409,N_4858,N_4634);
and UO_410 (O_410,N_4532,N_4794);
nor UO_411 (O_411,N_4988,N_4976);
nand UO_412 (O_412,N_4948,N_4714);
and UO_413 (O_413,N_4821,N_4613);
or UO_414 (O_414,N_4767,N_4522);
nand UO_415 (O_415,N_4820,N_4535);
nor UO_416 (O_416,N_4967,N_4820);
nand UO_417 (O_417,N_4854,N_4849);
nand UO_418 (O_418,N_4872,N_4687);
and UO_419 (O_419,N_4973,N_4937);
or UO_420 (O_420,N_4732,N_4717);
and UO_421 (O_421,N_4582,N_4971);
or UO_422 (O_422,N_4784,N_4529);
or UO_423 (O_423,N_4691,N_4661);
nor UO_424 (O_424,N_4738,N_4935);
nand UO_425 (O_425,N_4935,N_4602);
or UO_426 (O_426,N_4865,N_4630);
and UO_427 (O_427,N_4953,N_4926);
or UO_428 (O_428,N_4894,N_4863);
nor UO_429 (O_429,N_4816,N_4609);
nand UO_430 (O_430,N_4907,N_4545);
nand UO_431 (O_431,N_4954,N_4723);
and UO_432 (O_432,N_4753,N_4908);
and UO_433 (O_433,N_4637,N_4543);
and UO_434 (O_434,N_4932,N_4798);
or UO_435 (O_435,N_4534,N_4572);
nor UO_436 (O_436,N_4940,N_4933);
nand UO_437 (O_437,N_4816,N_4571);
and UO_438 (O_438,N_4788,N_4762);
nor UO_439 (O_439,N_4886,N_4554);
nor UO_440 (O_440,N_4945,N_4543);
and UO_441 (O_441,N_4831,N_4854);
nand UO_442 (O_442,N_4669,N_4782);
nor UO_443 (O_443,N_4610,N_4797);
or UO_444 (O_444,N_4936,N_4560);
or UO_445 (O_445,N_4949,N_4623);
nand UO_446 (O_446,N_4569,N_4945);
or UO_447 (O_447,N_4767,N_4604);
nand UO_448 (O_448,N_4571,N_4587);
xor UO_449 (O_449,N_4761,N_4971);
and UO_450 (O_450,N_4698,N_4958);
nor UO_451 (O_451,N_4986,N_4759);
nand UO_452 (O_452,N_4638,N_4662);
nand UO_453 (O_453,N_4942,N_4911);
and UO_454 (O_454,N_4811,N_4735);
nand UO_455 (O_455,N_4978,N_4569);
or UO_456 (O_456,N_4908,N_4987);
nand UO_457 (O_457,N_4716,N_4916);
and UO_458 (O_458,N_4579,N_4807);
nor UO_459 (O_459,N_4710,N_4505);
nor UO_460 (O_460,N_4666,N_4530);
and UO_461 (O_461,N_4820,N_4979);
nor UO_462 (O_462,N_4755,N_4939);
and UO_463 (O_463,N_4932,N_4958);
or UO_464 (O_464,N_4617,N_4755);
nor UO_465 (O_465,N_4778,N_4875);
and UO_466 (O_466,N_4756,N_4535);
and UO_467 (O_467,N_4692,N_4695);
or UO_468 (O_468,N_4793,N_4575);
and UO_469 (O_469,N_4991,N_4993);
and UO_470 (O_470,N_4924,N_4836);
or UO_471 (O_471,N_4672,N_4608);
or UO_472 (O_472,N_4507,N_4599);
and UO_473 (O_473,N_4857,N_4863);
and UO_474 (O_474,N_4619,N_4569);
or UO_475 (O_475,N_4811,N_4537);
nand UO_476 (O_476,N_4774,N_4564);
nor UO_477 (O_477,N_4971,N_4651);
and UO_478 (O_478,N_4775,N_4776);
or UO_479 (O_479,N_4850,N_4897);
and UO_480 (O_480,N_4857,N_4781);
nor UO_481 (O_481,N_4701,N_4572);
nor UO_482 (O_482,N_4686,N_4846);
and UO_483 (O_483,N_4990,N_4752);
nand UO_484 (O_484,N_4766,N_4560);
nor UO_485 (O_485,N_4625,N_4541);
xor UO_486 (O_486,N_4579,N_4837);
and UO_487 (O_487,N_4881,N_4648);
nand UO_488 (O_488,N_4681,N_4655);
nor UO_489 (O_489,N_4868,N_4732);
nor UO_490 (O_490,N_4652,N_4703);
nand UO_491 (O_491,N_4581,N_4565);
nor UO_492 (O_492,N_4884,N_4557);
nand UO_493 (O_493,N_4778,N_4914);
nand UO_494 (O_494,N_4682,N_4582);
nand UO_495 (O_495,N_4658,N_4688);
nand UO_496 (O_496,N_4983,N_4551);
and UO_497 (O_497,N_4823,N_4689);
nor UO_498 (O_498,N_4751,N_4882);
nor UO_499 (O_499,N_4554,N_4855);
and UO_500 (O_500,N_4671,N_4691);
xor UO_501 (O_501,N_4745,N_4935);
nor UO_502 (O_502,N_4504,N_4689);
nand UO_503 (O_503,N_4574,N_4875);
or UO_504 (O_504,N_4617,N_4897);
nor UO_505 (O_505,N_4505,N_4636);
and UO_506 (O_506,N_4921,N_4594);
and UO_507 (O_507,N_4637,N_4783);
and UO_508 (O_508,N_4647,N_4975);
or UO_509 (O_509,N_4865,N_4642);
nand UO_510 (O_510,N_4904,N_4682);
nor UO_511 (O_511,N_4614,N_4812);
or UO_512 (O_512,N_4794,N_4866);
nor UO_513 (O_513,N_4764,N_4683);
nand UO_514 (O_514,N_4749,N_4503);
nor UO_515 (O_515,N_4693,N_4717);
nor UO_516 (O_516,N_4753,N_4596);
nand UO_517 (O_517,N_4738,N_4696);
nand UO_518 (O_518,N_4532,N_4906);
nor UO_519 (O_519,N_4757,N_4504);
nor UO_520 (O_520,N_4768,N_4545);
nand UO_521 (O_521,N_4501,N_4840);
nor UO_522 (O_522,N_4622,N_4912);
nand UO_523 (O_523,N_4524,N_4655);
and UO_524 (O_524,N_4856,N_4548);
or UO_525 (O_525,N_4907,N_4524);
or UO_526 (O_526,N_4561,N_4735);
nand UO_527 (O_527,N_4793,N_4606);
or UO_528 (O_528,N_4760,N_4576);
nand UO_529 (O_529,N_4998,N_4779);
nor UO_530 (O_530,N_4652,N_4585);
nand UO_531 (O_531,N_4790,N_4922);
nor UO_532 (O_532,N_4854,N_4751);
and UO_533 (O_533,N_4846,N_4910);
and UO_534 (O_534,N_4677,N_4631);
nor UO_535 (O_535,N_4902,N_4875);
and UO_536 (O_536,N_4896,N_4899);
and UO_537 (O_537,N_4804,N_4705);
nor UO_538 (O_538,N_4900,N_4577);
nor UO_539 (O_539,N_4794,N_4786);
or UO_540 (O_540,N_4868,N_4884);
nor UO_541 (O_541,N_4647,N_4989);
nor UO_542 (O_542,N_4690,N_4603);
and UO_543 (O_543,N_4949,N_4809);
and UO_544 (O_544,N_4595,N_4645);
or UO_545 (O_545,N_4954,N_4556);
or UO_546 (O_546,N_4622,N_4803);
nand UO_547 (O_547,N_4781,N_4574);
nand UO_548 (O_548,N_4696,N_4632);
nand UO_549 (O_549,N_4855,N_4576);
or UO_550 (O_550,N_4711,N_4993);
and UO_551 (O_551,N_4747,N_4956);
nand UO_552 (O_552,N_4607,N_4756);
and UO_553 (O_553,N_4591,N_4883);
nor UO_554 (O_554,N_4764,N_4657);
or UO_555 (O_555,N_4504,N_4710);
nor UO_556 (O_556,N_4998,N_4661);
nor UO_557 (O_557,N_4892,N_4947);
nor UO_558 (O_558,N_4562,N_4686);
nor UO_559 (O_559,N_4828,N_4533);
and UO_560 (O_560,N_4922,N_4831);
nor UO_561 (O_561,N_4633,N_4846);
nor UO_562 (O_562,N_4623,N_4598);
nand UO_563 (O_563,N_4898,N_4726);
nand UO_564 (O_564,N_4935,N_4585);
or UO_565 (O_565,N_4640,N_4904);
nor UO_566 (O_566,N_4927,N_4672);
nand UO_567 (O_567,N_4809,N_4986);
nor UO_568 (O_568,N_4974,N_4671);
nor UO_569 (O_569,N_4893,N_4535);
nor UO_570 (O_570,N_4673,N_4682);
or UO_571 (O_571,N_4616,N_4888);
and UO_572 (O_572,N_4988,N_4746);
and UO_573 (O_573,N_4829,N_4547);
or UO_574 (O_574,N_4678,N_4509);
nand UO_575 (O_575,N_4942,N_4751);
nand UO_576 (O_576,N_4619,N_4824);
and UO_577 (O_577,N_4624,N_4515);
nor UO_578 (O_578,N_4765,N_4645);
nand UO_579 (O_579,N_4846,N_4967);
or UO_580 (O_580,N_4648,N_4942);
nor UO_581 (O_581,N_4915,N_4790);
and UO_582 (O_582,N_4977,N_4701);
nor UO_583 (O_583,N_4841,N_4552);
nor UO_584 (O_584,N_4864,N_4783);
nand UO_585 (O_585,N_4535,N_4560);
and UO_586 (O_586,N_4672,N_4940);
nor UO_587 (O_587,N_4917,N_4657);
nand UO_588 (O_588,N_4757,N_4964);
nand UO_589 (O_589,N_4701,N_4980);
nor UO_590 (O_590,N_4580,N_4745);
nand UO_591 (O_591,N_4950,N_4997);
and UO_592 (O_592,N_4995,N_4615);
nor UO_593 (O_593,N_4519,N_4509);
and UO_594 (O_594,N_4999,N_4924);
or UO_595 (O_595,N_4542,N_4503);
and UO_596 (O_596,N_4705,N_4695);
nor UO_597 (O_597,N_4923,N_4606);
nor UO_598 (O_598,N_4752,N_4608);
nand UO_599 (O_599,N_4931,N_4855);
nand UO_600 (O_600,N_4795,N_4550);
or UO_601 (O_601,N_4563,N_4769);
nand UO_602 (O_602,N_4913,N_4859);
nand UO_603 (O_603,N_4868,N_4503);
nor UO_604 (O_604,N_4624,N_4902);
or UO_605 (O_605,N_4946,N_4540);
nor UO_606 (O_606,N_4905,N_4750);
nand UO_607 (O_607,N_4527,N_4742);
and UO_608 (O_608,N_4978,N_4964);
or UO_609 (O_609,N_4690,N_4809);
nand UO_610 (O_610,N_4628,N_4537);
and UO_611 (O_611,N_4863,N_4747);
and UO_612 (O_612,N_4578,N_4835);
and UO_613 (O_613,N_4894,N_4972);
nor UO_614 (O_614,N_4599,N_4605);
nor UO_615 (O_615,N_4845,N_4586);
and UO_616 (O_616,N_4919,N_4810);
and UO_617 (O_617,N_4574,N_4512);
nor UO_618 (O_618,N_4949,N_4650);
nand UO_619 (O_619,N_4777,N_4564);
or UO_620 (O_620,N_4632,N_4911);
nand UO_621 (O_621,N_4733,N_4784);
or UO_622 (O_622,N_4759,N_4766);
or UO_623 (O_623,N_4900,N_4717);
and UO_624 (O_624,N_4881,N_4972);
or UO_625 (O_625,N_4654,N_4837);
and UO_626 (O_626,N_4663,N_4682);
or UO_627 (O_627,N_4645,N_4643);
or UO_628 (O_628,N_4713,N_4610);
and UO_629 (O_629,N_4889,N_4563);
and UO_630 (O_630,N_4540,N_4952);
nor UO_631 (O_631,N_4975,N_4539);
or UO_632 (O_632,N_4911,N_4912);
or UO_633 (O_633,N_4596,N_4545);
nand UO_634 (O_634,N_4917,N_4773);
nor UO_635 (O_635,N_4770,N_4525);
and UO_636 (O_636,N_4826,N_4951);
nand UO_637 (O_637,N_4590,N_4645);
nand UO_638 (O_638,N_4573,N_4706);
and UO_639 (O_639,N_4911,N_4699);
or UO_640 (O_640,N_4773,N_4947);
nor UO_641 (O_641,N_4996,N_4841);
nor UO_642 (O_642,N_4694,N_4936);
and UO_643 (O_643,N_4961,N_4979);
nor UO_644 (O_644,N_4937,N_4659);
or UO_645 (O_645,N_4913,N_4515);
nand UO_646 (O_646,N_4828,N_4856);
or UO_647 (O_647,N_4886,N_4813);
nor UO_648 (O_648,N_4547,N_4821);
nor UO_649 (O_649,N_4962,N_4870);
nand UO_650 (O_650,N_4656,N_4634);
and UO_651 (O_651,N_4992,N_4726);
nor UO_652 (O_652,N_4525,N_4613);
nor UO_653 (O_653,N_4828,N_4696);
nand UO_654 (O_654,N_4653,N_4732);
or UO_655 (O_655,N_4522,N_4516);
and UO_656 (O_656,N_4944,N_4755);
or UO_657 (O_657,N_4537,N_4855);
or UO_658 (O_658,N_4966,N_4600);
or UO_659 (O_659,N_4698,N_4682);
nor UO_660 (O_660,N_4823,N_4969);
nand UO_661 (O_661,N_4978,N_4522);
nor UO_662 (O_662,N_4656,N_4915);
nand UO_663 (O_663,N_4866,N_4861);
or UO_664 (O_664,N_4867,N_4622);
or UO_665 (O_665,N_4876,N_4586);
and UO_666 (O_666,N_4774,N_4685);
and UO_667 (O_667,N_4933,N_4587);
nor UO_668 (O_668,N_4868,N_4821);
nand UO_669 (O_669,N_4881,N_4927);
nand UO_670 (O_670,N_4943,N_4599);
and UO_671 (O_671,N_4992,N_4512);
and UO_672 (O_672,N_4854,N_4762);
and UO_673 (O_673,N_4920,N_4698);
nand UO_674 (O_674,N_4550,N_4660);
or UO_675 (O_675,N_4768,N_4708);
or UO_676 (O_676,N_4543,N_4781);
or UO_677 (O_677,N_4819,N_4579);
nand UO_678 (O_678,N_4546,N_4782);
nand UO_679 (O_679,N_4562,N_4767);
nor UO_680 (O_680,N_4940,N_4863);
and UO_681 (O_681,N_4514,N_4982);
nor UO_682 (O_682,N_4506,N_4653);
nand UO_683 (O_683,N_4722,N_4780);
nor UO_684 (O_684,N_4780,N_4597);
and UO_685 (O_685,N_4570,N_4594);
or UO_686 (O_686,N_4788,N_4823);
and UO_687 (O_687,N_4500,N_4671);
nor UO_688 (O_688,N_4711,N_4562);
nand UO_689 (O_689,N_4687,N_4863);
or UO_690 (O_690,N_4882,N_4929);
and UO_691 (O_691,N_4874,N_4988);
nand UO_692 (O_692,N_4745,N_4945);
and UO_693 (O_693,N_4724,N_4729);
nand UO_694 (O_694,N_4603,N_4980);
nor UO_695 (O_695,N_4935,N_4605);
xor UO_696 (O_696,N_4578,N_4561);
and UO_697 (O_697,N_4692,N_4840);
or UO_698 (O_698,N_4659,N_4758);
nor UO_699 (O_699,N_4758,N_4975);
nand UO_700 (O_700,N_4518,N_4656);
nor UO_701 (O_701,N_4847,N_4551);
or UO_702 (O_702,N_4764,N_4620);
nor UO_703 (O_703,N_4602,N_4942);
nand UO_704 (O_704,N_4860,N_4755);
nand UO_705 (O_705,N_4795,N_4894);
nor UO_706 (O_706,N_4782,N_4549);
or UO_707 (O_707,N_4947,N_4875);
nand UO_708 (O_708,N_4703,N_4590);
nor UO_709 (O_709,N_4935,N_4831);
and UO_710 (O_710,N_4593,N_4985);
nand UO_711 (O_711,N_4610,N_4594);
and UO_712 (O_712,N_4740,N_4551);
and UO_713 (O_713,N_4992,N_4940);
and UO_714 (O_714,N_4806,N_4908);
nor UO_715 (O_715,N_4833,N_4978);
and UO_716 (O_716,N_4843,N_4940);
nor UO_717 (O_717,N_4517,N_4679);
nand UO_718 (O_718,N_4814,N_4936);
and UO_719 (O_719,N_4535,N_4556);
nor UO_720 (O_720,N_4847,N_4502);
and UO_721 (O_721,N_4559,N_4535);
or UO_722 (O_722,N_4821,N_4701);
and UO_723 (O_723,N_4998,N_4502);
nand UO_724 (O_724,N_4888,N_4679);
nor UO_725 (O_725,N_4640,N_4811);
or UO_726 (O_726,N_4933,N_4614);
and UO_727 (O_727,N_4844,N_4930);
nand UO_728 (O_728,N_4832,N_4798);
nand UO_729 (O_729,N_4968,N_4879);
nand UO_730 (O_730,N_4992,N_4709);
nor UO_731 (O_731,N_4662,N_4696);
or UO_732 (O_732,N_4778,N_4799);
or UO_733 (O_733,N_4560,N_4688);
or UO_734 (O_734,N_4744,N_4980);
nand UO_735 (O_735,N_4857,N_4669);
and UO_736 (O_736,N_4811,N_4577);
and UO_737 (O_737,N_4874,N_4940);
and UO_738 (O_738,N_4568,N_4561);
nand UO_739 (O_739,N_4695,N_4501);
nor UO_740 (O_740,N_4959,N_4773);
nor UO_741 (O_741,N_4537,N_4863);
nor UO_742 (O_742,N_4708,N_4820);
and UO_743 (O_743,N_4578,N_4618);
and UO_744 (O_744,N_4939,N_4760);
and UO_745 (O_745,N_4726,N_4924);
nand UO_746 (O_746,N_4934,N_4570);
nor UO_747 (O_747,N_4570,N_4863);
and UO_748 (O_748,N_4500,N_4812);
nor UO_749 (O_749,N_4777,N_4673);
nor UO_750 (O_750,N_4633,N_4651);
nor UO_751 (O_751,N_4912,N_4963);
and UO_752 (O_752,N_4704,N_4846);
and UO_753 (O_753,N_4925,N_4839);
and UO_754 (O_754,N_4647,N_4858);
or UO_755 (O_755,N_4911,N_4757);
or UO_756 (O_756,N_4520,N_4923);
nand UO_757 (O_757,N_4886,N_4802);
and UO_758 (O_758,N_4847,N_4887);
nor UO_759 (O_759,N_4797,N_4857);
or UO_760 (O_760,N_4677,N_4589);
or UO_761 (O_761,N_4847,N_4637);
nor UO_762 (O_762,N_4719,N_4957);
and UO_763 (O_763,N_4652,N_4627);
nor UO_764 (O_764,N_4555,N_4836);
and UO_765 (O_765,N_4888,N_4538);
and UO_766 (O_766,N_4966,N_4627);
nand UO_767 (O_767,N_4977,N_4945);
xnor UO_768 (O_768,N_4882,N_4660);
nand UO_769 (O_769,N_4507,N_4659);
nand UO_770 (O_770,N_4895,N_4775);
nor UO_771 (O_771,N_4689,N_4520);
nand UO_772 (O_772,N_4599,N_4645);
and UO_773 (O_773,N_4734,N_4829);
nor UO_774 (O_774,N_4900,N_4897);
nand UO_775 (O_775,N_4756,N_4652);
nand UO_776 (O_776,N_4613,N_4854);
and UO_777 (O_777,N_4624,N_4771);
and UO_778 (O_778,N_4924,N_4553);
nand UO_779 (O_779,N_4694,N_4624);
and UO_780 (O_780,N_4856,N_4632);
and UO_781 (O_781,N_4569,N_4920);
or UO_782 (O_782,N_4980,N_4743);
nor UO_783 (O_783,N_4724,N_4691);
nor UO_784 (O_784,N_4813,N_4549);
and UO_785 (O_785,N_4683,N_4581);
and UO_786 (O_786,N_4839,N_4796);
nand UO_787 (O_787,N_4504,N_4700);
nor UO_788 (O_788,N_4913,N_4506);
nand UO_789 (O_789,N_4620,N_4927);
and UO_790 (O_790,N_4656,N_4566);
or UO_791 (O_791,N_4941,N_4712);
and UO_792 (O_792,N_4642,N_4632);
nand UO_793 (O_793,N_4951,N_4803);
and UO_794 (O_794,N_4780,N_4671);
nand UO_795 (O_795,N_4881,N_4669);
and UO_796 (O_796,N_4516,N_4730);
xor UO_797 (O_797,N_4615,N_4957);
nand UO_798 (O_798,N_4710,N_4862);
nand UO_799 (O_799,N_4860,N_4717);
nand UO_800 (O_800,N_4655,N_4591);
nand UO_801 (O_801,N_4870,N_4818);
and UO_802 (O_802,N_4844,N_4875);
nor UO_803 (O_803,N_4798,N_4734);
nor UO_804 (O_804,N_4528,N_4788);
nor UO_805 (O_805,N_4911,N_4621);
nor UO_806 (O_806,N_4521,N_4553);
or UO_807 (O_807,N_4663,N_4920);
nand UO_808 (O_808,N_4907,N_4612);
nor UO_809 (O_809,N_4537,N_4634);
and UO_810 (O_810,N_4578,N_4977);
nand UO_811 (O_811,N_4754,N_4957);
nand UO_812 (O_812,N_4912,N_4548);
nor UO_813 (O_813,N_4987,N_4771);
nand UO_814 (O_814,N_4511,N_4836);
or UO_815 (O_815,N_4843,N_4830);
nand UO_816 (O_816,N_4799,N_4720);
or UO_817 (O_817,N_4815,N_4742);
and UO_818 (O_818,N_4969,N_4607);
or UO_819 (O_819,N_4954,N_4568);
or UO_820 (O_820,N_4920,N_4824);
and UO_821 (O_821,N_4528,N_4725);
and UO_822 (O_822,N_4682,N_4691);
nand UO_823 (O_823,N_4654,N_4800);
and UO_824 (O_824,N_4723,N_4527);
or UO_825 (O_825,N_4567,N_4806);
or UO_826 (O_826,N_4553,N_4927);
or UO_827 (O_827,N_4990,N_4898);
or UO_828 (O_828,N_4886,N_4706);
or UO_829 (O_829,N_4751,N_4569);
nor UO_830 (O_830,N_4901,N_4761);
nand UO_831 (O_831,N_4930,N_4901);
and UO_832 (O_832,N_4847,N_4987);
and UO_833 (O_833,N_4686,N_4876);
nand UO_834 (O_834,N_4767,N_4817);
and UO_835 (O_835,N_4831,N_4943);
nand UO_836 (O_836,N_4766,N_4928);
nor UO_837 (O_837,N_4592,N_4902);
or UO_838 (O_838,N_4797,N_4794);
and UO_839 (O_839,N_4616,N_4958);
nand UO_840 (O_840,N_4720,N_4528);
nor UO_841 (O_841,N_4689,N_4883);
nand UO_842 (O_842,N_4879,N_4754);
xor UO_843 (O_843,N_4596,N_4936);
or UO_844 (O_844,N_4987,N_4830);
or UO_845 (O_845,N_4936,N_4850);
nor UO_846 (O_846,N_4749,N_4701);
and UO_847 (O_847,N_4774,N_4871);
and UO_848 (O_848,N_4776,N_4822);
and UO_849 (O_849,N_4756,N_4669);
nand UO_850 (O_850,N_4831,N_4669);
nor UO_851 (O_851,N_4720,N_4750);
or UO_852 (O_852,N_4516,N_4659);
or UO_853 (O_853,N_4819,N_4750);
or UO_854 (O_854,N_4972,N_4654);
nand UO_855 (O_855,N_4563,N_4722);
and UO_856 (O_856,N_4888,N_4519);
and UO_857 (O_857,N_4754,N_4772);
or UO_858 (O_858,N_4822,N_4709);
or UO_859 (O_859,N_4978,N_4637);
nor UO_860 (O_860,N_4741,N_4524);
and UO_861 (O_861,N_4643,N_4800);
nand UO_862 (O_862,N_4756,N_4547);
or UO_863 (O_863,N_4967,N_4996);
and UO_864 (O_864,N_4635,N_4744);
and UO_865 (O_865,N_4747,N_4698);
or UO_866 (O_866,N_4880,N_4696);
or UO_867 (O_867,N_4958,N_4771);
and UO_868 (O_868,N_4974,N_4555);
or UO_869 (O_869,N_4535,N_4540);
nand UO_870 (O_870,N_4785,N_4920);
nand UO_871 (O_871,N_4813,N_4555);
or UO_872 (O_872,N_4682,N_4749);
nand UO_873 (O_873,N_4967,N_4916);
nor UO_874 (O_874,N_4521,N_4827);
or UO_875 (O_875,N_4666,N_4972);
and UO_876 (O_876,N_4894,N_4688);
nand UO_877 (O_877,N_4857,N_4771);
and UO_878 (O_878,N_4771,N_4757);
nand UO_879 (O_879,N_4817,N_4966);
nand UO_880 (O_880,N_4872,N_4569);
and UO_881 (O_881,N_4673,N_4901);
nor UO_882 (O_882,N_4796,N_4911);
or UO_883 (O_883,N_4572,N_4618);
or UO_884 (O_884,N_4716,N_4678);
nand UO_885 (O_885,N_4994,N_4926);
nand UO_886 (O_886,N_4977,N_4736);
nor UO_887 (O_887,N_4749,N_4652);
and UO_888 (O_888,N_4730,N_4853);
or UO_889 (O_889,N_4624,N_4717);
nand UO_890 (O_890,N_4779,N_4745);
nor UO_891 (O_891,N_4511,N_4556);
and UO_892 (O_892,N_4952,N_4980);
and UO_893 (O_893,N_4893,N_4578);
nor UO_894 (O_894,N_4554,N_4875);
or UO_895 (O_895,N_4756,N_4933);
and UO_896 (O_896,N_4563,N_4578);
nor UO_897 (O_897,N_4618,N_4871);
nor UO_898 (O_898,N_4799,N_4758);
and UO_899 (O_899,N_4507,N_4990);
xor UO_900 (O_900,N_4852,N_4928);
and UO_901 (O_901,N_4923,N_4861);
and UO_902 (O_902,N_4654,N_4727);
nor UO_903 (O_903,N_4889,N_4547);
or UO_904 (O_904,N_4576,N_4603);
nor UO_905 (O_905,N_4513,N_4738);
or UO_906 (O_906,N_4876,N_4601);
and UO_907 (O_907,N_4952,N_4965);
nand UO_908 (O_908,N_4806,N_4804);
nor UO_909 (O_909,N_4519,N_4787);
or UO_910 (O_910,N_4638,N_4810);
nand UO_911 (O_911,N_4779,N_4648);
nand UO_912 (O_912,N_4810,N_4689);
or UO_913 (O_913,N_4905,N_4921);
nand UO_914 (O_914,N_4793,N_4799);
and UO_915 (O_915,N_4621,N_4878);
or UO_916 (O_916,N_4582,N_4799);
or UO_917 (O_917,N_4576,N_4546);
nor UO_918 (O_918,N_4867,N_4767);
nor UO_919 (O_919,N_4517,N_4675);
and UO_920 (O_920,N_4809,N_4893);
nor UO_921 (O_921,N_4895,N_4993);
nor UO_922 (O_922,N_4744,N_4625);
or UO_923 (O_923,N_4950,N_4827);
and UO_924 (O_924,N_4724,N_4647);
nor UO_925 (O_925,N_4711,N_4531);
or UO_926 (O_926,N_4587,N_4564);
xor UO_927 (O_927,N_4831,N_4861);
nand UO_928 (O_928,N_4955,N_4825);
or UO_929 (O_929,N_4864,N_4505);
and UO_930 (O_930,N_4839,N_4939);
xnor UO_931 (O_931,N_4900,N_4801);
nor UO_932 (O_932,N_4744,N_4580);
nand UO_933 (O_933,N_4690,N_4648);
or UO_934 (O_934,N_4642,N_4818);
nand UO_935 (O_935,N_4928,N_4584);
nor UO_936 (O_936,N_4689,N_4796);
nand UO_937 (O_937,N_4926,N_4657);
nand UO_938 (O_938,N_4948,N_4701);
nand UO_939 (O_939,N_4830,N_4895);
nor UO_940 (O_940,N_4872,N_4940);
nor UO_941 (O_941,N_4729,N_4749);
nand UO_942 (O_942,N_4629,N_4804);
nor UO_943 (O_943,N_4960,N_4731);
nor UO_944 (O_944,N_4783,N_4652);
nand UO_945 (O_945,N_4891,N_4764);
nor UO_946 (O_946,N_4954,N_4982);
and UO_947 (O_947,N_4895,N_4967);
and UO_948 (O_948,N_4595,N_4962);
nand UO_949 (O_949,N_4688,N_4532);
or UO_950 (O_950,N_4893,N_4754);
or UO_951 (O_951,N_4518,N_4598);
or UO_952 (O_952,N_4664,N_4965);
and UO_953 (O_953,N_4746,N_4662);
nand UO_954 (O_954,N_4721,N_4734);
nor UO_955 (O_955,N_4717,N_4742);
or UO_956 (O_956,N_4772,N_4589);
nand UO_957 (O_957,N_4902,N_4984);
and UO_958 (O_958,N_4603,N_4714);
nand UO_959 (O_959,N_4703,N_4525);
nand UO_960 (O_960,N_4615,N_4987);
nand UO_961 (O_961,N_4646,N_4905);
nand UO_962 (O_962,N_4608,N_4766);
nand UO_963 (O_963,N_4523,N_4891);
nor UO_964 (O_964,N_4750,N_4511);
and UO_965 (O_965,N_4504,N_4627);
and UO_966 (O_966,N_4661,N_4867);
nor UO_967 (O_967,N_4970,N_4544);
nand UO_968 (O_968,N_4729,N_4578);
or UO_969 (O_969,N_4631,N_4694);
nand UO_970 (O_970,N_4874,N_4566);
or UO_971 (O_971,N_4973,N_4866);
or UO_972 (O_972,N_4627,N_4611);
or UO_973 (O_973,N_4849,N_4769);
or UO_974 (O_974,N_4576,N_4989);
nand UO_975 (O_975,N_4891,N_4963);
or UO_976 (O_976,N_4779,N_4902);
nor UO_977 (O_977,N_4684,N_4681);
and UO_978 (O_978,N_4650,N_4813);
or UO_979 (O_979,N_4956,N_4704);
and UO_980 (O_980,N_4710,N_4589);
or UO_981 (O_981,N_4500,N_4572);
nand UO_982 (O_982,N_4821,N_4729);
or UO_983 (O_983,N_4552,N_4910);
nor UO_984 (O_984,N_4816,N_4669);
or UO_985 (O_985,N_4646,N_4588);
and UO_986 (O_986,N_4852,N_4776);
or UO_987 (O_987,N_4682,N_4602);
or UO_988 (O_988,N_4986,N_4524);
nand UO_989 (O_989,N_4580,N_4933);
or UO_990 (O_990,N_4616,N_4768);
nor UO_991 (O_991,N_4891,N_4873);
nand UO_992 (O_992,N_4911,N_4548);
nand UO_993 (O_993,N_4571,N_4981);
nand UO_994 (O_994,N_4664,N_4534);
xor UO_995 (O_995,N_4790,N_4735);
and UO_996 (O_996,N_4541,N_4999);
or UO_997 (O_997,N_4628,N_4677);
and UO_998 (O_998,N_4960,N_4802);
and UO_999 (O_999,N_4706,N_4876);
endmodule