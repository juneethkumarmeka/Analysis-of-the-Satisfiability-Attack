module basic_500_3000_500_40_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_397,In_76);
and U1 (N_1,In_325,In_479);
and U2 (N_2,In_320,In_136);
xnor U3 (N_3,In_321,In_208);
nand U4 (N_4,In_354,In_453);
nand U5 (N_5,In_34,In_295);
or U6 (N_6,In_350,In_499);
and U7 (N_7,In_251,In_171);
nand U8 (N_8,In_231,In_175);
nand U9 (N_9,In_126,In_240);
or U10 (N_10,In_299,In_108);
nor U11 (N_11,In_380,In_401);
nand U12 (N_12,In_406,In_264);
or U13 (N_13,In_75,In_496);
nor U14 (N_14,In_24,In_194);
and U15 (N_15,In_390,In_145);
nand U16 (N_16,In_253,In_13);
or U17 (N_17,In_296,In_464);
and U18 (N_18,In_210,In_166);
or U19 (N_19,In_116,In_167);
nand U20 (N_20,In_416,In_124);
nor U21 (N_21,In_329,In_310);
nand U22 (N_22,In_195,In_105);
nor U23 (N_23,In_54,In_213);
and U24 (N_24,In_92,In_254);
nand U25 (N_25,In_154,In_32);
nor U26 (N_26,In_478,In_368);
and U27 (N_27,In_130,In_435);
or U28 (N_28,In_66,In_217);
and U29 (N_29,In_104,In_50);
nand U30 (N_30,In_440,In_422);
or U31 (N_31,In_71,In_421);
nand U32 (N_32,In_138,In_59);
or U33 (N_33,In_163,In_311);
nor U34 (N_34,In_394,In_318);
nor U35 (N_35,In_375,In_257);
nor U36 (N_36,In_1,In_405);
or U37 (N_37,In_245,In_111);
nand U38 (N_38,In_176,In_216);
and U39 (N_39,In_330,In_449);
nand U40 (N_40,In_81,In_411);
nor U41 (N_41,In_234,In_441);
or U42 (N_42,In_414,In_140);
nand U43 (N_43,In_20,In_224);
nand U44 (N_44,In_308,In_336);
or U45 (N_45,In_309,In_369);
and U46 (N_46,In_121,In_474);
nor U47 (N_47,In_12,In_353);
and U48 (N_48,In_387,In_399);
nor U49 (N_49,In_278,In_112);
and U50 (N_50,In_101,In_8);
or U51 (N_51,In_347,In_383);
nor U52 (N_52,In_284,In_62);
nand U53 (N_53,In_495,In_333);
nand U54 (N_54,In_365,In_72);
or U55 (N_55,In_139,In_317);
nand U56 (N_56,In_212,In_226);
nor U57 (N_57,In_470,In_31);
nand U58 (N_58,In_243,In_425);
and U59 (N_59,In_300,In_388);
nand U60 (N_60,In_182,In_91);
or U61 (N_61,In_18,In_36);
or U62 (N_62,In_40,In_131);
and U63 (N_63,In_389,In_413);
nor U64 (N_64,In_274,In_491);
or U65 (N_65,In_181,In_94);
or U66 (N_66,In_52,In_261);
or U67 (N_67,In_385,In_438);
and U68 (N_68,In_476,In_444);
nor U69 (N_69,In_459,In_125);
nor U70 (N_70,In_146,In_291);
nor U71 (N_71,In_233,In_467);
and U72 (N_72,In_437,In_96);
and U73 (N_73,In_424,In_119);
or U74 (N_74,In_11,In_396);
and U75 (N_75,In_327,In_346);
nand U76 (N_76,In_358,In_481);
and U77 (N_77,N_7,In_69);
and U78 (N_78,In_99,In_16);
and U79 (N_79,In_279,In_48);
nand U80 (N_80,N_14,In_391);
and U81 (N_81,In_366,N_52);
nor U82 (N_82,N_70,In_219);
and U83 (N_83,In_443,In_103);
nor U84 (N_84,In_78,In_258);
nor U85 (N_85,In_335,In_79);
and U86 (N_86,In_22,In_83);
nor U87 (N_87,In_6,N_72);
nand U88 (N_88,In_307,In_410);
nor U89 (N_89,N_49,In_386);
nor U90 (N_90,In_46,N_12);
or U91 (N_91,In_169,In_41);
or U92 (N_92,In_316,In_74);
nand U93 (N_93,In_0,In_191);
and U94 (N_94,N_42,In_141);
and U95 (N_95,In_428,In_271);
and U96 (N_96,In_82,In_493);
and U97 (N_97,In_51,In_227);
or U98 (N_98,N_18,In_142);
nor U99 (N_99,In_482,In_2);
nand U100 (N_100,In_432,N_38);
and U101 (N_101,In_475,N_10);
nand U102 (N_102,In_306,In_262);
nor U103 (N_103,N_13,In_305);
nand U104 (N_104,N_60,In_361);
nand U105 (N_105,In_393,In_324);
nor U106 (N_106,In_42,In_415);
xnor U107 (N_107,In_448,In_352);
nor U108 (N_108,In_342,In_122);
and U109 (N_109,In_199,In_331);
nor U110 (N_110,N_20,In_268);
or U111 (N_111,In_447,In_137);
and U112 (N_112,In_345,N_58);
nor U113 (N_113,In_88,In_473);
nand U114 (N_114,In_466,In_497);
or U115 (N_115,N_51,In_289);
nor U116 (N_116,N_45,In_298);
nor U117 (N_117,In_149,N_16);
nor U118 (N_118,In_269,N_61);
nor U119 (N_119,In_86,In_285);
nand U120 (N_120,In_382,In_275);
and U121 (N_121,In_110,In_26);
or U122 (N_122,In_256,In_259);
nand U123 (N_123,In_168,In_209);
nor U124 (N_124,In_292,In_118);
or U125 (N_125,In_188,In_38);
nor U126 (N_126,N_25,In_148);
or U127 (N_127,In_374,In_419);
or U128 (N_128,In_402,In_370);
nand U129 (N_129,In_266,In_23);
and U130 (N_130,N_59,In_270);
and U131 (N_131,In_90,In_263);
nor U132 (N_132,N_19,In_356);
nor U133 (N_133,In_98,In_303);
xor U134 (N_134,In_60,In_328);
or U135 (N_135,In_472,In_37);
and U136 (N_136,N_71,In_102);
nand U137 (N_137,In_384,In_334);
nor U138 (N_138,In_326,In_283);
nand U139 (N_139,In_355,In_183);
nor U140 (N_140,In_107,In_128);
nor U141 (N_141,In_164,In_152);
nand U142 (N_142,In_35,In_85);
nand U143 (N_143,In_323,In_201);
nor U144 (N_144,In_132,In_290);
or U145 (N_145,In_160,In_127);
and U146 (N_146,In_73,In_357);
and U147 (N_147,In_403,In_109);
nand U148 (N_148,In_123,N_47);
and U149 (N_149,In_417,In_319);
nor U150 (N_150,In_172,In_407);
nor U151 (N_151,In_408,In_490);
nand U152 (N_152,N_105,In_49);
nand U153 (N_153,In_452,In_282);
and U154 (N_154,In_252,In_445);
and U155 (N_155,In_484,In_114);
nor U156 (N_156,N_145,N_112);
and U157 (N_157,In_376,N_115);
nand U158 (N_158,N_31,In_203);
nor U159 (N_159,N_56,In_486);
and U160 (N_160,N_15,In_398);
nand U161 (N_161,N_89,In_260);
nor U162 (N_162,In_161,In_492);
and U163 (N_163,N_131,In_426);
or U164 (N_164,In_10,In_280);
nand U165 (N_165,In_3,N_139);
and U166 (N_166,In_97,N_147);
or U167 (N_167,N_130,N_98);
nand U168 (N_168,N_63,N_96);
and U169 (N_169,N_35,In_221);
or U170 (N_170,In_429,In_273);
or U171 (N_171,N_62,N_81);
nor U172 (N_172,N_140,In_427);
or U173 (N_173,N_108,In_28);
or U174 (N_174,N_94,In_206);
or U175 (N_175,In_436,In_235);
nor U176 (N_176,N_82,In_272);
nand U177 (N_177,In_19,N_128);
or U178 (N_178,N_68,N_86);
or U179 (N_179,In_190,In_238);
nor U180 (N_180,In_373,N_32);
and U181 (N_181,N_67,In_187);
nand U182 (N_182,N_53,In_14);
nand U183 (N_183,In_115,In_93);
nor U184 (N_184,In_27,In_215);
nand U185 (N_185,In_379,N_84);
nand U186 (N_186,N_55,In_214);
nand U187 (N_187,In_430,N_74);
and U188 (N_188,In_313,N_33);
nand U189 (N_189,In_129,N_143);
nor U190 (N_190,N_36,In_43);
nor U191 (N_191,In_293,N_21);
and U192 (N_192,In_457,N_30);
nor U193 (N_193,In_232,In_371);
nand U194 (N_194,In_439,N_124);
nand U195 (N_195,N_107,N_148);
nand U196 (N_196,In_400,N_46);
nor U197 (N_197,In_134,In_343);
and U198 (N_198,N_134,In_67);
nor U199 (N_199,In_244,In_494);
or U200 (N_200,N_132,In_223);
nor U201 (N_201,In_367,In_162);
nor U202 (N_202,N_44,N_100);
nor U203 (N_203,In_225,In_468);
or U204 (N_204,N_113,In_360);
or U205 (N_205,N_138,N_95);
nor U206 (N_206,In_281,In_480);
nand U207 (N_207,N_29,In_30);
and U208 (N_208,In_159,In_246);
nor U209 (N_209,In_70,N_64);
and U210 (N_210,N_1,In_241);
nand U211 (N_211,N_57,In_184);
and U212 (N_212,In_409,In_193);
nand U213 (N_213,In_5,In_56);
nor U214 (N_214,In_442,In_192);
and U215 (N_215,N_104,In_53);
nor U216 (N_216,In_412,In_465);
or U217 (N_217,N_73,In_84);
and U218 (N_218,In_135,In_276);
nor U219 (N_219,In_211,N_39);
and U220 (N_220,In_456,N_0);
nand U221 (N_221,In_21,N_149);
and U222 (N_222,N_23,N_117);
and U223 (N_223,N_103,In_454);
nor U224 (N_224,In_338,In_301);
and U225 (N_225,In_242,N_34);
nand U226 (N_226,In_100,In_477);
or U227 (N_227,N_2,N_204);
nand U228 (N_228,N_209,N_121);
or U229 (N_229,N_198,N_159);
or U230 (N_230,In_351,In_58);
or U231 (N_231,N_90,In_200);
nor U232 (N_232,N_187,In_61);
or U233 (N_233,N_189,N_125);
and U234 (N_234,N_210,N_220);
and U235 (N_235,In_471,N_218);
and U236 (N_236,In_341,N_156);
and U237 (N_237,N_83,In_302);
nor U238 (N_238,N_177,In_158);
nand U239 (N_239,In_63,In_315);
nand U240 (N_240,N_120,In_377);
nor U241 (N_241,N_188,In_230);
nor U242 (N_242,In_277,N_6);
nor U243 (N_243,In_297,N_141);
nand U244 (N_244,In_25,In_489);
nand U245 (N_245,In_248,In_147);
or U246 (N_246,In_458,N_65);
and U247 (N_247,N_151,N_101);
and U248 (N_248,In_249,In_68);
nand U249 (N_249,N_150,In_485);
and U250 (N_250,In_332,In_95);
and U251 (N_251,N_182,In_434);
or U252 (N_252,In_173,N_91);
or U253 (N_253,N_163,N_178);
nor U254 (N_254,In_265,N_122);
and U255 (N_255,N_40,N_191);
and U256 (N_256,In_362,N_102);
or U257 (N_257,In_314,In_207);
nand U258 (N_258,N_223,N_222);
nand U259 (N_259,In_337,In_120);
nor U260 (N_260,N_4,In_55);
or U261 (N_261,In_446,N_106);
and U262 (N_262,N_79,N_11);
nor U263 (N_263,N_219,In_197);
and U264 (N_264,In_488,In_220);
nor U265 (N_265,In_487,N_26);
nand U266 (N_266,In_404,N_99);
nand U267 (N_267,N_54,N_166);
nor U268 (N_268,N_116,N_27);
nor U269 (N_269,N_206,In_287);
or U270 (N_270,N_216,In_144);
or U271 (N_271,In_179,N_123);
and U272 (N_272,N_66,In_15);
nor U273 (N_273,In_57,N_144);
nand U274 (N_274,In_177,In_395);
or U275 (N_275,In_433,In_178);
nand U276 (N_276,In_469,N_137);
nor U277 (N_277,N_162,N_168);
nand U278 (N_278,In_364,N_109);
or U279 (N_279,N_85,N_186);
nor U280 (N_280,In_204,In_418);
or U281 (N_281,N_152,In_113);
or U282 (N_282,N_142,N_78);
or U283 (N_283,N_224,N_114);
xor U284 (N_284,In_196,In_77);
or U285 (N_285,N_192,N_92);
and U286 (N_286,In_322,N_194);
nand U287 (N_287,In_267,In_420);
nor U288 (N_288,N_184,N_211);
nand U289 (N_289,N_172,N_154);
nor U290 (N_290,In_255,In_205);
nand U291 (N_291,N_213,In_312);
xnor U292 (N_292,In_156,In_228);
or U293 (N_293,N_202,N_76);
and U294 (N_294,N_190,In_185);
nand U295 (N_295,N_24,In_151);
or U296 (N_296,N_50,In_89);
nor U297 (N_297,N_3,N_153);
nand U298 (N_298,In_247,N_69);
xnor U299 (N_299,N_176,In_9);
nand U300 (N_300,In_339,N_256);
or U301 (N_301,N_127,In_239);
nor U302 (N_302,N_299,In_348);
and U303 (N_303,N_234,N_273);
nor U304 (N_304,N_93,N_249);
nor U305 (N_305,N_264,In_180);
and U306 (N_306,N_227,N_236);
nand U307 (N_307,N_285,In_143);
nand U308 (N_308,In_237,N_181);
or U309 (N_309,N_208,N_41);
nand U310 (N_310,N_239,N_158);
nor U311 (N_311,N_229,N_267);
nor U312 (N_312,In_150,In_381);
or U313 (N_313,In_106,In_202);
or U314 (N_314,In_236,N_258);
or U315 (N_315,N_246,In_64);
and U316 (N_316,In_483,N_231);
and U317 (N_317,In_47,N_262);
or U318 (N_318,N_157,In_392);
nor U319 (N_319,N_161,In_153);
or U320 (N_320,N_291,N_111);
nor U321 (N_321,N_110,N_173);
nand U322 (N_322,N_196,In_45);
and U323 (N_323,N_297,N_263);
nand U324 (N_324,In_157,In_431);
or U325 (N_325,In_498,N_243);
nand U326 (N_326,N_199,In_460);
nor U327 (N_327,N_217,In_250);
nand U328 (N_328,In_155,N_88);
nand U329 (N_329,N_203,N_221);
and U330 (N_330,N_225,N_293);
nand U331 (N_331,N_287,N_269);
or U332 (N_332,N_201,N_292);
nand U333 (N_333,N_87,N_242);
nor U334 (N_334,N_169,N_17);
nand U335 (N_335,In_65,N_241);
and U336 (N_336,N_226,N_215);
and U337 (N_337,N_245,N_228);
or U338 (N_338,N_167,In_165);
nor U339 (N_339,In_29,In_218);
nor U340 (N_340,In_39,N_237);
nor U341 (N_341,N_278,In_450);
and U342 (N_342,N_179,In_133);
nand U343 (N_343,In_359,N_260);
or U344 (N_344,N_97,N_193);
nor U345 (N_345,In_174,In_461);
or U346 (N_346,In_288,In_4);
nor U347 (N_347,N_270,In_117);
and U348 (N_348,N_37,N_268);
nand U349 (N_349,In_462,In_363);
and U350 (N_350,N_160,N_247);
nor U351 (N_351,N_272,N_135);
nand U352 (N_352,In_80,N_259);
nor U353 (N_353,In_222,N_180);
nand U354 (N_354,N_22,N_288);
or U355 (N_355,In_455,N_235);
nor U356 (N_356,N_295,N_279);
nand U357 (N_357,N_257,N_250);
or U358 (N_358,N_8,N_277);
or U359 (N_359,N_136,In_423);
or U360 (N_360,N_286,N_230);
or U361 (N_361,N_174,In_286);
or U362 (N_362,N_200,N_289);
and U363 (N_363,In_17,N_253);
nand U364 (N_364,In_198,In_451);
nand U365 (N_365,N_296,N_244);
and U366 (N_366,N_43,In_294);
and U367 (N_367,In_344,N_276);
and U368 (N_368,N_254,N_77);
or U369 (N_369,N_129,N_240);
nand U370 (N_370,N_183,N_5);
or U371 (N_371,N_251,In_340);
nand U372 (N_372,N_282,In_304);
nand U373 (N_373,N_146,N_274);
nor U374 (N_374,N_164,N_284);
xor U375 (N_375,N_248,N_294);
or U376 (N_376,N_255,N_283);
and U377 (N_377,N_342,N_333);
nand U378 (N_378,N_28,N_339);
nand U379 (N_379,N_175,N_366);
or U380 (N_380,N_352,N_361);
nand U381 (N_381,N_185,N_214);
or U382 (N_382,N_324,N_308);
and U383 (N_383,N_330,In_463);
and U384 (N_384,N_155,N_354);
and U385 (N_385,N_48,N_351);
nor U386 (N_386,N_368,N_290);
nand U387 (N_387,In_186,N_356);
or U388 (N_388,N_340,N_300);
or U389 (N_389,N_80,N_75);
and U390 (N_390,N_343,N_301);
and U391 (N_391,N_332,N_9);
and U392 (N_392,N_374,N_370);
nor U393 (N_393,N_266,N_281);
or U394 (N_394,N_170,N_310);
nand U395 (N_395,N_315,N_212);
or U396 (N_396,N_205,N_358);
nor U397 (N_397,N_252,N_197);
or U398 (N_398,N_207,N_319);
nand U399 (N_399,N_322,N_371);
nor U400 (N_400,N_298,In_33);
nand U401 (N_401,N_119,N_344);
or U402 (N_402,N_338,N_133);
xnor U403 (N_403,N_265,N_320);
or U404 (N_404,N_304,N_126);
nand U405 (N_405,In_170,N_334);
or U406 (N_406,In_189,N_327);
and U407 (N_407,In_87,N_331);
and U408 (N_408,N_346,N_305);
or U409 (N_409,N_321,N_365);
or U410 (N_410,N_311,N_364);
or U411 (N_411,N_316,N_233);
or U412 (N_412,In_44,N_373);
nor U413 (N_413,N_313,N_337);
nor U414 (N_414,N_306,N_335);
nor U415 (N_415,N_349,In_349);
nor U416 (N_416,N_232,N_307);
nor U417 (N_417,N_329,N_359);
and U418 (N_418,In_7,N_309);
or U419 (N_419,N_302,N_353);
and U420 (N_420,In_229,N_303);
and U421 (N_421,N_261,N_171);
or U422 (N_422,N_238,N_360);
nand U423 (N_423,N_323,N_345);
and U424 (N_424,N_326,N_312);
and U425 (N_425,N_362,N_271);
and U426 (N_426,N_341,N_328);
or U427 (N_427,N_275,N_350);
nor U428 (N_428,N_347,N_336);
or U429 (N_429,N_369,N_355);
xnor U430 (N_430,N_318,N_118);
and U431 (N_431,N_280,N_363);
or U432 (N_432,N_367,N_195);
nor U433 (N_433,N_357,In_372);
nand U434 (N_434,N_372,N_165);
nor U435 (N_435,In_378,N_325);
and U436 (N_436,N_317,N_314);
or U437 (N_437,N_348,N_118);
or U438 (N_438,N_311,N_355);
nor U439 (N_439,N_357,N_354);
nand U440 (N_440,N_319,N_175);
or U441 (N_441,N_175,N_365);
nand U442 (N_442,N_356,N_306);
nand U443 (N_443,N_336,N_238);
nand U444 (N_444,N_306,N_165);
nand U445 (N_445,In_44,N_214);
nand U446 (N_446,N_207,N_373);
nand U447 (N_447,In_189,N_369);
or U448 (N_448,N_337,N_265);
and U449 (N_449,N_316,N_126);
and U450 (N_450,N_433,N_419);
or U451 (N_451,N_394,N_408);
and U452 (N_452,N_415,N_427);
or U453 (N_453,N_379,N_384);
or U454 (N_454,N_436,N_414);
nor U455 (N_455,N_446,N_431);
or U456 (N_456,N_440,N_412);
nand U457 (N_457,N_399,N_441);
and U458 (N_458,N_396,N_432);
nor U459 (N_459,N_434,N_392);
and U460 (N_460,N_404,N_411);
nor U461 (N_461,N_390,N_443);
and U462 (N_462,N_410,N_435);
or U463 (N_463,N_389,N_377);
or U464 (N_464,N_449,N_423);
or U465 (N_465,N_420,N_421);
nor U466 (N_466,N_428,N_378);
or U467 (N_467,N_388,N_391);
and U468 (N_468,N_442,N_385);
and U469 (N_469,N_383,N_413);
and U470 (N_470,N_418,N_417);
nand U471 (N_471,N_381,N_448);
nor U472 (N_472,N_375,N_393);
nor U473 (N_473,N_445,N_407);
nand U474 (N_474,N_439,N_426);
or U475 (N_475,N_409,N_416);
or U476 (N_476,N_376,N_425);
nand U477 (N_477,N_437,N_398);
or U478 (N_478,N_430,N_395);
and U479 (N_479,N_444,N_438);
nand U480 (N_480,N_429,N_401);
nand U481 (N_481,N_382,N_405);
nor U482 (N_482,N_387,N_406);
and U483 (N_483,N_403,N_397);
nand U484 (N_484,N_424,N_422);
and U485 (N_485,N_386,N_400);
and U486 (N_486,N_402,N_447);
and U487 (N_487,N_380,N_424);
nor U488 (N_488,N_404,N_377);
or U489 (N_489,N_422,N_375);
nand U490 (N_490,N_376,N_446);
or U491 (N_491,N_429,N_403);
and U492 (N_492,N_436,N_444);
nand U493 (N_493,N_438,N_377);
nor U494 (N_494,N_389,N_411);
nor U495 (N_495,N_448,N_443);
or U496 (N_496,N_427,N_380);
nor U497 (N_497,N_382,N_442);
or U498 (N_498,N_385,N_408);
nand U499 (N_499,N_405,N_398);
nand U500 (N_500,N_424,N_445);
nor U501 (N_501,N_423,N_406);
and U502 (N_502,N_381,N_398);
or U503 (N_503,N_408,N_391);
nor U504 (N_504,N_394,N_402);
or U505 (N_505,N_395,N_402);
or U506 (N_506,N_430,N_415);
or U507 (N_507,N_400,N_380);
and U508 (N_508,N_439,N_430);
nand U509 (N_509,N_405,N_416);
or U510 (N_510,N_406,N_392);
and U511 (N_511,N_436,N_391);
nand U512 (N_512,N_397,N_398);
nor U513 (N_513,N_427,N_405);
or U514 (N_514,N_382,N_396);
or U515 (N_515,N_380,N_395);
and U516 (N_516,N_418,N_402);
and U517 (N_517,N_403,N_393);
nand U518 (N_518,N_444,N_449);
nor U519 (N_519,N_421,N_383);
nor U520 (N_520,N_435,N_424);
nand U521 (N_521,N_417,N_379);
or U522 (N_522,N_448,N_445);
nor U523 (N_523,N_430,N_434);
nor U524 (N_524,N_380,N_408);
and U525 (N_525,N_471,N_463);
or U526 (N_526,N_521,N_493);
or U527 (N_527,N_469,N_484);
and U528 (N_528,N_478,N_455);
and U529 (N_529,N_503,N_494);
and U530 (N_530,N_473,N_474);
or U531 (N_531,N_513,N_460);
nor U532 (N_532,N_495,N_482);
nor U533 (N_533,N_492,N_480);
nor U534 (N_534,N_458,N_477);
nor U535 (N_535,N_500,N_459);
nand U536 (N_536,N_456,N_487);
or U537 (N_537,N_466,N_517);
and U538 (N_538,N_481,N_467);
xor U539 (N_539,N_461,N_453);
and U540 (N_540,N_470,N_483);
nand U541 (N_541,N_504,N_515);
nand U542 (N_542,N_486,N_451);
and U543 (N_543,N_488,N_507);
nor U544 (N_544,N_514,N_464);
nor U545 (N_545,N_450,N_505);
nand U546 (N_546,N_485,N_491);
or U547 (N_547,N_479,N_496);
nor U548 (N_548,N_501,N_476);
and U549 (N_549,N_508,N_497);
or U550 (N_550,N_524,N_452);
nand U551 (N_551,N_489,N_502);
nand U552 (N_552,N_457,N_462);
nor U553 (N_553,N_518,N_523);
nand U554 (N_554,N_498,N_516);
and U555 (N_555,N_490,N_499);
nor U556 (N_556,N_510,N_519);
and U557 (N_557,N_468,N_475);
nor U558 (N_558,N_454,N_512);
or U559 (N_559,N_522,N_465);
nand U560 (N_560,N_520,N_506);
and U561 (N_561,N_511,N_472);
or U562 (N_562,N_509,N_459);
nor U563 (N_563,N_486,N_524);
or U564 (N_564,N_515,N_456);
nor U565 (N_565,N_464,N_490);
nor U566 (N_566,N_462,N_478);
nor U567 (N_567,N_493,N_505);
and U568 (N_568,N_475,N_481);
and U569 (N_569,N_518,N_503);
nor U570 (N_570,N_521,N_483);
nand U571 (N_571,N_454,N_453);
nand U572 (N_572,N_493,N_520);
nor U573 (N_573,N_454,N_460);
nor U574 (N_574,N_455,N_520);
or U575 (N_575,N_501,N_480);
or U576 (N_576,N_464,N_462);
nor U577 (N_577,N_513,N_508);
nor U578 (N_578,N_471,N_518);
nor U579 (N_579,N_487,N_515);
nor U580 (N_580,N_521,N_524);
or U581 (N_581,N_521,N_457);
or U582 (N_582,N_482,N_509);
and U583 (N_583,N_476,N_454);
or U584 (N_584,N_511,N_521);
nor U585 (N_585,N_486,N_487);
or U586 (N_586,N_524,N_450);
and U587 (N_587,N_522,N_477);
nand U588 (N_588,N_450,N_522);
nand U589 (N_589,N_520,N_497);
nor U590 (N_590,N_519,N_479);
nor U591 (N_591,N_461,N_493);
nand U592 (N_592,N_495,N_523);
nor U593 (N_593,N_517,N_472);
nand U594 (N_594,N_453,N_511);
nand U595 (N_595,N_486,N_484);
nor U596 (N_596,N_450,N_463);
nand U597 (N_597,N_507,N_496);
nor U598 (N_598,N_507,N_469);
nand U599 (N_599,N_498,N_453);
nand U600 (N_600,N_560,N_543);
and U601 (N_601,N_542,N_557);
nor U602 (N_602,N_528,N_565);
and U603 (N_603,N_561,N_529);
and U604 (N_604,N_527,N_536);
and U605 (N_605,N_526,N_531);
nor U606 (N_606,N_558,N_583);
nor U607 (N_607,N_530,N_555);
nand U608 (N_608,N_575,N_532);
and U609 (N_609,N_580,N_540);
nor U610 (N_610,N_576,N_598);
nand U611 (N_611,N_563,N_570);
and U612 (N_612,N_577,N_590);
and U613 (N_613,N_548,N_535);
or U614 (N_614,N_595,N_533);
or U615 (N_615,N_569,N_588);
and U616 (N_616,N_544,N_593);
nand U617 (N_617,N_549,N_559);
nand U618 (N_618,N_545,N_541);
nand U619 (N_619,N_538,N_594);
or U620 (N_620,N_596,N_556);
or U621 (N_621,N_525,N_567);
or U622 (N_622,N_572,N_550);
or U623 (N_623,N_551,N_578);
nor U624 (N_624,N_585,N_592);
or U625 (N_625,N_584,N_589);
or U626 (N_626,N_566,N_582);
nand U627 (N_627,N_547,N_568);
nand U628 (N_628,N_574,N_537);
or U629 (N_629,N_599,N_562);
or U630 (N_630,N_546,N_571);
nand U631 (N_631,N_597,N_554);
nor U632 (N_632,N_581,N_564);
or U633 (N_633,N_579,N_573);
or U634 (N_634,N_552,N_534);
and U635 (N_635,N_587,N_586);
nand U636 (N_636,N_591,N_553);
or U637 (N_637,N_539,N_575);
nor U638 (N_638,N_556,N_567);
or U639 (N_639,N_583,N_533);
or U640 (N_640,N_571,N_561);
nand U641 (N_641,N_594,N_541);
or U642 (N_642,N_575,N_584);
nand U643 (N_643,N_584,N_539);
nand U644 (N_644,N_535,N_558);
nor U645 (N_645,N_559,N_530);
nand U646 (N_646,N_539,N_548);
nand U647 (N_647,N_573,N_541);
and U648 (N_648,N_547,N_530);
and U649 (N_649,N_575,N_585);
and U650 (N_650,N_551,N_554);
nand U651 (N_651,N_596,N_586);
nand U652 (N_652,N_589,N_575);
or U653 (N_653,N_594,N_588);
and U654 (N_654,N_572,N_534);
and U655 (N_655,N_558,N_578);
and U656 (N_656,N_550,N_532);
and U657 (N_657,N_561,N_533);
nor U658 (N_658,N_533,N_554);
nor U659 (N_659,N_545,N_586);
and U660 (N_660,N_528,N_537);
nor U661 (N_661,N_583,N_560);
or U662 (N_662,N_552,N_590);
and U663 (N_663,N_569,N_594);
and U664 (N_664,N_590,N_589);
or U665 (N_665,N_585,N_567);
nor U666 (N_666,N_584,N_577);
nor U667 (N_667,N_546,N_552);
and U668 (N_668,N_559,N_578);
nand U669 (N_669,N_561,N_594);
or U670 (N_670,N_590,N_535);
nand U671 (N_671,N_577,N_544);
nor U672 (N_672,N_529,N_545);
and U673 (N_673,N_569,N_575);
nor U674 (N_674,N_580,N_556);
and U675 (N_675,N_615,N_610);
or U676 (N_676,N_632,N_664);
or U677 (N_677,N_625,N_642);
nand U678 (N_678,N_645,N_633);
and U679 (N_679,N_656,N_674);
or U680 (N_680,N_649,N_600);
nand U681 (N_681,N_662,N_672);
nor U682 (N_682,N_663,N_665);
nand U683 (N_683,N_660,N_648);
or U684 (N_684,N_602,N_670);
and U685 (N_685,N_655,N_669);
and U686 (N_686,N_641,N_629);
nand U687 (N_687,N_623,N_650);
and U688 (N_688,N_628,N_637);
nand U689 (N_689,N_661,N_604);
nand U690 (N_690,N_616,N_630);
nor U691 (N_691,N_653,N_638);
nand U692 (N_692,N_624,N_613);
or U693 (N_693,N_626,N_618);
or U694 (N_694,N_652,N_631);
or U695 (N_695,N_659,N_622);
nand U696 (N_696,N_608,N_601);
and U697 (N_697,N_657,N_639);
or U698 (N_698,N_607,N_612);
nor U699 (N_699,N_654,N_619);
nand U700 (N_700,N_667,N_636);
nor U701 (N_701,N_666,N_606);
nand U702 (N_702,N_646,N_658);
or U703 (N_703,N_634,N_640);
nand U704 (N_704,N_627,N_614);
or U705 (N_705,N_671,N_609);
nand U706 (N_706,N_621,N_668);
or U707 (N_707,N_635,N_644);
nor U708 (N_708,N_603,N_605);
or U709 (N_709,N_647,N_643);
nor U710 (N_710,N_620,N_617);
and U711 (N_711,N_673,N_611);
or U712 (N_712,N_651,N_619);
or U713 (N_713,N_650,N_603);
and U714 (N_714,N_669,N_630);
or U715 (N_715,N_674,N_615);
nand U716 (N_716,N_652,N_600);
nor U717 (N_717,N_610,N_600);
and U718 (N_718,N_616,N_621);
nor U719 (N_719,N_624,N_620);
nor U720 (N_720,N_658,N_643);
and U721 (N_721,N_613,N_665);
nand U722 (N_722,N_651,N_667);
nand U723 (N_723,N_643,N_673);
nor U724 (N_724,N_639,N_653);
nor U725 (N_725,N_620,N_630);
nand U726 (N_726,N_637,N_672);
or U727 (N_727,N_657,N_659);
and U728 (N_728,N_646,N_608);
and U729 (N_729,N_629,N_664);
and U730 (N_730,N_613,N_642);
or U731 (N_731,N_674,N_658);
or U732 (N_732,N_622,N_638);
and U733 (N_733,N_656,N_672);
nand U734 (N_734,N_656,N_673);
nor U735 (N_735,N_642,N_650);
and U736 (N_736,N_656,N_644);
and U737 (N_737,N_674,N_673);
nor U738 (N_738,N_649,N_647);
nor U739 (N_739,N_663,N_600);
nand U740 (N_740,N_632,N_668);
and U741 (N_741,N_639,N_669);
and U742 (N_742,N_609,N_618);
and U743 (N_743,N_656,N_606);
nand U744 (N_744,N_674,N_607);
nand U745 (N_745,N_619,N_648);
or U746 (N_746,N_603,N_611);
nor U747 (N_747,N_606,N_613);
or U748 (N_748,N_612,N_669);
nor U749 (N_749,N_605,N_661);
and U750 (N_750,N_748,N_684);
and U751 (N_751,N_726,N_716);
or U752 (N_752,N_723,N_729);
nand U753 (N_753,N_744,N_685);
or U754 (N_754,N_707,N_687);
and U755 (N_755,N_708,N_691);
nor U756 (N_756,N_703,N_705);
nor U757 (N_757,N_747,N_682);
nand U758 (N_758,N_735,N_722);
and U759 (N_759,N_737,N_749);
and U760 (N_760,N_734,N_740);
and U761 (N_761,N_746,N_741);
and U762 (N_762,N_679,N_690);
or U763 (N_763,N_720,N_695);
nand U764 (N_764,N_732,N_696);
nor U765 (N_765,N_715,N_704);
and U766 (N_766,N_698,N_713);
nor U767 (N_767,N_710,N_733);
and U768 (N_768,N_692,N_700);
nand U769 (N_769,N_681,N_743);
nor U770 (N_770,N_699,N_675);
nand U771 (N_771,N_727,N_714);
and U772 (N_772,N_736,N_725);
nand U773 (N_773,N_739,N_697);
nor U774 (N_774,N_738,N_745);
xnor U775 (N_775,N_688,N_728);
or U776 (N_776,N_680,N_712);
or U777 (N_777,N_742,N_702);
nor U778 (N_778,N_683,N_719);
and U779 (N_779,N_709,N_730);
or U780 (N_780,N_678,N_731);
nand U781 (N_781,N_706,N_694);
and U782 (N_782,N_711,N_676);
nand U783 (N_783,N_689,N_724);
and U784 (N_784,N_721,N_718);
and U785 (N_785,N_686,N_717);
or U786 (N_786,N_677,N_693);
nor U787 (N_787,N_701,N_677);
nor U788 (N_788,N_713,N_699);
nand U789 (N_789,N_735,N_740);
nor U790 (N_790,N_714,N_734);
and U791 (N_791,N_689,N_731);
nand U792 (N_792,N_679,N_721);
or U793 (N_793,N_690,N_744);
nor U794 (N_794,N_696,N_740);
nand U795 (N_795,N_729,N_745);
nand U796 (N_796,N_731,N_743);
nor U797 (N_797,N_685,N_742);
or U798 (N_798,N_713,N_680);
nand U799 (N_799,N_679,N_688);
and U800 (N_800,N_690,N_739);
or U801 (N_801,N_691,N_749);
nor U802 (N_802,N_694,N_738);
nand U803 (N_803,N_725,N_696);
nor U804 (N_804,N_728,N_709);
and U805 (N_805,N_690,N_697);
and U806 (N_806,N_730,N_735);
nor U807 (N_807,N_706,N_713);
nor U808 (N_808,N_692,N_714);
nand U809 (N_809,N_707,N_694);
nand U810 (N_810,N_690,N_695);
nand U811 (N_811,N_720,N_725);
and U812 (N_812,N_724,N_709);
and U813 (N_813,N_747,N_737);
or U814 (N_814,N_739,N_693);
or U815 (N_815,N_699,N_728);
nand U816 (N_816,N_742,N_696);
and U817 (N_817,N_745,N_694);
nor U818 (N_818,N_731,N_735);
nor U819 (N_819,N_691,N_719);
and U820 (N_820,N_732,N_715);
nor U821 (N_821,N_742,N_706);
nor U822 (N_822,N_712,N_744);
nor U823 (N_823,N_701,N_705);
or U824 (N_824,N_687,N_703);
and U825 (N_825,N_750,N_753);
and U826 (N_826,N_809,N_789);
or U827 (N_827,N_775,N_791);
nand U828 (N_828,N_767,N_822);
nor U829 (N_829,N_782,N_808);
nor U830 (N_830,N_821,N_798);
or U831 (N_831,N_824,N_762);
or U832 (N_832,N_751,N_803);
nand U833 (N_833,N_795,N_792);
nand U834 (N_834,N_759,N_760);
nor U835 (N_835,N_776,N_787);
nand U836 (N_836,N_756,N_768);
nand U837 (N_837,N_816,N_810);
or U838 (N_838,N_823,N_814);
nand U839 (N_839,N_770,N_769);
and U840 (N_840,N_806,N_793);
nor U841 (N_841,N_779,N_761);
nor U842 (N_842,N_784,N_799);
nand U843 (N_843,N_755,N_766);
nor U844 (N_844,N_774,N_752);
or U845 (N_845,N_807,N_772);
or U846 (N_846,N_758,N_771);
or U847 (N_847,N_763,N_818);
and U848 (N_848,N_817,N_813);
nor U849 (N_849,N_777,N_757);
or U850 (N_850,N_790,N_797);
nand U851 (N_851,N_794,N_819);
nor U852 (N_852,N_815,N_785);
or U853 (N_853,N_820,N_781);
nor U854 (N_854,N_754,N_796);
or U855 (N_855,N_801,N_812);
nor U856 (N_856,N_783,N_773);
or U857 (N_857,N_788,N_802);
and U858 (N_858,N_804,N_805);
nor U859 (N_859,N_780,N_765);
nand U860 (N_860,N_764,N_800);
nand U861 (N_861,N_778,N_786);
or U862 (N_862,N_811,N_799);
nor U863 (N_863,N_771,N_783);
and U864 (N_864,N_824,N_794);
and U865 (N_865,N_774,N_775);
and U866 (N_866,N_796,N_758);
nor U867 (N_867,N_819,N_817);
and U868 (N_868,N_752,N_764);
and U869 (N_869,N_769,N_791);
nand U870 (N_870,N_788,N_810);
nand U871 (N_871,N_760,N_798);
and U872 (N_872,N_779,N_781);
nor U873 (N_873,N_822,N_802);
or U874 (N_874,N_763,N_814);
nand U875 (N_875,N_765,N_824);
and U876 (N_876,N_784,N_805);
nor U877 (N_877,N_762,N_775);
or U878 (N_878,N_759,N_792);
nor U879 (N_879,N_819,N_776);
nor U880 (N_880,N_822,N_768);
or U881 (N_881,N_775,N_764);
or U882 (N_882,N_763,N_783);
nor U883 (N_883,N_765,N_794);
and U884 (N_884,N_789,N_775);
nor U885 (N_885,N_823,N_752);
nand U886 (N_886,N_821,N_789);
or U887 (N_887,N_764,N_791);
and U888 (N_888,N_823,N_803);
nor U889 (N_889,N_768,N_751);
nor U890 (N_890,N_821,N_788);
nand U891 (N_891,N_783,N_756);
and U892 (N_892,N_771,N_813);
and U893 (N_893,N_812,N_806);
and U894 (N_894,N_762,N_757);
nand U895 (N_895,N_806,N_815);
or U896 (N_896,N_771,N_774);
nor U897 (N_897,N_760,N_808);
nand U898 (N_898,N_820,N_764);
and U899 (N_899,N_751,N_822);
and U900 (N_900,N_863,N_849);
nor U901 (N_901,N_892,N_867);
and U902 (N_902,N_872,N_862);
and U903 (N_903,N_847,N_848);
nor U904 (N_904,N_875,N_885);
and U905 (N_905,N_853,N_858);
nor U906 (N_906,N_890,N_883);
or U907 (N_907,N_845,N_854);
and U908 (N_908,N_881,N_865);
nor U909 (N_909,N_864,N_869);
and U910 (N_910,N_846,N_878);
and U911 (N_911,N_899,N_832);
nor U912 (N_912,N_888,N_859);
or U913 (N_913,N_861,N_837);
and U914 (N_914,N_886,N_828);
xor U915 (N_915,N_884,N_839);
or U916 (N_916,N_838,N_827);
and U917 (N_917,N_893,N_830);
nor U918 (N_918,N_882,N_834);
or U919 (N_919,N_877,N_836);
or U920 (N_920,N_873,N_840);
and U921 (N_921,N_855,N_874);
nand U922 (N_922,N_835,N_895);
or U923 (N_923,N_879,N_829);
and U924 (N_924,N_851,N_826);
or U925 (N_925,N_843,N_844);
nor U926 (N_926,N_842,N_831);
nand U927 (N_927,N_860,N_868);
and U928 (N_928,N_894,N_870);
or U929 (N_929,N_880,N_866);
nand U930 (N_930,N_876,N_833);
nor U931 (N_931,N_871,N_896);
and U932 (N_932,N_856,N_887);
nor U933 (N_933,N_891,N_841);
nand U934 (N_934,N_889,N_825);
nand U935 (N_935,N_852,N_898);
xor U936 (N_936,N_857,N_897);
nand U937 (N_937,N_850,N_826);
nand U938 (N_938,N_898,N_883);
and U939 (N_939,N_870,N_876);
nor U940 (N_940,N_867,N_863);
nand U941 (N_941,N_899,N_885);
nand U942 (N_942,N_837,N_897);
nor U943 (N_943,N_833,N_896);
nor U944 (N_944,N_896,N_891);
nand U945 (N_945,N_861,N_875);
nor U946 (N_946,N_881,N_831);
nand U947 (N_947,N_879,N_834);
and U948 (N_948,N_826,N_835);
nand U949 (N_949,N_855,N_893);
nor U950 (N_950,N_856,N_826);
and U951 (N_951,N_844,N_873);
nand U952 (N_952,N_880,N_838);
or U953 (N_953,N_829,N_870);
nor U954 (N_954,N_845,N_852);
nand U955 (N_955,N_854,N_895);
and U956 (N_956,N_858,N_837);
nor U957 (N_957,N_830,N_863);
nand U958 (N_958,N_858,N_865);
nand U959 (N_959,N_891,N_898);
nor U960 (N_960,N_895,N_827);
or U961 (N_961,N_844,N_877);
nor U962 (N_962,N_898,N_830);
or U963 (N_963,N_850,N_897);
or U964 (N_964,N_885,N_848);
nand U965 (N_965,N_880,N_836);
nand U966 (N_966,N_855,N_870);
nor U967 (N_967,N_880,N_831);
and U968 (N_968,N_846,N_897);
or U969 (N_969,N_872,N_889);
and U970 (N_970,N_882,N_846);
nand U971 (N_971,N_832,N_845);
and U972 (N_972,N_862,N_843);
nor U973 (N_973,N_865,N_840);
or U974 (N_974,N_876,N_854);
and U975 (N_975,N_935,N_940);
and U976 (N_976,N_902,N_904);
nand U977 (N_977,N_901,N_954);
or U978 (N_978,N_907,N_928);
and U979 (N_979,N_934,N_958);
or U980 (N_980,N_944,N_953);
or U981 (N_981,N_906,N_945);
and U982 (N_982,N_922,N_970);
nand U983 (N_983,N_929,N_947);
or U984 (N_984,N_972,N_921);
and U985 (N_985,N_925,N_961);
and U986 (N_986,N_914,N_967);
nand U987 (N_987,N_938,N_943);
nand U988 (N_988,N_962,N_930);
or U989 (N_989,N_923,N_951);
and U990 (N_990,N_920,N_908);
and U991 (N_991,N_971,N_926);
nand U992 (N_992,N_941,N_910);
nand U993 (N_993,N_939,N_964);
nand U994 (N_994,N_927,N_932);
and U995 (N_995,N_973,N_905);
nor U996 (N_996,N_949,N_919);
nor U997 (N_997,N_955,N_912);
nand U998 (N_998,N_900,N_931);
and U999 (N_999,N_950,N_948);
and U1000 (N_1000,N_965,N_942);
or U1001 (N_1001,N_936,N_937);
or U1002 (N_1002,N_915,N_933);
and U1003 (N_1003,N_963,N_974);
nor U1004 (N_1004,N_968,N_917);
nor U1005 (N_1005,N_911,N_960);
nor U1006 (N_1006,N_913,N_969);
and U1007 (N_1007,N_959,N_903);
or U1008 (N_1008,N_924,N_918);
nor U1009 (N_1009,N_916,N_952);
or U1010 (N_1010,N_909,N_956);
nor U1011 (N_1011,N_957,N_946);
nand U1012 (N_1012,N_966,N_950);
and U1013 (N_1013,N_914,N_917);
nand U1014 (N_1014,N_965,N_958);
nand U1015 (N_1015,N_913,N_919);
nor U1016 (N_1016,N_973,N_922);
or U1017 (N_1017,N_937,N_974);
or U1018 (N_1018,N_957,N_965);
nor U1019 (N_1019,N_969,N_964);
nor U1020 (N_1020,N_958,N_929);
and U1021 (N_1021,N_934,N_940);
or U1022 (N_1022,N_974,N_935);
and U1023 (N_1023,N_930,N_947);
nor U1024 (N_1024,N_915,N_967);
nand U1025 (N_1025,N_929,N_915);
or U1026 (N_1026,N_937,N_915);
and U1027 (N_1027,N_952,N_970);
and U1028 (N_1028,N_950,N_955);
or U1029 (N_1029,N_913,N_922);
nor U1030 (N_1030,N_921,N_971);
nand U1031 (N_1031,N_963,N_932);
nand U1032 (N_1032,N_943,N_913);
nand U1033 (N_1033,N_900,N_959);
nor U1034 (N_1034,N_916,N_958);
or U1035 (N_1035,N_973,N_928);
nor U1036 (N_1036,N_956,N_920);
nand U1037 (N_1037,N_927,N_914);
or U1038 (N_1038,N_929,N_962);
or U1039 (N_1039,N_943,N_951);
and U1040 (N_1040,N_956,N_940);
and U1041 (N_1041,N_970,N_913);
nor U1042 (N_1042,N_913,N_927);
nand U1043 (N_1043,N_970,N_968);
or U1044 (N_1044,N_945,N_957);
nand U1045 (N_1045,N_907,N_972);
and U1046 (N_1046,N_933,N_923);
and U1047 (N_1047,N_921,N_926);
nor U1048 (N_1048,N_909,N_949);
nand U1049 (N_1049,N_969,N_910);
nor U1050 (N_1050,N_1016,N_978);
nand U1051 (N_1051,N_1048,N_1004);
nand U1052 (N_1052,N_1034,N_998);
nor U1053 (N_1053,N_979,N_1047);
and U1054 (N_1054,N_1039,N_1040);
and U1055 (N_1055,N_1044,N_996);
nand U1056 (N_1056,N_983,N_1037);
nor U1057 (N_1057,N_1018,N_988);
nor U1058 (N_1058,N_1036,N_1003);
or U1059 (N_1059,N_1026,N_993);
nand U1060 (N_1060,N_976,N_1024);
nor U1061 (N_1061,N_1027,N_997);
or U1062 (N_1062,N_977,N_1042);
nand U1063 (N_1063,N_1017,N_1049);
and U1064 (N_1064,N_985,N_1020);
nand U1065 (N_1065,N_1001,N_1012);
nor U1066 (N_1066,N_992,N_1009);
and U1067 (N_1067,N_1041,N_987);
or U1068 (N_1068,N_1022,N_1014);
or U1069 (N_1069,N_999,N_980);
nor U1070 (N_1070,N_1045,N_1013);
or U1071 (N_1071,N_1046,N_1032);
nor U1072 (N_1072,N_1043,N_1010);
or U1073 (N_1073,N_1028,N_1035);
or U1074 (N_1074,N_995,N_1011);
or U1075 (N_1075,N_1025,N_975);
nand U1076 (N_1076,N_986,N_1002);
nand U1077 (N_1077,N_1008,N_1019);
nor U1078 (N_1078,N_1005,N_982);
nand U1079 (N_1079,N_990,N_994);
or U1080 (N_1080,N_981,N_1015);
or U1081 (N_1081,N_1029,N_1006);
nand U1082 (N_1082,N_1038,N_991);
or U1083 (N_1083,N_1031,N_1000);
nor U1084 (N_1084,N_989,N_1033);
nand U1085 (N_1085,N_1007,N_1023);
and U1086 (N_1086,N_1021,N_984);
or U1087 (N_1087,N_1030,N_999);
or U1088 (N_1088,N_987,N_1018);
nand U1089 (N_1089,N_1009,N_1030);
and U1090 (N_1090,N_984,N_999);
nand U1091 (N_1091,N_996,N_1001);
nor U1092 (N_1092,N_1030,N_1036);
nand U1093 (N_1093,N_1000,N_1046);
nand U1094 (N_1094,N_990,N_1027);
or U1095 (N_1095,N_989,N_1042);
nand U1096 (N_1096,N_1033,N_991);
nor U1097 (N_1097,N_1011,N_998);
and U1098 (N_1098,N_1039,N_1037);
and U1099 (N_1099,N_1005,N_1018);
or U1100 (N_1100,N_1019,N_1037);
or U1101 (N_1101,N_1047,N_990);
nand U1102 (N_1102,N_1049,N_1031);
or U1103 (N_1103,N_1023,N_1013);
nand U1104 (N_1104,N_1023,N_995);
and U1105 (N_1105,N_984,N_1022);
or U1106 (N_1106,N_1047,N_1043);
or U1107 (N_1107,N_995,N_1005);
nand U1108 (N_1108,N_977,N_1048);
or U1109 (N_1109,N_1042,N_1025);
nor U1110 (N_1110,N_1007,N_1027);
nand U1111 (N_1111,N_1002,N_1041);
or U1112 (N_1112,N_1003,N_1015);
nand U1113 (N_1113,N_1037,N_1043);
and U1114 (N_1114,N_1011,N_1032);
and U1115 (N_1115,N_983,N_1021);
nor U1116 (N_1116,N_1040,N_1002);
nand U1117 (N_1117,N_986,N_1029);
and U1118 (N_1118,N_1029,N_1033);
or U1119 (N_1119,N_977,N_1008);
nor U1120 (N_1120,N_1006,N_1017);
nand U1121 (N_1121,N_984,N_978);
and U1122 (N_1122,N_994,N_979);
and U1123 (N_1123,N_1013,N_984);
xnor U1124 (N_1124,N_997,N_1018);
and U1125 (N_1125,N_1114,N_1108);
or U1126 (N_1126,N_1100,N_1103);
nand U1127 (N_1127,N_1062,N_1123);
nand U1128 (N_1128,N_1084,N_1056);
nand U1129 (N_1129,N_1051,N_1065);
and U1130 (N_1130,N_1055,N_1104);
and U1131 (N_1131,N_1119,N_1057);
and U1132 (N_1132,N_1080,N_1081);
or U1133 (N_1133,N_1111,N_1068);
or U1134 (N_1134,N_1106,N_1107);
or U1135 (N_1135,N_1096,N_1063);
nand U1136 (N_1136,N_1090,N_1079);
nand U1137 (N_1137,N_1085,N_1122);
nand U1138 (N_1138,N_1083,N_1101);
and U1139 (N_1139,N_1077,N_1121);
and U1140 (N_1140,N_1060,N_1117);
nand U1141 (N_1141,N_1124,N_1087);
nand U1142 (N_1142,N_1071,N_1078);
nor U1143 (N_1143,N_1058,N_1112);
nand U1144 (N_1144,N_1109,N_1053);
or U1145 (N_1145,N_1105,N_1088);
or U1146 (N_1146,N_1099,N_1089);
nor U1147 (N_1147,N_1095,N_1072);
or U1148 (N_1148,N_1098,N_1120);
nor U1149 (N_1149,N_1094,N_1061);
nor U1150 (N_1150,N_1115,N_1074);
nand U1151 (N_1151,N_1073,N_1093);
nand U1152 (N_1152,N_1097,N_1086);
or U1153 (N_1153,N_1102,N_1075);
or U1154 (N_1154,N_1116,N_1118);
xor U1155 (N_1155,N_1113,N_1066);
or U1156 (N_1156,N_1092,N_1069);
or U1157 (N_1157,N_1076,N_1091);
nor U1158 (N_1158,N_1070,N_1052);
or U1159 (N_1159,N_1110,N_1082);
and U1160 (N_1160,N_1064,N_1067);
nand U1161 (N_1161,N_1050,N_1054);
nor U1162 (N_1162,N_1059,N_1105);
nor U1163 (N_1163,N_1095,N_1085);
xnor U1164 (N_1164,N_1084,N_1089);
nand U1165 (N_1165,N_1113,N_1116);
xnor U1166 (N_1166,N_1053,N_1081);
or U1167 (N_1167,N_1080,N_1053);
nand U1168 (N_1168,N_1076,N_1064);
nor U1169 (N_1169,N_1053,N_1122);
and U1170 (N_1170,N_1091,N_1068);
nor U1171 (N_1171,N_1124,N_1104);
and U1172 (N_1172,N_1088,N_1094);
nand U1173 (N_1173,N_1115,N_1097);
nor U1174 (N_1174,N_1066,N_1106);
nor U1175 (N_1175,N_1065,N_1097);
nor U1176 (N_1176,N_1090,N_1060);
and U1177 (N_1177,N_1093,N_1089);
nand U1178 (N_1178,N_1108,N_1083);
nand U1179 (N_1179,N_1079,N_1097);
nor U1180 (N_1180,N_1112,N_1097);
nor U1181 (N_1181,N_1064,N_1123);
and U1182 (N_1182,N_1051,N_1091);
and U1183 (N_1183,N_1111,N_1121);
nand U1184 (N_1184,N_1065,N_1123);
and U1185 (N_1185,N_1107,N_1091);
nor U1186 (N_1186,N_1066,N_1114);
nor U1187 (N_1187,N_1092,N_1066);
or U1188 (N_1188,N_1050,N_1099);
and U1189 (N_1189,N_1072,N_1098);
and U1190 (N_1190,N_1073,N_1062);
nor U1191 (N_1191,N_1079,N_1082);
nand U1192 (N_1192,N_1058,N_1123);
nand U1193 (N_1193,N_1067,N_1071);
nor U1194 (N_1194,N_1069,N_1096);
nand U1195 (N_1195,N_1117,N_1113);
nor U1196 (N_1196,N_1053,N_1104);
nor U1197 (N_1197,N_1124,N_1099);
nor U1198 (N_1198,N_1071,N_1080);
and U1199 (N_1199,N_1055,N_1101);
or U1200 (N_1200,N_1188,N_1193);
or U1201 (N_1201,N_1159,N_1138);
nand U1202 (N_1202,N_1194,N_1127);
nand U1203 (N_1203,N_1152,N_1175);
or U1204 (N_1204,N_1148,N_1158);
nand U1205 (N_1205,N_1179,N_1198);
nand U1206 (N_1206,N_1182,N_1183);
nand U1207 (N_1207,N_1176,N_1170);
nor U1208 (N_1208,N_1162,N_1149);
nand U1209 (N_1209,N_1147,N_1143);
nand U1210 (N_1210,N_1191,N_1199);
or U1211 (N_1211,N_1155,N_1144);
nand U1212 (N_1212,N_1146,N_1136);
and U1213 (N_1213,N_1139,N_1151);
nor U1214 (N_1214,N_1184,N_1131);
nand U1215 (N_1215,N_1137,N_1186);
nor U1216 (N_1216,N_1140,N_1187);
nand U1217 (N_1217,N_1161,N_1141);
or U1218 (N_1218,N_1157,N_1180);
nor U1219 (N_1219,N_1132,N_1166);
or U1220 (N_1220,N_1142,N_1167);
or U1221 (N_1221,N_1195,N_1171);
or U1222 (N_1222,N_1134,N_1168);
nor U1223 (N_1223,N_1192,N_1196);
or U1224 (N_1224,N_1130,N_1154);
and U1225 (N_1225,N_1160,N_1150);
nor U1226 (N_1226,N_1165,N_1164);
and U1227 (N_1227,N_1125,N_1181);
nand U1228 (N_1228,N_1163,N_1128);
nand U1229 (N_1229,N_1129,N_1172);
nor U1230 (N_1230,N_1174,N_1178);
and U1231 (N_1231,N_1197,N_1185);
nor U1232 (N_1232,N_1177,N_1156);
or U1233 (N_1233,N_1169,N_1133);
nand U1234 (N_1234,N_1145,N_1190);
nand U1235 (N_1235,N_1189,N_1135);
nand U1236 (N_1236,N_1126,N_1153);
or U1237 (N_1237,N_1173,N_1129);
nor U1238 (N_1238,N_1165,N_1173);
nand U1239 (N_1239,N_1138,N_1144);
nand U1240 (N_1240,N_1197,N_1152);
or U1241 (N_1241,N_1138,N_1168);
or U1242 (N_1242,N_1167,N_1151);
and U1243 (N_1243,N_1139,N_1175);
nor U1244 (N_1244,N_1197,N_1142);
or U1245 (N_1245,N_1185,N_1180);
nor U1246 (N_1246,N_1133,N_1185);
or U1247 (N_1247,N_1164,N_1187);
nand U1248 (N_1248,N_1149,N_1161);
or U1249 (N_1249,N_1160,N_1149);
nor U1250 (N_1250,N_1145,N_1196);
nand U1251 (N_1251,N_1154,N_1161);
and U1252 (N_1252,N_1150,N_1196);
nand U1253 (N_1253,N_1162,N_1189);
nand U1254 (N_1254,N_1162,N_1130);
nand U1255 (N_1255,N_1187,N_1130);
xnor U1256 (N_1256,N_1139,N_1141);
nand U1257 (N_1257,N_1139,N_1146);
nand U1258 (N_1258,N_1196,N_1178);
nand U1259 (N_1259,N_1192,N_1168);
and U1260 (N_1260,N_1159,N_1184);
and U1261 (N_1261,N_1155,N_1197);
or U1262 (N_1262,N_1172,N_1188);
nand U1263 (N_1263,N_1183,N_1140);
nand U1264 (N_1264,N_1149,N_1153);
and U1265 (N_1265,N_1194,N_1162);
nor U1266 (N_1266,N_1153,N_1156);
nor U1267 (N_1267,N_1178,N_1136);
nand U1268 (N_1268,N_1132,N_1191);
and U1269 (N_1269,N_1164,N_1126);
nor U1270 (N_1270,N_1148,N_1170);
nor U1271 (N_1271,N_1148,N_1189);
and U1272 (N_1272,N_1174,N_1156);
nor U1273 (N_1273,N_1135,N_1179);
nand U1274 (N_1274,N_1171,N_1129);
and U1275 (N_1275,N_1265,N_1202);
nor U1276 (N_1276,N_1248,N_1271);
or U1277 (N_1277,N_1228,N_1206);
or U1278 (N_1278,N_1229,N_1211);
nor U1279 (N_1279,N_1230,N_1263);
nor U1280 (N_1280,N_1270,N_1221);
nor U1281 (N_1281,N_1269,N_1251);
or U1282 (N_1282,N_1255,N_1236);
and U1283 (N_1283,N_1258,N_1247);
nor U1284 (N_1284,N_1226,N_1253);
nand U1285 (N_1285,N_1240,N_1242);
nor U1286 (N_1286,N_1266,N_1220);
and U1287 (N_1287,N_1201,N_1231);
nand U1288 (N_1288,N_1264,N_1259);
nor U1289 (N_1289,N_1203,N_1207);
and U1290 (N_1290,N_1217,N_1239);
nor U1291 (N_1291,N_1254,N_1274);
nor U1292 (N_1292,N_1232,N_1235);
and U1293 (N_1293,N_1245,N_1219);
nor U1294 (N_1294,N_1273,N_1218);
and U1295 (N_1295,N_1214,N_1272);
nor U1296 (N_1296,N_1200,N_1249);
and U1297 (N_1297,N_1222,N_1243);
or U1298 (N_1298,N_1204,N_1257);
nor U1299 (N_1299,N_1210,N_1261);
and U1300 (N_1300,N_1238,N_1246);
nand U1301 (N_1301,N_1244,N_1227);
nand U1302 (N_1302,N_1213,N_1209);
nand U1303 (N_1303,N_1237,N_1260);
and U1304 (N_1304,N_1241,N_1224);
nor U1305 (N_1305,N_1205,N_1215);
nor U1306 (N_1306,N_1256,N_1225);
or U1307 (N_1307,N_1262,N_1250);
and U1308 (N_1308,N_1223,N_1268);
nor U1309 (N_1309,N_1212,N_1216);
or U1310 (N_1310,N_1267,N_1252);
or U1311 (N_1311,N_1208,N_1233);
nand U1312 (N_1312,N_1234,N_1210);
or U1313 (N_1313,N_1218,N_1209);
nor U1314 (N_1314,N_1257,N_1218);
nand U1315 (N_1315,N_1230,N_1214);
nor U1316 (N_1316,N_1207,N_1210);
or U1317 (N_1317,N_1223,N_1201);
and U1318 (N_1318,N_1266,N_1251);
nand U1319 (N_1319,N_1215,N_1269);
nor U1320 (N_1320,N_1210,N_1233);
or U1321 (N_1321,N_1268,N_1214);
nor U1322 (N_1322,N_1266,N_1256);
nor U1323 (N_1323,N_1257,N_1260);
or U1324 (N_1324,N_1245,N_1227);
nor U1325 (N_1325,N_1213,N_1270);
nand U1326 (N_1326,N_1241,N_1220);
and U1327 (N_1327,N_1231,N_1232);
and U1328 (N_1328,N_1245,N_1241);
nand U1329 (N_1329,N_1251,N_1261);
nor U1330 (N_1330,N_1231,N_1206);
nand U1331 (N_1331,N_1273,N_1203);
nand U1332 (N_1332,N_1227,N_1239);
nand U1333 (N_1333,N_1232,N_1220);
nor U1334 (N_1334,N_1208,N_1207);
nand U1335 (N_1335,N_1219,N_1265);
and U1336 (N_1336,N_1241,N_1267);
nand U1337 (N_1337,N_1220,N_1204);
nor U1338 (N_1338,N_1201,N_1235);
and U1339 (N_1339,N_1252,N_1204);
nand U1340 (N_1340,N_1231,N_1214);
and U1341 (N_1341,N_1205,N_1253);
or U1342 (N_1342,N_1248,N_1228);
or U1343 (N_1343,N_1245,N_1211);
or U1344 (N_1344,N_1250,N_1228);
or U1345 (N_1345,N_1245,N_1259);
or U1346 (N_1346,N_1224,N_1246);
nor U1347 (N_1347,N_1259,N_1266);
nor U1348 (N_1348,N_1249,N_1244);
nor U1349 (N_1349,N_1250,N_1266);
and U1350 (N_1350,N_1346,N_1331);
and U1351 (N_1351,N_1283,N_1342);
or U1352 (N_1352,N_1280,N_1344);
nor U1353 (N_1353,N_1315,N_1275);
or U1354 (N_1354,N_1335,N_1294);
or U1355 (N_1355,N_1298,N_1345);
and U1356 (N_1356,N_1328,N_1299);
or U1357 (N_1357,N_1301,N_1313);
nand U1358 (N_1358,N_1277,N_1293);
and U1359 (N_1359,N_1310,N_1326);
or U1360 (N_1360,N_1324,N_1305);
or U1361 (N_1361,N_1281,N_1291);
or U1362 (N_1362,N_1314,N_1312);
nor U1363 (N_1363,N_1336,N_1284);
and U1364 (N_1364,N_1279,N_1286);
and U1365 (N_1365,N_1289,N_1347);
or U1366 (N_1366,N_1318,N_1292);
or U1367 (N_1367,N_1341,N_1329);
nor U1368 (N_1368,N_1285,N_1332);
or U1369 (N_1369,N_1296,N_1311);
nand U1370 (N_1370,N_1316,N_1303);
nor U1371 (N_1371,N_1340,N_1323);
and U1372 (N_1372,N_1295,N_1278);
nor U1373 (N_1373,N_1349,N_1297);
or U1374 (N_1374,N_1304,N_1330);
or U1375 (N_1375,N_1327,N_1276);
or U1376 (N_1376,N_1287,N_1348);
and U1377 (N_1377,N_1321,N_1300);
nor U1378 (N_1378,N_1339,N_1334);
nor U1379 (N_1379,N_1308,N_1306);
nand U1380 (N_1380,N_1343,N_1333);
and U1381 (N_1381,N_1282,N_1337);
nand U1382 (N_1382,N_1302,N_1307);
nor U1383 (N_1383,N_1320,N_1290);
nor U1384 (N_1384,N_1325,N_1338);
and U1385 (N_1385,N_1317,N_1309);
and U1386 (N_1386,N_1322,N_1319);
and U1387 (N_1387,N_1288,N_1338);
nand U1388 (N_1388,N_1285,N_1326);
nand U1389 (N_1389,N_1276,N_1300);
and U1390 (N_1390,N_1313,N_1341);
nand U1391 (N_1391,N_1297,N_1280);
nor U1392 (N_1392,N_1314,N_1301);
nor U1393 (N_1393,N_1346,N_1320);
and U1394 (N_1394,N_1336,N_1288);
nand U1395 (N_1395,N_1325,N_1297);
nor U1396 (N_1396,N_1308,N_1282);
nand U1397 (N_1397,N_1288,N_1312);
nand U1398 (N_1398,N_1300,N_1345);
nor U1399 (N_1399,N_1289,N_1304);
and U1400 (N_1400,N_1324,N_1284);
or U1401 (N_1401,N_1349,N_1292);
nand U1402 (N_1402,N_1326,N_1331);
and U1403 (N_1403,N_1343,N_1293);
and U1404 (N_1404,N_1306,N_1322);
nand U1405 (N_1405,N_1341,N_1304);
and U1406 (N_1406,N_1295,N_1307);
nand U1407 (N_1407,N_1288,N_1300);
and U1408 (N_1408,N_1319,N_1348);
nand U1409 (N_1409,N_1329,N_1287);
nand U1410 (N_1410,N_1308,N_1281);
nor U1411 (N_1411,N_1325,N_1323);
nand U1412 (N_1412,N_1318,N_1335);
or U1413 (N_1413,N_1308,N_1342);
and U1414 (N_1414,N_1281,N_1296);
nor U1415 (N_1415,N_1294,N_1296);
or U1416 (N_1416,N_1275,N_1298);
nor U1417 (N_1417,N_1346,N_1343);
nand U1418 (N_1418,N_1301,N_1345);
or U1419 (N_1419,N_1342,N_1335);
or U1420 (N_1420,N_1323,N_1345);
or U1421 (N_1421,N_1334,N_1328);
nand U1422 (N_1422,N_1278,N_1339);
or U1423 (N_1423,N_1291,N_1345);
nor U1424 (N_1424,N_1336,N_1287);
nand U1425 (N_1425,N_1363,N_1406);
nand U1426 (N_1426,N_1386,N_1381);
or U1427 (N_1427,N_1411,N_1396);
nor U1428 (N_1428,N_1355,N_1359);
and U1429 (N_1429,N_1401,N_1416);
nor U1430 (N_1430,N_1391,N_1398);
nand U1431 (N_1431,N_1418,N_1421);
or U1432 (N_1432,N_1413,N_1387);
or U1433 (N_1433,N_1390,N_1392);
or U1434 (N_1434,N_1376,N_1384);
nand U1435 (N_1435,N_1415,N_1383);
or U1436 (N_1436,N_1400,N_1380);
and U1437 (N_1437,N_1373,N_1375);
or U1438 (N_1438,N_1368,N_1369);
nand U1439 (N_1439,N_1402,N_1361);
or U1440 (N_1440,N_1409,N_1422);
and U1441 (N_1441,N_1420,N_1372);
nor U1442 (N_1442,N_1352,N_1388);
or U1443 (N_1443,N_1407,N_1385);
and U1444 (N_1444,N_1389,N_1367);
or U1445 (N_1445,N_1357,N_1371);
or U1446 (N_1446,N_1365,N_1423);
nand U1447 (N_1447,N_1405,N_1412);
nor U1448 (N_1448,N_1410,N_1377);
nor U1449 (N_1449,N_1382,N_1393);
and U1450 (N_1450,N_1362,N_1414);
nor U1451 (N_1451,N_1424,N_1378);
or U1452 (N_1452,N_1358,N_1397);
or U1453 (N_1453,N_1350,N_1366);
or U1454 (N_1454,N_1399,N_1404);
nand U1455 (N_1455,N_1408,N_1417);
nor U1456 (N_1456,N_1403,N_1374);
nor U1457 (N_1457,N_1379,N_1360);
nand U1458 (N_1458,N_1354,N_1351);
nand U1459 (N_1459,N_1395,N_1356);
nand U1460 (N_1460,N_1370,N_1394);
or U1461 (N_1461,N_1364,N_1419);
nor U1462 (N_1462,N_1353,N_1377);
nor U1463 (N_1463,N_1404,N_1376);
and U1464 (N_1464,N_1420,N_1386);
nor U1465 (N_1465,N_1397,N_1411);
nand U1466 (N_1466,N_1355,N_1363);
nor U1467 (N_1467,N_1364,N_1407);
or U1468 (N_1468,N_1397,N_1391);
nor U1469 (N_1469,N_1351,N_1372);
nor U1470 (N_1470,N_1385,N_1384);
and U1471 (N_1471,N_1352,N_1401);
or U1472 (N_1472,N_1417,N_1422);
and U1473 (N_1473,N_1350,N_1410);
nor U1474 (N_1474,N_1398,N_1386);
or U1475 (N_1475,N_1392,N_1350);
nand U1476 (N_1476,N_1381,N_1424);
nand U1477 (N_1477,N_1417,N_1412);
nor U1478 (N_1478,N_1351,N_1422);
nand U1479 (N_1479,N_1355,N_1382);
or U1480 (N_1480,N_1406,N_1422);
or U1481 (N_1481,N_1366,N_1408);
and U1482 (N_1482,N_1362,N_1371);
nor U1483 (N_1483,N_1424,N_1365);
nand U1484 (N_1484,N_1360,N_1402);
nand U1485 (N_1485,N_1397,N_1419);
nor U1486 (N_1486,N_1380,N_1350);
nor U1487 (N_1487,N_1393,N_1379);
nand U1488 (N_1488,N_1369,N_1377);
nor U1489 (N_1489,N_1405,N_1371);
xor U1490 (N_1490,N_1366,N_1355);
and U1491 (N_1491,N_1420,N_1353);
nor U1492 (N_1492,N_1401,N_1366);
nor U1493 (N_1493,N_1366,N_1390);
or U1494 (N_1494,N_1391,N_1370);
nor U1495 (N_1495,N_1418,N_1350);
and U1496 (N_1496,N_1391,N_1360);
nand U1497 (N_1497,N_1382,N_1350);
or U1498 (N_1498,N_1409,N_1397);
or U1499 (N_1499,N_1405,N_1403);
nand U1500 (N_1500,N_1427,N_1492);
nand U1501 (N_1501,N_1486,N_1462);
and U1502 (N_1502,N_1442,N_1434);
nand U1503 (N_1503,N_1432,N_1474);
nand U1504 (N_1504,N_1477,N_1482);
nor U1505 (N_1505,N_1478,N_1438);
and U1506 (N_1506,N_1449,N_1458);
nor U1507 (N_1507,N_1448,N_1472);
nand U1508 (N_1508,N_1465,N_1476);
nand U1509 (N_1509,N_1431,N_1461);
nor U1510 (N_1510,N_1452,N_1490);
nand U1511 (N_1511,N_1495,N_1436);
and U1512 (N_1512,N_1426,N_1473);
nand U1513 (N_1513,N_1439,N_1450);
nor U1514 (N_1514,N_1466,N_1493);
nor U1515 (N_1515,N_1446,N_1491);
nor U1516 (N_1516,N_1484,N_1460);
nor U1517 (N_1517,N_1463,N_1430);
or U1518 (N_1518,N_1457,N_1459);
and U1519 (N_1519,N_1428,N_1468);
or U1520 (N_1520,N_1489,N_1487);
and U1521 (N_1521,N_1443,N_1455);
nand U1522 (N_1522,N_1437,N_1494);
or U1523 (N_1523,N_1425,N_1498);
or U1524 (N_1524,N_1456,N_1475);
nand U1525 (N_1525,N_1499,N_1470);
nor U1526 (N_1526,N_1471,N_1467);
nor U1527 (N_1527,N_1481,N_1435);
and U1528 (N_1528,N_1429,N_1444);
or U1529 (N_1529,N_1469,N_1454);
and U1530 (N_1530,N_1447,N_1451);
and U1531 (N_1531,N_1488,N_1483);
and U1532 (N_1532,N_1445,N_1433);
and U1533 (N_1533,N_1441,N_1479);
nor U1534 (N_1534,N_1464,N_1497);
and U1535 (N_1535,N_1496,N_1440);
nor U1536 (N_1536,N_1453,N_1485);
and U1537 (N_1537,N_1480,N_1461);
and U1538 (N_1538,N_1447,N_1432);
and U1539 (N_1539,N_1431,N_1434);
and U1540 (N_1540,N_1445,N_1436);
nor U1541 (N_1541,N_1460,N_1481);
or U1542 (N_1542,N_1458,N_1461);
nand U1543 (N_1543,N_1438,N_1441);
or U1544 (N_1544,N_1491,N_1464);
nor U1545 (N_1545,N_1490,N_1487);
or U1546 (N_1546,N_1469,N_1473);
and U1547 (N_1547,N_1471,N_1425);
nor U1548 (N_1548,N_1471,N_1438);
and U1549 (N_1549,N_1452,N_1499);
or U1550 (N_1550,N_1462,N_1434);
or U1551 (N_1551,N_1435,N_1474);
nand U1552 (N_1552,N_1487,N_1485);
or U1553 (N_1553,N_1452,N_1436);
or U1554 (N_1554,N_1441,N_1475);
nor U1555 (N_1555,N_1494,N_1444);
or U1556 (N_1556,N_1487,N_1444);
nand U1557 (N_1557,N_1492,N_1428);
xor U1558 (N_1558,N_1441,N_1486);
nor U1559 (N_1559,N_1496,N_1463);
and U1560 (N_1560,N_1480,N_1442);
or U1561 (N_1561,N_1479,N_1439);
or U1562 (N_1562,N_1474,N_1457);
or U1563 (N_1563,N_1469,N_1453);
nor U1564 (N_1564,N_1440,N_1481);
nor U1565 (N_1565,N_1473,N_1487);
nor U1566 (N_1566,N_1480,N_1427);
or U1567 (N_1567,N_1476,N_1474);
and U1568 (N_1568,N_1438,N_1488);
or U1569 (N_1569,N_1497,N_1448);
nand U1570 (N_1570,N_1498,N_1466);
and U1571 (N_1571,N_1431,N_1438);
nor U1572 (N_1572,N_1479,N_1477);
nor U1573 (N_1573,N_1480,N_1484);
nand U1574 (N_1574,N_1463,N_1443);
nor U1575 (N_1575,N_1572,N_1557);
and U1576 (N_1576,N_1534,N_1554);
nand U1577 (N_1577,N_1523,N_1556);
or U1578 (N_1578,N_1511,N_1555);
nor U1579 (N_1579,N_1569,N_1528);
nor U1580 (N_1580,N_1562,N_1500);
or U1581 (N_1581,N_1549,N_1573);
nand U1582 (N_1582,N_1529,N_1507);
nand U1583 (N_1583,N_1568,N_1544);
and U1584 (N_1584,N_1543,N_1503);
nand U1585 (N_1585,N_1564,N_1530);
or U1586 (N_1586,N_1552,N_1533);
nand U1587 (N_1587,N_1525,N_1535);
and U1588 (N_1588,N_1551,N_1548);
nor U1589 (N_1589,N_1515,N_1553);
nor U1590 (N_1590,N_1541,N_1524);
and U1591 (N_1591,N_1522,N_1514);
or U1592 (N_1592,N_1539,N_1558);
nand U1593 (N_1593,N_1542,N_1532);
or U1594 (N_1594,N_1537,N_1567);
and U1595 (N_1595,N_1570,N_1510);
or U1596 (N_1596,N_1559,N_1508);
nor U1597 (N_1597,N_1536,N_1563);
and U1598 (N_1598,N_1512,N_1571);
or U1599 (N_1599,N_1531,N_1546);
nor U1600 (N_1600,N_1509,N_1566);
nand U1601 (N_1601,N_1513,N_1520);
nor U1602 (N_1602,N_1506,N_1547);
nand U1603 (N_1603,N_1502,N_1565);
and U1604 (N_1604,N_1501,N_1550);
nor U1605 (N_1605,N_1560,N_1521);
nor U1606 (N_1606,N_1538,N_1504);
nor U1607 (N_1607,N_1527,N_1526);
and U1608 (N_1608,N_1561,N_1545);
or U1609 (N_1609,N_1516,N_1517);
nand U1610 (N_1610,N_1505,N_1519);
nor U1611 (N_1611,N_1540,N_1574);
and U1612 (N_1612,N_1518,N_1532);
nor U1613 (N_1613,N_1539,N_1534);
and U1614 (N_1614,N_1559,N_1557);
nor U1615 (N_1615,N_1529,N_1519);
nor U1616 (N_1616,N_1509,N_1504);
or U1617 (N_1617,N_1534,N_1558);
nor U1618 (N_1618,N_1532,N_1567);
nand U1619 (N_1619,N_1527,N_1574);
nand U1620 (N_1620,N_1515,N_1501);
nor U1621 (N_1621,N_1502,N_1513);
and U1622 (N_1622,N_1543,N_1509);
xor U1623 (N_1623,N_1500,N_1574);
nand U1624 (N_1624,N_1534,N_1567);
nand U1625 (N_1625,N_1564,N_1512);
nor U1626 (N_1626,N_1511,N_1539);
or U1627 (N_1627,N_1546,N_1555);
or U1628 (N_1628,N_1533,N_1546);
and U1629 (N_1629,N_1529,N_1509);
or U1630 (N_1630,N_1541,N_1560);
and U1631 (N_1631,N_1564,N_1538);
and U1632 (N_1632,N_1543,N_1538);
nor U1633 (N_1633,N_1525,N_1526);
and U1634 (N_1634,N_1559,N_1569);
nand U1635 (N_1635,N_1538,N_1568);
nand U1636 (N_1636,N_1507,N_1523);
or U1637 (N_1637,N_1545,N_1508);
nand U1638 (N_1638,N_1552,N_1531);
or U1639 (N_1639,N_1519,N_1542);
or U1640 (N_1640,N_1501,N_1530);
and U1641 (N_1641,N_1525,N_1539);
nand U1642 (N_1642,N_1539,N_1548);
nand U1643 (N_1643,N_1542,N_1500);
nor U1644 (N_1644,N_1523,N_1561);
nand U1645 (N_1645,N_1505,N_1571);
nand U1646 (N_1646,N_1555,N_1551);
nor U1647 (N_1647,N_1544,N_1560);
nand U1648 (N_1648,N_1500,N_1546);
or U1649 (N_1649,N_1548,N_1535);
nor U1650 (N_1650,N_1588,N_1613);
and U1651 (N_1651,N_1627,N_1620);
nor U1652 (N_1652,N_1575,N_1605);
nand U1653 (N_1653,N_1609,N_1630);
and U1654 (N_1654,N_1643,N_1612);
or U1655 (N_1655,N_1632,N_1600);
nand U1656 (N_1656,N_1611,N_1594);
or U1657 (N_1657,N_1598,N_1642);
and U1658 (N_1658,N_1602,N_1631);
nand U1659 (N_1659,N_1629,N_1633);
nand U1660 (N_1660,N_1649,N_1582);
nor U1661 (N_1661,N_1604,N_1621);
nand U1662 (N_1662,N_1576,N_1635);
nand U1663 (N_1663,N_1597,N_1590);
and U1664 (N_1664,N_1614,N_1638);
and U1665 (N_1665,N_1585,N_1636);
nand U1666 (N_1666,N_1644,N_1639);
nand U1667 (N_1667,N_1599,N_1616);
and U1668 (N_1668,N_1610,N_1592);
nor U1669 (N_1669,N_1618,N_1584);
or U1670 (N_1670,N_1617,N_1628);
and U1671 (N_1671,N_1577,N_1647);
nand U1672 (N_1672,N_1645,N_1586);
or U1673 (N_1673,N_1596,N_1640);
or U1674 (N_1674,N_1648,N_1591);
and U1675 (N_1675,N_1581,N_1637);
nor U1676 (N_1676,N_1641,N_1595);
or U1677 (N_1677,N_1603,N_1593);
and U1678 (N_1678,N_1578,N_1619);
nand U1679 (N_1679,N_1601,N_1579);
nor U1680 (N_1680,N_1587,N_1623);
nor U1681 (N_1681,N_1626,N_1622);
or U1682 (N_1682,N_1583,N_1646);
nor U1683 (N_1683,N_1615,N_1580);
nand U1684 (N_1684,N_1624,N_1606);
and U1685 (N_1685,N_1634,N_1589);
nand U1686 (N_1686,N_1608,N_1607);
and U1687 (N_1687,N_1625,N_1599);
or U1688 (N_1688,N_1582,N_1591);
and U1689 (N_1689,N_1635,N_1606);
or U1690 (N_1690,N_1637,N_1622);
or U1691 (N_1691,N_1606,N_1600);
and U1692 (N_1692,N_1607,N_1643);
nor U1693 (N_1693,N_1592,N_1622);
nor U1694 (N_1694,N_1644,N_1624);
and U1695 (N_1695,N_1619,N_1595);
nand U1696 (N_1696,N_1577,N_1643);
nor U1697 (N_1697,N_1580,N_1620);
nand U1698 (N_1698,N_1616,N_1604);
or U1699 (N_1699,N_1584,N_1644);
nand U1700 (N_1700,N_1646,N_1617);
or U1701 (N_1701,N_1586,N_1632);
and U1702 (N_1702,N_1626,N_1649);
nor U1703 (N_1703,N_1634,N_1613);
nor U1704 (N_1704,N_1639,N_1649);
or U1705 (N_1705,N_1620,N_1606);
and U1706 (N_1706,N_1611,N_1618);
nand U1707 (N_1707,N_1637,N_1607);
nand U1708 (N_1708,N_1591,N_1633);
nand U1709 (N_1709,N_1575,N_1611);
nor U1710 (N_1710,N_1634,N_1640);
nor U1711 (N_1711,N_1615,N_1607);
nor U1712 (N_1712,N_1617,N_1586);
or U1713 (N_1713,N_1619,N_1602);
or U1714 (N_1714,N_1623,N_1639);
or U1715 (N_1715,N_1642,N_1605);
and U1716 (N_1716,N_1616,N_1612);
or U1717 (N_1717,N_1632,N_1580);
or U1718 (N_1718,N_1630,N_1633);
nand U1719 (N_1719,N_1577,N_1623);
nor U1720 (N_1720,N_1601,N_1619);
or U1721 (N_1721,N_1624,N_1638);
or U1722 (N_1722,N_1603,N_1630);
or U1723 (N_1723,N_1628,N_1580);
nand U1724 (N_1724,N_1605,N_1625);
nor U1725 (N_1725,N_1690,N_1651);
or U1726 (N_1726,N_1684,N_1658);
or U1727 (N_1727,N_1657,N_1712);
or U1728 (N_1728,N_1694,N_1673);
nor U1729 (N_1729,N_1675,N_1655);
or U1730 (N_1730,N_1715,N_1706);
nand U1731 (N_1731,N_1654,N_1671);
or U1732 (N_1732,N_1722,N_1699);
and U1733 (N_1733,N_1714,N_1719);
nor U1734 (N_1734,N_1674,N_1701);
or U1735 (N_1735,N_1660,N_1666);
or U1736 (N_1736,N_1704,N_1689);
or U1737 (N_1737,N_1662,N_1724);
nand U1738 (N_1738,N_1672,N_1656);
nand U1739 (N_1739,N_1667,N_1650);
nand U1740 (N_1740,N_1696,N_1702);
nor U1741 (N_1741,N_1720,N_1653);
nor U1742 (N_1742,N_1669,N_1652);
or U1743 (N_1743,N_1686,N_1718);
and U1744 (N_1744,N_1677,N_1707);
nor U1745 (N_1745,N_1691,N_1692);
nand U1746 (N_1746,N_1668,N_1709);
xnor U1747 (N_1747,N_1700,N_1661);
or U1748 (N_1748,N_1711,N_1708);
nor U1749 (N_1749,N_1679,N_1678);
nor U1750 (N_1750,N_1665,N_1695);
nor U1751 (N_1751,N_1683,N_1705);
nand U1752 (N_1752,N_1716,N_1680);
and U1753 (N_1753,N_1670,N_1681);
nand U1754 (N_1754,N_1703,N_1698);
and U1755 (N_1755,N_1676,N_1697);
or U1756 (N_1756,N_1710,N_1685);
and U1757 (N_1757,N_1688,N_1717);
nor U1758 (N_1758,N_1687,N_1721);
or U1759 (N_1759,N_1664,N_1663);
xnor U1760 (N_1760,N_1682,N_1723);
and U1761 (N_1761,N_1713,N_1693);
nor U1762 (N_1762,N_1659,N_1672);
nor U1763 (N_1763,N_1685,N_1708);
nor U1764 (N_1764,N_1678,N_1708);
and U1765 (N_1765,N_1713,N_1690);
nand U1766 (N_1766,N_1705,N_1716);
and U1767 (N_1767,N_1658,N_1690);
nand U1768 (N_1768,N_1653,N_1682);
or U1769 (N_1769,N_1680,N_1695);
nand U1770 (N_1770,N_1665,N_1651);
or U1771 (N_1771,N_1699,N_1654);
nor U1772 (N_1772,N_1666,N_1655);
nand U1773 (N_1773,N_1676,N_1653);
or U1774 (N_1774,N_1709,N_1673);
nor U1775 (N_1775,N_1723,N_1659);
nor U1776 (N_1776,N_1697,N_1711);
or U1777 (N_1777,N_1682,N_1669);
nor U1778 (N_1778,N_1662,N_1652);
or U1779 (N_1779,N_1682,N_1709);
or U1780 (N_1780,N_1656,N_1651);
or U1781 (N_1781,N_1676,N_1686);
and U1782 (N_1782,N_1680,N_1683);
nor U1783 (N_1783,N_1693,N_1720);
or U1784 (N_1784,N_1665,N_1694);
and U1785 (N_1785,N_1721,N_1655);
or U1786 (N_1786,N_1716,N_1660);
nand U1787 (N_1787,N_1723,N_1708);
nand U1788 (N_1788,N_1652,N_1681);
and U1789 (N_1789,N_1660,N_1703);
nor U1790 (N_1790,N_1703,N_1677);
xor U1791 (N_1791,N_1677,N_1685);
nand U1792 (N_1792,N_1721,N_1682);
and U1793 (N_1793,N_1652,N_1674);
nor U1794 (N_1794,N_1655,N_1684);
nand U1795 (N_1795,N_1703,N_1659);
nand U1796 (N_1796,N_1683,N_1691);
nand U1797 (N_1797,N_1716,N_1653);
or U1798 (N_1798,N_1668,N_1671);
and U1799 (N_1799,N_1696,N_1664);
nand U1800 (N_1800,N_1731,N_1764);
nor U1801 (N_1801,N_1770,N_1741);
nor U1802 (N_1802,N_1777,N_1747);
nand U1803 (N_1803,N_1772,N_1771);
nor U1804 (N_1804,N_1760,N_1759);
or U1805 (N_1805,N_1796,N_1748);
and U1806 (N_1806,N_1785,N_1756);
or U1807 (N_1807,N_1793,N_1749);
and U1808 (N_1808,N_1790,N_1744);
and U1809 (N_1809,N_1799,N_1752);
or U1810 (N_1810,N_1735,N_1730);
or U1811 (N_1811,N_1774,N_1757);
nor U1812 (N_1812,N_1746,N_1789);
nand U1813 (N_1813,N_1732,N_1734);
nand U1814 (N_1814,N_1778,N_1728);
nor U1815 (N_1815,N_1750,N_1762);
and U1816 (N_1816,N_1780,N_1782);
and U1817 (N_1817,N_1792,N_1797);
nand U1818 (N_1818,N_1769,N_1738);
nand U1819 (N_1819,N_1776,N_1733);
nand U1820 (N_1820,N_1751,N_1740);
or U1821 (N_1821,N_1794,N_1737);
or U1822 (N_1822,N_1798,N_1726);
and U1823 (N_1823,N_1739,N_1781);
nor U1824 (N_1824,N_1761,N_1783);
and U1825 (N_1825,N_1729,N_1725);
nand U1826 (N_1826,N_1787,N_1745);
or U1827 (N_1827,N_1791,N_1775);
nor U1828 (N_1828,N_1767,N_1773);
nor U1829 (N_1829,N_1736,N_1753);
nand U1830 (N_1830,N_1784,N_1755);
nor U1831 (N_1831,N_1768,N_1765);
or U1832 (N_1832,N_1779,N_1788);
and U1833 (N_1833,N_1727,N_1763);
nand U1834 (N_1834,N_1758,N_1795);
nor U1835 (N_1835,N_1743,N_1766);
or U1836 (N_1836,N_1786,N_1742);
and U1837 (N_1837,N_1754,N_1782);
and U1838 (N_1838,N_1750,N_1741);
or U1839 (N_1839,N_1738,N_1735);
or U1840 (N_1840,N_1787,N_1744);
and U1841 (N_1841,N_1746,N_1750);
nand U1842 (N_1842,N_1760,N_1790);
nor U1843 (N_1843,N_1780,N_1776);
nor U1844 (N_1844,N_1766,N_1763);
nand U1845 (N_1845,N_1771,N_1738);
and U1846 (N_1846,N_1749,N_1768);
nor U1847 (N_1847,N_1757,N_1738);
and U1848 (N_1848,N_1765,N_1747);
nand U1849 (N_1849,N_1783,N_1742);
or U1850 (N_1850,N_1735,N_1765);
nor U1851 (N_1851,N_1799,N_1769);
nand U1852 (N_1852,N_1780,N_1781);
nor U1853 (N_1853,N_1746,N_1795);
nor U1854 (N_1854,N_1794,N_1744);
nor U1855 (N_1855,N_1789,N_1745);
or U1856 (N_1856,N_1752,N_1784);
nand U1857 (N_1857,N_1773,N_1729);
nand U1858 (N_1858,N_1770,N_1783);
and U1859 (N_1859,N_1779,N_1738);
or U1860 (N_1860,N_1763,N_1797);
nand U1861 (N_1861,N_1728,N_1754);
or U1862 (N_1862,N_1773,N_1778);
nor U1863 (N_1863,N_1762,N_1749);
nor U1864 (N_1864,N_1757,N_1765);
or U1865 (N_1865,N_1730,N_1774);
and U1866 (N_1866,N_1728,N_1759);
nor U1867 (N_1867,N_1732,N_1791);
and U1868 (N_1868,N_1745,N_1749);
nor U1869 (N_1869,N_1765,N_1789);
and U1870 (N_1870,N_1737,N_1781);
nor U1871 (N_1871,N_1767,N_1766);
and U1872 (N_1872,N_1760,N_1775);
or U1873 (N_1873,N_1793,N_1754);
nand U1874 (N_1874,N_1794,N_1799);
or U1875 (N_1875,N_1808,N_1835);
nand U1876 (N_1876,N_1847,N_1852);
nand U1877 (N_1877,N_1804,N_1817);
nor U1878 (N_1878,N_1857,N_1824);
and U1879 (N_1879,N_1805,N_1801);
nand U1880 (N_1880,N_1820,N_1812);
nand U1881 (N_1881,N_1838,N_1822);
nor U1882 (N_1882,N_1811,N_1819);
nand U1883 (N_1883,N_1871,N_1874);
nand U1884 (N_1884,N_1843,N_1806);
and U1885 (N_1885,N_1829,N_1826);
nor U1886 (N_1886,N_1807,N_1859);
nor U1887 (N_1887,N_1810,N_1803);
and U1888 (N_1888,N_1814,N_1813);
nand U1889 (N_1889,N_1872,N_1863);
nand U1890 (N_1890,N_1821,N_1869);
or U1891 (N_1891,N_1825,N_1828);
nand U1892 (N_1892,N_1860,N_1845);
nand U1893 (N_1893,N_1839,N_1830);
nor U1894 (N_1894,N_1816,N_1866);
or U1895 (N_1895,N_1864,N_1834);
xor U1896 (N_1896,N_1873,N_1846);
nor U1897 (N_1897,N_1823,N_1865);
nand U1898 (N_1898,N_1868,N_1870);
nor U1899 (N_1899,N_1851,N_1853);
or U1900 (N_1900,N_1809,N_1837);
or U1901 (N_1901,N_1831,N_1827);
or U1902 (N_1902,N_1842,N_1818);
nor U1903 (N_1903,N_1850,N_1844);
nor U1904 (N_1904,N_1836,N_1855);
nand U1905 (N_1905,N_1858,N_1862);
and U1906 (N_1906,N_1856,N_1802);
nor U1907 (N_1907,N_1861,N_1849);
nand U1908 (N_1908,N_1800,N_1841);
nor U1909 (N_1909,N_1854,N_1840);
nand U1910 (N_1910,N_1832,N_1867);
nor U1911 (N_1911,N_1833,N_1848);
nor U1912 (N_1912,N_1815,N_1802);
nor U1913 (N_1913,N_1854,N_1869);
nor U1914 (N_1914,N_1811,N_1826);
or U1915 (N_1915,N_1864,N_1832);
nor U1916 (N_1916,N_1833,N_1825);
and U1917 (N_1917,N_1827,N_1866);
nand U1918 (N_1918,N_1839,N_1816);
and U1919 (N_1919,N_1846,N_1867);
nor U1920 (N_1920,N_1851,N_1874);
or U1921 (N_1921,N_1844,N_1857);
nor U1922 (N_1922,N_1837,N_1844);
nand U1923 (N_1923,N_1805,N_1869);
or U1924 (N_1924,N_1847,N_1864);
nor U1925 (N_1925,N_1848,N_1811);
nand U1926 (N_1926,N_1813,N_1825);
or U1927 (N_1927,N_1804,N_1864);
nor U1928 (N_1928,N_1830,N_1863);
and U1929 (N_1929,N_1843,N_1857);
nand U1930 (N_1930,N_1811,N_1808);
and U1931 (N_1931,N_1821,N_1839);
nor U1932 (N_1932,N_1833,N_1859);
or U1933 (N_1933,N_1829,N_1864);
nand U1934 (N_1934,N_1854,N_1829);
and U1935 (N_1935,N_1850,N_1846);
nor U1936 (N_1936,N_1823,N_1858);
xor U1937 (N_1937,N_1811,N_1844);
or U1938 (N_1938,N_1831,N_1811);
and U1939 (N_1939,N_1860,N_1838);
or U1940 (N_1940,N_1804,N_1827);
nor U1941 (N_1941,N_1844,N_1863);
or U1942 (N_1942,N_1869,N_1853);
nor U1943 (N_1943,N_1806,N_1865);
nand U1944 (N_1944,N_1810,N_1841);
and U1945 (N_1945,N_1816,N_1801);
nand U1946 (N_1946,N_1869,N_1825);
and U1947 (N_1947,N_1825,N_1871);
or U1948 (N_1948,N_1858,N_1863);
nor U1949 (N_1949,N_1817,N_1829);
nand U1950 (N_1950,N_1902,N_1942);
nand U1951 (N_1951,N_1877,N_1901);
nand U1952 (N_1952,N_1932,N_1912);
nor U1953 (N_1953,N_1913,N_1937);
nor U1954 (N_1954,N_1888,N_1904);
or U1955 (N_1955,N_1949,N_1924);
or U1956 (N_1956,N_1929,N_1897);
and U1957 (N_1957,N_1923,N_1945);
and U1958 (N_1958,N_1914,N_1930);
nand U1959 (N_1959,N_1893,N_1946);
or U1960 (N_1960,N_1905,N_1938);
and U1961 (N_1961,N_1896,N_1907);
or U1962 (N_1962,N_1934,N_1879);
or U1963 (N_1963,N_1925,N_1889);
nor U1964 (N_1964,N_1891,N_1918);
nor U1965 (N_1965,N_1895,N_1920);
nor U1966 (N_1966,N_1875,N_1933);
nand U1967 (N_1967,N_1947,N_1927);
nand U1968 (N_1968,N_1926,N_1899);
nand U1969 (N_1969,N_1935,N_1919);
nor U1970 (N_1970,N_1892,N_1885);
nand U1971 (N_1971,N_1936,N_1883);
or U1972 (N_1972,N_1887,N_1906);
and U1973 (N_1973,N_1910,N_1948);
nor U1974 (N_1974,N_1915,N_1908);
and U1975 (N_1975,N_1911,N_1909);
or U1976 (N_1976,N_1890,N_1900);
nor U1977 (N_1977,N_1881,N_1944);
or U1978 (N_1978,N_1880,N_1941);
nand U1979 (N_1979,N_1922,N_1939);
and U1980 (N_1980,N_1940,N_1894);
xor U1981 (N_1981,N_1876,N_1878);
nand U1982 (N_1982,N_1917,N_1884);
and U1983 (N_1983,N_1882,N_1916);
or U1984 (N_1984,N_1886,N_1928);
nand U1985 (N_1985,N_1898,N_1943);
or U1986 (N_1986,N_1921,N_1931);
and U1987 (N_1987,N_1903,N_1929);
and U1988 (N_1988,N_1908,N_1875);
nand U1989 (N_1989,N_1875,N_1911);
or U1990 (N_1990,N_1919,N_1934);
and U1991 (N_1991,N_1925,N_1883);
and U1992 (N_1992,N_1928,N_1923);
and U1993 (N_1993,N_1907,N_1908);
or U1994 (N_1994,N_1894,N_1918);
and U1995 (N_1995,N_1923,N_1888);
nand U1996 (N_1996,N_1912,N_1911);
or U1997 (N_1997,N_1896,N_1884);
nand U1998 (N_1998,N_1945,N_1906);
or U1999 (N_1999,N_1931,N_1932);
and U2000 (N_2000,N_1924,N_1930);
and U2001 (N_2001,N_1887,N_1926);
nand U2002 (N_2002,N_1927,N_1928);
or U2003 (N_2003,N_1897,N_1940);
or U2004 (N_2004,N_1926,N_1943);
or U2005 (N_2005,N_1930,N_1906);
and U2006 (N_2006,N_1906,N_1933);
nand U2007 (N_2007,N_1914,N_1899);
and U2008 (N_2008,N_1943,N_1935);
nor U2009 (N_2009,N_1883,N_1879);
nand U2010 (N_2010,N_1912,N_1945);
or U2011 (N_2011,N_1907,N_1937);
and U2012 (N_2012,N_1910,N_1914);
nor U2013 (N_2013,N_1946,N_1943);
nand U2014 (N_2014,N_1928,N_1899);
and U2015 (N_2015,N_1943,N_1945);
and U2016 (N_2016,N_1883,N_1908);
or U2017 (N_2017,N_1945,N_1936);
and U2018 (N_2018,N_1931,N_1923);
or U2019 (N_2019,N_1902,N_1944);
nand U2020 (N_2020,N_1917,N_1913);
nor U2021 (N_2021,N_1902,N_1907);
nand U2022 (N_2022,N_1920,N_1947);
nand U2023 (N_2023,N_1936,N_1899);
nor U2024 (N_2024,N_1942,N_1896);
nand U2025 (N_2025,N_2012,N_2003);
or U2026 (N_2026,N_1972,N_1971);
nor U2027 (N_2027,N_1964,N_1958);
nor U2028 (N_2028,N_1996,N_1957);
or U2029 (N_2029,N_1967,N_1986);
and U2030 (N_2030,N_1960,N_1985);
and U2031 (N_2031,N_1981,N_2011);
nor U2032 (N_2032,N_1962,N_2024);
or U2033 (N_2033,N_1983,N_2018);
nor U2034 (N_2034,N_1982,N_2016);
nor U2035 (N_2035,N_1963,N_1979);
or U2036 (N_2036,N_1955,N_2013);
or U2037 (N_2037,N_1970,N_1966);
or U2038 (N_2038,N_2021,N_1961);
and U2039 (N_2039,N_1973,N_1976);
or U2040 (N_2040,N_2019,N_1974);
nor U2041 (N_2041,N_1995,N_1956);
nand U2042 (N_2042,N_1965,N_1988);
nand U2043 (N_2043,N_2000,N_2020);
or U2044 (N_2044,N_2010,N_1950);
nand U2045 (N_2045,N_1953,N_1994);
and U2046 (N_2046,N_1989,N_1969);
and U2047 (N_2047,N_2009,N_1997);
xor U2048 (N_2048,N_1987,N_1954);
or U2049 (N_2049,N_1951,N_1952);
nand U2050 (N_2050,N_2005,N_2017);
and U2051 (N_2051,N_1991,N_1992);
or U2052 (N_2052,N_2008,N_2015);
and U2053 (N_2053,N_1999,N_2022);
nor U2054 (N_2054,N_2001,N_1977);
nand U2055 (N_2055,N_1975,N_1980);
nand U2056 (N_2056,N_2004,N_1984);
nor U2057 (N_2057,N_2023,N_2002);
or U2058 (N_2058,N_2007,N_1993);
and U2059 (N_2059,N_2014,N_1990);
nor U2060 (N_2060,N_1998,N_1978);
and U2061 (N_2061,N_1968,N_2006);
or U2062 (N_2062,N_1959,N_1953);
and U2063 (N_2063,N_2005,N_2010);
nor U2064 (N_2064,N_2017,N_1993);
nand U2065 (N_2065,N_1997,N_2001);
and U2066 (N_2066,N_2000,N_2022);
nand U2067 (N_2067,N_1977,N_1972);
nand U2068 (N_2068,N_1990,N_2002);
nand U2069 (N_2069,N_1971,N_1950);
xor U2070 (N_2070,N_1962,N_1995);
and U2071 (N_2071,N_2005,N_1996);
and U2072 (N_2072,N_1973,N_1985);
nor U2073 (N_2073,N_1979,N_2023);
or U2074 (N_2074,N_1961,N_1974);
and U2075 (N_2075,N_1992,N_1960);
nor U2076 (N_2076,N_1981,N_1953);
and U2077 (N_2077,N_2014,N_2003);
nor U2078 (N_2078,N_1965,N_2012);
nor U2079 (N_2079,N_1952,N_2016);
and U2080 (N_2080,N_1950,N_1974);
nand U2081 (N_2081,N_1956,N_1976);
nand U2082 (N_2082,N_2003,N_1978);
or U2083 (N_2083,N_1979,N_2004);
and U2084 (N_2084,N_2009,N_2023);
and U2085 (N_2085,N_1985,N_1993);
or U2086 (N_2086,N_2014,N_2016);
nand U2087 (N_2087,N_1970,N_1950);
nor U2088 (N_2088,N_2017,N_2001);
nor U2089 (N_2089,N_1989,N_1987);
and U2090 (N_2090,N_2021,N_1979);
and U2091 (N_2091,N_1999,N_1951);
nand U2092 (N_2092,N_2017,N_1968);
nor U2093 (N_2093,N_1959,N_2006);
and U2094 (N_2094,N_1976,N_1990);
nand U2095 (N_2095,N_2024,N_1996);
nor U2096 (N_2096,N_1952,N_1999);
nor U2097 (N_2097,N_1961,N_1979);
nand U2098 (N_2098,N_1962,N_1950);
nor U2099 (N_2099,N_1970,N_1998);
nand U2100 (N_2100,N_2048,N_2075);
and U2101 (N_2101,N_2032,N_2027);
and U2102 (N_2102,N_2066,N_2097);
or U2103 (N_2103,N_2089,N_2096);
nand U2104 (N_2104,N_2069,N_2088);
and U2105 (N_2105,N_2033,N_2039);
or U2106 (N_2106,N_2070,N_2040);
nor U2107 (N_2107,N_2030,N_2068);
nor U2108 (N_2108,N_2093,N_2056);
nor U2109 (N_2109,N_2079,N_2092);
or U2110 (N_2110,N_2094,N_2065);
and U2111 (N_2111,N_2041,N_2051);
and U2112 (N_2112,N_2043,N_2080);
nand U2113 (N_2113,N_2083,N_2058);
nor U2114 (N_2114,N_2081,N_2029);
and U2115 (N_2115,N_2091,N_2098);
nor U2116 (N_2116,N_2074,N_2082);
nor U2117 (N_2117,N_2047,N_2077);
nand U2118 (N_2118,N_2076,N_2078);
nor U2119 (N_2119,N_2073,N_2060);
or U2120 (N_2120,N_2099,N_2045);
nor U2121 (N_2121,N_2046,N_2050);
and U2122 (N_2122,N_2071,N_2067);
xnor U2123 (N_2123,N_2038,N_2034);
or U2124 (N_2124,N_2052,N_2044);
or U2125 (N_2125,N_2084,N_2061);
or U2126 (N_2126,N_2055,N_2035);
and U2127 (N_2127,N_2095,N_2053);
nand U2128 (N_2128,N_2085,N_2054);
nor U2129 (N_2129,N_2031,N_2042);
nor U2130 (N_2130,N_2062,N_2026);
or U2131 (N_2131,N_2028,N_2057);
and U2132 (N_2132,N_2059,N_2087);
and U2133 (N_2133,N_2072,N_2064);
or U2134 (N_2134,N_2036,N_2049);
nor U2135 (N_2135,N_2090,N_2086);
nand U2136 (N_2136,N_2037,N_2025);
or U2137 (N_2137,N_2063,N_2042);
or U2138 (N_2138,N_2092,N_2051);
or U2139 (N_2139,N_2034,N_2096);
or U2140 (N_2140,N_2096,N_2079);
nand U2141 (N_2141,N_2055,N_2058);
or U2142 (N_2142,N_2070,N_2076);
and U2143 (N_2143,N_2080,N_2068);
nor U2144 (N_2144,N_2063,N_2043);
nand U2145 (N_2145,N_2033,N_2086);
nand U2146 (N_2146,N_2062,N_2092);
nand U2147 (N_2147,N_2054,N_2060);
nand U2148 (N_2148,N_2059,N_2085);
or U2149 (N_2149,N_2028,N_2036);
and U2150 (N_2150,N_2058,N_2085);
nor U2151 (N_2151,N_2080,N_2074);
nor U2152 (N_2152,N_2084,N_2080);
xor U2153 (N_2153,N_2094,N_2073);
and U2154 (N_2154,N_2081,N_2064);
and U2155 (N_2155,N_2094,N_2096);
nand U2156 (N_2156,N_2030,N_2083);
nor U2157 (N_2157,N_2090,N_2052);
and U2158 (N_2158,N_2077,N_2054);
and U2159 (N_2159,N_2034,N_2069);
and U2160 (N_2160,N_2072,N_2037);
or U2161 (N_2161,N_2073,N_2091);
and U2162 (N_2162,N_2088,N_2040);
nor U2163 (N_2163,N_2072,N_2044);
nand U2164 (N_2164,N_2053,N_2049);
and U2165 (N_2165,N_2070,N_2059);
or U2166 (N_2166,N_2042,N_2082);
nor U2167 (N_2167,N_2034,N_2071);
or U2168 (N_2168,N_2041,N_2059);
nand U2169 (N_2169,N_2041,N_2083);
nor U2170 (N_2170,N_2088,N_2083);
or U2171 (N_2171,N_2080,N_2078);
nor U2172 (N_2172,N_2061,N_2039);
nand U2173 (N_2173,N_2077,N_2051);
nor U2174 (N_2174,N_2041,N_2055);
nand U2175 (N_2175,N_2159,N_2167);
nand U2176 (N_2176,N_2151,N_2120);
nand U2177 (N_2177,N_2155,N_2135);
and U2178 (N_2178,N_2140,N_2145);
and U2179 (N_2179,N_2141,N_2109);
and U2180 (N_2180,N_2152,N_2146);
nand U2181 (N_2181,N_2100,N_2129);
or U2182 (N_2182,N_2110,N_2128);
nand U2183 (N_2183,N_2136,N_2126);
and U2184 (N_2184,N_2101,N_2142);
or U2185 (N_2185,N_2137,N_2154);
and U2186 (N_2186,N_2158,N_2130);
nand U2187 (N_2187,N_2122,N_2153);
nand U2188 (N_2188,N_2166,N_2127);
nor U2189 (N_2189,N_2156,N_2132);
and U2190 (N_2190,N_2115,N_2118);
nor U2191 (N_2191,N_2113,N_2134);
nand U2192 (N_2192,N_2147,N_2104);
or U2193 (N_2193,N_2131,N_2139);
nor U2194 (N_2194,N_2168,N_2174);
nand U2195 (N_2195,N_2163,N_2102);
nand U2196 (N_2196,N_2138,N_2172);
nand U2197 (N_2197,N_2112,N_2123);
nor U2198 (N_2198,N_2161,N_2111);
nor U2199 (N_2199,N_2125,N_2133);
nand U2200 (N_2200,N_2169,N_2157);
nand U2201 (N_2201,N_2162,N_2114);
nand U2202 (N_2202,N_2116,N_2165);
or U2203 (N_2203,N_2160,N_2124);
or U2204 (N_2204,N_2117,N_2121);
or U2205 (N_2205,N_2170,N_2106);
and U2206 (N_2206,N_2144,N_2143);
or U2207 (N_2207,N_2150,N_2103);
or U2208 (N_2208,N_2105,N_2107);
and U2209 (N_2209,N_2164,N_2149);
or U2210 (N_2210,N_2108,N_2148);
nand U2211 (N_2211,N_2173,N_2119);
or U2212 (N_2212,N_2171,N_2142);
and U2213 (N_2213,N_2173,N_2103);
nor U2214 (N_2214,N_2119,N_2146);
nand U2215 (N_2215,N_2156,N_2126);
nand U2216 (N_2216,N_2131,N_2129);
nor U2217 (N_2217,N_2114,N_2128);
nand U2218 (N_2218,N_2164,N_2150);
nand U2219 (N_2219,N_2161,N_2141);
nand U2220 (N_2220,N_2173,N_2115);
nand U2221 (N_2221,N_2124,N_2112);
nand U2222 (N_2222,N_2111,N_2172);
or U2223 (N_2223,N_2167,N_2155);
and U2224 (N_2224,N_2138,N_2152);
nor U2225 (N_2225,N_2160,N_2167);
nor U2226 (N_2226,N_2170,N_2119);
or U2227 (N_2227,N_2154,N_2103);
nor U2228 (N_2228,N_2159,N_2129);
or U2229 (N_2229,N_2162,N_2124);
nand U2230 (N_2230,N_2115,N_2120);
nand U2231 (N_2231,N_2112,N_2113);
or U2232 (N_2232,N_2169,N_2173);
xnor U2233 (N_2233,N_2160,N_2122);
or U2234 (N_2234,N_2111,N_2104);
nand U2235 (N_2235,N_2153,N_2109);
nand U2236 (N_2236,N_2114,N_2119);
nor U2237 (N_2237,N_2127,N_2105);
and U2238 (N_2238,N_2137,N_2145);
nor U2239 (N_2239,N_2169,N_2127);
and U2240 (N_2240,N_2114,N_2137);
nand U2241 (N_2241,N_2169,N_2103);
and U2242 (N_2242,N_2147,N_2169);
and U2243 (N_2243,N_2149,N_2131);
nand U2244 (N_2244,N_2136,N_2119);
xnor U2245 (N_2245,N_2112,N_2147);
and U2246 (N_2246,N_2170,N_2144);
nand U2247 (N_2247,N_2145,N_2151);
nor U2248 (N_2248,N_2171,N_2152);
nor U2249 (N_2249,N_2114,N_2147);
and U2250 (N_2250,N_2242,N_2189);
or U2251 (N_2251,N_2236,N_2245);
or U2252 (N_2252,N_2232,N_2199);
or U2253 (N_2253,N_2208,N_2187);
nor U2254 (N_2254,N_2179,N_2175);
or U2255 (N_2255,N_2231,N_2177);
nor U2256 (N_2256,N_2198,N_2209);
or U2257 (N_2257,N_2244,N_2203);
nand U2258 (N_2258,N_2190,N_2184);
or U2259 (N_2259,N_2228,N_2246);
or U2260 (N_2260,N_2235,N_2249);
nor U2261 (N_2261,N_2201,N_2219);
nand U2262 (N_2262,N_2225,N_2216);
nor U2263 (N_2263,N_2191,N_2196);
nor U2264 (N_2264,N_2218,N_2197);
nor U2265 (N_2265,N_2217,N_2188);
nor U2266 (N_2266,N_2240,N_2211);
and U2267 (N_2267,N_2210,N_2193);
nor U2268 (N_2268,N_2183,N_2215);
or U2269 (N_2269,N_2233,N_2247);
and U2270 (N_2270,N_2205,N_2234);
nand U2271 (N_2271,N_2181,N_2180);
nor U2272 (N_2272,N_2194,N_2238);
and U2273 (N_2273,N_2192,N_2248);
and U2274 (N_2274,N_2220,N_2226);
nor U2275 (N_2275,N_2237,N_2200);
nand U2276 (N_2276,N_2230,N_2241);
nor U2277 (N_2277,N_2221,N_2185);
nor U2278 (N_2278,N_2182,N_2213);
or U2279 (N_2279,N_2206,N_2176);
nand U2280 (N_2280,N_2224,N_2195);
or U2281 (N_2281,N_2178,N_2223);
or U2282 (N_2282,N_2227,N_2239);
nand U2283 (N_2283,N_2243,N_2186);
or U2284 (N_2284,N_2212,N_2204);
or U2285 (N_2285,N_2222,N_2207);
and U2286 (N_2286,N_2214,N_2229);
or U2287 (N_2287,N_2202,N_2179);
nand U2288 (N_2288,N_2239,N_2248);
nor U2289 (N_2289,N_2188,N_2203);
and U2290 (N_2290,N_2230,N_2177);
and U2291 (N_2291,N_2215,N_2240);
nand U2292 (N_2292,N_2247,N_2240);
nand U2293 (N_2293,N_2219,N_2224);
and U2294 (N_2294,N_2238,N_2190);
or U2295 (N_2295,N_2202,N_2244);
nor U2296 (N_2296,N_2199,N_2222);
or U2297 (N_2297,N_2179,N_2200);
or U2298 (N_2298,N_2198,N_2237);
or U2299 (N_2299,N_2246,N_2233);
nand U2300 (N_2300,N_2201,N_2217);
and U2301 (N_2301,N_2188,N_2185);
nand U2302 (N_2302,N_2184,N_2221);
nor U2303 (N_2303,N_2188,N_2191);
or U2304 (N_2304,N_2241,N_2216);
or U2305 (N_2305,N_2219,N_2233);
and U2306 (N_2306,N_2196,N_2215);
and U2307 (N_2307,N_2239,N_2187);
nand U2308 (N_2308,N_2189,N_2246);
nand U2309 (N_2309,N_2227,N_2187);
xnor U2310 (N_2310,N_2175,N_2185);
and U2311 (N_2311,N_2179,N_2228);
nor U2312 (N_2312,N_2220,N_2216);
nor U2313 (N_2313,N_2176,N_2177);
or U2314 (N_2314,N_2191,N_2195);
or U2315 (N_2315,N_2215,N_2245);
and U2316 (N_2316,N_2246,N_2195);
nand U2317 (N_2317,N_2223,N_2177);
nand U2318 (N_2318,N_2192,N_2175);
nor U2319 (N_2319,N_2244,N_2180);
and U2320 (N_2320,N_2208,N_2182);
and U2321 (N_2321,N_2190,N_2246);
nor U2322 (N_2322,N_2197,N_2219);
and U2323 (N_2323,N_2245,N_2235);
or U2324 (N_2324,N_2246,N_2232);
and U2325 (N_2325,N_2269,N_2280);
nor U2326 (N_2326,N_2291,N_2321);
nor U2327 (N_2327,N_2288,N_2273);
nand U2328 (N_2328,N_2252,N_2299);
and U2329 (N_2329,N_2251,N_2260);
nand U2330 (N_2330,N_2312,N_2315);
nor U2331 (N_2331,N_2305,N_2284);
nor U2332 (N_2332,N_2270,N_2254);
or U2333 (N_2333,N_2303,N_2268);
nor U2334 (N_2334,N_2263,N_2316);
nand U2335 (N_2335,N_2256,N_2253);
nor U2336 (N_2336,N_2287,N_2293);
or U2337 (N_2337,N_2322,N_2301);
and U2338 (N_2338,N_2313,N_2286);
nor U2339 (N_2339,N_2314,N_2283);
or U2340 (N_2340,N_2261,N_2289);
or U2341 (N_2341,N_2308,N_2309);
or U2342 (N_2342,N_2274,N_2304);
nand U2343 (N_2343,N_2324,N_2276);
nand U2344 (N_2344,N_2265,N_2294);
nand U2345 (N_2345,N_2282,N_2317);
nand U2346 (N_2346,N_2311,N_2266);
nor U2347 (N_2347,N_2300,N_2278);
nor U2348 (N_2348,N_2275,N_2306);
nand U2349 (N_2349,N_2277,N_2267);
nand U2350 (N_2350,N_2297,N_2298);
nand U2351 (N_2351,N_2292,N_2271);
and U2352 (N_2352,N_2250,N_2259);
nand U2353 (N_2353,N_2285,N_2323);
and U2354 (N_2354,N_2318,N_2320);
and U2355 (N_2355,N_2302,N_2258);
or U2356 (N_2356,N_2257,N_2255);
and U2357 (N_2357,N_2281,N_2262);
and U2358 (N_2358,N_2290,N_2279);
and U2359 (N_2359,N_2307,N_2264);
nand U2360 (N_2360,N_2319,N_2310);
nor U2361 (N_2361,N_2296,N_2295);
or U2362 (N_2362,N_2272,N_2284);
nand U2363 (N_2363,N_2289,N_2311);
or U2364 (N_2364,N_2322,N_2289);
nor U2365 (N_2365,N_2305,N_2269);
and U2366 (N_2366,N_2275,N_2314);
or U2367 (N_2367,N_2250,N_2311);
or U2368 (N_2368,N_2293,N_2273);
or U2369 (N_2369,N_2271,N_2258);
nand U2370 (N_2370,N_2258,N_2312);
nor U2371 (N_2371,N_2261,N_2298);
and U2372 (N_2372,N_2272,N_2258);
nor U2373 (N_2373,N_2310,N_2318);
nand U2374 (N_2374,N_2270,N_2315);
nor U2375 (N_2375,N_2281,N_2321);
or U2376 (N_2376,N_2312,N_2255);
nand U2377 (N_2377,N_2308,N_2263);
and U2378 (N_2378,N_2322,N_2277);
nor U2379 (N_2379,N_2299,N_2284);
or U2380 (N_2380,N_2265,N_2303);
or U2381 (N_2381,N_2259,N_2264);
and U2382 (N_2382,N_2297,N_2271);
or U2383 (N_2383,N_2299,N_2293);
or U2384 (N_2384,N_2254,N_2298);
nor U2385 (N_2385,N_2324,N_2280);
nor U2386 (N_2386,N_2293,N_2307);
or U2387 (N_2387,N_2294,N_2256);
nor U2388 (N_2388,N_2322,N_2303);
nand U2389 (N_2389,N_2296,N_2275);
nor U2390 (N_2390,N_2256,N_2323);
and U2391 (N_2391,N_2264,N_2289);
nor U2392 (N_2392,N_2254,N_2313);
nor U2393 (N_2393,N_2267,N_2288);
nand U2394 (N_2394,N_2287,N_2315);
or U2395 (N_2395,N_2279,N_2274);
and U2396 (N_2396,N_2275,N_2265);
nor U2397 (N_2397,N_2300,N_2265);
nor U2398 (N_2398,N_2298,N_2258);
nand U2399 (N_2399,N_2279,N_2317);
nand U2400 (N_2400,N_2367,N_2356);
and U2401 (N_2401,N_2351,N_2393);
nand U2402 (N_2402,N_2363,N_2333);
or U2403 (N_2403,N_2398,N_2346);
or U2404 (N_2404,N_2382,N_2329);
and U2405 (N_2405,N_2374,N_2392);
or U2406 (N_2406,N_2335,N_2353);
nor U2407 (N_2407,N_2381,N_2368);
and U2408 (N_2408,N_2332,N_2345);
or U2409 (N_2409,N_2331,N_2348);
or U2410 (N_2410,N_2357,N_2394);
or U2411 (N_2411,N_2395,N_2330);
nand U2412 (N_2412,N_2383,N_2341);
or U2413 (N_2413,N_2339,N_2390);
and U2414 (N_2414,N_2391,N_2380);
nor U2415 (N_2415,N_2354,N_2385);
and U2416 (N_2416,N_2386,N_2397);
or U2417 (N_2417,N_2342,N_2379);
or U2418 (N_2418,N_2359,N_2334);
nand U2419 (N_2419,N_2338,N_2364);
nand U2420 (N_2420,N_2349,N_2399);
and U2421 (N_2421,N_2362,N_2389);
nand U2422 (N_2422,N_2373,N_2336);
and U2423 (N_2423,N_2344,N_2384);
nand U2424 (N_2424,N_2361,N_2388);
nor U2425 (N_2425,N_2325,N_2358);
and U2426 (N_2426,N_2387,N_2378);
nand U2427 (N_2427,N_2337,N_2396);
or U2428 (N_2428,N_2343,N_2340);
nor U2429 (N_2429,N_2352,N_2328);
nor U2430 (N_2430,N_2347,N_2377);
nor U2431 (N_2431,N_2369,N_2372);
or U2432 (N_2432,N_2366,N_2355);
or U2433 (N_2433,N_2326,N_2365);
and U2434 (N_2434,N_2376,N_2370);
nor U2435 (N_2435,N_2350,N_2375);
nand U2436 (N_2436,N_2360,N_2371);
nand U2437 (N_2437,N_2327,N_2399);
or U2438 (N_2438,N_2330,N_2365);
nor U2439 (N_2439,N_2347,N_2391);
and U2440 (N_2440,N_2339,N_2362);
or U2441 (N_2441,N_2399,N_2333);
nor U2442 (N_2442,N_2391,N_2361);
nand U2443 (N_2443,N_2370,N_2392);
and U2444 (N_2444,N_2357,N_2362);
or U2445 (N_2445,N_2394,N_2340);
and U2446 (N_2446,N_2387,N_2393);
nand U2447 (N_2447,N_2390,N_2325);
or U2448 (N_2448,N_2393,N_2359);
and U2449 (N_2449,N_2327,N_2390);
nand U2450 (N_2450,N_2390,N_2349);
and U2451 (N_2451,N_2359,N_2338);
nand U2452 (N_2452,N_2388,N_2340);
nor U2453 (N_2453,N_2354,N_2327);
nand U2454 (N_2454,N_2361,N_2390);
nand U2455 (N_2455,N_2397,N_2326);
nand U2456 (N_2456,N_2331,N_2366);
nand U2457 (N_2457,N_2365,N_2397);
or U2458 (N_2458,N_2332,N_2344);
or U2459 (N_2459,N_2385,N_2327);
nand U2460 (N_2460,N_2382,N_2367);
and U2461 (N_2461,N_2341,N_2365);
or U2462 (N_2462,N_2349,N_2328);
and U2463 (N_2463,N_2388,N_2368);
nand U2464 (N_2464,N_2349,N_2370);
nand U2465 (N_2465,N_2346,N_2339);
nand U2466 (N_2466,N_2334,N_2339);
nand U2467 (N_2467,N_2342,N_2328);
nor U2468 (N_2468,N_2337,N_2381);
and U2469 (N_2469,N_2395,N_2373);
nand U2470 (N_2470,N_2375,N_2369);
and U2471 (N_2471,N_2384,N_2349);
and U2472 (N_2472,N_2358,N_2397);
or U2473 (N_2473,N_2378,N_2344);
and U2474 (N_2474,N_2391,N_2345);
and U2475 (N_2475,N_2423,N_2452);
or U2476 (N_2476,N_2449,N_2412);
and U2477 (N_2477,N_2441,N_2400);
and U2478 (N_2478,N_2424,N_2466);
or U2479 (N_2479,N_2434,N_2431);
nand U2480 (N_2480,N_2404,N_2447);
nand U2481 (N_2481,N_2468,N_2451);
nor U2482 (N_2482,N_2469,N_2446);
or U2483 (N_2483,N_2433,N_2444);
nor U2484 (N_2484,N_2470,N_2414);
or U2485 (N_2485,N_2472,N_2471);
nand U2486 (N_2486,N_2453,N_2457);
or U2487 (N_2487,N_2459,N_2437);
nand U2488 (N_2488,N_2438,N_2429);
and U2489 (N_2489,N_2416,N_2456);
or U2490 (N_2490,N_2426,N_2409);
and U2491 (N_2491,N_2418,N_2432);
nand U2492 (N_2492,N_2443,N_2407);
or U2493 (N_2493,N_2439,N_2455);
nor U2494 (N_2494,N_2458,N_2440);
nor U2495 (N_2495,N_2419,N_2442);
and U2496 (N_2496,N_2422,N_2417);
and U2497 (N_2497,N_2460,N_2461);
nand U2498 (N_2498,N_2445,N_2420);
nand U2499 (N_2499,N_2430,N_2401);
or U2500 (N_2500,N_2435,N_2473);
or U2501 (N_2501,N_2413,N_2428);
nand U2502 (N_2502,N_2463,N_2464);
and U2503 (N_2503,N_2474,N_2408);
and U2504 (N_2504,N_2450,N_2406);
nor U2505 (N_2505,N_2465,N_2425);
or U2506 (N_2506,N_2462,N_2454);
nor U2507 (N_2507,N_2410,N_2405);
nor U2508 (N_2508,N_2427,N_2402);
nand U2509 (N_2509,N_2411,N_2436);
or U2510 (N_2510,N_2448,N_2403);
or U2511 (N_2511,N_2421,N_2415);
nor U2512 (N_2512,N_2467,N_2400);
or U2513 (N_2513,N_2453,N_2408);
nand U2514 (N_2514,N_2406,N_2474);
nor U2515 (N_2515,N_2442,N_2409);
nor U2516 (N_2516,N_2422,N_2454);
nand U2517 (N_2517,N_2437,N_2402);
and U2518 (N_2518,N_2466,N_2405);
nand U2519 (N_2519,N_2421,N_2437);
nor U2520 (N_2520,N_2445,N_2474);
nor U2521 (N_2521,N_2439,N_2409);
nor U2522 (N_2522,N_2445,N_2468);
and U2523 (N_2523,N_2425,N_2457);
or U2524 (N_2524,N_2445,N_2408);
nor U2525 (N_2525,N_2435,N_2446);
nand U2526 (N_2526,N_2415,N_2462);
nor U2527 (N_2527,N_2431,N_2400);
nand U2528 (N_2528,N_2407,N_2453);
or U2529 (N_2529,N_2455,N_2469);
or U2530 (N_2530,N_2466,N_2437);
nand U2531 (N_2531,N_2440,N_2428);
or U2532 (N_2532,N_2443,N_2406);
and U2533 (N_2533,N_2419,N_2457);
nand U2534 (N_2534,N_2460,N_2402);
and U2535 (N_2535,N_2436,N_2415);
nand U2536 (N_2536,N_2449,N_2411);
nand U2537 (N_2537,N_2460,N_2462);
nor U2538 (N_2538,N_2434,N_2410);
nand U2539 (N_2539,N_2444,N_2451);
nand U2540 (N_2540,N_2470,N_2418);
and U2541 (N_2541,N_2454,N_2412);
nand U2542 (N_2542,N_2429,N_2453);
nand U2543 (N_2543,N_2453,N_2444);
and U2544 (N_2544,N_2436,N_2458);
or U2545 (N_2545,N_2443,N_2429);
or U2546 (N_2546,N_2446,N_2445);
nand U2547 (N_2547,N_2405,N_2461);
nor U2548 (N_2548,N_2419,N_2468);
nand U2549 (N_2549,N_2452,N_2438);
nand U2550 (N_2550,N_2481,N_2521);
nand U2551 (N_2551,N_2543,N_2515);
and U2552 (N_2552,N_2530,N_2545);
nor U2553 (N_2553,N_2502,N_2520);
nor U2554 (N_2554,N_2497,N_2536);
or U2555 (N_2555,N_2505,N_2510);
nor U2556 (N_2556,N_2507,N_2525);
or U2557 (N_2557,N_2504,N_2477);
and U2558 (N_2558,N_2526,N_2540);
nor U2559 (N_2559,N_2508,N_2522);
nor U2560 (N_2560,N_2482,N_2513);
nor U2561 (N_2561,N_2541,N_2548);
nand U2562 (N_2562,N_2489,N_2511);
nand U2563 (N_2563,N_2546,N_2542);
nor U2564 (N_2564,N_2498,N_2528);
or U2565 (N_2565,N_2537,N_2492);
or U2566 (N_2566,N_2514,N_2493);
nand U2567 (N_2567,N_2517,N_2488);
and U2568 (N_2568,N_2500,N_2523);
nand U2569 (N_2569,N_2547,N_2479);
nor U2570 (N_2570,N_2527,N_2509);
nor U2571 (N_2571,N_2539,N_2495);
or U2572 (N_2572,N_2501,N_2538);
nor U2573 (N_2573,N_2483,N_2529);
nor U2574 (N_2574,N_2478,N_2512);
or U2575 (N_2575,N_2519,N_2518);
xnor U2576 (N_2576,N_2496,N_2549);
nor U2577 (N_2577,N_2476,N_2531);
nand U2578 (N_2578,N_2486,N_2480);
or U2579 (N_2579,N_2491,N_2485);
nand U2580 (N_2580,N_2506,N_2532);
nor U2581 (N_2581,N_2484,N_2494);
nand U2582 (N_2582,N_2503,N_2490);
xor U2583 (N_2583,N_2516,N_2475);
nand U2584 (N_2584,N_2524,N_2544);
nand U2585 (N_2585,N_2487,N_2533);
nor U2586 (N_2586,N_2499,N_2535);
nand U2587 (N_2587,N_2534,N_2527);
nor U2588 (N_2588,N_2476,N_2538);
nand U2589 (N_2589,N_2495,N_2508);
nor U2590 (N_2590,N_2479,N_2549);
nand U2591 (N_2591,N_2484,N_2477);
and U2592 (N_2592,N_2525,N_2484);
and U2593 (N_2593,N_2480,N_2479);
nor U2594 (N_2594,N_2485,N_2493);
and U2595 (N_2595,N_2504,N_2502);
or U2596 (N_2596,N_2532,N_2496);
nor U2597 (N_2597,N_2538,N_2533);
and U2598 (N_2598,N_2485,N_2549);
and U2599 (N_2599,N_2530,N_2518);
nor U2600 (N_2600,N_2505,N_2497);
or U2601 (N_2601,N_2545,N_2491);
or U2602 (N_2602,N_2480,N_2533);
or U2603 (N_2603,N_2488,N_2522);
and U2604 (N_2604,N_2494,N_2508);
nand U2605 (N_2605,N_2546,N_2505);
nand U2606 (N_2606,N_2538,N_2532);
and U2607 (N_2607,N_2540,N_2511);
and U2608 (N_2608,N_2511,N_2503);
and U2609 (N_2609,N_2519,N_2509);
nor U2610 (N_2610,N_2523,N_2512);
and U2611 (N_2611,N_2511,N_2522);
nor U2612 (N_2612,N_2498,N_2521);
and U2613 (N_2613,N_2516,N_2508);
and U2614 (N_2614,N_2539,N_2510);
and U2615 (N_2615,N_2544,N_2481);
and U2616 (N_2616,N_2509,N_2493);
and U2617 (N_2617,N_2547,N_2526);
nor U2618 (N_2618,N_2501,N_2514);
or U2619 (N_2619,N_2533,N_2525);
nand U2620 (N_2620,N_2505,N_2529);
nor U2621 (N_2621,N_2493,N_2523);
nand U2622 (N_2622,N_2518,N_2482);
nand U2623 (N_2623,N_2511,N_2514);
and U2624 (N_2624,N_2502,N_2528);
or U2625 (N_2625,N_2569,N_2603);
nor U2626 (N_2626,N_2568,N_2621);
nand U2627 (N_2627,N_2615,N_2551);
and U2628 (N_2628,N_2573,N_2587);
nand U2629 (N_2629,N_2586,N_2622);
nand U2630 (N_2630,N_2620,N_2584);
or U2631 (N_2631,N_2578,N_2552);
or U2632 (N_2632,N_2598,N_2590);
or U2633 (N_2633,N_2588,N_2604);
nand U2634 (N_2634,N_2557,N_2567);
nand U2635 (N_2635,N_2606,N_2610);
or U2636 (N_2636,N_2563,N_2577);
or U2637 (N_2637,N_2599,N_2592);
nor U2638 (N_2638,N_2601,N_2614);
nor U2639 (N_2639,N_2561,N_2612);
xnor U2640 (N_2640,N_2560,N_2596);
or U2641 (N_2641,N_2575,N_2609);
nor U2642 (N_2642,N_2616,N_2623);
nor U2643 (N_2643,N_2576,N_2585);
nand U2644 (N_2644,N_2559,N_2555);
or U2645 (N_2645,N_2591,N_2564);
nand U2646 (N_2646,N_2571,N_2593);
and U2647 (N_2647,N_2583,N_2562);
nor U2648 (N_2648,N_2611,N_2618);
nor U2649 (N_2649,N_2608,N_2579);
nand U2650 (N_2650,N_2597,N_2589);
or U2651 (N_2651,N_2565,N_2550);
nand U2652 (N_2652,N_2617,N_2566);
nor U2653 (N_2653,N_2580,N_2595);
nand U2654 (N_2654,N_2607,N_2556);
nand U2655 (N_2655,N_2554,N_2619);
nand U2656 (N_2656,N_2574,N_2624);
nand U2657 (N_2657,N_2613,N_2594);
nor U2658 (N_2658,N_2558,N_2553);
nand U2659 (N_2659,N_2602,N_2582);
and U2660 (N_2660,N_2600,N_2581);
nor U2661 (N_2661,N_2570,N_2572);
nor U2662 (N_2662,N_2605,N_2590);
or U2663 (N_2663,N_2553,N_2551);
or U2664 (N_2664,N_2586,N_2588);
nand U2665 (N_2665,N_2618,N_2559);
or U2666 (N_2666,N_2609,N_2624);
xnor U2667 (N_2667,N_2560,N_2551);
and U2668 (N_2668,N_2578,N_2579);
nor U2669 (N_2669,N_2552,N_2550);
and U2670 (N_2670,N_2553,N_2550);
nand U2671 (N_2671,N_2567,N_2564);
and U2672 (N_2672,N_2607,N_2578);
nor U2673 (N_2673,N_2590,N_2621);
and U2674 (N_2674,N_2577,N_2610);
or U2675 (N_2675,N_2569,N_2576);
or U2676 (N_2676,N_2591,N_2570);
nand U2677 (N_2677,N_2584,N_2606);
and U2678 (N_2678,N_2564,N_2624);
nor U2679 (N_2679,N_2624,N_2584);
nor U2680 (N_2680,N_2613,N_2583);
xor U2681 (N_2681,N_2579,N_2551);
nand U2682 (N_2682,N_2612,N_2582);
nor U2683 (N_2683,N_2572,N_2591);
nand U2684 (N_2684,N_2614,N_2609);
and U2685 (N_2685,N_2580,N_2592);
nor U2686 (N_2686,N_2590,N_2570);
nor U2687 (N_2687,N_2579,N_2598);
or U2688 (N_2688,N_2575,N_2567);
nor U2689 (N_2689,N_2561,N_2565);
nor U2690 (N_2690,N_2589,N_2564);
and U2691 (N_2691,N_2554,N_2583);
or U2692 (N_2692,N_2563,N_2592);
xnor U2693 (N_2693,N_2582,N_2567);
nand U2694 (N_2694,N_2566,N_2587);
and U2695 (N_2695,N_2552,N_2622);
nor U2696 (N_2696,N_2550,N_2622);
and U2697 (N_2697,N_2568,N_2556);
nand U2698 (N_2698,N_2614,N_2584);
nand U2699 (N_2699,N_2591,N_2592);
nor U2700 (N_2700,N_2682,N_2664);
nor U2701 (N_2701,N_2628,N_2662);
or U2702 (N_2702,N_2696,N_2688);
nor U2703 (N_2703,N_2694,N_2690);
nor U2704 (N_2704,N_2669,N_2645);
nand U2705 (N_2705,N_2683,N_2698);
and U2706 (N_2706,N_2685,N_2625);
and U2707 (N_2707,N_2660,N_2686);
nor U2708 (N_2708,N_2678,N_2632);
nand U2709 (N_2709,N_2648,N_2674);
and U2710 (N_2710,N_2680,N_2647);
nand U2711 (N_2711,N_2659,N_2691);
or U2712 (N_2712,N_2644,N_2689);
and U2713 (N_2713,N_2675,N_2677);
nand U2714 (N_2714,N_2642,N_2697);
nor U2715 (N_2715,N_2641,N_2699);
nor U2716 (N_2716,N_2672,N_2657);
and U2717 (N_2717,N_2668,N_2654);
nand U2718 (N_2718,N_2646,N_2665);
nand U2719 (N_2719,N_2629,N_2666);
nor U2720 (N_2720,N_2663,N_2676);
or U2721 (N_2721,N_2635,N_2633);
nand U2722 (N_2722,N_2695,N_2653);
nor U2723 (N_2723,N_2679,N_2693);
nor U2724 (N_2724,N_2630,N_2636);
nor U2725 (N_2725,N_2638,N_2634);
nor U2726 (N_2726,N_2692,N_2652);
nand U2727 (N_2727,N_2627,N_2656);
and U2728 (N_2728,N_2687,N_2637);
nand U2729 (N_2729,N_2650,N_2640);
and U2730 (N_2730,N_2667,N_2626);
and U2731 (N_2731,N_2661,N_2631);
or U2732 (N_2732,N_2655,N_2681);
nand U2733 (N_2733,N_2643,N_2670);
or U2734 (N_2734,N_2658,N_2684);
nand U2735 (N_2735,N_2639,N_2673);
nor U2736 (N_2736,N_2651,N_2671);
nand U2737 (N_2737,N_2649,N_2633);
nand U2738 (N_2738,N_2656,N_2642);
or U2739 (N_2739,N_2693,N_2699);
nand U2740 (N_2740,N_2643,N_2651);
or U2741 (N_2741,N_2691,N_2699);
nor U2742 (N_2742,N_2664,N_2680);
or U2743 (N_2743,N_2638,N_2656);
nand U2744 (N_2744,N_2631,N_2656);
nand U2745 (N_2745,N_2645,N_2637);
nor U2746 (N_2746,N_2642,N_2644);
or U2747 (N_2747,N_2630,N_2657);
nor U2748 (N_2748,N_2638,N_2659);
nor U2749 (N_2749,N_2692,N_2685);
or U2750 (N_2750,N_2656,N_2650);
nand U2751 (N_2751,N_2646,N_2689);
xnor U2752 (N_2752,N_2684,N_2637);
nor U2753 (N_2753,N_2686,N_2676);
and U2754 (N_2754,N_2639,N_2628);
or U2755 (N_2755,N_2694,N_2650);
and U2756 (N_2756,N_2698,N_2681);
nor U2757 (N_2757,N_2668,N_2693);
and U2758 (N_2758,N_2666,N_2687);
or U2759 (N_2759,N_2689,N_2649);
and U2760 (N_2760,N_2670,N_2646);
nand U2761 (N_2761,N_2666,N_2641);
and U2762 (N_2762,N_2670,N_2655);
nor U2763 (N_2763,N_2694,N_2629);
nand U2764 (N_2764,N_2635,N_2662);
nor U2765 (N_2765,N_2655,N_2635);
or U2766 (N_2766,N_2641,N_2650);
and U2767 (N_2767,N_2649,N_2641);
or U2768 (N_2768,N_2654,N_2661);
nor U2769 (N_2769,N_2629,N_2633);
nand U2770 (N_2770,N_2641,N_2689);
and U2771 (N_2771,N_2693,N_2675);
and U2772 (N_2772,N_2671,N_2667);
nor U2773 (N_2773,N_2678,N_2629);
or U2774 (N_2774,N_2638,N_2664);
nor U2775 (N_2775,N_2734,N_2700);
nand U2776 (N_2776,N_2760,N_2747);
nor U2777 (N_2777,N_2744,N_2763);
or U2778 (N_2778,N_2758,N_2735);
and U2779 (N_2779,N_2733,N_2752);
and U2780 (N_2780,N_2739,N_2743);
and U2781 (N_2781,N_2759,N_2770);
nand U2782 (N_2782,N_2742,N_2745);
nand U2783 (N_2783,N_2772,N_2730);
nand U2784 (N_2784,N_2765,N_2709);
and U2785 (N_2785,N_2714,N_2726);
or U2786 (N_2786,N_2773,N_2713);
nor U2787 (N_2787,N_2728,N_2707);
nor U2788 (N_2788,N_2718,N_2704);
nor U2789 (N_2789,N_2725,N_2729);
or U2790 (N_2790,N_2757,N_2736);
and U2791 (N_2791,N_2762,N_2703);
nor U2792 (N_2792,N_2719,N_2767);
or U2793 (N_2793,N_2724,N_2740);
nand U2794 (N_2794,N_2755,N_2761);
nand U2795 (N_2795,N_2769,N_2701);
nand U2796 (N_2796,N_2723,N_2721);
nor U2797 (N_2797,N_2750,N_2722);
and U2798 (N_2798,N_2738,N_2753);
or U2799 (N_2799,N_2717,N_2708);
nand U2800 (N_2800,N_2766,N_2712);
or U2801 (N_2801,N_2749,N_2768);
nor U2802 (N_2802,N_2764,N_2727);
and U2803 (N_2803,N_2746,N_2771);
nand U2804 (N_2804,N_2710,N_2732);
or U2805 (N_2805,N_2720,N_2716);
and U2806 (N_2806,N_2774,N_2702);
and U2807 (N_2807,N_2748,N_2741);
or U2808 (N_2808,N_2731,N_2705);
xor U2809 (N_2809,N_2711,N_2751);
and U2810 (N_2810,N_2737,N_2706);
nand U2811 (N_2811,N_2756,N_2715);
xnor U2812 (N_2812,N_2754,N_2758);
or U2813 (N_2813,N_2736,N_2722);
and U2814 (N_2814,N_2702,N_2743);
and U2815 (N_2815,N_2715,N_2752);
nor U2816 (N_2816,N_2760,N_2702);
or U2817 (N_2817,N_2708,N_2710);
or U2818 (N_2818,N_2774,N_2747);
xnor U2819 (N_2819,N_2767,N_2762);
nor U2820 (N_2820,N_2701,N_2747);
nor U2821 (N_2821,N_2737,N_2773);
and U2822 (N_2822,N_2708,N_2735);
or U2823 (N_2823,N_2721,N_2757);
or U2824 (N_2824,N_2710,N_2740);
and U2825 (N_2825,N_2716,N_2703);
or U2826 (N_2826,N_2741,N_2710);
or U2827 (N_2827,N_2701,N_2723);
nand U2828 (N_2828,N_2730,N_2766);
or U2829 (N_2829,N_2744,N_2767);
or U2830 (N_2830,N_2733,N_2712);
or U2831 (N_2831,N_2774,N_2719);
nand U2832 (N_2832,N_2711,N_2762);
or U2833 (N_2833,N_2728,N_2744);
or U2834 (N_2834,N_2760,N_2767);
nor U2835 (N_2835,N_2732,N_2709);
nand U2836 (N_2836,N_2736,N_2730);
nand U2837 (N_2837,N_2730,N_2719);
and U2838 (N_2838,N_2708,N_2743);
and U2839 (N_2839,N_2706,N_2725);
or U2840 (N_2840,N_2763,N_2751);
nand U2841 (N_2841,N_2747,N_2753);
nand U2842 (N_2842,N_2742,N_2723);
and U2843 (N_2843,N_2714,N_2765);
nor U2844 (N_2844,N_2740,N_2726);
nand U2845 (N_2845,N_2748,N_2722);
and U2846 (N_2846,N_2747,N_2765);
or U2847 (N_2847,N_2722,N_2743);
and U2848 (N_2848,N_2714,N_2712);
nor U2849 (N_2849,N_2761,N_2709);
nand U2850 (N_2850,N_2817,N_2782);
nor U2851 (N_2851,N_2823,N_2842);
and U2852 (N_2852,N_2848,N_2839);
nand U2853 (N_2853,N_2776,N_2779);
or U2854 (N_2854,N_2814,N_2820);
nand U2855 (N_2855,N_2818,N_2808);
nor U2856 (N_2856,N_2780,N_2796);
nand U2857 (N_2857,N_2813,N_2788);
nand U2858 (N_2858,N_2834,N_2836);
or U2859 (N_2859,N_2821,N_2790);
nand U2860 (N_2860,N_2830,N_2806);
and U2861 (N_2861,N_2822,N_2811);
and U2862 (N_2862,N_2827,N_2843);
nand U2863 (N_2863,N_2802,N_2799);
nand U2864 (N_2864,N_2835,N_2792);
or U2865 (N_2865,N_2801,N_2837);
nor U2866 (N_2866,N_2825,N_2833);
nand U2867 (N_2867,N_2828,N_2778);
nand U2868 (N_2868,N_2805,N_2845);
or U2869 (N_2869,N_2812,N_2798);
nor U2870 (N_2870,N_2791,N_2777);
or U2871 (N_2871,N_2838,N_2829);
nand U2872 (N_2872,N_2844,N_2819);
and U2873 (N_2873,N_2831,N_2786);
xor U2874 (N_2874,N_2832,N_2840);
or U2875 (N_2875,N_2787,N_2815);
or U2876 (N_2876,N_2775,N_2816);
nand U2877 (N_2877,N_2794,N_2793);
nor U2878 (N_2878,N_2826,N_2797);
or U2879 (N_2879,N_2849,N_2841);
nand U2880 (N_2880,N_2803,N_2847);
nand U2881 (N_2881,N_2824,N_2785);
and U2882 (N_2882,N_2809,N_2810);
nand U2883 (N_2883,N_2807,N_2783);
or U2884 (N_2884,N_2789,N_2846);
xnor U2885 (N_2885,N_2804,N_2795);
and U2886 (N_2886,N_2784,N_2800);
or U2887 (N_2887,N_2781,N_2836);
nor U2888 (N_2888,N_2787,N_2781);
or U2889 (N_2889,N_2789,N_2836);
nand U2890 (N_2890,N_2841,N_2799);
and U2891 (N_2891,N_2839,N_2777);
or U2892 (N_2892,N_2799,N_2793);
nand U2893 (N_2893,N_2812,N_2808);
or U2894 (N_2894,N_2776,N_2789);
nor U2895 (N_2895,N_2822,N_2789);
and U2896 (N_2896,N_2831,N_2810);
nand U2897 (N_2897,N_2790,N_2833);
nand U2898 (N_2898,N_2809,N_2844);
or U2899 (N_2899,N_2838,N_2783);
nand U2900 (N_2900,N_2808,N_2776);
or U2901 (N_2901,N_2821,N_2820);
nand U2902 (N_2902,N_2835,N_2781);
nor U2903 (N_2903,N_2830,N_2808);
and U2904 (N_2904,N_2775,N_2788);
and U2905 (N_2905,N_2791,N_2810);
and U2906 (N_2906,N_2792,N_2800);
nand U2907 (N_2907,N_2816,N_2846);
nor U2908 (N_2908,N_2812,N_2819);
nor U2909 (N_2909,N_2836,N_2829);
nand U2910 (N_2910,N_2849,N_2779);
or U2911 (N_2911,N_2810,N_2844);
nor U2912 (N_2912,N_2800,N_2828);
and U2913 (N_2913,N_2814,N_2845);
nand U2914 (N_2914,N_2848,N_2811);
nand U2915 (N_2915,N_2845,N_2825);
or U2916 (N_2916,N_2835,N_2809);
and U2917 (N_2917,N_2788,N_2817);
nand U2918 (N_2918,N_2835,N_2811);
and U2919 (N_2919,N_2830,N_2835);
nor U2920 (N_2920,N_2832,N_2813);
nand U2921 (N_2921,N_2781,N_2818);
or U2922 (N_2922,N_2826,N_2780);
or U2923 (N_2923,N_2815,N_2835);
or U2924 (N_2924,N_2808,N_2825);
and U2925 (N_2925,N_2885,N_2870);
nor U2926 (N_2926,N_2865,N_2891);
nor U2927 (N_2927,N_2893,N_2867);
nor U2928 (N_2928,N_2854,N_2918);
nand U2929 (N_2929,N_2878,N_2859);
nor U2930 (N_2930,N_2880,N_2875);
and U2931 (N_2931,N_2905,N_2901);
and U2932 (N_2932,N_2889,N_2904);
nand U2933 (N_2933,N_2862,N_2913);
nor U2934 (N_2934,N_2886,N_2858);
and U2935 (N_2935,N_2884,N_2871);
and U2936 (N_2936,N_2908,N_2917);
or U2937 (N_2937,N_2922,N_2907);
and U2938 (N_2938,N_2890,N_2914);
nand U2939 (N_2939,N_2851,N_2912);
and U2940 (N_2940,N_2916,N_2911);
or U2941 (N_2941,N_2902,N_2877);
or U2942 (N_2942,N_2864,N_2900);
nor U2943 (N_2943,N_2883,N_2899);
and U2944 (N_2944,N_2903,N_2873);
and U2945 (N_2945,N_2898,N_2892);
or U2946 (N_2946,N_2909,N_2850);
and U2947 (N_2947,N_2872,N_2923);
nor U2948 (N_2948,N_2879,N_2882);
nor U2949 (N_2949,N_2915,N_2869);
nand U2950 (N_2950,N_2852,N_2857);
and U2951 (N_2951,N_2874,N_2921);
or U2952 (N_2952,N_2920,N_2861);
or U2953 (N_2953,N_2866,N_2856);
nand U2954 (N_2954,N_2863,N_2868);
or U2955 (N_2955,N_2906,N_2919);
or U2956 (N_2956,N_2881,N_2887);
nand U2957 (N_2957,N_2895,N_2924);
or U2958 (N_2958,N_2894,N_2896);
nor U2959 (N_2959,N_2876,N_2888);
or U2960 (N_2960,N_2860,N_2855);
or U2961 (N_2961,N_2910,N_2853);
or U2962 (N_2962,N_2897,N_2910);
or U2963 (N_2963,N_2899,N_2878);
and U2964 (N_2964,N_2901,N_2877);
and U2965 (N_2965,N_2887,N_2904);
nor U2966 (N_2966,N_2889,N_2885);
nand U2967 (N_2967,N_2866,N_2867);
or U2968 (N_2968,N_2852,N_2892);
nand U2969 (N_2969,N_2867,N_2858);
or U2970 (N_2970,N_2919,N_2907);
nor U2971 (N_2971,N_2892,N_2865);
and U2972 (N_2972,N_2875,N_2867);
and U2973 (N_2973,N_2905,N_2883);
or U2974 (N_2974,N_2923,N_2860);
or U2975 (N_2975,N_2857,N_2911);
nor U2976 (N_2976,N_2872,N_2870);
or U2977 (N_2977,N_2870,N_2906);
and U2978 (N_2978,N_2903,N_2866);
nand U2979 (N_2979,N_2871,N_2900);
or U2980 (N_2980,N_2894,N_2913);
nand U2981 (N_2981,N_2852,N_2916);
and U2982 (N_2982,N_2864,N_2866);
and U2983 (N_2983,N_2851,N_2889);
or U2984 (N_2984,N_2901,N_2872);
nand U2985 (N_2985,N_2859,N_2867);
or U2986 (N_2986,N_2901,N_2871);
nand U2987 (N_2987,N_2915,N_2881);
and U2988 (N_2988,N_2900,N_2907);
nand U2989 (N_2989,N_2870,N_2909);
and U2990 (N_2990,N_2896,N_2868);
or U2991 (N_2991,N_2863,N_2901);
or U2992 (N_2992,N_2856,N_2906);
or U2993 (N_2993,N_2872,N_2893);
or U2994 (N_2994,N_2850,N_2892);
or U2995 (N_2995,N_2904,N_2913);
and U2996 (N_2996,N_2895,N_2900);
nor U2997 (N_2997,N_2870,N_2868);
or U2998 (N_2998,N_2866,N_2888);
nor U2999 (N_2999,N_2866,N_2889);
nor UO_0 (O_0,N_2950,N_2996);
or UO_1 (O_1,N_2959,N_2969);
and UO_2 (O_2,N_2948,N_2986);
nand UO_3 (O_3,N_2975,N_2929);
and UO_4 (O_4,N_2983,N_2925);
and UO_5 (O_5,N_2928,N_2935);
nand UO_6 (O_6,N_2961,N_2943);
and UO_7 (O_7,N_2968,N_2990);
or UO_8 (O_8,N_2963,N_2953);
nand UO_9 (O_9,N_2973,N_2984);
nor UO_10 (O_10,N_2978,N_2998);
and UO_11 (O_11,N_2945,N_2992);
nor UO_12 (O_12,N_2966,N_2952);
or UO_13 (O_13,N_2988,N_2997);
and UO_14 (O_14,N_2937,N_2977);
and UO_15 (O_15,N_2960,N_2989);
and UO_16 (O_16,N_2930,N_2962);
or UO_17 (O_17,N_2934,N_2941);
nor UO_18 (O_18,N_2933,N_2931);
and UO_19 (O_19,N_2991,N_2995);
nand UO_20 (O_20,N_2985,N_2965);
nor UO_21 (O_21,N_2976,N_2944);
nand UO_22 (O_22,N_2993,N_2954);
or UO_23 (O_23,N_2932,N_2926);
xor UO_24 (O_24,N_2970,N_2946);
nand UO_25 (O_25,N_2964,N_2956);
nand UO_26 (O_26,N_2940,N_2936);
or UO_27 (O_27,N_2999,N_2974);
and UO_28 (O_28,N_2949,N_2955);
and UO_29 (O_29,N_2947,N_2927);
nor UO_30 (O_30,N_2979,N_2994);
nand UO_31 (O_31,N_2957,N_2942);
or UO_32 (O_32,N_2987,N_2951);
and UO_33 (O_33,N_2982,N_2972);
nand UO_34 (O_34,N_2967,N_2981);
nand UO_35 (O_35,N_2980,N_2938);
and UO_36 (O_36,N_2958,N_2971);
and UO_37 (O_37,N_2939,N_2964);
and UO_38 (O_38,N_2951,N_2941);
nand UO_39 (O_39,N_2962,N_2926);
nand UO_40 (O_40,N_2991,N_2982);
and UO_41 (O_41,N_2987,N_2954);
nor UO_42 (O_42,N_2981,N_2994);
nor UO_43 (O_43,N_2944,N_2980);
nor UO_44 (O_44,N_2941,N_2985);
or UO_45 (O_45,N_2982,N_2999);
and UO_46 (O_46,N_2965,N_2996);
nand UO_47 (O_47,N_2980,N_2987);
or UO_48 (O_48,N_2961,N_2997);
nor UO_49 (O_49,N_2981,N_2980);
nor UO_50 (O_50,N_2969,N_2970);
or UO_51 (O_51,N_2995,N_2975);
and UO_52 (O_52,N_2925,N_2940);
and UO_53 (O_53,N_2952,N_2967);
or UO_54 (O_54,N_2942,N_2993);
and UO_55 (O_55,N_2929,N_2946);
and UO_56 (O_56,N_2927,N_2971);
nor UO_57 (O_57,N_2972,N_2945);
or UO_58 (O_58,N_2977,N_2957);
or UO_59 (O_59,N_2944,N_2969);
and UO_60 (O_60,N_2951,N_2929);
or UO_61 (O_61,N_2932,N_2927);
nor UO_62 (O_62,N_2999,N_2927);
nor UO_63 (O_63,N_2964,N_2995);
nor UO_64 (O_64,N_2980,N_2940);
nand UO_65 (O_65,N_2986,N_2991);
or UO_66 (O_66,N_2999,N_2971);
nand UO_67 (O_67,N_2982,N_2973);
nand UO_68 (O_68,N_2994,N_2960);
nand UO_69 (O_69,N_2980,N_2925);
nor UO_70 (O_70,N_2941,N_2964);
nor UO_71 (O_71,N_2999,N_2979);
nor UO_72 (O_72,N_2971,N_2940);
or UO_73 (O_73,N_2947,N_2985);
nor UO_74 (O_74,N_2941,N_2961);
nand UO_75 (O_75,N_2996,N_2980);
xnor UO_76 (O_76,N_2975,N_2972);
or UO_77 (O_77,N_2955,N_2975);
and UO_78 (O_78,N_2998,N_2954);
and UO_79 (O_79,N_2944,N_2972);
or UO_80 (O_80,N_2989,N_2994);
nor UO_81 (O_81,N_2935,N_2957);
nor UO_82 (O_82,N_2980,N_2991);
xor UO_83 (O_83,N_2942,N_2943);
nand UO_84 (O_84,N_2998,N_2990);
or UO_85 (O_85,N_2948,N_2933);
and UO_86 (O_86,N_2988,N_2943);
and UO_87 (O_87,N_2971,N_2985);
nand UO_88 (O_88,N_2990,N_2949);
and UO_89 (O_89,N_2967,N_2928);
nor UO_90 (O_90,N_2948,N_2950);
nand UO_91 (O_91,N_2979,N_2963);
nor UO_92 (O_92,N_2926,N_2995);
nor UO_93 (O_93,N_2965,N_2983);
nor UO_94 (O_94,N_2981,N_2990);
nand UO_95 (O_95,N_2953,N_2999);
nand UO_96 (O_96,N_2947,N_2937);
nor UO_97 (O_97,N_2925,N_2953);
or UO_98 (O_98,N_2955,N_2992);
or UO_99 (O_99,N_2941,N_2960);
or UO_100 (O_100,N_2991,N_2937);
and UO_101 (O_101,N_2973,N_2956);
nand UO_102 (O_102,N_2994,N_2929);
nand UO_103 (O_103,N_2992,N_2944);
and UO_104 (O_104,N_2992,N_2959);
nor UO_105 (O_105,N_2958,N_2926);
or UO_106 (O_106,N_2953,N_2995);
nand UO_107 (O_107,N_2993,N_2985);
nor UO_108 (O_108,N_2987,N_2978);
nor UO_109 (O_109,N_2991,N_2927);
nand UO_110 (O_110,N_2936,N_2950);
xnor UO_111 (O_111,N_2935,N_2991);
or UO_112 (O_112,N_2928,N_2933);
nor UO_113 (O_113,N_2933,N_2966);
and UO_114 (O_114,N_2929,N_2995);
or UO_115 (O_115,N_2933,N_2932);
nand UO_116 (O_116,N_2968,N_2982);
and UO_117 (O_117,N_2974,N_2927);
or UO_118 (O_118,N_2951,N_2949);
nor UO_119 (O_119,N_2926,N_2950);
nand UO_120 (O_120,N_2987,N_2955);
or UO_121 (O_121,N_2997,N_2999);
nand UO_122 (O_122,N_2934,N_2955);
nand UO_123 (O_123,N_2930,N_2964);
and UO_124 (O_124,N_2957,N_2933);
nor UO_125 (O_125,N_2995,N_2959);
or UO_126 (O_126,N_2979,N_2993);
xnor UO_127 (O_127,N_2972,N_2942);
or UO_128 (O_128,N_2947,N_2970);
and UO_129 (O_129,N_2978,N_2938);
nor UO_130 (O_130,N_2964,N_2961);
nor UO_131 (O_131,N_2968,N_2987);
or UO_132 (O_132,N_2974,N_2992);
nor UO_133 (O_133,N_2994,N_2993);
nand UO_134 (O_134,N_2967,N_2942);
or UO_135 (O_135,N_2974,N_2987);
or UO_136 (O_136,N_2941,N_2995);
nand UO_137 (O_137,N_2931,N_2950);
and UO_138 (O_138,N_2999,N_2937);
and UO_139 (O_139,N_2996,N_2949);
nor UO_140 (O_140,N_2927,N_2930);
nor UO_141 (O_141,N_2939,N_2981);
nand UO_142 (O_142,N_2999,N_2930);
nor UO_143 (O_143,N_2973,N_2979);
or UO_144 (O_144,N_2997,N_2975);
nor UO_145 (O_145,N_2972,N_2991);
or UO_146 (O_146,N_2990,N_2985);
nor UO_147 (O_147,N_2991,N_2985);
nor UO_148 (O_148,N_2955,N_2969);
nor UO_149 (O_149,N_2991,N_2950);
or UO_150 (O_150,N_2950,N_2929);
or UO_151 (O_151,N_2972,N_2941);
and UO_152 (O_152,N_2944,N_2934);
nand UO_153 (O_153,N_2986,N_2972);
or UO_154 (O_154,N_2951,N_2984);
nor UO_155 (O_155,N_2994,N_2987);
or UO_156 (O_156,N_2996,N_2938);
nand UO_157 (O_157,N_2983,N_2962);
nor UO_158 (O_158,N_2979,N_2937);
nor UO_159 (O_159,N_2957,N_2928);
nor UO_160 (O_160,N_2993,N_2958);
and UO_161 (O_161,N_2936,N_2934);
nand UO_162 (O_162,N_2947,N_2990);
nor UO_163 (O_163,N_2936,N_2980);
nand UO_164 (O_164,N_2942,N_2963);
nand UO_165 (O_165,N_2993,N_2973);
nor UO_166 (O_166,N_2972,N_2952);
nand UO_167 (O_167,N_2945,N_2984);
nor UO_168 (O_168,N_2925,N_2973);
or UO_169 (O_169,N_2947,N_2981);
and UO_170 (O_170,N_2925,N_2952);
or UO_171 (O_171,N_2957,N_2999);
or UO_172 (O_172,N_2936,N_2973);
nand UO_173 (O_173,N_2984,N_2930);
nand UO_174 (O_174,N_2984,N_2971);
nand UO_175 (O_175,N_2925,N_2988);
nor UO_176 (O_176,N_2944,N_2968);
nor UO_177 (O_177,N_2936,N_2931);
nor UO_178 (O_178,N_2995,N_2961);
nor UO_179 (O_179,N_2999,N_2988);
and UO_180 (O_180,N_2979,N_2934);
nor UO_181 (O_181,N_2929,N_2942);
nor UO_182 (O_182,N_2926,N_2966);
and UO_183 (O_183,N_2938,N_2963);
nand UO_184 (O_184,N_2970,N_2994);
nor UO_185 (O_185,N_2979,N_2941);
nand UO_186 (O_186,N_2954,N_2928);
xor UO_187 (O_187,N_2961,N_2981);
and UO_188 (O_188,N_2952,N_2989);
or UO_189 (O_189,N_2946,N_2973);
nor UO_190 (O_190,N_2953,N_2954);
or UO_191 (O_191,N_2942,N_2938);
nand UO_192 (O_192,N_2973,N_2962);
nand UO_193 (O_193,N_2953,N_2980);
nand UO_194 (O_194,N_2957,N_2970);
nand UO_195 (O_195,N_2948,N_2966);
nor UO_196 (O_196,N_2979,N_2952);
or UO_197 (O_197,N_2937,N_2970);
nand UO_198 (O_198,N_2990,N_2927);
and UO_199 (O_199,N_2953,N_2943);
nor UO_200 (O_200,N_2940,N_2958);
or UO_201 (O_201,N_2974,N_2984);
and UO_202 (O_202,N_2976,N_2966);
and UO_203 (O_203,N_2977,N_2993);
nor UO_204 (O_204,N_2962,N_2946);
and UO_205 (O_205,N_2998,N_2993);
or UO_206 (O_206,N_2961,N_2984);
nor UO_207 (O_207,N_2955,N_2945);
nand UO_208 (O_208,N_2937,N_2958);
or UO_209 (O_209,N_2944,N_2993);
or UO_210 (O_210,N_2956,N_2972);
or UO_211 (O_211,N_2961,N_2925);
nor UO_212 (O_212,N_2994,N_2969);
nand UO_213 (O_213,N_2932,N_2962);
and UO_214 (O_214,N_2966,N_2985);
nand UO_215 (O_215,N_2981,N_2962);
or UO_216 (O_216,N_2959,N_2971);
and UO_217 (O_217,N_2937,N_2925);
or UO_218 (O_218,N_2930,N_2966);
or UO_219 (O_219,N_2966,N_2997);
and UO_220 (O_220,N_2987,N_2948);
nand UO_221 (O_221,N_2960,N_2927);
or UO_222 (O_222,N_2974,N_2972);
nor UO_223 (O_223,N_2953,N_2951);
nand UO_224 (O_224,N_2960,N_2943);
and UO_225 (O_225,N_2939,N_2994);
nor UO_226 (O_226,N_2982,N_2940);
xor UO_227 (O_227,N_2933,N_2951);
nor UO_228 (O_228,N_2932,N_2952);
nor UO_229 (O_229,N_2935,N_2974);
and UO_230 (O_230,N_2970,N_2953);
or UO_231 (O_231,N_2979,N_2990);
and UO_232 (O_232,N_2927,N_2929);
or UO_233 (O_233,N_2999,N_2956);
nor UO_234 (O_234,N_2943,N_2968);
nor UO_235 (O_235,N_2941,N_2994);
and UO_236 (O_236,N_2927,N_2942);
or UO_237 (O_237,N_2956,N_2949);
or UO_238 (O_238,N_2950,N_2979);
nor UO_239 (O_239,N_2955,N_2988);
nor UO_240 (O_240,N_2956,N_2994);
nand UO_241 (O_241,N_2961,N_2934);
nor UO_242 (O_242,N_2967,N_2970);
or UO_243 (O_243,N_2929,N_2933);
nand UO_244 (O_244,N_2951,N_2957);
nand UO_245 (O_245,N_2939,N_2942);
or UO_246 (O_246,N_2955,N_2938);
nor UO_247 (O_247,N_2991,N_2967);
and UO_248 (O_248,N_2960,N_2959);
nor UO_249 (O_249,N_2959,N_2985);
and UO_250 (O_250,N_2963,N_2990);
nand UO_251 (O_251,N_2982,N_2944);
or UO_252 (O_252,N_2977,N_2949);
nor UO_253 (O_253,N_2981,N_2949);
nor UO_254 (O_254,N_2980,N_2958);
or UO_255 (O_255,N_2978,N_2957);
nor UO_256 (O_256,N_2969,N_2940);
and UO_257 (O_257,N_2957,N_2996);
nand UO_258 (O_258,N_2998,N_2951);
and UO_259 (O_259,N_2950,N_2949);
and UO_260 (O_260,N_2942,N_2926);
and UO_261 (O_261,N_2947,N_2938);
and UO_262 (O_262,N_2956,N_2958);
nor UO_263 (O_263,N_2971,N_2974);
and UO_264 (O_264,N_2996,N_2930);
nand UO_265 (O_265,N_2956,N_2926);
and UO_266 (O_266,N_2991,N_2958);
or UO_267 (O_267,N_2996,N_2961);
nand UO_268 (O_268,N_2973,N_2967);
nor UO_269 (O_269,N_2993,N_2986);
nor UO_270 (O_270,N_2967,N_2959);
nand UO_271 (O_271,N_2988,N_2927);
nand UO_272 (O_272,N_2998,N_2977);
nor UO_273 (O_273,N_2953,N_2961);
or UO_274 (O_274,N_2975,N_2974);
nand UO_275 (O_275,N_2983,N_2985);
nand UO_276 (O_276,N_2949,N_2997);
and UO_277 (O_277,N_2987,N_2925);
nand UO_278 (O_278,N_2963,N_2996);
or UO_279 (O_279,N_2928,N_2960);
nand UO_280 (O_280,N_2927,N_2969);
or UO_281 (O_281,N_2965,N_2949);
and UO_282 (O_282,N_2943,N_2980);
and UO_283 (O_283,N_2998,N_2981);
or UO_284 (O_284,N_2989,N_2950);
and UO_285 (O_285,N_2980,N_2941);
or UO_286 (O_286,N_2963,N_2934);
nand UO_287 (O_287,N_2959,N_2941);
nor UO_288 (O_288,N_2931,N_2980);
nor UO_289 (O_289,N_2970,N_2996);
and UO_290 (O_290,N_2932,N_2971);
or UO_291 (O_291,N_2961,N_2957);
or UO_292 (O_292,N_2935,N_2994);
nor UO_293 (O_293,N_2942,N_2940);
and UO_294 (O_294,N_2936,N_2961);
nand UO_295 (O_295,N_2975,N_2935);
nand UO_296 (O_296,N_2983,N_2980);
or UO_297 (O_297,N_2982,N_2932);
nand UO_298 (O_298,N_2970,N_2983);
nand UO_299 (O_299,N_2999,N_2975);
and UO_300 (O_300,N_2926,N_2927);
and UO_301 (O_301,N_2994,N_2928);
or UO_302 (O_302,N_2988,N_2946);
nor UO_303 (O_303,N_2959,N_2932);
or UO_304 (O_304,N_2933,N_2982);
nor UO_305 (O_305,N_2938,N_2985);
nor UO_306 (O_306,N_2970,N_2931);
nor UO_307 (O_307,N_2968,N_2928);
or UO_308 (O_308,N_2955,N_2965);
nand UO_309 (O_309,N_2934,N_2965);
or UO_310 (O_310,N_2926,N_2967);
nand UO_311 (O_311,N_2960,N_2963);
nand UO_312 (O_312,N_2957,N_2986);
nor UO_313 (O_313,N_2944,N_2966);
or UO_314 (O_314,N_2994,N_2988);
nand UO_315 (O_315,N_2955,N_2968);
and UO_316 (O_316,N_2987,N_2999);
nand UO_317 (O_317,N_2935,N_2954);
nand UO_318 (O_318,N_2993,N_2928);
nand UO_319 (O_319,N_2949,N_2983);
or UO_320 (O_320,N_2943,N_2938);
and UO_321 (O_321,N_2988,N_2989);
or UO_322 (O_322,N_2943,N_2996);
and UO_323 (O_323,N_2941,N_2978);
nand UO_324 (O_324,N_2991,N_2932);
nand UO_325 (O_325,N_2993,N_2940);
nor UO_326 (O_326,N_2996,N_2962);
nand UO_327 (O_327,N_2971,N_2975);
or UO_328 (O_328,N_2929,N_2964);
nand UO_329 (O_329,N_2997,N_2992);
nand UO_330 (O_330,N_2977,N_2988);
nor UO_331 (O_331,N_2999,N_2934);
nand UO_332 (O_332,N_2931,N_2961);
nor UO_333 (O_333,N_2946,N_2998);
nor UO_334 (O_334,N_2934,N_2945);
or UO_335 (O_335,N_2929,N_2962);
nor UO_336 (O_336,N_2952,N_2999);
nand UO_337 (O_337,N_2977,N_2958);
nand UO_338 (O_338,N_2945,N_2953);
nand UO_339 (O_339,N_2927,N_2978);
and UO_340 (O_340,N_2940,N_2954);
or UO_341 (O_341,N_2962,N_2971);
nand UO_342 (O_342,N_2955,N_2952);
or UO_343 (O_343,N_2946,N_2953);
nand UO_344 (O_344,N_2989,N_2941);
nand UO_345 (O_345,N_2974,N_2952);
or UO_346 (O_346,N_2936,N_2978);
xnor UO_347 (O_347,N_2925,N_2954);
nor UO_348 (O_348,N_2949,N_2942);
nand UO_349 (O_349,N_2971,N_2969);
or UO_350 (O_350,N_2977,N_2946);
nand UO_351 (O_351,N_2937,N_2938);
and UO_352 (O_352,N_2972,N_2989);
and UO_353 (O_353,N_2979,N_2970);
nand UO_354 (O_354,N_2987,N_2950);
nor UO_355 (O_355,N_2978,N_2996);
nor UO_356 (O_356,N_2931,N_2951);
nor UO_357 (O_357,N_2950,N_2998);
nor UO_358 (O_358,N_2989,N_2953);
nor UO_359 (O_359,N_2991,N_2978);
nand UO_360 (O_360,N_2978,N_2989);
or UO_361 (O_361,N_2984,N_2939);
and UO_362 (O_362,N_2990,N_2991);
nand UO_363 (O_363,N_2993,N_2931);
and UO_364 (O_364,N_2956,N_2981);
nor UO_365 (O_365,N_2925,N_2930);
or UO_366 (O_366,N_2952,N_2993);
or UO_367 (O_367,N_2963,N_2969);
or UO_368 (O_368,N_2955,N_2974);
and UO_369 (O_369,N_2960,N_2926);
or UO_370 (O_370,N_2949,N_2953);
or UO_371 (O_371,N_2944,N_2994);
or UO_372 (O_372,N_2925,N_2965);
nor UO_373 (O_373,N_2951,N_2965);
nor UO_374 (O_374,N_2945,N_2944);
nand UO_375 (O_375,N_2953,N_2947);
nor UO_376 (O_376,N_2926,N_2961);
and UO_377 (O_377,N_2932,N_2998);
and UO_378 (O_378,N_2954,N_2931);
or UO_379 (O_379,N_2979,N_2945);
nor UO_380 (O_380,N_2986,N_2966);
nor UO_381 (O_381,N_2932,N_2968);
nor UO_382 (O_382,N_2940,N_2989);
nor UO_383 (O_383,N_2982,N_2927);
or UO_384 (O_384,N_2993,N_2950);
or UO_385 (O_385,N_2956,N_2960);
nor UO_386 (O_386,N_2940,N_2983);
or UO_387 (O_387,N_2967,N_2946);
nand UO_388 (O_388,N_2939,N_2961);
nor UO_389 (O_389,N_2987,N_2989);
and UO_390 (O_390,N_2926,N_2981);
or UO_391 (O_391,N_2986,N_2934);
and UO_392 (O_392,N_2992,N_2970);
nand UO_393 (O_393,N_2988,N_2963);
nor UO_394 (O_394,N_2989,N_2975);
and UO_395 (O_395,N_2978,N_2969);
nor UO_396 (O_396,N_2981,N_2973);
or UO_397 (O_397,N_2996,N_2982);
or UO_398 (O_398,N_2935,N_2944);
or UO_399 (O_399,N_2965,N_2973);
and UO_400 (O_400,N_2991,N_2976);
nor UO_401 (O_401,N_2940,N_2972);
nand UO_402 (O_402,N_2949,N_2993);
nand UO_403 (O_403,N_2999,N_2990);
or UO_404 (O_404,N_2969,N_2999);
or UO_405 (O_405,N_2941,N_2965);
nand UO_406 (O_406,N_2936,N_2942);
and UO_407 (O_407,N_2967,N_2929);
nand UO_408 (O_408,N_2953,N_2973);
or UO_409 (O_409,N_2965,N_2999);
or UO_410 (O_410,N_2928,N_2941);
or UO_411 (O_411,N_2978,N_2984);
or UO_412 (O_412,N_2982,N_2970);
and UO_413 (O_413,N_2993,N_2992);
nor UO_414 (O_414,N_2971,N_2925);
and UO_415 (O_415,N_2975,N_2984);
nor UO_416 (O_416,N_2965,N_2944);
and UO_417 (O_417,N_2926,N_2948);
nand UO_418 (O_418,N_2943,N_2925);
or UO_419 (O_419,N_2960,N_2951);
and UO_420 (O_420,N_2930,N_2998);
or UO_421 (O_421,N_2938,N_2969);
nand UO_422 (O_422,N_2949,N_2994);
or UO_423 (O_423,N_2952,N_2935);
nand UO_424 (O_424,N_2946,N_2984);
and UO_425 (O_425,N_2982,N_2960);
or UO_426 (O_426,N_2975,N_2956);
nand UO_427 (O_427,N_2927,N_2945);
nand UO_428 (O_428,N_2981,N_2930);
nand UO_429 (O_429,N_2947,N_2940);
and UO_430 (O_430,N_2977,N_2986);
and UO_431 (O_431,N_2988,N_2932);
nand UO_432 (O_432,N_2986,N_2946);
nand UO_433 (O_433,N_2984,N_2968);
or UO_434 (O_434,N_2950,N_2995);
nand UO_435 (O_435,N_2999,N_2948);
and UO_436 (O_436,N_2987,N_2942);
and UO_437 (O_437,N_2947,N_2951);
and UO_438 (O_438,N_2952,N_2971);
and UO_439 (O_439,N_2979,N_2943);
nor UO_440 (O_440,N_2978,N_2939);
and UO_441 (O_441,N_2955,N_2967);
nand UO_442 (O_442,N_2991,N_2925);
nor UO_443 (O_443,N_2999,N_2936);
and UO_444 (O_444,N_2927,N_2933);
and UO_445 (O_445,N_2959,N_2961);
nor UO_446 (O_446,N_2975,N_2960);
or UO_447 (O_447,N_2926,N_2952);
and UO_448 (O_448,N_2986,N_2944);
nand UO_449 (O_449,N_2931,N_2975);
and UO_450 (O_450,N_2963,N_2956);
nand UO_451 (O_451,N_2926,N_2945);
or UO_452 (O_452,N_2948,N_2951);
or UO_453 (O_453,N_2982,N_2935);
or UO_454 (O_454,N_2965,N_2939);
and UO_455 (O_455,N_2972,N_2963);
and UO_456 (O_456,N_2958,N_2925);
or UO_457 (O_457,N_2962,N_2925);
nand UO_458 (O_458,N_2936,N_2994);
and UO_459 (O_459,N_2934,N_2985);
nor UO_460 (O_460,N_2942,N_2989);
and UO_461 (O_461,N_2962,N_2974);
nor UO_462 (O_462,N_2934,N_2939);
or UO_463 (O_463,N_2978,N_2964);
and UO_464 (O_464,N_2970,N_2968);
nand UO_465 (O_465,N_2954,N_2973);
nand UO_466 (O_466,N_2948,N_2947);
nor UO_467 (O_467,N_2984,N_2963);
or UO_468 (O_468,N_2942,N_2934);
nand UO_469 (O_469,N_2969,N_2982);
nor UO_470 (O_470,N_2965,N_2972);
and UO_471 (O_471,N_2987,N_2943);
nand UO_472 (O_472,N_2973,N_2949);
nand UO_473 (O_473,N_2958,N_2976);
and UO_474 (O_474,N_2940,N_2977);
and UO_475 (O_475,N_2925,N_2939);
nand UO_476 (O_476,N_2980,N_2942);
and UO_477 (O_477,N_2931,N_2982);
xor UO_478 (O_478,N_2993,N_2945);
nor UO_479 (O_479,N_2985,N_2932);
or UO_480 (O_480,N_2958,N_2962);
or UO_481 (O_481,N_2925,N_2985);
nor UO_482 (O_482,N_2948,N_2971);
or UO_483 (O_483,N_2936,N_2966);
and UO_484 (O_484,N_2984,N_2991);
nor UO_485 (O_485,N_2981,N_2937);
or UO_486 (O_486,N_2942,N_2988);
or UO_487 (O_487,N_2988,N_2996);
nor UO_488 (O_488,N_2972,N_2962);
or UO_489 (O_489,N_2944,N_2930);
or UO_490 (O_490,N_2995,N_2978);
and UO_491 (O_491,N_2977,N_2952);
and UO_492 (O_492,N_2932,N_2977);
nand UO_493 (O_493,N_2999,N_2943);
or UO_494 (O_494,N_2996,N_2948);
and UO_495 (O_495,N_2938,N_2961);
nand UO_496 (O_496,N_2928,N_2970);
nand UO_497 (O_497,N_2930,N_2995);
and UO_498 (O_498,N_2930,N_2942);
or UO_499 (O_499,N_2970,N_2936);
endmodule