module basic_500_3000_500_4_levels_1xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_98,In_178);
and U1 (N_1,In_240,In_11);
and U2 (N_2,In_136,In_353);
nand U3 (N_3,In_358,In_313);
nor U4 (N_4,In_190,In_355);
xor U5 (N_5,In_46,In_328);
or U6 (N_6,In_309,In_182);
or U7 (N_7,In_51,In_440);
nand U8 (N_8,In_283,In_322);
and U9 (N_9,In_494,In_18);
or U10 (N_10,In_377,In_366);
nor U11 (N_11,In_157,In_67);
or U12 (N_12,In_38,In_277);
or U13 (N_13,In_387,In_122);
or U14 (N_14,In_85,In_155);
nor U15 (N_15,In_415,In_304);
nand U16 (N_16,In_274,In_249);
or U17 (N_17,In_180,In_315);
nor U18 (N_18,In_203,In_379);
nand U19 (N_19,In_497,In_158);
nand U20 (N_20,In_243,In_446);
nor U21 (N_21,In_252,In_345);
and U22 (N_22,In_334,In_204);
nand U23 (N_23,In_422,In_93);
and U24 (N_24,In_253,In_57);
or U25 (N_25,In_224,In_143);
nor U26 (N_26,In_15,In_97);
and U27 (N_27,In_34,In_110);
or U28 (N_28,In_194,In_431);
nor U29 (N_29,In_299,In_324);
nand U30 (N_30,In_295,In_221);
and U31 (N_31,In_326,In_305);
nor U32 (N_32,In_310,In_196);
or U33 (N_33,In_268,In_197);
and U34 (N_34,In_47,In_397);
and U35 (N_35,In_452,In_50);
and U36 (N_36,In_421,In_323);
nand U37 (N_37,In_73,In_453);
or U38 (N_38,In_33,In_375);
xor U39 (N_39,In_435,In_370);
nand U40 (N_40,In_43,In_383);
nor U41 (N_41,In_169,In_119);
or U42 (N_42,In_62,In_457);
and U43 (N_43,In_488,In_267);
nand U44 (N_44,In_361,In_402);
or U45 (N_45,In_76,In_20);
or U46 (N_46,In_29,In_384);
nand U47 (N_47,In_437,In_439);
and U48 (N_48,In_146,In_245);
nand U49 (N_49,In_92,In_469);
and U50 (N_50,In_430,In_137);
nand U51 (N_51,In_294,In_30);
and U52 (N_52,In_493,In_371);
or U53 (N_53,In_264,In_87);
and U54 (N_54,In_470,In_163);
or U55 (N_55,In_123,In_443);
and U56 (N_56,In_27,In_378);
or U57 (N_57,In_472,In_374);
nor U58 (N_58,In_212,In_22);
and U59 (N_59,In_399,In_392);
or U60 (N_60,In_239,In_306);
nand U61 (N_61,In_215,In_275);
and U62 (N_62,In_75,In_381);
nand U63 (N_63,In_236,In_428);
or U64 (N_64,In_247,In_201);
nor U65 (N_65,In_464,In_485);
and U66 (N_66,In_285,In_237);
nor U67 (N_67,In_71,In_346);
nand U68 (N_68,In_363,In_17);
nor U69 (N_69,In_219,In_260);
xnor U70 (N_70,In_362,In_226);
nand U71 (N_71,In_160,In_459);
nand U72 (N_72,In_386,In_466);
or U73 (N_73,In_429,In_126);
and U74 (N_74,In_96,In_26);
or U75 (N_75,In_179,In_108);
nor U76 (N_76,In_35,In_199);
nand U77 (N_77,In_52,In_241);
or U78 (N_78,In_175,In_1);
or U79 (N_79,In_10,In_231);
nor U80 (N_80,In_321,In_290);
nor U81 (N_81,In_418,In_438);
or U82 (N_82,In_13,In_32);
nand U83 (N_83,In_114,In_148);
nor U84 (N_84,In_28,In_341);
or U85 (N_85,In_282,In_495);
nand U86 (N_86,In_166,In_357);
or U87 (N_87,In_340,In_456);
nand U88 (N_88,In_468,In_273);
and U89 (N_89,In_351,In_214);
or U90 (N_90,In_106,In_188);
and U91 (N_91,In_218,In_410);
and U92 (N_92,In_380,In_484);
and U93 (N_93,In_296,In_339);
nand U94 (N_94,In_364,In_404);
nand U95 (N_95,In_481,In_40);
nand U96 (N_96,In_21,In_498);
or U97 (N_97,In_471,In_352);
nor U98 (N_98,In_4,In_293);
or U99 (N_99,In_256,In_189);
nor U100 (N_100,In_350,In_473);
and U101 (N_101,In_16,In_234);
and U102 (N_102,In_31,In_420);
or U103 (N_103,In_127,In_496);
nand U104 (N_104,In_91,In_129);
or U105 (N_105,In_69,In_263);
and U106 (N_106,In_265,In_138);
nand U107 (N_107,In_42,In_135);
or U108 (N_108,In_233,In_24);
and U109 (N_109,In_331,In_262);
nand U110 (N_110,In_90,In_45);
nand U111 (N_111,In_64,In_398);
or U112 (N_112,In_365,In_207);
nand U113 (N_113,In_60,In_349);
or U114 (N_114,In_213,In_133);
nand U115 (N_115,In_416,In_74);
nand U116 (N_116,In_112,In_205);
nand U117 (N_117,In_419,In_298);
or U118 (N_118,In_458,In_225);
and U119 (N_119,In_254,In_427);
nor U120 (N_120,In_195,In_316);
and U121 (N_121,In_44,In_217);
xor U122 (N_122,In_330,In_376);
nor U123 (N_123,In_99,In_385);
or U124 (N_124,In_132,In_107);
and U125 (N_125,In_423,In_342);
nor U126 (N_126,In_244,In_23);
nand U127 (N_127,In_144,In_159);
nor U128 (N_128,In_84,In_266);
or U129 (N_129,In_460,In_489);
and U130 (N_130,In_287,In_454);
nand U131 (N_131,In_368,In_373);
nor U132 (N_132,In_183,In_288);
nor U133 (N_133,In_156,In_72);
or U134 (N_134,In_173,In_436);
or U135 (N_135,In_449,In_68);
and U136 (N_136,In_113,In_65);
or U137 (N_137,In_327,In_396);
and U138 (N_138,In_486,In_289);
and U139 (N_139,In_425,In_367);
nor U140 (N_140,In_149,In_12);
nor U141 (N_141,In_162,In_434);
and U142 (N_142,In_147,In_280);
or U143 (N_143,In_128,In_391);
and U144 (N_144,In_0,In_115);
nand U145 (N_145,In_211,In_297);
or U146 (N_146,In_152,In_153);
and U147 (N_147,In_2,In_248);
nor U148 (N_148,In_389,In_462);
nand U149 (N_149,In_467,In_281);
or U150 (N_150,In_445,In_39);
nand U151 (N_151,In_54,In_192);
nor U152 (N_152,In_301,In_412);
or U153 (N_153,In_400,In_222);
nor U154 (N_154,In_176,In_270);
or U155 (N_155,In_82,In_455);
nand U156 (N_156,In_56,In_475);
nor U157 (N_157,In_118,In_154);
nor U158 (N_158,In_451,In_405);
and U159 (N_159,In_19,In_104);
or U160 (N_160,In_314,In_302);
nor U161 (N_161,In_272,In_48);
nor U162 (N_162,In_477,In_14);
xnor U163 (N_163,In_36,In_66);
nand U164 (N_164,In_284,In_325);
or U165 (N_165,In_77,In_450);
nor U166 (N_166,In_111,In_79);
nor U167 (N_167,In_292,In_390);
nand U168 (N_168,In_140,In_332);
nor U169 (N_169,In_177,In_480);
nor U170 (N_170,In_271,In_333);
nor U171 (N_171,In_220,In_347);
and U172 (N_172,In_441,In_409);
nor U173 (N_173,In_465,In_202);
and U174 (N_174,In_186,In_337);
and U175 (N_175,In_130,In_319);
nand U176 (N_176,In_109,In_318);
or U177 (N_177,In_250,In_417);
nor U178 (N_178,In_414,In_242);
nand U179 (N_179,In_388,In_229);
nand U180 (N_180,In_151,In_63);
or U181 (N_181,In_360,In_344);
or U182 (N_182,In_49,In_338);
and U183 (N_183,In_395,In_105);
or U184 (N_184,In_170,In_37);
xnor U185 (N_185,In_184,In_372);
or U186 (N_186,In_444,In_312);
nand U187 (N_187,In_230,In_100);
nand U188 (N_188,In_103,In_276);
or U189 (N_189,In_59,In_258);
and U190 (N_190,In_5,In_424);
nor U191 (N_191,In_235,In_139);
and U192 (N_192,In_102,In_246);
nand U193 (N_193,In_174,In_116);
nand U194 (N_194,In_145,In_131);
or U195 (N_195,In_492,In_474);
and U196 (N_196,In_279,In_70);
nand U197 (N_197,In_7,In_251);
nand U198 (N_198,In_191,In_53);
nand U199 (N_199,In_172,In_80);
nand U200 (N_200,In_78,In_483);
or U201 (N_201,In_369,In_134);
or U202 (N_202,In_257,In_426);
and U203 (N_203,In_8,In_117);
or U204 (N_204,In_165,In_300);
nand U205 (N_205,In_442,In_3);
nor U206 (N_206,In_403,In_329);
nor U207 (N_207,In_303,In_83);
nor U208 (N_208,In_150,In_89);
and U209 (N_209,In_88,In_81);
nor U210 (N_210,In_142,In_25);
nand U211 (N_211,In_359,In_406);
nand U212 (N_212,In_335,In_171);
and U213 (N_213,In_101,In_227);
nand U214 (N_214,In_187,In_286);
or U215 (N_215,In_308,In_6);
and U216 (N_216,In_478,In_141);
nor U217 (N_217,In_490,In_209);
and U218 (N_218,In_200,In_125);
nor U219 (N_219,In_121,In_413);
nor U220 (N_220,In_232,In_269);
nand U221 (N_221,In_491,In_9);
or U222 (N_222,In_476,In_185);
and U223 (N_223,In_447,In_448);
nor U224 (N_224,In_463,In_86);
nor U225 (N_225,In_261,In_317);
and U226 (N_226,In_161,In_228);
or U227 (N_227,In_487,In_482);
and U228 (N_228,In_278,In_198);
nor U229 (N_229,In_238,In_408);
and U230 (N_230,In_58,In_354);
nor U231 (N_231,In_61,In_167);
or U232 (N_232,In_164,In_168);
or U233 (N_233,In_461,In_401);
or U234 (N_234,In_216,In_291);
and U235 (N_235,In_41,In_336);
nand U236 (N_236,In_255,In_193);
and U237 (N_237,In_411,In_311);
or U238 (N_238,In_479,In_343);
and U239 (N_239,In_120,In_55);
and U240 (N_240,In_208,In_348);
or U241 (N_241,In_307,In_181);
and U242 (N_242,In_356,In_394);
and U243 (N_243,In_210,In_223);
nor U244 (N_244,In_433,In_382);
and U245 (N_245,In_206,In_95);
nand U246 (N_246,In_407,In_320);
nand U247 (N_247,In_94,In_259);
and U248 (N_248,In_393,In_432);
and U249 (N_249,In_499,In_124);
and U250 (N_250,In_174,In_251);
and U251 (N_251,In_323,In_207);
nand U252 (N_252,In_318,In_160);
or U253 (N_253,In_405,In_31);
or U254 (N_254,In_288,In_114);
nor U255 (N_255,In_65,In_46);
or U256 (N_256,In_93,In_255);
nor U257 (N_257,In_6,In_449);
nor U258 (N_258,In_69,In_43);
nand U259 (N_259,In_267,In_448);
nand U260 (N_260,In_226,In_215);
or U261 (N_261,In_458,In_83);
nand U262 (N_262,In_82,In_330);
nand U263 (N_263,In_222,In_16);
and U264 (N_264,In_91,In_432);
or U265 (N_265,In_112,In_225);
or U266 (N_266,In_112,In_53);
or U267 (N_267,In_326,In_320);
nand U268 (N_268,In_167,In_388);
and U269 (N_269,In_494,In_381);
or U270 (N_270,In_96,In_410);
and U271 (N_271,In_96,In_129);
and U272 (N_272,In_371,In_27);
or U273 (N_273,In_321,In_29);
or U274 (N_274,In_313,In_28);
and U275 (N_275,In_8,In_70);
nand U276 (N_276,In_73,In_416);
nand U277 (N_277,In_135,In_350);
nand U278 (N_278,In_313,In_181);
nand U279 (N_279,In_254,In_332);
and U280 (N_280,In_297,In_37);
nor U281 (N_281,In_220,In_231);
nand U282 (N_282,In_4,In_191);
or U283 (N_283,In_86,In_261);
nor U284 (N_284,In_167,In_72);
or U285 (N_285,In_452,In_183);
or U286 (N_286,In_4,In_57);
nor U287 (N_287,In_100,In_186);
or U288 (N_288,In_420,In_104);
and U289 (N_289,In_58,In_349);
and U290 (N_290,In_277,In_386);
or U291 (N_291,In_208,In_421);
nand U292 (N_292,In_390,In_436);
nand U293 (N_293,In_250,In_423);
and U294 (N_294,In_21,In_107);
and U295 (N_295,In_168,In_342);
nor U296 (N_296,In_40,In_384);
nor U297 (N_297,In_147,In_154);
and U298 (N_298,In_156,In_263);
nand U299 (N_299,In_453,In_373);
nor U300 (N_300,In_493,In_201);
nor U301 (N_301,In_81,In_194);
or U302 (N_302,In_170,In_262);
nor U303 (N_303,In_372,In_292);
or U304 (N_304,In_384,In_392);
nor U305 (N_305,In_228,In_33);
nor U306 (N_306,In_151,In_403);
nand U307 (N_307,In_223,In_12);
and U308 (N_308,In_305,In_489);
or U309 (N_309,In_390,In_147);
and U310 (N_310,In_73,In_430);
and U311 (N_311,In_314,In_397);
nor U312 (N_312,In_38,In_252);
nand U313 (N_313,In_130,In_5);
or U314 (N_314,In_170,In_232);
nand U315 (N_315,In_283,In_161);
nor U316 (N_316,In_292,In_351);
nand U317 (N_317,In_442,In_368);
and U318 (N_318,In_342,In_169);
nand U319 (N_319,In_51,In_354);
nor U320 (N_320,In_319,In_397);
and U321 (N_321,In_352,In_71);
nand U322 (N_322,In_457,In_418);
nor U323 (N_323,In_124,In_404);
or U324 (N_324,In_212,In_3);
and U325 (N_325,In_159,In_391);
and U326 (N_326,In_117,In_356);
or U327 (N_327,In_246,In_131);
or U328 (N_328,In_128,In_323);
nor U329 (N_329,In_170,In_226);
nor U330 (N_330,In_64,In_324);
nor U331 (N_331,In_298,In_166);
xor U332 (N_332,In_186,In_478);
xor U333 (N_333,In_107,In_313);
nand U334 (N_334,In_454,In_197);
nand U335 (N_335,In_222,In_426);
nor U336 (N_336,In_209,In_160);
nand U337 (N_337,In_358,In_55);
nor U338 (N_338,In_21,In_284);
nor U339 (N_339,In_484,In_44);
nor U340 (N_340,In_433,In_307);
and U341 (N_341,In_378,In_431);
nand U342 (N_342,In_164,In_326);
or U343 (N_343,In_161,In_446);
or U344 (N_344,In_423,In_17);
nand U345 (N_345,In_322,In_105);
and U346 (N_346,In_188,In_137);
nand U347 (N_347,In_473,In_189);
and U348 (N_348,In_286,In_151);
xor U349 (N_349,In_489,In_471);
nand U350 (N_350,In_459,In_45);
nor U351 (N_351,In_224,In_137);
and U352 (N_352,In_223,In_165);
and U353 (N_353,In_471,In_311);
nor U354 (N_354,In_160,In_327);
and U355 (N_355,In_409,In_496);
nand U356 (N_356,In_299,In_416);
or U357 (N_357,In_204,In_183);
nand U358 (N_358,In_163,In_174);
or U359 (N_359,In_398,In_182);
and U360 (N_360,In_473,In_455);
and U361 (N_361,In_22,In_173);
nand U362 (N_362,In_384,In_485);
nand U363 (N_363,In_211,In_69);
nand U364 (N_364,In_184,In_405);
or U365 (N_365,In_237,In_83);
or U366 (N_366,In_365,In_203);
nor U367 (N_367,In_462,In_55);
or U368 (N_368,In_303,In_222);
nor U369 (N_369,In_221,In_35);
or U370 (N_370,In_51,In_263);
nor U371 (N_371,In_105,In_95);
nand U372 (N_372,In_312,In_422);
and U373 (N_373,In_315,In_70);
and U374 (N_374,In_11,In_2);
or U375 (N_375,In_463,In_33);
or U376 (N_376,In_68,In_325);
nand U377 (N_377,In_131,In_265);
nand U378 (N_378,In_281,In_465);
nor U379 (N_379,In_114,In_475);
and U380 (N_380,In_36,In_444);
nand U381 (N_381,In_442,In_89);
nand U382 (N_382,In_267,In_290);
nor U383 (N_383,In_112,In_52);
nand U384 (N_384,In_351,In_291);
or U385 (N_385,In_444,In_112);
or U386 (N_386,In_283,In_121);
nand U387 (N_387,In_277,In_88);
and U388 (N_388,In_469,In_64);
nand U389 (N_389,In_469,In_483);
nand U390 (N_390,In_44,In_62);
or U391 (N_391,In_22,In_185);
and U392 (N_392,In_470,In_399);
nand U393 (N_393,In_272,In_75);
and U394 (N_394,In_36,In_233);
and U395 (N_395,In_286,In_184);
and U396 (N_396,In_268,In_420);
and U397 (N_397,In_77,In_394);
and U398 (N_398,In_234,In_252);
nand U399 (N_399,In_32,In_306);
and U400 (N_400,In_381,In_9);
nor U401 (N_401,In_448,In_145);
and U402 (N_402,In_345,In_101);
and U403 (N_403,In_353,In_441);
nor U404 (N_404,In_455,In_42);
and U405 (N_405,In_320,In_337);
xor U406 (N_406,In_355,In_0);
and U407 (N_407,In_189,In_449);
or U408 (N_408,In_353,In_17);
and U409 (N_409,In_98,In_73);
or U410 (N_410,In_0,In_37);
nor U411 (N_411,In_146,In_182);
nor U412 (N_412,In_417,In_249);
nor U413 (N_413,In_252,In_110);
or U414 (N_414,In_464,In_14);
nand U415 (N_415,In_294,In_169);
and U416 (N_416,In_203,In_121);
or U417 (N_417,In_147,In_236);
nor U418 (N_418,In_412,In_349);
nand U419 (N_419,In_339,In_434);
or U420 (N_420,In_145,In_263);
and U421 (N_421,In_78,In_193);
or U422 (N_422,In_198,In_181);
nand U423 (N_423,In_44,In_358);
and U424 (N_424,In_36,In_26);
or U425 (N_425,In_307,In_21);
nand U426 (N_426,In_133,In_231);
nor U427 (N_427,In_491,In_242);
or U428 (N_428,In_499,In_15);
nand U429 (N_429,In_499,In_250);
nand U430 (N_430,In_354,In_140);
nand U431 (N_431,In_494,In_108);
or U432 (N_432,In_12,In_254);
nor U433 (N_433,In_298,In_237);
or U434 (N_434,In_18,In_297);
nand U435 (N_435,In_351,In_289);
nor U436 (N_436,In_245,In_415);
nor U437 (N_437,In_239,In_14);
or U438 (N_438,In_486,In_98);
nand U439 (N_439,In_334,In_162);
and U440 (N_440,In_374,In_427);
nand U441 (N_441,In_431,In_261);
or U442 (N_442,In_208,In_438);
or U443 (N_443,In_282,In_455);
and U444 (N_444,In_355,In_399);
nand U445 (N_445,In_65,In_305);
and U446 (N_446,In_191,In_374);
or U447 (N_447,In_75,In_148);
nand U448 (N_448,In_453,In_333);
and U449 (N_449,In_419,In_62);
nor U450 (N_450,In_45,In_251);
nand U451 (N_451,In_363,In_286);
and U452 (N_452,In_283,In_345);
and U453 (N_453,In_42,In_438);
nand U454 (N_454,In_184,In_172);
nor U455 (N_455,In_436,In_141);
nor U456 (N_456,In_79,In_76);
or U457 (N_457,In_236,In_159);
nand U458 (N_458,In_349,In_403);
nand U459 (N_459,In_340,In_259);
or U460 (N_460,In_487,In_160);
or U461 (N_461,In_350,In_232);
nor U462 (N_462,In_122,In_389);
or U463 (N_463,In_178,In_405);
nor U464 (N_464,In_242,In_270);
nand U465 (N_465,In_322,In_94);
nor U466 (N_466,In_113,In_26);
or U467 (N_467,In_106,In_462);
and U468 (N_468,In_403,In_478);
nand U469 (N_469,In_286,In_158);
nand U470 (N_470,In_435,In_492);
and U471 (N_471,In_416,In_481);
nor U472 (N_472,In_27,In_34);
nor U473 (N_473,In_122,In_166);
nand U474 (N_474,In_237,In_491);
or U475 (N_475,In_52,In_270);
nor U476 (N_476,In_417,In_123);
and U477 (N_477,In_231,In_203);
and U478 (N_478,In_71,In_375);
or U479 (N_479,In_473,In_45);
nand U480 (N_480,In_306,In_132);
and U481 (N_481,In_97,In_187);
and U482 (N_482,In_31,In_478);
or U483 (N_483,In_213,In_425);
or U484 (N_484,In_70,In_488);
and U485 (N_485,In_226,In_151);
or U486 (N_486,In_164,In_331);
nor U487 (N_487,In_259,In_18);
or U488 (N_488,In_187,In_295);
or U489 (N_489,In_320,In_109);
or U490 (N_490,In_270,In_300);
or U491 (N_491,In_116,In_283);
or U492 (N_492,In_222,In_485);
and U493 (N_493,In_270,In_150);
nand U494 (N_494,In_117,In_101);
nor U495 (N_495,In_448,In_278);
and U496 (N_496,In_443,In_117);
nand U497 (N_497,In_411,In_105);
or U498 (N_498,In_63,In_152);
nand U499 (N_499,In_86,In_412);
or U500 (N_500,In_63,In_64);
nand U501 (N_501,In_36,In_149);
or U502 (N_502,In_167,In_189);
or U503 (N_503,In_22,In_293);
and U504 (N_504,In_401,In_497);
nor U505 (N_505,In_389,In_446);
or U506 (N_506,In_325,In_427);
and U507 (N_507,In_195,In_143);
nor U508 (N_508,In_278,In_469);
nor U509 (N_509,In_152,In_43);
xor U510 (N_510,In_230,In_154);
nand U511 (N_511,In_188,In_296);
nand U512 (N_512,In_50,In_3);
and U513 (N_513,In_184,In_496);
and U514 (N_514,In_122,In_372);
nand U515 (N_515,In_145,In_109);
nand U516 (N_516,In_474,In_320);
nor U517 (N_517,In_303,In_354);
and U518 (N_518,In_0,In_313);
nand U519 (N_519,In_190,In_217);
nand U520 (N_520,In_362,In_39);
or U521 (N_521,In_430,In_208);
nor U522 (N_522,In_10,In_234);
nand U523 (N_523,In_401,In_218);
and U524 (N_524,In_417,In_444);
nand U525 (N_525,In_387,In_212);
nor U526 (N_526,In_253,In_27);
or U527 (N_527,In_457,In_137);
nor U528 (N_528,In_396,In_282);
nor U529 (N_529,In_380,In_427);
and U530 (N_530,In_145,In_478);
nand U531 (N_531,In_474,In_358);
nor U532 (N_532,In_209,In_378);
nor U533 (N_533,In_467,In_52);
and U534 (N_534,In_89,In_485);
and U535 (N_535,In_291,In_73);
and U536 (N_536,In_340,In_75);
or U537 (N_537,In_439,In_499);
and U538 (N_538,In_66,In_443);
or U539 (N_539,In_412,In_103);
nor U540 (N_540,In_127,In_493);
nand U541 (N_541,In_195,In_315);
and U542 (N_542,In_338,In_309);
nand U543 (N_543,In_226,In_158);
and U544 (N_544,In_302,In_81);
nand U545 (N_545,In_124,In_384);
xnor U546 (N_546,In_308,In_312);
and U547 (N_547,In_332,In_94);
nor U548 (N_548,In_40,In_87);
nor U549 (N_549,In_390,In_41);
nor U550 (N_550,In_256,In_183);
or U551 (N_551,In_318,In_25);
and U552 (N_552,In_258,In_4);
nand U553 (N_553,In_160,In_290);
or U554 (N_554,In_458,In_219);
nor U555 (N_555,In_343,In_421);
nor U556 (N_556,In_416,In_380);
and U557 (N_557,In_124,In_334);
nor U558 (N_558,In_85,In_188);
or U559 (N_559,In_251,In_320);
or U560 (N_560,In_330,In_391);
nor U561 (N_561,In_442,In_113);
or U562 (N_562,In_457,In_211);
nand U563 (N_563,In_145,In_186);
nor U564 (N_564,In_169,In_429);
and U565 (N_565,In_41,In_325);
nand U566 (N_566,In_396,In_189);
nor U567 (N_567,In_42,In_264);
nor U568 (N_568,In_101,In_278);
nor U569 (N_569,In_296,In_389);
and U570 (N_570,In_442,In_104);
and U571 (N_571,In_440,In_22);
nor U572 (N_572,In_24,In_51);
and U573 (N_573,In_36,In_373);
or U574 (N_574,In_390,In_183);
and U575 (N_575,In_382,In_394);
and U576 (N_576,In_435,In_81);
and U577 (N_577,In_475,In_40);
nand U578 (N_578,In_403,In_46);
and U579 (N_579,In_218,In_443);
or U580 (N_580,In_293,In_130);
and U581 (N_581,In_317,In_262);
nand U582 (N_582,In_388,In_315);
and U583 (N_583,In_113,In_296);
and U584 (N_584,In_460,In_163);
and U585 (N_585,In_147,In_212);
or U586 (N_586,In_348,In_148);
nor U587 (N_587,In_341,In_342);
or U588 (N_588,In_240,In_155);
or U589 (N_589,In_234,In_218);
nand U590 (N_590,In_343,In_462);
and U591 (N_591,In_88,In_151);
nor U592 (N_592,In_462,In_100);
nor U593 (N_593,In_132,In_299);
nand U594 (N_594,In_86,In_71);
nor U595 (N_595,In_351,In_205);
and U596 (N_596,In_278,In_496);
nand U597 (N_597,In_35,In_266);
and U598 (N_598,In_136,In_442);
nand U599 (N_599,In_484,In_152);
nand U600 (N_600,In_404,In_345);
and U601 (N_601,In_20,In_18);
nand U602 (N_602,In_209,In_425);
or U603 (N_603,In_110,In_465);
nand U604 (N_604,In_490,In_282);
and U605 (N_605,In_73,In_76);
or U606 (N_606,In_371,In_362);
and U607 (N_607,In_178,In_390);
or U608 (N_608,In_15,In_348);
or U609 (N_609,In_82,In_281);
nor U610 (N_610,In_181,In_85);
nand U611 (N_611,In_462,In_424);
nand U612 (N_612,In_213,In_116);
nor U613 (N_613,In_415,In_478);
nor U614 (N_614,In_378,In_481);
or U615 (N_615,In_66,In_432);
nand U616 (N_616,In_332,In_454);
nor U617 (N_617,In_271,In_331);
or U618 (N_618,In_404,In_428);
or U619 (N_619,In_236,In_16);
or U620 (N_620,In_366,In_454);
or U621 (N_621,In_257,In_307);
and U622 (N_622,In_429,In_112);
or U623 (N_623,In_206,In_387);
or U624 (N_624,In_447,In_1);
or U625 (N_625,In_141,In_357);
and U626 (N_626,In_215,In_72);
nor U627 (N_627,In_411,In_267);
nor U628 (N_628,In_436,In_101);
and U629 (N_629,In_341,In_468);
and U630 (N_630,In_164,In_404);
nand U631 (N_631,In_114,In_431);
nor U632 (N_632,In_88,In_127);
nor U633 (N_633,In_284,In_179);
or U634 (N_634,In_348,In_470);
nor U635 (N_635,In_376,In_316);
and U636 (N_636,In_90,In_442);
or U637 (N_637,In_157,In_88);
or U638 (N_638,In_392,In_148);
or U639 (N_639,In_124,In_268);
nand U640 (N_640,In_116,In_361);
nand U641 (N_641,In_108,In_158);
nor U642 (N_642,In_69,In_492);
nand U643 (N_643,In_436,In_162);
nand U644 (N_644,In_358,In_170);
nor U645 (N_645,In_468,In_140);
nand U646 (N_646,In_138,In_177);
and U647 (N_647,In_11,In_408);
nor U648 (N_648,In_368,In_471);
nor U649 (N_649,In_429,In_6);
nor U650 (N_650,In_326,In_301);
or U651 (N_651,In_229,In_375);
nor U652 (N_652,In_279,In_392);
and U653 (N_653,In_410,In_489);
and U654 (N_654,In_382,In_116);
and U655 (N_655,In_409,In_262);
or U656 (N_656,In_77,In_1);
nand U657 (N_657,In_298,In_346);
nand U658 (N_658,In_123,In_465);
or U659 (N_659,In_408,In_147);
nor U660 (N_660,In_93,In_130);
or U661 (N_661,In_287,In_177);
nand U662 (N_662,In_13,In_320);
and U663 (N_663,In_463,In_331);
or U664 (N_664,In_425,In_260);
nor U665 (N_665,In_401,In_206);
nand U666 (N_666,In_216,In_177);
nand U667 (N_667,In_352,In_212);
or U668 (N_668,In_62,In_208);
nor U669 (N_669,In_58,In_128);
and U670 (N_670,In_253,In_2);
nand U671 (N_671,In_214,In_357);
nor U672 (N_672,In_274,In_484);
nor U673 (N_673,In_491,In_351);
and U674 (N_674,In_477,In_221);
and U675 (N_675,In_202,In_219);
and U676 (N_676,In_353,In_472);
nor U677 (N_677,In_72,In_319);
or U678 (N_678,In_65,In_304);
nand U679 (N_679,In_9,In_424);
or U680 (N_680,In_106,In_418);
and U681 (N_681,In_396,In_240);
nor U682 (N_682,In_276,In_429);
nor U683 (N_683,In_59,In_228);
or U684 (N_684,In_251,In_337);
nor U685 (N_685,In_72,In_345);
nand U686 (N_686,In_297,In_218);
nor U687 (N_687,In_498,In_144);
nand U688 (N_688,In_277,In_167);
or U689 (N_689,In_295,In_78);
nand U690 (N_690,In_427,In_27);
nor U691 (N_691,In_35,In_71);
or U692 (N_692,In_397,In_274);
nand U693 (N_693,In_269,In_318);
or U694 (N_694,In_439,In_132);
nor U695 (N_695,In_468,In_324);
or U696 (N_696,In_18,In_95);
nor U697 (N_697,In_348,In_299);
nor U698 (N_698,In_290,In_52);
nor U699 (N_699,In_274,In_340);
nand U700 (N_700,In_176,In_37);
nor U701 (N_701,In_345,In_11);
nor U702 (N_702,In_397,In_235);
nand U703 (N_703,In_252,In_480);
nor U704 (N_704,In_115,In_264);
nand U705 (N_705,In_446,In_181);
nor U706 (N_706,In_148,In_367);
nor U707 (N_707,In_140,In_69);
nand U708 (N_708,In_452,In_317);
nor U709 (N_709,In_30,In_222);
and U710 (N_710,In_195,In_3);
nor U711 (N_711,In_333,In_338);
or U712 (N_712,In_4,In_319);
nor U713 (N_713,In_395,In_44);
nand U714 (N_714,In_174,In_50);
and U715 (N_715,In_125,In_426);
nor U716 (N_716,In_268,In_151);
nor U717 (N_717,In_174,In_275);
nor U718 (N_718,In_226,In_445);
or U719 (N_719,In_336,In_203);
nor U720 (N_720,In_196,In_120);
and U721 (N_721,In_36,In_195);
nand U722 (N_722,In_436,In_461);
and U723 (N_723,In_408,In_383);
nand U724 (N_724,In_387,In_396);
or U725 (N_725,In_394,In_239);
and U726 (N_726,In_19,In_191);
nor U727 (N_727,In_140,In_185);
nor U728 (N_728,In_116,In_262);
nor U729 (N_729,In_499,In_134);
or U730 (N_730,In_462,In_282);
and U731 (N_731,In_301,In_203);
nand U732 (N_732,In_10,In_421);
or U733 (N_733,In_153,In_126);
or U734 (N_734,In_335,In_74);
or U735 (N_735,In_375,In_263);
nor U736 (N_736,In_17,In_493);
and U737 (N_737,In_276,In_3);
nand U738 (N_738,In_107,In_391);
xnor U739 (N_739,In_83,In_130);
nand U740 (N_740,In_272,In_330);
and U741 (N_741,In_319,In_470);
or U742 (N_742,In_3,In_68);
nor U743 (N_743,In_31,In_168);
or U744 (N_744,In_122,In_286);
and U745 (N_745,In_337,In_446);
nand U746 (N_746,In_57,In_410);
nand U747 (N_747,In_251,In_393);
nor U748 (N_748,In_187,In_244);
nor U749 (N_749,In_57,In_300);
nand U750 (N_750,N_456,N_575);
and U751 (N_751,N_26,N_21);
and U752 (N_752,N_682,N_547);
and U753 (N_753,N_233,N_182);
nor U754 (N_754,N_330,N_548);
or U755 (N_755,N_122,N_302);
nand U756 (N_756,N_345,N_157);
nor U757 (N_757,N_156,N_129);
or U758 (N_758,N_99,N_334);
nand U759 (N_759,N_744,N_535);
or U760 (N_760,N_662,N_183);
nor U761 (N_761,N_400,N_430);
nand U762 (N_762,N_423,N_609);
nand U763 (N_763,N_489,N_304);
and U764 (N_764,N_488,N_161);
and U765 (N_765,N_222,N_17);
nand U766 (N_766,N_601,N_331);
and U767 (N_767,N_446,N_409);
nand U768 (N_768,N_251,N_205);
nor U769 (N_769,N_697,N_214);
nor U770 (N_770,N_235,N_621);
or U771 (N_771,N_185,N_283);
and U772 (N_772,N_80,N_518);
nor U773 (N_773,N_350,N_741);
nor U774 (N_774,N_337,N_309);
or U775 (N_775,N_594,N_420);
nand U776 (N_776,N_730,N_435);
nand U777 (N_777,N_438,N_390);
nor U778 (N_778,N_708,N_629);
and U779 (N_779,N_33,N_7);
nand U780 (N_780,N_516,N_713);
nand U781 (N_781,N_360,N_363);
or U782 (N_782,N_656,N_478);
nor U783 (N_783,N_323,N_606);
or U784 (N_784,N_32,N_612);
nor U785 (N_785,N_212,N_449);
or U786 (N_786,N_76,N_696);
and U787 (N_787,N_325,N_492);
and U788 (N_788,N_568,N_515);
and U789 (N_789,N_496,N_630);
or U790 (N_790,N_148,N_109);
and U791 (N_791,N_270,N_69);
or U792 (N_792,N_211,N_158);
nand U793 (N_793,N_253,N_24);
or U794 (N_794,N_747,N_711);
and U795 (N_795,N_570,N_471);
xnor U796 (N_796,N_495,N_514);
and U797 (N_797,N_19,N_201);
or U798 (N_798,N_8,N_746);
or U799 (N_799,N_396,N_406);
and U800 (N_800,N_167,N_491);
nand U801 (N_801,N_57,N_384);
or U802 (N_802,N_417,N_245);
nand U803 (N_803,N_125,N_128);
and U804 (N_804,N_447,N_155);
and U805 (N_805,N_184,N_395);
and U806 (N_806,N_87,N_88);
and U807 (N_807,N_85,N_126);
or U808 (N_808,N_580,N_78);
nand U809 (N_809,N_238,N_241);
nor U810 (N_810,N_313,N_482);
nand U811 (N_811,N_610,N_294);
or U812 (N_812,N_694,N_149);
nor U813 (N_813,N_307,N_101);
nand U814 (N_814,N_346,N_692);
or U815 (N_815,N_4,N_550);
and U816 (N_816,N_297,N_506);
nor U817 (N_817,N_246,N_415);
or U818 (N_818,N_588,N_733);
and U819 (N_819,N_494,N_722);
nand U820 (N_820,N_193,N_555);
and U821 (N_821,N_450,N_532);
or U822 (N_822,N_187,N_1);
and U823 (N_823,N_68,N_596);
and U824 (N_824,N_95,N_45);
and U825 (N_825,N_476,N_521);
nor U826 (N_826,N_587,N_186);
or U827 (N_827,N_401,N_604);
and U828 (N_828,N_107,N_70);
nor U829 (N_829,N_556,N_481);
nor U830 (N_830,N_546,N_265);
or U831 (N_831,N_725,N_279);
and U832 (N_832,N_82,N_36);
nor U833 (N_833,N_705,N_695);
and U834 (N_834,N_90,N_105);
nor U835 (N_835,N_675,N_392);
nor U836 (N_836,N_616,N_94);
xnor U837 (N_837,N_732,N_252);
nand U838 (N_838,N_273,N_67);
nand U839 (N_839,N_698,N_584);
and U840 (N_840,N_457,N_333);
or U841 (N_841,N_40,N_593);
and U842 (N_842,N_727,N_370);
xor U843 (N_843,N_343,N_527);
and U844 (N_844,N_573,N_227);
or U845 (N_845,N_592,N_239);
or U846 (N_846,N_267,N_305);
and U847 (N_847,N_154,N_232);
nor U848 (N_848,N_354,N_531);
or U849 (N_849,N_719,N_647);
and U850 (N_850,N_320,N_269);
nand U851 (N_851,N_665,N_544);
nor U852 (N_852,N_586,N_284);
nand U853 (N_853,N_631,N_364);
nor U854 (N_854,N_502,N_558);
nor U855 (N_855,N_91,N_206);
nor U856 (N_856,N_106,N_344);
nand U857 (N_857,N_534,N_500);
and U858 (N_858,N_391,N_723);
and U859 (N_859,N_42,N_221);
nor U860 (N_860,N_191,N_683);
nand U861 (N_861,N_649,N_605);
nand U862 (N_862,N_460,N_164);
nor U863 (N_863,N_411,N_542);
nor U864 (N_864,N_275,N_266);
and U865 (N_865,N_299,N_296);
nor U866 (N_866,N_321,N_208);
and U867 (N_867,N_380,N_552);
or U868 (N_868,N_387,N_639);
and U869 (N_869,N_180,N_120);
and U870 (N_870,N_615,N_560);
nand U871 (N_871,N_30,N_640);
nor U872 (N_872,N_194,N_685);
nand U873 (N_873,N_369,N_318);
nor U874 (N_874,N_285,N_503);
or U875 (N_875,N_618,N_557);
or U876 (N_876,N_614,N_3);
or U877 (N_877,N_608,N_229);
or U878 (N_878,N_54,N_18);
nand U879 (N_879,N_43,N_452);
or U880 (N_880,N_382,N_104);
nor U881 (N_881,N_591,N_475);
or U882 (N_882,N_398,N_172);
nor U883 (N_883,N_427,N_748);
and U884 (N_884,N_490,N_376);
nor U885 (N_885,N_336,N_731);
nand U886 (N_886,N_429,N_451);
or U887 (N_887,N_530,N_600);
nand U888 (N_888,N_687,N_293);
or U889 (N_889,N_673,N_228);
or U890 (N_890,N_59,N_113);
and U891 (N_891,N_721,N_645);
xor U892 (N_892,N_700,N_611);
or U893 (N_893,N_300,N_140);
nor U894 (N_894,N_543,N_152);
and U895 (N_895,N_338,N_52);
or U896 (N_896,N_165,N_485);
or U897 (N_897,N_571,N_634);
nand U898 (N_898,N_133,N_301);
or U899 (N_899,N_2,N_466);
nand U900 (N_900,N_714,N_422);
or U901 (N_901,N_419,N_706);
nor U902 (N_902,N_536,N_327);
and U903 (N_903,N_402,N_539);
and U904 (N_904,N_204,N_443);
and U905 (N_905,N_486,N_190);
or U906 (N_906,N_358,N_249);
nand U907 (N_907,N_159,N_198);
nor U908 (N_908,N_513,N_432);
nor U909 (N_909,N_144,N_264);
and U910 (N_910,N_12,N_493);
and U911 (N_911,N_375,N_63);
nor U912 (N_912,N_329,N_220);
or U913 (N_913,N_386,N_244);
nor U914 (N_914,N_572,N_339);
or U915 (N_915,N_335,N_234);
nor U916 (N_916,N_124,N_366);
and U917 (N_917,N_463,N_703);
or U918 (N_918,N_373,N_315);
or U919 (N_919,N_507,N_114);
nand U920 (N_920,N_707,N_13);
and U921 (N_921,N_311,N_385);
xor U922 (N_922,N_35,N_174);
and U923 (N_923,N_347,N_117);
or U924 (N_924,N_738,N_579);
nand U925 (N_925,N_407,N_434);
nand U926 (N_926,N_661,N_316);
nand U927 (N_927,N_210,N_465);
and U928 (N_928,N_110,N_112);
and U929 (N_929,N_431,N_589);
nor U930 (N_930,N_559,N_178);
nor U931 (N_931,N_497,N_28);
nand U932 (N_932,N_209,N_218);
nor U933 (N_933,N_520,N_540);
nor U934 (N_934,N_393,N_508);
nor U935 (N_935,N_288,N_453);
xor U936 (N_936,N_278,N_84);
and U937 (N_937,N_282,N_720);
or U938 (N_938,N_16,N_260);
nand U939 (N_939,N_620,N_561);
nor U940 (N_940,N_403,N_365);
or U941 (N_941,N_501,N_53);
and U942 (N_942,N_525,N_710);
nand U943 (N_943,N_247,N_574);
nand U944 (N_944,N_290,N_567);
and U945 (N_945,N_439,N_121);
and U946 (N_946,N_65,N_74);
and U947 (N_947,N_213,N_276);
and U948 (N_948,N_308,N_268);
and U949 (N_949,N_664,N_135);
or U950 (N_950,N_134,N_170);
and U951 (N_951,N_348,N_289);
and U952 (N_952,N_189,N_29);
nand U953 (N_953,N_734,N_192);
or U954 (N_954,N_286,N_168);
nand U955 (N_955,N_92,N_641);
and U956 (N_956,N_404,N_737);
or U957 (N_957,N_689,N_340);
nand U958 (N_958,N_97,N_619);
nand U959 (N_959,N_468,N_145);
nor U960 (N_960,N_740,N_326);
or U961 (N_961,N_188,N_81);
nor U962 (N_962,N_702,N_693);
or U963 (N_963,N_440,N_71);
nor U964 (N_964,N_569,N_14);
and U965 (N_965,N_736,N_562);
xor U966 (N_966,N_196,N_362);
nand U967 (N_967,N_444,N_357);
nand U968 (N_968,N_424,N_622);
nor U969 (N_969,N_426,N_642);
and U970 (N_970,N_676,N_324);
nand U971 (N_971,N_62,N_226);
and U972 (N_972,N_653,N_116);
nand U973 (N_973,N_96,N_724);
or U974 (N_974,N_72,N_50);
nor U975 (N_975,N_255,N_9);
nand U976 (N_976,N_287,N_668);
or U977 (N_977,N_578,N_277);
or U978 (N_978,N_55,N_138);
nand U979 (N_979,N_652,N_577);
nand U980 (N_980,N_372,N_549);
and U981 (N_981,N_469,N_153);
or U982 (N_982,N_735,N_509);
or U983 (N_983,N_351,N_272);
nor U984 (N_984,N_51,N_510);
and U985 (N_985,N_505,N_659);
nand U986 (N_986,N_413,N_669);
nand U987 (N_987,N_627,N_623);
nor U988 (N_988,N_678,N_261);
or U989 (N_989,N_442,N_371);
nor U990 (N_990,N_565,N_139);
or U991 (N_991,N_256,N_31);
nor U992 (N_992,N_0,N_648);
or U993 (N_993,N_64,N_655);
or U994 (N_994,N_312,N_202);
and U995 (N_995,N_684,N_225);
nor U996 (N_996,N_504,N_461);
nor U997 (N_997,N_617,N_314);
or U998 (N_998,N_271,N_136);
nor U999 (N_999,N_717,N_729);
nand U1000 (N_1000,N_250,N_243);
nor U1001 (N_1001,N_10,N_203);
and U1002 (N_1002,N_454,N_131);
nor U1003 (N_1003,N_254,N_89);
nand U1004 (N_1004,N_526,N_353);
or U1005 (N_1005,N_437,N_46);
nor U1006 (N_1006,N_119,N_742);
nor U1007 (N_1007,N_433,N_58);
or U1008 (N_1008,N_47,N_34);
or U1009 (N_1009,N_484,N_699);
nand U1010 (N_1010,N_644,N_75);
nor U1011 (N_1011,N_108,N_436);
nor U1012 (N_1012,N_576,N_499);
and U1013 (N_1013,N_650,N_718);
and U1014 (N_1014,N_378,N_38);
and U1015 (N_1015,N_118,N_595);
nor U1016 (N_1016,N_498,N_200);
nand U1017 (N_1017,N_541,N_607);
nor U1018 (N_1018,N_77,N_688);
nand U1019 (N_1019,N_690,N_394);
nor U1020 (N_1020,N_230,N_459);
nand U1021 (N_1021,N_73,N_162);
nor U1022 (N_1022,N_679,N_712);
or U1023 (N_1023,N_680,N_11);
nand U1024 (N_1024,N_551,N_361);
or U1025 (N_1025,N_425,N_739);
nor U1026 (N_1026,N_632,N_480);
nand U1027 (N_1027,N_666,N_428);
or U1028 (N_1028,N_533,N_445);
or U1029 (N_1029,N_473,N_356);
and U1030 (N_1030,N_716,N_298);
and U1031 (N_1031,N_237,N_635);
or U1032 (N_1032,N_581,N_472);
nand U1033 (N_1033,N_388,N_412);
or U1034 (N_1034,N_553,N_389);
or U1035 (N_1035,N_538,N_274);
or U1036 (N_1036,N_474,N_585);
nand U1037 (N_1037,N_414,N_657);
and U1038 (N_1038,N_654,N_671);
nor U1039 (N_1039,N_519,N_704);
or U1040 (N_1040,N_150,N_217);
and U1041 (N_1041,N_637,N_399);
and U1042 (N_1042,N_280,N_524);
and U1043 (N_1043,N_599,N_60);
or U1044 (N_1044,N_410,N_236);
or U1045 (N_1045,N_563,N_691);
nand U1046 (N_1046,N_745,N_179);
nand U1047 (N_1047,N_102,N_670);
nand U1048 (N_1048,N_219,N_686);
or U1049 (N_1049,N_160,N_242);
or U1050 (N_1050,N_147,N_728);
nor U1051 (N_1051,N_146,N_352);
or U1052 (N_1052,N_663,N_259);
and U1053 (N_1053,N_467,N_175);
and U1054 (N_1054,N_177,N_332);
and U1055 (N_1055,N_15,N_636);
and U1056 (N_1056,N_651,N_529);
nor U1057 (N_1057,N_523,N_416);
nor U1058 (N_1058,N_625,N_528);
nand U1059 (N_1059,N_743,N_660);
or U1060 (N_1060,N_674,N_626);
nand U1061 (N_1061,N_281,N_143);
or U1062 (N_1062,N_405,N_22);
nor U1063 (N_1063,N_583,N_726);
nand U1064 (N_1064,N_643,N_263);
xor U1065 (N_1065,N_56,N_141);
or U1066 (N_1066,N_418,N_537);
and U1067 (N_1067,N_83,N_132);
and U1068 (N_1068,N_127,N_381);
nand U1069 (N_1069,N_582,N_441);
and U1070 (N_1070,N_166,N_672);
nor U1071 (N_1071,N_216,N_100);
nor U1072 (N_1072,N_566,N_715);
or U1073 (N_1073,N_368,N_163);
nor U1074 (N_1074,N_590,N_341);
nor U1075 (N_1075,N_199,N_319);
nand U1076 (N_1076,N_483,N_455);
nand U1077 (N_1077,N_598,N_39);
or U1078 (N_1078,N_262,N_6);
nor U1079 (N_1079,N_130,N_27);
nand U1080 (N_1080,N_115,N_367);
and U1081 (N_1081,N_379,N_240);
and U1082 (N_1082,N_171,N_303);
nand U1083 (N_1083,N_41,N_421);
nand U1084 (N_1084,N_310,N_61);
or U1085 (N_1085,N_383,N_342);
nand U1086 (N_1086,N_458,N_554);
and U1087 (N_1087,N_477,N_224);
or U1088 (N_1088,N_464,N_111);
nor U1089 (N_1089,N_295,N_677);
nor U1090 (N_1090,N_374,N_597);
and U1091 (N_1091,N_377,N_646);
nand U1092 (N_1092,N_667,N_98);
or U1093 (N_1093,N_151,N_603);
and U1094 (N_1094,N_355,N_223);
and U1095 (N_1095,N_44,N_602);
and U1096 (N_1096,N_215,N_169);
or U1097 (N_1097,N_462,N_49);
and U1098 (N_1098,N_633,N_79);
nor U1099 (N_1099,N_397,N_5);
or U1100 (N_1100,N_195,N_470);
nand U1101 (N_1101,N_628,N_142);
and U1102 (N_1102,N_197,N_176);
nor U1103 (N_1103,N_487,N_317);
and U1104 (N_1104,N_701,N_207);
and U1105 (N_1105,N_292,N_613);
nand U1106 (N_1106,N_48,N_103);
or U1107 (N_1107,N_23,N_749);
and U1108 (N_1108,N_258,N_512);
nand U1109 (N_1109,N_173,N_349);
nor U1110 (N_1110,N_248,N_231);
and U1111 (N_1111,N_479,N_291);
or U1112 (N_1112,N_322,N_37);
or U1113 (N_1113,N_257,N_20);
or U1114 (N_1114,N_328,N_137);
nand U1115 (N_1115,N_448,N_86);
and U1116 (N_1116,N_638,N_123);
nand U1117 (N_1117,N_709,N_564);
nand U1118 (N_1118,N_681,N_306);
or U1119 (N_1119,N_658,N_624);
or U1120 (N_1120,N_93,N_517);
nor U1121 (N_1121,N_408,N_66);
and U1122 (N_1122,N_522,N_359);
nand U1123 (N_1123,N_545,N_511);
or U1124 (N_1124,N_25,N_181);
nand U1125 (N_1125,N_700,N_277);
or U1126 (N_1126,N_38,N_736);
or U1127 (N_1127,N_299,N_160);
nor U1128 (N_1128,N_698,N_146);
or U1129 (N_1129,N_171,N_379);
nand U1130 (N_1130,N_85,N_48);
and U1131 (N_1131,N_553,N_618);
or U1132 (N_1132,N_132,N_98);
and U1133 (N_1133,N_112,N_34);
nor U1134 (N_1134,N_136,N_127);
nand U1135 (N_1135,N_412,N_12);
or U1136 (N_1136,N_236,N_152);
and U1137 (N_1137,N_46,N_638);
nand U1138 (N_1138,N_263,N_87);
nand U1139 (N_1139,N_392,N_419);
nand U1140 (N_1140,N_236,N_719);
xor U1141 (N_1141,N_491,N_498);
xor U1142 (N_1142,N_99,N_336);
and U1143 (N_1143,N_584,N_530);
nand U1144 (N_1144,N_481,N_68);
and U1145 (N_1145,N_275,N_81);
and U1146 (N_1146,N_96,N_652);
or U1147 (N_1147,N_181,N_29);
and U1148 (N_1148,N_410,N_146);
or U1149 (N_1149,N_484,N_727);
or U1150 (N_1150,N_655,N_182);
nor U1151 (N_1151,N_143,N_608);
nand U1152 (N_1152,N_720,N_335);
nand U1153 (N_1153,N_522,N_624);
nor U1154 (N_1154,N_625,N_194);
or U1155 (N_1155,N_71,N_20);
nor U1156 (N_1156,N_664,N_586);
or U1157 (N_1157,N_90,N_610);
or U1158 (N_1158,N_663,N_84);
and U1159 (N_1159,N_173,N_738);
or U1160 (N_1160,N_733,N_362);
nand U1161 (N_1161,N_266,N_713);
nor U1162 (N_1162,N_553,N_65);
and U1163 (N_1163,N_668,N_540);
nand U1164 (N_1164,N_497,N_103);
nand U1165 (N_1165,N_220,N_482);
nand U1166 (N_1166,N_306,N_204);
or U1167 (N_1167,N_526,N_189);
and U1168 (N_1168,N_556,N_723);
and U1169 (N_1169,N_125,N_568);
nand U1170 (N_1170,N_126,N_36);
xnor U1171 (N_1171,N_289,N_601);
or U1172 (N_1172,N_1,N_698);
and U1173 (N_1173,N_519,N_213);
nand U1174 (N_1174,N_738,N_361);
and U1175 (N_1175,N_579,N_309);
or U1176 (N_1176,N_85,N_228);
nand U1177 (N_1177,N_533,N_382);
nand U1178 (N_1178,N_591,N_316);
or U1179 (N_1179,N_666,N_374);
or U1180 (N_1180,N_231,N_14);
nand U1181 (N_1181,N_572,N_562);
nand U1182 (N_1182,N_210,N_40);
nand U1183 (N_1183,N_437,N_2);
nand U1184 (N_1184,N_201,N_226);
and U1185 (N_1185,N_204,N_626);
and U1186 (N_1186,N_554,N_192);
and U1187 (N_1187,N_70,N_463);
nor U1188 (N_1188,N_3,N_514);
or U1189 (N_1189,N_95,N_421);
nand U1190 (N_1190,N_634,N_393);
or U1191 (N_1191,N_314,N_425);
nor U1192 (N_1192,N_291,N_193);
nand U1193 (N_1193,N_736,N_307);
nor U1194 (N_1194,N_318,N_484);
nand U1195 (N_1195,N_105,N_687);
nand U1196 (N_1196,N_252,N_334);
nor U1197 (N_1197,N_319,N_382);
nand U1198 (N_1198,N_643,N_341);
nor U1199 (N_1199,N_540,N_379);
and U1200 (N_1200,N_435,N_21);
or U1201 (N_1201,N_267,N_486);
and U1202 (N_1202,N_620,N_87);
nor U1203 (N_1203,N_433,N_108);
or U1204 (N_1204,N_499,N_391);
or U1205 (N_1205,N_522,N_702);
nand U1206 (N_1206,N_581,N_590);
xnor U1207 (N_1207,N_692,N_696);
nor U1208 (N_1208,N_37,N_401);
nor U1209 (N_1209,N_677,N_348);
or U1210 (N_1210,N_316,N_689);
or U1211 (N_1211,N_201,N_116);
and U1212 (N_1212,N_412,N_628);
or U1213 (N_1213,N_512,N_132);
or U1214 (N_1214,N_98,N_595);
and U1215 (N_1215,N_605,N_691);
or U1216 (N_1216,N_408,N_301);
nand U1217 (N_1217,N_299,N_36);
nor U1218 (N_1218,N_57,N_190);
or U1219 (N_1219,N_137,N_559);
nand U1220 (N_1220,N_273,N_207);
nand U1221 (N_1221,N_412,N_109);
nor U1222 (N_1222,N_250,N_586);
xor U1223 (N_1223,N_294,N_489);
nor U1224 (N_1224,N_277,N_616);
nor U1225 (N_1225,N_669,N_432);
or U1226 (N_1226,N_59,N_748);
or U1227 (N_1227,N_297,N_91);
nand U1228 (N_1228,N_478,N_116);
nor U1229 (N_1229,N_445,N_543);
nand U1230 (N_1230,N_320,N_574);
or U1231 (N_1231,N_596,N_26);
nand U1232 (N_1232,N_458,N_164);
nand U1233 (N_1233,N_169,N_699);
and U1234 (N_1234,N_208,N_436);
nor U1235 (N_1235,N_674,N_305);
and U1236 (N_1236,N_587,N_385);
and U1237 (N_1237,N_506,N_507);
and U1238 (N_1238,N_652,N_52);
or U1239 (N_1239,N_177,N_20);
nor U1240 (N_1240,N_116,N_509);
or U1241 (N_1241,N_211,N_530);
nand U1242 (N_1242,N_15,N_595);
nand U1243 (N_1243,N_8,N_430);
or U1244 (N_1244,N_105,N_735);
and U1245 (N_1245,N_681,N_575);
nor U1246 (N_1246,N_640,N_485);
or U1247 (N_1247,N_61,N_363);
and U1248 (N_1248,N_321,N_603);
nand U1249 (N_1249,N_114,N_514);
nand U1250 (N_1250,N_313,N_90);
or U1251 (N_1251,N_167,N_186);
nor U1252 (N_1252,N_452,N_427);
nor U1253 (N_1253,N_14,N_103);
nor U1254 (N_1254,N_539,N_525);
and U1255 (N_1255,N_149,N_519);
nor U1256 (N_1256,N_118,N_422);
nand U1257 (N_1257,N_703,N_462);
nand U1258 (N_1258,N_252,N_165);
nand U1259 (N_1259,N_229,N_159);
or U1260 (N_1260,N_130,N_274);
and U1261 (N_1261,N_23,N_91);
nor U1262 (N_1262,N_687,N_605);
nor U1263 (N_1263,N_133,N_396);
or U1264 (N_1264,N_629,N_475);
nor U1265 (N_1265,N_726,N_318);
and U1266 (N_1266,N_697,N_123);
or U1267 (N_1267,N_728,N_592);
nand U1268 (N_1268,N_243,N_266);
nand U1269 (N_1269,N_622,N_209);
and U1270 (N_1270,N_673,N_508);
and U1271 (N_1271,N_534,N_75);
or U1272 (N_1272,N_246,N_575);
nand U1273 (N_1273,N_186,N_238);
nor U1274 (N_1274,N_142,N_26);
and U1275 (N_1275,N_704,N_732);
and U1276 (N_1276,N_738,N_158);
xnor U1277 (N_1277,N_286,N_705);
nor U1278 (N_1278,N_37,N_314);
nand U1279 (N_1279,N_299,N_308);
or U1280 (N_1280,N_279,N_334);
or U1281 (N_1281,N_399,N_33);
nand U1282 (N_1282,N_536,N_434);
nor U1283 (N_1283,N_585,N_45);
nor U1284 (N_1284,N_105,N_559);
and U1285 (N_1285,N_436,N_491);
xnor U1286 (N_1286,N_677,N_60);
or U1287 (N_1287,N_304,N_743);
nor U1288 (N_1288,N_401,N_115);
or U1289 (N_1289,N_704,N_457);
nand U1290 (N_1290,N_322,N_489);
and U1291 (N_1291,N_408,N_414);
or U1292 (N_1292,N_696,N_222);
nand U1293 (N_1293,N_305,N_298);
nand U1294 (N_1294,N_203,N_472);
nand U1295 (N_1295,N_319,N_738);
or U1296 (N_1296,N_399,N_496);
or U1297 (N_1297,N_653,N_705);
or U1298 (N_1298,N_133,N_669);
nand U1299 (N_1299,N_477,N_597);
or U1300 (N_1300,N_334,N_372);
nor U1301 (N_1301,N_428,N_390);
and U1302 (N_1302,N_548,N_466);
nor U1303 (N_1303,N_743,N_541);
and U1304 (N_1304,N_47,N_115);
nor U1305 (N_1305,N_131,N_518);
nand U1306 (N_1306,N_627,N_294);
nor U1307 (N_1307,N_295,N_43);
or U1308 (N_1308,N_327,N_521);
nand U1309 (N_1309,N_642,N_562);
or U1310 (N_1310,N_592,N_191);
or U1311 (N_1311,N_140,N_55);
and U1312 (N_1312,N_218,N_353);
and U1313 (N_1313,N_292,N_428);
nand U1314 (N_1314,N_115,N_16);
nand U1315 (N_1315,N_415,N_419);
nor U1316 (N_1316,N_747,N_17);
nand U1317 (N_1317,N_102,N_744);
or U1318 (N_1318,N_611,N_638);
and U1319 (N_1319,N_128,N_426);
and U1320 (N_1320,N_379,N_504);
nand U1321 (N_1321,N_310,N_264);
nor U1322 (N_1322,N_48,N_385);
nand U1323 (N_1323,N_663,N_680);
nand U1324 (N_1324,N_621,N_233);
nor U1325 (N_1325,N_369,N_62);
nand U1326 (N_1326,N_119,N_428);
nor U1327 (N_1327,N_196,N_228);
or U1328 (N_1328,N_101,N_125);
xor U1329 (N_1329,N_657,N_279);
nor U1330 (N_1330,N_178,N_63);
nand U1331 (N_1331,N_338,N_533);
nand U1332 (N_1332,N_459,N_369);
nor U1333 (N_1333,N_688,N_582);
nand U1334 (N_1334,N_725,N_292);
or U1335 (N_1335,N_18,N_111);
and U1336 (N_1336,N_702,N_184);
nor U1337 (N_1337,N_128,N_277);
or U1338 (N_1338,N_34,N_443);
nor U1339 (N_1339,N_421,N_82);
and U1340 (N_1340,N_571,N_585);
xnor U1341 (N_1341,N_130,N_433);
nand U1342 (N_1342,N_532,N_589);
nor U1343 (N_1343,N_412,N_182);
nand U1344 (N_1344,N_704,N_469);
or U1345 (N_1345,N_667,N_334);
nor U1346 (N_1346,N_652,N_547);
or U1347 (N_1347,N_399,N_657);
and U1348 (N_1348,N_369,N_656);
nand U1349 (N_1349,N_585,N_570);
nand U1350 (N_1350,N_277,N_33);
and U1351 (N_1351,N_356,N_634);
nor U1352 (N_1352,N_121,N_519);
nand U1353 (N_1353,N_481,N_54);
nor U1354 (N_1354,N_346,N_24);
or U1355 (N_1355,N_293,N_536);
or U1356 (N_1356,N_722,N_747);
or U1357 (N_1357,N_79,N_510);
or U1358 (N_1358,N_507,N_450);
and U1359 (N_1359,N_362,N_393);
nor U1360 (N_1360,N_71,N_583);
nor U1361 (N_1361,N_603,N_696);
and U1362 (N_1362,N_57,N_722);
or U1363 (N_1363,N_465,N_677);
or U1364 (N_1364,N_4,N_393);
xnor U1365 (N_1365,N_91,N_694);
nor U1366 (N_1366,N_604,N_93);
or U1367 (N_1367,N_675,N_342);
nand U1368 (N_1368,N_404,N_422);
or U1369 (N_1369,N_645,N_622);
or U1370 (N_1370,N_494,N_707);
and U1371 (N_1371,N_19,N_539);
nor U1372 (N_1372,N_649,N_234);
nand U1373 (N_1373,N_544,N_590);
or U1374 (N_1374,N_652,N_390);
nand U1375 (N_1375,N_212,N_13);
nor U1376 (N_1376,N_560,N_663);
or U1377 (N_1377,N_243,N_737);
nand U1378 (N_1378,N_342,N_264);
nand U1379 (N_1379,N_449,N_96);
or U1380 (N_1380,N_76,N_176);
nor U1381 (N_1381,N_479,N_353);
nand U1382 (N_1382,N_104,N_586);
or U1383 (N_1383,N_193,N_413);
nor U1384 (N_1384,N_579,N_495);
nand U1385 (N_1385,N_705,N_307);
nor U1386 (N_1386,N_670,N_219);
and U1387 (N_1387,N_216,N_260);
and U1388 (N_1388,N_177,N_229);
or U1389 (N_1389,N_462,N_587);
nor U1390 (N_1390,N_608,N_49);
and U1391 (N_1391,N_72,N_423);
and U1392 (N_1392,N_673,N_244);
or U1393 (N_1393,N_158,N_604);
or U1394 (N_1394,N_351,N_407);
nand U1395 (N_1395,N_420,N_432);
or U1396 (N_1396,N_156,N_630);
and U1397 (N_1397,N_336,N_183);
nand U1398 (N_1398,N_656,N_339);
and U1399 (N_1399,N_438,N_285);
nand U1400 (N_1400,N_322,N_48);
nand U1401 (N_1401,N_598,N_442);
or U1402 (N_1402,N_456,N_585);
or U1403 (N_1403,N_640,N_399);
nor U1404 (N_1404,N_746,N_391);
nor U1405 (N_1405,N_240,N_165);
and U1406 (N_1406,N_69,N_646);
and U1407 (N_1407,N_679,N_69);
nand U1408 (N_1408,N_330,N_46);
nand U1409 (N_1409,N_647,N_141);
nand U1410 (N_1410,N_274,N_197);
or U1411 (N_1411,N_367,N_24);
and U1412 (N_1412,N_642,N_390);
nor U1413 (N_1413,N_453,N_734);
xnor U1414 (N_1414,N_368,N_559);
nor U1415 (N_1415,N_247,N_387);
and U1416 (N_1416,N_175,N_676);
nor U1417 (N_1417,N_622,N_201);
nor U1418 (N_1418,N_401,N_17);
and U1419 (N_1419,N_111,N_707);
nand U1420 (N_1420,N_314,N_245);
nor U1421 (N_1421,N_289,N_386);
and U1422 (N_1422,N_280,N_424);
or U1423 (N_1423,N_101,N_29);
nor U1424 (N_1424,N_190,N_558);
nor U1425 (N_1425,N_397,N_393);
or U1426 (N_1426,N_305,N_434);
or U1427 (N_1427,N_412,N_491);
nand U1428 (N_1428,N_226,N_547);
nor U1429 (N_1429,N_370,N_498);
or U1430 (N_1430,N_183,N_579);
nand U1431 (N_1431,N_660,N_670);
nor U1432 (N_1432,N_60,N_195);
or U1433 (N_1433,N_531,N_429);
and U1434 (N_1434,N_499,N_91);
nor U1435 (N_1435,N_279,N_479);
or U1436 (N_1436,N_164,N_448);
and U1437 (N_1437,N_465,N_290);
and U1438 (N_1438,N_622,N_569);
nand U1439 (N_1439,N_622,N_367);
or U1440 (N_1440,N_579,N_518);
nor U1441 (N_1441,N_233,N_639);
nor U1442 (N_1442,N_257,N_85);
or U1443 (N_1443,N_674,N_533);
nor U1444 (N_1444,N_743,N_6);
nand U1445 (N_1445,N_131,N_255);
and U1446 (N_1446,N_516,N_335);
nor U1447 (N_1447,N_634,N_611);
nand U1448 (N_1448,N_368,N_83);
or U1449 (N_1449,N_746,N_144);
nor U1450 (N_1450,N_681,N_440);
or U1451 (N_1451,N_636,N_118);
and U1452 (N_1452,N_376,N_341);
nor U1453 (N_1453,N_712,N_39);
and U1454 (N_1454,N_384,N_634);
xnor U1455 (N_1455,N_434,N_249);
nand U1456 (N_1456,N_324,N_68);
nand U1457 (N_1457,N_414,N_688);
nand U1458 (N_1458,N_160,N_8);
and U1459 (N_1459,N_143,N_506);
nor U1460 (N_1460,N_6,N_117);
nand U1461 (N_1461,N_18,N_236);
nor U1462 (N_1462,N_45,N_506);
and U1463 (N_1463,N_518,N_526);
and U1464 (N_1464,N_320,N_232);
nor U1465 (N_1465,N_524,N_732);
and U1466 (N_1466,N_360,N_563);
nor U1467 (N_1467,N_442,N_570);
or U1468 (N_1468,N_290,N_56);
and U1469 (N_1469,N_319,N_673);
nor U1470 (N_1470,N_50,N_225);
or U1471 (N_1471,N_83,N_713);
xnor U1472 (N_1472,N_124,N_387);
xnor U1473 (N_1473,N_335,N_703);
nand U1474 (N_1474,N_651,N_121);
and U1475 (N_1475,N_362,N_123);
or U1476 (N_1476,N_716,N_190);
and U1477 (N_1477,N_410,N_618);
or U1478 (N_1478,N_557,N_519);
and U1479 (N_1479,N_137,N_234);
or U1480 (N_1480,N_678,N_42);
and U1481 (N_1481,N_137,N_546);
or U1482 (N_1482,N_286,N_502);
nand U1483 (N_1483,N_35,N_369);
or U1484 (N_1484,N_85,N_469);
and U1485 (N_1485,N_175,N_141);
and U1486 (N_1486,N_15,N_582);
or U1487 (N_1487,N_105,N_638);
and U1488 (N_1488,N_146,N_107);
or U1489 (N_1489,N_590,N_671);
or U1490 (N_1490,N_521,N_185);
or U1491 (N_1491,N_66,N_669);
or U1492 (N_1492,N_292,N_599);
nor U1493 (N_1493,N_582,N_555);
and U1494 (N_1494,N_652,N_206);
nand U1495 (N_1495,N_492,N_360);
nand U1496 (N_1496,N_677,N_27);
or U1497 (N_1497,N_176,N_604);
nand U1498 (N_1498,N_713,N_163);
nor U1499 (N_1499,N_42,N_106);
and U1500 (N_1500,N_853,N_1290);
nor U1501 (N_1501,N_1115,N_1236);
and U1502 (N_1502,N_1409,N_940);
or U1503 (N_1503,N_843,N_1403);
or U1504 (N_1504,N_1338,N_1034);
nand U1505 (N_1505,N_763,N_1367);
and U1506 (N_1506,N_1159,N_960);
and U1507 (N_1507,N_1248,N_1330);
nand U1508 (N_1508,N_1176,N_1272);
xor U1509 (N_1509,N_1323,N_1013);
nand U1510 (N_1510,N_954,N_1015);
and U1511 (N_1511,N_1244,N_1499);
xnor U1512 (N_1512,N_1360,N_1215);
or U1513 (N_1513,N_1408,N_1472);
and U1514 (N_1514,N_975,N_1405);
nor U1515 (N_1515,N_1186,N_1037);
nand U1516 (N_1516,N_1304,N_1436);
nor U1517 (N_1517,N_1368,N_1026);
nor U1518 (N_1518,N_1250,N_1233);
nand U1519 (N_1519,N_958,N_1181);
and U1520 (N_1520,N_1120,N_1006);
and U1521 (N_1521,N_1318,N_1163);
and U1522 (N_1522,N_1161,N_1375);
nand U1523 (N_1523,N_1298,N_1058);
nand U1524 (N_1524,N_1162,N_1216);
nor U1525 (N_1525,N_1397,N_849);
nor U1526 (N_1526,N_895,N_977);
nor U1527 (N_1527,N_1157,N_1112);
nor U1528 (N_1528,N_987,N_1458);
and U1529 (N_1529,N_1343,N_1035);
nor U1530 (N_1530,N_1200,N_1346);
or U1531 (N_1531,N_1363,N_781);
or U1532 (N_1532,N_850,N_1302);
nor U1533 (N_1533,N_817,N_1427);
nor U1534 (N_1534,N_1421,N_896);
or U1535 (N_1535,N_1151,N_756);
or U1536 (N_1536,N_1340,N_868);
or U1537 (N_1537,N_1428,N_1023);
and U1538 (N_1538,N_761,N_859);
or U1539 (N_1539,N_770,N_1217);
or U1540 (N_1540,N_950,N_1412);
nand U1541 (N_1541,N_797,N_886);
nor U1542 (N_1542,N_912,N_1169);
or U1543 (N_1543,N_905,N_762);
nor U1544 (N_1544,N_1135,N_996);
and U1545 (N_1545,N_1099,N_1122);
and U1546 (N_1546,N_885,N_786);
or U1547 (N_1547,N_1180,N_1241);
nand U1548 (N_1548,N_931,N_1148);
and U1549 (N_1549,N_1048,N_1075);
nand U1550 (N_1550,N_796,N_1106);
nand U1551 (N_1551,N_959,N_1275);
and U1552 (N_1552,N_1324,N_1240);
nor U1553 (N_1553,N_785,N_1086);
or U1554 (N_1554,N_754,N_1390);
and U1555 (N_1555,N_910,N_932);
or U1556 (N_1556,N_1172,N_1049);
and U1557 (N_1557,N_1213,N_1413);
nand U1558 (N_1558,N_1349,N_858);
nand U1559 (N_1559,N_1105,N_1144);
nor U1560 (N_1560,N_783,N_1039);
and U1561 (N_1561,N_1132,N_986);
nor U1562 (N_1562,N_840,N_1296);
nand U1563 (N_1563,N_1482,N_1104);
nor U1564 (N_1564,N_1228,N_1150);
nand U1565 (N_1565,N_1025,N_953);
nand U1566 (N_1566,N_1263,N_802);
and U1567 (N_1567,N_1459,N_1155);
nor U1568 (N_1568,N_1154,N_1254);
nand U1569 (N_1569,N_1022,N_1443);
nor U1570 (N_1570,N_1067,N_1014);
and U1571 (N_1571,N_1358,N_823);
nand U1572 (N_1572,N_983,N_1071);
nand U1573 (N_1573,N_1005,N_945);
nand U1574 (N_1574,N_1266,N_1429);
or U1575 (N_1575,N_946,N_1449);
nor U1576 (N_1576,N_1407,N_1274);
nand U1577 (N_1577,N_1052,N_964);
nor U1578 (N_1578,N_1268,N_978);
nand U1579 (N_1579,N_1383,N_1111);
nor U1580 (N_1580,N_1237,N_933);
nand U1581 (N_1581,N_1088,N_1433);
nand U1582 (N_1582,N_1199,N_821);
and U1583 (N_1583,N_1187,N_790);
or U1584 (N_1584,N_966,N_911);
nand U1585 (N_1585,N_1220,N_1142);
and U1586 (N_1586,N_877,N_1294);
nand U1587 (N_1587,N_962,N_1095);
nor U1588 (N_1588,N_1242,N_798);
or U1589 (N_1589,N_956,N_913);
and U1590 (N_1590,N_1072,N_1195);
or U1591 (N_1591,N_1327,N_1471);
nand U1592 (N_1592,N_982,N_1446);
or U1593 (N_1593,N_1083,N_1271);
or U1594 (N_1594,N_750,N_916);
or U1595 (N_1595,N_961,N_863);
nor U1596 (N_1596,N_1175,N_1054);
nor U1597 (N_1597,N_1129,N_1207);
or U1598 (N_1598,N_1357,N_1295);
nor U1599 (N_1599,N_1369,N_1399);
or U1600 (N_1600,N_908,N_759);
nor U1601 (N_1601,N_1125,N_872);
nor U1602 (N_1602,N_1189,N_1017);
nand U1603 (N_1603,N_1314,N_1174);
nor U1604 (N_1604,N_880,N_856);
nor U1605 (N_1605,N_1091,N_865);
and U1606 (N_1606,N_1377,N_1146);
or U1607 (N_1607,N_1425,N_1422);
nand U1608 (N_1608,N_1431,N_819);
nand U1609 (N_1609,N_909,N_1253);
nor U1610 (N_1610,N_775,N_963);
nor U1611 (N_1611,N_1096,N_1040);
xnor U1612 (N_1612,N_999,N_1496);
or U1613 (N_1613,N_902,N_936);
nand U1614 (N_1614,N_918,N_887);
or U1615 (N_1615,N_1158,N_1166);
or U1616 (N_1616,N_1074,N_1098);
and U1617 (N_1617,N_1444,N_794);
nand U1618 (N_1618,N_891,N_1398);
nand U1619 (N_1619,N_1029,N_1388);
nand U1620 (N_1620,N_1464,N_884);
nor U1621 (N_1621,N_1445,N_1261);
nand U1622 (N_1622,N_1251,N_1401);
nand U1623 (N_1623,N_989,N_1093);
nor U1624 (N_1624,N_1453,N_1494);
nand U1625 (N_1625,N_1103,N_1460);
nand U1626 (N_1626,N_969,N_1381);
and U1627 (N_1627,N_1416,N_813);
and U1628 (N_1628,N_947,N_1009);
nand U1629 (N_1629,N_1497,N_791);
nor U1630 (N_1630,N_1243,N_917);
and U1631 (N_1631,N_1454,N_1130);
or U1632 (N_1632,N_1140,N_1073);
nor U1633 (N_1633,N_1069,N_792);
and U1634 (N_1634,N_1010,N_997);
nand U1635 (N_1635,N_1117,N_772);
nor U1636 (N_1636,N_1041,N_1003);
and U1637 (N_1637,N_1031,N_1209);
nor U1638 (N_1638,N_1059,N_1267);
nor U1639 (N_1639,N_1487,N_1430);
nor U1640 (N_1640,N_1042,N_1448);
nor U1641 (N_1641,N_1177,N_767);
or U1642 (N_1642,N_1418,N_1400);
or U1643 (N_1643,N_1178,N_1288);
nor U1644 (N_1644,N_1291,N_1197);
or U1645 (N_1645,N_1223,N_1102);
or U1646 (N_1646,N_1203,N_1057);
nand U1647 (N_1647,N_1179,N_1018);
and U1648 (N_1648,N_780,N_1019);
and U1649 (N_1649,N_938,N_1404);
or U1650 (N_1650,N_1372,N_1204);
nor U1651 (N_1651,N_822,N_1109);
nor U1652 (N_1652,N_893,N_1392);
and U1653 (N_1653,N_1456,N_1475);
nand U1654 (N_1654,N_1118,N_846);
or U1655 (N_1655,N_1050,N_952);
or U1656 (N_1656,N_829,N_1366);
nor U1657 (N_1657,N_806,N_970);
nor U1658 (N_1658,N_837,N_758);
and U1659 (N_1659,N_1246,N_1045);
or U1660 (N_1660,N_1373,N_1007);
nand U1661 (N_1661,N_1085,N_1447);
and U1662 (N_1662,N_1114,N_1247);
nand U1663 (N_1663,N_839,N_1333);
nor U1664 (N_1664,N_1477,N_1198);
and U1665 (N_1665,N_1047,N_1352);
nor U1666 (N_1666,N_1440,N_1476);
nand U1667 (N_1667,N_1310,N_1024);
nor U1668 (N_1668,N_1082,N_1226);
and U1669 (N_1669,N_1299,N_922);
or U1670 (N_1670,N_991,N_1355);
nand U1671 (N_1671,N_1011,N_883);
nor U1672 (N_1672,N_984,N_1402);
nand U1673 (N_1673,N_1347,N_1001);
or U1674 (N_1674,N_1080,N_787);
and U1675 (N_1675,N_873,N_1280);
and U1676 (N_1676,N_1252,N_805);
or U1677 (N_1677,N_972,N_1386);
and U1678 (N_1678,N_1384,N_1002);
and U1679 (N_1679,N_824,N_779);
and U1680 (N_1680,N_1234,N_948);
nor U1681 (N_1681,N_1451,N_773);
or U1682 (N_1682,N_890,N_1332);
xor U1683 (N_1683,N_1311,N_1258);
and U1684 (N_1684,N_1235,N_942);
nor U1685 (N_1685,N_1124,N_1256);
nand U1686 (N_1686,N_1379,N_1165);
and U1687 (N_1687,N_860,N_1345);
nand U1688 (N_1688,N_1364,N_924);
and U1689 (N_1689,N_760,N_937);
nor U1690 (N_1690,N_1190,N_921);
nand U1691 (N_1691,N_1113,N_1393);
and U1692 (N_1692,N_1264,N_1208);
nor U1693 (N_1693,N_1322,N_930);
and U1694 (N_1694,N_1171,N_919);
nor U1695 (N_1695,N_1193,N_814);
nor U1696 (N_1696,N_1287,N_1182);
nand U1697 (N_1697,N_1336,N_1339);
or U1698 (N_1698,N_1479,N_1119);
nor U1699 (N_1699,N_1297,N_981);
and U1700 (N_1700,N_965,N_751);
nor U1701 (N_1701,N_1167,N_998);
or U1702 (N_1702,N_1206,N_1374);
or U1703 (N_1703,N_1143,N_799);
or U1704 (N_1704,N_808,N_1141);
nand U1705 (N_1705,N_1492,N_1282);
or U1706 (N_1706,N_776,N_1305);
or U1707 (N_1707,N_1152,N_826);
and U1708 (N_1708,N_1465,N_1222);
nand U1709 (N_1709,N_995,N_855);
nor U1710 (N_1710,N_1205,N_1016);
nand U1711 (N_1711,N_955,N_875);
nor U1712 (N_1712,N_1452,N_1278);
nand U1713 (N_1713,N_1480,N_1262);
nor U1714 (N_1714,N_1283,N_1396);
or U1715 (N_1715,N_985,N_1110);
nand U1716 (N_1716,N_1321,N_920);
nand U1717 (N_1717,N_769,N_828);
nor U1718 (N_1718,N_793,N_1128);
or U1719 (N_1719,N_845,N_1238);
nand U1720 (N_1720,N_1123,N_755);
and U1721 (N_1721,N_753,N_818);
or U1722 (N_1722,N_1079,N_1438);
nor U1723 (N_1723,N_1210,N_1131);
or U1724 (N_1724,N_1481,N_1435);
nand U1725 (N_1725,N_1326,N_1457);
or U1726 (N_1726,N_1353,N_1108);
nand U1727 (N_1727,N_1101,N_1196);
and U1728 (N_1728,N_1328,N_1491);
or U1729 (N_1729,N_1391,N_838);
nand U1730 (N_1730,N_1489,N_899);
nand U1731 (N_1731,N_1008,N_804);
and U1732 (N_1732,N_892,N_934);
and U1733 (N_1733,N_968,N_1212);
or U1734 (N_1734,N_980,N_1051);
or U1735 (N_1735,N_1076,N_1420);
and U1736 (N_1736,N_1473,N_1331);
nand U1737 (N_1737,N_1063,N_1192);
nor U1738 (N_1738,N_789,N_1012);
or U1739 (N_1739,N_1044,N_1320);
nor U1740 (N_1740,N_834,N_1149);
nor U1741 (N_1741,N_1419,N_854);
and U1742 (N_1742,N_1214,N_1317);
or U1743 (N_1743,N_1309,N_1257);
nand U1744 (N_1744,N_795,N_825);
nand U1745 (N_1745,N_1329,N_994);
nor U1746 (N_1746,N_1153,N_1084);
nand U1747 (N_1747,N_803,N_1273);
nand U1748 (N_1748,N_1313,N_1227);
and U1749 (N_1749,N_778,N_992);
nand U1750 (N_1750,N_862,N_1365);
nor U1751 (N_1751,N_784,N_1260);
and U1752 (N_1752,N_1188,N_1070);
nand U1753 (N_1753,N_1450,N_976);
or U1754 (N_1754,N_1232,N_766);
nand U1755 (N_1755,N_1078,N_1276);
or U1756 (N_1756,N_1437,N_1134);
nor U1757 (N_1757,N_1032,N_1285);
nor U1758 (N_1758,N_851,N_807);
nand U1759 (N_1759,N_842,N_1033);
or U1760 (N_1760,N_1127,N_1249);
or U1761 (N_1761,N_1133,N_1356);
and U1762 (N_1762,N_1376,N_871);
and U1763 (N_1763,N_1173,N_852);
nand U1764 (N_1764,N_1087,N_861);
and U1765 (N_1765,N_1462,N_801);
or U1766 (N_1766,N_988,N_1387);
and U1767 (N_1767,N_974,N_1020);
or U1768 (N_1768,N_1004,N_1493);
nand U1769 (N_1769,N_810,N_941);
and U1770 (N_1770,N_1255,N_1469);
and U1771 (N_1771,N_1036,N_882);
nand U1772 (N_1772,N_990,N_1461);
nand U1773 (N_1773,N_898,N_1194);
or U1774 (N_1774,N_1308,N_1414);
or U1775 (N_1775,N_1265,N_777);
nor U1776 (N_1776,N_1303,N_1350);
nand U1777 (N_1777,N_876,N_866);
and U1778 (N_1778,N_1139,N_1277);
nor U1779 (N_1779,N_904,N_1474);
or U1780 (N_1780,N_1498,N_1092);
or U1781 (N_1781,N_757,N_811);
and U1782 (N_1782,N_1245,N_881);
and U1783 (N_1783,N_1354,N_1359);
and U1784 (N_1784,N_1466,N_1486);
and U1785 (N_1785,N_894,N_830);
xor U1786 (N_1786,N_1426,N_879);
and U1787 (N_1787,N_1239,N_1056);
and U1788 (N_1788,N_1292,N_1286);
or U1789 (N_1789,N_1337,N_1306);
or U1790 (N_1790,N_1219,N_1455);
nand U1791 (N_1791,N_1185,N_993);
and U1792 (N_1792,N_809,N_820);
and U1793 (N_1793,N_889,N_1344);
and U1794 (N_1794,N_836,N_923);
and U1795 (N_1795,N_833,N_1341);
or U1796 (N_1796,N_815,N_1053);
nand U1797 (N_1797,N_870,N_1319);
or U1798 (N_1798,N_816,N_1370);
nand U1799 (N_1799,N_1293,N_1065);
and U1800 (N_1800,N_788,N_1230);
nand U1801 (N_1801,N_1046,N_1423);
nand U1802 (N_1802,N_928,N_1062);
or U1803 (N_1803,N_752,N_939);
or U1804 (N_1804,N_1229,N_1485);
or U1805 (N_1805,N_848,N_1385);
or U1806 (N_1806,N_1028,N_1279);
xnor U1807 (N_1807,N_1470,N_1147);
nand U1808 (N_1808,N_1417,N_1406);
or U1809 (N_1809,N_1439,N_927);
nor U1810 (N_1810,N_935,N_914);
and U1811 (N_1811,N_1378,N_1441);
nand U1812 (N_1812,N_1055,N_1170);
nor U1813 (N_1813,N_764,N_1027);
nand U1814 (N_1814,N_973,N_1424);
or U1815 (N_1815,N_1289,N_1410);
nand U1816 (N_1816,N_906,N_841);
and U1817 (N_1817,N_897,N_1183);
nor U1818 (N_1818,N_1259,N_857);
or U1819 (N_1819,N_1389,N_901);
and U1820 (N_1820,N_832,N_1312);
and U1821 (N_1821,N_957,N_1468);
nand U1822 (N_1822,N_771,N_925);
or U1823 (N_1823,N_1021,N_1483);
or U1824 (N_1824,N_1081,N_1371);
nor U1825 (N_1825,N_903,N_1066);
nand U1826 (N_1826,N_1201,N_782);
nand U1827 (N_1827,N_951,N_1488);
and U1828 (N_1828,N_1030,N_1038);
and U1829 (N_1829,N_827,N_1316);
nor U1830 (N_1830,N_1463,N_1484);
nor U1831 (N_1831,N_1335,N_1467);
nand U1832 (N_1832,N_765,N_1184);
or U1833 (N_1833,N_1315,N_900);
or U1834 (N_1834,N_1168,N_1351);
nand U1835 (N_1835,N_1334,N_1043);
nand U1836 (N_1836,N_1218,N_1432);
or U1837 (N_1837,N_874,N_1090);
xor U1838 (N_1838,N_1307,N_1270);
nand U1839 (N_1839,N_1068,N_800);
or U1840 (N_1840,N_1089,N_1225);
nand U1841 (N_1841,N_1284,N_979);
nor U1842 (N_1842,N_1121,N_943);
and U1843 (N_1843,N_1136,N_774);
and U1844 (N_1844,N_1301,N_864);
or U1845 (N_1845,N_1362,N_1160);
nor U1846 (N_1846,N_1211,N_1382);
nor U1847 (N_1847,N_967,N_1221);
nor U1848 (N_1848,N_847,N_1478);
and U1849 (N_1849,N_1490,N_1164);
and U1850 (N_1850,N_915,N_835);
or U1851 (N_1851,N_1000,N_1060);
and U1852 (N_1852,N_1094,N_1231);
and U1853 (N_1853,N_1061,N_1137);
nand U1854 (N_1854,N_1442,N_1415);
nor U1855 (N_1855,N_1380,N_1097);
and U1856 (N_1856,N_1224,N_1342);
nand U1857 (N_1857,N_768,N_1202);
or U1858 (N_1858,N_1495,N_1100);
or U1859 (N_1859,N_888,N_929);
nand U1860 (N_1860,N_1411,N_831);
nand U1861 (N_1861,N_812,N_878);
or U1862 (N_1862,N_1156,N_1191);
and U1863 (N_1863,N_1281,N_1138);
and U1864 (N_1864,N_926,N_971);
nand U1865 (N_1865,N_1434,N_1361);
and U1866 (N_1866,N_1348,N_1064);
nand U1867 (N_1867,N_1077,N_907);
nand U1868 (N_1868,N_1269,N_1116);
or U1869 (N_1869,N_949,N_1325);
or U1870 (N_1870,N_867,N_1395);
nor U1871 (N_1871,N_869,N_1300);
nand U1872 (N_1872,N_1145,N_1126);
or U1873 (N_1873,N_944,N_1394);
nand U1874 (N_1874,N_1107,N_844);
nor U1875 (N_1875,N_995,N_1393);
nand U1876 (N_1876,N_981,N_841);
nand U1877 (N_1877,N_1440,N_980);
or U1878 (N_1878,N_935,N_1223);
and U1879 (N_1879,N_1063,N_849);
and U1880 (N_1880,N_1077,N_822);
nor U1881 (N_1881,N_1365,N_1245);
and U1882 (N_1882,N_1225,N_1136);
and U1883 (N_1883,N_1037,N_1148);
and U1884 (N_1884,N_1353,N_1349);
and U1885 (N_1885,N_957,N_754);
or U1886 (N_1886,N_1290,N_1190);
or U1887 (N_1887,N_1374,N_758);
nor U1888 (N_1888,N_1126,N_1280);
nor U1889 (N_1889,N_969,N_1265);
and U1890 (N_1890,N_1022,N_1318);
nand U1891 (N_1891,N_1110,N_1174);
nor U1892 (N_1892,N_1237,N_914);
xnor U1893 (N_1893,N_1482,N_1313);
and U1894 (N_1894,N_825,N_1290);
nor U1895 (N_1895,N_1066,N_1446);
nor U1896 (N_1896,N_1344,N_868);
or U1897 (N_1897,N_1382,N_1463);
nor U1898 (N_1898,N_1193,N_1270);
nor U1899 (N_1899,N_806,N_1268);
or U1900 (N_1900,N_852,N_1179);
or U1901 (N_1901,N_890,N_1129);
or U1902 (N_1902,N_1468,N_1243);
nand U1903 (N_1903,N_895,N_1027);
and U1904 (N_1904,N_1284,N_1180);
nand U1905 (N_1905,N_864,N_813);
nand U1906 (N_1906,N_1085,N_835);
or U1907 (N_1907,N_1130,N_970);
nand U1908 (N_1908,N_1371,N_810);
nand U1909 (N_1909,N_1405,N_971);
and U1910 (N_1910,N_886,N_964);
or U1911 (N_1911,N_1103,N_1194);
nor U1912 (N_1912,N_829,N_1107);
nand U1913 (N_1913,N_1337,N_1324);
and U1914 (N_1914,N_1311,N_863);
nand U1915 (N_1915,N_1147,N_1233);
nand U1916 (N_1916,N_1181,N_804);
nor U1917 (N_1917,N_1475,N_1211);
and U1918 (N_1918,N_1070,N_754);
nor U1919 (N_1919,N_767,N_1450);
and U1920 (N_1920,N_1233,N_1430);
or U1921 (N_1921,N_776,N_1498);
nand U1922 (N_1922,N_1143,N_1413);
nor U1923 (N_1923,N_1143,N_1455);
and U1924 (N_1924,N_1222,N_1397);
and U1925 (N_1925,N_1135,N_1383);
nand U1926 (N_1926,N_963,N_1284);
nand U1927 (N_1927,N_1424,N_1164);
nand U1928 (N_1928,N_986,N_1035);
and U1929 (N_1929,N_1023,N_1392);
nand U1930 (N_1930,N_1332,N_1030);
nand U1931 (N_1931,N_1190,N_1282);
nand U1932 (N_1932,N_860,N_766);
nor U1933 (N_1933,N_1363,N_1044);
nand U1934 (N_1934,N_956,N_1200);
nor U1935 (N_1935,N_1053,N_790);
and U1936 (N_1936,N_926,N_1059);
nand U1937 (N_1937,N_1432,N_841);
or U1938 (N_1938,N_872,N_1005);
nand U1939 (N_1939,N_1238,N_784);
nor U1940 (N_1940,N_814,N_1323);
and U1941 (N_1941,N_751,N_1239);
and U1942 (N_1942,N_1178,N_1109);
nand U1943 (N_1943,N_1015,N_1275);
nor U1944 (N_1944,N_964,N_1088);
nor U1945 (N_1945,N_1282,N_1017);
nand U1946 (N_1946,N_1055,N_1200);
nor U1947 (N_1947,N_1093,N_1117);
nand U1948 (N_1948,N_834,N_1002);
nand U1949 (N_1949,N_782,N_1442);
nor U1950 (N_1950,N_1039,N_1030);
nor U1951 (N_1951,N_1193,N_875);
xnor U1952 (N_1952,N_1384,N_1000);
nor U1953 (N_1953,N_795,N_1202);
and U1954 (N_1954,N_1066,N_1327);
xnor U1955 (N_1955,N_1413,N_1117);
or U1956 (N_1956,N_1189,N_1366);
and U1957 (N_1957,N_1211,N_1194);
nor U1958 (N_1958,N_1430,N_1106);
or U1959 (N_1959,N_824,N_952);
or U1960 (N_1960,N_1251,N_1313);
or U1961 (N_1961,N_1343,N_986);
or U1962 (N_1962,N_1338,N_1092);
and U1963 (N_1963,N_1303,N_956);
or U1964 (N_1964,N_892,N_1138);
nand U1965 (N_1965,N_1466,N_969);
nor U1966 (N_1966,N_1282,N_948);
nor U1967 (N_1967,N_1179,N_1159);
and U1968 (N_1968,N_840,N_1445);
nor U1969 (N_1969,N_781,N_1282);
nor U1970 (N_1970,N_1228,N_812);
nor U1971 (N_1971,N_954,N_877);
or U1972 (N_1972,N_816,N_1059);
nor U1973 (N_1973,N_872,N_1251);
and U1974 (N_1974,N_991,N_1456);
or U1975 (N_1975,N_1198,N_1011);
nand U1976 (N_1976,N_1430,N_957);
or U1977 (N_1977,N_1235,N_1242);
nand U1978 (N_1978,N_1262,N_1462);
and U1979 (N_1979,N_1225,N_1470);
nor U1980 (N_1980,N_752,N_846);
nor U1981 (N_1981,N_1252,N_1111);
nand U1982 (N_1982,N_1447,N_1471);
nor U1983 (N_1983,N_1118,N_1226);
or U1984 (N_1984,N_1295,N_1400);
nor U1985 (N_1985,N_1215,N_1474);
or U1986 (N_1986,N_840,N_1223);
nand U1987 (N_1987,N_1024,N_754);
or U1988 (N_1988,N_814,N_1313);
nand U1989 (N_1989,N_1124,N_1248);
nand U1990 (N_1990,N_1231,N_1132);
nor U1991 (N_1991,N_781,N_1221);
and U1992 (N_1992,N_1226,N_879);
or U1993 (N_1993,N_1208,N_947);
nor U1994 (N_1994,N_1270,N_967);
nor U1995 (N_1995,N_1035,N_768);
nand U1996 (N_1996,N_1417,N_1211);
nand U1997 (N_1997,N_1311,N_1445);
nor U1998 (N_1998,N_1108,N_908);
nand U1999 (N_1999,N_1402,N_1457);
nand U2000 (N_2000,N_897,N_1436);
nor U2001 (N_2001,N_925,N_757);
and U2002 (N_2002,N_1103,N_954);
or U2003 (N_2003,N_765,N_1255);
nor U2004 (N_2004,N_820,N_1051);
nor U2005 (N_2005,N_1124,N_933);
and U2006 (N_2006,N_803,N_1487);
nand U2007 (N_2007,N_1030,N_1059);
nor U2008 (N_2008,N_1320,N_996);
and U2009 (N_2009,N_1406,N_944);
or U2010 (N_2010,N_1059,N_1350);
nand U2011 (N_2011,N_1216,N_1083);
and U2012 (N_2012,N_785,N_961);
or U2013 (N_2013,N_1132,N_1430);
or U2014 (N_2014,N_1223,N_1491);
nand U2015 (N_2015,N_892,N_1089);
nor U2016 (N_2016,N_835,N_1143);
xor U2017 (N_2017,N_1015,N_1345);
or U2018 (N_2018,N_1231,N_1328);
or U2019 (N_2019,N_1229,N_1140);
and U2020 (N_2020,N_1353,N_1249);
and U2021 (N_2021,N_1265,N_1369);
nand U2022 (N_2022,N_1343,N_1400);
and U2023 (N_2023,N_1070,N_804);
or U2024 (N_2024,N_841,N_1458);
and U2025 (N_2025,N_1185,N_868);
nand U2026 (N_2026,N_1158,N_840);
or U2027 (N_2027,N_1066,N_1185);
nand U2028 (N_2028,N_902,N_929);
nand U2029 (N_2029,N_894,N_1477);
and U2030 (N_2030,N_963,N_1039);
or U2031 (N_2031,N_1372,N_1474);
and U2032 (N_2032,N_1277,N_958);
or U2033 (N_2033,N_983,N_1299);
or U2034 (N_2034,N_1313,N_882);
nand U2035 (N_2035,N_1128,N_1455);
and U2036 (N_2036,N_1238,N_1220);
nand U2037 (N_2037,N_1452,N_1009);
nand U2038 (N_2038,N_1432,N_1197);
or U2039 (N_2039,N_1364,N_1276);
nor U2040 (N_2040,N_870,N_1469);
nand U2041 (N_2041,N_1198,N_929);
nor U2042 (N_2042,N_1349,N_971);
or U2043 (N_2043,N_966,N_1359);
or U2044 (N_2044,N_1044,N_1337);
and U2045 (N_2045,N_1007,N_1302);
nand U2046 (N_2046,N_947,N_1297);
and U2047 (N_2047,N_863,N_829);
and U2048 (N_2048,N_1475,N_1075);
or U2049 (N_2049,N_1207,N_1009);
xnor U2050 (N_2050,N_914,N_1418);
nand U2051 (N_2051,N_1438,N_1499);
or U2052 (N_2052,N_1029,N_991);
nor U2053 (N_2053,N_1144,N_973);
and U2054 (N_2054,N_766,N_1145);
xor U2055 (N_2055,N_928,N_1358);
nor U2056 (N_2056,N_959,N_1110);
and U2057 (N_2057,N_843,N_898);
nand U2058 (N_2058,N_764,N_851);
nand U2059 (N_2059,N_1446,N_855);
nand U2060 (N_2060,N_1173,N_1278);
and U2061 (N_2061,N_1033,N_1229);
nand U2062 (N_2062,N_1048,N_1481);
or U2063 (N_2063,N_1310,N_1480);
nor U2064 (N_2064,N_999,N_1190);
nor U2065 (N_2065,N_1199,N_971);
nand U2066 (N_2066,N_1250,N_1272);
and U2067 (N_2067,N_1357,N_1361);
nor U2068 (N_2068,N_1050,N_1315);
nor U2069 (N_2069,N_945,N_840);
and U2070 (N_2070,N_820,N_988);
or U2071 (N_2071,N_968,N_1458);
nor U2072 (N_2072,N_1242,N_871);
nand U2073 (N_2073,N_1450,N_908);
nand U2074 (N_2074,N_1015,N_921);
or U2075 (N_2075,N_1259,N_1050);
nand U2076 (N_2076,N_1183,N_905);
nand U2077 (N_2077,N_1294,N_1437);
or U2078 (N_2078,N_1028,N_864);
nor U2079 (N_2079,N_888,N_1054);
nand U2080 (N_2080,N_1162,N_1011);
or U2081 (N_2081,N_1142,N_1255);
nand U2082 (N_2082,N_1297,N_1075);
or U2083 (N_2083,N_873,N_1145);
and U2084 (N_2084,N_838,N_1277);
nand U2085 (N_2085,N_862,N_912);
nor U2086 (N_2086,N_871,N_1307);
nand U2087 (N_2087,N_916,N_1428);
nor U2088 (N_2088,N_1417,N_1252);
or U2089 (N_2089,N_1370,N_1379);
nand U2090 (N_2090,N_760,N_1246);
or U2091 (N_2091,N_1038,N_1394);
and U2092 (N_2092,N_1403,N_838);
or U2093 (N_2093,N_1038,N_1066);
or U2094 (N_2094,N_1175,N_1480);
or U2095 (N_2095,N_1383,N_1021);
or U2096 (N_2096,N_980,N_1340);
nor U2097 (N_2097,N_881,N_862);
and U2098 (N_2098,N_844,N_1478);
or U2099 (N_2099,N_1253,N_966);
nor U2100 (N_2100,N_775,N_1470);
nor U2101 (N_2101,N_1331,N_877);
or U2102 (N_2102,N_899,N_777);
and U2103 (N_2103,N_1383,N_1141);
nand U2104 (N_2104,N_900,N_1247);
and U2105 (N_2105,N_1157,N_982);
nand U2106 (N_2106,N_1219,N_1271);
nand U2107 (N_2107,N_899,N_1071);
or U2108 (N_2108,N_1039,N_1090);
and U2109 (N_2109,N_1195,N_1356);
and U2110 (N_2110,N_1300,N_803);
nor U2111 (N_2111,N_1024,N_989);
nor U2112 (N_2112,N_1266,N_771);
nor U2113 (N_2113,N_1192,N_873);
and U2114 (N_2114,N_1252,N_1381);
nor U2115 (N_2115,N_1106,N_873);
xnor U2116 (N_2116,N_862,N_1427);
nor U2117 (N_2117,N_1265,N_1390);
nor U2118 (N_2118,N_1167,N_789);
or U2119 (N_2119,N_1145,N_1494);
and U2120 (N_2120,N_1121,N_1220);
nand U2121 (N_2121,N_1079,N_1190);
or U2122 (N_2122,N_1475,N_1111);
or U2123 (N_2123,N_957,N_834);
and U2124 (N_2124,N_1316,N_1221);
and U2125 (N_2125,N_1429,N_1371);
nand U2126 (N_2126,N_1319,N_1183);
or U2127 (N_2127,N_1017,N_807);
and U2128 (N_2128,N_916,N_1310);
nand U2129 (N_2129,N_1203,N_1010);
or U2130 (N_2130,N_1395,N_1388);
and U2131 (N_2131,N_870,N_1095);
nor U2132 (N_2132,N_757,N_978);
and U2133 (N_2133,N_1187,N_1240);
and U2134 (N_2134,N_1271,N_878);
xnor U2135 (N_2135,N_1197,N_1326);
or U2136 (N_2136,N_1419,N_1268);
nor U2137 (N_2137,N_830,N_1356);
and U2138 (N_2138,N_1296,N_1328);
and U2139 (N_2139,N_871,N_750);
and U2140 (N_2140,N_819,N_1123);
nand U2141 (N_2141,N_1013,N_1449);
nor U2142 (N_2142,N_937,N_1326);
nand U2143 (N_2143,N_1054,N_1440);
nand U2144 (N_2144,N_785,N_1126);
nor U2145 (N_2145,N_1327,N_1465);
or U2146 (N_2146,N_1024,N_1162);
nor U2147 (N_2147,N_934,N_1027);
nor U2148 (N_2148,N_1098,N_982);
nor U2149 (N_2149,N_1298,N_1174);
nor U2150 (N_2150,N_917,N_1436);
nand U2151 (N_2151,N_961,N_1155);
nand U2152 (N_2152,N_900,N_1024);
and U2153 (N_2153,N_890,N_1120);
or U2154 (N_2154,N_1436,N_890);
and U2155 (N_2155,N_1341,N_758);
or U2156 (N_2156,N_1252,N_1341);
nand U2157 (N_2157,N_829,N_1029);
nor U2158 (N_2158,N_1359,N_1418);
or U2159 (N_2159,N_1033,N_1182);
and U2160 (N_2160,N_1022,N_762);
or U2161 (N_2161,N_1312,N_1015);
nor U2162 (N_2162,N_811,N_1332);
nand U2163 (N_2163,N_758,N_1293);
or U2164 (N_2164,N_1005,N_1343);
and U2165 (N_2165,N_1163,N_1342);
and U2166 (N_2166,N_1093,N_822);
and U2167 (N_2167,N_1053,N_1109);
or U2168 (N_2168,N_987,N_1244);
or U2169 (N_2169,N_1406,N_1032);
nand U2170 (N_2170,N_1014,N_810);
nor U2171 (N_2171,N_877,N_1491);
xnor U2172 (N_2172,N_788,N_1235);
or U2173 (N_2173,N_1201,N_1006);
and U2174 (N_2174,N_1277,N_1460);
nand U2175 (N_2175,N_1303,N_1411);
nor U2176 (N_2176,N_1430,N_1454);
and U2177 (N_2177,N_999,N_1402);
or U2178 (N_2178,N_1431,N_855);
nor U2179 (N_2179,N_1164,N_820);
and U2180 (N_2180,N_840,N_1339);
nor U2181 (N_2181,N_1323,N_1291);
and U2182 (N_2182,N_1066,N_1139);
nor U2183 (N_2183,N_1203,N_1462);
nand U2184 (N_2184,N_1060,N_904);
nand U2185 (N_2185,N_1039,N_1034);
nand U2186 (N_2186,N_942,N_856);
or U2187 (N_2187,N_1151,N_1092);
nor U2188 (N_2188,N_1330,N_1350);
nand U2189 (N_2189,N_1260,N_905);
and U2190 (N_2190,N_818,N_1022);
nand U2191 (N_2191,N_1401,N_1485);
or U2192 (N_2192,N_1215,N_1100);
nor U2193 (N_2193,N_890,N_1109);
nand U2194 (N_2194,N_1329,N_915);
or U2195 (N_2195,N_1431,N_1227);
xor U2196 (N_2196,N_1122,N_1443);
nand U2197 (N_2197,N_1467,N_786);
or U2198 (N_2198,N_1382,N_764);
nand U2199 (N_2199,N_817,N_1158);
and U2200 (N_2200,N_1461,N_914);
nor U2201 (N_2201,N_903,N_1405);
nor U2202 (N_2202,N_803,N_815);
nand U2203 (N_2203,N_914,N_1284);
nor U2204 (N_2204,N_1004,N_842);
and U2205 (N_2205,N_900,N_899);
nor U2206 (N_2206,N_1273,N_1135);
nor U2207 (N_2207,N_1034,N_1342);
nor U2208 (N_2208,N_1356,N_831);
or U2209 (N_2209,N_833,N_1072);
nor U2210 (N_2210,N_1102,N_1449);
nor U2211 (N_2211,N_1347,N_1228);
nand U2212 (N_2212,N_1068,N_1443);
nand U2213 (N_2213,N_1469,N_1389);
nor U2214 (N_2214,N_1446,N_1214);
and U2215 (N_2215,N_1458,N_883);
nand U2216 (N_2216,N_1394,N_1137);
or U2217 (N_2217,N_1077,N_984);
or U2218 (N_2218,N_1206,N_1283);
or U2219 (N_2219,N_778,N_1177);
or U2220 (N_2220,N_1302,N_1156);
or U2221 (N_2221,N_1184,N_1341);
nor U2222 (N_2222,N_1164,N_993);
xor U2223 (N_2223,N_1050,N_880);
nor U2224 (N_2224,N_869,N_1235);
nand U2225 (N_2225,N_1368,N_904);
or U2226 (N_2226,N_847,N_1345);
and U2227 (N_2227,N_959,N_931);
and U2228 (N_2228,N_969,N_1036);
nand U2229 (N_2229,N_1206,N_1186);
nand U2230 (N_2230,N_1322,N_788);
nand U2231 (N_2231,N_1125,N_888);
nor U2232 (N_2232,N_1215,N_1090);
nor U2233 (N_2233,N_1440,N_1367);
nor U2234 (N_2234,N_1226,N_981);
nand U2235 (N_2235,N_1246,N_1335);
and U2236 (N_2236,N_1317,N_815);
or U2237 (N_2237,N_1046,N_871);
nand U2238 (N_2238,N_1264,N_955);
and U2239 (N_2239,N_1305,N_1175);
or U2240 (N_2240,N_1167,N_897);
or U2241 (N_2241,N_1188,N_1113);
or U2242 (N_2242,N_773,N_1015);
or U2243 (N_2243,N_1314,N_992);
or U2244 (N_2244,N_989,N_892);
or U2245 (N_2245,N_784,N_920);
and U2246 (N_2246,N_1147,N_908);
or U2247 (N_2247,N_853,N_1469);
and U2248 (N_2248,N_869,N_1096);
nor U2249 (N_2249,N_1415,N_1026);
nand U2250 (N_2250,N_1926,N_2178);
nor U2251 (N_2251,N_2091,N_1662);
or U2252 (N_2252,N_2116,N_2108);
or U2253 (N_2253,N_2183,N_1761);
and U2254 (N_2254,N_1891,N_1777);
nor U2255 (N_2255,N_1687,N_1836);
nand U2256 (N_2256,N_1503,N_2002);
nor U2257 (N_2257,N_1530,N_1900);
nand U2258 (N_2258,N_1974,N_1847);
nand U2259 (N_2259,N_2149,N_2119);
or U2260 (N_2260,N_1760,N_2015);
nor U2261 (N_2261,N_1747,N_2135);
nand U2262 (N_2262,N_1507,N_1615);
nand U2263 (N_2263,N_2207,N_2208);
or U2264 (N_2264,N_1585,N_1800);
and U2265 (N_2265,N_1702,N_2033);
and U2266 (N_2266,N_1805,N_1816);
or U2267 (N_2267,N_1531,N_2113);
and U2268 (N_2268,N_1524,N_2234);
or U2269 (N_2269,N_2176,N_1655);
and U2270 (N_2270,N_1809,N_1521);
nand U2271 (N_2271,N_1882,N_1993);
and U2272 (N_2272,N_2164,N_1699);
nand U2273 (N_2273,N_1557,N_1877);
nand U2274 (N_2274,N_2014,N_2161);
nand U2275 (N_2275,N_2011,N_2030);
and U2276 (N_2276,N_1810,N_1784);
nand U2277 (N_2277,N_1646,N_2189);
nand U2278 (N_2278,N_1942,N_2168);
or U2279 (N_2279,N_1613,N_1617);
nor U2280 (N_2280,N_1846,N_2248);
or U2281 (N_2281,N_2105,N_2055);
nor U2282 (N_2282,N_1515,N_1685);
and U2283 (N_2283,N_1778,N_2231);
and U2284 (N_2284,N_1684,N_1929);
or U2285 (N_2285,N_1643,N_2124);
nor U2286 (N_2286,N_2196,N_2107);
or U2287 (N_2287,N_1916,N_1791);
and U2288 (N_2288,N_2089,N_1868);
nand U2289 (N_2289,N_2080,N_2115);
and U2290 (N_2290,N_1776,N_2146);
nor U2291 (N_2291,N_1710,N_1709);
nor U2292 (N_2292,N_1548,N_1894);
nor U2293 (N_2293,N_2134,N_2143);
or U2294 (N_2294,N_2102,N_1964);
or U2295 (N_2295,N_1682,N_1774);
and U2296 (N_2296,N_1647,N_2037);
nor U2297 (N_2297,N_1775,N_1696);
nor U2298 (N_2298,N_2040,N_2085);
nand U2299 (N_2299,N_2222,N_1580);
or U2300 (N_2300,N_1568,N_1952);
nand U2301 (N_2301,N_1915,N_1637);
nor U2302 (N_2302,N_1626,N_2050);
and U2303 (N_2303,N_1962,N_1931);
nand U2304 (N_2304,N_1554,N_1712);
or U2305 (N_2305,N_1513,N_1988);
nand U2306 (N_2306,N_1583,N_1560);
or U2307 (N_2307,N_1946,N_1725);
and U2308 (N_2308,N_2021,N_1860);
nor U2309 (N_2309,N_1551,N_1832);
nand U2310 (N_2310,N_1833,N_1787);
or U2311 (N_2311,N_1566,N_1971);
and U2312 (N_2312,N_1511,N_2086);
xnor U2313 (N_2313,N_2166,N_1883);
nand U2314 (N_2314,N_2063,N_1677);
nor U2315 (N_2315,N_2145,N_2126);
nor U2316 (N_2316,N_1622,N_2219);
and U2317 (N_2317,N_1855,N_1667);
and U2318 (N_2318,N_1674,N_2016);
and U2319 (N_2319,N_2000,N_1562);
or U2320 (N_2320,N_1576,N_1943);
nand U2321 (N_2321,N_1698,N_1893);
and U2322 (N_2322,N_2043,N_1895);
nand U2323 (N_2323,N_1748,N_2154);
nor U2324 (N_2324,N_1889,N_1992);
nand U2325 (N_2325,N_1796,N_1652);
and U2326 (N_2326,N_1595,N_2028);
nand U2327 (N_2327,N_1870,N_2090);
nand U2328 (N_2328,N_1506,N_1565);
nand U2329 (N_2329,N_1753,N_2203);
or U2330 (N_2330,N_2067,N_1913);
nand U2331 (N_2331,N_2026,N_1542);
nand U2332 (N_2332,N_1979,N_1851);
or U2333 (N_2333,N_2110,N_1885);
and U2334 (N_2334,N_1945,N_1737);
nor U2335 (N_2335,N_2204,N_2103);
nor U2336 (N_2336,N_1789,N_2242);
nor U2337 (N_2337,N_1909,N_1597);
or U2338 (N_2338,N_1839,N_1607);
nor U2339 (N_2339,N_2013,N_1648);
nor U2340 (N_2340,N_1938,N_1936);
nand U2341 (N_2341,N_2214,N_1547);
or U2342 (N_2342,N_1749,N_1518);
and U2343 (N_2343,N_2212,N_1624);
nor U2344 (N_2344,N_2081,N_1544);
nand U2345 (N_2345,N_2078,N_1584);
nand U2346 (N_2346,N_1865,N_2133);
nand U2347 (N_2347,N_2136,N_1527);
nor U2348 (N_2348,N_1975,N_1899);
nand U2349 (N_2349,N_1813,N_1766);
nand U2350 (N_2350,N_1944,N_1767);
and U2351 (N_2351,N_1733,N_1538);
nor U2352 (N_2352,N_1934,N_1969);
or U2353 (N_2353,N_1582,N_1999);
nor U2354 (N_2354,N_1540,N_2224);
or U2355 (N_2355,N_2087,N_1845);
and U2356 (N_2356,N_2047,N_1773);
and U2357 (N_2357,N_2093,N_1956);
nor U2358 (N_2358,N_1953,N_1740);
and U2359 (N_2359,N_2019,N_2174);
and U2360 (N_2360,N_1739,N_2117);
nor U2361 (N_2361,N_1627,N_2054);
or U2362 (N_2362,N_1780,N_1572);
and U2363 (N_2363,N_1676,N_2240);
xor U2364 (N_2364,N_2202,N_1982);
or U2365 (N_2365,N_1609,N_1922);
nor U2366 (N_2366,N_1686,N_2035);
nor U2367 (N_2367,N_2036,N_1605);
nand U2368 (N_2368,N_1857,N_1886);
nand U2369 (N_2369,N_1917,N_1879);
nand U2370 (N_2370,N_1995,N_1631);
and U2371 (N_2371,N_2144,N_1972);
or U2372 (N_2372,N_1821,N_1630);
or U2373 (N_2373,N_2139,N_2160);
or U2374 (N_2374,N_1587,N_2238);
or U2375 (N_2375,N_1859,N_1701);
or U2376 (N_2376,N_1850,N_2120);
nand U2377 (N_2377,N_2083,N_2150);
nand U2378 (N_2378,N_2111,N_1672);
or U2379 (N_2379,N_1644,N_2095);
or U2380 (N_2380,N_1723,N_1991);
or U2381 (N_2381,N_2209,N_2064);
nor U2382 (N_2382,N_2155,N_1835);
nor U2383 (N_2383,N_1711,N_2151);
and U2384 (N_2384,N_1724,N_2020);
nor U2385 (N_2385,N_1594,N_1755);
or U2386 (N_2386,N_1878,N_1692);
or U2387 (N_2387,N_2129,N_2073);
nor U2388 (N_2388,N_1681,N_1678);
nor U2389 (N_2389,N_1852,N_1892);
nand U2390 (N_2390,N_2058,N_1512);
nand U2391 (N_2391,N_1553,N_1657);
or U2392 (N_2392,N_1638,N_1951);
nand U2393 (N_2393,N_1793,N_2070);
nor U2394 (N_2394,N_2138,N_2235);
or U2395 (N_2395,N_1726,N_1700);
and U2396 (N_2396,N_1635,N_2186);
nor U2397 (N_2397,N_1887,N_2097);
or U2398 (N_2398,N_1798,N_1636);
nor U2399 (N_2399,N_1509,N_1939);
nor U2400 (N_2400,N_1842,N_1639);
nand U2401 (N_2401,N_1720,N_1785);
nand U2402 (N_2402,N_1792,N_1610);
nor U2403 (N_2403,N_2123,N_2236);
or U2404 (N_2404,N_1532,N_1935);
nand U2405 (N_2405,N_1732,N_1762);
nand U2406 (N_2406,N_2118,N_2101);
and U2407 (N_2407,N_1549,N_1574);
nor U2408 (N_2408,N_2059,N_2180);
and U2409 (N_2409,N_1522,N_1717);
nand U2410 (N_2410,N_1864,N_1693);
and U2411 (N_2411,N_1986,N_2132);
or U2412 (N_2412,N_2024,N_1754);
or U2413 (N_2413,N_2042,N_2092);
nand U2414 (N_2414,N_1608,N_1896);
nor U2415 (N_2415,N_1526,N_1640);
nand U2416 (N_2416,N_2072,N_2177);
or U2417 (N_2417,N_1914,N_2001);
and U2418 (N_2418,N_1559,N_1897);
and U2419 (N_2419,N_1653,N_1794);
or U2420 (N_2420,N_2074,N_1902);
nor U2421 (N_2421,N_1786,N_1694);
nor U2422 (N_2422,N_2084,N_1742);
nor U2423 (N_2423,N_1729,N_1884);
xnor U2424 (N_2424,N_1567,N_1820);
or U2425 (N_2425,N_1592,N_2034);
nor U2426 (N_2426,N_1843,N_1819);
nor U2427 (N_2427,N_2156,N_2220);
and U2428 (N_2428,N_1927,N_1933);
nor U2429 (N_2429,N_1603,N_1823);
or U2430 (N_2430,N_2025,N_1669);
nand U2431 (N_2431,N_1541,N_1660);
nor U2432 (N_2432,N_2049,N_1591);
and U2433 (N_2433,N_1704,N_1758);
nand U2434 (N_2434,N_1779,N_1598);
nand U2435 (N_2435,N_1683,N_2175);
nand U2436 (N_2436,N_1908,N_2159);
nand U2437 (N_2437,N_1705,N_1751);
nor U2438 (N_2438,N_1589,N_1966);
nand U2439 (N_2439,N_1930,N_2165);
nand U2440 (N_2440,N_2221,N_1604);
nand U2441 (N_2441,N_1750,N_1517);
and U2442 (N_2442,N_1960,N_2239);
and U2443 (N_2443,N_1659,N_1854);
nor U2444 (N_2444,N_1663,N_2065);
or U2445 (N_2445,N_2140,N_1921);
or U2446 (N_2446,N_1959,N_1826);
or U2447 (N_2447,N_1958,N_1715);
or U2448 (N_2448,N_1950,N_1872);
and U2449 (N_2449,N_2179,N_2184);
nand U2450 (N_2450,N_1937,N_1907);
nand U2451 (N_2451,N_1771,N_1856);
nand U2452 (N_2452,N_2162,N_1918);
or U2453 (N_2453,N_2247,N_2006);
nand U2454 (N_2454,N_1689,N_1756);
and U2455 (N_2455,N_2195,N_1623);
and U2456 (N_2456,N_1581,N_1871);
nor U2457 (N_2457,N_1695,N_2211);
or U2458 (N_2458,N_2096,N_2082);
nand U2459 (N_2459,N_1806,N_1743);
or U2460 (N_2460,N_1502,N_1781);
or U2461 (N_2461,N_1994,N_2171);
nand U2462 (N_2462,N_2125,N_2187);
and U2463 (N_2463,N_1911,N_1563);
nand U2464 (N_2464,N_2079,N_1713);
and U2465 (N_2465,N_1989,N_1963);
nor U2466 (N_2466,N_1601,N_2181);
nand U2467 (N_2467,N_2071,N_1831);
nor U2468 (N_2468,N_1814,N_1706);
nor U2469 (N_2469,N_2060,N_2018);
nand U2470 (N_2470,N_2010,N_2205);
or U2471 (N_2471,N_2007,N_1625);
or U2472 (N_2472,N_1973,N_1650);
nor U2473 (N_2473,N_1670,N_1874);
or U2474 (N_2474,N_1869,N_1984);
and U2475 (N_2475,N_2226,N_1998);
nor U2476 (N_2476,N_2163,N_2193);
or U2477 (N_2477,N_2029,N_2213);
nor U2478 (N_2478,N_1546,N_2228);
nor U2479 (N_2479,N_1519,N_1679);
nor U2480 (N_2480,N_1645,N_2056);
and U2481 (N_2481,N_1537,N_1719);
nor U2482 (N_2482,N_1664,N_1968);
and U2483 (N_2483,N_2022,N_2017);
nor U2484 (N_2484,N_2232,N_2053);
nor U2485 (N_2485,N_1783,N_1957);
nand U2486 (N_2486,N_2094,N_1703);
and U2487 (N_2487,N_2233,N_1803);
nand U2488 (N_2488,N_1673,N_2046);
nand U2489 (N_2489,N_1811,N_1641);
and U2490 (N_2490,N_2031,N_1508);
nand U2491 (N_2491,N_1578,N_2157);
nand U2492 (N_2492,N_2158,N_1634);
and U2493 (N_2493,N_1668,N_1661);
nand U2494 (N_2494,N_2199,N_1920);
or U2495 (N_2495,N_1718,N_2039);
and U2496 (N_2496,N_1525,N_1867);
and U2497 (N_2497,N_2147,N_1752);
and U2498 (N_2498,N_1649,N_1680);
xor U2499 (N_2499,N_2032,N_2023);
or U2500 (N_2500,N_2005,N_2173);
nor U2501 (N_2501,N_2137,N_1620);
nor U2502 (N_2502,N_1665,N_1500);
and U2503 (N_2503,N_1570,N_1690);
or U2504 (N_2504,N_1997,N_1834);
or U2505 (N_2505,N_1875,N_1797);
and U2506 (N_2506,N_1788,N_1577);
nor U2507 (N_2507,N_1782,N_2045);
and U2508 (N_2508,N_1504,N_2191);
and U2509 (N_2509,N_2122,N_2104);
nor U2510 (N_2510,N_1904,N_1925);
nand U2511 (N_2511,N_1545,N_1510);
or U2512 (N_2512,N_2077,N_1612);
nand U2513 (N_2513,N_1890,N_1849);
nand U2514 (N_2514,N_1881,N_1941);
or U2515 (N_2515,N_1799,N_2051);
nand U2516 (N_2516,N_2243,N_1656);
or U2517 (N_2517,N_2167,N_2185);
and U2518 (N_2518,N_1919,N_2112);
nand U2519 (N_2519,N_1817,N_2057);
nor U2520 (N_2520,N_1561,N_1880);
nand U2521 (N_2521,N_1822,N_1529);
xor U2522 (N_2522,N_1533,N_1731);
and U2523 (N_2523,N_1824,N_1523);
nor U2524 (N_2524,N_2172,N_1905);
nor U2525 (N_2525,N_2245,N_2201);
nand U2526 (N_2526,N_2061,N_1876);
and U2527 (N_2527,N_2062,N_1621);
nor U2528 (N_2528,N_1671,N_2197);
nand U2529 (N_2529,N_1837,N_1903);
nor U2530 (N_2530,N_2237,N_2027);
or U2531 (N_2531,N_1632,N_2200);
nand U2532 (N_2532,N_2215,N_1734);
and U2533 (N_2533,N_2246,N_2003);
or U2534 (N_2534,N_1516,N_2241);
and U2535 (N_2535,N_1539,N_1534);
and U2536 (N_2536,N_2148,N_2044);
and U2537 (N_2537,N_1770,N_1616);
or U2538 (N_2538,N_1602,N_1866);
nand U2539 (N_2539,N_1790,N_1716);
nor U2540 (N_2540,N_1741,N_2153);
or U2541 (N_2541,N_1815,N_2225);
nand U2542 (N_2542,N_1599,N_1745);
nand U2543 (N_2543,N_1901,N_1629);
nor U2544 (N_2544,N_1571,N_1688);
and U2545 (N_2545,N_1888,N_1848);
and U2546 (N_2546,N_1863,N_1965);
nand U2547 (N_2547,N_1593,N_1691);
or U2548 (N_2548,N_1873,N_1736);
or U2549 (N_2549,N_1569,N_1543);
and U2550 (N_2550,N_1768,N_1642);
and U2551 (N_2551,N_2008,N_1765);
nand U2552 (N_2552,N_1556,N_2009);
nor U2553 (N_2553,N_1853,N_2169);
or U2554 (N_2554,N_1552,N_1611);
nand U2555 (N_2555,N_2048,N_1746);
or U2556 (N_2556,N_2229,N_1708);
and U2557 (N_2557,N_1520,N_1619);
nand U2558 (N_2558,N_2041,N_2038);
or U2559 (N_2559,N_1714,N_1928);
nand U2560 (N_2560,N_1514,N_1600);
nor U2561 (N_2561,N_2142,N_2052);
and U2562 (N_2562,N_1721,N_1955);
and U2563 (N_2563,N_1802,N_2098);
nor U2564 (N_2564,N_1808,N_2012);
nor U2565 (N_2565,N_1590,N_1829);
and U2566 (N_2566,N_1618,N_1769);
and U2567 (N_2567,N_1633,N_1588);
and U2568 (N_2568,N_1772,N_1978);
nor U2569 (N_2569,N_1861,N_2152);
nand U2570 (N_2570,N_1697,N_1987);
or U2571 (N_2571,N_2099,N_1807);
and U2572 (N_2572,N_1801,N_1940);
nor U2573 (N_2573,N_2128,N_1967);
and U2574 (N_2574,N_1505,N_1949);
and U2575 (N_2575,N_1764,N_2131);
xor U2576 (N_2576,N_2206,N_1675);
nor U2577 (N_2577,N_1586,N_1830);
or U2578 (N_2578,N_2127,N_1932);
nand U2579 (N_2579,N_1898,N_2075);
nor U2580 (N_2580,N_2216,N_2068);
nand U2581 (N_2581,N_1727,N_2244);
and U2582 (N_2582,N_1757,N_1840);
or U2583 (N_2583,N_1906,N_1923);
nand U2584 (N_2584,N_2121,N_1985);
nand U2585 (N_2585,N_1825,N_1573);
and U2586 (N_2586,N_1795,N_1614);
or U2587 (N_2587,N_1738,N_1947);
or U2588 (N_2588,N_2218,N_1763);
nor U2589 (N_2589,N_1536,N_1961);
nor U2590 (N_2590,N_1970,N_2100);
nor U2591 (N_2591,N_1910,N_1759);
nand U2592 (N_2592,N_1924,N_2141);
nor U2593 (N_2593,N_2192,N_2194);
nand U2594 (N_2594,N_1735,N_1804);
nand U2595 (N_2595,N_1535,N_1980);
nor U2596 (N_2596,N_1841,N_2198);
or U2597 (N_2597,N_1628,N_1606);
nand U2598 (N_2598,N_1862,N_2182);
and U2599 (N_2599,N_1844,N_1744);
nand U2600 (N_2600,N_1555,N_1654);
nor U2601 (N_2601,N_1651,N_1707);
nor U2602 (N_2602,N_2227,N_1564);
nor U2603 (N_2603,N_1579,N_2114);
nand U2604 (N_2604,N_1730,N_2069);
or U2605 (N_2605,N_1954,N_1838);
nor U2606 (N_2606,N_1858,N_1990);
nor U2607 (N_2607,N_1981,N_2217);
or U2608 (N_2608,N_2106,N_1528);
or U2609 (N_2609,N_2210,N_1558);
and U2610 (N_2610,N_1666,N_1501);
nand U2611 (N_2611,N_2076,N_2066);
nand U2612 (N_2612,N_2230,N_1728);
and U2613 (N_2613,N_2130,N_1976);
nor U2614 (N_2614,N_1828,N_1722);
and U2615 (N_2615,N_2223,N_2190);
or U2616 (N_2616,N_1812,N_2109);
or U2617 (N_2617,N_1818,N_2004);
nor U2618 (N_2618,N_1977,N_1912);
nor U2619 (N_2619,N_2088,N_2170);
nor U2620 (N_2620,N_2249,N_1948);
and U2621 (N_2621,N_1658,N_1827);
nor U2622 (N_2622,N_1550,N_2188);
nor U2623 (N_2623,N_1996,N_1596);
or U2624 (N_2624,N_1983,N_1575);
nor U2625 (N_2625,N_1988,N_1690);
nand U2626 (N_2626,N_1507,N_2139);
and U2627 (N_2627,N_1741,N_1646);
or U2628 (N_2628,N_2088,N_1611);
or U2629 (N_2629,N_1600,N_1740);
nor U2630 (N_2630,N_1805,N_2107);
nor U2631 (N_2631,N_1819,N_1572);
nand U2632 (N_2632,N_1893,N_1631);
and U2633 (N_2633,N_1920,N_1916);
and U2634 (N_2634,N_1941,N_2103);
nor U2635 (N_2635,N_1988,N_2056);
or U2636 (N_2636,N_1736,N_1751);
nor U2637 (N_2637,N_1553,N_1530);
nand U2638 (N_2638,N_1924,N_1942);
xor U2639 (N_2639,N_1850,N_1977);
nand U2640 (N_2640,N_1807,N_1933);
and U2641 (N_2641,N_2073,N_2086);
and U2642 (N_2642,N_1545,N_1636);
and U2643 (N_2643,N_2243,N_1676);
nor U2644 (N_2644,N_1725,N_2231);
or U2645 (N_2645,N_1689,N_1787);
nand U2646 (N_2646,N_1991,N_1626);
nor U2647 (N_2647,N_1857,N_1646);
nand U2648 (N_2648,N_1637,N_1587);
or U2649 (N_2649,N_1610,N_1921);
nor U2650 (N_2650,N_1649,N_1544);
nand U2651 (N_2651,N_2131,N_2144);
and U2652 (N_2652,N_1749,N_2172);
and U2653 (N_2653,N_1754,N_2132);
and U2654 (N_2654,N_1611,N_1719);
or U2655 (N_2655,N_2226,N_1747);
and U2656 (N_2656,N_2229,N_1749);
and U2657 (N_2657,N_2133,N_2065);
or U2658 (N_2658,N_1671,N_1650);
nand U2659 (N_2659,N_1791,N_1756);
nand U2660 (N_2660,N_1947,N_2179);
and U2661 (N_2661,N_1781,N_1854);
or U2662 (N_2662,N_1746,N_2084);
nand U2663 (N_2663,N_1510,N_1953);
nand U2664 (N_2664,N_1858,N_1658);
nor U2665 (N_2665,N_1786,N_1569);
and U2666 (N_2666,N_2231,N_1927);
nor U2667 (N_2667,N_2228,N_2155);
nor U2668 (N_2668,N_2219,N_2109);
or U2669 (N_2669,N_1578,N_1793);
nor U2670 (N_2670,N_1679,N_1582);
nor U2671 (N_2671,N_2165,N_2076);
and U2672 (N_2672,N_1780,N_2236);
or U2673 (N_2673,N_1643,N_1983);
and U2674 (N_2674,N_1583,N_1523);
nand U2675 (N_2675,N_1650,N_1576);
and U2676 (N_2676,N_1689,N_1915);
nor U2677 (N_2677,N_1523,N_1530);
or U2678 (N_2678,N_2072,N_2069);
nor U2679 (N_2679,N_1654,N_1512);
nand U2680 (N_2680,N_1646,N_2131);
nand U2681 (N_2681,N_1984,N_2157);
and U2682 (N_2682,N_1684,N_2140);
or U2683 (N_2683,N_2093,N_2018);
and U2684 (N_2684,N_1969,N_2203);
and U2685 (N_2685,N_1803,N_2091);
nor U2686 (N_2686,N_2012,N_1956);
or U2687 (N_2687,N_1596,N_2025);
nand U2688 (N_2688,N_1994,N_1723);
nand U2689 (N_2689,N_2034,N_1801);
nor U2690 (N_2690,N_2125,N_1516);
nor U2691 (N_2691,N_2125,N_1865);
or U2692 (N_2692,N_2133,N_2016);
nor U2693 (N_2693,N_1931,N_2028);
nand U2694 (N_2694,N_1841,N_1684);
and U2695 (N_2695,N_1520,N_1840);
xor U2696 (N_2696,N_2082,N_1961);
and U2697 (N_2697,N_1898,N_2086);
and U2698 (N_2698,N_2002,N_1704);
or U2699 (N_2699,N_1503,N_1673);
nand U2700 (N_2700,N_2004,N_1736);
or U2701 (N_2701,N_1718,N_2105);
and U2702 (N_2702,N_1931,N_2181);
and U2703 (N_2703,N_2159,N_1741);
or U2704 (N_2704,N_1908,N_2115);
or U2705 (N_2705,N_1528,N_2185);
nand U2706 (N_2706,N_1784,N_1931);
nand U2707 (N_2707,N_2192,N_1722);
or U2708 (N_2708,N_1630,N_1782);
or U2709 (N_2709,N_2097,N_2048);
nand U2710 (N_2710,N_1850,N_1949);
and U2711 (N_2711,N_1567,N_1679);
and U2712 (N_2712,N_1585,N_2038);
nand U2713 (N_2713,N_2158,N_1887);
or U2714 (N_2714,N_2084,N_1540);
or U2715 (N_2715,N_1529,N_1955);
and U2716 (N_2716,N_2213,N_1705);
nand U2717 (N_2717,N_1827,N_1743);
and U2718 (N_2718,N_2121,N_1674);
or U2719 (N_2719,N_2097,N_1893);
nand U2720 (N_2720,N_1724,N_2049);
and U2721 (N_2721,N_1640,N_1676);
or U2722 (N_2722,N_2034,N_1661);
or U2723 (N_2723,N_2141,N_2246);
and U2724 (N_2724,N_1689,N_1592);
nand U2725 (N_2725,N_1664,N_1711);
nand U2726 (N_2726,N_1658,N_2031);
or U2727 (N_2727,N_2230,N_1718);
nor U2728 (N_2728,N_1647,N_1884);
or U2729 (N_2729,N_1844,N_1859);
nor U2730 (N_2730,N_2041,N_1677);
or U2731 (N_2731,N_2023,N_1885);
nand U2732 (N_2732,N_2140,N_1806);
nand U2733 (N_2733,N_1813,N_2085);
or U2734 (N_2734,N_1649,N_1546);
nand U2735 (N_2735,N_2153,N_1706);
nor U2736 (N_2736,N_2246,N_2091);
and U2737 (N_2737,N_1816,N_2078);
nor U2738 (N_2738,N_1614,N_1609);
nand U2739 (N_2739,N_1725,N_1797);
or U2740 (N_2740,N_1852,N_1768);
xnor U2741 (N_2741,N_1986,N_1978);
nand U2742 (N_2742,N_1703,N_2057);
and U2743 (N_2743,N_2008,N_1686);
or U2744 (N_2744,N_1860,N_1603);
or U2745 (N_2745,N_1657,N_2076);
nand U2746 (N_2746,N_1689,N_1769);
nor U2747 (N_2747,N_1918,N_2020);
and U2748 (N_2748,N_1756,N_2045);
nand U2749 (N_2749,N_1814,N_1811);
or U2750 (N_2750,N_1734,N_2177);
nor U2751 (N_2751,N_1819,N_2013);
and U2752 (N_2752,N_1620,N_1618);
nand U2753 (N_2753,N_1919,N_1888);
and U2754 (N_2754,N_2019,N_1747);
nor U2755 (N_2755,N_1778,N_2110);
or U2756 (N_2756,N_1871,N_1650);
or U2757 (N_2757,N_2175,N_1553);
or U2758 (N_2758,N_2051,N_1564);
nand U2759 (N_2759,N_2073,N_1703);
nand U2760 (N_2760,N_1956,N_1566);
nand U2761 (N_2761,N_1613,N_1776);
and U2762 (N_2762,N_1707,N_1548);
or U2763 (N_2763,N_2157,N_1712);
nor U2764 (N_2764,N_2189,N_1786);
nand U2765 (N_2765,N_1736,N_1948);
nor U2766 (N_2766,N_2244,N_2175);
nor U2767 (N_2767,N_2104,N_1531);
nand U2768 (N_2768,N_1564,N_2239);
nor U2769 (N_2769,N_2103,N_1866);
and U2770 (N_2770,N_2243,N_2028);
and U2771 (N_2771,N_1827,N_1947);
or U2772 (N_2772,N_1663,N_2055);
nor U2773 (N_2773,N_1900,N_1894);
or U2774 (N_2774,N_2032,N_2165);
and U2775 (N_2775,N_1630,N_1806);
nand U2776 (N_2776,N_2237,N_2161);
or U2777 (N_2777,N_1973,N_2188);
nor U2778 (N_2778,N_1687,N_1670);
and U2779 (N_2779,N_1532,N_2009);
nor U2780 (N_2780,N_1758,N_1863);
or U2781 (N_2781,N_2219,N_1542);
and U2782 (N_2782,N_2061,N_1552);
and U2783 (N_2783,N_1901,N_1538);
nor U2784 (N_2784,N_1713,N_2208);
and U2785 (N_2785,N_1673,N_2055);
nand U2786 (N_2786,N_2039,N_2091);
nor U2787 (N_2787,N_1758,N_1599);
nand U2788 (N_2788,N_1821,N_1796);
and U2789 (N_2789,N_2096,N_1861);
and U2790 (N_2790,N_1909,N_2023);
or U2791 (N_2791,N_1996,N_1612);
or U2792 (N_2792,N_2142,N_2237);
nor U2793 (N_2793,N_1693,N_1920);
xor U2794 (N_2794,N_1609,N_2234);
or U2795 (N_2795,N_1877,N_2100);
nand U2796 (N_2796,N_1700,N_1902);
nand U2797 (N_2797,N_1668,N_2199);
and U2798 (N_2798,N_2079,N_2043);
nand U2799 (N_2799,N_1649,N_1666);
and U2800 (N_2800,N_1611,N_1818);
nor U2801 (N_2801,N_2019,N_1619);
nor U2802 (N_2802,N_1906,N_2191);
and U2803 (N_2803,N_1861,N_1829);
and U2804 (N_2804,N_2164,N_1692);
nor U2805 (N_2805,N_2094,N_2157);
nor U2806 (N_2806,N_2192,N_2164);
xnor U2807 (N_2807,N_1769,N_1561);
and U2808 (N_2808,N_2074,N_1852);
nor U2809 (N_2809,N_2019,N_2017);
nor U2810 (N_2810,N_2033,N_2003);
nor U2811 (N_2811,N_1964,N_1647);
nand U2812 (N_2812,N_2229,N_2077);
or U2813 (N_2813,N_1702,N_1757);
nand U2814 (N_2814,N_2200,N_1672);
nand U2815 (N_2815,N_2151,N_1721);
and U2816 (N_2816,N_1875,N_1774);
and U2817 (N_2817,N_1967,N_1561);
nor U2818 (N_2818,N_1840,N_2172);
nor U2819 (N_2819,N_1772,N_1641);
nor U2820 (N_2820,N_1757,N_1512);
and U2821 (N_2821,N_1927,N_1908);
and U2822 (N_2822,N_1896,N_2001);
or U2823 (N_2823,N_1713,N_1961);
nor U2824 (N_2824,N_1814,N_1912);
nor U2825 (N_2825,N_1592,N_1928);
nand U2826 (N_2826,N_1676,N_1677);
nand U2827 (N_2827,N_1710,N_1560);
nor U2828 (N_2828,N_1671,N_1785);
and U2829 (N_2829,N_1514,N_1856);
nor U2830 (N_2830,N_1959,N_1816);
or U2831 (N_2831,N_1870,N_1539);
or U2832 (N_2832,N_1971,N_1625);
nand U2833 (N_2833,N_1817,N_2040);
and U2834 (N_2834,N_1711,N_1822);
nand U2835 (N_2835,N_1539,N_1666);
nor U2836 (N_2836,N_1688,N_1532);
and U2837 (N_2837,N_1710,N_2129);
or U2838 (N_2838,N_2137,N_1686);
and U2839 (N_2839,N_1971,N_2174);
and U2840 (N_2840,N_1967,N_1983);
nand U2841 (N_2841,N_1879,N_1840);
nor U2842 (N_2842,N_2240,N_2030);
and U2843 (N_2843,N_1927,N_2042);
and U2844 (N_2844,N_1837,N_2156);
nand U2845 (N_2845,N_2247,N_1583);
or U2846 (N_2846,N_1531,N_2098);
and U2847 (N_2847,N_1794,N_2243);
nor U2848 (N_2848,N_1973,N_1803);
or U2849 (N_2849,N_1689,N_2210);
nor U2850 (N_2850,N_1920,N_2090);
and U2851 (N_2851,N_1748,N_1790);
nand U2852 (N_2852,N_1890,N_2238);
nand U2853 (N_2853,N_1927,N_2169);
and U2854 (N_2854,N_1616,N_1753);
and U2855 (N_2855,N_1793,N_2083);
nand U2856 (N_2856,N_1946,N_2043);
nand U2857 (N_2857,N_1791,N_1769);
and U2858 (N_2858,N_1800,N_1685);
nand U2859 (N_2859,N_1720,N_1896);
nand U2860 (N_2860,N_2033,N_1541);
nand U2861 (N_2861,N_1525,N_1746);
or U2862 (N_2862,N_1538,N_1757);
and U2863 (N_2863,N_2142,N_1734);
and U2864 (N_2864,N_2021,N_2222);
nor U2865 (N_2865,N_1885,N_1844);
or U2866 (N_2866,N_1740,N_1945);
nand U2867 (N_2867,N_1928,N_2234);
or U2868 (N_2868,N_1537,N_2001);
and U2869 (N_2869,N_1551,N_2167);
and U2870 (N_2870,N_1859,N_1957);
and U2871 (N_2871,N_1584,N_1768);
nor U2872 (N_2872,N_1619,N_2249);
and U2873 (N_2873,N_2042,N_2086);
nor U2874 (N_2874,N_2219,N_2115);
or U2875 (N_2875,N_1566,N_1644);
nand U2876 (N_2876,N_1743,N_1791);
and U2877 (N_2877,N_2155,N_1907);
or U2878 (N_2878,N_2148,N_1966);
or U2879 (N_2879,N_2072,N_1601);
nand U2880 (N_2880,N_1610,N_1689);
and U2881 (N_2881,N_1994,N_1850);
and U2882 (N_2882,N_2210,N_1636);
nor U2883 (N_2883,N_1854,N_1859);
nor U2884 (N_2884,N_1686,N_1598);
nand U2885 (N_2885,N_1965,N_2235);
nor U2886 (N_2886,N_2138,N_1506);
xor U2887 (N_2887,N_2239,N_1834);
nor U2888 (N_2888,N_1643,N_1674);
nor U2889 (N_2889,N_2105,N_2192);
nor U2890 (N_2890,N_1757,N_2116);
nor U2891 (N_2891,N_2211,N_2155);
and U2892 (N_2892,N_1721,N_1893);
or U2893 (N_2893,N_1718,N_1879);
nand U2894 (N_2894,N_2075,N_2199);
nand U2895 (N_2895,N_2107,N_2109);
nand U2896 (N_2896,N_2068,N_1812);
and U2897 (N_2897,N_1811,N_2131);
xor U2898 (N_2898,N_1504,N_1690);
nor U2899 (N_2899,N_1766,N_1693);
and U2900 (N_2900,N_1817,N_1982);
nand U2901 (N_2901,N_1839,N_1979);
or U2902 (N_2902,N_2082,N_2068);
nor U2903 (N_2903,N_2002,N_1802);
nor U2904 (N_2904,N_1588,N_1974);
nor U2905 (N_2905,N_1508,N_1759);
or U2906 (N_2906,N_2120,N_1760);
or U2907 (N_2907,N_1831,N_2214);
and U2908 (N_2908,N_1527,N_1780);
or U2909 (N_2909,N_1906,N_1835);
nor U2910 (N_2910,N_2228,N_1992);
and U2911 (N_2911,N_1564,N_1610);
nand U2912 (N_2912,N_1860,N_2017);
nand U2913 (N_2913,N_1654,N_1943);
and U2914 (N_2914,N_1692,N_2228);
nand U2915 (N_2915,N_1819,N_1898);
nand U2916 (N_2916,N_1988,N_1845);
or U2917 (N_2917,N_2025,N_2190);
or U2918 (N_2918,N_1534,N_1976);
xor U2919 (N_2919,N_1632,N_1868);
nor U2920 (N_2920,N_1569,N_2208);
nand U2921 (N_2921,N_2227,N_1519);
nand U2922 (N_2922,N_1864,N_1593);
and U2923 (N_2923,N_2113,N_2198);
and U2924 (N_2924,N_2179,N_2232);
and U2925 (N_2925,N_1732,N_2041);
and U2926 (N_2926,N_1912,N_2152);
or U2927 (N_2927,N_1604,N_1851);
or U2928 (N_2928,N_1607,N_2199);
nand U2929 (N_2929,N_2172,N_1869);
and U2930 (N_2930,N_1703,N_1975);
or U2931 (N_2931,N_1525,N_1628);
nand U2932 (N_2932,N_1752,N_2052);
nor U2933 (N_2933,N_1538,N_1972);
and U2934 (N_2934,N_1905,N_2162);
nand U2935 (N_2935,N_1890,N_2178);
and U2936 (N_2936,N_1596,N_2155);
nand U2937 (N_2937,N_1597,N_1556);
nor U2938 (N_2938,N_2031,N_2212);
and U2939 (N_2939,N_1961,N_1821);
nor U2940 (N_2940,N_1728,N_1627);
nand U2941 (N_2941,N_1922,N_2128);
and U2942 (N_2942,N_2221,N_1996);
and U2943 (N_2943,N_2226,N_1666);
nand U2944 (N_2944,N_1511,N_1958);
and U2945 (N_2945,N_2209,N_2008);
nand U2946 (N_2946,N_1705,N_2126);
or U2947 (N_2947,N_2157,N_2241);
and U2948 (N_2948,N_1856,N_2033);
nand U2949 (N_2949,N_1766,N_2243);
nor U2950 (N_2950,N_2159,N_1605);
and U2951 (N_2951,N_1601,N_2021);
and U2952 (N_2952,N_1740,N_1984);
and U2953 (N_2953,N_2171,N_1842);
and U2954 (N_2954,N_1691,N_2216);
nand U2955 (N_2955,N_2209,N_2235);
and U2956 (N_2956,N_1823,N_1517);
nand U2957 (N_2957,N_1703,N_2084);
or U2958 (N_2958,N_2162,N_1986);
or U2959 (N_2959,N_1961,N_2210);
nor U2960 (N_2960,N_2194,N_2122);
and U2961 (N_2961,N_1971,N_1922);
nand U2962 (N_2962,N_1731,N_1726);
and U2963 (N_2963,N_2121,N_1895);
or U2964 (N_2964,N_1812,N_2204);
or U2965 (N_2965,N_1639,N_1834);
or U2966 (N_2966,N_1891,N_1836);
or U2967 (N_2967,N_2195,N_2066);
nand U2968 (N_2968,N_1724,N_2005);
nand U2969 (N_2969,N_1814,N_1846);
nand U2970 (N_2970,N_1852,N_1814);
nor U2971 (N_2971,N_2091,N_2052);
nand U2972 (N_2972,N_1632,N_1984);
or U2973 (N_2973,N_1812,N_1788);
or U2974 (N_2974,N_2139,N_2008);
nor U2975 (N_2975,N_1677,N_2149);
and U2976 (N_2976,N_1664,N_1645);
nand U2977 (N_2977,N_1923,N_1886);
nand U2978 (N_2978,N_2044,N_2069);
nor U2979 (N_2979,N_1778,N_2070);
and U2980 (N_2980,N_2031,N_2153);
and U2981 (N_2981,N_2157,N_1902);
nor U2982 (N_2982,N_1830,N_1771);
nand U2983 (N_2983,N_1750,N_1856);
and U2984 (N_2984,N_1656,N_1556);
or U2985 (N_2985,N_1549,N_1508);
and U2986 (N_2986,N_1952,N_1826);
nand U2987 (N_2987,N_1693,N_2197);
and U2988 (N_2988,N_1935,N_2086);
or U2989 (N_2989,N_2008,N_1655);
or U2990 (N_2990,N_2060,N_2089);
and U2991 (N_2991,N_1684,N_1586);
and U2992 (N_2992,N_2193,N_1657);
or U2993 (N_2993,N_1505,N_1576);
nor U2994 (N_2994,N_1969,N_1512);
and U2995 (N_2995,N_1554,N_1790);
or U2996 (N_2996,N_1784,N_2116);
nand U2997 (N_2997,N_1646,N_1584);
or U2998 (N_2998,N_2022,N_2132);
nor U2999 (N_2999,N_1931,N_2042);
nor UO_0 (O_0,N_2502,N_2867);
or UO_1 (O_1,N_2964,N_2656);
nor UO_2 (O_2,N_2564,N_2386);
or UO_3 (O_3,N_2920,N_2955);
or UO_4 (O_4,N_2724,N_2545);
and UO_5 (O_5,N_2938,N_2898);
and UO_6 (O_6,N_2276,N_2886);
or UO_7 (O_7,N_2852,N_2791);
or UO_8 (O_8,N_2485,N_2706);
and UO_9 (O_9,N_2625,N_2299);
xnor UO_10 (O_10,N_2712,N_2494);
and UO_11 (O_11,N_2830,N_2828);
nor UO_12 (O_12,N_2741,N_2322);
and UO_13 (O_13,N_2788,N_2780);
nand UO_14 (O_14,N_2650,N_2840);
or UO_15 (O_15,N_2398,N_2343);
nand UO_16 (O_16,N_2300,N_2407);
nor UO_17 (O_17,N_2691,N_2923);
nor UO_18 (O_18,N_2487,N_2874);
nand UO_19 (O_19,N_2423,N_2853);
nor UO_20 (O_20,N_2446,N_2538);
nor UO_21 (O_21,N_2293,N_2872);
and UO_22 (O_22,N_2355,N_2779);
or UO_23 (O_23,N_2353,N_2936);
and UO_24 (O_24,N_2774,N_2595);
nor UO_25 (O_25,N_2792,N_2908);
and UO_26 (O_26,N_2927,N_2399);
nor UO_27 (O_27,N_2611,N_2841);
nor UO_28 (O_28,N_2404,N_2555);
or UO_29 (O_29,N_2527,N_2847);
nor UO_30 (O_30,N_2848,N_2902);
and UO_31 (O_31,N_2272,N_2965);
or UO_32 (O_32,N_2713,N_2888);
nand UO_33 (O_33,N_2464,N_2419);
or UO_34 (O_34,N_2345,N_2462);
nand UO_35 (O_35,N_2914,N_2668);
or UO_36 (O_36,N_2410,N_2806);
or UO_37 (O_37,N_2534,N_2716);
nand UO_38 (O_38,N_2444,N_2893);
or UO_39 (O_39,N_2636,N_2903);
and UO_40 (O_40,N_2844,N_2510);
and UO_41 (O_41,N_2319,N_2929);
nor UO_42 (O_42,N_2687,N_2829);
and UO_43 (O_43,N_2470,N_2866);
nor UO_44 (O_44,N_2352,N_2403);
nand UO_45 (O_45,N_2744,N_2646);
and UO_46 (O_46,N_2381,N_2608);
and UO_47 (O_47,N_2537,N_2270);
or UO_48 (O_48,N_2569,N_2439);
and UO_49 (O_49,N_2368,N_2676);
nor UO_50 (O_50,N_2359,N_2428);
nand UO_51 (O_51,N_2489,N_2890);
and UO_52 (O_52,N_2473,N_2523);
nand UO_53 (O_53,N_2605,N_2918);
nor UO_54 (O_54,N_2394,N_2642);
and UO_55 (O_55,N_2580,N_2651);
nor UO_56 (O_56,N_2518,N_2887);
or UO_57 (O_57,N_2937,N_2686);
or UO_58 (O_58,N_2800,N_2274);
and UO_59 (O_59,N_2333,N_2296);
nor UO_60 (O_60,N_2305,N_2496);
nor UO_61 (O_61,N_2863,N_2568);
nand UO_62 (O_62,N_2254,N_2412);
nor UO_63 (O_63,N_2490,N_2382);
xor UO_64 (O_64,N_2397,N_2856);
and UO_65 (O_65,N_2973,N_2384);
nor UO_66 (O_66,N_2358,N_2837);
nand UO_67 (O_67,N_2786,N_2962);
or UO_68 (O_68,N_2543,N_2635);
nor UO_69 (O_69,N_2776,N_2777);
and UO_70 (O_70,N_2430,N_2609);
nor UO_71 (O_71,N_2435,N_2836);
nor UO_72 (O_72,N_2324,N_2804);
nand UO_73 (O_73,N_2453,N_2339);
nor UO_74 (O_74,N_2869,N_2730);
and UO_75 (O_75,N_2793,N_2375);
nor UO_76 (O_76,N_2680,N_2935);
nand UO_77 (O_77,N_2986,N_2311);
and UO_78 (O_78,N_2501,N_2586);
nor UO_79 (O_79,N_2910,N_2495);
or UO_80 (O_80,N_2732,N_2572);
or UO_81 (O_81,N_2374,N_2729);
and UO_82 (O_82,N_2942,N_2400);
nor UO_83 (O_83,N_2811,N_2778);
and UO_84 (O_84,N_2924,N_2907);
nor UO_85 (O_85,N_2463,N_2758);
or UO_86 (O_86,N_2912,N_2885);
and UO_87 (O_87,N_2309,N_2413);
or UO_88 (O_88,N_2367,N_2648);
or UO_89 (O_89,N_2633,N_2566);
nand UO_90 (O_90,N_2548,N_2693);
nor UO_91 (O_91,N_2775,N_2554);
nor UO_92 (O_92,N_2892,N_2748);
or UO_93 (O_93,N_2610,N_2431);
nand UO_94 (O_94,N_2972,N_2292);
and UO_95 (O_95,N_2768,N_2736);
and UO_96 (O_96,N_2370,N_2369);
or UO_97 (O_97,N_2275,N_2544);
or UO_98 (O_98,N_2714,N_2858);
and UO_99 (O_99,N_2959,N_2969);
nand UO_100 (O_100,N_2700,N_2773);
nor UO_101 (O_101,N_2406,N_2875);
and UO_102 (O_102,N_2949,N_2402);
and UO_103 (O_103,N_2993,N_2436);
or UO_104 (O_104,N_2575,N_2612);
nor UO_105 (O_105,N_2963,N_2817);
or UO_106 (O_106,N_2926,N_2469);
nor UO_107 (O_107,N_2366,N_2442);
or UO_108 (O_108,N_2497,N_2287);
nand UO_109 (O_109,N_2522,N_2316);
nor UO_110 (O_110,N_2432,N_2392);
nand UO_111 (O_111,N_2873,N_2931);
and UO_112 (O_112,N_2842,N_2956);
and UO_113 (O_113,N_2916,N_2958);
nand UO_114 (O_114,N_2573,N_2721);
nor UO_115 (O_115,N_2337,N_2878);
or UO_116 (O_116,N_2579,N_2813);
nand UO_117 (O_117,N_2868,N_2928);
and UO_118 (O_118,N_2801,N_2647);
xor UO_119 (O_119,N_2720,N_2905);
and UO_120 (O_120,N_2770,N_2754);
and UO_121 (O_121,N_2722,N_2289);
or UO_122 (O_122,N_2306,N_2944);
nand UO_123 (O_123,N_2894,N_2461);
nor UO_124 (O_124,N_2536,N_2393);
or UO_125 (O_125,N_2483,N_2695);
nor UO_126 (O_126,N_2663,N_2506);
nand UO_127 (O_127,N_2269,N_2378);
nand UO_128 (O_128,N_2356,N_2600);
nand UO_129 (O_129,N_2940,N_2984);
nor UO_130 (O_130,N_2354,N_2547);
or UO_131 (O_131,N_2328,N_2468);
nand UO_132 (O_132,N_2643,N_2477);
or UO_133 (O_133,N_2622,N_2734);
and UO_134 (O_134,N_2499,N_2696);
or UO_135 (O_135,N_2661,N_2298);
nand UO_136 (O_136,N_2290,N_2717);
nand UO_137 (O_137,N_2562,N_2532);
or UO_138 (O_138,N_2932,N_2278);
and UO_139 (O_139,N_2342,N_2785);
nand UO_140 (O_140,N_2346,N_2851);
nand UO_141 (O_141,N_2698,N_2360);
nor UO_142 (O_142,N_2531,N_2953);
or UO_143 (O_143,N_2565,N_2616);
or UO_144 (O_144,N_2911,N_2479);
nor UO_145 (O_145,N_2409,N_2808);
nand UO_146 (O_146,N_2880,N_2769);
nand UO_147 (O_147,N_2816,N_2447);
and UO_148 (O_148,N_2618,N_2558);
or UO_149 (O_149,N_2728,N_2560);
nand UO_150 (O_150,N_2747,N_2471);
nand UO_151 (O_151,N_2528,N_2980);
nor UO_152 (O_152,N_2753,N_2443);
nand UO_153 (O_153,N_2985,N_2974);
nand UO_154 (O_154,N_2649,N_2725);
nor UO_155 (O_155,N_2677,N_2438);
and UO_156 (O_156,N_2831,N_2624);
and UO_157 (O_157,N_2755,N_2373);
and UO_158 (O_158,N_2365,N_2396);
nor UO_159 (O_159,N_2904,N_2970);
and UO_160 (O_160,N_2604,N_2833);
and UO_161 (O_161,N_2301,N_2699);
nor UO_162 (O_162,N_2348,N_2906);
nand UO_163 (O_163,N_2826,N_2584);
or UO_164 (O_164,N_2883,N_2781);
nand UO_165 (O_165,N_2790,N_2784);
nand UO_166 (O_166,N_2996,N_2645);
or UO_167 (O_167,N_2433,N_2332);
and UO_168 (O_168,N_2976,N_2417);
and UO_169 (O_169,N_2617,N_2827);
or UO_170 (O_170,N_2783,N_2933);
or UO_171 (O_171,N_2665,N_2256);
nand UO_172 (O_172,N_2947,N_2388);
or UO_173 (O_173,N_2684,N_2669);
nand UO_174 (O_174,N_2524,N_2987);
nor UO_175 (O_175,N_2945,N_2594);
or UO_176 (O_176,N_2839,N_2563);
and UO_177 (O_177,N_2678,N_2327);
xnor UO_178 (O_178,N_2702,N_2719);
nor UO_179 (O_179,N_2990,N_2310);
and UO_180 (O_180,N_2750,N_2284);
and UO_181 (O_181,N_2825,N_2637);
nor UO_182 (O_182,N_2641,N_2796);
nand UO_183 (O_183,N_2556,N_2731);
or UO_184 (O_184,N_2621,N_2530);
and UO_185 (O_185,N_2606,N_2859);
nor UO_186 (O_186,N_2260,N_2930);
nor UO_187 (O_187,N_2653,N_2862);
or UO_188 (O_188,N_2474,N_2456);
nand UO_189 (O_189,N_2427,N_2807);
nor UO_190 (O_190,N_2762,N_2657);
and UO_191 (O_191,N_2480,N_2585);
nor UO_192 (O_192,N_2897,N_2514);
nor UO_193 (O_193,N_2401,N_2557);
or UO_194 (O_194,N_2598,N_2420);
nand UO_195 (O_195,N_2593,N_2913);
and UO_196 (O_196,N_2297,N_2835);
nand UO_197 (O_197,N_2268,N_2395);
nor UO_198 (O_198,N_2338,N_2330);
or UO_199 (O_199,N_2692,N_2457);
or UO_200 (O_200,N_2441,N_2711);
nor UO_201 (O_201,N_2448,N_2267);
nor UO_202 (O_202,N_2861,N_2476);
nand UO_203 (O_203,N_2659,N_2739);
nor UO_204 (O_204,N_2992,N_2542);
and UO_205 (O_205,N_2772,N_2820);
nor UO_206 (O_206,N_2467,N_2818);
and UO_207 (O_207,N_2574,N_2449);
and UO_208 (O_208,N_2418,N_2946);
nand UO_209 (O_209,N_2282,N_2597);
or UO_210 (O_210,N_2708,N_2798);
or UO_211 (O_211,N_2896,N_2794);
nand UO_212 (O_212,N_2387,N_2602);
and UO_213 (O_213,N_2782,N_2252);
nand UO_214 (O_214,N_2824,N_2361);
nand UO_215 (O_215,N_2630,N_2989);
nor UO_216 (O_216,N_2553,N_2492);
nand UO_217 (O_217,N_2607,N_2408);
nand UO_218 (O_218,N_2482,N_2849);
nand UO_219 (O_219,N_2265,N_2389);
nand UO_220 (O_220,N_2321,N_2667);
and UO_221 (O_221,N_2909,N_2957);
and UO_222 (O_222,N_2505,N_2812);
nor UO_223 (O_223,N_2682,N_2662);
nand UO_224 (O_224,N_2516,N_2701);
nor UO_225 (O_225,N_2644,N_2364);
or UO_226 (O_226,N_2726,N_2982);
or UO_227 (O_227,N_2884,N_2414);
nor UO_228 (O_228,N_2437,N_2968);
nand UO_229 (O_229,N_2279,N_2629);
and UO_230 (O_230,N_2672,N_2704);
or UO_231 (O_231,N_2426,N_2761);
nor UO_232 (O_232,N_2411,N_2727);
nand UO_233 (O_233,N_2280,N_2951);
and UO_234 (O_234,N_2967,N_2960);
and UO_235 (O_235,N_2379,N_2658);
nor UO_236 (O_236,N_2978,N_2660);
and UO_237 (O_237,N_2765,N_2351);
nand UO_238 (O_238,N_2493,N_2941);
nor UO_239 (O_239,N_2362,N_2899);
nor UO_240 (O_240,N_2317,N_2690);
nand UO_241 (O_241,N_2742,N_2440);
and UO_242 (O_242,N_2498,N_2294);
or UO_243 (O_243,N_2623,N_2854);
nand UO_244 (O_244,N_2683,N_2329);
nand UO_245 (O_245,N_2582,N_2881);
nor UO_246 (O_246,N_2981,N_2255);
nor UO_247 (O_247,N_2504,N_2259);
nand UO_248 (O_248,N_2846,N_2533);
nor UO_249 (O_249,N_2797,N_2451);
nand UO_250 (O_250,N_2771,N_2925);
and UO_251 (O_251,N_2738,N_2288);
or UO_252 (O_252,N_2535,N_2634);
nand UO_253 (O_253,N_2655,N_2587);
nor UO_254 (O_254,N_2559,N_2710);
or UO_255 (O_255,N_2455,N_2478);
nand UO_256 (O_256,N_2261,N_2994);
nor UO_257 (O_257,N_2258,N_2703);
and UO_258 (O_258,N_2705,N_2503);
nor UO_259 (O_259,N_2879,N_2921);
nand UO_260 (O_260,N_2266,N_2484);
or UO_261 (O_261,N_2652,N_2285);
and UO_262 (O_262,N_2519,N_2517);
nor UO_263 (O_263,N_2977,N_2809);
nand UO_264 (O_264,N_2640,N_2340);
and UO_265 (O_265,N_2315,N_2995);
nor UO_266 (O_266,N_2459,N_2472);
or UO_267 (O_267,N_2901,N_2380);
and UO_268 (O_268,N_2341,N_2371);
nor UO_269 (O_269,N_2307,N_2520);
and UO_270 (O_270,N_2749,N_2803);
or UO_271 (O_271,N_2694,N_2567);
or UO_272 (O_272,N_2740,N_2745);
and UO_273 (O_273,N_2834,N_2723);
nand UO_274 (O_274,N_2253,N_2281);
and UO_275 (O_275,N_2632,N_2671);
or UO_276 (O_276,N_2283,N_2971);
nor UO_277 (O_277,N_2666,N_2999);
and UO_278 (O_278,N_2639,N_2615);
and UO_279 (O_279,N_2424,N_2948);
and UO_280 (O_280,N_2857,N_2549);
and UO_281 (O_281,N_2760,N_2344);
and UO_282 (O_282,N_2756,N_2377);
and UO_283 (O_283,N_2500,N_2795);
nor UO_284 (O_284,N_2277,N_2347);
nand UO_285 (O_285,N_2900,N_2541);
nand UO_286 (O_286,N_2746,N_2383);
nor UO_287 (O_287,N_2814,N_2917);
and UO_288 (O_288,N_2561,N_2591);
or UO_289 (O_289,N_2805,N_2821);
nand UO_290 (O_290,N_2581,N_2654);
or UO_291 (O_291,N_2675,N_2876);
nand UO_292 (O_292,N_2743,N_2546);
nand UO_293 (O_293,N_2583,N_2822);
or UO_294 (O_294,N_2737,N_2870);
nor UO_295 (O_295,N_2318,N_2515);
nor UO_296 (O_296,N_2871,N_2787);
or UO_297 (O_297,N_2466,N_2421);
or UO_298 (O_298,N_2864,N_2312);
or UO_299 (O_299,N_2759,N_2295);
and UO_300 (O_300,N_2718,N_2855);
and UO_301 (O_301,N_2975,N_2934);
nor UO_302 (O_302,N_2313,N_2308);
nand UO_303 (O_303,N_2303,N_2257);
or UO_304 (O_304,N_2460,N_2810);
nor UO_305 (O_305,N_2320,N_2326);
nand UO_306 (O_306,N_2334,N_2550);
nand UO_307 (O_307,N_2915,N_2815);
and UO_308 (O_308,N_2961,N_2619);
or UO_309 (O_309,N_2458,N_2922);
or UO_310 (O_310,N_2664,N_2997);
nand UO_311 (O_311,N_2952,N_2983);
or UO_312 (O_312,N_2590,N_2425);
nor UO_313 (O_313,N_2465,N_2709);
or UO_314 (O_314,N_2521,N_2697);
nor UO_315 (O_315,N_2764,N_2488);
and UO_316 (O_316,N_2454,N_2434);
nor UO_317 (O_317,N_2481,N_2707);
nand UO_318 (O_318,N_2601,N_2843);
nand UO_319 (O_319,N_2513,N_2823);
or UO_320 (O_320,N_2349,N_2877);
nand UO_321 (O_321,N_2620,N_2507);
nand UO_322 (O_322,N_2626,N_2551);
nand UO_323 (O_323,N_2895,N_2350);
or UO_324 (O_324,N_2273,N_2263);
nand UO_325 (O_325,N_2405,N_2674);
nand UO_326 (O_326,N_2250,N_2331);
or UO_327 (O_327,N_2966,N_2571);
nor UO_328 (O_328,N_2628,N_2577);
or UO_329 (O_329,N_2850,N_2592);
nor UO_330 (O_330,N_2589,N_2681);
nor UO_331 (O_331,N_2670,N_2264);
nor UO_332 (O_332,N_2529,N_2673);
and UO_333 (O_333,N_2271,N_2845);
or UO_334 (O_334,N_2304,N_2939);
or UO_335 (O_335,N_2357,N_2372);
or UO_336 (O_336,N_2596,N_2512);
nor UO_337 (O_337,N_2751,N_2576);
nand UO_338 (O_338,N_2415,N_2631);
nand UO_339 (O_339,N_2552,N_2979);
nor UO_340 (O_340,N_2599,N_2613);
nand UO_341 (O_341,N_2511,N_2486);
nor UO_342 (O_342,N_2733,N_2335);
and UO_343 (O_343,N_2422,N_2508);
and UO_344 (O_344,N_2865,N_2323);
nor UO_345 (O_345,N_2588,N_2688);
nor UO_346 (O_346,N_2391,N_2789);
nor UO_347 (O_347,N_2627,N_2325);
and UO_348 (O_348,N_2509,N_2891);
nor UO_349 (O_349,N_2526,N_2882);
nand UO_350 (O_350,N_2838,N_2919);
nand UO_351 (O_351,N_2286,N_2539);
and UO_352 (O_352,N_2638,N_2679);
nand UO_353 (O_353,N_2376,N_2685);
or UO_354 (O_354,N_2998,N_2262);
or UO_355 (O_355,N_2416,N_2954);
or UO_356 (O_356,N_2943,N_2450);
nand UO_357 (O_357,N_2475,N_2735);
nand UO_358 (O_358,N_2689,N_2715);
and UO_359 (O_359,N_2757,N_2570);
and UO_360 (O_360,N_2767,N_2445);
or UO_361 (O_361,N_2819,N_2832);
nand UO_362 (O_362,N_2603,N_2752);
nand UO_363 (O_363,N_2336,N_2578);
and UO_364 (O_364,N_2991,N_2766);
or UO_365 (O_365,N_2988,N_2291);
nor UO_366 (O_366,N_2302,N_2763);
nand UO_367 (O_367,N_2390,N_2429);
or UO_368 (O_368,N_2314,N_2889);
and UO_369 (O_369,N_2614,N_2802);
or UO_370 (O_370,N_2452,N_2950);
nand UO_371 (O_371,N_2540,N_2251);
nand UO_372 (O_372,N_2860,N_2385);
nor UO_373 (O_373,N_2491,N_2363);
or UO_374 (O_374,N_2799,N_2525);
and UO_375 (O_375,N_2322,N_2992);
nor UO_376 (O_376,N_2670,N_2376);
and UO_377 (O_377,N_2894,N_2560);
nand UO_378 (O_378,N_2333,N_2809);
nand UO_379 (O_379,N_2530,N_2636);
nand UO_380 (O_380,N_2425,N_2353);
or UO_381 (O_381,N_2395,N_2507);
and UO_382 (O_382,N_2968,N_2518);
nand UO_383 (O_383,N_2978,N_2439);
and UO_384 (O_384,N_2814,N_2534);
nor UO_385 (O_385,N_2880,N_2998);
nor UO_386 (O_386,N_2547,N_2416);
nor UO_387 (O_387,N_2921,N_2835);
nor UO_388 (O_388,N_2948,N_2684);
nand UO_389 (O_389,N_2941,N_2520);
nor UO_390 (O_390,N_2374,N_2688);
nor UO_391 (O_391,N_2620,N_2710);
and UO_392 (O_392,N_2579,N_2708);
nand UO_393 (O_393,N_2270,N_2822);
or UO_394 (O_394,N_2354,N_2631);
or UO_395 (O_395,N_2756,N_2626);
and UO_396 (O_396,N_2761,N_2412);
or UO_397 (O_397,N_2690,N_2469);
nor UO_398 (O_398,N_2314,N_2919);
or UO_399 (O_399,N_2604,N_2470);
and UO_400 (O_400,N_2947,N_2408);
and UO_401 (O_401,N_2739,N_2872);
or UO_402 (O_402,N_2734,N_2337);
or UO_403 (O_403,N_2856,N_2737);
and UO_404 (O_404,N_2283,N_2302);
or UO_405 (O_405,N_2617,N_2673);
nand UO_406 (O_406,N_2251,N_2668);
or UO_407 (O_407,N_2975,N_2292);
xnor UO_408 (O_408,N_2842,N_2657);
and UO_409 (O_409,N_2413,N_2340);
nand UO_410 (O_410,N_2742,N_2341);
or UO_411 (O_411,N_2479,N_2509);
nor UO_412 (O_412,N_2997,N_2407);
nor UO_413 (O_413,N_2782,N_2376);
nor UO_414 (O_414,N_2261,N_2521);
nor UO_415 (O_415,N_2964,N_2973);
nand UO_416 (O_416,N_2505,N_2621);
and UO_417 (O_417,N_2344,N_2289);
and UO_418 (O_418,N_2937,N_2634);
nand UO_419 (O_419,N_2335,N_2847);
and UO_420 (O_420,N_2475,N_2317);
or UO_421 (O_421,N_2687,N_2485);
nor UO_422 (O_422,N_2858,N_2626);
and UO_423 (O_423,N_2639,N_2772);
and UO_424 (O_424,N_2883,N_2274);
or UO_425 (O_425,N_2393,N_2915);
nor UO_426 (O_426,N_2532,N_2963);
and UO_427 (O_427,N_2579,N_2544);
and UO_428 (O_428,N_2302,N_2270);
or UO_429 (O_429,N_2501,N_2754);
nand UO_430 (O_430,N_2620,N_2821);
and UO_431 (O_431,N_2527,N_2801);
and UO_432 (O_432,N_2643,N_2824);
nor UO_433 (O_433,N_2784,N_2961);
nand UO_434 (O_434,N_2908,N_2692);
and UO_435 (O_435,N_2853,N_2326);
and UO_436 (O_436,N_2811,N_2937);
or UO_437 (O_437,N_2428,N_2565);
nor UO_438 (O_438,N_2790,N_2950);
and UO_439 (O_439,N_2932,N_2513);
nand UO_440 (O_440,N_2988,N_2379);
nor UO_441 (O_441,N_2272,N_2617);
nand UO_442 (O_442,N_2754,N_2333);
and UO_443 (O_443,N_2984,N_2858);
and UO_444 (O_444,N_2367,N_2327);
nor UO_445 (O_445,N_2587,N_2929);
nor UO_446 (O_446,N_2853,N_2907);
and UO_447 (O_447,N_2602,N_2870);
nor UO_448 (O_448,N_2662,N_2644);
and UO_449 (O_449,N_2724,N_2317);
nand UO_450 (O_450,N_2691,N_2798);
nor UO_451 (O_451,N_2450,N_2472);
or UO_452 (O_452,N_2506,N_2320);
or UO_453 (O_453,N_2275,N_2655);
nand UO_454 (O_454,N_2289,N_2675);
or UO_455 (O_455,N_2954,N_2588);
nor UO_456 (O_456,N_2854,N_2794);
nand UO_457 (O_457,N_2264,N_2444);
nand UO_458 (O_458,N_2417,N_2574);
nor UO_459 (O_459,N_2300,N_2666);
or UO_460 (O_460,N_2870,N_2449);
and UO_461 (O_461,N_2279,N_2705);
or UO_462 (O_462,N_2874,N_2471);
or UO_463 (O_463,N_2618,N_2976);
nor UO_464 (O_464,N_2647,N_2298);
or UO_465 (O_465,N_2298,N_2890);
nor UO_466 (O_466,N_2357,N_2689);
xor UO_467 (O_467,N_2503,N_2425);
nor UO_468 (O_468,N_2672,N_2899);
or UO_469 (O_469,N_2452,N_2312);
nor UO_470 (O_470,N_2890,N_2742);
nor UO_471 (O_471,N_2343,N_2675);
or UO_472 (O_472,N_2455,N_2985);
nor UO_473 (O_473,N_2541,N_2831);
nor UO_474 (O_474,N_2329,N_2502);
nor UO_475 (O_475,N_2285,N_2866);
nand UO_476 (O_476,N_2419,N_2294);
or UO_477 (O_477,N_2861,N_2343);
and UO_478 (O_478,N_2654,N_2349);
nand UO_479 (O_479,N_2387,N_2331);
and UO_480 (O_480,N_2581,N_2415);
nor UO_481 (O_481,N_2895,N_2640);
or UO_482 (O_482,N_2790,N_2775);
and UO_483 (O_483,N_2944,N_2826);
and UO_484 (O_484,N_2518,N_2321);
nand UO_485 (O_485,N_2574,N_2359);
nand UO_486 (O_486,N_2522,N_2804);
nor UO_487 (O_487,N_2376,N_2902);
and UO_488 (O_488,N_2881,N_2967);
nor UO_489 (O_489,N_2268,N_2482);
nand UO_490 (O_490,N_2708,N_2403);
nand UO_491 (O_491,N_2350,N_2945);
nand UO_492 (O_492,N_2291,N_2310);
and UO_493 (O_493,N_2705,N_2807);
nand UO_494 (O_494,N_2573,N_2807);
nand UO_495 (O_495,N_2538,N_2817);
nor UO_496 (O_496,N_2943,N_2335);
nor UO_497 (O_497,N_2878,N_2745);
or UO_498 (O_498,N_2365,N_2250);
and UO_499 (O_499,N_2892,N_2774);
endmodule