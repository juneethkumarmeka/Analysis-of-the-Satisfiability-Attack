module basic_1500_15000_2000_30_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_460,In_955);
nand U1 (N_1,In_499,In_599);
or U2 (N_2,In_1485,In_56);
xnor U3 (N_3,In_223,In_1246);
and U4 (N_4,In_1341,In_754);
nand U5 (N_5,In_1271,In_583);
or U6 (N_6,In_119,In_1380);
nand U7 (N_7,In_1188,In_463);
and U8 (N_8,In_769,In_1074);
nand U9 (N_9,In_1263,In_743);
and U10 (N_10,In_71,In_1312);
or U11 (N_11,In_1295,In_932);
and U12 (N_12,In_938,In_778);
nor U13 (N_13,In_1267,In_246);
and U14 (N_14,In_814,In_190);
nor U15 (N_15,In_22,In_103);
nor U16 (N_16,In_594,In_236);
and U17 (N_17,In_1165,In_1107);
nor U18 (N_18,In_189,In_1307);
or U19 (N_19,In_967,In_986);
and U20 (N_20,In_1310,In_588);
nor U21 (N_21,In_1181,In_289);
or U22 (N_22,In_355,In_1000);
or U23 (N_23,In_1477,In_812);
and U24 (N_24,In_603,In_903);
nand U25 (N_25,In_1489,In_653);
and U26 (N_26,In_996,In_1190);
and U27 (N_27,In_1409,In_751);
nor U28 (N_28,In_1261,In_1306);
nand U29 (N_29,In_701,In_447);
nand U30 (N_30,In_529,In_1143);
or U31 (N_31,In_284,In_1138);
nand U32 (N_32,In_712,In_937);
and U33 (N_33,In_893,In_997);
xnor U34 (N_34,In_1134,In_448);
and U35 (N_35,In_477,In_440);
nor U36 (N_36,In_143,In_1493);
and U37 (N_37,In_62,In_979);
nand U38 (N_38,In_241,In_1168);
or U39 (N_39,In_136,In_558);
nand U40 (N_40,In_293,In_641);
xor U41 (N_41,In_395,In_157);
nand U42 (N_42,In_1484,In_1416);
nor U43 (N_43,In_1297,In_930);
nand U44 (N_44,In_1483,In_1226);
xor U45 (N_45,In_1251,In_128);
nand U46 (N_46,In_1137,In_1317);
and U47 (N_47,In_1432,In_584);
or U48 (N_48,In_179,In_753);
or U49 (N_49,In_309,In_580);
and U50 (N_50,In_1050,In_1240);
nor U51 (N_51,In_1058,In_647);
nor U52 (N_52,In_908,In_153);
or U53 (N_53,In_147,In_557);
nor U54 (N_54,In_1196,In_1304);
nor U55 (N_55,In_1334,In_708);
and U56 (N_56,In_44,In_474);
or U57 (N_57,In_631,In_1055);
xnor U58 (N_58,In_1260,In_634);
nand U59 (N_59,In_679,In_678);
nand U60 (N_60,In_1346,In_1252);
nand U61 (N_61,In_418,In_97);
xnor U62 (N_62,In_1434,In_1017);
nor U63 (N_63,In_1289,In_670);
and U64 (N_64,In_855,In_1335);
nand U65 (N_65,In_59,In_135);
or U66 (N_66,In_1407,In_628);
xnor U67 (N_67,In_1216,In_704);
nand U68 (N_68,In_363,In_951);
xnor U69 (N_69,In_184,In_1418);
nor U70 (N_70,In_1343,In_734);
or U71 (N_71,In_1466,In_1440);
nor U72 (N_72,In_799,In_315);
xnor U73 (N_73,In_1233,In_816);
xnor U74 (N_74,In_655,In_795);
and U75 (N_75,In_1430,In_1047);
or U76 (N_76,In_919,In_430);
or U77 (N_77,In_498,In_64);
or U78 (N_78,In_493,In_632);
nand U79 (N_79,In_569,In_730);
nand U80 (N_80,In_1098,In_74);
nand U81 (N_81,In_702,In_526);
nor U82 (N_82,In_695,In_1223);
nor U83 (N_83,In_683,In_784);
xnor U84 (N_84,In_1090,In_1109);
or U85 (N_85,In_619,In_1102);
nor U86 (N_86,In_1243,In_544);
or U87 (N_87,In_456,In_661);
nand U88 (N_88,In_0,In_70);
or U89 (N_89,In_694,In_706);
nor U90 (N_90,In_481,In_1482);
nor U91 (N_91,In_860,In_509);
and U92 (N_92,In_1202,In_643);
xor U93 (N_93,In_332,In_212);
xnor U94 (N_94,In_671,In_335);
nand U95 (N_95,In_1395,In_100);
and U96 (N_96,In_608,In_791);
and U97 (N_97,In_1139,In_65);
or U98 (N_98,In_707,In_1420);
or U99 (N_99,In_1149,In_394);
and U100 (N_100,In_1160,In_371);
and U101 (N_101,In_1285,In_1022);
nand U102 (N_102,In_566,In_487);
nor U103 (N_103,In_1378,In_843);
nor U104 (N_104,In_361,In_1305);
nand U105 (N_105,In_271,In_765);
or U106 (N_106,In_16,In_1488);
nor U107 (N_107,In_862,In_453);
or U108 (N_108,In_519,In_1377);
nor U109 (N_109,In_1023,In_1433);
and U110 (N_110,In_177,In_251);
nor U111 (N_111,In_1207,In_727);
nor U112 (N_112,In_372,In_1172);
or U113 (N_113,In_299,In_504);
nor U114 (N_114,In_1257,In_102);
or U115 (N_115,In_1414,In_160);
nor U116 (N_116,In_1281,In_344);
and U117 (N_117,In_1401,In_1481);
or U118 (N_118,In_1259,In_113);
nor U119 (N_119,In_181,In_1410);
and U120 (N_120,In_1024,In_195);
or U121 (N_121,In_1099,In_749);
nand U122 (N_122,In_947,In_773);
nand U123 (N_123,In_384,In_449);
or U124 (N_124,In_388,In_1062);
nand U125 (N_125,In_970,In_601);
or U126 (N_126,In_78,In_736);
and U127 (N_127,In_85,In_1372);
nand U128 (N_128,In_870,In_511);
nand U129 (N_129,In_1404,In_1179);
nand U130 (N_130,In_681,In_1120);
and U131 (N_131,In_374,In_971);
nor U132 (N_132,In_120,In_1136);
nor U133 (N_133,In_1486,In_1406);
and U134 (N_134,In_972,In_609);
and U135 (N_135,In_1332,In_851);
nand U136 (N_136,In_1490,In_370);
and U137 (N_137,In_1464,In_15);
and U138 (N_138,In_911,In_572);
nor U139 (N_139,In_1158,In_890);
nor U140 (N_140,In_1326,In_775);
nor U141 (N_141,In_1142,In_1135);
nor U142 (N_142,In_1122,In_494);
or U143 (N_143,In_396,In_7);
nand U144 (N_144,In_1412,In_1431);
and U145 (N_145,In_1105,In_1044);
nor U146 (N_146,In_35,In_1153);
and U147 (N_147,In_1316,In_338);
nor U148 (N_148,In_1474,In_770);
or U149 (N_149,In_469,In_148);
nand U150 (N_150,In_127,In_1092);
or U151 (N_151,In_484,In_693);
or U152 (N_152,In_1319,In_222);
or U153 (N_153,In_1428,In_151);
nor U154 (N_154,In_844,In_443);
and U155 (N_155,In_1364,In_1290);
and U156 (N_156,In_1163,In_464);
and U157 (N_157,In_1441,In_1070);
nor U158 (N_158,In_316,In_1169);
or U159 (N_159,In_1480,In_400);
or U160 (N_160,In_1390,In_403);
and U161 (N_161,In_774,In_1133);
xnor U162 (N_162,In_1038,In_571);
nor U163 (N_163,In_660,In_605);
and U164 (N_164,In_386,In_1444);
nor U165 (N_165,In_506,In_1187);
or U166 (N_166,In_760,In_427);
nor U167 (N_167,In_573,In_146);
nor U168 (N_168,In_772,In_854);
xnor U169 (N_169,In_429,In_815);
and U170 (N_170,In_1173,In_1167);
nand U171 (N_171,In_1497,In_729);
xor U172 (N_172,In_959,In_404);
and U173 (N_173,In_436,In_1104);
and U174 (N_174,In_393,In_883);
nor U175 (N_175,In_1039,In_1438);
and U176 (N_176,In_1358,In_607);
or U177 (N_177,In_901,In_822);
nor U178 (N_178,In_1119,In_1094);
or U179 (N_179,In_1209,In_1427);
xor U180 (N_180,In_61,In_648);
nand U181 (N_181,In_1132,In_204);
xor U182 (N_182,In_672,In_629);
and U183 (N_183,In_360,In_806);
and U184 (N_184,In_1494,In_999);
or U185 (N_185,In_1291,In_907);
and U186 (N_186,In_1386,In_516);
and U187 (N_187,In_1191,In_615);
and U188 (N_188,In_1336,In_644);
and U189 (N_189,In_1029,In_1303);
nand U190 (N_190,In_483,In_140);
nor U191 (N_191,In_1415,In_96);
nor U192 (N_192,In_534,In_423);
or U193 (N_193,In_902,In_824);
and U194 (N_194,In_383,In_688);
or U195 (N_195,In_894,In_1073);
xnor U196 (N_196,In_1126,In_802);
or U197 (N_197,In_412,In_538);
or U198 (N_198,In_542,In_1349);
nor U199 (N_199,In_662,In_548);
and U200 (N_200,In_921,In_1324);
xor U201 (N_201,In_820,In_718);
nand U202 (N_202,In_45,In_1200);
nand U203 (N_203,In_827,In_742);
and U204 (N_204,In_776,In_1338);
nor U205 (N_205,In_726,In_1076);
and U206 (N_206,In_459,In_1183);
xnor U207 (N_207,In_1159,In_1046);
nor U208 (N_208,In_658,In_111);
or U209 (N_209,In_1387,In_1091);
or U210 (N_210,In_788,In_1476);
nor U211 (N_211,In_1048,In_748);
nor U212 (N_212,In_790,In_848);
and U213 (N_213,In_507,In_831);
and U214 (N_214,In_130,In_89);
nor U215 (N_215,In_771,In_20);
nand U216 (N_216,In_968,In_438);
and U217 (N_217,In_1473,In_166);
nor U218 (N_218,In_1041,In_1366);
nor U219 (N_219,In_684,In_207);
nand U220 (N_220,In_1337,In_1175);
xnor U221 (N_221,In_900,In_275);
nor U222 (N_222,In_431,In_203);
nor U223 (N_223,In_735,In_1237);
nand U224 (N_224,In_437,In_666);
xnor U225 (N_225,In_547,In_406);
xor U226 (N_226,In_164,In_1388);
xor U227 (N_227,In_1061,In_191);
nand U228 (N_228,In_523,In_110);
nand U229 (N_229,In_1330,In_1156);
or U230 (N_230,In_837,In_874);
nor U231 (N_231,In_624,In_37);
or U232 (N_232,In_1286,In_556);
nand U233 (N_233,In_1262,In_40);
or U234 (N_234,In_1154,In_918);
and U235 (N_235,In_1193,In_485);
nor U236 (N_236,In_257,In_692);
or U237 (N_237,In_1006,In_1278);
and U238 (N_238,In_966,In_23);
nor U239 (N_239,In_1323,In_1370);
or U240 (N_240,In_6,In_479);
and U241 (N_241,In_528,In_243);
nand U242 (N_242,In_1322,In_1342);
nand U243 (N_243,In_1315,In_280);
or U244 (N_244,In_336,In_1195);
and U245 (N_245,In_1115,In_1491);
nor U246 (N_246,In_1344,In_1405);
or U247 (N_247,In_567,In_869);
nor U248 (N_248,In_1222,In_537);
and U249 (N_249,In_656,In_1421);
nand U250 (N_250,In_623,In_1462);
nand U251 (N_251,In_746,In_413);
nand U252 (N_252,In_109,In_1081);
nor U253 (N_253,In_709,In_645);
nor U254 (N_254,In_1258,In_1273);
nor U255 (N_255,In_940,In_800);
nor U256 (N_256,In_1066,In_1340);
nand U257 (N_257,In_321,In_410);
xor U258 (N_258,In_324,In_1383);
nand U259 (N_259,In_86,In_1247);
and U260 (N_260,In_905,In_333);
nand U261 (N_261,In_1446,In_347);
nand U262 (N_262,In_156,In_1220);
nand U263 (N_263,In_714,In_287);
or U264 (N_264,In_1368,In_115);
and U265 (N_265,In_180,In_737);
nand U266 (N_266,In_1253,In_1314);
xnor U267 (N_267,In_107,In_741);
nor U268 (N_268,In_1455,In_131);
or U269 (N_269,In_221,In_31);
and U270 (N_270,In_554,In_540);
or U271 (N_271,In_175,In_1208);
xnor U272 (N_272,In_781,In_1425);
and U273 (N_273,In_1363,In_2);
and U274 (N_274,In_432,In_1284);
or U275 (N_275,In_1325,In_270);
or U276 (N_276,In_421,In_382);
nor U277 (N_277,In_1351,In_250);
nor U278 (N_278,In_1205,In_733);
or U279 (N_279,In_1032,In_873);
or U280 (N_280,In_724,In_878);
or U281 (N_281,In_428,In_1020);
or U282 (N_282,In_941,In_486);
xnor U283 (N_283,In_1096,In_1472);
nor U284 (N_284,In_740,In_444);
and U285 (N_285,In_3,In_398);
or U286 (N_286,In_43,In_777);
nor U287 (N_287,In_810,In_1007);
nand U288 (N_288,In_1011,In_232);
and U289 (N_289,In_452,In_864);
nand U290 (N_290,In_904,In_272);
or U291 (N_291,In_1111,In_466);
xor U292 (N_292,In_357,In_291);
xnor U293 (N_293,In_665,In_24);
and U294 (N_294,In_57,In_1225);
or U295 (N_295,In_260,In_916);
and U296 (N_296,In_622,In_1460);
xnor U297 (N_297,In_1113,In_297);
or U298 (N_298,In_1034,In_269);
and U299 (N_299,In_636,In_351);
or U300 (N_300,In_134,In_14);
nor U301 (N_301,In_1492,In_419);
xor U302 (N_302,In_168,In_705);
nor U303 (N_303,In_1069,In_1054);
nand U304 (N_304,In_762,In_1308);
and U305 (N_305,In_314,In_1221);
or U306 (N_306,In_104,In_885);
nand U307 (N_307,In_652,In_1013);
nor U308 (N_308,In_301,In_687);
nor U309 (N_309,In_1461,In_1213);
nor U310 (N_310,In_1059,In_1277);
or U311 (N_311,In_1382,In_876);
xor U312 (N_312,In_892,In_350);
nor U313 (N_313,In_161,In_501);
nand U314 (N_314,In_353,In_711);
nand U315 (N_315,In_1052,In_9);
nor U316 (N_316,In_989,In_171);
xor U317 (N_317,In_359,In_294);
and U318 (N_318,In_473,In_1043);
or U319 (N_319,In_285,In_305);
nor U320 (N_320,In_924,In_721);
nor U321 (N_321,In_958,In_266);
nor U322 (N_322,In_1176,In_974);
nor U323 (N_323,In_1385,In_560);
and U324 (N_324,In_41,In_1311);
nor U325 (N_325,In_1174,In_1235);
nand U326 (N_326,In_1203,In_201);
nand U327 (N_327,In_682,In_896);
nor U328 (N_328,In_1309,In_183);
and U329 (N_329,In_1117,In_302);
and U330 (N_330,In_1384,In_227);
and U331 (N_331,In_1140,In_833);
xnor U332 (N_332,In_1033,In_1301);
nand U333 (N_333,In_123,In_1009);
or U334 (N_334,In_719,In_1199);
nand U335 (N_335,In_10,In_492);
xnor U336 (N_336,In_1145,In_1361);
and U337 (N_337,In_206,In_1180);
nor U338 (N_338,In_318,In_633);
nor U339 (N_339,In_818,In_377);
nor U340 (N_340,In_186,In_1238);
xnor U341 (N_341,In_759,In_376);
or U342 (N_342,In_87,In_317);
nand U343 (N_343,In_764,In_155);
and U344 (N_344,In_756,In_1411);
nand U345 (N_345,In_879,In_998);
or U346 (N_346,In_984,In_1211);
xnor U347 (N_347,In_245,In_1030);
nor U348 (N_348,In_458,In_929);
nor U349 (N_349,In_461,In_1391);
and U350 (N_350,In_913,In_1178);
and U351 (N_351,In_165,In_259);
nor U352 (N_352,In_789,In_530);
nand U353 (N_353,In_574,In_1345);
and U354 (N_354,In_320,In_1272);
nor U355 (N_355,In_72,In_988);
or U356 (N_356,In_262,In_1302);
nor U357 (N_357,In_1450,In_193);
nor U358 (N_358,In_1467,In_365);
nand U359 (N_359,In_821,In_792);
nand U360 (N_360,In_239,In_1212);
nor U361 (N_361,In_322,In_1083);
xor U362 (N_362,In_1292,In_1078);
xor U363 (N_363,In_1085,In_1114);
nor U364 (N_364,In_17,In_1242);
nand U365 (N_365,In_1177,In_53);
or U366 (N_366,In_496,In_1417);
nor U367 (N_367,In_312,In_308);
or U368 (N_368,In_1400,In_1360);
nor U369 (N_369,In_793,In_829);
nand U370 (N_370,In_1454,In_337);
nand U371 (N_371,In_1451,In_553);
nor U372 (N_372,In_228,In_1164);
xnor U373 (N_373,In_597,In_216);
nor U374 (N_374,In_639,In_875);
and U375 (N_375,In_373,In_1146);
or U376 (N_376,In_490,In_1356);
nand U377 (N_377,In_48,In_1331);
and U378 (N_378,In_564,In_539);
and U379 (N_379,In_1230,In_578);
or U380 (N_380,In_273,In_887);
or U381 (N_381,In_731,In_68);
nand U382 (N_382,In_1125,In_853);
xor U383 (N_383,In_981,In_991);
and U384 (N_384,In_313,In_627);
nor U385 (N_385,In_1184,In_367);
nor U386 (N_386,In_238,In_253);
and U387 (N_387,In_1015,In_969);
and U388 (N_388,In_910,In_75);
nand U389 (N_389,In_1131,In_559);
or U390 (N_390,In_1192,In_1014);
and U391 (N_391,In_895,In_1110);
and U392 (N_392,In_994,In_993);
and U393 (N_393,In_422,In_797);
and U394 (N_394,In_150,In_691);
nand U395 (N_395,In_975,In_1496);
nand U396 (N_396,In_1250,In_1171);
and U397 (N_397,In_750,In_1475);
and U398 (N_398,In_390,In_654);
nand U399 (N_399,In_139,In_1287);
nand U400 (N_400,In_1049,In_478);
nand U401 (N_401,In_1270,In_116);
nor U402 (N_402,In_12,In_836);
and U403 (N_403,In_1403,In_214);
and U404 (N_404,In_354,In_163);
xnor U405 (N_405,In_1453,In_328);
nand U406 (N_406,In_828,In_897);
nand U407 (N_407,In_713,In_230);
xnor U408 (N_408,In_1408,In_592);
and U409 (N_409,In_304,In_364);
nand U410 (N_410,In_1274,In_1353);
nand U411 (N_411,In_782,In_39);
or U412 (N_412,In_1328,In_1379);
or U413 (N_413,In_745,In_757);
or U414 (N_414,In_582,In_618);
nor U415 (N_415,In_1027,In_274);
or U416 (N_416,In_1498,In_407);
nor U417 (N_417,In_980,In_1327);
or U418 (N_418,In_761,In_1350);
or U419 (N_419,In_640,In_1352);
nand U420 (N_420,In_915,In_1318);
nand U421 (N_421,In_295,In_1084);
or U422 (N_422,In_1296,In_1123);
and U423 (N_423,In_866,In_149);
and U424 (N_424,In_1419,In_1101);
nand U425 (N_425,In_258,In_1231);
nor U426 (N_426,In_521,In_616);
nor U427 (N_427,In_79,In_524);
nor U428 (N_428,In_861,In_1465);
and U429 (N_429,In_723,In_217);
nor U430 (N_430,In_926,In_300);
nor U431 (N_431,In_1067,In_69);
nor U432 (N_432,In_1201,In_1021);
nor U433 (N_433,In_1320,In_651);
nor U434 (N_434,In_55,In_612);
nor U435 (N_435,In_141,In_489);
xor U436 (N_436,In_669,In_898);
nand U437 (N_437,In_1437,In_249);
or U438 (N_438,In_1264,In_1219);
and U439 (N_439,In_747,In_311);
xnor U440 (N_440,In_132,In_326);
nand U441 (N_441,In_330,In_1227);
and U442 (N_442,In_1280,In_956);
nand U443 (N_443,In_689,In_604);
and U444 (N_444,In_659,In_199);
and U445 (N_445,In_176,In_1002);
or U446 (N_446,In_664,In_495);
nand U447 (N_447,In_935,In_1339);
nand U448 (N_448,In_809,In_767);
nand U449 (N_449,In_783,In_1300);
nand U450 (N_450,In_420,In_699);
xor U451 (N_451,In_933,In_106);
nand U452 (N_452,In_581,In_889);
nand U453 (N_453,In_555,In_167);
and U454 (N_454,In_405,In_1151);
or U455 (N_455,In_1095,In_535);
or U456 (N_456,In_158,In_346);
nand U457 (N_457,In_391,In_81);
and U458 (N_458,In_415,In_948);
nor U459 (N_459,In_804,In_152);
nor U460 (N_460,In_247,In_1127);
nand U461 (N_461,In_345,In_823);
nand U462 (N_462,In_863,In_533);
and U463 (N_463,In_626,In_133);
xor U464 (N_464,In_1072,In_1026);
nor U465 (N_465,In_1255,In_1371);
nor U466 (N_466,In_1008,In_244);
and U467 (N_467,In_1244,In_82);
nor U468 (N_468,In_38,In_1071);
and U469 (N_469,In_595,In_1313);
nor U470 (N_470,In_471,In_210);
or U471 (N_471,In_331,In_482);
xnor U472 (N_472,In_1376,In_198);
or U473 (N_473,In_1116,In_242);
nand U474 (N_474,In_219,In_457);
and U475 (N_475,In_1079,In_42);
and U476 (N_476,In_282,In_596);
nand U477 (N_477,In_579,In_117);
xnor U478 (N_478,In_1001,In_1224);
and U479 (N_479,In_1229,In_568);
nand U480 (N_480,In_976,In_218);
nand U481 (N_481,In_1354,In_196);
nand U482 (N_482,In_953,In_450);
or U483 (N_483,In_1282,In_1161);
xor U484 (N_484,In_550,In_832);
and U485 (N_485,In_235,In_1012);
and U486 (N_486,In_715,In_614);
xor U487 (N_487,In_352,In_1045);
or U488 (N_488,In_1124,In_442);
nand U489 (N_489,In_178,In_1357);
and U490 (N_490,In_1499,In_173);
or U491 (N_491,In_637,In_488);
xnor U492 (N_492,In_66,In_32);
or U493 (N_493,In_19,In_891);
nand U494 (N_494,In_943,In_545);
nor U495 (N_495,In_920,In_26);
nand U496 (N_496,In_475,In_886);
nand U497 (N_497,In_1355,In_392);
nand U498 (N_498,In_142,In_591);
nor U499 (N_499,In_1359,In_1394);
nand U500 (N_500,N_345,In_1194);
or U501 (N_501,N_348,In_1003);
nand U502 (N_502,In_188,In_950);
nor U503 (N_503,N_457,In_1369);
nor U504 (N_504,In_1398,In_752);
and U505 (N_505,N_445,N_341);
nor U506 (N_506,N_4,In_587);
nor U507 (N_507,N_326,In_663);
nor U508 (N_508,N_375,In_497);
xor U509 (N_509,N_449,N_151);
or U510 (N_510,N_67,N_26);
nand U511 (N_511,In_1077,N_300);
nor U512 (N_512,N_158,In_755);
xnor U513 (N_513,In_77,N_5);
and U514 (N_514,N_388,In_5);
or U515 (N_515,In_67,N_132);
and U516 (N_516,In_543,In_18);
nor U517 (N_517,N_135,N_57);
or U518 (N_518,N_70,N_200);
or U519 (N_519,In_1463,In_1087);
and U520 (N_520,N_32,In_1204);
and U521 (N_521,In_716,In_859);
nand U522 (N_522,N_352,N_19);
and U523 (N_523,N_193,In_1035);
and U524 (N_524,N_426,In_1130);
nor U525 (N_525,N_31,N_44);
or U526 (N_526,N_157,N_84);
nor U527 (N_527,In_1080,In_387);
or U528 (N_528,N_337,N_383);
nand U529 (N_529,In_162,In_825);
and U530 (N_530,N_212,In_906);
or U531 (N_531,N_185,In_399);
and U532 (N_532,In_598,In_728);
and U533 (N_533,In_472,In_798);
and U534 (N_534,In_698,In_1298);
and U535 (N_535,N_101,N_374);
nor U536 (N_536,In_1458,N_228);
and U537 (N_537,N_149,N_78);
xor U538 (N_538,In_194,In_1333);
or U539 (N_539,In_1197,In_435);
and U540 (N_540,In_356,N_480);
and U541 (N_541,In_586,In_1396);
xor U542 (N_542,In_613,N_358);
and U543 (N_543,In_341,N_125);
nand U544 (N_544,In_909,N_114);
nor U545 (N_545,In_276,N_233);
xnor U546 (N_546,N_33,In_288);
or U547 (N_547,N_77,In_541);
nand U548 (N_548,N_197,N_203);
or U549 (N_549,N_239,In_794);
nand U550 (N_550,N_387,N_169);
nor U551 (N_551,In_277,N_361);
nand U552 (N_552,In_467,N_258);
xor U553 (N_553,N_418,N_310);
and U554 (N_554,N_397,In_114);
or U555 (N_555,N_21,In_983);
xnor U556 (N_556,N_286,N_376);
nand U557 (N_557,N_188,N_313);
nand U558 (N_558,In_676,N_97);
or U559 (N_559,In_122,In_508);
xor U560 (N_560,In_888,In_620);
and U561 (N_561,N_131,N_141);
or U562 (N_562,N_332,N_398);
and U563 (N_563,N_40,In_368);
and U564 (N_564,In_732,In_434);
nor U565 (N_565,In_197,In_677);
nand U566 (N_566,N_285,In_884);
nand U567 (N_567,N_194,N_400);
nand U568 (N_568,N_325,N_53);
nor U569 (N_569,N_246,In_170);
or U570 (N_570,In_606,In_54);
or U571 (N_571,N_353,In_517);
nand U572 (N_572,In_237,In_1108);
nor U573 (N_573,In_1217,N_349);
nand U574 (N_574,N_408,In_446);
nand U575 (N_575,In_402,In_1299);
or U576 (N_576,In_840,N_218);
nor U577 (N_577,N_92,N_162);
or U578 (N_578,In_995,In_872);
nor U579 (N_579,N_362,N_432);
and U580 (N_580,N_106,In_914);
and U581 (N_581,N_227,In_1106);
or U582 (N_582,N_2,N_304);
or U583 (N_583,N_396,N_223);
or U584 (N_584,N_11,N_458);
or U585 (N_585,N_221,In_455);
or U586 (N_586,In_265,N_461);
nand U587 (N_587,N_459,In_510);
or U588 (N_588,In_1402,In_1060);
and U589 (N_589,In_409,In_1389);
and U590 (N_590,In_1249,N_271);
nor U591 (N_591,N_406,In_625);
nand U592 (N_592,N_253,N_69);
nand U593 (N_593,N_257,N_302);
xor U594 (N_594,N_93,In_73);
or U595 (N_595,In_642,N_45);
and U596 (N_596,In_842,N_10);
nand U597 (N_597,N_421,In_108);
or U598 (N_598,In_84,In_813);
and U599 (N_599,In_381,In_536);
nand U600 (N_600,N_210,N_323);
nand U601 (N_601,N_49,N_455);
and U602 (N_602,N_448,In_899);
nand U603 (N_603,N_235,In_1283);
and U604 (N_604,N_321,N_288);
nor U605 (N_605,N_205,N_399);
nand U606 (N_606,N_184,N_66);
xor U607 (N_607,N_41,In_47);
or U608 (N_608,In_549,In_340);
nand U609 (N_609,In_424,In_1469);
nand U610 (N_610,N_363,In_650);
nor U611 (N_611,N_404,N_198);
nor U612 (N_612,In_965,In_36);
nand U613 (N_613,In_768,In_675);
nand U614 (N_614,In_515,In_1186);
nand U615 (N_615,In_25,In_830);
or U616 (N_616,N_433,In_1215);
or U617 (N_617,N_424,N_122);
or U618 (N_618,N_127,N_120);
or U619 (N_619,N_483,N_307);
xnor U620 (N_620,N_301,N_96);
nand U621 (N_621,N_390,N_168);
xor U622 (N_622,In_1097,N_425);
nand U623 (N_623,N_442,N_278);
nand U624 (N_624,In_1265,In_1198);
or U625 (N_625,In_414,N_75);
nor U626 (N_626,N_306,In_505);
nand U627 (N_627,N_324,N_140);
nor U628 (N_628,N_264,In_454);
or U629 (N_629,N_444,In_1064);
nand U630 (N_630,N_42,In_1443);
nor U631 (N_631,In_1082,In_942);
nor U632 (N_632,In_1445,N_56);
nand U633 (N_633,N_110,N_137);
and U634 (N_634,In_451,N_454);
and U635 (N_635,In_80,N_220);
nor U636 (N_636,In_281,N_378);
nand U637 (N_637,N_136,N_12);
nand U638 (N_638,N_269,In_1189);
or U639 (N_639,In_846,N_208);
nor U640 (N_640,In_1152,N_279);
nor U641 (N_641,In_1275,N_354);
and U642 (N_642,N_466,N_54);
nor U643 (N_643,In_610,In_378);
nor U644 (N_644,N_187,N_86);
nand U645 (N_645,N_266,In_600);
and U646 (N_646,N_3,N_283);
nor U647 (N_647,In_358,N_419);
or U648 (N_648,In_174,N_393);
nand U649 (N_649,N_386,In_1144);
or U650 (N_650,In_101,In_1457);
and U651 (N_651,N_76,In_91);
and U652 (N_652,In_593,N_416);
and U653 (N_653,In_1293,N_477);
nand U654 (N_654,N_402,In_635);
and U655 (N_655,N_417,In_826);
or U656 (N_656,In_306,In_1241);
nand U657 (N_657,In_787,N_366);
nor U658 (N_658,N_292,N_451);
nand U659 (N_659,In_1276,N_71);
and U660 (N_660,In_835,N_335);
nand U661 (N_661,N_290,In_590);
nand U662 (N_662,In_1374,N_117);
nand U663 (N_663,In_99,In_200);
xnor U664 (N_664,In_225,N_103);
nand U665 (N_665,N_344,N_409);
xor U666 (N_666,N_81,N_379);
and U667 (N_667,In_1348,In_118);
nor U668 (N_668,In_1112,In_231);
xor U669 (N_669,In_514,In_1214);
and U670 (N_670,In_520,In_268);
or U671 (N_671,In_339,N_190);
xnor U672 (N_672,N_38,In_657);
nor U673 (N_673,N_265,In_379);
nand U674 (N_674,In_685,N_104);
and U675 (N_675,N_371,N_231);
and U676 (N_676,In_1182,In_310);
nand U677 (N_677,In_264,In_298);
xor U678 (N_678,N_1,N_327);
xnor U679 (N_679,N_145,In_1397);
and U680 (N_680,In_945,In_763);
or U681 (N_681,N_146,N_333);
nand U682 (N_682,N_488,N_452);
nor U683 (N_683,In_856,N_294);
and U684 (N_684,N_360,N_309);
and U685 (N_685,In_858,In_21);
or U686 (N_686,N_238,In_1236);
and U687 (N_687,In_503,N_384);
nor U688 (N_688,N_412,N_394);
or U689 (N_689,In_690,N_315);
and U690 (N_690,N_329,N_119);
and U691 (N_691,In_1468,N_201);
or U692 (N_692,In_95,N_16);
and U693 (N_693,In_577,N_133);
and U694 (N_694,In_60,In_710);
or U695 (N_695,In_1288,In_720);
nand U696 (N_696,N_282,In_1147);
nand U697 (N_697,N_211,In_563);
nor U698 (N_698,In_13,N_144);
nor U699 (N_699,In_852,In_292);
and U700 (N_700,N_217,In_1037);
and U701 (N_701,N_22,In_1367);
or U702 (N_702,In_912,N_389);
and U703 (N_703,N_216,N_256);
nor U704 (N_704,In_849,N_153);
or U705 (N_705,N_474,N_191);
nor U706 (N_706,In_94,In_697);
and U707 (N_707,In_1452,In_226);
nand U708 (N_708,In_255,N_263);
and U709 (N_709,N_90,N_367);
nand U710 (N_710,N_50,N_27);
nand U711 (N_711,In_476,N_165);
and U712 (N_712,N_296,N_202);
nand U713 (N_713,N_34,N_139);
nand U714 (N_714,N_17,In_1166);
and U715 (N_715,In_925,In_575);
nand U716 (N_716,N_160,In_973);
and U717 (N_717,N_475,In_187);
nor U718 (N_718,N_484,In_1429);
and U719 (N_719,N_150,N_413);
and U720 (N_720,In_375,In_290);
xor U721 (N_721,In_502,N_199);
and U722 (N_722,N_155,In_389);
or U723 (N_723,N_450,N_275);
nor U724 (N_724,In_1393,In_1093);
nor U725 (N_725,In_411,N_178);
xnor U726 (N_726,In_936,In_1329);
nor U727 (N_727,N_338,N_443);
or U728 (N_728,In_1157,In_50);
or U729 (N_729,In_192,N_63);
nor U730 (N_730,In_1362,N_303);
nand U731 (N_731,N_317,N_312);
nor U732 (N_732,In_125,N_195);
nor U733 (N_733,In_307,In_680);
and U734 (N_734,In_1248,In_1051);
nor U735 (N_735,In_348,N_368);
xor U736 (N_736,In_939,In_1239);
nor U737 (N_737,N_252,N_147);
and U738 (N_738,In_1065,N_322);
and U739 (N_739,In_252,In_839);
and U740 (N_740,N_245,N_364);
nor U741 (N_741,In_93,N_230);
and U742 (N_742,N_83,N_420);
nor U743 (N_743,N_369,In_725);
nor U744 (N_744,In_1053,N_438);
or U745 (N_745,In_248,In_961);
nand U746 (N_746,In_267,In_240);
nor U747 (N_747,N_95,In_1103);
and U748 (N_748,In_213,In_1075);
or U749 (N_749,N_357,In_808);
nand U750 (N_750,N_112,N_126);
and U751 (N_751,N_196,N_251);
or U752 (N_752,In_1426,In_779);
nand U753 (N_753,N_336,In_1005);
nor U754 (N_754,N_18,N_460);
or U755 (N_755,In_1459,In_185);
nor U756 (N_756,N_249,N_355);
xnor U757 (N_757,N_28,N_89);
or U758 (N_758,In_1004,N_102);
nor U759 (N_759,In_877,In_978);
nand U760 (N_760,In_1399,In_1118);
or U761 (N_761,In_445,In_1042);
or U762 (N_762,In_1162,In_722);
nand U763 (N_763,In_169,N_113);
nor U764 (N_764,N_206,N_318);
and U765 (N_765,N_207,In_425);
nand U766 (N_766,In_1449,N_331);
xor U767 (N_767,In_1019,In_1170);
nor U768 (N_768,In_982,In_985);
nand U769 (N_769,N_43,In_145);
nor U770 (N_770,In_1040,N_308);
nor U771 (N_771,N_260,In_834);
and U772 (N_772,N_172,N_163);
xnor U773 (N_773,In_949,N_213);
and U774 (N_774,In_838,In_1245);
and U775 (N_775,N_61,N_489);
nor U776 (N_776,N_422,N_177);
and U777 (N_777,In_334,In_585);
nor U778 (N_778,In_465,N_35);
nor U779 (N_779,In_931,In_229);
xnor U780 (N_780,N_287,In_1057);
nor U781 (N_781,N_154,In_805);
nand U782 (N_782,N_431,N_343);
and U783 (N_783,N_470,N_250);
nand U784 (N_784,N_129,In_286);
and U785 (N_785,In_1185,In_1294);
or U786 (N_786,In_927,In_881);
or U787 (N_787,In_88,In_977);
nor U788 (N_788,In_11,In_1256);
nand U789 (N_789,N_68,N_274);
nor U790 (N_790,N_224,N_347);
nor U791 (N_791,N_128,In_850);
nor U792 (N_792,N_243,In_1025);
and U793 (N_793,In_686,N_340);
or U794 (N_794,N_237,In_1);
nand U795 (N_795,In_1228,N_365);
nor U796 (N_796,In_527,In_327);
nand U797 (N_797,N_39,In_934);
or U798 (N_798,In_112,In_946);
nand U799 (N_799,In_865,In_92);
nor U800 (N_800,In_646,N_52);
or U801 (N_801,In_532,In_963);
nand U802 (N_802,N_456,N_319);
and U803 (N_803,In_964,In_667);
xor U804 (N_804,In_211,N_65);
nand U805 (N_805,N_330,N_91);
or U806 (N_806,In_1129,N_342);
xor U807 (N_807,In_278,In_1375);
or U808 (N_808,N_118,N_58);
and U809 (N_809,N_62,N_20);
nand U810 (N_810,In_1210,In_63);
and U811 (N_811,In_1088,In_1056);
or U812 (N_812,In_882,N_124);
nand U813 (N_813,In_1155,In_703);
nand U814 (N_814,N_7,In_342);
nand U815 (N_815,N_48,In_738);
nor U816 (N_816,In_923,N_234);
and U817 (N_817,In_868,N_289);
and U818 (N_818,N_94,N_116);
nor U819 (N_819,In_1010,N_247);
and U820 (N_820,N_491,In_233);
xnor U821 (N_821,N_423,In_928);
or U822 (N_822,N_439,In_1148);
or U823 (N_823,In_630,In_992);
or U824 (N_824,N_166,N_204);
and U825 (N_825,In_397,In_917);
or U826 (N_826,N_123,N_430);
and U827 (N_827,N_23,N_293);
nor U828 (N_828,N_464,N_351);
nand U829 (N_829,N_15,In_1365);
and U830 (N_830,In_1268,N_64);
and U831 (N_831,N_175,N_192);
and U832 (N_832,N_407,In_871);
or U833 (N_833,In_1206,In_46);
xor U834 (N_834,In_739,In_462);
nand U835 (N_835,N_280,N_471);
and U836 (N_836,In_649,N_295);
and U837 (N_837,In_1471,In_744);
nand U838 (N_838,In_159,In_1381);
or U839 (N_839,In_34,In_1422);
nand U840 (N_840,N_100,In_780);
nor U841 (N_841,In_990,N_435);
and U842 (N_842,N_105,N_427);
nor U843 (N_843,In_1018,In_785);
nand U844 (N_844,N_30,In_366);
and U845 (N_845,In_385,In_4);
nand U846 (N_846,N_469,N_229);
and U847 (N_847,N_254,In_786);
nand U848 (N_848,N_415,In_1436);
or U849 (N_849,In_441,In_668);
and U850 (N_850,N_180,N_46);
and U851 (N_851,N_380,N_29);
xnor U852 (N_852,In_1128,N_79);
nand U853 (N_853,N_262,In_960);
or U854 (N_854,In_182,In_144);
or U855 (N_855,In_129,N_385);
or U856 (N_856,In_561,N_414);
or U857 (N_857,N_225,N_88);
nand U858 (N_858,N_72,N_121);
nor U859 (N_859,N_182,N_99);
or U860 (N_860,In_1068,N_176);
nor U861 (N_861,N_496,N_284);
or U862 (N_862,In_1063,In_638);
nor U863 (N_863,N_0,In_962);
nor U864 (N_864,In_416,In_329);
xnor U865 (N_865,In_673,In_28);
and U866 (N_866,In_380,In_343);
nand U867 (N_867,In_796,In_674);
and U868 (N_868,In_857,N_219);
nor U869 (N_869,N_391,N_472);
nand U870 (N_870,N_311,In_138);
and U871 (N_871,In_49,In_518);
and U872 (N_872,N_299,N_328);
nor U873 (N_873,N_339,In_261);
xnor U874 (N_874,In_480,N_405);
nand U875 (N_875,In_1373,N_473);
nand U876 (N_876,In_349,N_181);
nor U877 (N_877,N_372,N_268);
nor U878 (N_878,N_261,N_370);
and U879 (N_879,N_51,N_148);
nor U880 (N_880,In_1456,In_1232);
or U881 (N_881,In_602,N_356);
nor U882 (N_882,N_248,N_13);
or U883 (N_883,N_73,N_446);
xnor U884 (N_884,In_215,In_1495);
nand U885 (N_885,In_296,In_1423);
and U886 (N_886,N_60,N_9);
and U887 (N_887,N_495,In_1234);
nand U888 (N_888,N_215,In_408);
nor U889 (N_889,N_236,N_259);
and U890 (N_890,N_437,In_52);
and U891 (N_891,In_1347,N_179);
or U892 (N_892,In_1269,In_1435);
nand U893 (N_893,In_83,In_700);
nor U894 (N_894,N_411,In_90);
or U895 (N_895,In_303,In_512);
nand U896 (N_896,In_433,In_1478);
nand U897 (N_897,In_1086,N_277);
nand U898 (N_898,N_107,In_439);
nor U899 (N_899,N_214,In_766);
nand U900 (N_900,N_109,In_263);
or U901 (N_901,In_208,In_126);
nor U902 (N_902,N_314,N_115);
and U903 (N_903,N_25,N_6);
nor U904 (N_904,In_1031,N_183);
or U905 (N_905,N_47,In_811);
and U906 (N_906,N_174,N_55);
nand U907 (N_907,N_171,In_807);
or U908 (N_908,N_226,N_382);
and U909 (N_909,N_481,In_254);
or U910 (N_910,In_105,N_152);
nand U911 (N_911,N_494,N_142);
and U912 (N_912,N_395,In_1266);
nor U913 (N_913,In_154,N_403);
and U914 (N_914,In_1424,N_320);
and U915 (N_915,N_463,N_130);
xnor U916 (N_916,In_954,In_1479);
nor U917 (N_917,N_453,In_58);
nor U918 (N_918,N_441,N_74);
nor U919 (N_919,In_817,In_417);
and U920 (N_920,N_476,N_487);
xnor U921 (N_921,N_232,N_281);
nor U922 (N_922,N_436,In_803);
or U923 (N_923,In_137,In_845);
nand U924 (N_924,In_717,N_222);
or U925 (N_925,N_359,N_291);
or U926 (N_926,N_161,N_316);
nand U927 (N_927,N_429,In_525);
nand U928 (N_928,N_298,In_1439);
nor U929 (N_929,In_202,In_1036);
nor U930 (N_930,N_462,N_467);
nor U931 (N_931,In_1413,In_551);
nor U932 (N_932,N_485,In_362);
nand U933 (N_933,In_522,N_392);
nor U934 (N_934,N_82,In_546);
nor U935 (N_935,N_241,N_173);
nor U936 (N_936,N_434,N_240);
and U937 (N_937,In_758,In_500);
nand U938 (N_938,In_224,N_346);
nor U939 (N_939,In_51,N_186);
and U940 (N_940,In_801,N_410);
and U941 (N_941,N_272,In_98);
nand U942 (N_942,In_1254,In_880);
or U943 (N_943,In_283,In_1121);
nor U944 (N_944,In_491,In_1448);
or U945 (N_945,N_244,In_8);
nand U946 (N_946,N_209,N_493);
or U947 (N_947,In_944,In_234);
and U948 (N_948,In_33,In_957);
xnor U949 (N_949,N_497,N_98);
and U950 (N_950,N_377,N_350);
nor U951 (N_951,N_428,In_847);
nor U952 (N_952,In_1321,N_170);
nand U953 (N_953,N_87,In_256);
and U954 (N_954,In_841,In_76);
nor U955 (N_955,N_276,In_1016);
or U956 (N_956,In_867,N_111);
nand U957 (N_957,N_270,In_27);
or U958 (N_958,N_498,N_242);
and U959 (N_959,N_108,In_220);
nand U960 (N_960,In_1218,N_297);
and U961 (N_961,N_80,N_499);
and U962 (N_962,In_987,N_255);
nor U963 (N_963,In_1392,In_1487);
nand U964 (N_964,In_589,N_486);
nor U965 (N_965,N_267,N_14);
or U966 (N_966,In_121,In_209);
nor U967 (N_967,In_124,N_36);
or U968 (N_968,N_273,N_305);
nand U969 (N_969,In_621,N_85);
and U970 (N_970,N_334,In_369);
or U971 (N_971,N_373,In_319);
or U972 (N_972,In_1447,In_1150);
nor U973 (N_973,In_819,In_576);
and U974 (N_974,N_440,In_617);
nor U975 (N_975,In_1442,In_279);
nor U976 (N_976,In_696,In_1141);
or U977 (N_977,In_468,In_922);
nor U978 (N_978,N_465,N_381);
nand U979 (N_979,In_1470,In_323);
and U980 (N_980,N_134,In_205);
nand U981 (N_981,In_470,N_401);
and U982 (N_982,N_490,In_562);
xor U983 (N_983,N_138,In_1089);
and U984 (N_984,N_164,In_1100);
nand U985 (N_985,N_143,N_37);
nor U986 (N_986,N_447,In_611);
or U987 (N_987,N_478,N_24);
or U988 (N_988,In_325,N_8);
nand U989 (N_989,N_167,In_30);
nor U990 (N_990,In_426,In_29);
or U991 (N_991,N_159,N_479);
and U992 (N_992,In_570,In_531);
and U993 (N_993,In_952,N_482);
nor U994 (N_994,In_1028,In_401);
nor U995 (N_995,N_468,N_156);
xor U996 (N_996,In_552,In_1279);
and U997 (N_997,In_513,N_189);
xor U998 (N_998,N_492,In_172);
nor U999 (N_999,In_565,N_59);
xor U1000 (N_1000,N_638,N_545);
and U1001 (N_1001,N_729,N_682);
and U1002 (N_1002,N_990,N_580);
or U1003 (N_1003,N_736,N_964);
and U1004 (N_1004,N_853,N_702);
nor U1005 (N_1005,N_868,N_516);
or U1006 (N_1006,N_769,N_630);
or U1007 (N_1007,N_741,N_835);
or U1008 (N_1008,N_517,N_629);
or U1009 (N_1009,N_695,N_713);
and U1010 (N_1010,N_855,N_807);
nand U1011 (N_1011,N_792,N_989);
nand U1012 (N_1012,N_616,N_982);
or U1013 (N_1013,N_543,N_970);
and U1014 (N_1014,N_582,N_579);
or U1015 (N_1015,N_932,N_960);
nand U1016 (N_1016,N_951,N_896);
xor U1017 (N_1017,N_997,N_717);
xnor U1018 (N_1018,N_594,N_965);
or U1019 (N_1019,N_824,N_968);
or U1020 (N_1020,N_919,N_798);
and U1021 (N_1021,N_830,N_722);
nor U1022 (N_1022,N_565,N_825);
xor U1023 (N_1023,N_753,N_512);
nor U1024 (N_1024,N_891,N_870);
or U1025 (N_1025,N_791,N_762);
nor U1026 (N_1026,N_694,N_971);
xnor U1027 (N_1027,N_884,N_881);
or U1028 (N_1028,N_833,N_981);
or U1029 (N_1029,N_535,N_999);
and U1030 (N_1030,N_504,N_759);
and U1031 (N_1031,N_773,N_693);
and U1032 (N_1032,N_784,N_572);
xor U1033 (N_1033,N_635,N_644);
xor U1034 (N_1034,N_715,N_622);
or U1035 (N_1035,N_618,N_612);
xor U1036 (N_1036,N_969,N_872);
or U1037 (N_1037,N_901,N_885);
nor U1038 (N_1038,N_856,N_812);
nand U1039 (N_1039,N_666,N_567);
and U1040 (N_1040,N_863,N_734);
and U1041 (N_1041,N_506,N_542);
xor U1042 (N_1042,N_811,N_879);
or U1043 (N_1043,N_847,N_794);
nor U1044 (N_1044,N_749,N_514);
nand U1045 (N_1045,N_831,N_529);
nor U1046 (N_1046,N_846,N_684);
and U1047 (N_1047,N_934,N_966);
and U1048 (N_1048,N_710,N_692);
nor U1049 (N_1049,N_946,N_866);
nor U1050 (N_1050,N_748,N_574);
and U1051 (N_1051,N_728,N_568);
xor U1052 (N_1052,N_661,N_549);
nor U1053 (N_1053,N_887,N_813);
nor U1054 (N_1054,N_850,N_700);
or U1055 (N_1055,N_918,N_699);
and U1056 (N_1056,N_920,N_701);
nor U1057 (N_1057,N_680,N_716);
or U1058 (N_1058,N_554,N_986);
xor U1059 (N_1059,N_652,N_520);
nand U1060 (N_1060,N_895,N_928);
and U1061 (N_1061,N_834,N_528);
nand U1062 (N_1062,N_510,N_826);
nand U1063 (N_1063,N_585,N_735);
and U1064 (N_1064,N_795,N_774);
nor U1065 (N_1065,N_977,N_770);
nor U1066 (N_1066,N_783,N_503);
nor U1067 (N_1067,N_952,N_800);
nor U1068 (N_1068,N_511,N_653);
nand U1069 (N_1069,N_765,N_975);
or U1070 (N_1070,N_533,N_696);
xor U1071 (N_1071,N_739,N_842);
nor U1072 (N_1072,N_558,N_609);
nor U1073 (N_1073,N_610,N_808);
xor U1074 (N_1074,N_818,N_714);
nor U1075 (N_1075,N_524,N_843);
nand U1076 (N_1076,N_522,N_737);
nand U1077 (N_1077,N_780,N_740);
or U1078 (N_1078,N_756,N_598);
nand U1079 (N_1079,N_844,N_996);
xor U1080 (N_1080,N_561,N_976);
or U1081 (N_1081,N_892,N_793);
or U1082 (N_1082,N_651,N_669);
nor U1083 (N_1083,N_987,N_851);
xor U1084 (N_1084,N_963,N_782);
xnor U1085 (N_1085,N_867,N_913);
and U1086 (N_1086,N_679,N_910);
nand U1087 (N_1087,N_502,N_576);
nand U1088 (N_1088,N_967,N_665);
nor U1089 (N_1089,N_615,N_778);
nor U1090 (N_1090,N_926,N_933);
or U1091 (N_1091,N_556,N_859);
nor U1092 (N_1092,N_925,N_861);
or U1093 (N_1093,N_608,N_704);
or U1094 (N_1094,N_633,N_553);
nor U1095 (N_1095,N_840,N_927);
and U1096 (N_1096,N_530,N_632);
nand U1097 (N_1097,N_537,N_779);
or U1098 (N_1098,N_688,N_540);
xnor U1099 (N_1099,N_691,N_600);
or U1100 (N_1100,N_660,N_555);
nand U1101 (N_1101,N_930,N_950);
or U1102 (N_1102,N_854,N_974);
nand U1103 (N_1103,N_822,N_874);
nor U1104 (N_1104,N_973,N_804);
nand U1105 (N_1105,N_828,N_601);
and U1106 (N_1106,N_698,N_689);
and U1107 (N_1107,N_532,N_864);
nor U1108 (N_1108,N_501,N_742);
and U1109 (N_1109,N_876,N_978);
nor U1110 (N_1110,N_738,N_519);
and U1111 (N_1111,N_873,N_938);
and U1112 (N_1112,N_706,N_655);
nand U1113 (N_1113,N_577,N_726);
nor U1114 (N_1114,N_531,N_709);
nand U1115 (N_1115,N_668,N_639);
nand U1116 (N_1116,N_823,N_958);
and U1117 (N_1117,N_733,N_602);
and U1118 (N_1118,N_562,N_569);
nand U1119 (N_1119,N_755,N_827);
nor U1120 (N_1120,N_637,N_687);
nor U1121 (N_1121,N_607,N_546);
xnor U1122 (N_1122,N_536,N_659);
or U1123 (N_1123,N_515,N_583);
nand U1124 (N_1124,N_908,N_788);
or U1125 (N_1125,N_882,N_747);
nor U1126 (N_1126,N_586,N_525);
xor U1127 (N_1127,N_905,N_673);
nor U1128 (N_1128,N_810,N_648);
and U1129 (N_1129,N_513,N_760);
or U1130 (N_1130,N_604,N_595);
or U1131 (N_1131,N_566,N_838);
nand U1132 (N_1132,N_758,N_957);
nand U1133 (N_1133,N_898,N_647);
nand U1134 (N_1134,N_781,N_708);
or U1135 (N_1135,N_605,N_730);
nor U1136 (N_1136,N_954,N_785);
and U1137 (N_1137,N_814,N_761);
xor U1138 (N_1138,N_750,N_658);
nor U1139 (N_1139,N_771,N_902);
or U1140 (N_1140,N_796,N_538);
nand U1141 (N_1141,N_937,N_571);
nor U1142 (N_1142,N_912,N_945);
xnor U1143 (N_1143,N_640,N_563);
and U1144 (N_1144,N_596,N_707);
and U1145 (N_1145,N_862,N_900);
nor U1146 (N_1146,N_766,N_819);
xnor U1147 (N_1147,N_581,N_929);
or U1148 (N_1148,N_797,N_685);
nand U1149 (N_1149,N_805,N_712);
nand U1150 (N_1150,N_994,N_664);
xnor U1151 (N_1151,N_552,N_832);
nand U1152 (N_1152,N_956,N_718);
xor U1153 (N_1153,N_817,N_625);
nand U1154 (N_1154,N_526,N_559);
nand U1155 (N_1155,N_676,N_993);
nor U1156 (N_1156,N_939,N_723);
and U1157 (N_1157,N_907,N_806);
nor U1158 (N_1158,N_578,N_899);
or U1159 (N_1159,N_654,N_829);
and U1160 (N_1160,N_816,N_962);
nor U1161 (N_1161,N_650,N_720);
and U1162 (N_1162,N_935,N_683);
xor U1163 (N_1163,N_943,N_801);
nor U1164 (N_1164,N_507,N_906);
nor U1165 (N_1165,N_949,N_877);
and U1166 (N_1166,N_948,N_705);
or U1167 (N_1167,N_849,N_777);
nor U1168 (N_1168,N_883,N_621);
or U1169 (N_1169,N_955,N_623);
and U1170 (N_1170,N_626,N_799);
nor U1171 (N_1171,N_772,N_551);
and U1172 (N_1172,N_988,N_611);
and U1173 (N_1173,N_697,N_643);
or U1174 (N_1174,N_865,N_848);
xor U1175 (N_1175,N_603,N_686);
and U1176 (N_1176,N_983,N_992);
and U1177 (N_1177,N_936,N_869);
and U1178 (N_1178,N_509,N_893);
nand U1179 (N_1179,N_672,N_878);
or U1180 (N_1180,N_790,N_678);
or U1181 (N_1181,N_575,N_809);
or U1182 (N_1182,N_570,N_593);
nand U1183 (N_1183,N_991,N_727);
nor U1184 (N_1184,N_539,N_518);
and U1185 (N_1185,N_914,N_550);
or U1186 (N_1186,N_573,N_663);
and U1187 (N_1187,N_627,N_961);
xor U1188 (N_1188,N_886,N_703);
nor U1189 (N_1189,N_624,N_557);
nor U1190 (N_1190,N_613,N_751);
nor U1191 (N_1191,N_721,N_942);
nand U1192 (N_1192,N_821,N_634);
xor U1193 (N_1193,N_614,N_764);
xor U1194 (N_1194,N_754,N_860);
and U1195 (N_1195,N_897,N_921);
and U1196 (N_1196,N_786,N_591);
and U1197 (N_1197,N_670,N_953);
nand U1198 (N_1198,N_675,N_662);
xor U1199 (N_1199,N_922,N_959);
nand U1200 (N_1200,N_521,N_836);
and U1201 (N_1201,N_592,N_674);
nand U1202 (N_1202,N_589,N_903);
and U1203 (N_1203,N_857,N_984);
nor U1204 (N_1204,N_636,N_619);
or U1205 (N_1205,N_995,N_845);
nand U1206 (N_1206,N_657,N_776);
or U1207 (N_1207,N_890,N_888);
and U1208 (N_1208,N_858,N_852);
and U1209 (N_1209,N_587,N_931);
nor U1210 (N_1210,N_719,N_839);
nor U1211 (N_1211,N_642,N_646);
nor U1212 (N_1212,N_671,N_924);
xnor U1213 (N_1213,N_880,N_606);
or U1214 (N_1214,N_775,N_641);
nand U1215 (N_1215,N_767,N_911);
or U1216 (N_1216,N_746,N_590);
and U1217 (N_1217,N_972,N_544);
nor U1218 (N_1218,N_894,N_889);
xnor U1219 (N_1219,N_711,N_789);
or U1220 (N_1220,N_527,N_505);
or U1221 (N_1221,N_547,N_820);
nor U1222 (N_1222,N_617,N_763);
nand U1223 (N_1223,N_560,N_677);
and U1224 (N_1224,N_998,N_523);
nor U1225 (N_1225,N_985,N_916);
nand U1226 (N_1226,N_667,N_744);
nand U1227 (N_1227,N_944,N_875);
nand U1228 (N_1228,N_815,N_752);
nor U1229 (N_1229,N_909,N_841);
xnor U1230 (N_1230,N_500,N_731);
or U1231 (N_1231,N_725,N_588);
nor U1232 (N_1232,N_917,N_548);
and U1233 (N_1233,N_979,N_940);
nand U1234 (N_1234,N_947,N_802);
or U1235 (N_1235,N_923,N_904);
xnor U1236 (N_1236,N_980,N_620);
and U1237 (N_1237,N_599,N_941);
nand U1238 (N_1238,N_745,N_564);
or U1239 (N_1239,N_915,N_787);
nor U1240 (N_1240,N_628,N_534);
and U1241 (N_1241,N_597,N_690);
or U1242 (N_1242,N_757,N_508);
or U1243 (N_1243,N_743,N_681);
and U1244 (N_1244,N_656,N_871);
xnor U1245 (N_1245,N_732,N_649);
or U1246 (N_1246,N_645,N_837);
or U1247 (N_1247,N_803,N_768);
nand U1248 (N_1248,N_631,N_584);
nand U1249 (N_1249,N_541,N_724);
and U1250 (N_1250,N_579,N_981);
nor U1251 (N_1251,N_855,N_621);
xor U1252 (N_1252,N_535,N_801);
xor U1253 (N_1253,N_939,N_731);
or U1254 (N_1254,N_826,N_608);
nand U1255 (N_1255,N_539,N_619);
or U1256 (N_1256,N_698,N_832);
or U1257 (N_1257,N_895,N_986);
and U1258 (N_1258,N_700,N_885);
nor U1259 (N_1259,N_783,N_784);
nand U1260 (N_1260,N_974,N_896);
or U1261 (N_1261,N_569,N_752);
and U1262 (N_1262,N_819,N_561);
nand U1263 (N_1263,N_666,N_947);
or U1264 (N_1264,N_876,N_633);
or U1265 (N_1265,N_993,N_771);
or U1266 (N_1266,N_913,N_921);
nand U1267 (N_1267,N_523,N_536);
nor U1268 (N_1268,N_507,N_934);
and U1269 (N_1269,N_607,N_702);
nand U1270 (N_1270,N_526,N_797);
or U1271 (N_1271,N_558,N_821);
or U1272 (N_1272,N_538,N_614);
nand U1273 (N_1273,N_582,N_923);
and U1274 (N_1274,N_922,N_592);
nor U1275 (N_1275,N_604,N_675);
nor U1276 (N_1276,N_753,N_823);
and U1277 (N_1277,N_675,N_986);
and U1278 (N_1278,N_993,N_519);
nand U1279 (N_1279,N_938,N_708);
nand U1280 (N_1280,N_701,N_821);
nand U1281 (N_1281,N_578,N_963);
xor U1282 (N_1282,N_952,N_662);
and U1283 (N_1283,N_981,N_544);
nand U1284 (N_1284,N_877,N_559);
xnor U1285 (N_1285,N_610,N_884);
or U1286 (N_1286,N_673,N_816);
or U1287 (N_1287,N_882,N_656);
and U1288 (N_1288,N_904,N_903);
xnor U1289 (N_1289,N_911,N_682);
or U1290 (N_1290,N_549,N_876);
or U1291 (N_1291,N_520,N_911);
and U1292 (N_1292,N_751,N_810);
or U1293 (N_1293,N_882,N_596);
nor U1294 (N_1294,N_823,N_764);
or U1295 (N_1295,N_901,N_569);
nand U1296 (N_1296,N_797,N_961);
or U1297 (N_1297,N_745,N_922);
xnor U1298 (N_1298,N_520,N_951);
and U1299 (N_1299,N_500,N_590);
and U1300 (N_1300,N_575,N_840);
or U1301 (N_1301,N_508,N_676);
and U1302 (N_1302,N_621,N_919);
and U1303 (N_1303,N_964,N_567);
nand U1304 (N_1304,N_604,N_872);
or U1305 (N_1305,N_670,N_509);
xnor U1306 (N_1306,N_712,N_568);
nand U1307 (N_1307,N_925,N_619);
and U1308 (N_1308,N_617,N_972);
nand U1309 (N_1309,N_826,N_928);
or U1310 (N_1310,N_903,N_550);
and U1311 (N_1311,N_658,N_564);
nand U1312 (N_1312,N_663,N_714);
or U1313 (N_1313,N_989,N_577);
nor U1314 (N_1314,N_715,N_996);
or U1315 (N_1315,N_866,N_805);
nor U1316 (N_1316,N_716,N_964);
nand U1317 (N_1317,N_785,N_673);
and U1318 (N_1318,N_845,N_747);
or U1319 (N_1319,N_577,N_719);
and U1320 (N_1320,N_867,N_799);
nand U1321 (N_1321,N_695,N_791);
and U1322 (N_1322,N_786,N_931);
nor U1323 (N_1323,N_654,N_608);
nand U1324 (N_1324,N_749,N_844);
and U1325 (N_1325,N_947,N_808);
nor U1326 (N_1326,N_831,N_740);
or U1327 (N_1327,N_885,N_946);
xor U1328 (N_1328,N_905,N_621);
or U1329 (N_1329,N_869,N_906);
or U1330 (N_1330,N_900,N_752);
nor U1331 (N_1331,N_860,N_874);
nand U1332 (N_1332,N_897,N_827);
nand U1333 (N_1333,N_966,N_672);
nor U1334 (N_1334,N_735,N_806);
nand U1335 (N_1335,N_822,N_935);
and U1336 (N_1336,N_536,N_508);
nand U1337 (N_1337,N_983,N_719);
and U1338 (N_1338,N_941,N_894);
or U1339 (N_1339,N_512,N_802);
nor U1340 (N_1340,N_598,N_787);
nand U1341 (N_1341,N_598,N_788);
and U1342 (N_1342,N_756,N_741);
and U1343 (N_1343,N_974,N_791);
and U1344 (N_1344,N_785,N_925);
or U1345 (N_1345,N_577,N_812);
nand U1346 (N_1346,N_792,N_882);
nand U1347 (N_1347,N_789,N_523);
and U1348 (N_1348,N_501,N_588);
and U1349 (N_1349,N_941,N_983);
nor U1350 (N_1350,N_993,N_968);
or U1351 (N_1351,N_556,N_997);
and U1352 (N_1352,N_873,N_687);
nand U1353 (N_1353,N_925,N_743);
or U1354 (N_1354,N_844,N_508);
and U1355 (N_1355,N_770,N_763);
nor U1356 (N_1356,N_832,N_912);
and U1357 (N_1357,N_609,N_987);
or U1358 (N_1358,N_995,N_938);
nand U1359 (N_1359,N_817,N_672);
or U1360 (N_1360,N_501,N_733);
or U1361 (N_1361,N_546,N_705);
nor U1362 (N_1362,N_749,N_842);
nor U1363 (N_1363,N_927,N_714);
nor U1364 (N_1364,N_560,N_945);
and U1365 (N_1365,N_748,N_779);
or U1366 (N_1366,N_951,N_550);
and U1367 (N_1367,N_853,N_546);
or U1368 (N_1368,N_981,N_691);
nor U1369 (N_1369,N_954,N_850);
or U1370 (N_1370,N_773,N_701);
nor U1371 (N_1371,N_998,N_606);
and U1372 (N_1372,N_676,N_573);
or U1373 (N_1373,N_809,N_815);
and U1374 (N_1374,N_945,N_572);
nand U1375 (N_1375,N_691,N_910);
nor U1376 (N_1376,N_699,N_786);
or U1377 (N_1377,N_611,N_980);
nand U1378 (N_1378,N_669,N_779);
nor U1379 (N_1379,N_732,N_841);
nand U1380 (N_1380,N_598,N_941);
nor U1381 (N_1381,N_626,N_504);
nand U1382 (N_1382,N_627,N_508);
and U1383 (N_1383,N_837,N_948);
and U1384 (N_1384,N_820,N_744);
nor U1385 (N_1385,N_806,N_749);
nor U1386 (N_1386,N_553,N_790);
or U1387 (N_1387,N_965,N_933);
nand U1388 (N_1388,N_984,N_572);
and U1389 (N_1389,N_666,N_713);
nor U1390 (N_1390,N_975,N_605);
nand U1391 (N_1391,N_523,N_989);
and U1392 (N_1392,N_996,N_974);
or U1393 (N_1393,N_505,N_661);
and U1394 (N_1394,N_921,N_605);
and U1395 (N_1395,N_505,N_993);
nor U1396 (N_1396,N_942,N_786);
xor U1397 (N_1397,N_808,N_886);
nor U1398 (N_1398,N_985,N_674);
and U1399 (N_1399,N_929,N_689);
or U1400 (N_1400,N_686,N_994);
nor U1401 (N_1401,N_814,N_893);
nor U1402 (N_1402,N_646,N_985);
or U1403 (N_1403,N_804,N_925);
nor U1404 (N_1404,N_931,N_657);
nor U1405 (N_1405,N_514,N_664);
nand U1406 (N_1406,N_534,N_710);
nand U1407 (N_1407,N_508,N_690);
nor U1408 (N_1408,N_586,N_507);
nor U1409 (N_1409,N_896,N_569);
or U1410 (N_1410,N_807,N_645);
and U1411 (N_1411,N_629,N_573);
or U1412 (N_1412,N_563,N_871);
nand U1413 (N_1413,N_895,N_513);
nand U1414 (N_1414,N_528,N_593);
nor U1415 (N_1415,N_808,N_965);
nor U1416 (N_1416,N_799,N_598);
and U1417 (N_1417,N_699,N_681);
nor U1418 (N_1418,N_984,N_528);
or U1419 (N_1419,N_729,N_517);
nand U1420 (N_1420,N_844,N_976);
or U1421 (N_1421,N_772,N_767);
or U1422 (N_1422,N_638,N_744);
and U1423 (N_1423,N_540,N_774);
nor U1424 (N_1424,N_895,N_749);
nor U1425 (N_1425,N_712,N_638);
and U1426 (N_1426,N_784,N_525);
nor U1427 (N_1427,N_612,N_578);
or U1428 (N_1428,N_664,N_797);
nand U1429 (N_1429,N_519,N_942);
and U1430 (N_1430,N_812,N_876);
and U1431 (N_1431,N_693,N_910);
or U1432 (N_1432,N_815,N_502);
and U1433 (N_1433,N_638,N_826);
and U1434 (N_1434,N_932,N_733);
xor U1435 (N_1435,N_504,N_569);
nor U1436 (N_1436,N_983,N_751);
and U1437 (N_1437,N_571,N_810);
nand U1438 (N_1438,N_826,N_625);
or U1439 (N_1439,N_679,N_593);
and U1440 (N_1440,N_762,N_953);
or U1441 (N_1441,N_754,N_865);
and U1442 (N_1442,N_875,N_521);
and U1443 (N_1443,N_811,N_576);
or U1444 (N_1444,N_628,N_822);
or U1445 (N_1445,N_578,N_587);
nor U1446 (N_1446,N_550,N_818);
nand U1447 (N_1447,N_563,N_789);
nand U1448 (N_1448,N_767,N_574);
or U1449 (N_1449,N_650,N_940);
xor U1450 (N_1450,N_904,N_583);
and U1451 (N_1451,N_851,N_948);
or U1452 (N_1452,N_636,N_923);
nand U1453 (N_1453,N_797,N_780);
nor U1454 (N_1454,N_624,N_586);
nor U1455 (N_1455,N_915,N_742);
or U1456 (N_1456,N_809,N_879);
nor U1457 (N_1457,N_747,N_994);
xnor U1458 (N_1458,N_853,N_870);
xnor U1459 (N_1459,N_576,N_601);
nor U1460 (N_1460,N_930,N_702);
nor U1461 (N_1461,N_876,N_891);
or U1462 (N_1462,N_775,N_631);
and U1463 (N_1463,N_953,N_761);
or U1464 (N_1464,N_853,N_975);
nor U1465 (N_1465,N_680,N_766);
nand U1466 (N_1466,N_681,N_819);
nand U1467 (N_1467,N_695,N_661);
nand U1468 (N_1468,N_890,N_721);
nor U1469 (N_1469,N_745,N_578);
nor U1470 (N_1470,N_820,N_644);
nor U1471 (N_1471,N_578,N_681);
nand U1472 (N_1472,N_905,N_854);
nand U1473 (N_1473,N_676,N_911);
nand U1474 (N_1474,N_993,N_963);
nand U1475 (N_1475,N_602,N_569);
nor U1476 (N_1476,N_809,N_764);
xor U1477 (N_1477,N_897,N_814);
nor U1478 (N_1478,N_886,N_977);
nand U1479 (N_1479,N_881,N_792);
and U1480 (N_1480,N_981,N_830);
or U1481 (N_1481,N_588,N_975);
nor U1482 (N_1482,N_797,N_775);
or U1483 (N_1483,N_710,N_920);
and U1484 (N_1484,N_959,N_807);
xnor U1485 (N_1485,N_706,N_996);
nand U1486 (N_1486,N_739,N_585);
nand U1487 (N_1487,N_978,N_913);
nor U1488 (N_1488,N_974,N_917);
and U1489 (N_1489,N_740,N_715);
nand U1490 (N_1490,N_909,N_643);
and U1491 (N_1491,N_964,N_706);
or U1492 (N_1492,N_976,N_842);
nor U1493 (N_1493,N_811,N_850);
or U1494 (N_1494,N_824,N_772);
or U1495 (N_1495,N_740,N_750);
or U1496 (N_1496,N_896,N_528);
and U1497 (N_1497,N_728,N_658);
nor U1498 (N_1498,N_824,N_885);
and U1499 (N_1499,N_558,N_594);
and U1500 (N_1500,N_1019,N_1077);
and U1501 (N_1501,N_1225,N_1091);
nand U1502 (N_1502,N_1229,N_1390);
nand U1503 (N_1503,N_1158,N_1072);
or U1504 (N_1504,N_1369,N_1307);
nand U1505 (N_1505,N_1032,N_1367);
nor U1506 (N_1506,N_1472,N_1220);
nor U1507 (N_1507,N_1011,N_1110);
nand U1508 (N_1508,N_1435,N_1421);
and U1509 (N_1509,N_1499,N_1012);
xnor U1510 (N_1510,N_1335,N_1079);
and U1511 (N_1511,N_1192,N_1135);
or U1512 (N_1512,N_1062,N_1164);
or U1513 (N_1513,N_1493,N_1191);
nand U1514 (N_1514,N_1174,N_1278);
nor U1515 (N_1515,N_1219,N_1046);
and U1516 (N_1516,N_1213,N_1450);
or U1517 (N_1517,N_1461,N_1061);
or U1518 (N_1518,N_1494,N_1363);
nand U1519 (N_1519,N_1113,N_1121);
xnor U1520 (N_1520,N_1156,N_1232);
nand U1521 (N_1521,N_1392,N_1495);
nand U1522 (N_1522,N_1427,N_1207);
or U1523 (N_1523,N_1333,N_1200);
nor U1524 (N_1524,N_1463,N_1237);
nor U1525 (N_1525,N_1180,N_1107);
or U1526 (N_1526,N_1394,N_1096);
or U1527 (N_1527,N_1184,N_1370);
and U1528 (N_1528,N_1210,N_1028);
nand U1529 (N_1529,N_1144,N_1029);
or U1530 (N_1530,N_1141,N_1197);
nor U1531 (N_1531,N_1134,N_1150);
or U1532 (N_1532,N_1424,N_1422);
nand U1533 (N_1533,N_1052,N_1477);
and U1534 (N_1534,N_1224,N_1290);
nor U1535 (N_1535,N_1188,N_1301);
nor U1536 (N_1536,N_1471,N_1397);
nor U1537 (N_1537,N_1273,N_1000);
and U1538 (N_1538,N_1337,N_1438);
nand U1539 (N_1539,N_1086,N_1124);
or U1540 (N_1540,N_1255,N_1389);
and U1541 (N_1541,N_1095,N_1442);
and U1542 (N_1542,N_1068,N_1020);
and U1543 (N_1543,N_1283,N_1221);
and U1544 (N_1544,N_1069,N_1203);
nand U1545 (N_1545,N_1492,N_1445);
or U1546 (N_1546,N_1168,N_1355);
nor U1547 (N_1547,N_1385,N_1145);
nor U1548 (N_1548,N_1300,N_1329);
and U1549 (N_1549,N_1374,N_1284);
nand U1550 (N_1550,N_1447,N_1256);
and U1551 (N_1551,N_1309,N_1230);
or U1552 (N_1552,N_1308,N_1119);
or U1553 (N_1553,N_1295,N_1194);
or U1554 (N_1554,N_1112,N_1280);
xor U1555 (N_1555,N_1212,N_1142);
nand U1556 (N_1556,N_1294,N_1281);
and U1557 (N_1557,N_1264,N_1274);
or U1558 (N_1558,N_1393,N_1449);
and U1559 (N_1559,N_1265,N_1382);
and U1560 (N_1560,N_1381,N_1328);
xnor U1561 (N_1561,N_1451,N_1259);
xor U1562 (N_1562,N_1462,N_1245);
nand U1563 (N_1563,N_1253,N_1338);
nor U1564 (N_1564,N_1303,N_1360);
xnor U1565 (N_1565,N_1478,N_1371);
and U1566 (N_1566,N_1423,N_1404);
and U1567 (N_1567,N_1227,N_1146);
or U1568 (N_1568,N_1205,N_1117);
or U1569 (N_1569,N_1130,N_1101);
nand U1570 (N_1570,N_1099,N_1088);
nor U1571 (N_1571,N_1400,N_1260);
and U1572 (N_1572,N_1023,N_1453);
or U1573 (N_1573,N_1272,N_1064);
nand U1574 (N_1574,N_1045,N_1487);
and U1575 (N_1575,N_1185,N_1004);
or U1576 (N_1576,N_1042,N_1143);
nor U1577 (N_1577,N_1330,N_1017);
and U1578 (N_1578,N_1286,N_1152);
xnor U1579 (N_1579,N_1054,N_1199);
nand U1580 (N_1580,N_1001,N_1246);
and U1581 (N_1581,N_1165,N_1342);
nand U1582 (N_1582,N_1109,N_1341);
nand U1583 (N_1583,N_1196,N_1456);
nor U1584 (N_1584,N_1208,N_1187);
nand U1585 (N_1585,N_1271,N_1037);
and U1586 (N_1586,N_1178,N_1258);
nand U1587 (N_1587,N_1345,N_1356);
or U1588 (N_1588,N_1351,N_1340);
xnor U1589 (N_1589,N_1008,N_1314);
and U1590 (N_1590,N_1395,N_1282);
nor U1591 (N_1591,N_1407,N_1151);
nand U1592 (N_1592,N_1074,N_1252);
nand U1593 (N_1593,N_1455,N_1129);
or U1594 (N_1594,N_1263,N_1240);
or U1595 (N_1595,N_1201,N_1365);
and U1596 (N_1596,N_1261,N_1093);
nand U1597 (N_1597,N_1209,N_1234);
nand U1598 (N_1598,N_1031,N_1076);
xnor U1599 (N_1599,N_1033,N_1327);
and U1600 (N_1600,N_1376,N_1247);
nor U1601 (N_1601,N_1161,N_1378);
or U1602 (N_1602,N_1318,N_1211);
and U1603 (N_1603,N_1235,N_1458);
and U1604 (N_1604,N_1304,N_1386);
and U1605 (N_1605,N_1412,N_1484);
nor U1606 (N_1606,N_1090,N_1018);
nand U1607 (N_1607,N_1025,N_1444);
xnor U1608 (N_1608,N_1324,N_1436);
or U1609 (N_1609,N_1137,N_1277);
or U1610 (N_1610,N_1287,N_1040);
or U1611 (N_1611,N_1114,N_1270);
nor U1612 (N_1612,N_1396,N_1359);
or U1613 (N_1613,N_1080,N_1266);
or U1614 (N_1614,N_1454,N_1116);
xnor U1615 (N_1615,N_1047,N_1497);
and U1616 (N_1616,N_1010,N_1343);
and U1617 (N_1617,N_1071,N_1094);
and U1618 (N_1618,N_1036,N_1167);
nor U1619 (N_1619,N_1122,N_1108);
xnor U1620 (N_1620,N_1014,N_1348);
and U1621 (N_1621,N_1157,N_1315);
xnor U1622 (N_1622,N_1479,N_1408);
or U1623 (N_1623,N_1440,N_1291);
and U1624 (N_1624,N_1457,N_1489);
and U1625 (N_1625,N_1417,N_1391);
nor U1626 (N_1626,N_1366,N_1419);
and U1627 (N_1627,N_1048,N_1005);
nand U1628 (N_1628,N_1089,N_1060);
or U1629 (N_1629,N_1331,N_1002);
or U1630 (N_1630,N_1193,N_1027);
or U1631 (N_1631,N_1081,N_1092);
xnor U1632 (N_1632,N_1206,N_1214);
or U1633 (N_1633,N_1349,N_1443);
nor U1634 (N_1634,N_1352,N_1414);
nor U1635 (N_1635,N_1358,N_1323);
nor U1636 (N_1636,N_1043,N_1083);
nand U1637 (N_1637,N_1222,N_1486);
and U1638 (N_1638,N_1420,N_1175);
and U1639 (N_1639,N_1465,N_1297);
or U1640 (N_1640,N_1415,N_1131);
nand U1641 (N_1641,N_1115,N_1148);
nand U1642 (N_1642,N_1321,N_1262);
and U1643 (N_1643,N_1267,N_1428);
nor U1644 (N_1644,N_1411,N_1357);
and U1645 (N_1645,N_1215,N_1183);
nor U1646 (N_1646,N_1310,N_1302);
xnor U1647 (N_1647,N_1228,N_1039);
nor U1648 (N_1648,N_1172,N_1276);
or U1649 (N_1649,N_1067,N_1053);
or U1650 (N_1650,N_1241,N_1179);
nand U1651 (N_1651,N_1133,N_1292);
nor U1652 (N_1652,N_1078,N_1459);
nor U1653 (N_1653,N_1306,N_1496);
nor U1654 (N_1654,N_1485,N_1413);
nand U1655 (N_1655,N_1147,N_1446);
nor U1656 (N_1656,N_1339,N_1476);
or U1657 (N_1657,N_1429,N_1473);
nand U1658 (N_1658,N_1403,N_1138);
nor U1659 (N_1659,N_1474,N_1176);
nor U1660 (N_1660,N_1275,N_1038);
or U1661 (N_1661,N_1195,N_1383);
and U1662 (N_1662,N_1250,N_1132);
nand U1663 (N_1663,N_1401,N_1475);
and U1664 (N_1664,N_1136,N_1063);
and U1665 (N_1665,N_1439,N_1239);
or U1666 (N_1666,N_1013,N_1312);
nor U1667 (N_1667,N_1057,N_1123);
xnor U1668 (N_1668,N_1384,N_1084);
nand U1669 (N_1669,N_1313,N_1464);
and U1670 (N_1670,N_1171,N_1059);
nand U1671 (N_1671,N_1326,N_1467);
or U1672 (N_1672,N_1433,N_1249);
nor U1673 (N_1673,N_1223,N_1051);
and U1674 (N_1674,N_1181,N_1035);
nand U1675 (N_1675,N_1202,N_1434);
nor U1676 (N_1676,N_1127,N_1009);
nand U1677 (N_1677,N_1418,N_1402);
or U1678 (N_1678,N_1106,N_1006);
xnor U1679 (N_1679,N_1490,N_1163);
and U1680 (N_1680,N_1041,N_1377);
xor U1681 (N_1681,N_1007,N_1254);
or U1682 (N_1682,N_1350,N_1320);
nor U1683 (N_1683,N_1398,N_1388);
nand U1684 (N_1684,N_1347,N_1379);
and U1685 (N_1685,N_1325,N_1003);
and U1686 (N_1686,N_1100,N_1026);
or U1687 (N_1687,N_1154,N_1097);
nor U1688 (N_1688,N_1128,N_1034);
or U1689 (N_1689,N_1288,N_1087);
nand U1690 (N_1690,N_1498,N_1044);
nor U1691 (N_1691,N_1336,N_1296);
nand U1692 (N_1692,N_1311,N_1480);
or U1693 (N_1693,N_1149,N_1437);
and U1694 (N_1694,N_1120,N_1217);
nor U1695 (N_1695,N_1066,N_1431);
nor U1696 (N_1696,N_1452,N_1021);
and U1697 (N_1697,N_1242,N_1022);
or U1698 (N_1698,N_1375,N_1073);
and U1699 (N_1699,N_1441,N_1160);
nand U1700 (N_1700,N_1102,N_1139);
and U1701 (N_1701,N_1125,N_1346);
and U1702 (N_1702,N_1056,N_1104);
nand U1703 (N_1703,N_1024,N_1016);
or U1704 (N_1704,N_1155,N_1353);
nand U1705 (N_1705,N_1070,N_1049);
and U1706 (N_1706,N_1460,N_1236);
and U1707 (N_1707,N_1238,N_1362);
or U1708 (N_1708,N_1305,N_1162);
nand U1709 (N_1709,N_1166,N_1298);
or U1710 (N_1710,N_1285,N_1416);
or U1711 (N_1711,N_1468,N_1082);
or U1712 (N_1712,N_1448,N_1491);
nor U1713 (N_1713,N_1153,N_1105);
xnor U1714 (N_1714,N_1322,N_1425);
xnor U1715 (N_1715,N_1204,N_1248);
xor U1716 (N_1716,N_1186,N_1354);
and U1717 (N_1717,N_1190,N_1111);
or U1718 (N_1718,N_1364,N_1103);
xnor U1719 (N_1719,N_1482,N_1483);
nor U1720 (N_1720,N_1399,N_1216);
nor U1721 (N_1721,N_1319,N_1030);
nor U1722 (N_1722,N_1481,N_1289);
or U1723 (N_1723,N_1269,N_1470);
and U1724 (N_1724,N_1177,N_1055);
nand U1725 (N_1725,N_1243,N_1182);
and U1726 (N_1726,N_1231,N_1466);
or U1727 (N_1727,N_1426,N_1244);
nor U1728 (N_1728,N_1334,N_1058);
or U1729 (N_1729,N_1218,N_1373);
and U1730 (N_1730,N_1198,N_1118);
and U1731 (N_1731,N_1380,N_1361);
or U1732 (N_1732,N_1406,N_1251);
or U1733 (N_1733,N_1344,N_1410);
xnor U1734 (N_1734,N_1317,N_1257);
or U1735 (N_1735,N_1098,N_1488);
or U1736 (N_1736,N_1065,N_1293);
nand U1737 (N_1737,N_1368,N_1169);
nor U1738 (N_1738,N_1430,N_1189);
nor U1739 (N_1739,N_1140,N_1372);
or U1740 (N_1740,N_1332,N_1226);
nand U1741 (N_1741,N_1015,N_1387);
nand U1742 (N_1742,N_1316,N_1469);
and U1743 (N_1743,N_1050,N_1432);
or U1744 (N_1744,N_1085,N_1233);
nand U1745 (N_1745,N_1268,N_1075);
or U1746 (N_1746,N_1279,N_1405);
nand U1747 (N_1747,N_1126,N_1159);
nor U1748 (N_1748,N_1409,N_1173);
nand U1749 (N_1749,N_1170,N_1299);
or U1750 (N_1750,N_1062,N_1131);
nand U1751 (N_1751,N_1073,N_1424);
or U1752 (N_1752,N_1483,N_1354);
nand U1753 (N_1753,N_1156,N_1170);
nand U1754 (N_1754,N_1357,N_1427);
nor U1755 (N_1755,N_1154,N_1100);
and U1756 (N_1756,N_1020,N_1054);
nor U1757 (N_1757,N_1342,N_1230);
or U1758 (N_1758,N_1377,N_1494);
and U1759 (N_1759,N_1455,N_1088);
nor U1760 (N_1760,N_1497,N_1089);
and U1761 (N_1761,N_1257,N_1172);
nor U1762 (N_1762,N_1475,N_1031);
or U1763 (N_1763,N_1415,N_1311);
and U1764 (N_1764,N_1241,N_1001);
and U1765 (N_1765,N_1140,N_1346);
or U1766 (N_1766,N_1341,N_1354);
nor U1767 (N_1767,N_1053,N_1007);
nand U1768 (N_1768,N_1276,N_1259);
or U1769 (N_1769,N_1318,N_1383);
or U1770 (N_1770,N_1166,N_1284);
and U1771 (N_1771,N_1459,N_1211);
or U1772 (N_1772,N_1222,N_1403);
and U1773 (N_1773,N_1119,N_1391);
and U1774 (N_1774,N_1489,N_1460);
or U1775 (N_1775,N_1292,N_1361);
or U1776 (N_1776,N_1304,N_1155);
nor U1777 (N_1777,N_1383,N_1042);
or U1778 (N_1778,N_1147,N_1461);
nand U1779 (N_1779,N_1371,N_1108);
nor U1780 (N_1780,N_1399,N_1087);
or U1781 (N_1781,N_1249,N_1458);
and U1782 (N_1782,N_1344,N_1114);
nand U1783 (N_1783,N_1314,N_1427);
or U1784 (N_1784,N_1278,N_1215);
nor U1785 (N_1785,N_1388,N_1357);
and U1786 (N_1786,N_1079,N_1314);
nand U1787 (N_1787,N_1240,N_1439);
nand U1788 (N_1788,N_1070,N_1143);
or U1789 (N_1789,N_1260,N_1072);
nand U1790 (N_1790,N_1329,N_1033);
nand U1791 (N_1791,N_1066,N_1127);
and U1792 (N_1792,N_1257,N_1274);
and U1793 (N_1793,N_1024,N_1051);
xnor U1794 (N_1794,N_1218,N_1083);
or U1795 (N_1795,N_1479,N_1451);
nor U1796 (N_1796,N_1369,N_1419);
nor U1797 (N_1797,N_1252,N_1066);
nand U1798 (N_1798,N_1351,N_1239);
xnor U1799 (N_1799,N_1391,N_1017);
or U1800 (N_1800,N_1048,N_1340);
and U1801 (N_1801,N_1147,N_1023);
or U1802 (N_1802,N_1276,N_1113);
or U1803 (N_1803,N_1445,N_1414);
and U1804 (N_1804,N_1291,N_1101);
and U1805 (N_1805,N_1139,N_1073);
and U1806 (N_1806,N_1400,N_1266);
nand U1807 (N_1807,N_1190,N_1438);
xnor U1808 (N_1808,N_1044,N_1355);
nor U1809 (N_1809,N_1397,N_1373);
nand U1810 (N_1810,N_1084,N_1250);
nor U1811 (N_1811,N_1044,N_1095);
nand U1812 (N_1812,N_1386,N_1147);
xnor U1813 (N_1813,N_1292,N_1166);
and U1814 (N_1814,N_1487,N_1267);
and U1815 (N_1815,N_1158,N_1059);
nand U1816 (N_1816,N_1433,N_1221);
or U1817 (N_1817,N_1465,N_1477);
or U1818 (N_1818,N_1486,N_1049);
and U1819 (N_1819,N_1466,N_1017);
and U1820 (N_1820,N_1065,N_1369);
xor U1821 (N_1821,N_1336,N_1470);
and U1822 (N_1822,N_1493,N_1008);
nor U1823 (N_1823,N_1193,N_1052);
nor U1824 (N_1824,N_1422,N_1249);
and U1825 (N_1825,N_1493,N_1063);
nand U1826 (N_1826,N_1265,N_1429);
xnor U1827 (N_1827,N_1438,N_1495);
and U1828 (N_1828,N_1458,N_1015);
xnor U1829 (N_1829,N_1290,N_1377);
nor U1830 (N_1830,N_1099,N_1174);
nor U1831 (N_1831,N_1203,N_1235);
nor U1832 (N_1832,N_1130,N_1369);
nand U1833 (N_1833,N_1495,N_1116);
and U1834 (N_1834,N_1213,N_1227);
nand U1835 (N_1835,N_1028,N_1495);
and U1836 (N_1836,N_1436,N_1297);
or U1837 (N_1837,N_1301,N_1461);
or U1838 (N_1838,N_1155,N_1083);
and U1839 (N_1839,N_1251,N_1305);
or U1840 (N_1840,N_1431,N_1056);
nor U1841 (N_1841,N_1144,N_1373);
nor U1842 (N_1842,N_1300,N_1302);
nor U1843 (N_1843,N_1367,N_1374);
or U1844 (N_1844,N_1334,N_1069);
or U1845 (N_1845,N_1221,N_1368);
nand U1846 (N_1846,N_1121,N_1419);
and U1847 (N_1847,N_1492,N_1280);
or U1848 (N_1848,N_1042,N_1102);
nor U1849 (N_1849,N_1371,N_1305);
nand U1850 (N_1850,N_1181,N_1410);
and U1851 (N_1851,N_1422,N_1037);
xor U1852 (N_1852,N_1367,N_1113);
and U1853 (N_1853,N_1084,N_1368);
nand U1854 (N_1854,N_1399,N_1294);
nand U1855 (N_1855,N_1156,N_1468);
nand U1856 (N_1856,N_1055,N_1431);
nor U1857 (N_1857,N_1230,N_1281);
and U1858 (N_1858,N_1138,N_1291);
and U1859 (N_1859,N_1000,N_1123);
nand U1860 (N_1860,N_1490,N_1285);
or U1861 (N_1861,N_1390,N_1246);
or U1862 (N_1862,N_1301,N_1330);
nor U1863 (N_1863,N_1353,N_1235);
nor U1864 (N_1864,N_1113,N_1219);
xnor U1865 (N_1865,N_1258,N_1395);
or U1866 (N_1866,N_1431,N_1260);
and U1867 (N_1867,N_1262,N_1446);
nor U1868 (N_1868,N_1373,N_1340);
and U1869 (N_1869,N_1395,N_1307);
and U1870 (N_1870,N_1491,N_1328);
and U1871 (N_1871,N_1481,N_1288);
nor U1872 (N_1872,N_1052,N_1028);
xor U1873 (N_1873,N_1479,N_1427);
and U1874 (N_1874,N_1188,N_1051);
or U1875 (N_1875,N_1282,N_1090);
nor U1876 (N_1876,N_1411,N_1082);
or U1877 (N_1877,N_1487,N_1226);
nor U1878 (N_1878,N_1248,N_1286);
nor U1879 (N_1879,N_1363,N_1296);
nor U1880 (N_1880,N_1232,N_1394);
nand U1881 (N_1881,N_1469,N_1151);
or U1882 (N_1882,N_1413,N_1143);
xnor U1883 (N_1883,N_1189,N_1063);
or U1884 (N_1884,N_1490,N_1140);
xnor U1885 (N_1885,N_1110,N_1425);
nor U1886 (N_1886,N_1395,N_1198);
or U1887 (N_1887,N_1137,N_1402);
nand U1888 (N_1888,N_1264,N_1097);
nor U1889 (N_1889,N_1165,N_1402);
and U1890 (N_1890,N_1239,N_1402);
nor U1891 (N_1891,N_1022,N_1320);
and U1892 (N_1892,N_1378,N_1142);
and U1893 (N_1893,N_1418,N_1369);
and U1894 (N_1894,N_1434,N_1085);
xor U1895 (N_1895,N_1321,N_1048);
nor U1896 (N_1896,N_1097,N_1306);
and U1897 (N_1897,N_1068,N_1001);
and U1898 (N_1898,N_1263,N_1362);
and U1899 (N_1899,N_1056,N_1030);
or U1900 (N_1900,N_1366,N_1180);
or U1901 (N_1901,N_1340,N_1074);
nand U1902 (N_1902,N_1408,N_1216);
and U1903 (N_1903,N_1473,N_1302);
nand U1904 (N_1904,N_1482,N_1154);
nand U1905 (N_1905,N_1079,N_1356);
and U1906 (N_1906,N_1463,N_1133);
and U1907 (N_1907,N_1343,N_1232);
nor U1908 (N_1908,N_1358,N_1398);
xor U1909 (N_1909,N_1449,N_1098);
nor U1910 (N_1910,N_1065,N_1346);
or U1911 (N_1911,N_1433,N_1499);
or U1912 (N_1912,N_1355,N_1198);
or U1913 (N_1913,N_1214,N_1209);
nand U1914 (N_1914,N_1482,N_1399);
or U1915 (N_1915,N_1089,N_1331);
nor U1916 (N_1916,N_1359,N_1033);
xor U1917 (N_1917,N_1177,N_1007);
and U1918 (N_1918,N_1117,N_1168);
and U1919 (N_1919,N_1131,N_1221);
nand U1920 (N_1920,N_1423,N_1109);
nor U1921 (N_1921,N_1352,N_1377);
nor U1922 (N_1922,N_1270,N_1466);
nor U1923 (N_1923,N_1098,N_1211);
nand U1924 (N_1924,N_1208,N_1283);
xnor U1925 (N_1925,N_1184,N_1461);
nor U1926 (N_1926,N_1159,N_1133);
nor U1927 (N_1927,N_1119,N_1108);
or U1928 (N_1928,N_1201,N_1354);
nor U1929 (N_1929,N_1384,N_1479);
or U1930 (N_1930,N_1357,N_1202);
nor U1931 (N_1931,N_1081,N_1247);
nand U1932 (N_1932,N_1457,N_1088);
or U1933 (N_1933,N_1221,N_1450);
nand U1934 (N_1934,N_1271,N_1410);
nor U1935 (N_1935,N_1337,N_1374);
or U1936 (N_1936,N_1149,N_1483);
nand U1937 (N_1937,N_1210,N_1394);
xnor U1938 (N_1938,N_1455,N_1443);
or U1939 (N_1939,N_1442,N_1283);
xnor U1940 (N_1940,N_1235,N_1220);
and U1941 (N_1941,N_1250,N_1234);
xnor U1942 (N_1942,N_1172,N_1345);
or U1943 (N_1943,N_1478,N_1036);
or U1944 (N_1944,N_1303,N_1481);
nor U1945 (N_1945,N_1297,N_1190);
or U1946 (N_1946,N_1373,N_1189);
or U1947 (N_1947,N_1467,N_1166);
nand U1948 (N_1948,N_1241,N_1307);
and U1949 (N_1949,N_1068,N_1417);
nor U1950 (N_1950,N_1466,N_1210);
and U1951 (N_1951,N_1175,N_1310);
and U1952 (N_1952,N_1175,N_1022);
nor U1953 (N_1953,N_1002,N_1118);
or U1954 (N_1954,N_1479,N_1480);
or U1955 (N_1955,N_1374,N_1416);
nor U1956 (N_1956,N_1249,N_1322);
nor U1957 (N_1957,N_1457,N_1362);
and U1958 (N_1958,N_1044,N_1281);
xor U1959 (N_1959,N_1006,N_1369);
and U1960 (N_1960,N_1253,N_1111);
and U1961 (N_1961,N_1224,N_1367);
or U1962 (N_1962,N_1161,N_1011);
or U1963 (N_1963,N_1039,N_1369);
and U1964 (N_1964,N_1321,N_1375);
nor U1965 (N_1965,N_1477,N_1366);
nand U1966 (N_1966,N_1260,N_1459);
nor U1967 (N_1967,N_1217,N_1384);
nor U1968 (N_1968,N_1428,N_1355);
or U1969 (N_1969,N_1234,N_1088);
or U1970 (N_1970,N_1485,N_1387);
and U1971 (N_1971,N_1025,N_1323);
nand U1972 (N_1972,N_1330,N_1047);
nand U1973 (N_1973,N_1102,N_1306);
nor U1974 (N_1974,N_1488,N_1191);
nand U1975 (N_1975,N_1259,N_1201);
nor U1976 (N_1976,N_1391,N_1130);
xor U1977 (N_1977,N_1155,N_1147);
nand U1978 (N_1978,N_1040,N_1417);
nand U1979 (N_1979,N_1330,N_1238);
xor U1980 (N_1980,N_1464,N_1317);
xor U1981 (N_1981,N_1212,N_1107);
and U1982 (N_1982,N_1189,N_1048);
or U1983 (N_1983,N_1290,N_1073);
nor U1984 (N_1984,N_1350,N_1075);
nand U1985 (N_1985,N_1135,N_1064);
nor U1986 (N_1986,N_1415,N_1087);
or U1987 (N_1987,N_1104,N_1204);
and U1988 (N_1988,N_1481,N_1053);
or U1989 (N_1989,N_1354,N_1345);
xor U1990 (N_1990,N_1232,N_1141);
xnor U1991 (N_1991,N_1180,N_1047);
or U1992 (N_1992,N_1364,N_1382);
or U1993 (N_1993,N_1180,N_1241);
nor U1994 (N_1994,N_1363,N_1098);
nand U1995 (N_1995,N_1218,N_1286);
nand U1996 (N_1996,N_1263,N_1467);
and U1997 (N_1997,N_1260,N_1409);
nor U1998 (N_1998,N_1387,N_1314);
nand U1999 (N_1999,N_1328,N_1126);
nor U2000 (N_2000,N_1905,N_1550);
nand U2001 (N_2001,N_1881,N_1712);
and U2002 (N_2002,N_1955,N_1853);
and U2003 (N_2003,N_1738,N_1925);
nand U2004 (N_2004,N_1721,N_1632);
and U2005 (N_2005,N_1743,N_1602);
or U2006 (N_2006,N_1787,N_1578);
nor U2007 (N_2007,N_1669,N_1848);
xor U2008 (N_2008,N_1623,N_1840);
and U2009 (N_2009,N_1614,N_1637);
nor U2010 (N_2010,N_1872,N_1768);
nand U2011 (N_2011,N_1877,N_1554);
and U2012 (N_2012,N_1819,N_1635);
or U2013 (N_2013,N_1907,N_1826);
nand U2014 (N_2014,N_1603,N_1668);
or U2015 (N_2015,N_1571,N_1938);
nor U2016 (N_2016,N_1735,N_1770);
nor U2017 (N_2017,N_1854,N_1715);
nand U2018 (N_2018,N_1551,N_1744);
nor U2019 (N_2019,N_1675,N_1720);
or U2020 (N_2020,N_1884,N_1564);
or U2021 (N_2021,N_1645,N_1761);
nand U2022 (N_2022,N_1994,N_1508);
and U2023 (N_2023,N_1555,N_1656);
and U2024 (N_2024,N_1788,N_1689);
xor U2025 (N_2025,N_1500,N_1811);
or U2026 (N_2026,N_1902,N_1882);
or U2027 (N_2027,N_1654,N_1847);
or U2028 (N_2028,N_1983,N_1958);
nor U2029 (N_2029,N_1749,N_1501);
and U2030 (N_2030,N_1934,N_1783);
nand U2031 (N_2031,N_1676,N_1965);
nand U2032 (N_2032,N_1827,N_1923);
or U2033 (N_2033,N_1940,N_1653);
and U2034 (N_2034,N_1651,N_1672);
nor U2035 (N_2035,N_1541,N_1652);
or U2036 (N_2036,N_1893,N_1575);
or U2037 (N_2037,N_1560,N_1778);
nand U2038 (N_2038,N_1939,N_1937);
and U2039 (N_2039,N_1906,N_1506);
nand U2040 (N_2040,N_1512,N_1729);
nor U2041 (N_2041,N_1953,N_1998);
nor U2042 (N_2042,N_1982,N_1582);
nor U2043 (N_2043,N_1693,N_1756);
or U2044 (N_2044,N_1518,N_1918);
or U2045 (N_2045,N_1869,N_1849);
nand U2046 (N_2046,N_1973,N_1642);
and U2047 (N_2047,N_1775,N_1910);
and U2048 (N_2048,N_1886,N_1935);
nor U2049 (N_2049,N_1640,N_1921);
xor U2050 (N_2050,N_1839,N_1584);
nor U2051 (N_2051,N_1926,N_1966);
xnor U2052 (N_2052,N_1596,N_1810);
nor U2053 (N_2053,N_1972,N_1750);
nor U2054 (N_2054,N_1682,N_1838);
nand U2055 (N_2055,N_1821,N_1532);
xnor U2056 (N_2056,N_1539,N_1798);
or U2057 (N_2057,N_1647,N_1719);
nor U2058 (N_2058,N_1597,N_1694);
nand U2059 (N_2059,N_1969,N_1540);
nand U2060 (N_2060,N_1618,N_1981);
or U2061 (N_2061,N_1638,N_1894);
nand U2062 (N_2062,N_1552,N_1570);
xnor U2063 (N_2063,N_1948,N_1780);
or U2064 (N_2064,N_1785,N_1858);
xnor U2065 (N_2065,N_1663,N_1723);
and U2066 (N_2066,N_1643,N_1852);
and U2067 (N_2067,N_1868,N_1874);
nor U2068 (N_2068,N_1888,N_1836);
nor U2069 (N_2069,N_1559,N_1714);
and U2070 (N_2070,N_1547,N_1957);
or U2071 (N_2071,N_1863,N_1701);
xor U2072 (N_2072,N_1624,N_1943);
and U2073 (N_2073,N_1776,N_1542);
nor U2074 (N_2074,N_1724,N_1519);
and U2075 (N_2075,N_1753,N_1802);
nand U2076 (N_2076,N_1699,N_1931);
nor U2077 (N_2077,N_1598,N_1583);
xor U2078 (N_2078,N_1686,N_1862);
and U2079 (N_2079,N_1646,N_1534);
xnor U2080 (N_2080,N_1612,N_1851);
nand U2081 (N_2081,N_1708,N_1565);
and U2082 (N_2082,N_1580,N_1890);
nor U2083 (N_2083,N_1625,N_1870);
or U2084 (N_2084,N_1837,N_1691);
nand U2085 (N_2085,N_1610,N_1748);
xnor U2086 (N_2086,N_1704,N_1795);
and U2087 (N_2087,N_1977,N_1760);
nor U2088 (N_2088,N_1845,N_1641);
and U2089 (N_2089,N_1590,N_1628);
and U2090 (N_2090,N_1562,N_1967);
nor U2091 (N_2091,N_1791,N_1667);
nor U2092 (N_2092,N_1546,N_1855);
nand U2093 (N_2093,N_1589,N_1947);
or U2094 (N_2094,N_1573,N_1746);
and U2095 (N_2095,N_1620,N_1703);
nor U2096 (N_2096,N_1657,N_1754);
nand U2097 (N_2097,N_1767,N_1803);
nand U2098 (N_2098,N_1685,N_1569);
nor U2099 (N_2099,N_1912,N_1524);
or U2100 (N_2100,N_1961,N_1717);
nor U2101 (N_2101,N_1889,N_1666);
or U2102 (N_2102,N_1526,N_1670);
or U2103 (N_2103,N_1974,N_1528);
nor U2104 (N_2104,N_1509,N_1636);
xnor U2105 (N_2105,N_1777,N_1914);
nor U2106 (N_2106,N_1794,N_1960);
and U2107 (N_2107,N_1711,N_1850);
nor U2108 (N_2108,N_1956,N_1728);
and U2109 (N_2109,N_1639,N_1825);
nor U2110 (N_2110,N_1739,N_1997);
nand U2111 (N_2111,N_1502,N_1504);
xor U2112 (N_2112,N_1747,N_1660);
or U2113 (N_2113,N_1986,N_1913);
and U2114 (N_2114,N_1873,N_1740);
nor U2115 (N_2115,N_1678,N_1805);
nor U2116 (N_2116,N_1959,N_1616);
and U2117 (N_2117,N_1710,N_1979);
xnor U2118 (N_2118,N_1769,N_1915);
nor U2119 (N_2119,N_1741,N_1976);
nand U2120 (N_2120,N_1800,N_1844);
nand U2121 (N_2121,N_1820,N_1615);
and U2122 (N_2122,N_1520,N_1722);
nor U2123 (N_2123,N_1503,N_1942);
and U2124 (N_2124,N_1930,N_1698);
nand U2125 (N_2125,N_1878,N_1813);
xor U2126 (N_2126,N_1807,N_1527);
or U2127 (N_2127,N_1865,N_1680);
nand U2128 (N_2128,N_1557,N_1814);
and U2129 (N_2129,N_1924,N_1815);
nand U2130 (N_2130,N_1611,N_1988);
nor U2131 (N_2131,N_1592,N_1606);
nand U2132 (N_2132,N_1707,N_1970);
and U2133 (N_2133,N_1688,N_1841);
xor U2134 (N_2134,N_1548,N_1644);
nor U2135 (N_2135,N_1594,N_1538);
nand U2136 (N_2136,N_1861,N_1655);
xnor U2137 (N_2137,N_1898,N_1608);
and U2138 (N_2138,N_1619,N_1659);
nand U2139 (N_2139,N_1731,N_1876);
or U2140 (N_2140,N_1909,N_1556);
nor U2141 (N_2141,N_1954,N_1936);
or U2142 (N_2142,N_1545,N_1897);
xnor U2143 (N_2143,N_1816,N_1808);
and U2144 (N_2144,N_1543,N_1757);
nand U2145 (N_2145,N_1662,N_1842);
and U2146 (N_2146,N_1919,N_1763);
xnor U2147 (N_2147,N_1859,N_1971);
nor U2148 (N_2148,N_1607,N_1864);
nor U2149 (N_2149,N_1629,N_1829);
nand U2150 (N_2150,N_1745,N_1515);
nand U2151 (N_2151,N_1984,N_1823);
nor U2152 (N_2152,N_1797,N_1649);
and U2153 (N_2153,N_1774,N_1895);
nor U2154 (N_2154,N_1796,N_1516);
nand U2155 (N_2155,N_1593,N_1790);
and U2156 (N_2156,N_1922,N_1674);
nor U2157 (N_2157,N_1736,N_1764);
or U2158 (N_2158,N_1630,N_1834);
nor U2159 (N_2159,N_1762,N_1987);
nand U2160 (N_2160,N_1963,N_1950);
nand U2161 (N_2161,N_1705,N_1581);
nand U2162 (N_2162,N_1991,N_1650);
or U2163 (N_2163,N_1732,N_1968);
or U2164 (N_2164,N_1944,N_1951);
nand U2165 (N_2165,N_1574,N_1759);
nor U2166 (N_2166,N_1946,N_1900);
nor U2167 (N_2167,N_1985,N_1737);
and U2168 (N_2168,N_1692,N_1779);
nand U2169 (N_2169,N_1846,N_1832);
and U2170 (N_2170,N_1673,N_1941);
or U2171 (N_2171,N_1999,N_1681);
xnor U2172 (N_2172,N_1978,N_1585);
xnor U2173 (N_2173,N_1995,N_1697);
and U2174 (N_2174,N_1742,N_1773);
xnor U2175 (N_2175,N_1713,N_1792);
and U2176 (N_2176,N_1758,N_1505);
nor U2177 (N_2177,N_1822,N_1989);
nand U2178 (N_2178,N_1591,N_1733);
xnor U2179 (N_2179,N_1522,N_1525);
or U2180 (N_2180,N_1806,N_1595);
xor U2181 (N_2181,N_1734,N_1600);
or U2182 (N_2182,N_1782,N_1605);
or U2183 (N_2183,N_1700,N_1871);
nand U2184 (N_2184,N_1752,N_1784);
and U2185 (N_2185,N_1599,N_1875);
or U2186 (N_2186,N_1601,N_1609);
nor U2187 (N_2187,N_1626,N_1665);
and U2188 (N_2188,N_1771,N_1521);
and U2189 (N_2189,N_1828,N_1949);
and U2190 (N_2190,N_1671,N_1661);
or U2191 (N_2191,N_1843,N_1772);
nor U2192 (N_2192,N_1812,N_1725);
nand U2193 (N_2193,N_1726,N_1892);
nand U2194 (N_2194,N_1709,N_1730);
nor U2195 (N_2195,N_1511,N_1572);
or U2196 (N_2196,N_1765,N_1718);
and U2197 (N_2197,N_1517,N_1818);
and U2198 (N_2198,N_1627,N_1945);
or U2199 (N_2199,N_1833,N_1690);
nor U2200 (N_2200,N_1677,N_1980);
and U2201 (N_2201,N_1604,N_1523);
nand U2202 (N_2202,N_1679,N_1824);
nand U2203 (N_2203,N_1755,N_1916);
and U2204 (N_2204,N_1896,N_1904);
nand U2205 (N_2205,N_1695,N_1567);
xnor U2206 (N_2206,N_1860,N_1766);
nand U2207 (N_2207,N_1835,N_1579);
nor U2208 (N_2208,N_1529,N_1558);
nand U2209 (N_2209,N_1634,N_1561);
xor U2210 (N_2210,N_1993,N_1587);
nor U2211 (N_2211,N_1856,N_1533);
or U2212 (N_2212,N_1866,N_1544);
nor U2213 (N_2213,N_1648,N_1952);
xnor U2214 (N_2214,N_1867,N_1751);
nand U2215 (N_2215,N_1996,N_1887);
nor U2216 (N_2216,N_1901,N_1831);
nand U2217 (N_2217,N_1588,N_1549);
nand U2218 (N_2218,N_1927,N_1563);
and U2219 (N_2219,N_1990,N_1879);
or U2220 (N_2220,N_1929,N_1553);
nor U2221 (N_2221,N_1536,N_1799);
xnor U2222 (N_2222,N_1566,N_1804);
nand U2223 (N_2223,N_1793,N_1622);
nand U2224 (N_2224,N_1917,N_1911);
nor U2225 (N_2225,N_1535,N_1880);
nand U2226 (N_2226,N_1903,N_1928);
nand U2227 (N_2227,N_1891,N_1617);
xnor U2228 (N_2228,N_1706,N_1537);
or U2229 (N_2229,N_1883,N_1781);
or U2230 (N_2230,N_1687,N_1530);
nand U2231 (N_2231,N_1716,N_1908);
and U2232 (N_2232,N_1920,N_1830);
and U2233 (N_2233,N_1586,N_1696);
nor U2234 (N_2234,N_1513,N_1568);
nor U2235 (N_2235,N_1817,N_1789);
nor U2236 (N_2236,N_1885,N_1633);
nand U2237 (N_2237,N_1857,N_1664);
nand U2238 (N_2238,N_1683,N_1975);
and U2239 (N_2239,N_1658,N_1631);
and U2240 (N_2240,N_1576,N_1507);
or U2241 (N_2241,N_1727,N_1684);
nand U2242 (N_2242,N_1531,N_1510);
xnor U2243 (N_2243,N_1809,N_1621);
or U2244 (N_2244,N_1964,N_1613);
nor U2245 (N_2245,N_1702,N_1932);
or U2246 (N_2246,N_1577,N_1933);
nand U2247 (N_2247,N_1801,N_1962);
nand U2248 (N_2248,N_1514,N_1899);
nor U2249 (N_2249,N_1786,N_1992);
nor U2250 (N_2250,N_1845,N_1698);
nor U2251 (N_2251,N_1547,N_1895);
nor U2252 (N_2252,N_1546,N_1501);
nand U2253 (N_2253,N_1615,N_1800);
nand U2254 (N_2254,N_1516,N_1752);
and U2255 (N_2255,N_1831,N_1722);
nor U2256 (N_2256,N_1862,N_1620);
nor U2257 (N_2257,N_1723,N_1644);
and U2258 (N_2258,N_1930,N_1882);
and U2259 (N_2259,N_1624,N_1511);
or U2260 (N_2260,N_1674,N_1958);
nor U2261 (N_2261,N_1855,N_1964);
and U2262 (N_2262,N_1536,N_1872);
or U2263 (N_2263,N_1813,N_1948);
or U2264 (N_2264,N_1677,N_1781);
nor U2265 (N_2265,N_1811,N_1576);
nand U2266 (N_2266,N_1943,N_1942);
and U2267 (N_2267,N_1877,N_1511);
or U2268 (N_2268,N_1901,N_1501);
xnor U2269 (N_2269,N_1863,N_1970);
nor U2270 (N_2270,N_1505,N_1868);
xor U2271 (N_2271,N_1712,N_1967);
and U2272 (N_2272,N_1760,N_1596);
and U2273 (N_2273,N_1914,N_1996);
nand U2274 (N_2274,N_1873,N_1520);
nand U2275 (N_2275,N_1706,N_1599);
nor U2276 (N_2276,N_1989,N_1790);
nand U2277 (N_2277,N_1516,N_1675);
xor U2278 (N_2278,N_1968,N_1748);
and U2279 (N_2279,N_1669,N_1574);
and U2280 (N_2280,N_1671,N_1862);
or U2281 (N_2281,N_1615,N_1933);
and U2282 (N_2282,N_1669,N_1766);
and U2283 (N_2283,N_1729,N_1561);
nor U2284 (N_2284,N_1910,N_1741);
nor U2285 (N_2285,N_1550,N_1980);
or U2286 (N_2286,N_1614,N_1589);
and U2287 (N_2287,N_1865,N_1858);
xor U2288 (N_2288,N_1777,N_1589);
nand U2289 (N_2289,N_1879,N_1942);
nor U2290 (N_2290,N_1840,N_1538);
or U2291 (N_2291,N_1885,N_1514);
nand U2292 (N_2292,N_1955,N_1719);
and U2293 (N_2293,N_1594,N_1990);
nor U2294 (N_2294,N_1879,N_1596);
nor U2295 (N_2295,N_1993,N_1808);
nor U2296 (N_2296,N_1753,N_1930);
xor U2297 (N_2297,N_1833,N_1879);
nand U2298 (N_2298,N_1738,N_1657);
nor U2299 (N_2299,N_1578,N_1666);
and U2300 (N_2300,N_1678,N_1742);
and U2301 (N_2301,N_1604,N_1881);
and U2302 (N_2302,N_1644,N_1565);
nor U2303 (N_2303,N_1893,N_1737);
and U2304 (N_2304,N_1598,N_1712);
or U2305 (N_2305,N_1631,N_1601);
nor U2306 (N_2306,N_1779,N_1600);
or U2307 (N_2307,N_1805,N_1919);
and U2308 (N_2308,N_1739,N_1762);
xor U2309 (N_2309,N_1960,N_1674);
nor U2310 (N_2310,N_1792,N_1920);
nor U2311 (N_2311,N_1681,N_1763);
nor U2312 (N_2312,N_1984,N_1738);
and U2313 (N_2313,N_1508,N_1874);
and U2314 (N_2314,N_1600,N_1852);
nor U2315 (N_2315,N_1869,N_1987);
nand U2316 (N_2316,N_1583,N_1641);
and U2317 (N_2317,N_1534,N_1945);
nor U2318 (N_2318,N_1970,N_1621);
or U2319 (N_2319,N_1759,N_1851);
nor U2320 (N_2320,N_1528,N_1556);
or U2321 (N_2321,N_1797,N_1922);
nor U2322 (N_2322,N_1741,N_1723);
and U2323 (N_2323,N_1695,N_1531);
nor U2324 (N_2324,N_1822,N_1833);
or U2325 (N_2325,N_1774,N_1870);
nor U2326 (N_2326,N_1714,N_1838);
or U2327 (N_2327,N_1825,N_1615);
xor U2328 (N_2328,N_1638,N_1735);
xnor U2329 (N_2329,N_1728,N_1834);
and U2330 (N_2330,N_1948,N_1754);
nor U2331 (N_2331,N_1818,N_1727);
and U2332 (N_2332,N_1735,N_1567);
or U2333 (N_2333,N_1938,N_1801);
nand U2334 (N_2334,N_1577,N_1701);
nand U2335 (N_2335,N_1949,N_1565);
xnor U2336 (N_2336,N_1552,N_1930);
and U2337 (N_2337,N_1735,N_1566);
and U2338 (N_2338,N_1723,N_1829);
or U2339 (N_2339,N_1835,N_1692);
nand U2340 (N_2340,N_1623,N_1527);
and U2341 (N_2341,N_1622,N_1516);
nand U2342 (N_2342,N_1665,N_1984);
and U2343 (N_2343,N_1951,N_1565);
or U2344 (N_2344,N_1551,N_1993);
nand U2345 (N_2345,N_1999,N_1543);
or U2346 (N_2346,N_1732,N_1952);
xnor U2347 (N_2347,N_1906,N_1658);
nor U2348 (N_2348,N_1650,N_1866);
xor U2349 (N_2349,N_1586,N_1686);
nand U2350 (N_2350,N_1537,N_1897);
and U2351 (N_2351,N_1866,N_1586);
nor U2352 (N_2352,N_1846,N_1870);
nor U2353 (N_2353,N_1752,N_1961);
nor U2354 (N_2354,N_1859,N_1597);
nand U2355 (N_2355,N_1872,N_1614);
nor U2356 (N_2356,N_1611,N_1905);
nor U2357 (N_2357,N_1758,N_1988);
and U2358 (N_2358,N_1752,N_1967);
or U2359 (N_2359,N_1576,N_1705);
xor U2360 (N_2360,N_1794,N_1735);
and U2361 (N_2361,N_1554,N_1581);
or U2362 (N_2362,N_1990,N_1829);
or U2363 (N_2363,N_1527,N_1879);
or U2364 (N_2364,N_1944,N_1520);
or U2365 (N_2365,N_1536,N_1994);
or U2366 (N_2366,N_1503,N_1643);
nor U2367 (N_2367,N_1840,N_1665);
and U2368 (N_2368,N_1805,N_1637);
xnor U2369 (N_2369,N_1885,N_1521);
nor U2370 (N_2370,N_1830,N_1898);
or U2371 (N_2371,N_1649,N_1604);
or U2372 (N_2372,N_1965,N_1728);
xor U2373 (N_2373,N_1637,N_1532);
and U2374 (N_2374,N_1984,N_1573);
nor U2375 (N_2375,N_1600,N_1961);
and U2376 (N_2376,N_1706,N_1937);
xor U2377 (N_2377,N_1635,N_1782);
nor U2378 (N_2378,N_1871,N_1562);
nor U2379 (N_2379,N_1819,N_1671);
or U2380 (N_2380,N_1824,N_1837);
or U2381 (N_2381,N_1981,N_1800);
nor U2382 (N_2382,N_1515,N_1743);
xor U2383 (N_2383,N_1582,N_1707);
and U2384 (N_2384,N_1539,N_1643);
nand U2385 (N_2385,N_1929,N_1770);
and U2386 (N_2386,N_1769,N_1799);
nand U2387 (N_2387,N_1682,N_1515);
or U2388 (N_2388,N_1730,N_1529);
nor U2389 (N_2389,N_1592,N_1689);
nand U2390 (N_2390,N_1817,N_1961);
or U2391 (N_2391,N_1859,N_1573);
nor U2392 (N_2392,N_1557,N_1826);
nand U2393 (N_2393,N_1950,N_1543);
and U2394 (N_2394,N_1863,N_1756);
nor U2395 (N_2395,N_1571,N_1816);
xnor U2396 (N_2396,N_1753,N_1719);
nor U2397 (N_2397,N_1669,N_1534);
and U2398 (N_2398,N_1632,N_1560);
and U2399 (N_2399,N_1582,N_1566);
or U2400 (N_2400,N_1627,N_1992);
and U2401 (N_2401,N_1812,N_1622);
or U2402 (N_2402,N_1913,N_1836);
or U2403 (N_2403,N_1688,N_1894);
nand U2404 (N_2404,N_1736,N_1834);
or U2405 (N_2405,N_1583,N_1964);
nand U2406 (N_2406,N_1884,N_1737);
and U2407 (N_2407,N_1788,N_1971);
nor U2408 (N_2408,N_1625,N_1857);
and U2409 (N_2409,N_1868,N_1519);
nor U2410 (N_2410,N_1651,N_1762);
or U2411 (N_2411,N_1557,N_1654);
and U2412 (N_2412,N_1939,N_1523);
or U2413 (N_2413,N_1777,N_1750);
nor U2414 (N_2414,N_1692,N_1964);
and U2415 (N_2415,N_1789,N_1886);
and U2416 (N_2416,N_1723,N_1976);
nand U2417 (N_2417,N_1796,N_1651);
or U2418 (N_2418,N_1823,N_1700);
or U2419 (N_2419,N_1924,N_1526);
nand U2420 (N_2420,N_1562,N_1541);
nand U2421 (N_2421,N_1819,N_1661);
and U2422 (N_2422,N_1666,N_1811);
or U2423 (N_2423,N_1531,N_1846);
nor U2424 (N_2424,N_1665,N_1728);
and U2425 (N_2425,N_1642,N_1640);
xor U2426 (N_2426,N_1744,N_1980);
nand U2427 (N_2427,N_1644,N_1511);
nand U2428 (N_2428,N_1763,N_1576);
nand U2429 (N_2429,N_1719,N_1538);
nand U2430 (N_2430,N_1535,N_1706);
nand U2431 (N_2431,N_1844,N_1662);
nor U2432 (N_2432,N_1730,N_1933);
or U2433 (N_2433,N_1567,N_1628);
or U2434 (N_2434,N_1969,N_1558);
or U2435 (N_2435,N_1826,N_1503);
nor U2436 (N_2436,N_1704,N_1505);
nand U2437 (N_2437,N_1528,N_1770);
and U2438 (N_2438,N_1509,N_1976);
nand U2439 (N_2439,N_1854,N_1884);
nor U2440 (N_2440,N_1599,N_1632);
and U2441 (N_2441,N_1653,N_1854);
and U2442 (N_2442,N_1608,N_1707);
or U2443 (N_2443,N_1587,N_1743);
nand U2444 (N_2444,N_1550,N_1565);
nand U2445 (N_2445,N_1699,N_1666);
nor U2446 (N_2446,N_1624,N_1541);
or U2447 (N_2447,N_1517,N_1879);
or U2448 (N_2448,N_1731,N_1986);
nand U2449 (N_2449,N_1887,N_1649);
nand U2450 (N_2450,N_1813,N_1812);
nand U2451 (N_2451,N_1583,N_1704);
nand U2452 (N_2452,N_1866,N_1501);
nor U2453 (N_2453,N_1968,N_1509);
xnor U2454 (N_2454,N_1970,N_1942);
xnor U2455 (N_2455,N_1765,N_1630);
and U2456 (N_2456,N_1577,N_1690);
and U2457 (N_2457,N_1952,N_1688);
or U2458 (N_2458,N_1713,N_1692);
or U2459 (N_2459,N_1862,N_1865);
xnor U2460 (N_2460,N_1561,N_1833);
and U2461 (N_2461,N_1988,N_1901);
or U2462 (N_2462,N_1775,N_1696);
nand U2463 (N_2463,N_1831,N_1798);
and U2464 (N_2464,N_1769,N_1968);
or U2465 (N_2465,N_1758,N_1525);
and U2466 (N_2466,N_1812,N_1995);
and U2467 (N_2467,N_1797,N_1812);
and U2468 (N_2468,N_1967,N_1512);
or U2469 (N_2469,N_1980,N_1839);
xnor U2470 (N_2470,N_1723,N_1970);
xnor U2471 (N_2471,N_1728,N_1589);
nand U2472 (N_2472,N_1772,N_1961);
nor U2473 (N_2473,N_1686,N_1879);
nor U2474 (N_2474,N_1940,N_1970);
and U2475 (N_2475,N_1836,N_1628);
nor U2476 (N_2476,N_1851,N_1579);
and U2477 (N_2477,N_1511,N_1785);
nand U2478 (N_2478,N_1808,N_1889);
or U2479 (N_2479,N_1940,N_1508);
nand U2480 (N_2480,N_1677,N_1818);
nor U2481 (N_2481,N_1979,N_1931);
nand U2482 (N_2482,N_1866,N_1618);
or U2483 (N_2483,N_1936,N_1760);
or U2484 (N_2484,N_1971,N_1792);
or U2485 (N_2485,N_1892,N_1689);
nand U2486 (N_2486,N_1966,N_1560);
or U2487 (N_2487,N_1612,N_1530);
xor U2488 (N_2488,N_1692,N_1608);
xnor U2489 (N_2489,N_1651,N_1648);
or U2490 (N_2490,N_1599,N_1997);
and U2491 (N_2491,N_1713,N_1983);
or U2492 (N_2492,N_1947,N_1638);
nand U2493 (N_2493,N_1925,N_1667);
nand U2494 (N_2494,N_1569,N_1688);
nor U2495 (N_2495,N_1553,N_1630);
nor U2496 (N_2496,N_1664,N_1643);
and U2497 (N_2497,N_1838,N_1589);
xor U2498 (N_2498,N_1851,N_1737);
nor U2499 (N_2499,N_1731,N_1640);
or U2500 (N_2500,N_2166,N_2315);
or U2501 (N_2501,N_2255,N_2041);
and U2502 (N_2502,N_2269,N_2175);
nor U2503 (N_2503,N_2251,N_2256);
nor U2504 (N_2504,N_2063,N_2361);
nor U2505 (N_2505,N_2123,N_2425);
or U2506 (N_2506,N_2356,N_2272);
or U2507 (N_2507,N_2039,N_2016);
nor U2508 (N_2508,N_2142,N_2342);
nand U2509 (N_2509,N_2216,N_2132);
nor U2510 (N_2510,N_2057,N_2185);
nor U2511 (N_2511,N_2150,N_2127);
nand U2512 (N_2512,N_2431,N_2261);
and U2513 (N_2513,N_2253,N_2310);
nor U2514 (N_2514,N_2217,N_2452);
nor U2515 (N_2515,N_2260,N_2349);
nor U2516 (N_2516,N_2043,N_2080);
or U2517 (N_2517,N_2324,N_2090);
nor U2518 (N_2518,N_2116,N_2044);
or U2519 (N_2519,N_2104,N_2005);
nand U2520 (N_2520,N_2240,N_2199);
nor U2521 (N_2521,N_2456,N_2494);
and U2522 (N_2522,N_2226,N_2164);
or U2523 (N_2523,N_2141,N_2233);
or U2524 (N_2524,N_2493,N_2239);
nor U2525 (N_2525,N_2284,N_2131);
or U2526 (N_2526,N_2443,N_2085);
or U2527 (N_2527,N_2320,N_2314);
and U2528 (N_2528,N_2335,N_2479);
or U2529 (N_2529,N_2299,N_2464);
nor U2530 (N_2530,N_2024,N_2028);
and U2531 (N_2531,N_2487,N_2343);
nor U2532 (N_2532,N_2082,N_2145);
or U2533 (N_2533,N_2154,N_2405);
nor U2534 (N_2534,N_2196,N_2308);
and U2535 (N_2535,N_2197,N_2302);
or U2536 (N_2536,N_2355,N_2176);
or U2537 (N_2537,N_2473,N_2222);
xnor U2538 (N_2538,N_2103,N_2388);
and U2539 (N_2539,N_2397,N_2428);
and U2540 (N_2540,N_2004,N_2088);
or U2541 (N_2541,N_2219,N_2440);
nand U2542 (N_2542,N_2481,N_2377);
nor U2543 (N_2543,N_2421,N_2432);
and U2544 (N_2544,N_2488,N_2186);
or U2545 (N_2545,N_2097,N_2159);
or U2546 (N_2546,N_2084,N_2398);
or U2547 (N_2547,N_2466,N_2411);
or U2548 (N_2548,N_2322,N_2409);
and U2549 (N_2549,N_2068,N_2160);
nand U2550 (N_2550,N_2205,N_2200);
nor U2551 (N_2551,N_2304,N_2072);
nor U2552 (N_2552,N_2029,N_2204);
or U2553 (N_2553,N_2404,N_2376);
nor U2554 (N_2554,N_2179,N_2275);
nand U2555 (N_2555,N_2012,N_2455);
or U2556 (N_2556,N_2054,N_2457);
nor U2557 (N_2557,N_2348,N_2424);
xor U2558 (N_2558,N_2468,N_2340);
and U2559 (N_2559,N_2143,N_2282);
nor U2560 (N_2560,N_2156,N_2357);
nand U2561 (N_2561,N_2098,N_2292);
xnor U2562 (N_2562,N_2379,N_2265);
xnor U2563 (N_2563,N_2483,N_2394);
nor U2564 (N_2564,N_2120,N_2025);
nand U2565 (N_2565,N_2445,N_2076);
nand U2566 (N_2566,N_2060,N_2318);
xor U2567 (N_2567,N_2095,N_2300);
nand U2568 (N_2568,N_2223,N_2105);
or U2569 (N_2569,N_2247,N_2259);
xor U2570 (N_2570,N_2218,N_2415);
and U2571 (N_2571,N_2181,N_2050);
nor U2572 (N_2572,N_2056,N_2283);
nor U2573 (N_2573,N_2371,N_2130);
or U2574 (N_2574,N_2389,N_2306);
nor U2575 (N_2575,N_2451,N_2401);
or U2576 (N_2576,N_2289,N_2110);
and U2577 (N_2577,N_2002,N_2426);
and U2578 (N_2578,N_2350,N_2212);
nand U2579 (N_2579,N_2046,N_2430);
nand U2580 (N_2580,N_2066,N_2037);
nand U2581 (N_2581,N_2263,N_2301);
nor U2582 (N_2582,N_2383,N_2158);
and U2583 (N_2583,N_2395,N_2450);
or U2584 (N_2584,N_2258,N_2385);
or U2585 (N_2585,N_2317,N_2359);
xnor U2586 (N_2586,N_2184,N_2246);
nor U2587 (N_2587,N_2210,N_2111);
or U2588 (N_2588,N_2091,N_2250);
nand U2589 (N_2589,N_2243,N_2168);
and U2590 (N_2590,N_2003,N_2345);
nand U2591 (N_2591,N_2262,N_2047);
or U2592 (N_2592,N_2071,N_2173);
nor U2593 (N_2593,N_2436,N_2209);
nand U2594 (N_2594,N_2416,N_2417);
nand U2595 (N_2595,N_2391,N_2220);
xor U2596 (N_2596,N_2434,N_2126);
or U2597 (N_2597,N_2378,N_2448);
nand U2598 (N_2598,N_2121,N_2172);
nand U2599 (N_2599,N_2491,N_2033);
xor U2600 (N_2600,N_2155,N_2297);
and U2601 (N_2601,N_2285,N_2387);
or U2602 (N_2602,N_2366,N_2169);
nor U2603 (N_2603,N_2045,N_2178);
and U2604 (N_2604,N_2118,N_2406);
and U2605 (N_2605,N_2369,N_2267);
nor U2606 (N_2606,N_2399,N_2058);
and U2607 (N_2607,N_2419,N_2472);
nand U2608 (N_2608,N_2461,N_2462);
nand U2609 (N_2609,N_2276,N_2278);
xor U2610 (N_2610,N_2174,N_2469);
nand U2611 (N_2611,N_2372,N_2193);
and U2612 (N_2612,N_2053,N_2007);
nor U2613 (N_2613,N_2000,N_2038);
nor U2614 (N_2614,N_2274,N_2454);
and U2615 (N_2615,N_2484,N_2157);
and U2616 (N_2616,N_2013,N_2362);
nand U2617 (N_2617,N_2192,N_2089);
and U2618 (N_2618,N_2138,N_2224);
or U2619 (N_2619,N_2319,N_2167);
and U2620 (N_2620,N_2069,N_2100);
nor U2621 (N_2621,N_2380,N_2374);
and U2622 (N_2622,N_2485,N_2460);
and U2623 (N_2623,N_2190,N_2093);
xor U2624 (N_2624,N_2497,N_2444);
and U2625 (N_2625,N_2286,N_2107);
and U2626 (N_2626,N_2202,N_2009);
nand U2627 (N_2627,N_2271,N_2227);
nand U2628 (N_2628,N_2042,N_2295);
nand U2629 (N_2629,N_2248,N_2006);
nor U2630 (N_2630,N_2489,N_2235);
nor U2631 (N_2631,N_2073,N_2188);
xor U2632 (N_2632,N_2402,N_2498);
and U2633 (N_2633,N_2102,N_2153);
and U2634 (N_2634,N_2242,N_2144);
or U2635 (N_2635,N_2403,N_2017);
and U2636 (N_2636,N_2108,N_2331);
or U2637 (N_2637,N_2467,N_2139);
nor U2638 (N_2638,N_2215,N_2270);
nor U2639 (N_2639,N_2393,N_2115);
or U2640 (N_2640,N_2026,N_2273);
nand U2641 (N_2641,N_2277,N_2040);
or U2642 (N_2642,N_2070,N_2293);
nand U2643 (N_2643,N_2344,N_2207);
and U2644 (N_2644,N_2392,N_2321);
nor U2645 (N_2645,N_2151,N_2477);
xor U2646 (N_2646,N_2470,N_2427);
or U2647 (N_2647,N_2458,N_2208);
nand U2648 (N_2648,N_2162,N_2294);
or U2649 (N_2649,N_2206,N_2305);
and U2650 (N_2650,N_2117,N_2365);
and U2651 (N_2651,N_2177,N_2133);
xor U2652 (N_2652,N_2211,N_2447);
nand U2653 (N_2653,N_2480,N_2171);
nand U2654 (N_2654,N_2059,N_2113);
nand U2655 (N_2655,N_2136,N_2030);
nand U2656 (N_2656,N_2413,N_2079);
and U2657 (N_2657,N_2170,N_2364);
nand U2658 (N_2658,N_2373,N_2396);
or U2659 (N_2659,N_2400,N_2386);
or U2660 (N_2660,N_2360,N_2307);
or U2661 (N_2661,N_2441,N_2119);
nor U2662 (N_2662,N_2412,N_2092);
nor U2663 (N_2663,N_2384,N_2252);
nand U2664 (N_2664,N_2244,N_2309);
and U2665 (N_2665,N_2475,N_2064);
nor U2666 (N_2666,N_2109,N_2194);
nor U2667 (N_2667,N_2074,N_2165);
or U2668 (N_2668,N_2241,N_2325);
or U2669 (N_2669,N_2279,N_2125);
nand U2670 (N_2670,N_2327,N_2333);
or U2671 (N_2671,N_2124,N_2140);
nor U2672 (N_2672,N_2015,N_2203);
and U2673 (N_2673,N_2099,N_2254);
nand U2674 (N_2674,N_2198,N_2474);
nor U2675 (N_2675,N_2330,N_2414);
and U2676 (N_2676,N_2363,N_2326);
xor U2677 (N_2677,N_2316,N_2490);
nor U2678 (N_2678,N_2429,N_2303);
xor U2679 (N_2679,N_2281,N_2449);
and U2680 (N_2680,N_2049,N_2328);
and U2681 (N_2681,N_2021,N_2332);
nor U2682 (N_2682,N_2237,N_2129);
nand U2683 (N_2683,N_2087,N_2423);
and U2684 (N_2684,N_2266,N_2478);
and U2685 (N_2685,N_2228,N_2354);
xor U2686 (N_2686,N_2114,N_2433);
nor U2687 (N_2687,N_2018,N_2336);
nor U2688 (N_2688,N_2358,N_2230);
nand U2689 (N_2689,N_2214,N_2347);
or U2690 (N_2690,N_2191,N_2137);
nor U2691 (N_2691,N_2337,N_2086);
nor U2692 (N_2692,N_2065,N_2075);
nor U2693 (N_2693,N_2496,N_2180);
and U2694 (N_2694,N_2339,N_2368);
nand U2695 (N_2695,N_2051,N_2189);
nor U2696 (N_2696,N_2135,N_2161);
or U2697 (N_2697,N_2268,N_2035);
or U2698 (N_2698,N_2311,N_2329);
and U2699 (N_2699,N_2234,N_2375);
or U2700 (N_2700,N_2463,N_2408);
and U2701 (N_2701,N_2020,N_2410);
or U2702 (N_2702,N_2122,N_2492);
or U2703 (N_2703,N_2081,N_2287);
nand U2704 (N_2704,N_2486,N_2232);
and U2705 (N_2705,N_2249,N_2078);
nor U2706 (N_2706,N_2312,N_2439);
nand U2707 (N_2707,N_2482,N_2438);
nor U2708 (N_2708,N_2465,N_2148);
nand U2709 (N_2709,N_2163,N_2229);
and U2710 (N_2710,N_2225,N_2221);
and U2711 (N_2711,N_2257,N_2435);
or U2712 (N_2712,N_2442,N_2201);
and U2713 (N_2713,N_2067,N_2338);
or U2714 (N_2714,N_2367,N_2476);
nor U2715 (N_2715,N_2027,N_2146);
or U2716 (N_2716,N_2055,N_2048);
and U2717 (N_2717,N_2022,N_2418);
nor U2718 (N_2718,N_2471,N_2236);
xnor U2719 (N_2719,N_2149,N_2370);
nor U2720 (N_2720,N_2019,N_2014);
xnor U2721 (N_2721,N_2062,N_2446);
and U2722 (N_2722,N_2052,N_2382);
or U2723 (N_2723,N_2183,N_2390);
or U2724 (N_2724,N_2381,N_2323);
nand U2725 (N_2725,N_2499,N_2453);
nand U2726 (N_2726,N_2341,N_2264);
or U2727 (N_2727,N_2152,N_2437);
nor U2728 (N_2728,N_2112,N_2407);
nor U2729 (N_2729,N_2008,N_2238);
and U2730 (N_2730,N_2288,N_2032);
nand U2731 (N_2731,N_2134,N_2023);
or U2732 (N_2732,N_2459,N_2034);
and U2733 (N_2733,N_2353,N_2245);
or U2734 (N_2734,N_2106,N_2346);
and U2735 (N_2735,N_2298,N_2077);
or U2736 (N_2736,N_2495,N_2187);
nor U2737 (N_2737,N_2296,N_2213);
and U2738 (N_2738,N_2101,N_2420);
xor U2739 (N_2739,N_2128,N_2036);
nand U2740 (N_2740,N_2313,N_2011);
and U2741 (N_2741,N_2290,N_2422);
or U2742 (N_2742,N_2280,N_2351);
and U2743 (N_2743,N_2031,N_2147);
nand U2744 (N_2744,N_2231,N_2195);
or U2745 (N_2745,N_2061,N_2096);
or U2746 (N_2746,N_2291,N_2334);
or U2747 (N_2747,N_2352,N_2001);
nand U2748 (N_2748,N_2083,N_2182);
xor U2749 (N_2749,N_2094,N_2010);
nand U2750 (N_2750,N_2121,N_2436);
or U2751 (N_2751,N_2240,N_2252);
nor U2752 (N_2752,N_2287,N_2033);
nand U2753 (N_2753,N_2134,N_2271);
nand U2754 (N_2754,N_2319,N_2456);
and U2755 (N_2755,N_2039,N_2421);
or U2756 (N_2756,N_2063,N_2354);
or U2757 (N_2757,N_2247,N_2015);
nand U2758 (N_2758,N_2110,N_2345);
nor U2759 (N_2759,N_2176,N_2363);
or U2760 (N_2760,N_2039,N_2195);
nor U2761 (N_2761,N_2323,N_2102);
nor U2762 (N_2762,N_2052,N_2186);
and U2763 (N_2763,N_2082,N_2301);
or U2764 (N_2764,N_2127,N_2032);
or U2765 (N_2765,N_2250,N_2368);
nand U2766 (N_2766,N_2033,N_2452);
nor U2767 (N_2767,N_2410,N_2083);
and U2768 (N_2768,N_2375,N_2305);
and U2769 (N_2769,N_2397,N_2422);
and U2770 (N_2770,N_2271,N_2035);
nand U2771 (N_2771,N_2066,N_2306);
and U2772 (N_2772,N_2458,N_2129);
and U2773 (N_2773,N_2488,N_2459);
and U2774 (N_2774,N_2266,N_2193);
and U2775 (N_2775,N_2140,N_2367);
or U2776 (N_2776,N_2407,N_2234);
and U2777 (N_2777,N_2237,N_2478);
nor U2778 (N_2778,N_2251,N_2197);
or U2779 (N_2779,N_2272,N_2111);
nand U2780 (N_2780,N_2467,N_2499);
nand U2781 (N_2781,N_2423,N_2089);
or U2782 (N_2782,N_2260,N_2382);
or U2783 (N_2783,N_2066,N_2370);
or U2784 (N_2784,N_2378,N_2427);
and U2785 (N_2785,N_2113,N_2233);
or U2786 (N_2786,N_2150,N_2418);
nand U2787 (N_2787,N_2263,N_2016);
nand U2788 (N_2788,N_2168,N_2459);
or U2789 (N_2789,N_2012,N_2489);
or U2790 (N_2790,N_2356,N_2259);
nand U2791 (N_2791,N_2216,N_2218);
nor U2792 (N_2792,N_2292,N_2167);
and U2793 (N_2793,N_2363,N_2478);
nand U2794 (N_2794,N_2097,N_2260);
nand U2795 (N_2795,N_2236,N_2089);
nor U2796 (N_2796,N_2290,N_2079);
or U2797 (N_2797,N_2226,N_2210);
and U2798 (N_2798,N_2145,N_2454);
or U2799 (N_2799,N_2144,N_2367);
or U2800 (N_2800,N_2015,N_2052);
and U2801 (N_2801,N_2423,N_2083);
or U2802 (N_2802,N_2129,N_2121);
nand U2803 (N_2803,N_2167,N_2300);
nand U2804 (N_2804,N_2482,N_2032);
xor U2805 (N_2805,N_2366,N_2298);
nor U2806 (N_2806,N_2128,N_2315);
xnor U2807 (N_2807,N_2285,N_2489);
nor U2808 (N_2808,N_2356,N_2053);
or U2809 (N_2809,N_2092,N_2104);
nor U2810 (N_2810,N_2389,N_2335);
and U2811 (N_2811,N_2031,N_2354);
or U2812 (N_2812,N_2188,N_2039);
or U2813 (N_2813,N_2437,N_2430);
and U2814 (N_2814,N_2127,N_2082);
nand U2815 (N_2815,N_2038,N_2488);
nor U2816 (N_2816,N_2168,N_2364);
nand U2817 (N_2817,N_2306,N_2134);
or U2818 (N_2818,N_2163,N_2131);
and U2819 (N_2819,N_2430,N_2045);
or U2820 (N_2820,N_2040,N_2298);
or U2821 (N_2821,N_2121,N_2438);
and U2822 (N_2822,N_2474,N_2197);
and U2823 (N_2823,N_2213,N_2324);
or U2824 (N_2824,N_2254,N_2054);
xnor U2825 (N_2825,N_2125,N_2247);
and U2826 (N_2826,N_2030,N_2388);
and U2827 (N_2827,N_2477,N_2369);
xor U2828 (N_2828,N_2248,N_2070);
or U2829 (N_2829,N_2488,N_2065);
or U2830 (N_2830,N_2424,N_2040);
or U2831 (N_2831,N_2309,N_2054);
and U2832 (N_2832,N_2211,N_2472);
and U2833 (N_2833,N_2389,N_2454);
and U2834 (N_2834,N_2167,N_2433);
and U2835 (N_2835,N_2178,N_2249);
and U2836 (N_2836,N_2375,N_2351);
and U2837 (N_2837,N_2101,N_2362);
or U2838 (N_2838,N_2421,N_2364);
nand U2839 (N_2839,N_2064,N_2034);
nand U2840 (N_2840,N_2486,N_2442);
or U2841 (N_2841,N_2039,N_2142);
and U2842 (N_2842,N_2275,N_2236);
nor U2843 (N_2843,N_2135,N_2204);
nor U2844 (N_2844,N_2215,N_2340);
or U2845 (N_2845,N_2099,N_2158);
or U2846 (N_2846,N_2016,N_2097);
nor U2847 (N_2847,N_2307,N_2395);
nor U2848 (N_2848,N_2299,N_2139);
nand U2849 (N_2849,N_2195,N_2026);
nand U2850 (N_2850,N_2471,N_2122);
and U2851 (N_2851,N_2496,N_2044);
or U2852 (N_2852,N_2400,N_2097);
and U2853 (N_2853,N_2489,N_2181);
and U2854 (N_2854,N_2253,N_2121);
and U2855 (N_2855,N_2208,N_2229);
and U2856 (N_2856,N_2487,N_2234);
nand U2857 (N_2857,N_2128,N_2296);
nand U2858 (N_2858,N_2083,N_2273);
xor U2859 (N_2859,N_2306,N_2421);
and U2860 (N_2860,N_2067,N_2341);
or U2861 (N_2861,N_2227,N_2307);
nand U2862 (N_2862,N_2066,N_2025);
xnor U2863 (N_2863,N_2233,N_2379);
nand U2864 (N_2864,N_2001,N_2436);
or U2865 (N_2865,N_2467,N_2063);
or U2866 (N_2866,N_2191,N_2176);
nand U2867 (N_2867,N_2394,N_2359);
or U2868 (N_2868,N_2235,N_2106);
or U2869 (N_2869,N_2124,N_2137);
xor U2870 (N_2870,N_2142,N_2108);
nand U2871 (N_2871,N_2064,N_2037);
nand U2872 (N_2872,N_2254,N_2261);
xor U2873 (N_2873,N_2374,N_2318);
nand U2874 (N_2874,N_2430,N_2301);
nand U2875 (N_2875,N_2025,N_2492);
xnor U2876 (N_2876,N_2251,N_2009);
or U2877 (N_2877,N_2372,N_2267);
nand U2878 (N_2878,N_2143,N_2475);
nor U2879 (N_2879,N_2372,N_2412);
and U2880 (N_2880,N_2412,N_2316);
nand U2881 (N_2881,N_2006,N_2426);
xor U2882 (N_2882,N_2309,N_2168);
and U2883 (N_2883,N_2419,N_2346);
or U2884 (N_2884,N_2429,N_2336);
or U2885 (N_2885,N_2412,N_2351);
and U2886 (N_2886,N_2385,N_2167);
nor U2887 (N_2887,N_2214,N_2406);
nand U2888 (N_2888,N_2439,N_2222);
nor U2889 (N_2889,N_2200,N_2192);
or U2890 (N_2890,N_2336,N_2372);
or U2891 (N_2891,N_2156,N_2199);
or U2892 (N_2892,N_2198,N_2359);
and U2893 (N_2893,N_2067,N_2238);
or U2894 (N_2894,N_2485,N_2116);
nor U2895 (N_2895,N_2034,N_2074);
or U2896 (N_2896,N_2092,N_2224);
and U2897 (N_2897,N_2264,N_2430);
or U2898 (N_2898,N_2400,N_2188);
nor U2899 (N_2899,N_2171,N_2008);
or U2900 (N_2900,N_2152,N_2256);
or U2901 (N_2901,N_2295,N_2050);
or U2902 (N_2902,N_2354,N_2469);
and U2903 (N_2903,N_2454,N_2003);
or U2904 (N_2904,N_2339,N_2401);
nor U2905 (N_2905,N_2227,N_2329);
or U2906 (N_2906,N_2319,N_2362);
nand U2907 (N_2907,N_2128,N_2251);
or U2908 (N_2908,N_2482,N_2151);
nor U2909 (N_2909,N_2316,N_2168);
nand U2910 (N_2910,N_2273,N_2405);
nor U2911 (N_2911,N_2203,N_2348);
and U2912 (N_2912,N_2006,N_2430);
or U2913 (N_2913,N_2206,N_2096);
xnor U2914 (N_2914,N_2265,N_2239);
nor U2915 (N_2915,N_2237,N_2271);
or U2916 (N_2916,N_2216,N_2490);
and U2917 (N_2917,N_2065,N_2012);
nor U2918 (N_2918,N_2415,N_2094);
nor U2919 (N_2919,N_2080,N_2085);
nor U2920 (N_2920,N_2064,N_2349);
and U2921 (N_2921,N_2028,N_2482);
xnor U2922 (N_2922,N_2435,N_2415);
nand U2923 (N_2923,N_2406,N_2462);
xnor U2924 (N_2924,N_2297,N_2257);
nor U2925 (N_2925,N_2459,N_2276);
nand U2926 (N_2926,N_2322,N_2057);
and U2927 (N_2927,N_2469,N_2326);
and U2928 (N_2928,N_2301,N_2159);
and U2929 (N_2929,N_2492,N_2317);
nand U2930 (N_2930,N_2386,N_2040);
or U2931 (N_2931,N_2463,N_2015);
nor U2932 (N_2932,N_2140,N_2197);
nand U2933 (N_2933,N_2074,N_2135);
or U2934 (N_2934,N_2098,N_2267);
nor U2935 (N_2935,N_2465,N_2262);
nor U2936 (N_2936,N_2217,N_2159);
or U2937 (N_2937,N_2319,N_2364);
xor U2938 (N_2938,N_2184,N_2073);
and U2939 (N_2939,N_2119,N_2154);
or U2940 (N_2940,N_2276,N_2091);
nand U2941 (N_2941,N_2410,N_2158);
xor U2942 (N_2942,N_2336,N_2433);
or U2943 (N_2943,N_2481,N_2429);
xnor U2944 (N_2944,N_2435,N_2062);
or U2945 (N_2945,N_2224,N_2125);
nor U2946 (N_2946,N_2080,N_2372);
xor U2947 (N_2947,N_2404,N_2064);
nor U2948 (N_2948,N_2267,N_2415);
or U2949 (N_2949,N_2118,N_2001);
nor U2950 (N_2950,N_2341,N_2114);
or U2951 (N_2951,N_2012,N_2148);
nor U2952 (N_2952,N_2420,N_2162);
xor U2953 (N_2953,N_2081,N_2003);
or U2954 (N_2954,N_2051,N_2029);
nand U2955 (N_2955,N_2434,N_2149);
nor U2956 (N_2956,N_2324,N_2007);
nor U2957 (N_2957,N_2096,N_2299);
or U2958 (N_2958,N_2484,N_2391);
or U2959 (N_2959,N_2209,N_2351);
or U2960 (N_2960,N_2153,N_2470);
or U2961 (N_2961,N_2480,N_2456);
nor U2962 (N_2962,N_2324,N_2124);
nand U2963 (N_2963,N_2391,N_2049);
and U2964 (N_2964,N_2005,N_2290);
xnor U2965 (N_2965,N_2344,N_2330);
nor U2966 (N_2966,N_2192,N_2250);
nor U2967 (N_2967,N_2158,N_2412);
and U2968 (N_2968,N_2125,N_2005);
nand U2969 (N_2969,N_2453,N_2490);
xnor U2970 (N_2970,N_2152,N_2485);
nand U2971 (N_2971,N_2015,N_2069);
nand U2972 (N_2972,N_2197,N_2342);
nor U2973 (N_2973,N_2115,N_2073);
and U2974 (N_2974,N_2261,N_2009);
nor U2975 (N_2975,N_2235,N_2236);
nand U2976 (N_2976,N_2317,N_2292);
or U2977 (N_2977,N_2274,N_2032);
nand U2978 (N_2978,N_2148,N_2456);
xnor U2979 (N_2979,N_2483,N_2303);
and U2980 (N_2980,N_2108,N_2240);
nor U2981 (N_2981,N_2092,N_2471);
and U2982 (N_2982,N_2254,N_2386);
nor U2983 (N_2983,N_2047,N_2482);
nand U2984 (N_2984,N_2239,N_2311);
nand U2985 (N_2985,N_2167,N_2220);
nor U2986 (N_2986,N_2139,N_2382);
and U2987 (N_2987,N_2330,N_2433);
nor U2988 (N_2988,N_2426,N_2483);
xor U2989 (N_2989,N_2223,N_2122);
and U2990 (N_2990,N_2473,N_2049);
nand U2991 (N_2991,N_2106,N_2051);
nor U2992 (N_2992,N_2380,N_2440);
or U2993 (N_2993,N_2305,N_2333);
or U2994 (N_2994,N_2433,N_2466);
or U2995 (N_2995,N_2079,N_2308);
and U2996 (N_2996,N_2170,N_2262);
nand U2997 (N_2997,N_2044,N_2154);
nand U2998 (N_2998,N_2251,N_2103);
and U2999 (N_2999,N_2276,N_2182);
nor U3000 (N_3000,N_2733,N_2760);
and U3001 (N_3001,N_2938,N_2655);
nor U3002 (N_3002,N_2557,N_2587);
xor U3003 (N_3003,N_2770,N_2727);
nor U3004 (N_3004,N_2973,N_2577);
nor U3005 (N_3005,N_2786,N_2520);
nor U3006 (N_3006,N_2966,N_2512);
and U3007 (N_3007,N_2685,N_2796);
nand U3008 (N_3008,N_2679,N_2736);
or U3009 (N_3009,N_2551,N_2570);
or U3010 (N_3010,N_2673,N_2827);
or U3011 (N_3011,N_2549,N_2757);
or U3012 (N_3012,N_2672,N_2730);
or U3013 (N_3013,N_2921,N_2614);
nand U3014 (N_3014,N_2874,N_2741);
nand U3015 (N_3015,N_2771,N_2682);
nor U3016 (N_3016,N_2828,N_2660);
nand U3017 (N_3017,N_2891,N_2889);
nand U3018 (N_3018,N_2969,N_2820);
nor U3019 (N_3019,N_2962,N_2508);
nor U3020 (N_3020,N_2693,N_2531);
and U3021 (N_3021,N_2671,N_2575);
or U3022 (N_3022,N_2644,N_2562);
nand U3023 (N_3023,N_2568,N_2896);
nand U3024 (N_3024,N_2576,N_2871);
or U3025 (N_3025,N_2635,N_2588);
nand U3026 (N_3026,N_2959,N_2803);
nor U3027 (N_3027,N_2911,N_2968);
or U3028 (N_3028,N_2734,N_2610);
or U3029 (N_3029,N_2514,N_2815);
xnor U3030 (N_3030,N_2952,N_2790);
or U3031 (N_3031,N_2802,N_2859);
xnor U3032 (N_3032,N_2882,N_2768);
nand U3033 (N_3033,N_2515,N_2849);
or U3034 (N_3034,N_2611,N_2728);
and U3035 (N_3035,N_2552,N_2954);
nand U3036 (N_3036,N_2868,N_2569);
nor U3037 (N_3037,N_2763,N_2967);
nor U3038 (N_3038,N_2503,N_2941);
nor U3039 (N_3039,N_2913,N_2524);
and U3040 (N_3040,N_2980,N_2683);
or U3041 (N_3041,N_2637,N_2586);
xor U3042 (N_3042,N_2627,N_2659);
nor U3043 (N_3043,N_2535,N_2858);
nor U3044 (N_3044,N_2695,N_2979);
or U3045 (N_3045,N_2948,N_2875);
nor U3046 (N_3046,N_2582,N_2521);
or U3047 (N_3047,N_2777,N_2840);
nand U3048 (N_3048,N_2804,N_2821);
and U3049 (N_3049,N_2624,N_2657);
nor U3050 (N_3050,N_2932,N_2971);
or U3051 (N_3051,N_2755,N_2940);
xnor U3052 (N_3052,N_2834,N_2511);
nand U3053 (N_3053,N_2878,N_2870);
xor U3054 (N_3054,N_2850,N_2958);
or U3055 (N_3055,N_2539,N_2523);
or U3056 (N_3056,N_2662,N_2795);
nor U3057 (N_3057,N_2892,N_2572);
xor U3058 (N_3058,N_2640,N_2784);
nand U3059 (N_3059,N_2935,N_2960);
or U3060 (N_3060,N_2553,N_2951);
and U3061 (N_3061,N_2782,N_2706);
or U3062 (N_3062,N_2584,N_2857);
and U3063 (N_3063,N_2731,N_2591);
or U3064 (N_3064,N_2925,N_2594);
nor U3065 (N_3065,N_2788,N_2708);
and U3066 (N_3066,N_2919,N_2613);
nor U3067 (N_3067,N_2642,N_2526);
and U3068 (N_3068,N_2534,N_2583);
xnor U3069 (N_3069,N_2801,N_2985);
nand U3070 (N_3070,N_2630,N_2717);
nor U3071 (N_3071,N_2724,N_2691);
or U3072 (N_3072,N_2918,N_2527);
nand U3073 (N_3073,N_2792,N_2654);
xor U3074 (N_3074,N_2785,N_2933);
or U3075 (N_3075,N_2716,N_2965);
nand U3076 (N_3076,N_2797,N_2519);
and U3077 (N_3077,N_2615,N_2603);
nor U3078 (N_3078,N_2560,N_2990);
nor U3079 (N_3079,N_2653,N_2686);
nand U3080 (N_3080,N_2988,N_2561);
and U3081 (N_3081,N_2843,N_2559);
or U3082 (N_3082,N_2664,N_2543);
or U3083 (N_3083,N_2629,N_2705);
nand U3084 (N_3084,N_2643,N_2684);
nor U3085 (N_3085,N_2722,N_2528);
xor U3086 (N_3086,N_2749,N_2608);
nand U3087 (N_3087,N_2818,N_2983);
nor U3088 (N_3088,N_2548,N_2981);
nor U3089 (N_3089,N_2928,N_2595);
or U3090 (N_3090,N_2725,N_2856);
nand U3091 (N_3091,N_2670,N_2977);
and U3092 (N_3092,N_2620,N_2754);
or U3093 (N_3093,N_2929,N_2863);
and U3094 (N_3094,N_2982,N_2632);
or U3095 (N_3095,N_2937,N_2813);
or U3096 (N_3096,N_2530,N_2694);
or U3097 (N_3097,N_2502,N_2590);
and U3098 (N_3098,N_2837,N_2602);
and U3099 (N_3099,N_2574,N_2809);
nor U3100 (N_3100,N_2573,N_2905);
or U3101 (N_3101,N_2677,N_2789);
xnor U3102 (N_3102,N_2961,N_2793);
nand U3103 (N_3103,N_2645,N_2712);
and U3104 (N_3104,N_2661,N_2752);
xnor U3105 (N_3105,N_2510,N_2646);
nand U3106 (N_3106,N_2914,N_2832);
nor U3107 (N_3107,N_2987,N_2893);
nor U3108 (N_3108,N_2970,N_2751);
and U3109 (N_3109,N_2810,N_2864);
or U3110 (N_3110,N_2920,N_2545);
or U3111 (N_3111,N_2869,N_2668);
nand U3112 (N_3112,N_2743,N_2887);
xnor U3113 (N_3113,N_2989,N_2541);
and U3114 (N_3114,N_2773,N_2689);
xnor U3115 (N_3115,N_2996,N_2634);
nand U3116 (N_3116,N_2740,N_2908);
xnor U3117 (N_3117,N_2579,N_2723);
and U3118 (N_3118,N_2844,N_2702);
and U3119 (N_3119,N_2852,N_2778);
nand U3120 (N_3120,N_2907,N_2978);
nand U3121 (N_3121,N_2604,N_2711);
xor U3122 (N_3122,N_2715,N_2898);
nor U3123 (N_3123,N_2862,N_2639);
xnor U3124 (N_3124,N_2881,N_2822);
and U3125 (N_3125,N_2894,N_2794);
nor U3126 (N_3126,N_2533,N_2589);
xnor U3127 (N_3127,N_2936,N_2550);
nor U3128 (N_3128,N_2994,N_2900);
nand U3129 (N_3129,N_2816,N_2769);
nand U3130 (N_3130,N_2904,N_2872);
or U3131 (N_3131,N_2963,N_2903);
nor U3132 (N_3132,N_2934,N_2578);
nor U3133 (N_3133,N_2707,N_2890);
and U3134 (N_3134,N_2866,N_2943);
nor U3135 (N_3135,N_2565,N_2955);
and U3136 (N_3136,N_2732,N_2656);
and U3137 (N_3137,N_2747,N_2580);
nor U3138 (N_3138,N_2688,N_2667);
and U3139 (N_3139,N_2901,N_2621);
or U3140 (N_3140,N_2529,N_2687);
or U3141 (N_3141,N_2525,N_2842);
or U3142 (N_3142,N_2623,N_2719);
or U3143 (N_3143,N_2501,N_2504);
and U3144 (N_3144,N_2993,N_2616);
nand U3145 (N_3145,N_2759,N_2556);
and U3146 (N_3146,N_2819,N_2532);
nand U3147 (N_3147,N_2841,N_2945);
and U3148 (N_3148,N_2772,N_2617);
or U3149 (N_3149,N_2947,N_2555);
or U3150 (N_3150,N_2665,N_2876);
or U3151 (N_3151,N_2593,N_2867);
nand U3152 (N_3152,N_2697,N_2956);
or U3153 (N_3153,N_2991,N_2767);
or U3154 (N_3154,N_2780,N_2814);
or U3155 (N_3155,N_2998,N_2571);
xor U3156 (N_3156,N_2839,N_2781);
nand U3157 (N_3157,N_2746,N_2944);
nor U3158 (N_3158,N_2618,N_2651);
nor U3159 (N_3159,N_2883,N_2600);
and U3160 (N_3160,N_2675,N_2817);
and U3161 (N_3161,N_2748,N_2704);
or U3162 (N_3162,N_2585,N_2681);
and U3163 (N_3163,N_2917,N_2544);
or U3164 (N_3164,N_2791,N_2811);
and U3165 (N_3165,N_2984,N_2765);
nor U3166 (N_3166,N_2674,N_2631);
and U3167 (N_3167,N_2753,N_2877);
and U3168 (N_3168,N_2658,N_2606);
or U3169 (N_3169,N_2676,N_2564);
nand U3170 (N_3170,N_2592,N_2879);
xnor U3171 (N_3171,N_2729,N_2536);
xor U3172 (N_3172,N_2601,N_2666);
nand U3173 (N_3173,N_2692,N_2957);
nand U3174 (N_3174,N_2546,N_2513);
or U3175 (N_3175,N_2720,N_2829);
xnor U3176 (N_3176,N_2902,N_2854);
nor U3177 (N_3177,N_2847,N_2974);
and U3178 (N_3178,N_2744,N_2783);
xnor U3179 (N_3179,N_2507,N_2709);
and U3180 (N_3180,N_2516,N_2915);
nand U3181 (N_3181,N_2779,N_2718);
or U3182 (N_3182,N_2865,N_2848);
nor U3183 (N_3183,N_2846,N_2851);
or U3184 (N_3184,N_2800,N_2946);
or U3185 (N_3185,N_2949,N_2537);
or U3186 (N_3186,N_2899,N_2505);
nand U3187 (N_3187,N_2517,N_2652);
nor U3188 (N_3188,N_2897,N_2776);
nor U3189 (N_3189,N_2999,N_2647);
or U3190 (N_3190,N_2500,N_2823);
or U3191 (N_3191,N_2703,N_2745);
nand U3192 (N_3192,N_2597,N_2906);
nor U3193 (N_3193,N_2599,N_2638);
xnor U3194 (N_3194,N_2563,N_2538);
nand U3195 (N_3195,N_2805,N_2622);
or U3196 (N_3196,N_2806,N_2607);
nand U3197 (N_3197,N_2895,N_2710);
nor U3198 (N_3198,N_2787,N_2721);
or U3199 (N_3199,N_2542,N_2737);
nand U3200 (N_3200,N_2626,N_2714);
nand U3201 (N_3201,N_2700,N_2910);
or U3202 (N_3202,N_2750,N_2649);
nand U3203 (N_3203,N_2764,N_2888);
nand U3204 (N_3204,N_2986,N_2761);
or U3205 (N_3205,N_2880,N_2742);
or U3206 (N_3206,N_2824,N_2884);
nand U3207 (N_3207,N_2738,N_2964);
and U3208 (N_3208,N_2726,N_2581);
nor U3209 (N_3209,N_2633,N_2833);
xnor U3210 (N_3210,N_2855,N_2663);
nor U3211 (N_3211,N_2930,N_2845);
xnor U3212 (N_3212,N_2812,N_2598);
and U3213 (N_3213,N_2506,N_2554);
or U3214 (N_3214,N_2836,N_2774);
or U3215 (N_3215,N_2873,N_2923);
xnor U3216 (N_3216,N_2972,N_2926);
or U3217 (N_3217,N_2636,N_2853);
and U3218 (N_3218,N_2558,N_2838);
xnor U3219 (N_3219,N_2825,N_2912);
and U3220 (N_3220,N_2885,N_2950);
or U3221 (N_3221,N_2758,N_2808);
nor U3222 (N_3222,N_2830,N_2775);
and U3223 (N_3223,N_2690,N_2975);
or U3224 (N_3224,N_2916,N_2992);
or U3225 (N_3225,N_2861,N_2995);
or U3226 (N_3226,N_2713,N_2518);
or U3227 (N_3227,N_2680,N_2567);
or U3228 (N_3228,N_2669,N_2924);
and U3229 (N_3229,N_2596,N_2698);
xor U3230 (N_3230,N_2927,N_2735);
or U3231 (N_3231,N_2701,N_2547);
or U3232 (N_3232,N_2997,N_2609);
nor U3233 (N_3233,N_2766,N_2619);
or U3234 (N_3234,N_2831,N_2566);
or U3235 (N_3235,N_2605,N_2886);
or U3236 (N_3236,N_2909,N_2931);
and U3237 (N_3237,N_2860,N_2678);
nand U3238 (N_3238,N_2942,N_2699);
nor U3239 (N_3239,N_2762,N_2540);
and U3240 (N_3240,N_2826,N_2798);
nor U3241 (N_3241,N_2628,N_2522);
nand U3242 (N_3242,N_2648,N_2953);
nor U3243 (N_3243,N_2939,N_2976);
nor U3244 (N_3244,N_2641,N_2650);
nand U3245 (N_3245,N_2922,N_2807);
nand U3246 (N_3246,N_2612,N_2756);
or U3247 (N_3247,N_2799,N_2696);
xnor U3248 (N_3248,N_2625,N_2509);
and U3249 (N_3249,N_2739,N_2835);
and U3250 (N_3250,N_2678,N_2796);
or U3251 (N_3251,N_2575,N_2844);
or U3252 (N_3252,N_2866,N_2732);
nand U3253 (N_3253,N_2770,N_2761);
or U3254 (N_3254,N_2967,N_2907);
or U3255 (N_3255,N_2546,N_2686);
nand U3256 (N_3256,N_2611,N_2703);
xor U3257 (N_3257,N_2991,N_2546);
nand U3258 (N_3258,N_2624,N_2980);
nand U3259 (N_3259,N_2932,N_2661);
nand U3260 (N_3260,N_2588,N_2798);
and U3261 (N_3261,N_2712,N_2961);
nand U3262 (N_3262,N_2580,N_2533);
or U3263 (N_3263,N_2714,N_2713);
or U3264 (N_3264,N_2588,N_2611);
nand U3265 (N_3265,N_2901,N_2724);
xnor U3266 (N_3266,N_2966,N_2636);
and U3267 (N_3267,N_2745,N_2657);
xnor U3268 (N_3268,N_2678,N_2741);
nor U3269 (N_3269,N_2599,N_2661);
nand U3270 (N_3270,N_2924,N_2532);
nor U3271 (N_3271,N_2805,N_2726);
xnor U3272 (N_3272,N_2574,N_2969);
and U3273 (N_3273,N_2996,N_2714);
nor U3274 (N_3274,N_2801,N_2678);
nand U3275 (N_3275,N_2815,N_2905);
nor U3276 (N_3276,N_2522,N_2990);
or U3277 (N_3277,N_2777,N_2984);
nor U3278 (N_3278,N_2656,N_2696);
and U3279 (N_3279,N_2685,N_2873);
nor U3280 (N_3280,N_2891,N_2951);
nand U3281 (N_3281,N_2659,N_2501);
or U3282 (N_3282,N_2655,N_2840);
nor U3283 (N_3283,N_2858,N_2821);
xnor U3284 (N_3284,N_2964,N_2691);
nor U3285 (N_3285,N_2728,N_2988);
nand U3286 (N_3286,N_2607,N_2781);
nand U3287 (N_3287,N_2663,N_2804);
or U3288 (N_3288,N_2671,N_2916);
xnor U3289 (N_3289,N_2643,N_2681);
or U3290 (N_3290,N_2845,N_2679);
nand U3291 (N_3291,N_2994,N_2899);
nor U3292 (N_3292,N_2954,N_2844);
and U3293 (N_3293,N_2611,N_2857);
xor U3294 (N_3294,N_2687,N_2614);
or U3295 (N_3295,N_2575,N_2517);
or U3296 (N_3296,N_2609,N_2773);
xor U3297 (N_3297,N_2582,N_2748);
and U3298 (N_3298,N_2603,N_2706);
nor U3299 (N_3299,N_2598,N_2871);
or U3300 (N_3300,N_2977,N_2766);
nand U3301 (N_3301,N_2906,N_2691);
and U3302 (N_3302,N_2947,N_2752);
nor U3303 (N_3303,N_2570,N_2502);
or U3304 (N_3304,N_2818,N_2740);
and U3305 (N_3305,N_2831,N_2527);
nor U3306 (N_3306,N_2508,N_2868);
nand U3307 (N_3307,N_2781,N_2566);
nand U3308 (N_3308,N_2644,N_2982);
nor U3309 (N_3309,N_2814,N_2545);
and U3310 (N_3310,N_2734,N_2862);
xnor U3311 (N_3311,N_2585,N_2997);
and U3312 (N_3312,N_2966,N_2699);
or U3313 (N_3313,N_2550,N_2883);
or U3314 (N_3314,N_2981,N_2858);
nand U3315 (N_3315,N_2950,N_2542);
nor U3316 (N_3316,N_2656,N_2510);
nor U3317 (N_3317,N_2813,N_2849);
or U3318 (N_3318,N_2788,N_2682);
nor U3319 (N_3319,N_2668,N_2865);
nand U3320 (N_3320,N_2766,N_2740);
and U3321 (N_3321,N_2542,N_2999);
or U3322 (N_3322,N_2895,N_2965);
and U3323 (N_3323,N_2599,N_2554);
nand U3324 (N_3324,N_2897,N_2600);
nand U3325 (N_3325,N_2998,N_2890);
or U3326 (N_3326,N_2573,N_2999);
and U3327 (N_3327,N_2868,N_2557);
or U3328 (N_3328,N_2589,N_2510);
and U3329 (N_3329,N_2940,N_2769);
or U3330 (N_3330,N_2542,N_2543);
xnor U3331 (N_3331,N_2702,N_2982);
nor U3332 (N_3332,N_2896,N_2645);
nor U3333 (N_3333,N_2572,N_2885);
nand U3334 (N_3334,N_2923,N_2918);
nor U3335 (N_3335,N_2757,N_2854);
nor U3336 (N_3336,N_2892,N_2650);
or U3337 (N_3337,N_2626,N_2775);
or U3338 (N_3338,N_2807,N_2517);
or U3339 (N_3339,N_2591,N_2578);
nand U3340 (N_3340,N_2676,N_2602);
and U3341 (N_3341,N_2724,N_2508);
or U3342 (N_3342,N_2675,N_2983);
or U3343 (N_3343,N_2854,N_2977);
nand U3344 (N_3344,N_2608,N_2542);
or U3345 (N_3345,N_2971,N_2883);
nand U3346 (N_3346,N_2765,N_2565);
nor U3347 (N_3347,N_2592,N_2718);
nand U3348 (N_3348,N_2966,N_2506);
nor U3349 (N_3349,N_2619,N_2627);
nand U3350 (N_3350,N_2665,N_2799);
xor U3351 (N_3351,N_2874,N_2887);
nand U3352 (N_3352,N_2613,N_2907);
nand U3353 (N_3353,N_2637,N_2866);
and U3354 (N_3354,N_2626,N_2533);
or U3355 (N_3355,N_2762,N_2895);
nor U3356 (N_3356,N_2884,N_2631);
or U3357 (N_3357,N_2796,N_2562);
nand U3358 (N_3358,N_2913,N_2683);
nor U3359 (N_3359,N_2886,N_2638);
nor U3360 (N_3360,N_2875,N_2637);
or U3361 (N_3361,N_2663,N_2737);
and U3362 (N_3362,N_2873,N_2517);
nand U3363 (N_3363,N_2986,N_2700);
xor U3364 (N_3364,N_2971,N_2927);
nor U3365 (N_3365,N_2820,N_2587);
xnor U3366 (N_3366,N_2935,N_2782);
or U3367 (N_3367,N_2830,N_2932);
nor U3368 (N_3368,N_2942,N_2951);
nand U3369 (N_3369,N_2863,N_2744);
nand U3370 (N_3370,N_2782,N_2984);
xor U3371 (N_3371,N_2787,N_2567);
or U3372 (N_3372,N_2953,N_2852);
and U3373 (N_3373,N_2578,N_2839);
or U3374 (N_3374,N_2829,N_2708);
or U3375 (N_3375,N_2983,N_2902);
or U3376 (N_3376,N_2876,N_2592);
or U3377 (N_3377,N_2514,N_2862);
nand U3378 (N_3378,N_2994,N_2993);
and U3379 (N_3379,N_2738,N_2537);
or U3380 (N_3380,N_2906,N_2942);
nand U3381 (N_3381,N_2853,N_2563);
and U3382 (N_3382,N_2643,N_2670);
nand U3383 (N_3383,N_2575,N_2775);
nor U3384 (N_3384,N_2542,N_2586);
nor U3385 (N_3385,N_2833,N_2988);
nor U3386 (N_3386,N_2860,N_2517);
and U3387 (N_3387,N_2521,N_2686);
xnor U3388 (N_3388,N_2546,N_2886);
and U3389 (N_3389,N_2793,N_2594);
and U3390 (N_3390,N_2860,N_2560);
nand U3391 (N_3391,N_2924,N_2732);
or U3392 (N_3392,N_2768,N_2536);
nand U3393 (N_3393,N_2550,N_2623);
or U3394 (N_3394,N_2571,N_2510);
or U3395 (N_3395,N_2750,N_2677);
or U3396 (N_3396,N_2835,N_2726);
and U3397 (N_3397,N_2598,N_2650);
or U3398 (N_3398,N_2831,N_2645);
nor U3399 (N_3399,N_2972,N_2736);
or U3400 (N_3400,N_2928,N_2955);
or U3401 (N_3401,N_2553,N_2955);
nand U3402 (N_3402,N_2709,N_2516);
and U3403 (N_3403,N_2716,N_2955);
nor U3404 (N_3404,N_2984,N_2885);
nor U3405 (N_3405,N_2920,N_2608);
nor U3406 (N_3406,N_2849,N_2627);
nor U3407 (N_3407,N_2943,N_2869);
xnor U3408 (N_3408,N_2610,N_2926);
nand U3409 (N_3409,N_2681,N_2937);
and U3410 (N_3410,N_2856,N_2655);
and U3411 (N_3411,N_2771,N_2607);
or U3412 (N_3412,N_2547,N_2662);
nor U3413 (N_3413,N_2523,N_2679);
nand U3414 (N_3414,N_2785,N_2637);
nor U3415 (N_3415,N_2772,N_2663);
nand U3416 (N_3416,N_2712,N_2673);
or U3417 (N_3417,N_2935,N_2649);
nor U3418 (N_3418,N_2540,N_2881);
nand U3419 (N_3419,N_2639,N_2642);
or U3420 (N_3420,N_2670,N_2828);
xor U3421 (N_3421,N_2851,N_2741);
nand U3422 (N_3422,N_2869,N_2786);
xnor U3423 (N_3423,N_2907,N_2656);
nor U3424 (N_3424,N_2868,N_2948);
nand U3425 (N_3425,N_2831,N_2658);
nor U3426 (N_3426,N_2696,N_2562);
and U3427 (N_3427,N_2919,N_2850);
or U3428 (N_3428,N_2761,N_2795);
xor U3429 (N_3429,N_2717,N_2521);
nor U3430 (N_3430,N_2517,N_2653);
nor U3431 (N_3431,N_2875,N_2651);
and U3432 (N_3432,N_2675,N_2796);
and U3433 (N_3433,N_2669,N_2713);
and U3434 (N_3434,N_2661,N_2911);
nor U3435 (N_3435,N_2904,N_2661);
nor U3436 (N_3436,N_2693,N_2566);
nand U3437 (N_3437,N_2891,N_2586);
and U3438 (N_3438,N_2936,N_2543);
and U3439 (N_3439,N_2849,N_2918);
and U3440 (N_3440,N_2706,N_2929);
nand U3441 (N_3441,N_2669,N_2749);
xor U3442 (N_3442,N_2808,N_2599);
nand U3443 (N_3443,N_2745,N_2674);
nor U3444 (N_3444,N_2872,N_2978);
nor U3445 (N_3445,N_2903,N_2740);
nor U3446 (N_3446,N_2653,N_2730);
or U3447 (N_3447,N_2645,N_2515);
nor U3448 (N_3448,N_2708,N_2742);
xnor U3449 (N_3449,N_2873,N_2701);
and U3450 (N_3450,N_2791,N_2874);
and U3451 (N_3451,N_2843,N_2543);
nor U3452 (N_3452,N_2892,N_2668);
or U3453 (N_3453,N_2925,N_2915);
nand U3454 (N_3454,N_2982,N_2760);
or U3455 (N_3455,N_2932,N_2621);
nand U3456 (N_3456,N_2618,N_2615);
nand U3457 (N_3457,N_2712,N_2519);
and U3458 (N_3458,N_2910,N_2716);
nand U3459 (N_3459,N_2694,N_2830);
or U3460 (N_3460,N_2744,N_2993);
nand U3461 (N_3461,N_2853,N_2728);
nand U3462 (N_3462,N_2889,N_2656);
nand U3463 (N_3463,N_2757,N_2874);
or U3464 (N_3464,N_2793,N_2843);
nand U3465 (N_3465,N_2986,N_2963);
nor U3466 (N_3466,N_2881,N_2621);
and U3467 (N_3467,N_2795,N_2826);
or U3468 (N_3468,N_2645,N_2646);
or U3469 (N_3469,N_2944,N_2965);
nand U3470 (N_3470,N_2775,N_2609);
or U3471 (N_3471,N_2942,N_2554);
nor U3472 (N_3472,N_2891,N_2697);
or U3473 (N_3473,N_2879,N_2905);
nor U3474 (N_3474,N_2901,N_2924);
or U3475 (N_3475,N_2748,N_2568);
nand U3476 (N_3476,N_2774,N_2807);
nor U3477 (N_3477,N_2698,N_2785);
and U3478 (N_3478,N_2841,N_2809);
nor U3479 (N_3479,N_2995,N_2531);
nand U3480 (N_3480,N_2932,N_2736);
nor U3481 (N_3481,N_2584,N_2707);
or U3482 (N_3482,N_2835,N_2931);
xnor U3483 (N_3483,N_2894,N_2679);
and U3484 (N_3484,N_2854,N_2692);
or U3485 (N_3485,N_2934,N_2748);
nand U3486 (N_3486,N_2891,N_2917);
and U3487 (N_3487,N_2944,N_2733);
nand U3488 (N_3488,N_2794,N_2603);
or U3489 (N_3489,N_2793,N_2526);
nor U3490 (N_3490,N_2986,N_2550);
nand U3491 (N_3491,N_2698,N_2806);
and U3492 (N_3492,N_2693,N_2842);
or U3493 (N_3493,N_2522,N_2502);
nor U3494 (N_3494,N_2597,N_2957);
nor U3495 (N_3495,N_2664,N_2751);
nand U3496 (N_3496,N_2967,N_2552);
and U3497 (N_3497,N_2513,N_2601);
xnor U3498 (N_3498,N_2707,N_2624);
nor U3499 (N_3499,N_2966,N_2663);
nand U3500 (N_3500,N_3011,N_3353);
nand U3501 (N_3501,N_3199,N_3080);
or U3502 (N_3502,N_3132,N_3244);
nor U3503 (N_3503,N_3002,N_3072);
or U3504 (N_3504,N_3198,N_3492);
and U3505 (N_3505,N_3335,N_3484);
or U3506 (N_3506,N_3041,N_3166);
and U3507 (N_3507,N_3315,N_3326);
nor U3508 (N_3508,N_3396,N_3471);
and U3509 (N_3509,N_3025,N_3460);
and U3510 (N_3510,N_3454,N_3228);
nor U3511 (N_3511,N_3232,N_3048);
and U3512 (N_3512,N_3256,N_3393);
nand U3513 (N_3513,N_3026,N_3230);
and U3514 (N_3514,N_3224,N_3445);
nand U3515 (N_3515,N_3419,N_3434);
xnor U3516 (N_3516,N_3075,N_3014);
xor U3517 (N_3517,N_3069,N_3307);
nand U3518 (N_3518,N_3033,N_3358);
or U3519 (N_3519,N_3062,N_3263);
nor U3520 (N_3520,N_3451,N_3091);
nand U3521 (N_3521,N_3010,N_3064);
nor U3522 (N_3522,N_3212,N_3137);
nand U3523 (N_3523,N_3438,N_3389);
or U3524 (N_3524,N_3397,N_3238);
or U3525 (N_3525,N_3104,N_3441);
or U3526 (N_3526,N_3371,N_3270);
or U3527 (N_3527,N_3117,N_3017);
nand U3528 (N_3528,N_3098,N_3233);
or U3529 (N_3529,N_3257,N_3405);
nand U3530 (N_3530,N_3314,N_3465);
or U3531 (N_3531,N_3400,N_3290);
nand U3532 (N_3532,N_3184,N_3413);
and U3533 (N_3533,N_3076,N_3443);
and U3534 (N_3534,N_3142,N_3071);
or U3535 (N_3535,N_3031,N_3399);
and U3536 (N_3536,N_3188,N_3096);
and U3537 (N_3537,N_3032,N_3466);
nor U3538 (N_3538,N_3209,N_3280);
nor U3539 (N_3539,N_3266,N_3177);
nor U3540 (N_3540,N_3324,N_3346);
nand U3541 (N_3541,N_3052,N_3255);
nand U3542 (N_3542,N_3489,N_3424);
and U3543 (N_3543,N_3126,N_3455);
or U3544 (N_3544,N_3370,N_3106);
or U3545 (N_3545,N_3007,N_3412);
or U3546 (N_3546,N_3247,N_3368);
or U3547 (N_3547,N_3302,N_3019);
or U3548 (N_3548,N_3216,N_3361);
xnor U3549 (N_3549,N_3388,N_3356);
or U3550 (N_3550,N_3220,N_3201);
and U3551 (N_3551,N_3488,N_3254);
nor U3552 (N_3552,N_3057,N_3494);
or U3553 (N_3553,N_3428,N_3487);
nor U3554 (N_3554,N_3380,N_3322);
and U3555 (N_3555,N_3083,N_3248);
or U3556 (N_3556,N_3284,N_3016);
nand U3557 (N_3557,N_3459,N_3359);
and U3558 (N_3558,N_3447,N_3294);
nor U3559 (N_3559,N_3024,N_3340);
xor U3560 (N_3560,N_3476,N_3360);
nand U3561 (N_3561,N_3190,N_3196);
or U3562 (N_3562,N_3470,N_3114);
or U3563 (N_3563,N_3179,N_3097);
nand U3564 (N_3564,N_3279,N_3180);
nand U3565 (N_3565,N_3474,N_3036);
nand U3566 (N_3566,N_3049,N_3246);
nand U3567 (N_3567,N_3486,N_3274);
or U3568 (N_3568,N_3392,N_3418);
and U3569 (N_3569,N_3289,N_3386);
nand U3570 (N_3570,N_3009,N_3185);
nor U3571 (N_3571,N_3429,N_3108);
nor U3572 (N_3572,N_3350,N_3176);
or U3573 (N_3573,N_3136,N_3181);
and U3574 (N_3574,N_3164,N_3303);
or U3575 (N_3575,N_3194,N_3433);
nand U3576 (N_3576,N_3450,N_3008);
nand U3577 (N_3577,N_3165,N_3205);
xor U3578 (N_3578,N_3195,N_3367);
nor U3579 (N_3579,N_3403,N_3141);
or U3580 (N_3580,N_3125,N_3401);
nor U3581 (N_3581,N_3312,N_3225);
or U3582 (N_3582,N_3309,N_3021);
nand U3583 (N_3583,N_3050,N_3187);
nand U3584 (N_3584,N_3480,N_3300);
or U3585 (N_3585,N_3219,N_3310);
nand U3586 (N_3586,N_3102,N_3252);
nor U3587 (N_3587,N_3223,N_3366);
nand U3588 (N_3588,N_3497,N_3332);
and U3589 (N_3589,N_3153,N_3053);
and U3590 (N_3590,N_3395,N_3373);
nor U3591 (N_3591,N_3063,N_3375);
or U3592 (N_3592,N_3409,N_3065);
or U3593 (N_3593,N_3156,N_3134);
nor U3594 (N_3594,N_3160,N_3140);
and U3595 (N_3595,N_3426,N_3382);
and U3596 (N_3596,N_3234,N_3264);
and U3597 (N_3597,N_3121,N_3200);
xnor U3598 (N_3598,N_3155,N_3088);
nand U3599 (N_3599,N_3059,N_3038);
nand U3600 (N_3600,N_3079,N_3328);
nand U3601 (N_3601,N_3407,N_3425);
and U3602 (N_3602,N_3214,N_3092);
nand U3603 (N_3603,N_3319,N_3211);
or U3604 (N_3604,N_3369,N_3437);
nand U3605 (N_3605,N_3068,N_3472);
or U3606 (N_3606,N_3491,N_3272);
and U3607 (N_3607,N_3404,N_3352);
nor U3608 (N_3608,N_3464,N_3111);
nand U3609 (N_3609,N_3456,N_3498);
nand U3610 (N_3610,N_3336,N_3318);
or U3611 (N_3611,N_3215,N_3051);
nor U3612 (N_3612,N_3151,N_3414);
xnor U3613 (N_3613,N_3305,N_3005);
xnor U3614 (N_3614,N_3182,N_3150);
nor U3615 (N_3615,N_3135,N_3422);
and U3616 (N_3616,N_3331,N_3448);
nand U3617 (N_3617,N_3202,N_3093);
and U3618 (N_3618,N_3119,N_3210);
nand U3619 (N_3619,N_3139,N_3327);
xor U3620 (N_3620,N_3285,N_3461);
nand U3621 (N_3621,N_3301,N_3431);
and U3622 (N_3622,N_3192,N_3143);
and U3623 (N_3623,N_3056,N_3261);
nor U3624 (N_3624,N_3090,N_3226);
nor U3625 (N_3625,N_3169,N_3073);
or U3626 (N_3626,N_3325,N_3145);
or U3627 (N_3627,N_3457,N_3020);
and U3628 (N_3628,N_3162,N_3415);
or U3629 (N_3629,N_3377,N_3197);
and U3630 (N_3630,N_3341,N_3376);
and U3631 (N_3631,N_3402,N_3094);
or U3632 (N_3632,N_3107,N_3082);
nor U3633 (N_3633,N_3317,N_3449);
and U3634 (N_3634,N_3446,N_3178);
nor U3635 (N_3635,N_3334,N_3030);
nand U3636 (N_3636,N_3243,N_3027);
nor U3637 (N_3637,N_3146,N_3453);
or U3638 (N_3638,N_3235,N_3439);
or U3639 (N_3639,N_3384,N_3183);
or U3640 (N_3640,N_3269,N_3262);
xnor U3641 (N_3641,N_3138,N_3365);
nand U3642 (N_3642,N_3168,N_3105);
and U3643 (N_3643,N_3206,N_3089);
nand U3644 (N_3644,N_3112,N_3163);
or U3645 (N_3645,N_3251,N_3042);
xnor U3646 (N_3646,N_3440,N_3004);
xnor U3647 (N_3647,N_3203,N_3249);
nand U3648 (N_3648,N_3286,N_3193);
and U3649 (N_3649,N_3171,N_3159);
or U3650 (N_3650,N_3046,N_3345);
xor U3651 (N_3651,N_3043,N_3174);
nor U3652 (N_3652,N_3333,N_3385);
nand U3653 (N_3653,N_3374,N_3351);
or U3654 (N_3654,N_3283,N_3311);
or U3655 (N_3655,N_3070,N_3158);
nor U3656 (N_3656,N_3003,N_3291);
and U3657 (N_3657,N_3394,N_3013);
nor U3658 (N_3658,N_3320,N_3250);
or U3659 (N_3659,N_3410,N_3085);
or U3660 (N_3660,N_3330,N_3271);
and U3661 (N_3661,N_3006,N_3306);
xor U3662 (N_3662,N_3287,N_3344);
nand U3663 (N_3663,N_3435,N_3436);
and U3664 (N_3664,N_3095,N_3278);
nand U3665 (N_3665,N_3242,N_3275);
nand U3666 (N_3666,N_3044,N_3313);
nand U3667 (N_3667,N_3118,N_3276);
nor U3668 (N_3668,N_3468,N_3147);
nor U3669 (N_3669,N_3122,N_3040);
nand U3670 (N_3670,N_3478,N_3084);
or U3671 (N_3671,N_3288,N_3390);
nand U3672 (N_3672,N_3229,N_3028);
and U3673 (N_3673,N_3175,N_3208);
nor U3674 (N_3674,N_3423,N_3308);
or U3675 (N_3675,N_3259,N_3293);
or U3676 (N_3676,N_3129,N_3124);
nand U3677 (N_3677,N_3000,N_3152);
xnor U3678 (N_3678,N_3265,N_3037);
or U3679 (N_3679,N_3001,N_3022);
nand U3680 (N_3680,N_3035,N_3482);
nand U3681 (N_3681,N_3128,N_3061);
nand U3682 (N_3682,N_3496,N_3100);
nor U3683 (N_3683,N_3493,N_3387);
xnor U3684 (N_3684,N_3477,N_3469);
nand U3685 (N_3685,N_3338,N_3191);
or U3686 (N_3686,N_3292,N_3499);
nor U3687 (N_3687,N_3149,N_3329);
nor U3688 (N_3688,N_3029,N_3207);
and U3689 (N_3689,N_3458,N_3054);
nand U3690 (N_3690,N_3161,N_3495);
and U3691 (N_3691,N_3120,N_3258);
nor U3692 (N_3692,N_3170,N_3227);
nor U3693 (N_3693,N_3239,N_3167);
or U3694 (N_3694,N_3157,N_3267);
or U3695 (N_3695,N_3012,N_3347);
xor U3696 (N_3696,N_3273,N_3357);
nor U3697 (N_3697,N_3115,N_3066);
xor U3698 (N_3698,N_3463,N_3427);
or U3699 (N_3699,N_3099,N_3133);
nand U3700 (N_3700,N_3372,N_3067);
or U3701 (N_3701,N_3483,N_3213);
xor U3702 (N_3702,N_3343,N_3381);
or U3703 (N_3703,N_3110,N_3236);
and U3704 (N_3704,N_3131,N_3296);
nor U3705 (N_3705,N_3481,N_3268);
or U3706 (N_3706,N_3354,N_3045);
nor U3707 (N_3707,N_3241,N_3060);
or U3708 (N_3708,N_3467,N_3015);
and U3709 (N_3709,N_3101,N_3408);
xnor U3710 (N_3710,N_3452,N_3047);
nand U3711 (N_3711,N_3485,N_3023);
and U3712 (N_3712,N_3087,N_3339);
or U3713 (N_3713,N_3420,N_3416);
or U3714 (N_3714,N_3034,N_3245);
nand U3715 (N_3715,N_3282,N_3074);
nor U3716 (N_3716,N_3154,N_3109);
or U3717 (N_3717,N_3260,N_3406);
nor U3718 (N_3718,N_3304,N_3417);
nor U3719 (N_3719,N_3081,N_3411);
nor U3720 (N_3720,N_3173,N_3475);
nand U3721 (N_3721,N_3355,N_3362);
nand U3722 (N_3722,N_3363,N_3473);
nor U3723 (N_3723,N_3444,N_3297);
nor U3724 (N_3724,N_3172,N_3337);
xnor U3725 (N_3725,N_3295,N_3123);
xnor U3726 (N_3726,N_3432,N_3113);
or U3727 (N_3727,N_3349,N_3421);
nor U3728 (N_3728,N_3391,N_3442);
nand U3729 (N_3729,N_3018,N_3221);
or U3730 (N_3730,N_3144,N_3058);
nor U3731 (N_3731,N_3237,N_3342);
xor U3732 (N_3732,N_3379,N_3298);
or U3733 (N_3733,N_3148,N_3231);
nor U3734 (N_3734,N_3316,N_3086);
and U3735 (N_3735,N_3490,N_3217);
nor U3736 (N_3736,N_3055,N_3116);
and U3737 (N_3737,N_3383,N_3321);
xnor U3738 (N_3738,N_3039,N_3398);
nand U3739 (N_3739,N_3078,N_3103);
or U3740 (N_3740,N_3299,N_3240);
or U3741 (N_3741,N_3204,N_3323);
nand U3742 (N_3742,N_3430,N_3130);
nand U3743 (N_3743,N_3186,N_3462);
or U3744 (N_3744,N_3378,N_3281);
nor U3745 (N_3745,N_3277,N_3218);
nor U3746 (N_3746,N_3348,N_3364);
and U3747 (N_3747,N_3253,N_3127);
and U3748 (N_3748,N_3189,N_3479);
and U3749 (N_3749,N_3222,N_3077);
or U3750 (N_3750,N_3033,N_3365);
nor U3751 (N_3751,N_3149,N_3074);
and U3752 (N_3752,N_3193,N_3141);
nor U3753 (N_3753,N_3472,N_3016);
and U3754 (N_3754,N_3421,N_3109);
nand U3755 (N_3755,N_3184,N_3032);
and U3756 (N_3756,N_3290,N_3197);
nand U3757 (N_3757,N_3424,N_3047);
or U3758 (N_3758,N_3383,N_3297);
nand U3759 (N_3759,N_3306,N_3322);
or U3760 (N_3760,N_3014,N_3170);
nor U3761 (N_3761,N_3050,N_3436);
xnor U3762 (N_3762,N_3310,N_3287);
or U3763 (N_3763,N_3179,N_3165);
nor U3764 (N_3764,N_3173,N_3471);
nand U3765 (N_3765,N_3254,N_3394);
nor U3766 (N_3766,N_3280,N_3303);
and U3767 (N_3767,N_3144,N_3320);
nor U3768 (N_3768,N_3360,N_3198);
xor U3769 (N_3769,N_3274,N_3039);
nor U3770 (N_3770,N_3022,N_3470);
nor U3771 (N_3771,N_3076,N_3178);
nand U3772 (N_3772,N_3479,N_3153);
and U3773 (N_3773,N_3168,N_3155);
nor U3774 (N_3774,N_3290,N_3258);
xor U3775 (N_3775,N_3232,N_3121);
nor U3776 (N_3776,N_3341,N_3466);
or U3777 (N_3777,N_3262,N_3145);
xnor U3778 (N_3778,N_3154,N_3438);
xor U3779 (N_3779,N_3143,N_3306);
and U3780 (N_3780,N_3381,N_3111);
or U3781 (N_3781,N_3082,N_3390);
nand U3782 (N_3782,N_3134,N_3380);
or U3783 (N_3783,N_3172,N_3432);
and U3784 (N_3784,N_3149,N_3000);
nor U3785 (N_3785,N_3275,N_3217);
nor U3786 (N_3786,N_3293,N_3329);
nor U3787 (N_3787,N_3421,N_3083);
nor U3788 (N_3788,N_3488,N_3420);
or U3789 (N_3789,N_3448,N_3362);
nand U3790 (N_3790,N_3141,N_3245);
nor U3791 (N_3791,N_3397,N_3030);
xnor U3792 (N_3792,N_3056,N_3149);
nor U3793 (N_3793,N_3253,N_3392);
nor U3794 (N_3794,N_3357,N_3271);
or U3795 (N_3795,N_3477,N_3087);
or U3796 (N_3796,N_3004,N_3464);
nor U3797 (N_3797,N_3287,N_3404);
and U3798 (N_3798,N_3147,N_3015);
and U3799 (N_3799,N_3065,N_3449);
or U3800 (N_3800,N_3223,N_3166);
or U3801 (N_3801,N_3092,N_3332);
nand U3802 (N_3802,N_3356,N_3465);
and U3803 (N_3803,N_3404,N_3471);
nor U3804 (N_3804,N_3367,N_3318);
xor U3805 (N_3805,N_3466,N_3467);
xor U3806 (N_3806,N_3326,N_3051);
nor U3807 (N_3807,N_3119,N_3158);
or U3808 (N_3808,N_3300,N_3301);
and U3809 (N_3809,N_3265,N_3146);
nand U3810 (N_3810,N_3241,N_3467);
or U3811 (N_3811,N_3376,N_3103);
and U3812 (N_3812,N_3207,N_3312);
nor U3813 (N_3813,N_3328,N_3163);
nor U3814 (N_3814,N_3066,N_3422);
or U3815 (N_3815,N_3062,N_3235);
nand U3816 (N_3816,N_3046,N_3316);
nand U3817 (N_3817,N_3384,N_3268);
nand U3818 (N_3818,N_3165,N_3237);
xor U3819 (N_3819,N_3297,N_3412);
and U3820 (N_3820,N_3161,N_3393);
or U3821 (N_3821,N_3433,N_3120);
nor U3822 (N_3822,N_3009,N_3405);
nor U3823 (N_3823,N_3374,N_3011);
or U3824 (N_3824,N_3072,N_3230);
or U3825 (N_3825,N_3178,N_3132);
and U3826 (N_3826,N_3065,N_3003);
and U3827 (N_3827,N_3014,N_3079);
or U3828 (N_3828,N_3377,N_3003);
nor U3829 (N_3829,N_3401,N_3135);
and U3830 (N_3830,N_3338,N_3263);
nor U3831 (N_3831,N_3305,N_3113);
nor U3832 (N_3832,N_3073,N_3387);
nor U3833 (N_3833,N_3397,N_3103);
nor U3834 (N_3834,N_3008,N_3179);
or U3835 (N_3835,N_3201,N_3134);
nand U3836 (N_3836,N_3025,N_3235);
or U3837 (N_3837,N_3003,N_3007);
and U3838 (N_3838,N_3312,N_3251);
and U3839 (N_3839,N_3076,N_3194);
nor U3840 (N_3840,N_3265,N_3466);
and U3841 (N_3841,N_3353,N_3125);
or U3842 (N_3842,N_3460,N_3001);
and U3843 (N_3843,N_3401,N_3075);
and U3844 (N_3844,N_3192,N_3460);
nor U3845 (N_3845,N_3004,N_3068);
and U3846 (N_3846,N_3218,N_3392);
and U3847 (N_3847,N_3030,N_3257);
and U3848 (N_3848,N_3304,N_3477);
xor U3849 (N_3849,N_3196,N_3232);
nor U3850 (N_3850,N_3114,N_3163);
xnor U3851 (N_3851,N_3378,N_3432);
nor U3852 (N_3852,N_3005,N_3499);
xnor U3853 (N_3853,N_3437,N_3337);
or U3854 (N_3854,N_3374,N_3174);
or U3855 (N_3855,N_3321,N_3029);
and U3856 (N_3856,N_3084,N_3359);
or U3857 (N_3857,N_3382,N_3060);
or U3858 (N_3858,N_3454,N_3318);
nor U3859 (N_3859,N_3084,N_3402);
nor U3860 (N_3860,N_3036,N_3089);
xnor U3861 (N_3861,N_3473,N_3325);
nand U3862 (N_3862,N_3287,N_3386);
nand U3863 (N_3863,N_3091,N_3277);
nand U3864 (N_3864,N_3173,N_3095);
and U3865 (N_3865,N_3406,N_3111);
nand U3866 (N_3866,N_3118,N_3248);
and U3867 (N_3867,N_3486,N_3179);
xor U3868 (N_3868,N_3145,N_3235);
and U3869 (N_3869,N_3496,N_3161);
nand U3870 (N_3870,N_3420,N_3472);
or U3871 (N_3871,N_3367,N_3346);
nor U3872 (N_3872,N_3396,N_3336);
or U3873 (N_3873,N_3432,N_3413);
or U3874 (N_3874,N_3190,N_3193);
nor U3875 (N_3875,N_3245,N_3183);
or U3876 (N_3876,N_3282,N_3218);
xor U3877 (N_3877,N_3177,N_3300);
xnor U3878 (N_3878,N_3144,N_3479);
or U3879 (N_3879,N_3367,N_3457);
xor U3880 (N_3880,N_3132,N_3311);
and U3881 (N_3881,N_3031,N_3379);
xnor U3882 (N_3882,N_3093,N_3475);
xor U3883 (N_3883,N_3286,N_3060);
and U3884 (N_3884,N_3417,N_3252);
and U3885 (N_3885,N_3278,N_3371);
or U3886 (N_3886,N_3050,N_3459);
and U3887 (N_3887,N_3096,N_3434);
xor U3888 (N_3888,N_3246,N_3310);
or U3889 (N_3889,N_3327,N_3163);
or U3890 (N_3890,N_3251,N_3293);
nor U3891 (N_3891,N_3452,N_3283);
nor U3892 (N_3892,N_3129,N_3309);
nor U3893 (N_3893,N_3067,N_3225);
nor U3894 (N_3894,N_3383,N_3327);
nand U3895 (N_3895,N_3330,N_3257);
or U3896 (N_3896,N_3038,N_3105);
or U3897 (N_3897,N_3348,N_3285);
and U3898 (N_3898,N_3130,N_3420);
nand U3899 (N_3899,N_3007,N_3275);
nor U3900 (N_3900,N_3498,N_3340);
and U3901 (N_3901,N_3052,N_3452);
nor U3902 (N_3902,N_3003,N_3294);
nand U3903 (N_3903,N_3110,N_3360);
and U3904 (N_3904,N_3064,N_3380);
nor U3905 (N_3905,N_3234,N_3408);
xnor U3906 (N_3906,N_3225,N_3404);
nand U3907 (N_3907,N_3375,N_3228);
and U3908 (N_3908,N_3198,N_3164);
xor U3909 (N_3909,N_3022,N_3105);
and U3910 (N_3910,N_3255,N_3469);
or U3911 (N_3911,N_3498,N_3056);
and U3912 (N_3912,N_3089,N_3073);
or U3913 (N_3913,N_3498,N_3020);
xor U3914 (N_3914,N_3146,N_3389);
nand U3915 (N_3915,N_3447,N_3256);
or U3916 (N_3916,N_3257,N_3055);
or U3917 (N_3917,N_3343,N_3227);
and U3918 (N_3918,N_3427,N_3499);
nand U3919 (N_3919,N_3171,N_3143);
or U3920 (N_3920,N_3478,N_3421);
nor U3921 (N_3921,N_3345,N_3337);
or U3922 (N_3922,N_3272,N_3486);
nand U3923 (N_3923,N_3287,N_3336);
and U3924 (N_3924,N_3458,N_3221);
xnor U3925 (N_3925,N_3174,N_3285);
and U3926 (N_3926,N_3354,N_3037);
or U3927 (N_3927,N_3473,N_3421);
or U3928 (N_3928,N_3461,N_3478);
or U3929 (N_3929,N_3371,N_3243);
and U3930 (N_3930,N_3222,N_3083);
xnor U3931 (N_3931,N_3256,N_3235);
or U3932 (N_3932,N_3334,N_3456);
and U3933 (N_3933,N_3388,N_3425);
nand U3934 (N_3934,N_3424,N_3263);
or U3935 (N_3935,N_3369,N_3427);
nand U3936 (N_3936,N_3409,N_3313);
and U3937 (N_3937,N_3220,N_3436);
xnor U3938 (N_3938,N_3350,N_3490);
or U3939 (N_3939,N_3304,N_3004);
nor U3940 (N_3940,N_3131,N_3248);
nand U3941 (N_3941,N_3180,N_3309);
nor U3942 (N_3942,N_3359,N_3330);
nand U3943 (N_3943,N_3129,N_3431);
and U3944 (N_3944,N_3465,N_3303);
or U3945 (N_3945,N_3239,N_3307);
and U3946 (N_3946,N_3070,N_3128);
xnor U3947 (N_3947,N_3425,N_3027);
and U3948 (N_3948,N_3229,N_3147);
nand U3949 (N_3949,N_3372,N_3331);
or U3950 (N_3950,N_3328,N_3282);
and U3951 (N_3951,N_3024,N_3483);
and U3952 (N_3952,N_3021,N_3436);
and U3953 (N_3953,N_3356,N_3404);
nor U3954 (N_3954,N_3346,N_3489);
nand U3955 (N_3955,N_3130,N_3393);
nand U3956 (N_3956,N_3218,N_3113);
or U3957 (N_3957,N_3123,N_3046);
or U3958 (N_3958,N_3156,N_3061);
and U3959 (N_3959,N_3251,N_3280);
or U3960 (N_3960,N_3058,N_3390);
or U3961 (N_3961,N_3086,N_3222);
or U3962 (N_3962,N_3440,N_3354);
nand U3963 (N_3963,N_3246,N_3004);
nand U3964 (N_3964,N_3049,N_3014);
nand U3965 (N_3965,N_3265,N_3450);
nor U3966 (N_3966,N_3282,N_3274);
and U3967 (N_3967,N_3328,N_3122);
or U3968 (N_3968,N_3287,N_3135);
xnor U3969 (N_3969,N_3454,N_3021);
or U3970 (N_3970,N_3230,N_3311);
nand U3971 (N_3971,N_3067,N_3481);
and U3972 (N_3972,N_3431,N_3022);
and U3973 (N_3973,N_3330,N_3278);
or U3974 (N_3974,N_3358,N_3497);
and U3975 (N_3975,N_3012,N_3378);
or U3976 (N_3976,N_3163,N_3185);
nand U3977 (N_3977,N_3245,N_3417);
and U3978 (N_3978,N_3149,N_3052);
nand U3979 (N_3979,N_3410,N_3005);
nor U3980 (N_3980,N_3084,N_3225);
nor U3981 (N_3981,N_3499,N_3146);
nor U3982 (N_3982,N_3488,N_3423);
nand U3983 (N_3983,N_3170,N_3375);
nand U3984 (N_3984,N_3264,N_3225);
or U3985 (N_3985,N_3340,N_3439);
nor U3986 (N_3986,N_3429,N_3022);
nand U3987 (N_3987,N_3023,N_3273);
nor U3988 (N_3988,N_3417,N_3366);
nand U3989 (N_3989,N_3452,N_3367);
nor U3990 (N_3990,N_3492,N_3261);
nand U3991 (N_3991,N_3422,N_3197);
and U3992 (N_3992,N_3082,N_3040);
nand U3993 (N_3993,N_3185,N_3195);
nand U3994 (N_3994,N_3301,N_3188);
and U3995 (N_3995,N_3250,N_3149);
nand U3996 (N_3996,N_3316,N_3221);
and U3997 (N_3997,N_3458,N_3081);
nor U3998 (N_3998,N_3142,N_3438);
or U3999 (N_3999,N_3297,N_3462);
xor U4000 (N_4000,N_3505,N_3644);
and U4001 (N_4001,N_3612,N_3533);
nor U4002 (N_4002,N_3960,N_3677);
nor U4003 (N_4003,N_3899,N_3849);
and U4004 (N_4004,N_3866,N_3536);
or U4005 (N_4005,N_3743,N_3572);
nor U4006 (N_4006,N_3887,N_3624);
nand U4007 (N_4007,N_3750,N_3812);
or U4008 (N_4008,N_3756,N_3645);
or U4009 (N_4009,N_3813,N_3882);
and U4010 (N_4010,N_3664,N_3651);
nand U4011 (N_4011,N_3772,N_3800);
or U4012 (N_4012,N_3716,N_3563);
and U4013 (N_4013,N_3749,N_3891);
and U4014 (N_4014,N_3604,N_3809);
and U4015 (N_4015,N_3641,N_3917);
and U4016 (N_4016,N_3930,N_3957);
and U4017 (N_4017,N_3778,N_3981);
nor U4018 (N_4018,N_3737,N_3646);
nor U4019 (N_4019,N_3504,N_3995);
nor U4020 (N_4020,N_3875,N_3517);
or U4021 (N_4021,N_3864,N_3652);
nand U4022 (N_4022,N_3782,N_3876);
nand U4023 (N_4023,N_3923,N_3924);
or U4024 (N_4024,N_3835,N_3852);
nor U4025 (N_4025,N_3633,N_3661);
xor U4026 (N_4026,N_3821,N_3710);
and U4027 (N_4027,N_3636,N_3647);
and U4028 (N_4028,N_3690,N_3593);
nor U4029 (N_4029,N_3993,N_3968);
nand U4030 (N_4030,N_3831,N_3523);
nor U4031 (N_4031,N_3587,N_3983);
or U4032 (N_4032,N_3600,N_3739);
nand U4033 (N_4033,N_3599,N_3579);
nand U4034 (N_4034,N_3574,N_3794);
nand U4035 (N_4035,N_3860,N_3971);
or U4036 (N_4036,N_3807,N_3975);
nor U4037 (N_4037,N_3718,N_3655);
xnor U4038 (N_4038,N_3781,N_3817);
nand U4039 (N_4039,N_3705,N_3642);
nor U4040 (N_4040,N_3793,N_3902);
and U4041 (N_4041,N_3659,N_3557);
and U4042 (N_4042,N_3826,N_3613);
nand U4043 (N_4043,N_3699,N_3906);
or U4044 (N_4044,N_3823,N_3900);
nand U4045 (N_4045,N_3685,N_3639);
nor U4046 (N_4046,N_3627,N_3700);
nand U4047 (N_4047,N_3577,N_3903);
or U4048 (N_4048,N_3684,N_3952);
and U4049 (N_4049,N_3565,N_3569);
and U4050 (N_4050,N_3571,N_3506);
or U4051 (N_4051,N_3632,N_3741);
xnor U4052 (N_4052,N_3789,N_3996);
nand U4053 (N_4053,N_3561,N_3970);
nor U4054 (N_4054,N_3736,N_3539);
or U4055 (N_4055,N_3522,N_3942);
nor U4056 (N_4056,N_3583,N_3769);
nand U4057 (N_4057,N_3724,N_3631);
and U4058 (N_4058,N_3745,N_3703);
nand U4059 (N_4059,N_3621,N_3767);
nand U4060 (N_4060,N_3878,N_3886);
or U4061 (N_4061,N_3735,N_3824);
nor U4062 (N_4062,N_3846,N_3618);
xnor U4063 (N_4063,N_3681,N_3568);
nor U4064 (N_4064,N_3722,N_3582);
nor U4065 (N_4065,N_3626,N_3799);
or U4066 (N_4066,N_3758,N_3606);
and U4067 (N_4067,N_3529,N_3992);
and U4068 (N_4068,N_3680,N_3501);
nand U4069 (N_4069,N_3775,N_3802);
nand U4070 (N_4070,N_3939,N_3988);
and U4071 (N_4071,N_3963,N_3698);
and U4072 (N_4072,N_3512,N_3546);
or U4073 (N_4073,N_3801,N_3511);
and U4074 (N_4074,N_3721,N_3667);
and U4075 (N_4075,N_3711,N_3640);
nand U4076 (N_4076,N_3602,N_3714);
nor U4077 (N_4077,N_3715,N_3603);
and U4078 (N_4078,N_3972,N_3895);
nor U4079 (N_4079,N_3610,N_3933);
or U4080 (N_4080,N_3945,N_3670);
nor U4081 (N_4081,N_3570,N_3842);
nor U4082 (N_4082,N_3986,N_3682);
nor U4083 (N_4083,N_3768,N_3978);
and U4084 (N_4084,N_3907,N_3779);
nor U4085 (N_4085,N_3752,N_3958);
nor U4086 (N_4086,N_3607,N_3982);
xor U4087 (N_4087,N_3845,N_3701);
or U4088 (N_4088,N_3910,N_3798);
nand U4089 (N_4089,N_3947,N_3530);
nor U4090 (N_4090,N_3921,N_3719);
or U4091 (N_4091,N_3863,N_3908);
nand U4092 (N_4092,N_3591,N_3580);
nor U4093 (N_4093,N_3815,N_3709);
nand U4094 (N_4094,N_3774,N_3980);
or U4095 (N_4095,N_3893,N_3785);
nor U4096 (N_4096,N_3656,N_3814);
nand U4097 (N_4097,N_3611,N_3560);
and U4098 (N_4098,N_3760,N_3989);
and U4099 (N_4099,N_3796,N_3726);
and U4100 (N_4100,N_3829,N_3609);
or U4101 (N_4101,N_3788,N_3585);
nor U4102 (N_4102,N_3623,N_3643);
xnor U4103 (N_4103,N_3990,N_3567);
nor U4104 (N_4104,N_3833,N_3732);
nand U4105 (N_4105,N_3562,N_3855);
nand U4106 (N_4106,N_3578,N_3552);
or U4107 (N_4107,N_3649,N_3666);
nor U4108 (N_4108,N_3940,N_3538);
nand U4109 (N_4109,N_3524,N_3730);
xnor U4110 (N_4110,N_3733,N_3912);
xor U4111 (N_4111,N_3590,N_3843);
nor U4112 (N_4112,N_3566,N_3979);
or U4113 (N_4113,N_3507,N_3897);
nor U4114 (N_4114,N_3548,N_3707);
and U4115 (N_4115,N_3559,N_3994);
nand U4116 (N_4116,N_3728,N_3783);
nor U4117 (N_4117,N_3770,N_3601);
and U4118 (N_4118,N_3965,N_3911);
nand U4119 (N_4119,N_3625,N_3803);
nor U4120 (N_4120,N_3605,N_3747);
and U4121 (N_4121,N_3985,N_3766);
or U4122 (N_4122,N_3915,N_3731);
and U4123 (N_4123,N_3776,N_3959);
or U4124 (N_4124,N_3576,N_3927);
or U4125 (N_4125,N_3874,N_3628);
and U4126 (N_4126,N_3790,N_3634);
xnor U4127 (N_4127,N_3532,N_3780);
or U4128 (N_4128,N_3695,N_3820);
or U4129 (N_4129,N_3848,N_3870);
nand U4130 (N_4130,N_3859,N_3521);
nand U4131 (N_4131,N_3660,N_3668);
nand U4132 (N_4132,N_3811,N_3616);
nor U4133 (N_4133,N_3762,N_3808);
nor U4134 (N_4134,N_3748,N_3810);
or U4135 (N_4135,N_3961,N_3503);
nor U4136 (N_4136,N_3854,N_3950);
nor U4137 (N_4137,N_3754,N_3637);
and U4138 (N_4138,N_3653,N_3595);
or U4139 (N_4139,N_3828,N_3551);
nor U4140 (N_4140,N_3687,N_3549);
and U4141 (N_4141,N_3584,N_3837);
or U4142 (N_4142,N_3884,N_3851);
nand U4143 (N_4143,N_3956,N_3784);
nand U4144 (N_4144,N_3615,N_3658);
nand U4145 (N_4145,N_3706,N_3871);
nand U4146 (N_4146,N_3806,N_3954);
and U4147 (N_4147,N_3597,N_3555);
nand U4148 (N_4148,N_3725,N_3712);
nand U4149 (N_4149,N_3937,N_3541);
or U4150 (N_4150,N_3825,N_3525);
nor U4151 (N_4151,N_3713,N_3973);
nand U4152 (N_4152,N_3941,N_3573);
and U4153 (N_4153,N_3753,N_3929);
and U4154 (N_4154,N_3827,N_3673);
nand U4155 (N_4155,N_3751,N_3764);
or U4156 (N_4156,N_3918,N_3598);
nand U4157 (N_4157,N_3868,N_3676);
or U4158 (N_4158,N_3925,N_3763);
nor U4159 (N_4159,N_3894,N_3922);
nand U4160 (N_4160,N_3861,N_3969);
nand U4161 (N_4161,N_3999,N_3696);
xnor U4162 (N_4162,N_3596,N_3535);
or U4163 (N_4163,N_3967,N_3746);
or U4164 (N_4164,N_3856,N_3686);
and U4165 (N_4165,N_3890,N_3558);
xor U4166 (N_4166,N_3987,N_3926);
nand U4167 (N_4167,N_3689,N_3594);
nand U4168 (N_4168,N_3509,N_3759);
nor U4169 (N_4169,N_3830,N_3883);
and U4170 (N_4170,N_3669,N_3932);
or U4171 (N_4171,N_3919,N_3955);
or U4172 (N_4172,N_3547,N_3635);
nor U4173 (N_4173,N_3966,N_3510);
and U4174 (N_4174,N_3951,N_3905);
or U4175 (N_4175,N_3672,N_3519);
nand U4176 (N_4176,N_3836,N_3832);
or U4177 (N_4177,N_3998,N_3885);
nand U4178 (N_4178,N_3528,N_3976);
or U4179 (N_4179,N_3761,N_3526);
nand U4180 (N_4180,N_3822,N_3543);
nor U4181 (N_4181,N_3888,N_3777);
nand U4182 (N_4182,N_3857,N_3755);
nor U4183 (N_4183,N_3935,N_3841);
nand U4184 (N_4184,N_3928,N_3791);
nand U4185 (N_4185,N_3675,N_3554);
nand U4186 (N_4186,N_3542,N_3638);
or U4187 (N_4187,N_3729,N_3974);
and U4188 (N_4188,N_3513,N_3630);
and U4189 (N_4189,N_3520,N_3662);
xor U4190 (N_4190,N_3697,N_3740);
and U4191 (N_4191,N_3962,N_3514);
and U4192 (N_4192,N_3744,N_3792);
nor U4193 (N_4193,N_3946,N_3614);
nor U4194 (N_4194,N_3518,N_3867);
nor U4195 (N_4195,N_3723,N_3914);
and U4196 (N_4196,N_3704,N_3622);
nor U4197 (N_4197,N_3742,N_3818);
nor U4198 (N_4198,N_3620,N_3869);
nand U4199 (N_4199,N_3515,N_3692);
and U4200 (N_4200,N_3944,N_3765);
or U4201 (N_4201,N_3516,N_3581);
nand U4202 (N_4202,N_3589,N_3805);
nand U4203 (N_4203,N_3839,N_3502);
nand U4204 (N_4204,N_3920,N_3537);
or U4205 (N_4205,N_3702,N_3545);
or U4206 (N_4206,N_3657,N_3949);
and U4207 (N_4207,N_3916,N_3691);
nand U4208 (N_4208,N_3880,N_3889);
or U4209 (N_4209,N_3934,N_3877);
nand U4210 (N_4210,N_3720,N_3938);
nand U4211 (N_4211,N_3683,N_3865);
xnor U4212 (N_4212,N_3564,N_3738);
nand U4213 (N_4213,N_3892,N_3953);
xor U4214 (N_4214,N_3586,N_3575);
or U4215 (N_4215,N_3617,N_3619);
and U4216 (N_4216,N_3786,N_3663);
nor U4217 (N_4217,N_3654,N_3534);
nor U4218 (N_4218,N_3508,N_3862);
nand U4219 (N_4219,N_3688,N_3679);
nand U4220 (N_4220,N_3819,N_3879);
nand U4221 (N_4221,N_3853,N_3629);
nor U4222 (N_4222,N_3881,N_3909);
xor U4223 (N_4223,N_3674,N_3838);
nor U4224 (N_4224,N_3795,N_3977);
or U4225 (N_4225,N_3734,N_3991);
nor U4226 (N_4226,N_3872,N_3904);
and U4227 (N_4227,N_3500,N_3678);
or U4228 (N_4228,N_3847,N_3901);
nor U4229 (N_4229,N_3665,N_3694);
or U4230 (N_4230,N_3840,N_3693);
nor U4231 (N_4231,N_3913,N_3943);
nand U4232 (N_4232,N_3771,N_3588);
nand U4233 (N_4233,N_3717,N_3787);
and U4234 (N_4234,N_3592,N_3708);
and U4235 (N_4235,N_3816,N_3648);
or U4236 (N_4236,N_3556,N_3553);
nor U4237 (N_4237,N_3931,N_3773);
xor U4238 (N_4238,N_3858,N_3540);
nor U4239 (N_4239,N_3727,N_3550);
and U4240 (N_4240,N_3850,N_3898);
or U4241 (N_4241,N_3608,N_3757);
or U4242 (N_4242,N_3873,N_3650);
and U4243 (N_4243,N_3671,N_3797);
xor U4244 (N_4244,N_3804,N_3936);
nand U4245 (N_4245,N_3948,N_3544);
nor U4246 (N_4246,N_3527,N_3984);
nand U4247 (N_4247,N_3844,N_3964);
and U4248 (N_4248,N_3896,N_3834);
or U4249 (N_4249,N_3531,N_3997);
nand U4250 (N_4250,N_3865,N_3720);
nor U4251 (N_4251,N_3862,N_3524);
xnor U4252 (N_4252,N_3721,N_3982);
or U4253 (N_4253,N_3766,N_3699);
and U4254 (N_4254,N_3920,N_3908);
nor U4255 (N_4255,N_3673,N_3799);
or U4256 (N_4256,N_3524,N_3654);
or U4257 (N_4257,N_3821,N_3781);
nor U4258 (N_4258,N_3538,N_3963);
or U4259 (N_4259,N_3725,N_3673);
or U4260 (N_4260,N_3766,N_3576);
nor U4261 (N_4261,N_3951,N_3796);
nand U4262 (N_4262,N_3832,N_3999);
nor U4263 (N_4263,N_3700,N_3997);
or U4264 (N_4264,N_3853,N_3680);
and U4265 (N_4265,N_3854,N_3569);
and U4266 (N_4266,N_3740,N_3578);
and U4267 (N_4267,N_3561,N_3741);
or U4268 (N_4268,N_3800,N_3766);
nand U4269 (N_4269,N_3533,N_3548);
or U4270 (N_4270,N_3867,N_3514);
xnor U4271 (N_4271,N_3605,N_3709);
or U4272 (N_4272,N_3662,N_3764);
and U4273 (N_4273,N_3948,N_3947);
nor U4274 (N_4274,N_3778,N_3539);
nor U4275 (N_4275,N_3728,N_3761);
and U4276 (N_4276,N_3775,N_3857);
or U4277 (N_4277,N_3904,N_3945);
or U4278 (N_4278,N_3574,N_3528);
or U4279 (N_4279,N_3684,N_3959);
or U4280 (N_4280,N_3694,N_3659);
nand U4281 (N_4281,N_3562,N_3739);
or U4282 (N_4282,N_3857,N_3885);
nand U4283 (N_4283,N_3721,N_3733);
nor U4284 (N_4284,N_3762,N_3927);
nand U4285 (N_4285,N_3918,N_3612);
xnor U4286 (N_4286,N_3760,N_3796);
xor U4287 (N_4287,N_3648,N_3864);
or U4288 (N_4288,N_3934,N_3736);
or U4289 (N_4289,N_3843,N_3823);
nand U4290 (N_4290,N_3984,N_3760);
or U4291 (N_4291,N_3924,N_3993);
xor U4292 (N_4292,N_3749,N_3825);
nand U4293 (N_4293,N_3979,N_3832);
nor U4294 (N_4294,N_3662,N_3700);
and U4295 (N_4295,N_3686,N_3949);
nand U4296 (N_4296,N_3643,N_3736);
nor U4297 (N_4297,N_3776,N_3833);
or U4298 (N_4298,N_3580,N_3930);
nor U4299 (N_4299,N_3554,N_3528);
or U4300 (N_4300,N_3647,N_3645);
or U4301 (N_4301,N_3510,N_3970);
nand U4302 (N_4302,N_3877,N_3952);
nand U4303 (N_4303,N_3830,N_3744);
xor U4304 (N_4304,N_3800,N_3951);
and U4305 (N_4305,N_3585,N_3795);
nand U4306 (N_4306,N_3761,N_3859);
nor U4307 (N_4307,N_3863,N_3675);
and U4308 (N_4308,N_3949,N_3633);
and U4309 (N_4309,N_3544,N_3695);
or U4310 (N_4310,N_3590,N_3508);
or U4311 (N_4311,N_3640,N_3503);
nand U4312 (N_4312,N_3662,N_3725);
nor U4313 (N_4313,N_3668,N_3858);
or U4314 (N_4314,N_3853,N_3601);
nand U4315 (N_4315,N_3942,N_3974);
xnor U4316 (N_4316,N_3684,N_3978);
or U4317 (N_4317,N_3816,N_3825);
nor U4318 (N_4318,N_3912,N_3864);
or U4319 (N_4319,N_3868,N_3561);
nand U4320 (N_4320,N_3823,N_3905);
nor U4321 (N_4321,N_3629,N_3589);
or U4322 (N_4322,N_3591,N_3854);
nor U4323 (N_4323,N_3716,N_3970);
or U4324 (N_4324,N_3535,N_3785);
and U4325 (N_4325,N_3652,N_3622);
nand U4326 (N_4326,N_3605,N_3919);
and U4327 (N_4327,N_3821,N_3703);
nor U4328 (N_4328,N_3736,N_3593);
and U4329 (N_4329,N_3697,N_3943);
xnor U4330 (N_4330,N_3698,N_3674);
or U4331 (N_4331,N_3661,N_3968);
or U4332 (N_4332,N_3500,N_3507);
and U4333 (N_4333,N_3572,N_3584);
nand U4334 (N_4334,N_3842,N_3515);
and U4335 (N_4335,N_3629,N_3715);
and U4336 (N_4336,N_3852,N_3798);
or U4337 (N_4337,N_3762,N_3783);
or U4338 (N_4338,N_3710,N_3827);
or U4339 (N_4339,N_3593,N_3890);
or U4340 (N_4340,N_3520,N_3599);
nor U4341 (N_4341,N_3672,N_3942);
and U4342 (N_4342,N_3636,N_3828);
nor U4343 (N_4343,N_3838,N_3810);
nand U4344 (N_4344,N_3881,N_3525);
nand U4345 (N_4345,N_3510,N_3723);
nand U4346 (N_4346,N_3564,N_3799);
nand U4347 (N_4347,N_3817,N_3893);
nor U4348 (N_4348,N_3882,N_3830);
nor U4349 (N_4349,N_3781,N_3770);
and U4350 (N_4350,N_3864,N_3878);
and U4351 (N_4351,N_3838,N_3966);
nor U4352 (N_4352,N_3810,N_3517);
or U4353 (N_4353,N_3752,N_3516);
nand U4354 (N_4354,N_3930,N_3533);
nand U4355 (N_4355,N_3646,N_3949);
nand U4356 (N_4356,N_3557,N_3723);
and U4357 (N_4357,N_3670,N_3543);
or U4358 (N_4358,N_3543,N_3802);
and U4359 (N_4359,N_3924,N_3508);
xnor U4360 (N_4360,N_3664,N_3848);
or U4361 (N_4361,N_3947,N_3847);
nor U4362 (N_4362,N_3607,N_3610);
xor U4363 (N_4363,N_3708,N_3711);
nand U4364 (N_4364,N_3741,N_3885);
or U4365 (N_4365,N_3577,N_3632);
and U4366 (N_4366,N_3723,N_3580);
nand U4367 (N_4367,N_3893,N_3951);
nor U4368 (N_4368,N_3732,N_3584);
or U4369 (N_4369,N_3731,N_3761);
nor U4370 (N_4370,N_3669,N_3686);
and U4371 (N_4371,N_3597,N_3819);
nor U4372 (N_4372,N_3705,N_3854);
and U4373 (N_4373,N_3759,N_3565);
nor U4374 (N_4374,N_3540,N_3965);
nand U4375 (N_4375,N_3658,N_3512);
nor U4376 (N_4376,N_3613,N_3959);
nor U4377 (N_4377,N_3646,N_3597);
or U4378 (N_4378,N_3599,N_3751);
or U4379 (N_4379,N_3713,N_3789);
or U4380 (N_4380,N_3513,N_3985);
or U4381 (N_4381,N_3630,N_3949);
nor U4382 (N_4382,N_3643,N_3831);
nor U4383 (N_4383,N_3831,N_3666);
nand U4384 (N_4384,N_3590,N_3666);
nor U4385 (N_4385,N_3727,N_3715);
nor U4386 (N_4386,N_3599,N_3902);
nand U4387 (N_4387,N_3512,N_3771);
or U4388 (N_4388,N_3969,N_3818);
nor U4389 (N_4389,N_3886,N_3978);
or U4390 (N_4390,N_3926,N_3779);
and U4391 (N_4391,N_3521,N_3867);
nand U4392 (N_4392,N_3642,N_3841);
nand U4393 (N_4393,N_3619,N_3849);
or U4394 (N_4394,N_3623,N_3572);
nand U4395 (N_4395,N_3943,N_3832);
or U4396 (N_4396,N_3703,N_3557);
nor U4397 (N_4397,N_3739,N_3628);
or U4398 (N_4398,N_3724,N_3553);
nor U4399 (N_4399,N_3635,N_3941);
xor U4400 (N_4400,N_3962,N_3999);
nor U4401 (N_4401,N_3972,N_3906);
and U4402 (N_4402,N_3750,N_3712);
xnor U4403 (N_4403,N_3991,N_3530);
and U4404 (N_4404,N_3504,N_3740);
and U4405 (N_4405,N_3837,N_3742);
nor U4406 (N_4406,N_3766,N_3880);
nand U4407 (N_4407,N_3565,N_3600);
or U4408 (N_4408,N_3918,N_3992);
nor U4409 (N_4409,N_3880,N_3854);
xnor U4410 (N_4410,N_3966,N_3822);
nor U4411 (N_4411,N_3783,N_3575);
or U4412 (N_4412,N_3644,N_3655);
and U4413 (N_4413,N_3520,N_3740);
and U4414 (N_4414,N_3752,N_3676);
xor U4415 (N_4415,N_3983,N_3762);
and U4416 (N_4416,N_3602,N_3859);
or U4417 (N_4417,N_3924,N_3526);
and U4418 (N_4418,N_3732,N_3748);
or U4419 (N_4419,N_3670,N_3725);
or U4420 (N_4420,N_3861,N_3560);
or U4421 (N_4421,N_3924,N_3603);
nor U4422 (N_4422,N_3507,N_3601);
nand U4423 (N_4423,N_3581,N_3662);
xnor U4424 (N_4424,N_3730,N_3670);
or U4425 (N_4425,N_3717,N_3601);
nand U4426 (N_4426,N_3826,N_3641);
or U4427 (N_4427,N_3791,N_3930);
or U4428 (N_4428,N_3980,N_3609);
xnor U4429 (N_4429,N_3910,N_3822);
nor U4430 (N_4430,N_3797,N_3835);
and U4431 (N_4431,N_3552,N_3820);
nand U4432 (N_4432,N_3818,N_3962);
xor U4433 (N_4433,N_3519,N_3847);
and U4434 (N_4434,N_3760,N_3699);
and U4435 (N_4435,N_3822,N_3668);
nand U4436 (N_4436,N_3954,N_3559);
or U4437 (N_4437,N_3765,N_3998);
xnor U4438 (N_4438,N_3553,N_3624);
nand U4439 (N_4439,N_3876,N_3912);
nor U4440 (N_4440,N_3759,N_3545);
nand U4441 (N_4441,N_3653,N_3611);
and U4442 (N_4442,N_3626,N_3555);
nor U4443 (N_4443,N_3586,N_3576);
nand U4444 (N_4444,N_3790,N_3982);
or U4445 (N_4445,N_3697,N_3623);
nand U4446 (N_4446,N_3695,N_3801);
and U4447 (N_4447,N_3654,N_3908);
nor U4448 (N_4448,N_3902,N_3910);
nand U4449 (N_4449,N_3602,N_3932);
or U4450 (N_4450,N_3839,N_3516);
nand U4451 (N_4451,N_3616,N_3540);
nor U4452 (N_4452,N_3528,N_3529);
nand U4453 (N_4453,N_3679,N_3887);
or U4454 (N_4454,N_3815,N_3884);
nor U4455 (N_4455,N_3888,N_3641);
and U4456 (N_4456,N_3728,N_3678);
nor U4457 (N_4457,N_3867,N_3968);
and U4458 (N_4458,N_3690,N_3615);
or U4459 (N_4459,N_3660,N_3854);
xor U4460 (N_4460,N_3599,N_3590);
and U4461 (N_4461,N_3750,N_3931);
and U4462 (N_4462,N_3740,N_3736);
nand U4463 (N_4463,N_3955,N_3786);
or U4464 (N_4464,N_3803,N_3921);
nand U4465 (N_4465,N_3965,N_3578);
xnor U4466 (N_4466,N_3831,N_3603);
and U4467 (N_4467,N_3917,N_3852);
nor U4468 (N_4468,N_3882,N_3966);
nand U4469 (N_4469,N_3778,N_3692);
or U4470 (N_4470,N_3663,N_3941);
nor U4471 (N_4471,N_3875,N_3942);
and U4472 (N_4472,N_3758,N_3872);
nor U4473 (N_4473,N_3524,N_3863);
nand U4474 (N_4474,N_3685,N_3673);
or U4475 (N_4475,N_3766,N_3879);
xnor U4476 (N_4476,N_3818,N_3799);
and U4477 (N_4477,N_3591,N_3622);
nand U4478 (N_4478,N_3617,N_3634);
nor U4479 (N_4479,N_3877,N_3896);
and U4480 (N_4480,N_3650,N_3976);
nand U4481 (N_4481,N_3935,N_3502);
nand U4482 (N_4482,N_3686,N_3788);
nor U4483 (N_4483,N_3640,N_3517);
nor U4484 (N_4484,N_3826,N_3567);
nand U4485 (N_4485,N_3696,N_3631);
or U4486 (N_4486,N_3989,N_3833);
or U4487 (N_4487,N_3528,N_3726);
or U4488 (N_4488,N_3600,N_3932);
nor U4489 (N_4489,N_3982,N_3639);
or U4490 (N_4490,N_3532,N_3944);
and U4491 (N_4491,N_3806,N_3768);
and U4492 (N_4492,N_3514,N_3955);
nor U4493 (N_4493,N_3742,N_3934);
or U4494 (N_4494,N_3944,N_3801);
and U4495 (N_4495,N_3755,N_3571);
xnor U4496 (N_4496,N_3566,N_3859);
or U4497 (N_4497,N_3623,N_3515);
and U4498 (N_4498,N_3636,N_3625);
and U4499 (N_4499,N_3974,N_3583);
nor U4500 (N_4500,N_4087,N_4370);
or U4501 (N_4501,N_4310,N_4332);
nor U4502 (N_4502,N_4004,N_4009);
or U4503 (N_4503,N_4448,N_4053);
nor U4504 (N_4504,N_4207,N_4463);
or U4505 (N_4505,N_4286,N_4269);
or U4506 (N_4506,N_4368,N_4294);
or U4507 (N_4507,N_4001,N_4139);
or U4508 (N_4508,N_4261,N_4265);
nor U4509 (N_4509,N_4033,N_4318);
nand U4510 (N_4510,N_4467,N_4345);
or U4511 (N_4511,N_4330,N_4169);
nor U4512 (N_4512,N_4088,N_4275);
and U4513 (N_4513,N_4222,N_4324);
nor U4514 (N_4514,N_4414,N_4117);
and U4515 (N_4515,N_4451,N_4406);
nor U4516 (N_4516,N_4454,N_4431);
xor U4517 (N_4517,N_4236,N_4135);
nand U4518 (N_4518,N_4389,N_4060);
and U4519 (N_4519,N_4335,N_4128);
or U4520 (N_4520,N_4258,N_4072);
nand U4521 (N_4521,N_4348,N_4358);
nor U4522 (N_4522,N_4405,N_4290);
or U4523 (N_4523,N_4172,N_4472);
xnor U4524 (N_4524,N_4442,N_4006);
nand U4525 (N_4525,N_4347,N_4134);
and U4526 (N_4526,N_4400,N_4056);
nand U4527 (N_4527,N_4132,N_4148);
or U4528 (N_4528,N_4364,N_4447);
or U4529 (N_4529,N_4082,N_4440);
xor U4530 (N_4530,N_4080,N_4177);
nand U4531 (N_4531,N_4255,N_4031);
nor U4532 (N_4532,N_4316,N_4349);
and U4533 (N_4533,N_4107,N_4126);
or U4534 (N_4534,N_4159,N_4297);
nand U4535 (N_4535,N_4045,N_4312);
nand U4536 (N_4536,N_4016,N_4422);
nor U4537 (N_4537,N_4254,N_4231);
and U4538 (N_4538,N_4064,N_4250);
nor U4539 (N_4539,N_4057,N_4011);
or U4540 (N_4540,N_4327,N_4227);
or U4541 (N_4541,N_4449,N_4311);
nand U4542 (N_4542,N_4339,N_4419);
or U4543 (N_4543,N_4380,N_4163);
nor U4544 (N_4544,N_4421,N_4167);
or U4545 (N_4545,N_4424,N_4302);
and U4546 (N_4546,N_4019,N_4040);
nor U4547 (N_4547,N_4284,N_4085);
and U4548 (N_4548,N_4136,N_4003);
nor U4549 (N_4549,N_4032,N_4241);
or U4550 (N_4550,N_4027,N_4049);
nor U4551 (N_4551,N_4300,N_4109);
xor U4552 (N_4552,N_4147,N_4257);
or U4553 (N_4553,N_4476,N_4051);
nor U4554 (N_4554,N_4252,N_4341);
nor U4555 (N_4555,N_4041,N_4202);
nand U4556 (N_4556,N_4281,N_4029);
or U4557 (N_4557,N_4112,N_4156);
and U4558 (N_4558,N_4306,N_4133);
nand U4559 (N_4559,N_4480,N_4425);
or U4560 (N_4560,N_4168,N_4403);
and U4561 (N_4561,N_4268,N_4193);
and U4562 (N_4562,N_4489,N_4307);
nand U4563 (N_4563,N_4313,N_4234);
and U4564 (N_4564,N_4475,N_4283);
nand U4565 (N_4565,N_4468,N_4428);
or U4566 (N_4566,N_4038,N_4015);
or U4567 (N_4567,N_4378,N_4247);
and U4568 (N_4568,N_4384,N_4012);
and U4569 (N_4569,N_4140,N_4355);
xor U4570 (N_4570,N_4196,N_4399);
nor U4571 (N_4571,N_4151,N_4209);
and U4572 (N_4572,N_4430,N_4484);
nand U4573 (N_4573,N_4195,N_4095);
and U4574 (N_4574,N_4483,N_4150);
or U4575 (N_4575,N_4093,N_4065);
nor U4576 (N_4576,N_4402,N_4305);
and U4577 (N_4577,N_4259,N_4342);
xnor U4578 (N_4578,N_4477,N_4433);
nor U4579 (N_4579,N_4071,N_4097);
and U4580 (N_4580,N_4044,N_4473);
xnor U4581 (N_4581,N_4081,N_4069);
or U4582 (N_4582,N_4233,N_4469);
nor U4583 (N_4583,N_4392,N_4223);
and U4584 (N_4584,N_4287,N_4180);
xnor U4585 (N_4585,N_4170,N_4372);
and U4586 (N_4586,N_4164,N_4459);
nand U4587 (N_4587,N_4017,N_4420);
xor U4588 (N_4588,N_4130,N_4187);
nand U4589 (N_4589,N_4343,N_4217);
and U4590 (N_4590,N_4353,N_4350);
nand U4591 (N_4591,N_4220,N_4018);
or U4592 (N_4592,N_4116,N_4188);
xor U4593 (N_4593,N_4435,N_4121);
or U4594 (N_4594,N_4374,N_4411);
and U4595 (N_4595,N_4418,N_4314);
and U4596 (N_4596,N_4340,N_4062);
and U4597 (N_4597,N_4212,N_4118);
and U4598 (N_4598,N_4205,N_4079);
nor U4599 (N_4599,N_4386,N_4367);
nand U4600 (N_4600,N_4333,N_4216);
nor U4601 (N_4601,N_4161,N_4211);
nor U4602 (N_4602,N_4299,N_4194);
or U4603 (N_4603,N_4393,N_4007);
and U4604 (N_4604,N_4200,N_4113);
nor U4605 (N_4605,N_4185,N_4096);
or U4606 (N_4606,N_4086,N_4471);
nand U4607 (N_4607,N_4171,N_4490);
xnor U4608 (N_4608,N_4068,N_4478);
nand U4609 (N_4609,N_4103,N_4398);
and U4610 (N_4610,N_4091,N_4249);
or U4611 (N_4611,N_4083,N_4423);
and U4612 (N_4612,N_4042,N_4179);
or U4613 (N_4613,N_4174,N_4479);
nor U4614 (N_4614,N_4201,N_4025);
nand U4615 (N_4615,N_4266,N_4120);
xor U4616 (N_4616,N_4090,N_4050);
nand U4617 (N_4617,N_4465,N_4142);
or U4618 (N_4618,N_4323,N_4391);
and U4619 (N_4619,N_4183,N_4395);
and U4620 (N_4620,N_4052,N_4273);
and U4621 (N_4621,N_4450,N_4125);
nand U4622 (N_4622,N_4496,N_4158);
nor U4623 (N_4623,N_4228,N_4146);
nor U4624 (N_4624,N_4439,N_4417);
or U4625 (N_4625,N_4214,N_4073);
nand U4626 (N_4626,N_4315,N_4010);
nand U4627 (N_4627,N_4282,N_4326);
nor U4628 (N_4628,N_4138,N_4360);
nor U4629 (N_4629,N_4055,N_4206);
or U4630 (N_4630,N_4022,N_4381);
or U4631 (N_4631,N_4396,N_4337);
nor U4632 (N_4632,N_4232,N_4144);
nand U4633 (N_4633,N_4488,N_4092);
nor U4634 (N_4634,N_4352,N_4020);
or U4635 (N_4635,N_4320,N_4461);
and U4636 (N_4636,N_4365,N_4485);
nand U4637 (N_4637,N_4089,N_4239);
and U4638 (N_4638,N_4497,N_4149);
or U4639 (N_4639,N_4457,N_4426);
xnor U4640 (N_4640,N_4427,N_4304);
or U4641 (N_4641,N_4184,N_4295);
nor U4642 (N_4642,N_4429,N_4262);
nor U4643 (N_4643,N_4387,N_4076);
xnor U4644 (N_4644,N_4409,N_4240);
or U4645 (N_4645,N_4204,N_4043);
nor U4646 (N_4646,N_4100,N_4308);
and U4647 (N_4647,N_4376,N_4369);
and U4648 (N_4648,N_4474,N_4493);
nand U4649 (N_4649,N_4309,N_4165);
nor U4650 (N_4650,N_4014,N_4470);
nor U4651 (N_4651,N_4190,N_4008);
xnor U4652 (N_4652,N_4410,N_4145);
nand U4653 (N_4653,N_4155,N_4357);
and U4654 (N_4654,N_4110,N_4182);
or U4655 (N_4655,N_4013,N_4385);
or U4656 (N_4656,N_4263,N_4293);
nor U4657 (N_4657,N_4383,N_4203);
nor U4658 (N_4658,N_4119,N_4215);
nor U4659 (N_4659,N_4413,N_4063);
or U4660 (N_4660,N_4181,N_4296);
nand U4661 (N_4661,N_4289,N_4037);
nor U4662 (N_4662,N_4157,N_4363);
nor U4663 (N_4663,N_4084,N_4344);
and U4664 (N_4664,N_4066,N_4054);
and U4665 (N_4665,N_4225,N_4176);
or U4666 (N_4666,N_4034,N_4453);
or U4667 (N_4667,N_4359,N_4021);
xnor U4668 (N_4668,N_4198,N_4213);
nor U4669 (N_4669,N_4226,N_4114);
and U4670 (N_4670,N_4141,N_4035);
nor U4671 (N_4671,N_4288,N_4229);
or U4672 (N_4672,N_4303,N_4432);
xor U4673 (N_4673,N_4373,N_4000);
or U4674 (N_4674,N_4271,N_4407);
and U4675 (N_4675,N_4351,N_4274);
and U4676 (N_4676,N_4058,N_4030);
xor U4677 (N_4677,N_4074,N_4199);
nand U4678 (N_4678,N_4094,N_4238);
nor U4679 (N_4679,N_4434,N_4191);
xnor U4680 (N_4680,N_4482,N_4221);
nand U4681 (N_4681,N_4317,N_4278);
nor U4682 (N_4682,N_4248,N_4105);
or U4683 (N_4683,N_4319,N_4067);
or U4684 (N_4684,N_4346,N_4444);
nand U4685 (N_4685,N_4127,N_4106);
nand U4686 (N_4686,N_4059,N_4464);
nand U4687 (N_4687,N_4285,N_4443);
xor U4688 (N_4688,N_4277,N_4111);
or U4689 (N_4689,N_4371,N_4329);
nand U4690 (N_4690,N_4356,N_4280);
nand U4691 (N_4691,N_4460,N_4197);
nand U4692 (N_4692,N_4338,N_4377);
nand U4693 (N_4693,N_4301,N_4235);
or U4694 (N_4694,N_4218,N_4436);
nand U4695 (N_4695,N_4166,N_4244);
and U4696 (N_4696,N_4026,N_4331);
nor U4697 (N_4697,N_4466,N_4173);
and U4698 (N_4698,N_4242,N_4124);
nand U4699 (N_4699,N_4481,N_4245);
or U4700 (N_4700,N_4192,N_4415);
nor U4701 (N_4701,N_4230,N_4078);
nor U4702 (N_4702,N_4388,N_4491);
or U4703 (N_4703,N_4494,N_4492);
or U4704 (N_4704,N_4375,N_4256);
or U4705 (N_4705,N_4322,N_4189);
xnor U4706 (N_4706,N_4390,N_4382);
nand U4707 (N_4707,N_4099,N_4246);
nor U4708 (N_4708,N_4272,N_4153);
nand U4709 (N_4709,N_4404,N_4048);
or U4710 (N_4710,N_4366,N_4115);
nand U4711 (N_4711,N_4224,N_4361);
xor U4712 (N_4712,N_4005,N_4098);
nand U4713 (N_4713,N_4328,N_4276);
xnor U4714 (N_4714,N_4160,N_4321);
nand U4715 (N_4715,N_4495,N_4446);
and U4716 (N_4716,N_4104,N_4270);
or U4717 (N_4717,N_4186,N_4208);
or U4718 (N_4718,N_4024,N_4251);
or U4719 (N_4719,N_4458,N_4137);
nor U4720 (N_4720,N_4210,N_4260);
or U4721 (N_4721,N_4237,N_4129);
and U4722 (N_4722,N_4264,N_4416);
nand U4723 (N_4723,N_4047,N_4023);
and U4724 (N_4724,N_4456,N_4070);
or U4725 (N_4725,N_4379,N_4292);
or U4726 (N_4726,N_4455,N_4412);
and U4727 (N_4727,N_4445,N_4028);
or U4728 (N_4728,N_4101,N_4401);
nand U4729 (N_4729,N_4131,N_4108);
xnor U4730 (N_4730,N_4498,N_4122);
nor U4731 (N_4731,N_4162,N_4354);
and U4732 (N_4732,N_4325,N_4438);
or U4733 (N_4733,N_4362,N_4486);
or U4734 (N_4734,N_4397,N_4039);
and U4735 (N_4735,N_4143,N_4462);
nand U4736 (N_4736,N_4499,N_4046);
or U4737 (N_4737,N_4253,N_4336);
nor U4738 (N_4738,N_4002,N_4487);
nor U4739 (N_4739,N_4291,N_4154);
or U4740 (N_4740,N_4077,N_4298);
or U4741 (N_4741,N_4437,N_4441);
nor U4742 (N_4742,N_4243,N_4102);
xnor U4743 (N_4743,N_4334,N_4452);
nand U4744 (N_4744,N_4061,N_4394);
or U4745 (N_4745,N_4123,N_4075);
nand U4746 (N_4746,N_4267,N_4408);
nor U4747 (N_4747,N_4219,N_4178);
and U4748 (N_4748,N_4036,N_4175);
nor U4749 (N_4749,N_4152,N_4279);
nand U4750 (N_4750,N_4344,N_4139);
or U4751 (N_4751,N_4488,N_4238);
xor U4752 (N_4752,N_4309,N_4362);
nand U4753 (N_4753,N_4190,N_4083);
nor U4754 (N_4754,N_4498,N_4391);
and U4755 (N_4755,N_4444,N_4130);
nand U4756 (N_4756,N_4306,N_4104);
nand U4757 (N_4757,N_4331,N_4255);
and U4758 (N_4758,N_4044,N_4426);
or U4759 (N_4759,N_4253,N_4366);
or U4760 (N_4760,N_4324,N_4105);
nor U4761 (N_4761,N_4212,N_4203);
nor U4762 (N_4762,N_4396,N_4423);
or U4763 (N_4763,N_4053,N_4132);
nand U4764 (N_4764,N_4105,N_4411);
or U4765 (N_4765,N_4208,N_4163);
nor U4766 (N_4766,N_4139,N_4448);
or U4767 (N_4767,N_4261,N_4146);
nor U4768 (N_4768,N_4198,N_4495);
nor U4769 (N_4769,N_4227,N_4128);
nand U4770 (N_4770,N_4477,N_4227);
nand U4771 (N_4771,N_4422,N_4213);
nor U4772 (N_4772,N_4058,N_4150);
or U4773 (N_4773,N_4368,N_4199);
or U4774 (N_4774,N_4353,N_4462);
nor U4775 (N_4775,N_4066,N_4304);
and U4776 (N_4776,N_4150,N_4227);
xnor U4777 (N_4777,N_4368,N_4404);
or U4778 (N_4778,N_4177,N_4009);
nor U4779 (N_4779,N_4077,N_4174);
and U4780 (N_4780,N_4022,N_4493);
nand U4781 (N_4781,N_4132,N_4474);
and U4782 (N_4782,N_4364,N_4346);
or U4783 (N_4783,N_4212,N_4233);
or U4784 (N_4784,N_4223,N_4175);
nand U4785 (N_4785,N_4174,N_4455);
nor U4786 (N_4786,N_4189,N_4273);
or U4787 (N_4787,N_4348,N_4106);
nand U4788 (N_4788,N_4113,N_4147);
xnor U4789 (N_4789,N_4350,N_4421);
nand U4790 (N_4790,N_4283,N_4155);
xnor U4791 (N_4791,N_4025,N_4490);
and U4792 (N_4792,N_4153,N_4348);
nand U4793 (N_4793,N_4082,N_4369);
or U4794 (N_4794,N_4294,N_4175);
or U4795 (N_4795,N_4419,N_4123);
or U4796 (N_4796,N_4013,N_4082);
nand U4797 (N_4797,N_4192,N_4207);
or U4798 (N_4798,N_4176,N_4449);
nor U4799 (N_4799,N_4251,N_4472);
xor U4800 (N_4800,N_4076,N_4456);
xor U4801 (N_4801,N_4166,N_4009);
nor U4802 (N_4802,N_4059,N_4351);
nor U4803 (N_4803,N_4480,N_4355);
nor U4804 (N_4804,N_4192,N_4007);
xnor U4805 (N_4805,N_4452,N_4251);
nor U4806 (N_4806,N_4215,N_4151);
and U4807 (N_4807,N_4028,N_4214);
nor U4808 (N_4808,N_4455,N_4492);
nand U4809 (N_4809,N_4330,N_4120);
or U4810 (N_4810,N_4019,N_4036);
and U4811 (N_4811,N_4391,N_4377);
and U4812 (N_4812,N_4464,N_4167);
or U4813 (N_4813,N_4177,N_4184);
and U4814 (N_4814,N_4087,N_4315);
and U4815 (N_4815,N_4424,N_4020);
and U4816 (N_4816,N_4318,N_4164);
or U4817 (N_4817,N_4044,N_4361);
xor U4818 (N_4818,N_4104,N_4310);
and U4819 (N_4819,N_4184,N_4429);
and U4820 (N_4820,N_4218,N_4259);
nor U4821 (N_4821,N_4099,N_4351);
or U4822 (N_4822,N_4185,N_4177);
or U4823 (N_4823,N_4294,N_4231);
nor U4824 (N_4824,N_4405,N_4276);
and U4825 (N_4825,N_4303,N_4135);
and U4826 (N_4826,N_4434,N_4150);
nand U4827 (N_4827,N_4374,N_4209);
nor U4828 (N_4828,N_4211,N_4308);
or U4829 (N_4829,N_4067,N_4189);
and U4830 (N_4830,N_4403,N_4379);
and U4831 (N_4831,N_4229,N_4442);
nor U4832 (N_4832,N_4023,N_4265);
xnor U4833 (N_4833,N_4145,N_4209);
and U4834 (N_4834,N_4147,N_4123);
or U4835 (N_4835,N_4089,N_4455);
nor U4836 (N_4836,N_4466,N_4067);
or U4837 (N_4837,N_4389,N_4167);
or U4838 (N_4838,N_4172,N_4230);
or U4839 (N_4839,N_4402,N_4286);
or U4840 (N_4840,N_4019,N_4071);
nand U4841 (N_4841,N_4238,N_4366);
nand U4842 (N_4842,N_4419,N_4026);
or U4843 (N_4843,N_4026,N_4499);
nor U4844 (N_4844,N_4373,N_4399);
nor U4845 (N_4845,N_4055,N_4204);
or U4846 (N_4846,N_4135,N_4025);
and U4847 (N_4847,N_4175,N_4299);
and U4848 (N_4848,N_4059,N_4271);
nor U4849 (N_4849,N_4422,N_4426);
or U4850 (N_4850,N_4166,N_4295);
nand U4851 (N_4851,N_4250,N_4045);
and U4852 (N_4852,N_4431,N_4357);
or U4853 (N_4853,N_4320,N_4192);
xnor U4854 (N_4854,N_4297,N_4275);
nor U4855 (N_4855,N_4031,N_4109);
nand U4856 (N_4856,N_4422,N_4386);
and U4857 (N_4857,N_4398,N_4259);
nand U4858 (N_4858,N_4007,N_4229);
xor U4859 (N_4859,N_4316,N_4086);
nor U4860 (N_4860,N_4303,N_4322);
nor U4861 (N_4861,N_4132,N_4411);
nand U4862 (N_4862,N_4419,N_4062);
nor U4863 (N_4863,N_4098,N_4150);
and U4864 (N_4864,N_4205,N_4416);
nand U4865 (N_4865,N_4446,N_4473);
or U4866 (N_4866,N_4056,N_4349);
and U4867 (N_4867,N_4446,N_4490);
or U4868 (N_4868,N_4357,N_4375);
and U4869 (N_4869,N_4356,N_4414);
or U4870 (N_4870,N_4199,N_4399);
and U4871 (N_4871,N_4381,N_4310);
nor U4872 (N_4872,N_4339,N_4314);
or U4873 (N_4873,N_4057,N_4186);
and U4874 (N_4874,N_4327,N_4408);
xnor U4875 (N_4875,N_4499,N_4221);
xor U4876 (N_4876,N_4006,N_4380);
or U4877 (N_4877,N_4472,N_4233);
nor U4878 (N_4878,N_4027,N_4385);
and U4879 (N_4879,N_4099,N_4251);
and U4880 (N_4880,N_4055,N_4405);
nand U4881 (N_4881,N_4195,N_4210);
nor U4882 (N_4882,N_4338,N_4264);
nor U4883 (N_4883,N_4007,N_4196);
or U4884 (N_4884,N_4061,N_4147);
or U4885 (N_4885,N_4318,N_4187);
or U4886 (N_4886,N_4280,N_4338);
nor U4887 (N_4887,N_4440,N_4436);
or U4888 (N_4888,N_4356,N_4218);
and U4889 (N_4889,N_4239,N_4206);
nand U4890 (N_4890,N_4390,N_4479);
or U4891 (N_4891,N_4046,N_4232);
or U4892 (N_4892,N_4094,N_4275);
xor U4893 (N_4893,N_4060,N_4132);
or U4894 (N_4894,N_4185,N_4206);
or U4895 (N_4895,N_4292,N_4354);
or U4896 (N_4896,N_4220,N_4359);
or U4897 (N_4897,N_4004,N_4019);
or U4898 (N_4898,N_4058,N_4085);
and U4899 (N_4899,N_4127,N_4293);
xnor U4900 (N_4900,N_4382,N_4277);
or U4901 (N_4901,N_4149,N_4405);
nor U4902 (N_4902,N_4435,N_4125);
or U4903 (N_4903,N_4003,N_4313);
or U4904 (N_4904,N_4394,N_4242);
nand U4905 (N_4905,N_4413,N_4016);
nor U4906 (N_4906,N_4285,N_4348);
and U4907 (N_4907,N_4119,N_4326);
and U4908 (N_4908,N_4267,N_4205);
xnor U4909 (N_4909,N_4194,N_4205);
and U4910 (N_4910,N_4084,N_4343);
nor U4911 (N_4911,N_4409,N_4051);
and U4912 (N_4912,N_4426,N_4258);
or U4913 (N_4913,N_4286,N_4220);
nor U4914 (N_4914,N_4245,N_4373);
nand U4915 (N_4915,N_4262,N_4484);
and U4916 (N_4916,N_4404,N_4120);
and U4917 (N_4917,N_4366,N_4285);
or U4918 (N_4918,N_4313,N_4442);
nor U4919 (N_4919,N_4317,N_4295);
nand U4920 (N_4920,N_4058,N_4433);
nor U4921 (N_4921,N_4097,N_4426);
and U4922 (N_4922,N_4435,N_4106);
xor U4923 (N_4923,N_4012,N_4356);
xnor U4924 (N_4924,N_4082,N_4128);
xnor U4925 (N_4925,N_4084,N_4360);
nand U4926 (N_4926,N_4481,N_4095);
nand U4927 (N_4927,N_4065,N_4089);
and U4928 (N_4928,N_4121,N_4227);
or U4929 (N_4929,N_4452,N_4064);
nor U4930 (N_4930,N_4484,N_4077);
and U4931 (N_4931,N_4421,N_4046);
and U4932 (N_4932,N_4134,N_4282);
nand U4933 (N_4933,N_4309,N_4181);
or U4934 (N_4934,N_4131,N_4176);
nor U4935 (N_4935,N_4429,N_4264);
and U4936 (N_4936,N_4172,N_4414);
nor U4937 (N_4937,N_4163,N_4271);
and U4938 (N_4938,N_4382,N_4294);
and U4939 (N_4939,N_4150,N_4199);
or U4940 (N_4940,N_4236,N_4419);
nor U4941 (N_4941,N_4107,N_4303);
nand U4942 (N_4942,N_4081,N_4001);
nor U4943 (N_4943,N_4034,N_4215);
nor U4944 (N_4944,N_4432,N_4319);
nor U4945 (N_4945,N_4450,N_4071);
xor U4946 (N_4946,N_4191,N_4240);
nand U4947 (N_4947,N_4401,N_4005);
and U4948 (N_4948,N_4146,N_4014);
and U4949 (N_4949,N_4027,N_4345);
or U4950 (N_4950,N_4462,N_4416);
and U4951 (N_4951,N_4108,N_4114);
or U4952 (N_4952,N_4399,N_4197);
nor U4953 (N_4953,N_4386,N_4120);
or U4954 (N_4954,N_4394,N_4355);
or U4955 (N_4955,N_4307,N_4289);
and U4956 (N_4956,N_4329,N_4450);
xor U4957 (N_4957,N_4287,N_4353);
xnor U4958 (N_4958,N_4230,N_4363);
xnor U4959 (N_4959,N_4154,N_4442);
nor U4960 (N_4960,N_4385,N_4114);
and U4961 (N_4961,N_4182,N_4368);
or U4962 (N_4962,N_4154,N_4155);
and U4963 (N_4963,N_4128,N_4071);
xnor U4964 (N_4964,N_4456,N_4150);
and U4965 (N_4965,N_4322,N_4180);
and U4966 (N_4966,N_4355,N_4495);
or U4967 (N_4967,N_4065,N_4353);
nor U4968 (N_4968,N_4014,N_4253);
nand U4969 (N_4969,N_4405,N_4234);
and U4970 (N_4970,N_4483,N_4306);
and U4971 (N_4971,N_4109,N_4479);
or U4972 (N_4972,N_4491,N_4497);
or U4973 (N_4973,N_4405,N_4040);
and U4974 (N_4974,N_4278,N_4107);
or U4975 (N_4975,N_4243,N_4193);
nand U4976 (N_4976,N_4453,N_4380);
and U4977 (N_4977,N_4082,N_4088);
and U4978 (N_4978,N_4270,N_4143);
nand U4979 (N_4979,N_4024,N_4398);
or U4980 (N_4980,N_4270,N_4276);
nor U4981 (N_4981,N_4185,N_4247);
nand U4982 (N_4982,N_4430,N_4220);
nand U4983 (N_4983,N_4445,N_4447);
nand U4984 (N_4984,N_4045,N_4275);
nor U4985 (N_4985,N_4283,N_4158);
nor U4986 (N_4986,N_4223,N_4475);
and U4987 (N_4987,N_4329,N_4449);
nor U4988 (N_4988,N_4393,N_4378);
nor U4989 (N_4989,N_4445,N_4023);
or U4990 (N_4990,N_4354,N_4330);
nand U4991 (N_4991,N_4133,N_4031);
or U4992 (N_4992,N_4189,N_4456);
xor U4993 (N_4993,N_4088,N_4097);
and U4994 (N_4994,N_4045,N_4103);
or U4995 (N_4995,N_4482,N_4408);
and U4996 (N_4996,N_4031,N_4163);
and U4997 (N_4997,N_4147,N_4290);
nand U4998 (N_4998,N_4102,N_4066);
nor U4999 (N_4999,N_4495,N_4426);
or U5000 (N_5000,N_4854,N_4538);
nand U5001 (N_5001,N_4666,N_4693);
xnor U5002 (N_5002,N_4741,N_4550);
or U5003 (N_5003,N_4851,N_4535);
nor U5004 (N_5004,N_4995,N_4711);
nor U5005 (N_5005,N_4793,N_4542);
nor U5006 (N_5006,N_4546,N_4732);
nor U5007 (N_5007,N_4824,N_4888);
or U5008 (N_5008,N_4744,N_4799);
nand U5009 (N_5009,N_4841,N_4567);
or U5010 (N_5010,N_4961,N_4707);
nor U5011 (N_5011,N_4844,N_4846);
nor U5012 (N_5012,N_4768,N_4674);
nand U5013 (N_5013,N_4624,N_4733);
nand U5014 (N_5014,N_4684,N_4808);
or U5015 (N_5015,N_4689,N_4729);
and U5016 (N_5016,N_4900,N_4775);
or U5017 (N_5017,N_4529,N_4970);
and U5018 (N_5018,N_4797,N_4985);
or U5019 (N_5019,N_4734,N_4918);
nand U5020 (N_5020,N_4610,N_4556);
and U5021 (N_5021,N_4620,N_4770);
nand U5022 (N_5022,N_4524,N_4941);
and U5023 (N_5023,N_4518,N_4613);
nor U5024 (N_5024,N_4834,N_4944);
nor U5025 (N_5025,N_4719,N_4783);
and U5026 (N_5026,N_4519,N_4974);
nor U5027 (N_5027,N_4656,N_4581);
nand U5028 (N_5028,N_4641,N_4776);
nor U5029 (N_5029,N_4644,N_4560);
or U5030 (N_5030,N_4767,N_4902);
and U5031 (N_5031,N_4833,N_4738);
and U5032 (N_5032,N_4779,N_4572);
nor U5033 (N_5033,N_4747,N_4587);
and U5034 (N_5034,N_4688,N_4790);
and U5035 (N_5035,N_4821,N_4825);
xnor U5036 (N_5036,N_4883,N_4607);
or U5037 (N_5037,N_4751,N_4817);
or U5038 (N_5038,N_4971,N_4969);
or U5039 (N_5039,N_4862,N_4919);
nor U5040 (N_5040,N_4989,N_4810);
nor U5041 (N_5041,N_4715,N_4891);
or U5042 (N_5042,N_4530,N_4822);
or U5043 (N_5043,N_4877,N_4875);
nor U5044 (N_5044,N_4921,N_4925);
nor U5045 (N_5045,N_4811,N_4651);
nor U5046 (N_5046,N_4664,N_4690);
and U5047 (N_5047,N_4720,N_4762);
xor U5048 (N_5048,N_4743,N_4653);
nor U5049 (N_5049,N_4668,N_4692);
and U5050 (N_5050,N_4894,N_4864);
nand U5051 (N_5051,N_4574,N_4643);
nor U5052 (N_5052,N_4927,N_4831);
or U5053 (N_5053,N_4827,N_4706);
and U5054 (N_5054,N_4951,N_4952);
nor U5055 (N_5055,N_4502,N_4739);
or U5056 (N_5056,N_4874,N_4604);
nor U5057 (N_5057,N_4848,N_4594);
or U5058 (N_5058,N_4920,N_4922);
nor U5059 (N_5059,N_4721,N_4893);
nor U5060 (N_5060,N_4553,N_4716);
xnor U5061 (N_5061,N_4953,N_4508);
nand U5062 (N_5062,N_4507,N_4677);
nor U5063 (N_5063,N_4724,N_4740);
and U5064 (N_5064,N_4788,N_4980);
nand U5065 (N_5065,N_4742,N_4512);
nand U5066 (N_5066,N_4837,N_4596);
xnor U5067 (N_5067,N_4615,N_4531);
nand U5068 (N_5068,N_4806,N_4930);
xnor U5069 (N_5069,N_4622,N_4801);
nand U5070 (N_5070,N_4557,N_4761);
and U5071 (N_5071,N_4785,N_4540);
nor U5072 (N_5072,N_4517,N_4547);
nor U5073 (N_5073,N_4972,N_4682);
and U5074 (N_5074,N_4936,N_4601);
and U5075 (N_5075,N_4552,N_4781);
and U5076 (N_5076,N_4598,N_4608);
nand U5077 (N_5077,N_4662,N_4988);
or U5078 (N_5078,N_4544,N_4857);
or U5079 (N_5079,N_4654,N_4994);
nor U5080 (N_5080,N_4513,N_4606);
and U5081 (N_5081,N_4726,N_4898);
xor U5082 (N_5082,N_4561,N_4536);
or U5083 (N_5083,N_4939,N_4670);
or U5084 (N_5084,N_4959,N_4655);
nor U5085 (N_5085,N_4566,N_4709);
nand U5086 (N_5086,N_4573,N_4990);
xor U5087 (N_5087,N_4602,N_4886);
xnor U5088 (N_5088,N_4605,N_4982);
nor U5089 (N_5089,N_4943,N_4603);
nand U5090 (N_5090,N_4926,N_4816);
nor U5091 (N_5091,N_4820,N_4755);
nand U5092 (N_5092,N_4847,N_4996);
nand U5093 (N_5093,N_4881,N_4619);
xnor U5094 (N_5094,N_4850,N_4583);
nor U5095 (N_5095,N_4954,N_4597);
and U5096 (N_5096,N_4599,N_4828);
and U5097 (N_5097,N_4766,N_4876);
and U5098 (N_5098,N_4955,N_4510);
or U5099 (N_5099,N_4647,N_4749);
nor U5100 (N_5100,N_4983,N_4814);
nand U5101 (N_5101,N_4646,N_4802);
nand U5102 (N_5102,N_4813,N_4906);
and U5103 (N_5103,N_4873,N_4782);
and U5104 (N_5104,N_4504,N_4697);
or U5105 (N_5105,N_4549,N_4748);
nor U5106 (N_5106,N_4687,N_4777);
nor U5107 (N_5107,N_4611,N_4703);
or U5108 (N_5108,N_4609,N_4616);
or U5109 (N_5109,N_4992,N_4849);
nor U5110 (N_5110,N_4853,N_4946);
nor U5111 (N_5111,N_4856,N_4924);
nor U5112 (N_5112,N_4855,N_4842);
nor U5113 (N_5113,N_4570,N_4691);
nand U5114 (N_5114,N_4780,N_4869);
and U5115 (N_5115,N_4913,N_4578);
or U5116 (N_5116,N_4577,N_4750);
nand U5117 (N_5117,N_4548,N_4859);
and U5118 (N_5118,N_4640,N_4576);
or U5119 (N_5119,N_4503,N_4683);
or U5120 (N_5120,N_4628,N_4696);
nor U5121 (N_5121,N_4589,N_4977);
nor U5122 (N_5122,N_4963,N_4809);
or U5123 (N_5123,N_4635,N_4978);
nand U5124 (N_5124,N_4966,N_4673);
or U5125 (N_5125,N_4665,N_4658);
nand U5126 (N_5126,N_4541,N_4812);
or U5127 (N_5127,N_4889,N_4559);
or U5128 (N_5128,N_4865,N_4890);
nor U5129 (N_5129,N_4752,N_4554);
nand U5130 (N_5130,N_4829,N_4964);
or U5131 (N_5131,N_4736,N_4975);
nand U5132 (N_5132,N_4958,N_4705);
nor U5133 (N_5133,N_4579,N_4884);
and U5134 (N_5134,N_4712,N_4642);
nor U5135 (N_5135,N_4872,N_4648);
xnor U5136 (N_5136,N_4725,N_4614);
nand U5137 (N_5137,N_4746,N_4999);
or U5138 (N_5138,N_4632,N_4979);
and U5139 (N_5139,N_4997,N_4626);
and U5140 (N_5140,N_4882,N_4933);
or U5141 (N_5141,N_4571,N_4823);
or U5142 (N_5142,N_4534,N_4835);
and U5143 (N_5143,N_4595,N_4678);
nor U5144 (N_5144,N_4652,N_4986);
or U5145 (N_5145,N_4600,N_4672);
nand U5146 (N_5146,N_4764,N_4686);
nor U5147 (N_5147,N_4700,N_4965);
nor U5148 (N_5148,N_4545,N_4588);
and U5149 (N_5149,N_4500,N_4501);
nand U5150 (N_5150,N_4937,N_4843);
nand U5151 (N_5151,N_4629,N_4657);
nand U5152 (N_5152,N_4520,N_4984);
nor U5153 (N_5153,N_4962,N_4634);
and U5154 (N_5154,N_4774,N_4728);
nor U5155 (N_5155,N_4526,N_4798);
or U5156 (N_5156,N_4525,N_4815);
nor U5157 (N_5157,N_4956,N_4592);
and U5158 (N_5158,N_4722,N_4704);
or U5159 (N_5159,N_4830,N_4586);
nand U5160 (N_5160,N_4879,N_4617);
and U5161 (N_5161,N_4660,N_4866);
xnor U5162 (N_5162,N_4940,N_4568);
nand U5163 (N_5163,N_4923,N_4805);
nand U5164 (N_5164,N_4532,N_4543);
nand U5165 (N_5165,N_4772,N_4905);
nand U5166 (N_5166,N_4717,N_4645);
xor U5167 (N_5167,N_4737,N_4511);
and U5168 (N_5168,N_4950,N_4506);
and U5169 (N_5169,N_4897,N_4911);
nor U5170 (N_5170,N_4659,N_4671);
nand U5171 (N_5171,N_4695,N_4917);
nor U5172 (N_5172,N_4794,N_4967);
and U5173 (N_5173,N_4727,N_4871);
nor U5174 (N_5174,N_4533,N_4714);
nand U5175 (N_5175,N_4908,N_4760);
nand U5176 (N_5176,N_4580,N_4957);
nand U5177 (N_5177,N_4915,N_4590);
nor U5178 (N_5178,N_4934,N_4896);
nor U5179 (N_5179,N_4522,N_4991);
nand U5180 (N_5180,N_4998,N_4636);
nor U5181 (N_5181,N_4637,N_4753);
or U5182 (N_5182,N_4555,N_4591);
xor U5183 (N_5183,N_4968,N_4558);
nand U5184 (N_5184,N_4885,N_4718);
and U5185 (N_5185,N_4551,N_4675);
and U5186 (N_5186,N_4904,N_4702);
nor U5187 (N_5187,N_4796,N_4639);
and U5188 (N_5188,N_4912,N_4633);
xor U5189 (N_5189,N_4771,N_4505);
or U5190 (N_5190,N_4840,N_4987);
nor U5191 (N_5191,N_4903,N_4778);
or U5192 (N_5192,N_4993,N_4701);
or U5193 (N_5193,N_4731,N_4887);
and U5194 (N_5194,N_4839,N_4563);
and U5195 (N_5195,N_4769,N_4773);
and U5196 (N_5196,N_4523,N_4763);
or U5197 (N_5197,N_4676,N_4756);
or U5198 (N_5198,N_4860,N_4757);
nand U5199 (N_5199,N_4521,N_4758);
xnor U5200 (N_5200,N_4537,N_4575);
nand U5201 (N_5201,N_4623,N_4612);
nand U5202 (N_5202,N_4784,N_4932);
and U5203 (N_5203,N_4618,N_4981);
nor U5204 (N_5204,N_4680,N_4907);
and U5205 (N_5205,N_4945,N_4514);
and U5206 (N_5206,N_4928,N_4949);
or U5207 (N_5207,N_4650,N_4527);
and U5208 (N_5208,N_4807,N_4792);
nand U5209 (N_5209,N_4787,N_4858);
nor U5210 (N_5210,N_4948,N_4867);
or U5211 (N_5211,N_4745,N_4832);
nor U5212 (N_5212,N_4562,N_4661);
and U5213 (N_5213,N_4649,N_4730);
or U5214 (N_5214,N_4870,N_4947);
and U5215 (N_5215,N_4786,N_4931);
or U5216 (N_5216,N_4698,N_4723);
nand U5217 (N_5217,N_4679,N_4804);
and U5218 (N_5218,N_4838,N_4789);
and U5219 (N_5219,N_4515,N_4667);
nand U5220 (N_5220,N_4892,N_4584);
nor U5221 (N_5221,N_4909,N_4929);
and U5222 (N_5222,N_4569,N_4735);
nor U5223 (N_5223,N_4935,N_4819);
nor U5224 (N_5224,N_4539,N_4916);
or U5225 (N_5225,N_4630,N_4868);
xnor U5226 (N_5226,N_4826,N_4976);
nand U5227 (N_5227,N_4694,N_4631);
and U5228 (N_5228,N_4910,N_4516);
and U5229 (N_5229,N_4509,N_4759);
or U5230 (N_5230,N_4528,N_4914);
and U5231 (N_5231,N_4564,N_4699);
and U5232 (N_5232,N_4836,N_4818);
nand U5233 (N_5233,N_4663,N_4582);
nand U5234 (N_5234,N_4973,N_4852);
or U5235 (N_5235,N_4861,N_4625);
nand U5236 (N_5236,N_4585,N_4845);
nand U5237 (N_5237,N_4795,N_4713);
nand U5238 (N_5238,N_4638,N_4895);
nand U5239 (N_5239,N_4565,N_4710);
nor U5240 (N_5240,N_4765,N_4938);
or U5241 (N_5241,N_4878,N_4942);
and U5242 (N_5242,N_4627,N_4863);
or U5243 (N_5243,N_4681,N_4669);
nand U5244 (N_5244,N_4791,N_4800);
nor U5245 (N_5245,N_4708,N_4685);
nor U5246 (N_5246,N_4803,N_4593);
and U5247 (N_5247,N_4754,N_4880);
or U5248 (N_5248,N_4621,N_4901);
or U5249 (N_5249,N_4960,N_4899);
nor U5250 (N_5250,N_4697,N_4633);
xor U5251 (N_5251,N_4686,N_4960);
and U5252 (N_5252,N_4545,N_4607);
or U5253 (N_5253,N_4597,N_4696);
and U5254 (N_5254,N_4763,N_4917);
nand U5255 (N_5255,N_4685,N_4858);
or U5256 (N_5256,N_4741,N_4901);
and U5257 (N_5257,N_4627,N_4689);
nand U5258 (N_5258,N_4958,N_4923);
or U5259 (N_5259,N_4976,N_4564);
and U5260 (N_5260,N_4673,N_4701);
or U5261 (N_5261,N_4673,N_4831);
nand U5262 (N_5262,N_4924,N_4717);
xor U5263 (N_5263,N_4923,N_4797);
and U5264 (N_5264,N_4951,N_4767);
or U5265 (N_5265,N_4590,N_4933);
or U5266 (N_5266,N_4610,N_4648);
and U5267 (N_5267,N_4772,N_4940);
nand U5268 (N_5268,N_4911,N_4678);
nor U5269 (N_5269,N_4602,N_4507);
and U5270 (N_5270,N_4521,N_4957);
xnor U5271 (N_5271,N_4719,N_4856);
nand U5272 (N_5272,N_4529,N_4692);
nand U5273 (N_5273,N_4808,N_4675);
xnor U5274 (N_5274,N_4666,N_4967);
nor U5275 (N_5275,N_4979,N_4973);
xor U5276 (N_5276,N_4543,N_4953);
nor U5277 (N_5277,N_4567,N_4636);
nand U5278 (N_5278,N_4601,N_4726);
nor U5279 (N_5279,N_4850,N_4972);
nand U5280 (N_5280,N_4763,N_4581);
or U5281 (N_5281,N_4902,N_4885);
xor U5282 (N_5282,N_4864,N_4918);
and U5283 (N_5283,N_4735,N_4934);
and U5284 (N_5284,N_4872,N_4798);
nand U5285 (N_5285,N_4541,N_4794);
and U5286 (N_5286,N_4902,N_4512);
nor U5287 (N_5287,N_4595,N_4694);
nor U5288 (N_5288,N_4688,N_4859);
nor U5289 (N_5289,N_4990,N_4936);
xnor U5290 (N_5290,N_4700,N_4768);
or U5291 (N_5291,N_4942,N_4971);
nor U5292 (N_5292,N_4995,N_4899);
xor U5293 (N_5293,N_4779,N_4976);
xnor U5294 (N_5294,N_4927,N_4993);
nor U5295 (N_5295,N_4718,N_4762);
nor U5296 (N_5296,N_4509,N_4622);
nor U5297 (N_5297,N_4970,N_4564);
or U5298 (N_5298,N_4703,N_4841);
and U5299 (N_5299,N_4759,N_4857);
nor U5300 (N_5300,N_4652,N_4605);
or U5301 (N_5301,N_4509,N_4981);
nor U5302 (N_5302,N_4536,N_4706);
or U5303 (N_5303,N_4934,N_4973);
nor U5304 (N_5304,N_4973,N_4816);
and U5305 (N_5305,N_4810,N_4748);
or U5306 (N_5306,N_4628,N_4844);
nand U5307 (N_5307,N_4738,N_4977);
or U5308 (N_5308,N_4622,N_4684);
nor U5309 (N_5309,N_4737,N_4748);
nor U5310 (N_5310,N_4993,N_4788);
nor U5311 (N_5311,N_4985,N_4737);
nand U5312 (N_5312,N_4820,N_4925);
nand U5313 (N_5313,N_4598,N_4766);
or U5314 (N_5314,N_4841,N_4808);
nand U5315 (N_5315,N_4572,N_4723);
and U5316 (N_5316,N_4526,N_4705);
nand U5317 (N_5317,N_4907,N_4990);
nand U5318 (N_5318,N_4792,N_4829);
nand U5319 (N_5319,N_4631,N_4733);
or U5320 (N_5320,N_4751,N_4598);
nand U5321 (N_5321,N_4605,N_4998);
or U5322 (N_5322,N_4846,N_4915);
nand U5323 (N_5323,N_4809,N_4853);
and U5324 (N_5324,N_4909,N_4901);
nand U5325 (N_5325,N_4916,N_4871);
and U5326 (N_5326,N_4677,N_4567);
nand U5327 (N_5327,N_4845,N_4688);
or U5328 (N_5328,N_4631,N_4593);
or U5329 (N_5329,N_4677,N_4758);
nand U5330 (N_5330,N_4969,N_4555);
and U5331 (N_5331,N_4591,N_4552);
and U5332 (N_5332,N_4564,N_4615);
nor U5333 (N_5333,N_4961,N_4581);
and U5334 (N_5334,N_4816,N_4920);
nor U5335 (N_5335,N_4536,N_4947);
nand U5336 (N_5336,N_4846,N_4954);
or U5337 (N_5337,N_4787,N_4774);
and U5338 (N_5338,N_4702,N_4691);
and U5339 (N_5339,N_4510,N_4900);
nand U5340 (N_5340,N_4912,N_4743);
or U5341 (N_5341,N_4864,N_4951);
nor U5342 (N_5342,N_4557,N_4649);
nor U5343 (N_5343,N_4540,N_4640);
nand U5344 (N_5344,N_4634,N_4813);
or U5345 (N_5345,N_4946,N_4767);
xor U5346 (N_5346,N_4809,N_4808);
and U5347 (N_5347,N_4788,N_4675);
xor U5348 (N_5348,N_4672,N_4942);
nor U5349 (N_5349,N_4706,N_4757);
nor U5350 (N_5350,N_4843,N_4583);
and U5351 (N_5351,N_4540,N_4738);
nand U5352 (N_5352,N_4585,N_4526);
nor U5353 (N_5353,N_4643,N_4612);
xor U5354 (N_5354,N_4583,N_4704);
and U5355 (N_5355,N_4541,N_4607);
nor U5356 (N_5356,N_4790,N_4725);
or U5357 (N_5357,N_4931,N_4654);
and U5358 (N_5358,N_4632,N_4676);
and U5359 (N_5359,N_4907,N_4976);
xor U5360 (N_5360,N_4870,N_4708);
or U5361 (N_5361,N_4827,N_4653);
nor U5362 (N_5362,N_4861,N_4653);
or U5363 (N_5363,N_4551,N_4688);
or U5364 (N_5364,N_4704,N_4506);
xor U5365 (N_5365,N_4778,N_4571);
or U5366 (N_5366,N_4961,N_4921);
nor U5367 (N_5367,N_4626,N_4858);
nor U5368 (N_5368,N_4652,N_4763);
xnor U5369 (N_5369,N_4700,N_4931);
nor U5370 (N_5370,N_4622,N_4737);
or U5371 (N_5371,N_4818,N_4832);
or U5372 (N_5372,N_4883,N_4804);
xor U5373 (N_5373,N_4747,N_4779);
nand U5374 (N_5374,N_4836,N_4547);
xor U5375 (N_5375,N_4707,N_4993);
nand U5376 (N_5376,N_4937,N_4697);
xnor U5377 (N_5377,N_4587,N_4577);
nor U5378 (N_5378,N_4658,N_4979);
and U5379 (N_5379,N_4824,N_4565);
xor U5380 (N_5380,N_4891,N_4996);
nor U5381 (N_5381,N_4911,N_4877);
or U5382 (N_5382,N_4566,N_4857);
nand U5383 (N_5383,N_4568,N_4730);
nand U5384 (N_5384,N_4512,N_4895);
or U5385 (N_5385,N_4666,N_4676);
or U5386 (N_5386,N_4971,N_4986);
or U5387 (N_5387,N_4686,N_4693);
and U5388 (N_5388,N_4866,N_4713);
nor U5389 (N_5389,N_4840,N_4699);
and U5390 (N_5390,N_4572,N_4888);
nand U5391 (N_5391,N_4958,N_4681);
nand U5392 (N_5392,N_4755,N_4568);
nand U5393 (N_5393,N_4847,N_4674);
and U5394 (N_5394,N_4845,N_4530);
nor U5395 (N_5395,N_4828,N_4879);
nor U5396 (N_5396,N_4910,N_4927);
and U5397 (N_5397,N_4928,N_4901);
xor U5398 (N_5398,N_4815,N_4855);
nand U5399 (N_5399,N_4758,N_4889);
nand U5400 (N_5400,N_4624,N_4889);
or U5401 (N_5401,N_4855,N_4776);
nand U5402 (N_5402,N_4883,N_4999);
nand U5403 (N_5403,N_4539,N_4991);
and U5404 (N_5404,N_4528,N_4545);
nand U5405 (N_5405,N_4883,N_4577);
nor U5406 (N_5406,N_4999,N_4993);
nor U5407 (N_5407,N_4956,N_4941);
nor U5408 (N_5408,N_4642,N_4890);
nand U5409 (N_5409,N_4656,N_4873);
nor U5410 (N_5410,N_4895,N_4535);
or U5411 (N_5411,N_4524,N_4690);
nor U5412 (N_5412,N_4947,N_4815);
nor U5413 (N_5413,N_4956,N_4888);
nand U5414 (N_5414,N_4827,N_4865);
and U5415 (N_5415,N_4576,N_4968);
nand U5416 (N_5416,N_4555,N_4835);
xnor U5417 (N_5417,N_4707,N_4904);
nor U5418 (N_5418,N_4823,N_4738);
or U5419 (N_5419,N_4514,N_4693);
nand U5420 (N_5420,N_4930,N_4977);
nand U5421 (N_5421,N_4767,N_4795);
or U5422 (N_5422,N_4900,N_4822);
nand U5423 (N_5423,N_4866,N_4856);
and U5424 (N_5424,N_4885,N_4737);
or U5425 (N_5425,N_4618,N_4918);
and U5426 (N_5426,N_4951,N_4520);
nor U5427 (N_5427,N_4764,N_4821);
nor U5428 (N_5428,N_4920,N_4649);
or U5429 (N_5429,N_4754,N_4530);
nand U5430 (N_5430,N_4584,N_4833);
nand U5431 (N_5431,N_4807,N_4865);
nand U5432 (N_5432,N_4542,N_4963);
nor U5433 (N_5433,N_4715,N_4945);
xor U5434 (N_5434,N_4809,N_4953);
nand U5435 (N_5435,N_4513,N_4860);
nor U5436 (N_5436,N_4947,N_4727);
nand U5437 (N_5437,N_4583,N_4913);
xor U5438 (N_5438,N_4524,N_4699);
nor U5439 (N_5439,N_4855,N_4783);
nand U5440 (N_5440,N_4762,N_4619);
nor U5441 (N_5441,N_4696,N_4719);
nand U5442 (N_5442,N_4899,N_4554);
nor U5443 (N_5443,N_4668,N_4539);
and U5444 (N_5444,N_4948,N_4610);
nand U5445 (N_5445,N_4795,N_4832);
and U5446 (N_5446,N_4515,N_4870);
or U5447 (N_5447,N_4557,N_4743);
or U5448 (N_5448,N_4596,N_4707);
or U5449 (N_5449,N_4780,N_4797);
or U5450 (N_5450,N_4800,N_4958);
or U5451 (N_5451,N_4947,N_4608);
and U5452 (N_5452,N_4709,N_4796);
and U5453 (N_5453,N_4862,N_4509);
or U5454 (N_5454,N_4887,N_4809);
nand U5455 (N_5455,N_4689,N_4839);
nand U5456 (N_5456,N_4561,N_4905);
xor U5457 (N_5457,N_4666,N_4872);
or U5458 (N_5458,N_4686,N_4609);
or U5459 (N_5459,N_4749,N_4885);
nor U5460 (N_5460,N_4746,N_4885);
nor U5461 (N_5461,N_4824,N_4790);
nor U5462 (N_5462,N_4584,N_4715);
nor U5463 (N_5463,N_4749,N_4768);
xnor U5464 (N_5464,N_4809,N_4855);
nor U5465 (N_5465,N_4942,N_4891);
or U5466 (N_5466,N_4776,N_4843);
nand U5467 (N_5467,N_4860,N_4941);
or U5468 (N_5468,N_4831,N_4983);
and U5469 (N_5469,N_4674,N_4539);
nor U5470 (N_5470,N_4811,N_4710);
and U5471 (N_5471,N_4827,N_4671);
or U5472 (N_5472,N_4681,N_4528);
xor U5473 (N_5473,N_4885,N_4632);
nand U5474 (N_5474,N_4786,N_4697);
or U5475 (N_5475,N_4762,N_4792);
or U5476 (N_5476,N_4792,N_4734);
nor U5477 (N_5477,N_4933,N_4787);
nor U5478 (N_5478,N_4601,N_4792);
and U5479 (N_5479,N_4737,N_4732);
nor U5480 (N_5480,N_4866,N_4604);
or U5481 (N_5481,N_4866,N_4844);
nor U5482 (N_5482,N_4834,N_4671);
xnor U5483 (N_5483,N_4997,N_4758);
nand U5484 (N_5484,N_4685,N_4953);
and U5485 (N_5485,N_4917,N_4506);
nand U5486 (N_5486,N_4801,N_4981);
and U5487 (N_5487,N_4844,N_4551);
or U5488 (N_5488,N_4616,N_4706);
nand U5489 (N_5489,N_4746,N_4961);
nand U5490 (N_5490,N_4973,N_4766);
nand U5491 (N_5491,N_4769,N_4842);
and U5492 (N_5492,N_4714,N_4607);
or U5493 (N_5493,N_4827,N_4577);
nand U5494 (N_5494,N_4578,N_4575);
nand U5495 (N_5495,N_4552,N_4939);
nand U5496 (N_5496,N_4804,N_4938);
and U5497 (N_5497,N_4748,N_4618);
nor U5498 (N_5498,N_4645,N_4593);
nand U5499 (N_5499,N_4728,N_4737);
nor U5500 (N_5500,N_5154,N_5273);
xnor U5501 (N_5501,N_5019,N_5416);
nand U5502 (N_5502,N_5294,N_5405);
or U5503 (N_5503,N_5151,N_5399);
or U5504 (N_5504,N_5099,N_5062);
nand U5505 (N_5505,N_5125,N_5469);
nand U5506 (N_5506,N_5331,N_5404);
nand U5507 (N_5507,N_5045,N_5353);
and U5508 (N_5508,N_5270,N_5395);
nor U5509 (N_5509,N_5021,N_5356);
or U5510 (N_5510,N_5265,N_5417);
and U5511 (N_5511,N_5166,N_5298);
nor U5512 (N_5512,N_5106,N_5279);
or U5513 (N_5513,N_5187,N_5016);
and U5514 (N_5514,N_5182,N_5177);
and U5515 (N_5515,N_5079,N_5025);
nor U5516 (N_5516,N_5179,N_5233);
and U5517 (N_5517,N_5336,N_5198);
or U5518 (N_5518,N_5303,N_5199);
or U5519 (N_5519,N_5332,N_5058);
xor U5520 (N_5520,N_5367,N_5039);
nand U5521 (N_5521,N_5114,N_5387);
nand U5522 (N_5522,N_5436,N_5357);
xor U5523 (N_5523,N_5118,N_5388);
and U5524 (N_5524,N_5171,N_5197);
or U5525 (N_5525,N_5359,N_5204);
nor U5526 (N_5526,N_5061,N_5278);
or U5527 (N_5527,N_5013,N_5479);
xnor U5528 (N_5528,N_5004,N_5186);
nand U5529 (N_5529,N_5443,N_5433);
nor U5530 (N_5530,N_5059,N_5421);
nand U5531 (N_5531,N_5373,N_5306);
nand U5532 (N_5532,N_5441,N_5254);
or U5533 (N_5533,N_5223,N_5425);
or U5534 (N_5534,N_5091,N_5145);
xnor U5535 (N_5535,N_5320,N_5050);
nor U5536 (N_5536,N_5028,N_5261);
nand U5537 (N_5537,N_5322,N_5364);
or U5538 (N_5538,N_5159,N_5398);
nand U5539 (N_5539,N_5499,N_5007);
nand U5540 (N_5540,N_5326,N_5232);
or U5541 (N_5541,N_5474,N_5108);
nand U5542 (N_5542,N_5227,N_5253);
nor U5543 (N_5543,N_5147,N_5299);
and U5544 (N_5544,N_5445,N_5415);
or U5545 (N_5545,N_5226,N_5496);
or U5546 (N_5546,N_5170,N_5066);
and U5547 (N_5547,N_5112,N_5313);
nand U5548 (N_5548,N_5252,N_5117);
nor U5549 (N_5549,N_5491,N_5456);
nor U5550 (N_5550,N_5480,N_5259);
nand U5551 (N_5551,N_5427,N_5375);
and U5552 (N_5552,N_5140,N_5082);
nor U5553 (N_5553,N_5296,N_5494);
nand U5554 (N_5554,N_5408,N_5422);
nand U5555 (N_5555,N_5195,N_5161);
or U5556 (N_5556,N_5192,N_5003);
nor U5557 (N_5557,N_5263,N_5418);
or U5558 (N_5558,N_5208,N_5428);
or U5559 (N_5559,N_5053,N_5096);
nor U5560 (N_5560,N_5384,N_5123);
nand U5561 (N_5561,N_5219,N_5142);
and U5562 (N_5562,N_5409,N_5430);
and U5563 (N_5563,N_5344,N_5495);
or U5564 (N_5564,N_5368,N_5318);
xor U5565 (N_5565,N_5075,N_5287);
nand U5566 (N_5566,N_5295,N_5153);
nor U5567 (N_5567,N_5293,N_5215);
or U5568 (N_5568,N_5150,N_5349);
nand U5569 (N_5569,N_5401,N_5483);
nor U5570 (N_5570,N_5184,N_5243);
and U5571 (N_5571,N_5010,N_5221);
nor U5572 (N_5572,N_5037,N_5244);
and U5573 (N_5573,N_5248,N_5202);
nor U5574 (N_5574,N_5193,N_5334);
nor U5575 (N_5575,N_5435,N_5167);
or U5576 (N_5576,N_5354,N_5319);
nor U5577 (N_5577,N_5222,N_5157);
nor U5578 (N_5578,N_5042,N_5097);
or U5579 (N_5579,N_5001,N_5070);
or U5580 (N_5580,N_5292,N_5149);
or U5581 (N_5581,N_5277,N_5385);
nor U5582 (N_5582,N_5046,N_5341);
xnor U5583 (N_5583,N_5172,N_5266);
nor U5584 (N_5584,N_5146,N_5251);
nor U5585 (N_5585,N_5498,N_5009);
nand U5586 (N_5586,N_5458,N_5047);
nor U5587 (N_5587,N_5185,N_5086);
and U5588 (N_5588,N_5238,N_5486);
or U5589 (N_5589,N_5450,N_5429);
nor U5590 (N_5590,N_5181,N_5413);
nor U5591 (N_5591,N_5081,N_5139);
nor U5592 (N_5592,N_5453,N_5020);
or U5593 (N_5593,N_5236,N_5459);
or U5594 (N_5594,N_5497,N_5345);
nor U5595 (N_5595,N_5103,N_5271);
and U5596 (N_5596,N_5328,N_5214);
nand U5597 (N_5597,N_5262,N_5347);
or U5598 (N_5598,N_5481,N_5390);
nand U5599 (N_5599,N_5023,N_5454);
and U5600 (N_5600,N_5035,N_5311);
nand U5601 (N_5601,N_5281,N_5191);
and U5602 (N_5602,N_5131,N_5457);
xnor U5603 (N_5603,N_5463,N_5230);
nand U5604 (N_5604,N_5340,N_5006);
and U5605 (N_5605,N_5231,N_5174);
and U5606 (N_5606,N_5471,N_5464);
and U5607 (N_5607,N_5370,N_5069);
or U5608 (N_5608,N_5073,N_5462);
and U5609 (N_5609,N_5129,N_5064);
xnor U5610 (N_5610,N_5475,N_5235);
xor U5611 (N_5611,N_5011,N_5485);
nor U5612 (N_5612,N_5107,N_5228);
and U5613 (N_5613,N_5285,N_5310);
nand U5614 (N_5614,N_5164,N_5284);
and U5615 (N_5615,N_5120,N_5424);
xor U5616 (N_5616,N_5201,N_5488);
nand U5617 (N_5617,N_5031,N_5196);
and U5618 (N_5618,N_5054,N_5321);
or U5619 (N_5619,N_5000,N_5268);
nor U5620 (N_5620,N_5034,N_5030);
or U5621 (N_5621,N_5329,N_5297);
and U5622 (N_5622,N_5205,N_5363);
or U5623 (N_5623,N_5478,N_5178);
nor U5624 (N_5624,N_5074,N_5324);
xnor U5625 (N_5625,N_5314,N_5100);
or U5626 (N_5626,N_5124,N_5432);
xnor U5627 (N_5627,N_5440,N_5209);
and U5628 (N_5628,N_5304,N_5465);
or U5629 (N_5629,N_5141,N_5048);
or U5630 (N_5630,N_5126,N_5451);
xor U5631 (N_5631,N_5335,N_5206);
or U5632 (N_5632,N_5234,N_5378);
nand U5633 (N_5633,N_5449,N_5121);
nor U5634 (N_5634,N_5043,N_5022);
nand U5635 (N_5635,N_5267,N_5275);
and U5636 (N_5636,N_5105,N_5240);
xor U5637 (N_5637,N_5029,N_5122);
nand U5638 (N_5638,N_5323,N_5249);
xor U5639 (N_5639,N_5274,N_5360);
nand U5640 (N_5640,N_5063,N_5438);
nor U5641 (N_5641,N_5346,N_5183);
nor U5642 (N_5642,N_5207,N_5246);
nor U5643 (N_5643,N_5049,N_5308);
xnor U5644 (N_5644,N_5439,N_5392);
and U5645 (N_5645,N_5325,N_5283);
or U5646 (N_5646,N_5127,N_5110);
nor U5647 (N_5647,N_5036,N_5180);
nand U5648 (N_5648,N_5256,N_5468);
and U5649 (N_5649,N_5374,N_5213);
nor U5650 (N_5650,N_5113,N_5437);
xnor U5651 (N_5651,N_5302,N_5290);
nand U5652 (N_5652,N_5255,N_5348);
nand U5653 (N_5653,N_5057,N_5426);
or U5654 (N_5654,N_5410,N_5490);
nor U5655 (N_5655,N_5229,N_5225);
nor U5656 (N_5656,N_5095,N_5338);
nand U5657 (N_5657,N_5212,N_5472);
or U5658 (N_5658,N_5237,N_5394);
and U5659 (N_5659,N_5317,N_5067);
nand U5660 (N_5660,N_5026,N_5333);
xor U5661 (N_5661,N_5420,N_5291);
nor U5662 (N_5662,N_5444,N_5239);
or U5663 (N_5663,N_5211,N_5330);
nand U5664 (N_5664,N_5210,N_5188);
nor U5665 (N_5665,N_5300,N_5130);
or U5666 (N_5666,N_5241,N_5093);
nand U5667 (N_5667,N_5406,N_5250);
and U5668 (N_5668,N_5305,N_5258);
and U5669 (N_5669,N_5447,N_5379);
and U5670 (N_5670,N_5156,N_5102);
nand U5671 (N_5671,N_5245,N_5381);
and U5672 (N_5672,N_5111,N_5286);
or U5673 (N_5673,N_5339,N_5247);
or U5674 (N_5674,N_5411,N_5396);
xnor U5675 (N_5675,N_5158,N_5203);
or U5676 (N_5676,N_5423,N_5018);
nor U5677 (N_5677,N_5041,N_5155);
and U5678 (N_5678,N_5090,N_5312);
or U5679 (N_5679,N_5040,N_5493);
or U5680 (N_5680,N_5301,N_5175);
and U5681 (N_5681,N_5165,N_5482);
or U5682 (N_5682,N_5466,N_5460);
nor U5683 (N_5683,N_5055,N_5077);
nor U5684 (N_5684,N_5136,N_5389);
and U5685 (N_5685,N_5065,N_5138);
xnor U5686 (N_5686,N_5143,N_5358);
and U5687 (N_5687,N_5056,N_5327);
nand U5688 (N_5688,N_5288,N_5008);
nand U5689 (N_5689,N_5380,N_5242);
nand U5690 (N_5690,N_5220,N_5137);
nand U5691 (N_5691,N_5104,N_5448);
and U5692 (N_5692,N_5487,N_5098);
or U5693 (N_5693,N_5078,N_5393);
nand U5694 (N_5694,N_5072,N_5269);
xor U5695 (N_5695,N_5119,N_5272);
xor U5696 (N_5696,N_5309,N_5033);
nand U5697 (N_5697,N_5015,N_5024);
xnor U5698 (N_5698,N_5163,N_5361);
nand U5699 (N_5699,N_5160,N_5094);
and U5700 (N_5700,N_5128,N_5386);
xnor U5701 (N_5701,N_5190,N_5038);
nor U5702 (N_5702,N_5473,N_5350);
or U5703 (N_5703,N_5371,N_5032);
nor U5704 (N_5704,N_5397,N_5071);
and U5705 (N_5705,N_5017,N_5085);
nand U5706 (N_5706,N_5307,N_5005);
and U5707 (N_5707,N_5135,N_5431);
or U5708 (N_5708,N_5101,N_5084);
or U5709 (N_5709,N_5376,N_5200);
nor U5710 (N_5710,N_5052,N_5218);
and U5711 (N_5711,N_5148,N_5173);
nand U5712 (N_5712,N_5144,N_5383);
nand U5713 (N_5713,N_5083,N_5316);
or U5714 (N_5714,N_5060,N_5168);
nor U5715 (N_5715,N_5068,N_5264);
and U5716 (N_5716,N_5470,N_5362);
nor U5717 (N_5717,N_5109,N_5044);
nor U5718 (N_5718,N_5372,N_5169);
nand U5719 (N_5719,N_5369,N_5134);
and U5720 (N_5720,N_5484,N_5391);
nor U5721 (N_5721,N_5224,N_5051);
or U5722 (N_5722,N_5257,N_5115);
nand U5723 (N_5723,N_5152,N_5092);
and U5724 (N_5724,N_5434,N_5282);
nand U5725 (N_5725,N_5116,N_5133);
nand U5726 (N_5726,N_5012,N_5217);
or U5727 (N_5727,N_5176,N_5461);
xnor U5728 (N_5728,N_5189,N_5088);
xnor U5729 (N_5729,N_5452,N_5489);
and U5730 (N_5730,N_5407,N_5492);
or U5731 (N_5731,N_5352,N_5076);
and U5732 (N_5732,N_5467,N_5476);
nand U5733 (N_5733,N_5355,N_5027);
or U5734 (N_5734,N_5446,N_5343);
nor U5735 (N_5735,N_5442,N_5280);
and U5736 (N_5736,N_5342,N_5132);
or U5737 (N_5737,N_5315,N_5477);
or U5738 (N_5738,N_5366,N_5419);
or U5739 (N_5739,N_5377,N_5382);
nor U5740 (N_5740,N_5412,N_5194);
or U5741 (N_5741,N_5276,N_5403);
and U5742 (N_5742,N_5080,N_5365);
or U5743 (N_5743,N_5014,N_5162);
and U5744 (N_5744,N_5289,N_5337);
nand U5745 (N_5745,N_5455,N_5089);
nand U5746 (N_5746,N_5087,N_5414);
nand U5747 (N_5747,N_5351,N_5216);
nand U5748 (N_5748,N_5400,N_5402);
and U5749 (N_5749,N_5260,N_5002);
or U5750 (N_5750,N_5478,N_5067);
nand U5751 (N_5751,N_5224,N_5048);
nor U5752 (N_5752,N_5009,N_5332);
and U5753 (N_5753,N_5253,N_5260);
nor U5754 (N_5754,N_5178,N_5258);
or U5755 (N_5755,N_5050,N_5435);
nand U5756 (N_5756,N_5389,N_5191);
nor U5757 (N_5757,N_5366,N_5256);
or U5758 (N_5758,N_5180,N_5384);
nor U5759 (N_5759,N_5380,N_5196);
nor U5760 (N_5760,N_5452,N_5273);
nand U5761 (N_5761,N_5250,N_5447);
nor U5762 (N_5762,N_5499,N_5085);
nand U5763 (N_5763,N_5190,N_5095);
or U5764 (N_5764,N_5411,N_5433);
nand U5765 (N_5765,N_5372,N_5468);
nor U5766 (N_5766,N_5046,N_5139);
and U5767 (N_5767,N_5293,N_5147);
nand U5768 (N_5768,N_5105,N_5027);
or U5769 (N_5769,N_5112,N_5315);
nor U5770 (N_5770,N_5222,N_5053);
or U5771 (N_5771,N_5176,N_5434);
nand U5772 (N_5772,N_5025,N_5114);
xor U5773 (N_5773,N_5099,N_5355);
nor U5774 (N_5774,N_5389,N_5309);
or U5775 (N_5775,N_5090,N_5005);
or U5776 (N_5776,N_5041,N_5251);
and U5777 (N_5777,N_5025,N_5173);
xnor U5778 (N_5778,N_5434,N_5349);
nand U5779 (N_5779,N_5000,N_5462);
nor U5780 (N_5780,N_5478,N_5453);
or U5781 (N_5781,N_5134,N_5059);
and U5782 (N_5782,N_5422,N_5285);
xnor U5783 (N_5783,N_5316,N_5068);
nor U5784 (N_5784,N_5043,N_5447);
nor U5785 (N_5785,N_5346,N_5461);
or U5786 (N_5786,N_5287,N_5274);
or U5787 (N_5787,N_5047,N_5161);
or U5788 (N_5788,N_5454,N_5049);
and U5789 (N_5789,N_5139,N_5205);
nand U5790 (N_5790,N_5060,N_5405);
or U5791 (N_5791,N_5332,N_5417);
or U5792 (N_5792,N_5408,N_5069);
xor U5793 (N_5793,N_5344,N_5120);
nor U5794 (N_5794,N_5352,N_5362);
nor U5795 (N_5795,N_5362,N_5037);
or U5796 (N_5796,N_5030,N_5333);
nand U5797 (N_5797,N_5418,N_5048);
nand U5798 (N_5798,N_5352,N_5097);
and U5799 (N_5799,N_5097,N_5439);
or U5800 (N_5800,N_5101,N_5479);
nor U5801 (N_5801,N_5224,N_5286);
nand U5802 (N_5802,N_5218,N_5032);
nor U5803 (N_5803,N_5416,N_5239);
and U5804 (N_5804,N_5238,N_5317);
xnor U5805 (N_5805,N_5446,N_5235);
nor U5806 (N_5806,N_5299,N_5003);
and U5807 (N_5807,N_5405,N_5019);
or U5808 (N_5808,N_5429,N_5150);
nor U5809 (N_5809,N_5200,N_5024);
nor U5810 (N_5810,N_5437,N_5420);
nand U5811 (N_5811,N_5004,N_5281);
and U5812 (N_5812,N_5177,N_5251);
nand U5813 (N_5813,N_5132,N_5021);
or U5814 (N_5814,N_5057,N_5284);
xnor U5815 (N_5815,N_5140,N_5341);
and U5816 (N_5816,N_5462,N_5441);
nor U5817 (N_5817,N_5258,N_5401);
xnor U5818 (N_5818,N_5003,N_5061);
and U5819 (N_5819,N_5237,N_5336);
and U5820 (N_5820,N_5433,N_5076);
nor U5821 (N_5821,N_5056,N_5100);
nand U5822 (N_5822,N_5355,N_5452);
nand U5823 (N_5823,N_5237,N_5325);
and U5824 (N_5824,N_5101,N_5242);
xnor U5825 (N_5825,N_5465,N_5359);
nand U5826 (N_5826,N_5448,N_5161);
nor U5827 (N_5827,N_5432,N_5066);
or U5828 (N_5828,N_5339,N_5464);
nand U5829 (N_5829,N_5100,N_5362);
nor U5830 (N_5830,N_5022,N_5131);
or U5831 (N_5831,N_5072,N_5341);
xnor U5832 (N_5832,N_5304,N_5054);
xor U5833 (N_5833,N_5315,N_5365);
xor U5834 (N_5834,N_5016,N_5242);
and U5835 (N_5835,N_5108,N_5154);
nand U5836 (N_5836,N_5084,N_5385);
or U5837 (N_5837,N_5211,N_5255);
or U5838 (N_5838,N_5379,N_5025);
nor U5839 (N_5839,N_5274,N_5488);
or U5840 (N_5840,N_5091,N_5215);
and U5841 (N_5841,N_5198,N_5142);
or U5842 (N_5842,N_5064,N_5263);
and U5843 (N_5843,N_5035,N_5196);
nor U5844 (N_5844,N_5334,N_5303);
nand U5845 (N_5845,N_5389,N_5046);
and U5846 (N_5846,N_5427,N_5352);
nor U5847 (N_5847,N_5446,N_5282);
nand U5848 (N_5848,N_5250,N_5487);
or U5849 (N_5849,N_5074,N_5415);
nand U5850 (N_5850,N_5420,N_5346);
nor U5851 (N_5851,N_5275,N_5483);
and U5852 (N_5852,N_5242,N_5312);
or U5853 (N_5853,N_5432,N_5341);
and U5854 (N_5854,N_5138,N_5317);
nor U5855 (N_5855,N_5394,N_5151);
nand U5856 (N_5856,N_5151,N_5031);
and U5857 (N_5857,N_5449,N_5237);
and U5858 (N_5858,N_5426,N_5431);
and U5859 (N_5859,N_5309,N_5461);
nand U5860 (N_5860,N_5265,N_5150);
and U5861 (N_5861,N_5019,N_5127);
xnor U5862 (N_5862,N_5250,N_5404);
or U5863 (N_5863,N_5161,N_5116);
and U5864 (N_5864,N_5107,N_5262);
or U5865 (N_5865,N_5168,N_5316);
and U5866 (N_5866,N_5325,N_5402);
nand U5867 (N_5867,N_5393,N_5432);
and U5868 (N_5868,N_5255,N_5400);
or U5869 (N_5869,N_5336,N_5169);
and U5870 (N_5870,N_5104,N_5056);
nand U5871 (N_5871,N_5484,N_5049);
and U5872 (N_5872,N_5336,N_5358);
and U5873 (N_5873,N_5194,N_5135);
or U5874 (N_5874,N_5440,N_5254);
nand U5875 (N_5875,N_5496,N_5458);
nor U5876 (N_5876,N_5442,N_5447);
xnor U5877 (N_5877,N_5277,N_5160);
nor U5878 (N_5878,N_5230,N_5179);
or U5879 (N_5879,N_5332,N_5218);
nand U5880 (N_5880,N_5269,N_5391);
or U5881 (N_5881,N_5200,N_5212);
or U5882 (N_5882,N_5268,N_5156);
nand U5883 (N_5883,N_5139,N_5426);
xor U5884 (N_5884,N_5445,N_5199);
and U5885 (N_5885,N_5464,N_5390);
nand U5886 (N_5886,N_5461,N_5037);
xnor U5887 (N_5887,N_5482,N_5002);
nand U5888 (N_5888,N_5110,N_5118);
and U5889 (N_5889,N_5280,N_5031);
nor U5890 (N_5890,N_5272,N_5336);
and U5891 (N_5891,N_5375,N_5248);
and U5892 (N_5892,N_5055,N_5323);
and U5893 (N_5893,N_5162,N_5287);
or U5894 (N_5894,N_5362,N_5355);
or U5895 (N_5895,N_5434,N_5188);
nand U5896 (N_5896,N_5324,N_5161);
and U5897 (N_5897,N_5393,N_5157);
nand U5898 (N_5898,N_5249,N_5105);
nand U5899 (N_5899,N_5410,N_5012);
nor U5900 (N_5900,N_5250,N_5378);
and U5901 (N_5901,N_5262,N_5334);
or U5902 (N_5902,N_5326,N_5241);
nor U5903 (N_5903,N_5426,N_5045);
or U5904 (N_5904,N_5304,N_5148);
or U5905 (N_5905,N_5276,N_5495);
and U5906 (N_5906,N_5462,N_5076);
nand U5907 (N_5907,N_5005,N_5096);
xor U5908 (N_5908,N_5062,N_5233);
nor U5909 (N_5909,N_5461,N_5163);
nand U5910 (N_5910,N_5439,N_5456);
nor U5911 (N_5911,N_5487,N_5351);
or U5912 (N_5912,N_5274,N_5459);
and U5913 (N_5913,N_5192,N_5251);
or U5914 (N_5914,N_5192,N_5173);
nand U5915 (N_5915,N_5230,N_5052);
nand U5916 (N_5916,N_5377,N_5091);
or U5917 (N_5917,N_5317,N_5009);
or U5918 (N_5918,N_5450,N_5224);
or U5919 (N_5919,N_5493,N_5016);
or U5920 (N_5920,N_5389,N_5217);
and U5921 (N_5921,N_5112,N_5395);
xnor U5922 (N_5922,N_5400,N_5241);
xnor U5923 (N_5923,N_5208,N_5004);
or U5924 (N_5924,N_5313,N_5360);
and U5925 (N_5925,N_5238,N_5262);
nor U5926 (N_5926,N_5075,N_5309);
nand U5927 (N_5927,N_5132,N_5217);
and U5928 (N_5928,N_5319,N_5490);
nor U5929 (N_5929,N_5112,N_5378);
xor U5930 (N_5930,N_5197,N_5064);
or U5931 (N_5931,N_5389,N_5037);
xor U5932 (N_5932,N_5158,N_5206);
or U5933 (N_5933,N_5256,N_5194);
and U5934 (N_5934,N_5225,N_5489);
nor U5935 (N_5935,N_5314,N_5398);
nand U5936 (N_5936,N_5286,N_5484);
nor U5937 (N_5937,N_5289,N_5101);
or U5938 (N_5938,N_5007,N_5027);
or U5939 (N_5939,N_5210,N_5119);
or U5940 (N_5940,N_5249,N_5224);
and U5941 (N_5941,N_5209,N_5068);
or U5942 (N_5942,N_5252,N_5112);
or U5943 (N_5943,N_5367,N_5142);
nand U5944 (N_5944,N_5122,N_5226);
or U5945 (N_5945,N_5009,N_5377);
and U5946 (N_5946,N_5083,N_5304);
and U5947 (N_5947,N_5456,N_5257);
xor U5948 (N_5948,N_5423,N_5137);
and U5949 (N_5949,N_5037,N_5349);
nor U5950 (N_5950,N_5391,N_5436);
nand U5951 (N_5951,N_5162,N_5161);
nand U5952 (N_5952,N_5484,N_5059);
nand U5953 (N_5953,N_5342,N_5110);
xor U5954 (N_5954,N_5251,N_5314);
xor U5955 (N_5955,N_5053,N_5018);
xor U5956 (N_5956,N_5288,N_5039);
nand U5957 (N_5957,N_5464,N_5124);
and U5958 (N_5958,N_5028,N_5456);
and U5959 (N_5959,N_5172,N_5454);
nand U5960 (N_5960,N_5098,N_5140);
nor U5961 (N_5961,N_5477,N_5336);
nor U5962 (N_5962,N_5203,N_5161);
nand U5963 (N_5963,N_5452,N_5221);
xnor U5964 (N_5964,N_5401,N_5333);
nor U5965 (N_5965,N_5462,N_5483);
or U5966 (N_5966,N_5167,N_5446);
and U5967 (N_5967,N_5094,N_5355);
or U5968 (N_5968,N_5255,N_5043);
nand U5969 (N_5969,N_5308,N_5309);
nor U5970 (N_5970,N_5027,N_5421);
or U5971 (N_5971,N_5415,N_5148);
xor U5972 (N_5972,N_5116,N_5400);
nand U5973 (N_5973,N_5304,N_5293);
and U5974 (N_5974,N_5284,N_5154);
or U5975 (N_5975,N_5155,N_5146);
or U5976 (N_5976,N_5380,N_5132);
nand U5977 (N_5977,N_5215,N_5465);
nor U5978 (N_5978,N_5043,N_5163);
nor U5979 (N_5979,N_5304,N_5221);
nand U5980 (N_5980,N_5008,N_5304);
nand U5981 (N_5981,N_5008,N_5387);
and U5982 (N_5982,N_5408,N_5476);
or U5983 (N_5983,N_5173,N_5215);
xnor U5984 (N_5984,N_5352,N_5411);
nand U5985 (N_5985,N_5119,N_5121);
or U5986 (N_5986,N_5371,N_5261);
nor U5987 (N_5987,N_5102,N_5013);
nor U5988 (N_5988,N_5181,N_5263);
nand U5989 (N_5989,N_5022,N_5399);
or U5990 (N_5990,N_5214,N_5366);
xor U5991 (N_5991,N_5314,N_5473);
nand U5992 (N_5992,N_5003,N_5039);
xor U5993 (N_5993,N_5214,N_5428);
nor U5994 (N_5994,N_5477,N_5208);
nor U5995 (N_5995,N_5319,N_5288);
nand U5996 (N_5996,N_5061,N_5425);
and U5997 (N_5997,N_5377,N_5084);
or U5998 (N_5998,N_5275,N_5005);
or U5999 (N_5999,N_5020,N_5462);
or U6000 (N_6000,N_5932,N_5955);
nor U6001 (N_6001,N_5541,N_5858);
and U6002 (N_6002,N_5765,N_5997);
nor U6003 (N_6003,N_5806,N_5700);
and U6004 (N_6004,N_5526,N_5937);
nor U6005 (N_6005,N_5785,N_5877);
nor U6006 (N_6006,N_5843,N_5857);
or U6007 (N_6007,N_5738,N_5945);
nor U6008 (N_6008,N_5555,N_5989);
or U6009 (N_6009,N_5626,N_5925);
nor U6010 (N_6010,N_5698,N_5732);
and U6011 (N_6011,N_5856,N_5661);
nand U6012 (N_6012,N_5602,N_5846);
nand U6013 (N_6013,N_5531,N_5999);
nor U6014 (N_6014,N_5548,N_5904);
and U6015 (N_6015,N_5728,N_5560);
and U6016 (N_6016,N_5618,N_5998);
nand U6017 (N_6017,N_5851,N_5978);
nand U6018 (N_6018,N_5687,N_5537);
and U6019 (N_6019,N_5591,N_5990);
or U6020 (N_6020,N_5791,N_5612);
nand U6021 (N_6021,N_5686,N_5762);
nand U6022 (N_6022,N_5772,N_5505);
or U6023 (N_6023,N_5640,N_5819);
nand U6024 (N_6024,N_5500,N_5717);
and U6025 (N_6025,N_5939,N_5809);
nand U6026 (N_6026,N_5615,N_5694);
or U6027 (N_6027,N_5664,N_5563);
or U6028 (N_6028,N_5834,N_5679);
and U6029 (N_6029,N_5893,N_5701);
and U6030 (N_6030,N_5572,N_5807);
and U6031 (N_6031,N_5777,N_5524);
xnor U6032 (N_6032,N_5817,N_5745);
or U6033 (N_6033,N_5642,N_5523);
nor U6034 (N_6034,N_5684,N_5677);
nor U6035 (N_6035,N_5909,N_5719);
nand U6036 (N_6036,N_5780,N_5658);
nor U6037 (N_6037,N_5993,N_5900);
or U6038 (N_6038,N_5963,N_5656);
nor U6039 (N_6039,N_5603,N_5530);
or U6040 (N_6040,N_5597,N_5695);
or U6041 (N_6041,N_5580,N_5634);
nand U6042 (N_6042,N_5767,N_5914);
nand U6043 (N_6043,N_5960,N_5730);
nand U6044 (N_6044,N_5586,N_5923);
nor U6045 (N_6045,N_5986,N_5880);
or U6046 (N_6046,N_5666,N_5828);
or U6047 (N_6047,N_5693,N_5912);
nand U6048 (N_6048,N_5619,N_5891);
nor U6049 (N_6049,N_5561,N_5910);
nor U6050 (N_6050,N_5558,N_5575);
nand U6051 (N_6051,N_5752,N_5611);
or U6052 (N_6052,N_5798,N_5559);
and U6053 (N_6053,N_5567,N_5689);
and U6054 (N_6054,N_5742,N_5646);
or U6055 (N_6055,N_5840,N_5797);
and U6056 (N_6056,N_5959,N_5546);
or U6057 (N_6057,N_5595,N_5926);
nor U6058 (N_6058,N_5502,N_5643);
nand U6059 (N_6059,N_5660,N_5746);
nor U6060 (N_6060,N_5631,N_5763);
xnor U6061 (N_6061,N_5885,N_5953);
or U6062 (N_6062,N_5744,N_5985);
or U6063 (N_6063,N_5655,N_5758);
nand U6064 (N_6064,N_5929,N_5831);
nand U6065 (N_6065,N_5715,N_5731);
and U6066 (N_6066,N_5652,N_5933);
nor U6067 (N_6067,N_5621,N_5753);
and U6068 (N_6068,N_5610,N_5570);
or U6069 (N_6069,N_5888,N_5915);
or U6070 (N_6070,N_5599,N_5883);
or U6071 (N_6071,N_5871,N_5971);
or U6072 (N_6072,N_5855,N_5995);
xnor U6073 (N_6073,N_5924,N_5839);
nand U6074 (N_6074,N_5515,N_5680);
nor U6075 (N_6075,N_5585,N_5829);
xnor U6076 (N_6076,N_5952,N_5635);
nand U6077 (N_6077,N_5670,N_5562);
nor U6078 (N_6078,N_5943,N_5950);
and U6079 (N_6079,N_5946,N_5659);
nand U6080 (N_6080,N_5847,N_5941);
and U6081 (N_6081,N_5761,N_5632);
nor U6082 (N_6082,N_5508,N_5882);
nand U6083 (N_6083,N_5514,N_5906);
nand U6084 (N_6084,N_5868,N_5630);
xnor U6085 (N_6085,N_5581,N_5844);
nand U6086 (N_6086,N_5557,N_5781);
xor U6087 (N_6087,N_5638,N_5723);
nand U6088 (N_6088,N_5981,N_5633);
or U6089 (N_6089,N_5543,N_5651);
nand U6090 (N_6090,N_5872,N_5734);
nor U6091 (N_6091,N_5881,N_5759);
and U6092 (N_6092,N_5574,N_5783);
or U6093 (N_6093,N_5890,N_5653);
nor U6094 (N_6094,N_5850,N_5928);
xnor U6095 (N_6095,N_5962,N_5671);
nand U6096 (N_6096,N_5907,N_5566);
and U6097 (N_6097,N_5968,N_5613);
or U6098 (N_6098,N_5875,N_5866);
or U6099 (N_6099,N_5848,N_5965);
xnor U6100 (N_6100,N_5992,N_5678);
nand U6101 (N_6101,N_5617,N_5533);
nand U6102 (N_6102,N_5803,N_5813);
nor U6103 (N_6103,N_5628,N_5725);
nor U6104 (N_6104,N_5908,N_5865);
and U6105 (N_6105,N_5886,N_5788);
and U6106 (N_6106,N_5710,N_5535);
nand U6107 (N_6107,N_5683,N_5836);
xnor U6108 (N_6108,N_5782,N_5564);
nor U6109 (N_6109,N_5573,N_5709);
nor U6110 (N_6110,N_5938,N_5596);
nor U6111 (N_6111,N_5905,N_5808);
and U6112 (N_6112,N_5930,N_5849);
nor U6113 (N_6113,N_5716,N_5811);
nand U6114 (N_6114,N_5947,N_5810);
or U6115 (N_6115,N_5690,N_5571);
nand U6116 (N_6116,N_5793,N_5815);
nand U6117 (N_6117,N_5973,N_5835);
nor U6118 (N_6118,N_5936,N_5956);
xnor U6119 (N_6119,N_5902,N_5521);
nand U6120 (N_6120,N_5665,N_5601);
or U6121 (N_6121,N_5837,N_5688);
nand U6122 (N_6122,N_5887,N_5896);
or U6123 (N_6123,N_5587,N_5708);
and U6124 (N_6124,N_5736,N_5727);
nand U6125 (N_6125,N_5940,N_5650);
xnor U6126 (N_6126,N_5534,N_5739);
nor U6127 (N_6127,N_5920,N_5894);
nand U6128 (N_6128,N_5954,N_5787);
nand U6129 (N_6129,N_5721,N_5553);
or U6130 (N_6130,N_5697,N_5802);
or U6131 (N_6131,N_5771,N_5876);
or U6132 (N_6132,N_5584,N_5672);
or U6133 (N_6133,N_5980,N_5545);
nand U6134 (N_6134,N_5794,N_5796);
nor U6135 (N_6135,N_5784,N_5507);
nand U6136 (N_6136,N_5822,N_5898);
or U6137 (N_6137,N_5773,N_5676);
nand U6138 (N_6138,N_5801,N_5862);
nand U6139 (N_6139,N_5977,N_5895);
nor U6140 (N_6140,N_5516,N_5692);
and U6141 (N_6141,N_5504,N_5942);
or U6142 (N_6142,N_5712,N_5713);
or U6143 (N_6143,N_5616,N_5774);
and U6144 (N_6144,N_5565,N_5639);
or U6145 (N_6145,N_5852,N_5961);
or U6146 (N_6146,N_5576,N_5826);
or U6147 (N_6147,N_5931,N_5593);
or U6148 (N_6148,N_5779,N_5503);
nor U6149 (N_6149,N_5623,N_5922);
xnor U6150 (N_6150,N_5550,N_5824);
nand U6151 (N_6151,N_5705,N_5812);
nor U6152 (N_6152,N_5799,N_5751);
or U6153 (N_6153,N_5927,N_5854);
xor U6154 (N_6154,N_5789,N_5598);
nor U6155 (N_6155,N_5892,N_5805);
and U6156 (N_6156,N_5870,N_5590);
and U6157 (N_6157,N_5766,N_5832);
nor U6158 (N_6158,N_5790,N_5775);
and U6159 (N_6159,N_5726,N_5889);
and U6160 (N_6160,N_5919,N_5629);
nor U6161 (N_6161,N_5704,N_5921);
or U6162 (N_6162,N_5913,N_5528);
nor U6163 (N_6163,N_5583,N_5951);
or U6164 (N_6164,N_5525,N_5673);
and U6165 (N_6165,N_5662,N_5833);
xnor U6166 (N_6166,N_5976,N_5722);
and U6167 (N_6167,N_5879,N_5668);
nor U6168 (N_6168,N_5750,N_5800);
xor U6169 (N_6169,N_5568,N_5991);
and U6170 (N_6170,N_5510,N_5869);
or U6171 (N_6171,N_5996,N_5768);
nand U6172 (N_6172,N_5506,N_5624);
nand U6173 (N_6173,N_5641,N_5703);
or U6174 (N_6174,N_5600,N_5608);
nor U6175 (N_6175,N_5970,N_5756);
nand U6176 (N_6176,N_5592,N_5748);
or U6177 (N_6177,N_5527,N_5518);
or U6178 (N_6178,N_5884,N_5972);
nand U6179 (N_6179,N_5737,N_5609);
and U6180 (N_6180,N_5823,N_5522);
nand U6181 (N_6181,N_5792,N_5982);
or U6182 (N_6182,N_5691,N_5669);
and U6183 (N_6183,N_5589,N_5682);
nand U6184 (N_6184,N_5720,N_5544);
or U6185 (N_6185,N_5821,N_5594);
and U6186 (N_6186,N_5604,N_5983);
nor U6187 (N_6187,N_5724,N_5577);
nand U6188 (N_6188,N_5873,N_5964);
nor U6189 (N_6189,N_5867,N_5649);
nor U6190 (N_6190,N_5675,N_5606);
nor U6191 (N_6191,N_5949,N_5974);
nor U6192 (N_6192,N_5786,N_5764);
nand U6193 (N_6193,N_5743,N_5899);
and U6194 (N_6194,N_5536,N_5863);
nand U6195 (N_6195,N_5979,N_5778);
nand U6196 (N_6196,N_5551,N_5944);
nand U6197 (N_6197,N_5707,N_5532);
xor U6198 (N_6198,N_5674,N_5511);
or U6199 (N_6199,N_5554,N_5818);
or U6200 (N_6200,N_5864,N_5859);
nand U6201 (N_6201,N_5816,N_5733);
xnor U6202 (N_6202,N_5814,N_5654);
or U6203 (N_6203,N_5770,N_5582);
nor U6204 (N_6204,N_5520,N_5696);
nor U6205 (N_6205,N_5718,N_5699);
and U6206 (N_6206,N_5841,N_5614);
nor U6207 (N_6207,N_5512,N_5769);
nor U6208 (N_6208,N_5637,N_5605);
and U6209 (N_6209,N_5827,N_5776);
nor U6210 (N_6210,N_5644,N_5509);
or U6211 (N_6211,N_5754,N_5711);
nand U6212 (N_6212,N_5513,N_5579);
nand U6213 (N_6213,N_5934,N_5625);
nor U6214 (N_6214,N_5622,N_5842);
nand U6215 (N_6215,N_5911,N_5917);
xnor U6216 (N_6216,N_5607,N_5681);
nand U6217 (N_6217,N_5757,N_5918);
and U6218 (N_6218,N_5588,N_5663);
nor U6219 (N_6219,N_5552,N_5760);
and U6220 (N_6220,N_5667,N_5547);
or U6221 (N_6221,N_5549,N_5648);
nand U6222 (N_6222,N_5702,N_5519);
nor U6223 (N_6223,N_5966,N_5517);
and U6224 (N_6224,N_5749,N_5501);
nand U6225 (N_6225,N_5948,N_5878);
and U6226 (N_6226,N_5657,N_5825);
and U6227 (N_6227,N_5755,N_5556);
nand U6228 (N_6228,N_5706,N_5569);
nor U6229 (N_6229,N_5935,N_5957);
nor U6230 (N_6230,N_5861,N_5838);
nand U6231 (N_6231,N_5542,N_5685);
xnor U6232 (N_6232,N_5795,N_5860);
or U6233 (N_6233,N_5897,N_5747);
xnor U6234 (N_6234,N_5539,N_5830);
and U6235 (N_6235,N_5804,N_5538);
or U6236 (N_6236,N_5820,N_5903);
or U6237 (N_6237,N_5578,N_5916);
nor U6238 (N_6238,N_5741,N_5969);
xor U6239 (N_6239,N_5845,N_5729);
and U6240 (N_6240,N_5987,N_5975);
or U6241 (N_6241,N_5988,N_5645);
and U6242 (N_6242,N_5984,N_5994);
and U6243 (N_6243,N_5647,N_5529);
and U6244 (N_6244,N_5735,N_5627);
nand U6245 (N_6245,N_5714,N_5620);
and U6246 (N_6246,N_5540,N_5740);
xnor U6247 (N_6247,N_5636,N_5853);
or U6248 (N_6248,N_5874,N_5901);
nand U6249 (N_6249,N_5967,N_5958);
and U6250 (N_6250,N_5880,N_5833);
and U6251 (N_6251,N_5768,N_5607);
xnor U6252 (N_6252,N_5892,N_5944);
or U6253 (N_6253,N_5525,N_5748);
or U6254 (N_6254,N_5636,N_5517);
and U6255 (N_6255,N_5910,N_5598);
and U6256 (N_6256,N_5967,N_5813);
or U6257 (N_6257,N_5909,N_5969);
or U6258 (N_6258,N_5623,N_5912);
nand U6259 (N_6259,N_5528,N_5650);
and U6260 (N_6260,N_5501,N_5877);
nand U6261 (N_6261,N_5968,N_5537);
and U6262 (N_6262,N_5899,N_5727);
nor U6263 (N_6263,N_5626,N_5883);
nor U6264 (N_6264,N_5538,N_5641);
and U6265 (N_6265,N_5633,N_5747);
xnor U6266 (N_6266,N_5702,N_5957);
and U6267 (N_6267,N_5957,N_5605);
and U6268 (N_6268,N_5819,N_5990);
and U6269 (N_6269,N_5983,N_5832);
or U6270 (N_6270,N_5566,N_5999);
xnor U6271 (N_6271,N_5532,N_5870);
and U6272 (N_6272,N_5884,N_5625);
and U6273 (N_6273,N_5525,N_5937);
and U6274 (N_6274,N_5676,N_5663);
nand U6275 (N_6275,N_5826,N_5961);
or U6276 (N_6276,N_5725,N_5564);
nand U6277 (N_6277,N_5905,N_5525);
or U6278 (N_6278,N_5900,N_5806);
nand U6279 (N_6279,N_5595,N_5932);
nor U6280 (N_6280,N_5893,N_5612);
nor U6281 (N_6281,N_5646,N_5912);
nor U6282 (N_6282,N_5561,N_5898);
and U6283 (N_6283,N_5900,N_5516);
nand U6284 (N_6284,N_5576,N_5725);
and U6285 (N_6285,N_5964,N_5659);
or U6286 (N_6286,N_5684,N_5554);
nand U6287 (N_6287,N_5753,N_5636);
nor U6288 (N_6288,N_5828,N_5525);
xor U6289 (N_6289,N_5721,N_5802);
and U6290 (N_6290,N_5867,N_5781);
xnor U6291 (N_6291,N_5654,N_5794);
and U6292 (N_6292,N_5763,N_5840);
nand U6293 (N_6293,N_5576,N_5957);
nand U6294 (N_6294,N_5527,N_5703);
xor U6295 (N_6295,N_5981,N_5678);
or U6296 (N_6296,N_5712,N_5626);
nand U6297 (N_6297,N_5742,N_5544);
and U6298 (N_6298,N_5955,N_5693);
or U6299 (N_6299,N_5694,N_5752);
or U6300 (N_6300,N_5612,N_5829);
nand U6301 (N_6301,N_5507,N_5707);
nand U6302 (N_6302,N_5650,N_5928);
nand U6303 (N_6303,N_5521,N_5538);
or U6304 (N_6304,N_5663,N_5503);
and U6305 (N_6305,N_5942,N_5522);
and U6306 (N_6306,N_5547,N_5622);
nand U6307 (N_6307,N_5602,N_5818);
nor U6308 (N_6308,N_5786,N_5796);
nor U6309 (N_6309,N_5831,N_5756);
and U6310 (N_6310,N_5711,N_5894);
nor U6311 (N_6311,N_5750,N_5627);
nand U6312 (N_6312,N_5525,N_5809);
nand U6313 (N_6313,N_5561,N_5685);
nor U6314 (N_6314,N_5698,N_5679);
nand U6315 (N_6315,N_5636,N_5709);
and U6316 (N_6316,N_5891,N_5763);
and U6317 (N_6317,N_5686,N_5775);
or U6318 (N_6318,N_5925,N_5814);
and U6319 (N_6319,N_5946,N_5976);
nand U6320 (N_6320,N_5624,N_5851);
nor U6321 (N_6321,N_5590,N_5731);
and U6322 (N_6322,N_5834,N_5672);
nor U6323 (N_6323,N_5550,N_5858);
nor U6324 (N_6324,N_5580,N_5696);
xor U6325 (N_6325,N_5700,N_5585);
and U6326 (N_6326,N_5526,N_5722);
nand U6327 (N_6327,N_5783,N_5593);
nor U6328 (N_6328,N_5946,N_5601);
nand U6329 (N_6329,N_5513,N_5835);
xor U6330 (N_6330,N_5669,N_5519);
or U6331 (N_6331,N_5573,N_5707);
nor U6332 (N_6332,N_5819,N_5863);
nand U6333 (N_6333,N_5840,N_5890);
and U6334 (N_6334,N_5917,N_5932);
nand U6335 (N_6335,N_5990,N_5725);
nor U6336 (N_6336,N_5971,N_5783);
and U6337 (N_6337,N_5595,N_5940);
and U6338 (N_6338,N_5536,N_5817);
nand U6339 (N_6339,N_5945,N_5917);
nor U6340 (N_6340,N_5698,N_5914);
and U6341 (N_6341,N_5583,N_5946);
nand U6342 (N_6342,N_5586,N_5948);
xnor U6343 (N_6343,N_5901,N_5745);
and U6344 (N_6344,N_5610,N_5802);
xnor U6345 (N_6345,N_5923,N_5899);
nand U6346 (N_6346,N_5570,N_5916);
or U6347 (N_6347,N_5543,N_5994);
or U6348 (N_6348,N_5640,N_5846);
nor U6349 (N_6349,N_5500,N_5674);
xor U6350 (N_6350,N_5992,N_5764);
or U6351 (N_6351,N_5622,N_5557);
or U6352 (N_6352,N_5607,N_5591);
xor U6353 (N_6353,N_5637,N_5554);
xor U6354 (N_6354,N_5914,N_5614);
nand U6355 (N_6355,N_5853,N_5623);
or U6356 (N_6356,N_5796,N_5976);
nand U6357 (N_6357,N_5576,N_5794);
nor U6358 (N_6358,N_5973,N_5870);
nor U6359 (N_6359,N_5850,N_5760);
xnor U6360 (N_6360,N_5689,N_5990);
or U6361 (N_6361,N_5774,N_5521);
nand U6362 (N_6362,N_5525,N_5644);
xor U6363 (N_6363,N_5672,N_5982);
and U6364 (N_6364,N_5652,N_5876);
nor U6365 (N_6365,N_5857,N_5676);
nor U6366 (N_6366,N_5854,N_5838);
nand U6367 (N_6367,N_5769,N_5704);
xor U6368 (N_6368,N_5871,N_5669);
and U6369 (N_6369,N_5811,N_5651);
and U6370 (N_6370,N_5965,N_5798);
or U6371 (N_6371,N_5586,N_5951);
and U6372 (N_6372,N_5651,N_5974);
and U6373 (N_6373,N_5597,N_5675);
nand U6374 (N_6374,N_5877,N_5870);
and U6375 (N_6375,N_5867,N_5594);
and U6376 (N_6376,N_5542,N_5813);
and U6377 (N_6377,N_5884,N_5504);
nor U6378 (N_6378,N_5944,N_5813);
nand U6379 (N_6379,N_5676,N_5788);
nand U6380 (N_6380,N_5556,N_5658);
and U6381 (N_6381,N_5930,N_5711);
xnor U6382 (N_6382,N_5850,N_5877);
and U6383 (N_6383,N_5604,N_5958);
nand U6384 (N_6384,N_5970,N_5728);
nor U6385 (N_6385,N_5848,N_5515);
and U6386 (N_6386,N_5621,N_5657);
or U6387 (N_6387,N_5572,N_5684);
nor U6388 (N_6388,N_5766,N_5507);
nand U6389 (N_6389,N_5602,N_5668);
nor U6390 (N_6390,N_5992,N_5717);
or U6391 (N_6391,N_5747,N_5889);
or U6392 (N_6392,N_5837,N_5903);
xnor U6393 (N_6393,N_5722,N_5847);
or U6394 (N_6394,N_5757,N_5577);
nor U6395 (N_6395,N_5956,N_5764);
nor U6396 (N_6396,N_5901,N_5821);
nand U6397 (N_6397,N_5907,N_5758);
nand U6398 (N_6398,N_5997,N_5929);
nand U6399 (N_6399,N_5749,N_5703);
or U6400 (N_6400,N_5514,N_5984);
and U6401 (N_6401,N_5705,N_5721);
nor U6402 (N_6402,N_5555,N_5537);
xnor U6403 (N_6403,N_5566,N_5547);
or U6404 (N_6404,N_5780,N_5762);
and U6405 (N_6405,N_5935,N_5528);
or U6406 (N_6406,N_5573,N_5866);
nand U6407 (N_6407,N_5804,N_5806);
nor U6408 (N_6408,N_5591,N_5652);
xor U6409 (N_6409,N_5748,N_5912);
nand U6410 (N_6410,N_5644,N_5821);
nor U6411 (N_6411,N_5672,N_5842);
and U6412 (N_6412,N_5967,N_5505);
and U6413 (N_6413,N_5557,N_5979);
and U6414 (N_6414,N_5728,N_5828);
nand U6415 (N_6415,N_5505,N_5731);
nor U6416 (N_6416,N_5615,N_5757);
nand U6417 (N_6417,N_5906,N_5552);
nand U6418 (N_6418,N_5592,N_5656);
or U6419 (N_6419,N_5855,N_5940);
or U6420 (N_6420,N_5809,N_5544);
and U6421 (N_6421,N_5986,N_5783);
nor U6422 (N_6422,N_5540,N_5962);
or U6423 (N_6423,N_5503,N_5877);
xnor U6424 (N_6424,N_5699,N_5891);
and U6425 (N_6425,N_5765,N_5921);
nor U6426 (N_6426,N_5511,N_5597);
and U6427 (N_6427,N_5991,N_5760);
xnor U6428 (N_6428,N_5827,N_5550);
nor U6429 (N_6429,N_5642,N_5660);
xor U6430 (N_6430,N_5683,N_5779);
or U6431 (N_6431,N_5953,N_5563);
nand U6432 (N_6432,N_5618,N_5542);
and U6433 (N_6433,N_5681,N_5711);
nor U6434 (N_6434,N_5777,N_5928);
nand U6435 (N_6435,N_5912,N_5511);
nand U6436 (N_6436,N_5851,N_5901);
and U6437 (N_6437,N_5501,N_5766);
xor U6438 (N_6438,N_5624,N_5924);
and U6439 (N_6439,N_5856,N_5596);
nand U6440 (N_6440,N_5700,N_5543);
or U6441 (N_6441,N_5901,N_5565);
nor U6442 (N_6442,N_5773,N_5946);
nor U6443 (N_6443,N_5616,N_5710);
nand U6444 (N_6444,N_5709,N_5716);
and U6445 (N_6445,N_5769,N_5913);
nand U6446 (N_6446,N_5923,N_5794);
and U6447 (N_6447,N_5688,N_5702);
xnor U6448 (N_6448,N_5776,N_5985);
or U6449 (N_6449,N_5719,N_5915);
or U6450 (N_6450,N_5608,N_5790);
and U6451 (N_6451,N_5547,N_5540);
and U6452 (N_6452,N_5670,N_5985);
or U6453 (N_6453,N_5902,N_5665);
or U6454 (N_6454,N_5714,N_5979);
nand U6455 (N_6455,N_5643,N_5628);
xnor U6456 (N_6456,N_5545,N_5735);
or U6457 (N_6457,N_5556,N_5863);
nand U6458 (N_6458,N_5805,N_5528);
xor U6459 (N_6459,N_5949,N_5903);
nand U6460 (N_6460,N_5703,N_5570);
nor U6461 (N_6461,N_5867,N_5539);
or U6462 (N_6462,N_5674,N_5532);
nand U6463 (N_6463,N_5650,N_5817);
nand U6464 (N_6464,N_5694,N_5571);
nand U6465 (N_6465,N_5689,N_5690);
nand U6466 (N_6466,N_5740,N_5689);
nor U6467 (N_6467,N_5687,N_5560);
xor U6468 (N_6468,N_5886,N_5599);
nor U6469 (N_6469,N_5562,N_5595);
nand U6470 (N_6470,N_5616,N_5958);
or U6471 (N_6471,N_5862,N_5583);
nor U6472 (N_6472,N_5949,N_5628);
nor U6473 (N_6473,N_5968,N_5938);
and U6474 (N_6474,N_5979,N_5598);
nor U6475 (N_6475,N_5716,N_5526);
nor U6476 (N_6476,N_5857,N_5919);
and U6477 (N_6477,N_5626,N_5771);
and U6478 (N_6478,N_5820,N_5636);
and U6479 (N_6479,N_5722,N_5672);
nor U6480 (N_6480,N_5596,N_5822);
nand U6481 (N_6481,N_5894,N_5646);
or U6482 (N_6482,N_5842,N_5943);
nand U6483 (N_6483,N_5774,N_5554);
and U6484 (N_6484,N_5680,N_5960);
and U6485 (N_6485,N_5685,N_5597);
or U6486 (N_6486,N_5967,N_5829);
and U6487 (N_6487,N_5878,N_5873);
and U6488 (N_6488,N_5655,N_5669);
or U6489 (N_6489,N_5728,N_5789);
xnor U6490 (N_6490,N_5925,N_5873);
and U6491 (N_6491,N_5799,N_5698);
and U6492 (N_6492,N_5719,N_5794);
or U6493 (N_6493,N_5557,N_5767);
nor U6494 (N_6494,N_5714,N_5588);
or U6495 (N_6495,N_5961,N_5744);
nor U6496 (N_6496,N_5656,N_5661);
nand U6497 (N_6497,N_5530,N_5920);
nor U6498 (N_6498,N_5573,N_5520);
or U6499 (N_6499,N_5948,N_5981);
nand U6500 (N_6500,N_6081,N_6429);
nor U6501 (N_6501,N_6310,N_6440);
nand U6502 (N_6502,N_6161,N_6162);
nand U6503 (N_6503,N_6441,N_6196);
nor U6504 (N_6504,N_6139,N_6017);
nor U6505 (N_6505,N_6490,N_6381);
and U6506 (N_6506,N_6221,N_6027);
nand U6507 (N_6507,N_6459,N_6167);
nand U6508 (N_6508,N_6028,N_6464);
and U6509 (N_6509,N_6222,N_6488);
and U6510 (N_6510,N_6389,N_6402);
or U6511 (N_6511,N_6304,N_6447);
or U6512 (N_6512,N_6187,N_6358);
xnor U6513 (N_6513,N_6226,N_6120);
nor U6514 (N_6514,N_6181,N_6386);
and U6515 (N_6515,N_6078,N_6307);
nand U6516 (N_6516,N_6416,N_6320);
and U6517 (N_6517,N_6036,N_6461);
nor U6518 (N_6518,N_6173,N_6007);
or U6519 (N_6519,N_6319,N_6029);
and U6520 (N_6520,N_6008,N_6018);
or U6521 (N_6521,N_6413,N_6475);
nand U6522 (N_6522,N_6457,N_6095);
nand U6523 (N_6523,N_6092,N_6335);
nand U6524 (N_6524,N_6483,N_6170);
and U6525 (N_6525,N_6052,N_6171);
or U6526 (N_6526,N_6494,N_6063);
nand U6527 (N_6527,N_6420,N_6444);
and U6528 (N_6528,N_6022,N_6409);
and U6529 (N_6529,N_6426,N_6435);
nor U6530 (N_6530,N_6012,N_6143);
or U6531 (N_6531,N_6131,N_6314);
and U6532 (N_6532,N_6214,N_6127);
nand U6533 (N_6533,N_6054,N_6013);
xnor U6534 (N_6534,N_6244,N_6313);
nor U6535 (N_6535,N_6371,N_6376);
nor U6536 (N_6536,N_6390,N_6000);
nor U6537 (N_6537,N_6168,N_6098);
xnor U6538 (N_6538,N_6086,N_6145);
and U6539 (N_6539,N_6303,N_6257);
or U6540 (N_6540,N_6034,N_6346);
or U6541 (N_6541,N_6469,N_6123);
nor U6542 (N_6542,N_6190,N_6116);
and U6543 (N_6543,N_6010,N_6020);
nand U6544 (N_6544,N_6067,N_6178);
and U6545 (N_6545,N_6436,N_6341);
and U6546 (N_6546,N_6014,N_6284);
nand U6547 (N_6547,N_6258,N_6198);
nand U6548 (N_6548,N_6419,N_6138);
nand U6549 (N_6549,N_6135,N_6043);
nand U6550 (N_6550,N_6427,N_6184);
nor U6551 (N_6551,N_6312,N_6249);
nand U6552 (N_6552,N_6180,N_6451);
nor U6553 (N_6553,N_6251,N_6431);
nand U6554 (N_6554,N_6348,N_6262);
and U6555 (N_6555,N_6481,N_6282);
and U6556 (N_6556,N_6388,N_6003);
or U6557 (N_6557,N_6468,N_6188);
or U6558 (N_6558,N_6033,N_6082);
or U6559 (N_6559,N_6405,N_6480);
nor U6560 (N_6560,N_6418,N_6422);
nand U6561 (N_6561,N_6204,N_6300);
or U6562 (N_6562,N_6492,N_6317);
nor U6563 (N_6563,N_6351,N_6298);
or U6564 (N_6564,N_6268,N_6212);
nand U6565 (N_6565,N_6292,N_6087);
or U6566 (N_6566,N_6477,N_6438);
and U6567 (N_6567,N_6215,N_6201);
nor U6568 (N_6568,N_6216,N_6159);
and U6569 (N_6569,N_6015,N_6295);
nand U6570 (N_6570,N_6446,N_6001);
nand U6571 (N_6571,N_6164,N_6125);
or U6572 (N_6572,N_6174,N_6232);
and U6573 (N_6573,N_6255,N_6278);
or U6574 (N_6574,N_6456,N_6247);
or U6575 (N_6575,N_6316,N_6263);
nand U6576 (N_6576,N_6177,N_6210);
and U6577 (N_6577,N_6336,N_6152);
nand U6578 (N_6578,N_6458,N_6073);
nand U6579 (N_6579,N_6434,N_6045);
or U6580 (N_6580,N_6193,N_6349);
or U6581 (N_6581,N_6285,N_6404);
nor U6582 (N_6582,N_6025,N_6023);
and U6583 (N_6583,N_6423,N_6071);
or U6584 (N_6584,N_6096,N_6110);
nand U6585 (N_6585,N_6396,N_6279);
nor U6586 (N_6586,N_6217,N_6403);
or U6587 (N_6587,N_6021,N_6175);
and U6588 (N_6588,N_6191,N_6286);
and U6589 (N_6589,N_6484,N_6172);
nand U6590 (N_6590,N_6373,N_6097);
or U6591 (N_6591,N_6118,N_6450);
and U6592 (N_6592,N_6084,N_6274);
or U6593 (N_6593,N_6267,N_6377);
nor U6594 (N_6594,N_6070,N_6189);
nor U6595 (N_6595,N_6315,N_6301);
nor U6596 (N_6596,N_6041,N_6364);
or U6597 (N_6597,N_6385,N_6103);
nand U6598 (N_6598,N_6410,N_6151);
and U6599 (N_6599,N_6337,N_6047);
or U6600 (N_6600,N_6383,N_6107);
nand U6601 (N_6601,N_6366,N_6155);
nor U6602 (N_6602,N_6424,N_6487);
xor U6603 (N_6603,N_6203,N_6100);
nor U6604 (N_6604,N_6032,N_6250);
nor U6605 (N_6605,N_6368,N_6328);
nand U6606 (N_6606,N_6037,N_6342);
nand U6607 (N_6607,N_6160,N_6259);
nor U6608 (N_6608,N_6064,N_6121);
nor U6609 (N_6609,N_6030,N_6365);
nor U6610 (N_6610,N_6239,N_6372);
or U6611 (N_6611,N_6290,N_6219);
nand U6612 (N_6612,N_6202,N_6088);
nand U6613 (N_6613,N_6115,N_6209);
or U6614 (N_6614,N_6367,N_6261);
nor U6615 (N_6615,N_6192,N_6142);
nor U6616 (N_6616,N_6331,N_6050);
or U6617 (N_6617,N_6399,N_6472);
or U6618 (N_6618,N_6004,N_6166);
nor U6619 (N_6619,N_6325,N_6207);
or U6620 (N_6620,N_6421,N_6387);
nand U6621 (N_6621,N_6147,N_6074);
and U6622 (N_6622,N_6197,N_6499);
or U6623 (N_6623,N_6374,N_6256);
nand U6624 (N_6624,N_6400,N_6350);
and U6625 (N_6625,N_6417,N_6306);
xor U6626 (N_6626,N_6061,N_6498);
nand U6627 (N_6627,N_6104,N_6114);
or U6628 (N_6628,N_6042,N_6153);
or U6629 (N_6629,N_6075,N_6449);
xor U6630 (N_6630,N_6370,N_6362);
or U6631 (N_6631,N_6452,N_6146);
nor U6632 (N_6632,N_6493,N_6384);
nand U6633 (N_6633,N_6165,N_6194);
nor U6634 (N_6634,N_6243,N_6056);
and U6635 (N_6635,N_6156,N_6357);
nor U6636 (N_6636,N_6225,N_6065);
and U6637 (N_6637,N_6218,N_6398);
nand U6638 (N_6638,N_6085,N_6124);
or U6639 (N_6639,N_6106,N_6462);
nor U6640 (N_6640,N_6133,N_6090);
xnor U6641 (N_6641,N_6158,N_6169);
and U6642 (N_6642,N_6471,N_6235);
nor U6643 (N_6643,N_6375,N_6051);
nor U6644 (N_6644,N_6111,N_6496);
nor U6645 (N_6645,N_6266,N_6199);
nand U6646 (N_6646,N_6411,N_6294);
nor U6647 (N_6647,N_6253,N_6289);
nand U6648 (N_6648,N_6011,N_6318);
nor U6649 (N_6649,N_6016,N_6269);
and U6650 (N_6650,N_6252,N_6430);
and U6651 (N_6651,N_6345,N_6476);
and U6652 (N_6652,N_6283,N_6068);
nor U6653 (N_6653,N_6254,N_6273);
nand U6654 (N_6654,N_6080,N_6059);
and U6655 (N_6655,N_6240,N_6465);
nand U6656 (N_6656,N_6182,N_6454);
nor U6657 (N_6657,N_6428,N_6058);
nor U6658 (N_6658,N_6136,N_6489);
or U6659 (N_6659,N_6048,N_6205);
nor U6660 (N_6660,N_6455,N_6122);
xnor U6661 (N_6661,N_6329,N_6270);
or U6662 (N_6662,N_6265,N_6150);
or U6663 (N_6663,N_6149,N_6333);
and U6664 (N_6664,N_6089,N_6291);
xnor U6665 (N_6665,N_6072,N_6211);
or U6666 (N_6666,N_6332,N_6006);
nor U6667 (N_6667,N_6439,N_6176);
and U6668 (N_6668,N_6393,N_6183);
and U6669 (N_6669,N_6397,N_6031);
and U6670 (N_6670,N_6060,N_6272);
nor U6671 (N_6671,N_6237,N_6354);
and U6672 (N_6672,N_6276,N_6236);
nand U6673 (N_6673,N_6361,N_6378);
or U6674 (N_6674,N_6395,N_6049);
and U6675 (N_6675,N_6356,N_6414);
nand U6676 (N_6676,N_6005,N_6343);
nand U6677 (N_6677,N_6412,N_6230);
or U6678 (N_6678,N_6287,N_6486);
or U6679 (N_6679,N_6264,N_6069);
nand U6680 (N_6680,N_6093,N_6140);
or U6681 (N_6681,N_6246,N_6478);
nor U6682 (N_6682,N_6026,N_6200);
or U6683 (N_6683,N_6208,N_6248);
or U6684 (N_6684,N_6280,N_6433);
nor U6685 (N_6685,N_6002,N_6297);
nand U6686 (N_6686,N_6079,N_6077);
or U6687 (N_6687,N_6293,N_6359);
nor U6688 (N_6688,N_6101,N_6445);
nor U6689 (N_6689,N_6392,N_6238);
nor U6690 (N_6690,N_6224,N_6302);
nand U6691 (N_6691,N_6046,N_6326);
nor U6692 (N_6692,N_6195,N_6380);
nand U6693 (N_6693,N_6227,N_6442);
nor U6694 (N_6694,N_6401,N_6479);
xor U6695 (N_6695,N_6223,N_6154);
nand U6696 (N_6696,N_6330,N_6432);
nand U6697 (N_6697,N_6425,N_6474);
nor U6698 (N_6698,N_6113,N_6220);
or U6699 (N_6699,N_6019,N_6338);
or U6700 (N_6700,N_6382,N_6231);
and U6701 (N_6701,N_6355,N_6055);
and U6702 (N_6702,N_6406,N_6296);
and U6703 (N_6703,N_6141,N_6179);
xnor U6704 (N_6704,N_6213,N_6497);
nand U6705 (N_6705,N_6044,N_6009);
or U6706 (N_6706,N_6245,N_6408);
or U6707 (N_6707,N_6137,N_6039);
nand U6708 (N_6708,N_6144,N_6407);
nor U6709 (N_6709,N_6229,N_6470);
and U6710 (N_6710,N_6467,N_6062);
xor U6711 (N_6711,N_6437,N_6271);
xnor U6712 (N_6712,N_6066,N_6130);
xnor U6713 (N_6713,N_6347,N_6308);
or U6714 (N_6714,N_6091,N_6228);
and U6715 (N_6715,N_6234,N_6117);
and U6716 (N_6716,N_6109,N_6360);
nor U6717 (N_6717,N_6344,N_6305);
nor U6718 (N_6718,N_6053,N_6102);
and U6719 (N_6719,N_6327,N_6186);
xnor U6720 (N_6720,N_6394,N_6040);
nand U6721 (N_6721,N_6391,N_6057);
xor U6722 (N_6722,N_6323,N_6353);
and U6723 (N_6723,N_6321,N_6163);
and U6724 (N_6724,N_6132,N_6038);
or U6725 (N_6725,N_6185,N_6340);
and U6726 (N_6726,N_6024,N_6105);
and U6727 (N_6727,N_6288,N_6339);
or U6728 (N_6728,N_6322,N_6157);
nor U6729 (N_6729,N_6112,N_6277);
nand U6730 (N_6730,N_6108,N_6309);
nor U6731 (N_6731,N_6281,N_6094);
or U6732 (N_6732,N_6099,N_6242);
nor U6733 (N_6733,N_6148,N_6126);
nor U6734 (N_6734,N_6443,N_6275);
xnor U6735 (N_6735,N_6334,N_6128);
nor U6736 (N_6736,N_6453,N_6460);
and U6737 (N_6737,N_6369,N_6119);
and U6738 (N_6738,N_6352,N_6241);
xor U6739 (N_6739,N_6485,N_6379);
nor U6740 (N_6740,N_6482,N_6466);
and U6741 (N_6741,N_6083,N_6448);
nand U6742 (N_6742,N_6463,N_6233);
nor U6743 (N_6743,N_6415,N_6206);
nand U6744 (N_6744,N_6076,N_6299);
and U6745 (N_6745,N_6495,N_6035);
and U6746 (N_6746,N_6134,N_6311);
and U6747 (N_6747,N_6129,N_6473);
and U6748 (N_6748,N_6324,N_6260);
or U6749 (N_6749,N_6363,N_6491);
nand U6750 (N_6750,N_6363,N_6093);
and U6751 (N_6751,N_6499,N_6488);
nor U6752 (N_6752,N_6200,N_6202);
or U6753 (N_6753,N_6117,N_6328);
or U6754 (N_6754,N_6059,N_6275);
nor U6755 (N_6755,N_6015,N_6147);
or U6756 (N_6756,N_6157,N_6312);
and U6757 (N_6757,N_6387,N_6498);
xnor U6758 (N_6758,N_6364,N_6177);
or U6759 (N_6759,N_6396,N_6144);
and U6760 (N_6760,N_6174,N_6055);
nor U6761 (N_6761,N_6433,N_6320);
nand U6762 (N_6762,N_6263,N_6000);
nand U6763 (N_6763,N_6217,N_6376);
nand U6764 (N_6764,N_6431,N_6433);
nor U6765 (N_6765,N_6343,N_6083);
or U6766 (N_6766,N_6432,N_6216);
nor U6767 (N_6767,N_6322,N_6342);
and U6768 (N_6768,N_6183,N_6190);
nor U6769 (N_6769,N_6493,N_6284);
xor U6770 (N_6770,N_6127,N_6005);
nor U6771 (N_6771,N_6419,N_6130);
nor U6772 (N_6772,N_6011,N_6113);
nor U6773 (N_6773,N_6146,N_6361);
nor U6774 (N_6774,N_6255,N_6157);
or U6775 (N_6775,N_6211,N_6141);
or U6776 (N_6776,N_6475,N_6149);
and U6777 (N_6777,N_6441,N_6161);
and U6778 (N_6778,N_6242,N_6396);
xor U6779 (N_6779,N_6075,N_6134);
and U6780 (N_6780,N_6437,N_6377);
or U6781 (N_6781,N_6466,N_6182);
nand U6782 (N_6782,N_6451,N_6248);
and U6783 (N_6783,N_6371,N_6020);
and U6784 (N_6784,N_6425,N_6459);
and U6785 (N_6785,N_6203,N_6035);
nand U6786 (N_6786,N_6270,N_6088);
nor U6787 (N_6787,N_6130,N_6293);
nand U6788 (N_6788,N_6045,N_6093);
nand U6789 (N_6789,N_6381,N_6103);
xnor U6790 (N_6790,N_6181,N_6254);
nor U6791 (N_6791,N_6040,N_6205);
or U6792 (N_6792,N_6452,N_6010);
nand U6793 (N_6793,N_6384,N_6311);
nor U6794 (N_6794,N_6148,N_6363);
nand U6795 (N_6795,N_6099,N_6337);
and U6796 (N_6796,N_6079,N_6092);
or U6797 (N_6797,N_6371,N_6315);
xor U6798 (N_6798,N_6218,N_6476);
nor U6799 (N_6799,N_6471,N_6447);
nand U6800 (N_6800,N_6382,N_6172);
xor U6801 (N_6801,N_6061,N_6097);
and U6802 (N_6802,N_6350,N_6101);
nor U6803 (N_6803,N_6110,N_6467);
nand U6804 (N_6804,N_6306,N_6130);
nor U6805 (N_6805,N_6058,N_6416);
or U6806 (N_6806,N_6440,N_6032);
nor U6807 (N_6807,N_6416,N_6101);
and U6808 (N_6808,N_6319,N_6471);
xor U6809 (N_6809,N_6441,N_6404);
nor U6810 (N_6810,N_6282,N_6178);
xnor U6811 (N_6811,N_6106,N_6133);
and U6812 (N_6812,N_6232,N_6113);
nand U6813 (N_6813,N_6495,N_6011);
or U6814 (N_6814,N_6031,N_6210);
nor U6815 (N_6815,N_6065,N_6335);
and U6816 (N_6816,N_6204,N_6444);
or U6817 (N_6817,N_6433,N_6271);
nor U6818 (N_6818,N_6061,N_6058);
nand U6819 (N_6819,N_6019,N_6357);
and U6820 (N_6820,N_6488,N_6214);
and U6821 (N_6821,N_6144,N_6355);
and U6822 (N_6822,N_6072,N_6239);
and U6823 (N_6823,N_6123,N_6102);
and U6824 (N_6824,N_6138,N_6373);
nor U6825 (N_6825,N_6209,N_6463);
nand U6826 (N_6826,N_6156,N_6381);
and U6827 (N_6827,N_6068,N_6104);
nor U6828 (N_6828,N_6212,N_6165);
nand U6829 (N_6829,N_6265,N_6229);
and U6830 (N_6830,N_6076,N_6258);
or U6831 (N_6831,N_6110,N_6291);
or U6832 (N_6832,N_6311,N_6330);
nand U6833 (N_6833,N_6012,N_6263);
nor U6834 (N_6834,N_6475,N_6408);
or U6835 (N_6835,N_6132,N_6118);
nand U6836 (N_6836,N_6246,N_6243);
or U6837 (N_6837,N_6488,N_6074);
nand U6838 (N_6838,N_6270,N_6334);
nor U6839 (N_6839,N_6498,N_6473);
nor U6840 (N_6840,N_6455,N_6040);
xor U6841 (N_6841,N_6062,N_6213);
nand U6842 (N_6842,N_6198,N_6207);
xnor U6843 (N_6843,N_6044,N_6442);
nand U6844 (N_6844,N_6264,N_6414);
nand U6845 (N_6845,N_6181,N_6287);
and U6846 (N_6846,N_6232,N_6327);
nor U6847 (N_6847,N_6248,N_6309);
nand U6848 (N_6848,N_6221,N_6087);
nor U6849 (N_6849,N_6005,N_6189);
nand U6850 (N_6850,N_6293,N_6361);
nor U6851 (N_6851,N_6021,N_6217);
xnor U6852 (N_6852,N_6281,N_6393);
nand U6853 (N_6853,N_6120,N_6066);
or U6854 (N_6854,N_6040,N_6317);
nand U6855 (N_6855,N_6482,N_6371);
and U6856 (N_6856,N_6060,N_6102);
and U6857 (N_6857,N_6080,N_6419);
and U6858 (N_6858,N_6461,N_6052);
nand U6859 (N_6859,N_6152,N_6399);
nand U6860 (N_6860,N_6418,N_6276);
or U6861 (N_6861,N_6042,N_6363);
nor U6862 (N_6862,N_6142,N_6487);
nand U6863 (N_6863,N_6082,N_6443);
or U6864 (N_6864,N_6219,N_6137);
and U6865 (N_6865,N_6022,N_6159);
and U6866 (N_6866,N_6176,N_6023);
or U6867 (N_6867,N_6479,N_6102);
and U6868 (N_6868,N_6282,N_6436);
and U6869 (N_6869,N_6292,N_6128);
nor U6870 (N_6870,N_6241,N_6356);
or U6871 (N_6871,N_6310,N_6149);
xnor U6872 (N_6872,N_6212,N_6177);
or U6873 (N_6873,N_6254,N_6302);
or U6874 (N_6874,N_6146,N_6366);
xor U6875 (N_6875,N_6160,N_6375);
or U6876 (N_6876,N_6225,N_6355);
or U6877 (N_6877,N_6349,N_6378);
nor U6878 (N_6878,N_6394,N_6164);
nor U6879 (N_6879,N_6061,N_6395);
or U6880 (N_6880,N_6121,N_6127);
or U6881 (N_6881,N_6160,N_6411);
xnor U6882 (N_6882,N_6297,N_6388);
and U6883 (N_6883,N_6129,N_6166);
xnor U6884 (N_6884,N_6207,N_6409);
or U6885 (N_6885,N_6212,N_6029);
or U6886 (N_6886,N_6390,N_6470);
nor U6887 (N_6887,N_6013,N_6378);
nor U6888 (N_6888,N_6397,N_6105);
nand U6889 (N_6889,N_6157,N_6348);
nand U6890 (N_6890,N_6101,N_6431);
nand U6891 (N_6891,N_6060,N_6200);
and U6892 (N_6892,N_6289,N_6480);
nand U6893 (N_6893,N_6354,N_6160);
or U6894 (N_6894,N_6148,N_6415);
and U6895 (N_6895,N_6391,N_6467);
or U6896 (N_6896,N_6211,N_6297);
and U6897 (N_6897,N_6060,N_6031);
nand U6898 (N_6898,N_6166,N_6294);
or U6899 (N_6899,N_6293,N_6060);
nand U6900 (N_6900,N_6182,N_6375);
or U6901 (N_6901,N_6142,N_6480);
or U6902 (N_6902,N_6396,N_6444);
and U6903 (N_6903,N_6022,N_6254);
or U6904 (N_6904,N_6224,N_6404);
and U6905 (N_6905,N_6290,N_6050);
and U6906 (N_6906,N_6264,N_6269);
and U6907 (N_6907,N_6388,N_6351);
nor U6908 (N_6908,N_6362,N_6185);
nor U6909 (N_6909,N_6190,N_6112);
and U6910 (N_6910,N_6053,N_6091);
or U6911 (N_6911,N_6104,N_6128);
and U6912 (N_6912,N_6222,N_6163);
or U6913 (N_6913,N_6224,N_6231);
nor U6914 (N_6914,N_6396,N_6476);
or U6915 (N_6915,N_6078,N_6021);
or U6916 (N_6916,N_6048,N_6108);
nor U6917 (N_6917,N_6167,N_6200);
nor U6918 (N_6918,N_6466,N_6167);
xor U6919 (N_6919,N_6396,N_6070);
xnor U6920 (N_6920,N_6129,N_6262);
nor U6921 (N_6921,N_6150,N_6475);
xnor U6922 (N_6922,N_6358,N_6182);
nand U6923 (N_6923,N_6000,N_6197);
nand U6924 (N_6924,N_6077,N_6271);
nand U6925 (N_6925,N_6480,N_6091);
nand U6926 (N_6926,N_6437,N_6297);
or U6927 (N_6927,N_6262,N_6258);
or U6928 (N_6928,N_6454,N_6263);
or U6929 (N_6929,N_6309,N_6189);
nor U6930 (N_6930,N_6463,N_6461);
nor U6931 (N_6931,N_6007,N_6286);
nand U6932 (N_6932,N_6000,N_6355);
nor U6933 (N_6933,N_6323,N_6029);
and U6934 (N_6934,N_6269,N_6274);
and U6935 (N_6935,N_6347,N_6423);
xor U6936 (N_6936,N_6166,N_6258);
nor U6937 (N_6937,N_6109,N_6400);
and U6938 (N_6938,N_6192,N_6362);
nand U6939 (N_6939,N_6355,N_6410);
nor U6940 (N_6940,N_6116,N_6226);
and U6941 (N_6941,N_6164,N_6057);
or U6942 (N_6942,N_6183,N_6293);
nor U6943 (N_6943,N_6155,N_6100);
and U6944 (N_6944,N_6217,N_6387);
and U6945 (N_6945,N_6062,N_6283);
nor U6946 (N_6946,N_6089,N_6181);
and U6947 (N_6947,N_6013,N_6443);
nand U6948 (N_6948,N_6050,N_6272);
or U6949 (N_6949,N_6432,N_6052);
xnor U6950 (N_6950,N_6094,N_6464);
and U6951 (N_6951,N_6394,N_6482);
and U6952 (N_6952,N_6065,N_6337);
nor U6953 (N_6953,N_6299,N_6072);
nor U6954 (N_6954,N_6118,N_6050);
xor U6955 (N_6955,N_6064,N_6324);
or U6956 (N_6956,N_6302,N_6012);
or U6957 (N_6957,N_6473,N_6165);
nor U6958 (N_6958,N_6084,N_6200);
or U6959 (N_6959,N_6140,N_6214);
or U6960 (N_6960,N_6119,N_6461);
nor U6961 (N_6961,N_6004,N_6278);
nand U6962 (N_6962,N_6229,N_6284);
nand U6963 (N_6963,N_6192,N_6401);
xor U6964 (N_6964,N_6322,N_6039);
nand U6965 (N_6965,N_6242,N_6171);
nor U6966 (N_6966,N_6190,N_6424);
nor U6967 (N_6967,N_6167,N_6159);
nor U6968 (N_6968,N_6340,N_6119);
nor U6969 (N_6969,N_6364,N_6052);
nand U6970 (N_6970,N_6226,N_6143);
and U6971 (N_6971,N_6465,N_6478);
and U6972 (N_6972,N_6429,N_6048);
and U6973 (N_6973,N_6366,N_6220);
nand U6974 (N_6974,N_6445,N_6389);
nor U6975 (N_6975,N_6248,N_6380);
nor U6976 (N_6976,N_6350,N_6087);
xnor U6977 (N_6977,N_6447,N_6084);
or U6978 (N_6978,N_6168,N_6210);
and U6979 (N_6979,N_6070,N_6311);
nor U6980 (N_6980,N_6239,N_6293);
xor U6981 (N_6981,N_6454,N_6399);
or U6982 (N_6982,N_6365,N_6105);
nand U6983 (N_6983,N_6136,N_6410);
and U6984 (N_6984,N_6347,N_6338);
nand U6985 (N_6985,N_6291,N_6173);
nor U6986 (N_6986,N_6013,N_6372);
nor U6987 (N_6987,N_6187,N_6255);
nor U6988 (N_6988,N_6384,N_6178);
or U6989 (N_6989,N_6308,N_6354);
nand U6990 (N_6990,N_6431,N_6451);
nand U6991 (N_6991,N_6297,N_6013);
or U6992 (N_6992,N_6213,N_6439);
or U6993 (N_6993,N_6374,N_6432);
and U6994 (N_6994,N_6043,N_6402);
or U6995 (N_6995,N_6114,N_6396);
nor U6996 (N_6996,N_6372,N_6288);
nor U6997 (N_6997,N_6119,N_6241);
nand U6998 (N_6998,N_6298,N_6074);
xor U6999 (N_6999,N_6402,N_6218);
or U7000 (N_7000,N_6669,N_6830);
xnor U7001 (N_7001,N_6832,N_6820);
and U7002 (N_7002,N_6732,N_6535);
nor U7003 (N_7003,N_6545,N_6653);
nor U7004 (N_7004,N_6597,N_6739);
nor U7005 (N_7005,N_6549,N_6918);
or U7006 (N_7006,N_6601,N_6897);
nand U7007 (N_7007,N_6706,N_6623);
and U7008 (N_7008,N_6812,N_6514);
nor U7009 (N_7009,N_6756,N_6734);
xor U7010 (N_7010,N_6504,N_6560);
nand U7011 (N_7011,N_6961,N_6677);
or U7012 (N_7012,N_6843,N_6840);
nor U7013 (N_7013,N_6640,N_6748);
or U7014 (N_7014,N_6893,N_6891);
xor U7015 (N_7015,N_6860,N_6790);
or U7016 (N_7016,N_6511,N_6884);
or U7017 (N_7017,N_6707,N_6651);
or U7018 (N_7018,N_6526,N_6510);
nor U7019 (N_7019,N_6829,N_6762);
nand U7020 (N_7020,N_6655,N_6740);
and U7021 (N_7021,N_6696,N_6589);
nor U7022 (N_7022,N_6742,N_6834);
xor U7023 (N_7023,N_6544,N_6555);
and U7024 (N_7024,N_6925,N_6733);
nand U7025 (N_7025,N_6920,N_6643);
nor U7026 (N_7026,N_6596,N_6780);
or U7027 (N_7027,N_6794,N_6939);
nor U7028 (N_7028,N_6695,N_6629);
nor U7029 (N_7029,N_6890,N_6573);
nand U7030 (N_7030,N_6808,N_6804);
nor U7031 (N_7031,N_6693,N_6703);
nor U7032 (N_7032,N_6697,N_6684);
nor U7033 (N_7033,N_6758,N_6996);
nand U7034 (N_7034,N_6543,N_6809);
nor U7035 (N_7035,N_6667,N_6969);
or U7036 (N_7036,N_6691,N_6936);
xor U7037 (N_7037,N_6644,N_6753);
or U7038 (N_7038,N_6594,N_6883);
and U7039 (N_7039,N_6611,N_6675);
nand U7040 (N_7040,N_6531,N_6855);
nor U7041 (N_7041,N_6750,N_6802);
nand U7042 (N_7042,N_6519,N_6507);
nand U7043 (N_7043,N_6603,N_6977);
nand U7044 (N_7044,N_6735,N_6945);
nand U7045 (N_7045,N_6679,N_6767);
and U7046 (N_7046,N_6769,N_6631);
or U7047 (N_7047,N_6971,N_6870);
or U7048 (N_7048,N_6805,N_6578);
xnor U7049 (N_7049,N_6737,N_6931);
nor U7050 (N_7050,N_6888,N_6725);
nor U7051 (N_7051,N_6659,N_6877);
xnor U7052 (N_7052,N_6865,N_6701);
and U7053 (N_7053,N_6646,N_6714);
xor U7054 (N_7054,N_6937,N_6751);
nand U7055 (N_7055,N_6906,N_6574);
or U7056 (N_7056,N_6983,N_6537);
or U7057 (N_7057,N_6953,N_6921);
and U7058 (N_7058,N_6881,N_6728);
or U7059 (N_7059,N_6604,N_6817);
nand U7060 (N_7060,N_6503,N_6729);
or U7061 (N_7061,N_6869,N_6513);
nand U7062 (N_7062,N_6943,N_6582);
nor U7063 (N_7063,N_6864,N_6664);
and U7064 (N_7064,N_6642,N_6871);
xor U7065 (N_7065,N_6827,N_6911);
nor U7066 (N_7066,N_6878,N_6766);
xnor U7067 (N_7067,N_6520,N_6889);
nand U7068 (N_7068,N_6521,N_6894);
nand U7069 (N_7069,N_6602,N_6689);
or U7070 (N_7070,N_6968,N_6502);
nor U7071 (N_7071,N_6821,N_6579);
and U7072 (N_7072,N_6874,N_6856);
nor U7073 (N_7073,N_6956,N_6610);
nor U7074 (N_7074,N_6775,N_6752);
and U7075 (N_7075,N_6654,N_6831);
and U7076 (N_7076,N_6731,N_6588);
nor U7077 (N_7077,N_6622,N_6556);
and U7078 (N_7078,N_6929,N_6710);
nor U7079 (N_7079,N_6959,N_6946);
and U7080 (N_7080,N_6845,N_6630);
nand U7081 (N_7081,N_6786,N_6999);
nand U7082 (N_7082,N_6803,N_6720);
nand U7083 (N_7083,N_6641,N_6847);
or U7084 (N_7084,N_6564,N_6744);
nand U7085 (N_7085,N_6711,N_6719);
nand U7086 (N_7086,N_6846,N_6614);
nor U7087 (N_7087,N_6776,N_6960);
nand U7088 (N_7088,N_6913,N_6987);
nand U7089 (N_7089,N_6765,N_6822);
and U7090 (N_7090,N_6976,N_6620);
nor U7091 (N_7091,N_6958,N_6721);
nand U7092 (N_7092,N_6788,N_6715);
nor U7093 (N_7093,N_6542,N_6798);
or U7094 (N_7094,N_6599,N_6837);
nor U7095 (N_7095,N_6963,N_6523);
xor U7096 (N_7096,N_6704,N_6508);
nor U7097 (N_7097,N_6981,N_6824);
nor U7098 (N_7098,N_6718,N_6974);
nor U7099 (N_7099,N_6928,N_6687);
or U7100 (N_7100,N_6815,N_6896);
and U7101 (N_7101,N_6636,N_6778);
and U7102 (N_7102,N_6652,N_6517);
nand U7103 (N_7103,N_6559,N_6650);
xor U7104 (N_7104,N_6932,N_6858);
nand U7105 (N_7105,N_6944,N_6593);
nand U7106 (N_7106,N_6852,N_6992);
and U7107 (N_7107,N_6626,N_6606);
and U7108 (N_7108,N_6527,N_6685);
and U7109 (N_7109,N_6850,N_6998);
and U7110 (N_7110,N_6909,N_6712);
nor U7111 (N_7111,N_6518,N_6532);
and U7112 (N_7112,N_6615,N_6668);
nand U7113 (N_7113,N_6577,N_6863);
nand U7114 (N_7114,N_6682,N_6791);
nand U7115 (N_7115,N_6793,N_6773);
or U7116 (N_7116,N_6759,N_6634);
nor U7117 (N_7117,N_6568,N_6940);
and U7118 (N_7118,N_6592,N_6967);
or U7119 (N_7119,N_6616,N_6567);
nor U7120 (N_7120,N_6917,N_6900);
nand U7121 (N_7121,N_6548,N_6880);
nor U7122 (N_7122,N_6576,N_6624);
nor U7123 (N_7123,N_6700,N_6638);
and U7124 (N_7124,N_6617,N_6690);
nor U7125 (N_7125,N_6529,N_6885);
or U7126 (N_7126,N_6770,N_6534);
nand U7127 (N_7127,N_6660,N_6747);
nor U7128 (N_7128,N_6670,N_6661);
nor U7129 (N_7129,N_6970,N_6980);
or U7130 (N_7130,N_6908,N_6882);
nand U7131 (N_7131,N_6924,N_6746);
nor U7132 (N_7132,N_6922,N_6605);
or U7133 (N_7133,N_6783,N_6819);
nor U7134 (N_7134,N_6554,N_6949);
nor U7135 (N_7135,N_6835,N_6525);
or U7136 (N_7136,N_6760,N_6528);
or U7137 (N_7137,N_6892,N_6671);
nand U7138 (N_7138,N_6901,N_6823);
or U7139 (N_7139,N_6886,N_6797);
or U7140 (N_7140,N_6947,N_6982);
and U7141 (N_7141,N_6795,N_6935);
and U7142 (N_7142,N_6930,N_6694);
nand U7143 (N_7143,N_6879,N_6875);
nand U7144 (N_7144,N_6512,N_6853);
xnor U7145 (N_7145,N_6903,N_6699);
or U7146 (N_7146,N_6657,N_6816);
and U7147 (N_7147,N_6645,N_6738);
nand U7148 (N_7148,N_6619,N_6942);
nor U7149 (N_7149,N_6923,N_6779);
and U7150 (N_7150,N_6648,N_6562);
nor U7151 (N_7151,N_6698,N_6515);
nor U7152 (N_7152,N_6872,N_6551);
nand U7153 (N_7153,N_6964,N_6806);
nand U7154 (N_7154,N_6771,N_6800);
and U7155 (N_7155,N_6663,N_6912);
and U7156 (N_7156,N_6849,N_6565);
or U7157 (N_7157,N_6833,N_6566);
nor U7158 (N_7158,N_6867,N_6975);
or U7159 (N_7159,N_6557,N_6989);
xnor U7160 (N_7160,N_6763,N_6647);
and U7161 (N_7161,N_6919,N_6506);
nand U7162 (N_7162,N_6501,N_6625);
and U7163 (N_7163,N_6635,N_6723);
nand U7164 (N_7164,N_6789,N_6941);
nor U7165 (N_7165,N_6524,N_6590);
and U7166 (N_7166,N_6768,N_6536);
nor U7167 (N_7167,N_6705,N_6990);
or U7168 (N_7168,N_6522,N_6627);
xnor U7169 (N_7169,N_6965,N_6632);
xnor U7170 (N_7170,N_6836,N_6757);
and U7171 (N_7171,N_6995,N_6633);
and U7172 (N_7172,N_6584,N_6637);
nor U7173 (N_7173,N_6954,N_6814);
nor U7174 (N_7174,N_6844,N_6674);
or U7175 (N_7175,N_6583,N_6828);
nand U7176 (N_7176,N_6957,N_6541);
nor U7177 (N_7177,N_6859,N_6955);
nor U7178 (N_7178,N_6561,N_6618);
nor U7179 (N_7179,N_6799,N_6796);
xnor U7180 (N_7180,N_6962,N_6952);
xor U7181 (N_7181,N_6785,N_6581);
and U7182 (N_7182,N_6585,N_6772);
nor U7183 (N_7183,N_6571,N_6997);
nand U7184 (N_7184,N_6727,N_6774);
and U7185 (N_7185,N_6781,N_6966);
or U7186 (N_7186,N_6726,N_6902);
and U7187 (N_7187,N_6683,N_6713);
and U7188 (N_7188,N_6716,N_6777);
xor U7189 (N_7189,N_6842,N_6741);
nand U7190 (N_7190,N_6672,N_6658);
nor U7191 (N_7191,N_6587,N_6708);
or U7192 (N_7192,N_6991,N_6933);
or U7193 (N_7193,N_6784,N_6628);
and U7194 (N_7194,N_6826,N_6916);
nand U7195 (N_7195,N_6595,N_6782);
and U7196 (N_7196,N_6973,N_6533);
nand U7197 (N_7197,N_6539,N_6538);
nor U7198 (N_7198,N_6563,N_6607);
nand U7199 (N_7199,N_6612,N_6938);
and U7200 (N_7200,N_6818,N_6761);
nor U7201 (N_7201,N_6702,N_6950);
xor U7202 (N_7202,N_6993,N_6979);
or U7203 (N_7203,N_6730,N_6540);
or U7204 (N_7204,N_6861,N_6811);
or U7205 (N_7205,N_6792,N_6907);
or U7206 (N_7206,N_6866,N_6807);
nand U7207 (N_7207,N_6686,N_6580);
nand U7208 (N_7208,N_6899,N_6810);
nand U7209 (N_7209,N_6665,N_6500);
and U7210 (N_7210,N_6552,N_6984);
nor U7211 (N_7211,N_6673,N_6986);
nand U7212 (N_7212,N_6621,N_6898);
nand U7213 (N_7213,N_6745,N_6988);
and U7214 (N_7214,N_6609,N_6600);
nor U7215 (N_7215,N_6724,N_6895);
nor U7216 (N_7216,N_6680,N_6951);
nand U7217 (N_7217,N_6676,N_6586);
xnor U7218 (N_7218,N_6550,N_6915);
nand U7219 (N_7219,N_6857,N_6755);
and U7220 (N_7220,N_6553,N_6509);
or U7221 (N_7221,N_6978,N_6910);
and U7222 (N_7222,N_6516,N_6838);
xor U7223 (N_7223,N_6743,N_6887);
nand U7224 (N_7224,N_6764,N_6591);
nor U7225 (N_7225,N_6905,N_6570);
nor U7226 (N_7226,N_6613,N_6547);
nor U7227 (N_7227,N_6749,N_6688);
nand U7228 (N_7228,N_6927,N_6575);
or U7229 (N_7229,N_6558,N_6972);
nand U7230 (N_7230,N_6569,N_6656);
and U7231 (N_7231,N_6505,N_6868);
nand U7232 (N_7232,N_6994,N_6862);
and U7233 (N_7233,N_6722,N_6598);
and U7234 (N_7234,N_6639,N_6926);
and U7235 (N_7235,N_6985,N_6662);
and U7236 (N_7236,N_6934,N_6848);
nand U7237 (N_7237,N_6914,N_6546);
xor U7238 (N_7238,N_6572,N_6709);
xor U7239 (N_7239,N_6841,N_6904);
nor U7240 (N_7240,N_6876,N_6851);
nand U7241 (N_7241,N_6678,N_6530);
nand U7242 (N_7242,N_6948,N_6787);
nand U7243 (N_7243,N_6736,N_6754);
nand U7244 (N_7244,N_6825,N_6873);
and U7245 (N_7245,N_6692,N_6666);
nor U7246 (N_7246,N_6854,N_6649);
or U7247 (N_7247,N_6717,N_6608);
nand U7248 (N_7248,N_6839,N_6813);
nor U7249 (N_7249,N_6801,N_6681);
nor U7250 (N_7250,N_6512,N_6710);
and U7251 (N_7251,N_6782,N_6621);
xor U7252 (N_7252,N_6707,N_6660);
xnor U7253 (N_7253,N_6882,N_6548);
xor U7254 (N_7254,N_6786,N_6856);
nand U7255 (N_7255,N_6852,N_6832);
or U7256 (N_7256,N_6598,N_6607);
and U7257 (N_7257,N_6543,N_6596);
xnor U7258 (N_7258,N_6752,N_6899);
nor U7259 (N_7259,N_6739,N_6795);
or U7260 (N_7260,N_6704,N_6793);
or U7261 (N_7261,N_6666,N_6688);
xor U7262 (N_7262,N_6876,N_6937);
nand U7263 (N_7263,N_6611,N_6801);
or U7264 (N_7264,N_6669,N_6699);
nand U7265 (N_7265,N_6997,N_6655);
or U7266 (N_7266,N_6922,N_6545);
and U7267 (N_7267,N_6855,N_6548);
nor U7268 (N_7268,N_6923,N_6880);
nand U7269 (N_7269,N_6779,N_6788);
and U7270 (N_7270,N_6642,N_6823);
nor U7271 (N_7271,N_6655,N_6994);
or U7272 (N_7272,N_6516,N_6541);
and U7273 (N_7273,N_6636,N_6707);
nand U7274 (N_7274,N_6983,N_6688);
nor U7275 (N_7275,N_6919,N_6813);
and U7276 (N_7276,N_6848,N_6916);
nor U7277 (N_7277,N_6833,N_6776);
nand U7278 (N_7278,N_6714,N_6835);
nand U7279 (N_7279,N_6809,N_6799);
and U7280 (N_7280,N_6789,N_6643);
and U7281 (N_7281,N_6820,N_6959);
nand U7282 (N_7282,N_6863,N_6751);
nand U7283 (N_7283,N_6833,N_6693);
nand U7284 (N_7284,N_6852,N_6829);
nor U7285 (N_7285,N_6949,N_6607);
and U7286 (N_7286,N_6824,N_6677);
or U7287 (N_7287,N_6635,N_6654);
and U7288 (N_7288,N_6873,N_6626);
xnor U7289 (N_7289,N_6752,N_6527);
and U7290 (N_7290,N_6935,N_6753);
and U7291 (N_7291,N_6796,N_6671);
nand U7292 (N_7292,N_6571,N_6919);
and U7293 (N_7293,N_6975,N_6724);
nor U7294 (N_7294,N_6862,N_6945);
nor U7295 (N_7295,N_6795,N_6806);
nor U7296 (N_7296,N_6930,N_6663);
nand U7297 (N_7297,N_6927,N_6673);
or U7298 (N_7298,N_6564,N_6529);
nand U7299 (N_7299,N_6727,N_6709);
and U7300 (N_7300,N_6849,N_6626);
nor U7301 (N_7301,N_6943,N_6659);
xnor U7302 (N_7302,N_6501,N_6872);
nor U7303 (N_7303,N_6721,N_6807);
and U7304 (N_7304,N_6723,N_6616);
nand U7305 (N_7305,N_6849,N_6797);
nand U7306 (N_7306,N_6971,N_6562);
nor U7307 (N_7307,N_6587,N_6832);
and U7308 (N_7308,N_6795,N_6577);
nor U7309 (N_7309,N_6895,N_6598);
nor U7310 (N_7310,N_6750,N_6785);
and U7311 (N_7311,N_6856,N_6729);
and U7312 (N_7312,N_6604,N_6924);
or U7313 (N_7313,N_6526,N_6750);
nor U7314 (N_7314,N_6619,N_6936);
nor U7315 (N_7315,N_6847,N_6721);
and U7316 (N_7316,N_6799,N_6645);
or U7317 (N_7317,N_6797,N_6572);
and U7318 (N_7318,N_6727,N_6570);
nor U7319 (N_7319,N_6858,N_6962);
xnor U7320 (N_7320,N_6982,N_6801);
xnor U7321 (N_7321,N_6739,N_6634);
nor U7322 (N_7322,N_6532,N_6634);
and U7323 (N_7323,N_6529,N_6600);
and U7324 (N_7324,N_6710,N_6621);
and U7325 (N_7325,N_6716,N_6666);
or U7326 (N_7326,N_6594,N_6505);
and U7327 (N_7327,N_6952,N_6747);
or U7328 (N_7328,N_6722,N_6833);
nor U7329 (N_7329,N_6783,N_6820);
nand U7330 (N_7330,N_6569,N_6923);
nand U7331 (N_7331,N_6729,N_6540);
or U7332 (N_7332,N_6771,N_6835);
or U7333 (N_7333,N_6593,N_6557);
nand U7334 (N_7334,N_6710,N_6938);
or U7335 (N_7335,N_6698,N_6520);
and U7336 (N_7336,N_6604,N_6914);
nand U7337 (N_7337,N_6933,N_6574);
and U7338 (N_7338,N_6731,N_6760);
or U7339 (N_7339,N_6721,N_6914);
and U7340 (N_7340,N_6697,N_6746);
and U7341 (N_7341,N_6937,N_6790);
and U7342 (N_7342,N_6987,N_6740);
or U7343 (N_7343,N_6927,N_6657);
nand U7344 (N_7344,N_6590,N_6737);
nor U7345 (N_7345,N_6743,N_6812);
nor U7346 (N_7346,N_6864,N_6899);
and U7347 (N_7347,N_6953,N_6582);
or U7348 (N_7348,N_6768,N_6861);
nor U7349 (N_7349,N_6538,N_6523);
xor U7350 (N_7350,N_6832,N_6616);
and U7351 (N_7351,N_6609,N_6755);
and U7352 (N_7352,N_6587,N_6983);
xnor U7353 (N_7353,N_6532,N_6732);
nand U7354 (N_7354,N_6616,N_6852);
or U7355 (N_7355,N_6978,N_6902);
and U7356 (N_7356,N_6904,N_6839);
xnor U7357 (N_7357,N_6686,N_6534);
or U7358 (N_7358,N_6890,N_6814);
or U7359 (N_7359,N_6919,N_6860);
nand U7360 (N_7360,N_6968,N_6769);
or U7361 (N_7361,N_6665,N_6543);
nand U7362 (N_7362,N_6762,N_6865);
nand U7363 (N_7363,N_6683,N_6624);
xnor U7364 (N_7364,N_6756,N_6689);
or U7365 (N_7365,N_6905,N_6641);
or U7366 (N_7366,N_6641,N_6643);
nand U7367 (N_7367,N_6581,N_6812);
or U7368 (N_7368,N_6899,N_6974);
nor U7369 (N_7369,N_6981,N_6781);
and U7370 (N_7370,N_6826,N_6871);
xnor U7371 (N_7371,N_6695,N_6693);
xor U7372 (N_7372,N_6548,N_6644);
and U7373 (N_7373,N_6828,N_6996);
xnor U7374 (N_7374,N_6965,N_6709);
and U7375 (N_7375,N_6765,N_6810);
xnor U7376 (N_7376,N_6872,N_6537);
and U7377 (N_7377,N_6978,N_6809);
xor U7378 (N_7378,N_6811,N_6760);
xnor U7379 (N_7379,N_6883,N_6652);
nand U7380 (N_7380,N_6909,N_6876);
xor U7381 (N_7381,N_6852,N_6567);
and U7382 (N_7382,N_6931,N_6640);
nor U7383 (N_7383,N_6964,N_6686);
or U7384 (N_7384,N_6551,N_6528);
and U7385 (N_7385,N_6690,N_6685);
or U7386 (N_7386,N_6634,N_6824);
or U7387 (N_7387,N_6838,N_6893);
or U7388 (N_7388,N_6811,N_6599);
nand U7389 (N_7389,N_6522,N_6703);
or U7390 (N_7390,N_6623,N_6590);
nor U7391 (N_7391,N_6861,N_6525);
nand U7392 (N_7392,N_6710,N_6767);
nor U7393 (N_7393,N_6801,N_6553);
and U7394 (N_7394,N_6915,N_6922);
nor U7395 (N_7395,N_6865,N_6604);
xor U7396 (N_7396,N_6901,N_6697);
nor U7397 (N_7397,N_6986,N_6702);
nand U7398 (N_7398,N_6991,N_6927);
xor U7399 (N_7399,N_6989,N_6791);
and U7400 (N_7400,N_6796,N_6724);
or U7401 (N_7401,N_6812,N_6724);
nand U7402 (N_7402,N_6913,N_6545);
nor U7403 (N_7403,N_6764,N_6996);
nand U7404 (N_7404,N_6935,N_6803);
or U7405 (N_7405,N_6569,N_6852);
nand U7406 (N_7406,N_6860,N_6772);
nand U7407 (N_7407,N_6531,N_6992);
or U7408 (N_7408,N_6650,N_6748);
xor U7409 (N_7409,N_6805,N_6658);
xnor U7410 (N_7410,N_6753,N_6870);
or U7411 (N_7411,N_6707,N_6653);
or U7412 (N_7412,N_6670,N_6593);
nor U7413 (N_7413,N_6771,N_6996);
nor U7414 (N_7414,N_6932,N_6936);
or U7415 (N_7415,N_6687,N_6868);
nand U7416 (N_7416,N_6906,N_6826);
xnor U7417 (N_7417,N_6620,N_6946);
nand U7418 (N_7418,N_6936,N_6604);
or U7419 (N_7419,N_6949,N_6781);
and U7420 (N_7420,N_6502,N_6855);
or U7421 (N_7421,N_6981,N_6830);
or U7422 (N_7422,N_6821,N_6521);
nand U7423 (N_7423,N_6942,N_6895);
and U7424 (N_7424,N_6816,N_6569);
nor U7425 (N_7425,N_6590,N_6865);
and U7426 (N_7426,N_6767,N_6714);
or U7427 (N_7427,N_6559,N_6838);
nor U7428 (N_7428,N_6881,N_6978);
nand U7429 (N_7429,N_6876,N_6510);
nand U7430 (N_7430,N_6558,N_6769);
nand U7431 (N_7431,N_6984,N_6769);
or U7432 (N_7432,N_6522,N_6922);
and U7433 (N_7433,N_6523,N_6714);
nor U7434 (N_7434,N_6756,N_6706);
and U7435 (N_7435,N_6604,N_6886);
nor U7436 (N_7436,N_6822,N_6839);
or U7437 (N_7437,N_6817,N_6779);
nand U7438 (N_7438,N_6671,N_6504);
and U7439 (N_7439,N_6720,N_6832);
and U7440 (N_7440,N_6582,N_6778);
or U7441 (N_7441,N_6919,N_6582);
nand U7442 (N_7442,N_6743,N_6537);
xnor U7443 (N_7443,N_6552,N_6943);
nor U7444 (N_7444,N_6757,N_6707);
or U7445 (N_7445,N_6601,N_6890);
or U7446 (N_7446,N_6601,N_6706);
or U7447 (N_7447,N_6894,N_6751);
nor U7448 (N_7448,N_6638,N_6691);
and U7449 (N_7449,N_6803,N_6957);
or U7450 (N_7450,N_6660,N_6556);
and U7451 (N_7451,N_6937,N_6846);
and U7452 (N_7452,N_6898,N_6789);
xor U7453 (N_7453,N_6555,N_6530);
nand U7454 (N_7454,N_6728,N_6769);
nor U7455 (N_7455,N_6680,N_6941);
nand U7456 (N_7456,N_6925,N_6697);
and U7457 (N_7457,N_6576,N_6517);
nor U7458 (N_7458,N_6624,N_6942);
or U7459 (N_7459,N_6836,N_6615);
nand U7460 (N_7460,N_6782,N_6760);
nand U7461 (N_7461,N_6646,N_6516);
and U7462 (N_7462,N_6679,N_6535);
nor U7463 (N_7463,N_6891,N_6915);
nand U7464 (N_7464,N_6911,N_6698);
or U7465 (N_7465,N_6792,N_6962);
xnor U7466 (N_7466,N_6836,N_6600);
and U7467 (N_7467,N_6730,N_6524);
and U7468 (N_7468,N_6827,N_6969);
or U7469 (N_7469,N_6922,N_6626);
and U7470 (N_7470,N_6533,N_6551);
or U7471 (N_7471,N_6600,N_6613);
nor U7472 (N_7472,N_6844,N_6662);
and U7473 (N_7473,N_6957,N_6976);
xor U7474 (N_7474,N_6741,N_6758);
nand U7475 (N_7475,N_6833,N_6548);
nand U7476 (N_7476,N_6701,N_6762);
and U7477 (N_7477,N_6511,N_6817);
nor U7478 (N_7478,N_6834,N_6795);
xnor U7479 (N_7479,N_6971,N_6811);
or U7480 (N_7480,N_6589,N_6953);
nor U7481 (N_7481,N_6517,N_6698);
and U7482 (N_7482,N_6991,N_6706);
nand U7483 (N_7483,N_6643,N_6700);
nor U7484 (N_7484,N_6721,N_6573);
nand U7485 (N_7485,N_6572,N_6670);
nor U7486 (N_7486,N_6517,N_6781);
or U7487 (N_7487,N_6713,N_6754);
and U7488 (N_7488,N_6652,N_6769);
or U7489 (N_7489,N_6856,N_6508);
and U7490 (N_7490,N_6779,N_6724);
nor U7491 (N_7491,N_6512,N_6951);
or U7492 (N_7492,N_6685,N_6662);
or U7493 (N_7493,N_6918,N_6972);
nor U7494 (N_7494,N_6661,N_6805);
or U7495 (N_7495,N_6653,N_6898);
or U7496 (N_7496,N_6517,N_6792);
and U7497 (N_7497,N_6909,N_6967);
nor U7498 (N_7498,N_6701,N_6924);
and U7499 (N_7499,N_6809,N_6662);
nor U7500 (N_7500,N_7221,N_7007);
nor U7501 (N_7501,N_7137,N_7302);
nor U7502 (N_7502,N_7293,N_7349);
nor U7503 (N_7503,N_7224,N_7359);
nand U7504 (N_7504,N_7257,N_7499);
nand U7505 (N_7505,N_7134,N_7121);
and U7506 (N_7506,N_7182,N_7026);
nor U7507 (N_7507,N_7114,N_7415);
nor U7508 (N_7508,N_7020,N_7384);
or U7509 (N_7509,N_7033,N_7338);
nor U7510 (N_7510,N_7309,N_7089);
nand U7511 (N_7511,N_7198,N_7436);
nor U7512 (N_7512,N_7276,N_7018);
or U7513 (N_7513,N_7393,N_7312);
or U7514 (N_7514,N_7357,N_7178);
nand U7515 (N_7515,N_7373,N_7076);
nand U7516 (N_7516,N_7377,N_7285);
and U7517 (N_7517,N_7070,N_7380);
or U7518 (N_7518,N_7253,N_7159);
xnor U7519 (N_7519,N_7484,N_7064);
and U7520 (N_7520,N_7081,N_7039);
and U7521 (N_7521,N_7466,N_7152);
nand U7522 (N_7522,N_7196,N_7268);
nand U7523 (N_7523,N_7270,N_7244);
and U7524 (N_7524,N_7497,N_7226);
and U7525 (N_7525,N_7489,N_7455);
nor U7526 (N_7526,N_7037,N_7399);
and U7527 (N_7527,N_7019,N_7414);
xor U7528 (N_7528,N_7487,N_7108);
nor U7529 (N_7529,N_7119,N_7311);
nand U7530 (N_7530,N_7124,N_7163);
nor U7531 (N_7531,N_7468,N_7223);
or U7532 (N_7532,N_7021,N_7128);
and U7533 (N_7533,N_7061,N_7122);
and U7534 (N_7534,N_7008,N_7336);
nand U7535 (N_7535,N_7150,N_7495);
and U7536 (N_7536,N_7191,N_7088);
nor U7537 (N_7537,N_7387,N_7168);
nor U7538 (N_7538,N_7104,N_7181);
or U7539 (N_7539,N_7464,N_7188);
and U7540 (N_7540,N_7381,N_7147);
nor U7541 (N_7541,N_7494,N_7288);
and U7542 (N_7542,N_7190,N_7115);
or U7543 (N_7543,N_7162,N_7169);
and U7544 (N_7544,N_7485,N_7421);
and U7545 (N_7545,N_7165,N_7125);
or U7546 (N_7546,N_7245,N_7301);
nand U7547 (N_7547,N_7470,N_7049);
or U7548 (N_7548,N_7011,N_7400);
or U7549 (N_7549,N_7351,N_7475);
nand U7550 (N_7550,N_7457,N_7427);
nand U7551 (N_7551,N_7036,N_7303);
and U7552 (N_7552,N_7207,N_7238);
nor U7553 (N_7553,N_7118,N_7051);
nor U7554 (N_7554,N_7004,N_7385);
or U7555 (N_7555,N_7342,N_7157);
nor U7556 (N_7556,N_7447,N_7291);
nand U7557 (N_7557,N_7363,N_7286);
nand U7558 (N_7558,N_7180,N_7326);
nand U7559 (N_7559,N_7325,N_7106);
and U7560 (N_7560,N_7407,N_7438);
nor U7561 (N_7561,N_7046,N_7452);
nor U7562 (N_7562,N_7343,N_7153);
and U7563 (N_7563,N_7120,N_7142);
or U7564 (N_7564,N_7173,N_7480);
or U7565 (N_7565,N_7298,N_7278);
xor U7566 (N_7566,N_7282,N_7014);
xor U7567 (N_7567,N_7172,N_7174);
or U7568 (N_7568,N_7496,N_7112);
nand U7569 (N_7569,N_7215,N_7237);
and U7570 (N_7570,N_7445,N_7091);
or U7571 (N_7571,N_7056,N_7059);
and U7572 (N_7572,N_7378,N_7320);
and U7573 (N_7573,N_7395,N_7424);
xnor U7574 (N_7574,N_7440,N_7283);
xor U7575 (N_7575,N_7044,N_7100);
or U7576 (N_7576,N_7294,N_7355);
nand U7577 (N_7577,N_7354,N_7360);
nor U7578 (N_7578,N_7366,N_7139);
or U7579 (N_7579,N_7315,N_7473);
nand U7580 (N_7580,N_7346,N_7306);
nand U7581 (N_7581,N_7454,N_7146);
and U7582 (N_7582,N_7166,N_7030);
nand U7583 (N_7583,N_7322,N_7032);
nand U7584 (N_7584,N_7477,N_7370);
nand U7585 (N_7585,N_7175,N_7206);
or U7586 (N_7586,N_7113,N_7193);
nor U7587 (N_7587,N_7300,N_7067);
nand U7588 (N_7588,N_7000,N_7284);
or U7589 (N_7589,N_7231,N_7465);
or U7590 (N_7590,N_7383,N_7358);
nor U7591 (N_7591,N_7154,N_7098);
or U7592 (N_7592,N_7047,N_7161);
and U7593 (N_7593,N_7367,N_7195);
nand U7594 (N_7594,N_7048,N_7390);
or U7595 (N_7595,N_7176,N_7023);
nor U7596 (N_7596,N_7411,N_7187);
xnor U7597 (N_7597,N_7167,N_7469);
xnor U7598 (N_7598,N_7318,N_7218);
or U7599 (N_7599,N_7261,N_7001);
xnor U7600 (N_7600,N_7398,N_7273);
and U7601 (N_7601,N_7297,N_7092);
nand U7602 (N_7602,N_7344,N_7164);
or U7603 (N_7603,N_7027,N_7256);
nand U7604 (N_7604,N_7327,N_7086);
xnor U7605 (N_7605,N_7158,N_7230);
nor U7606 (N_7606,N_7423,N_7266);
nand U7607 (N_7607,N_7317,N_7015);
nand U7608 (N_7608,N_7375,N_7361);
nor U7609 (N_7609,N_7319,N_7127);
xnor U7610 (N_7610,N_7308,N_7107);
and U7611 (N_7611,N_7246,N_7132);
nor U7612 (N_7612,N_7459,N_7211);
and U7613 (N_7613,N_7087,N_7305);
nand U7614 (N_7614,N_7442,N_7332);
nand U7615 (N_7615,N_7350,N_7258);
nand U7616 (N_7616,N_7079,N_7295);
nor U7617 (N_7617,N_7212,N_7434);
nand U7618 (N_7618,N_7274,N_7126);
and U7619 (N_7619,N_7374,N_7210);
or U7620 (N_7620,N_7450,N_7456);
and U7621 (N_7621,N_7394,N_7252);
or U7622 (N_7622,N_7448,N_7209);
nand U7623 (N_7623,N_7225,N_7328);
nand U7624 (N_7624,N_7177,N_7289);
or U7625 (N_7625,N_7202,N_7053);
nand U7626 (N_7626,N_7060,N_7247);
and U7627 (N_7627,N_7123,N_7371);
and U7628 (N_7628,N_7310,N_7185);
nand U7629 (N_7629,N_7203,N_7478);
nor U7630 (N_7630,N_7144,N_7192);
xnor U7631 (N_7631,N_7304,N_7432);
nor U7632 (N_7632,N_7376,N_7262);
nand U7633 (N_7633,N_7280,N_7337);
nor U7634 (N_7634,N_7189,N_7405);
nand U7635 (N_7635,N_7151,N_7419);
nand U7636 (N_7636,N_7422,N_7105);
and U7637 (N_7637,N_7052,N_7229);
and U7638 (N_7638,N_7017,N_7420);
nor U7639 (N_7639,N_7041,N_7009);
nand U7640 (N_7640,N_7233,N_7254);
nor U7641 (N_7641,N_7458,N_7461);
nand U7642 (N_7642,N_7364,N_7208);
xnor U7643 (N_7643,N_7435,N_7271);
nand U7644 (N_7644,N_7031,N_7005);
xnor U7645 (N_7645,N_7382,N_7409);
or U7646 (N_7646,N_7141,N_7038);
nor U7647 (N_7647,N_7186,N_7130);
nand U7648 (N_7648,N_7267,N_7082);
or U7649 (N_7649,N_7093,N_7369);
xor U7650 (N_7650,N_7034,N_7071);
nor U7651 (N_7651,N_7431,N_7340);
and U7652 (N_7652,N_7408,N_7083);
nand U7653 (N_7653,N_7260,N_7022);
nand U7654 (N_7654,N_7402,N_7063);
nor U7655 (N_7655,N_7331,N_7449);
and U7656 (N_7656,N_7073,N_7028);
nand U7657 (N_7657,N_7220,N_7418);
nor U7658 (N_7658,N_7265,N_7428);
nor U7659 (N_7659,N_7148,N_7471);
xor U7660 (N_7660,N_7498,N_7013);
nor U7661 (N_7661,N_7090,N_7010);
nand U7662 (N_7662,N_7437,N_7232);
or U7663 (N_7663,N_7269,N_7216);
and U7664 (N_7664,N_7353,N_7433);
nand U7665 (N_7665,N_7386,N_7099);
nand U7666 (N_7666,N_7149,N_7334);
nand U7667 (N_7667,N_7463,N_7095);
or U7668 (N_7668,N_7429,N_7406);
nand U7669 (N_7669,N_7365,N_7251);
nand U7670 (N_7670,N_7110,N_7129);
nor U7671 (N_7671,N_7050,N_7441);
and U7672 (N_7672,N_7392,N_7102);
xnor U7673 (N_7673,N_7138,N_7016);
nand U7674 (N_7674,N_7314,N_7057);
xor U7675 (N_7675,N_7479,N_7228);
and U7676 (N_7676,N_7025,N_7404);
nor U7677 (N_7677,N_7329,N_7410);
nor U7678 (N_7678,N_7054,N_7179);
nand U7679 (N_7679,N_7263,N_7239);
nor U7680 (N_7680,N_7323,N_7307);
xor U7681 (N_7681,N_7109,N_7277);
and U7682 (N_7682,N_7199,N_7281);
nor U7683 (N_7683,N_7234,N_7012);
and U7684 (N_7684,N_7481,N_7094);
nor U7685 (N_7685,N_7474,N_7096);
or U7686 (N_7686,N_7065,N_7460);
or U7687 (N_7687,N_7476,N_7111);
nor U7688 (N_7688,N_7488,N_7117);
nand U7689 (N_7689,N_7029,N_7486);
nand U7690 (N_7690,N_7439,N_7133);
nand U7691 (N_7691,N_7242,N_7024);
and U7692 (N_7692,N_7313,N_7492);
or U7693 (N_7693,N_7356,N_7483);
nand U7694 (N_7694,N_7101,N_7035);
and U7695 (N_7695,N_7074,N_7401);
or U7696 (N_7696,N_7379,N_7058);
and U7697 (N_7697,N_7170,N_7084);
or U7698 (N_7698,N_7335,N_7068);
or U7699 (N_7699,N_7240,N_7145);
and U7700 (N_7700,N_7131,N_7347);
and U7701 (N_7701,N_7491,N_7482);
or U7702 (N_7702,N_7264,N_7416);
xnor U7703 (N_7703,N_7160,N_7201);
nand U7704 (N_7704,N_7316,N_7391);
nand U7705 (N_7705,N_7430,N_7243);
nor U7706 (N_7706,N_7080,N_7200);
or U7707 (N_7707,N_7227,N_7446);
and U7708 (N_7708,N_7287,N_7040);
nor U7709 (N_7709,N_7472,N_7451);
and U7710 (N_7710,N_7235,N_7417);
nand U7711 (N_7711,N_7426,N_7072);
nor U7712 (N_7712,N_7248,N_7236);
or U7713 (N_7713,N_7339,N_7213);
nor U7714 (N_7714,N_7043,N_7171);
or U7715 (N_7715,N_7292,N_7183);
nand U7716 (N_7716,N_7204,N_7413);
nor U7717 (N_7717,N_7066,N_7156);
and U7718 (N_7718,N_7241,N_7042);
or U7719 (N_7719,N_7348,N_7194);
nor U7720 (N_7720,N_7279,N_7321);
and U7721 (N_7721,N_7249,N_7467);
or U7722 (N_7722,N_7324,N_7214);
nor U7723 (N_7723,N_7205,N_7362);
and U7724 (N_7724,N_7062,N_7003);
and U7725 (N_7725,N_7250,N_7155);
nand U7726 (N_7726,N_7184,N_7345);
nand U7727 (N_7727,N_7259,N_7143);
and U7728 (N_7728,N_7290,N_7403);
and U7729 (N_7729,N_7006,N_7490);
nor U7730 (N_7730,N_7368,N_7272);
xnor U7731 (N_7731,N_7352,N_7299);
nor U7732 (N_7732,N_7135,N_7085);
xnor U7733 (N_7733,N_7219,N_7002);
or U7734 (N_7734,N_7140,N_7330);
nand U7735 (N_7735,N_7136,N_7397);
nand U7736 (N_7736,N_7296,N_7493);
xor U7737 (N_7737,N_7217,N_7255);
nand U7738 (N_7738,N_7389,N_7462);
and U7739 (N_7739,N_7078,N_7077);
or U7740 (N_7740,N_7396,N_7453);
or U7741 (N_7741,N_7097,N_7275);
nand U7742 (N_7742,N_7333,N_7444);
and U7743 (N_7743,N_7412,N_7055);
xor U7744 (N_7744,N_7069,N_7045);
and U7745 (N_7745,N_7103,N_7372);
and U7746 (N_7746,N_7075,N_7388);
and U7747 (N_7747,N_7443,N_7341);
xnor U7748 (N_7748,N_7222,N_7116);
xnor U7749 (N_7749,N_7197,N_7425);
nor U7750 (N_7750,N_7437,N_7339);
or U7751 (N_7751,N_7154,N_7271);
and U7752 (N_7752,N_7119,N_7299);
nand U7753 (N_7753,N_7078,N_7148);
nand U7754 (N_7754,N_7167,N_7272);
xnor U7755 (N_7755,N_7427,N_7451);
nand U7756 (N_7756,N_7164,N_7493);
and U7757 (N_7757,N_7385,N_7104);
and U7758 (N_7758,N_7119,N_7496);
nand U7759 (N_7759,N_7266,N_7254);
and U7760 (N_7760,N_7486,N_7408);
nand U7761 (N_7761,N_7208,N_7187);
and U7762 (N_7762,N_7397,N_7012);
and U7763 (N_7763,N_7032,N_7101);
nor U7764 (N_7764,N_7442,N_7464);
and U7765 (N_7765,N_7373,N_7137);
nor U7766 (N_7766,N_7378,N_7115);
or U7767 (N_7767,N_7385,N_7015);
nor U7768 (N_7768,N_7033,N_7002);
nor U7769 (N_7769,N_7482,N_7180);
nor U7770 (N_7770,N_7453,N_7408);
nand U7771 (N_7771,N_7092,N_7309);
and U7772 (N_7772,N_7151,N_7307);
nand U7773 (N_7773,N_7288,N_7379);
nor U7774 (N_7774,N_7442,N_7077);
or U7775 (N_7775,N_7147,N_7060);
nand U7776 (N_7776,N_7026,N_7155);
and U7777 (N_7777,N_7078,N_7324);
or U7778 (N_7778,N_7053,N_7304);
xnor U7779 (N_7779,N_7096,N_7290);
or U7780 (N_7780,N_7007,N_7213);
xor U7781 (N_7781,N_7195,N_7313);
nand U7782 (N_7782,N_7059,N_7304);
nor U7783 (N_7783,N_7426,N_7077);
and U7784 (N_7784,N_7325,N_7285);
nand U7785 (N_7785,N_7489,N_7441);
or U7786 (N_7786,N_7299,N_7089);
and U7787 (N_7787,N_7088,N_7103);
nand U7788 (N_7788,N_7374,N_7366);
and U7789 (N_7789,N_7367,N_7379);
nand U7790 (N_7790,N_7306,N_7060);
nor U7791 (N_7791,N_7251,N_7441);
nand U7792 (N_7792,N_7295,N_7320);
or U7793 (N_7793,N_7072,N_7027);
xnor U7794 (N_7794,N_7324,N_7028);
and U7795 (N_7795,N_7151,N_7056);
nand U7796 (N_7796,N_7005,N_7286);
or U7797 (N_7797,N_7094,N_7351);
nand U7798 (N_7798,N_7013,N_7286);
nand U7799 (N_7799,N_7105,N_7162);
or U7800 (N_7800,N_7229,N_7220);
nor U7801 (N_7801,N_7282,N_7194);
or U7802 (N_7802,N_7233,N_7392);
nand U7803 (N_7803,N_7343,N_7209);
nand U7804 (N_7804,N_7216,N_7198);
nor U7805 (N_7805,N_7481,N_7381);
nand U7806 (N_7806,N_7029,N_7206);
and U7807 (N_7807,N_7048,N_7218);
or U7808 (N_7808,N_7442,N_7297);
nor U7809 (N_7809,N_7308,N_7048);
and U7810 (N_7810,N_7343,N_7039);
nand U7811 (N_7811,N_7118,N_7488);
or U7812 (N_7812,N_7350,N_7352);
nor U7813 (N_7813,N_7219,N_7487);
nor U7814 (N_7814,N_7448,N_7227);
nand U7815 (N_7815,N_7338,N_7413);
nor U7816 (N_7816,N_7013,N_7180);
nand U7817 (N_7817,N_7176,N_7035);
xnor U7818 (N_7818,N_7312,N_7246);
nand U7819 (N_7819,N_7377,N_7176);
or U7820 (N_7820,N_7188,N_7402);
nor U7821 (N_7821,N_7288,N_7144);
nand U7822 (N_7822,N_7265,N_7073);
or U7823 (N_7823,N_7309,N_7294);
and U7824 (N_7824,N_7023,N_7471);
nand U7825 (N_7825,N_7337,N_7164);
xnor U7826 (N_7826,N_7128,N_7110);
or U7827 (N_7827,N_7172,N_7473);
or U7828 (N_7828,N_7384,N_7114);
or U7829 (N_7829,N_7029,N_7189);
xnor U7830 (N_7830,N_7431,N_7280);
or U7831 (N_7831,N_7476,N_7423);
or U7832 (N_7832,N_7304,N_7411);
nand U7833 (N_7833,N_7371,N_7068);
and U7834 (N_7834,N_7215,N_7433);
nor U7835 (N_7835,N_7047,N_7329);
nor U7836 (N_7836,N_7228,N_7445);
nand U7837 (N_7837,N_7257,N_7428);
nand U7838 (N_7838,N_7097,N_7047);
or U7839 (N_7839,N_7037,N_7186);
and U7840 (N_7840,N_7366,N_7424);
xnor U7841 (N_7841,N_7032,N_7078);
or U7842 (N_7842,N_7302,N_7374);
and U7843 (N_7843,N_7402,N_7271);
and U7844 (N_7844,N_7028,N_7398);
or U7845 (N_7845,N_7230,N_7409);
nor U7846 (N_7846,N_7073,N_7449);
nand U7847 (N_7847,N_7368,N_7254);
nor U7848 (N_7848,N_7497,N_7359);
nor U7849 (N_7849,N_7282,N_7276);
xnor U7850 (N_7850,N_7415,N_7012);
and U7851 (N_7851,N_7174,N_7330);
nor U7852 (N_7852,N_7296,N_7418);
nor U7853 (N_7853,N_7499,N_7222);
nor U7854 (N_7854,N_7159,N_7241);
or U7855 (N_7855,N_7300,N_7237);
and U7856 (N_7856,N_7427,N_7486);
or U7857 (N_7857,N_7025,N_7044);
or U7858 (N_7858,N_7331,N_7041);
and U7859 (N_7859,N_7092,N_7257);
or U7860 (N_7860,N_7074,N_7259);
and U7861 (N_7861,N_7317,N_7452);
and U7862 (N_7862,N_7290,N_7381);
nand U7863 (N_7863,N_7497,N_7408);
nor U7864 (N_7864,N_7410,N_7241);
nand U7865 (N_7865,N_7358,N_7269);
nor U7866 (N_7866,N_7289,N_7426);
nand U7867 (N_7867,N_7429,N_7030);
or U7868 (N_7868,N_7057,N_7109);
nor U7869 (N_7869,N_7398,N_7435);
and U7870 (N_7870,N_7273,N_7427);
nand U7871 (N_7871,N_7348,N_7336);
xnor U7872 (N_7872,N_7296,N_7263);
nor U7873 (N_7873,N_7121,N_7009);
nand U7874 (N_7874,N_7461,N_7381);
nor U7875 (N_7875,N_7310,N_7354);
and U7876 (N_7876,N_7045,N_7061);
and U7877 (N_7877,N_7235,N_7415);
nand U7878 (N_7878,N_7389,N_7272);
nand U7879 (N_7879,N_7154,N_7099);
nor U7880 (N_7880,N_7096,N_7423);
or U7881 (N_7881,N_7474,N_7357);
or U7882 (N_7882,N_7164,N_7096);
nor U7883 (N_7883,N_7237,N_7268);
and U7884 (N_7884,N_7283,N_7163);
nand U7885 (N_7885,N_7425,N_7118);
and U7886 (N_7886,N_7182,N_7480);
or U7887 (N_7887,N_7017,N_7075);
and U7888 (N_7888,N_7188,N_7309);
xnor U7889 (N_7889,N_7369,N_7491);
nand U7890 (N_7890,N_7483,N_7096);
nand U7891 (N_7891,N_7494,N_7072);
nand U7892 (N_7892,N_7111,N_7365);
or U7893 (N_7893,N_7258,N_7163);
nand U7894 (N_7894,N_7477,N_7155);
and U7895 (N_7895,N_7383,N_7114);
nand U7896 (N_7896,N_7345,N_7005);
or U7897 (N_7897,N_7455,N_7403);
and U7898 (N_7898,N_7117,N_7375);
or U7899 (N_7899,N_7059,N_7385);
nand U7900 (N_7900,N_7181,N_7036);
and U7901 (N_7901,N_7131,N_7135);
and U7902 (N_7902,N_7451,N_7187);
nor U7903 (N_7903,N_7102,N_7415);
nor U7904 (N_7904,N_7449,N_7071);
nand U7905 (N_7905,N_7012,N_7243);
and U7906 (N_7906,N_7441,N_7020);
nor U7907 (N_7907,N_7246,N_7327);
nand U7908 (N_7908,N_7360,N_7461);
and U7909 (N_7909,N_7375,N_7153);
or U7910 (N_7910,N_7405,N_7391);
nor U7911 (N_7911,N_7300,N_7273);
and U7912 (N_7912,N_7346,N_7403);
and U7913 (N_7913,N_7391,N_7177);
nand U7914 (N_7914,N_7024,N_7365);
nand U7915 (N_7915,N_7434,N_7447);
nand U7916 (N_7916,N_7257,N_7401);
xor U7917 (N_7917,N_7205,N_7324);
or U7918 (N_7918,N_7229,N_7079);
and U7919 (N_7919,N_7485,N_7231);
nor U7920 (N_7920,N_7418,N_7330);
nand U7921 (N_7921,N_7253,N_7049);
xnor U7922 (N_7922,N_7476,N_7138);
or U7923 (N_7923,N_7385,N_7414);
nor U7924 (N_7924,N_7398,N_7197);
xor U7925 (N_7925,N_7022,N_7159);
or U7926 (N_7926,N_7141,N_7002);
nand U7927 (N_7927,N_7307,N_7088);
nand U7928 (N_7928,N_7241,N_7261);
nand U7929 (N_7929,N_7151,N_7322);
nor U7930 (N_7930,N_7442,N_7066);
or U7931 (N_7931,N_7211,N_7329);
and U7932 (N_7932,N_7459,N_7037);
nand U7933 (N_7933,N_7240,N_7108);
or U7934 (N_7934,N_7121,N_7109);
nand U7935 (N_7935,N_7217,N_7408);
or U7936 (N_7936,N_7335,N_7352);
nor U7937 (N_7937,N_7459,N_7297);
xnor U7938 (N_7938,N_7026,N_7135);
nor U7939 (N_7939,N_7141,N_7027);
or U7940 (N_7940,N_7332,N_7344);
and U7941 (N_7941,N_7000,N_7184);
and U7942 (N_7942,N_7148,N_7376);
nor U7943 (N_7943,N_7063,N_7202);
nand U7944 (N_7944,N_7143,N_7291);
or U7945 (N_7945,N_7313,N_7436);
or U7946 (N_7946,N_7030,N_7250);
nor U7947 (N_7947,N_7233,N_7265);
or U7948 (N_7948,N_7459,N_7327);
nor U7949 (N_7949,N_7134,N_7196);
xor U7950 (N_7950,N_7468,N_7261);
xor U7951 (N_7951,N_7127,N_7233);
and U7952 (N_7952,N_7286,N_7205);
and U7953 (N_7953,N_7242,N_7109);
or U7954 (N_7954,N_7306,N_7454);
and U7955 (N_7955,N_7319,N_7171);
nand U7956 (N_7956,N_7459,N_7452);
xor U7957 (N_7957,N_7490,N_7275);
nor U7958 (N_7958,N_7343,N_7116);
or U7959 (N_7959,N_7342,N_7356);
xor U7960 (N_7960,N_7298,N_7444);
nand U7961 (N_7961,N_7361,N_7406);
or U7962 (N_7962,N_7125,N_7149);
or U7963 (N_7963,N_7433,N_7118);
or U7964 (N_7964,N_7051,N_7097);
and U7965 (N_7965,N_7459,N_7241);
nor U7966 (N_7966,N_7391,N_7460);
nand U7967 (N_7967,N_7494,N_7368);
or U7968 (N_7968,N_7316,N_7090);
nor U7969 (N_7969,N_7192,N_7401);
nor U7970 (N_7970,N_7354,N_7494);
or U7971 (N_7971,N_7416,N_7354);
xnor U7972 (N_7972,N_7237,N_7131);
and U7973 (N_7973,N_7367,N_7349);
nor U7974 (N_7974,N_7165,N_7462);
or U7975 (N_7975,N_7039,N_7192);
nand U7976 (N_7976,N_7176,N_7302);
or U7977 (N_7977,N_7410,N_7369);
and U7978 (N_7978,N_7070,N_7179);
nor U7979 (N_7979,N_7229,N_7300);
and U7980 (N_7980,N_7070,N_7096);
nor U7981 (N_7981,N_7069,N_7087);
and U7982 (N_7982,N_7468,N_7295);
nor U7983 (N_7983,N_7420,N_7426);
and U7984 (N_7984,N_7015,N_7118);
or U7985 (N_7985,N_7127,N_7055);
or U7986 (N_7986,N_7375,N_7440);
nand U7987 (N_7987,N_7181,N_7425);
nand U7988 (N_7988,N_7252,N_7269);
or U7989 (N_7989,N_7087,N_7044);
nor U7990 (N_7990,N_7119,N_7464);
nand U7991 (N_7991,N_7217,N_7207);
nand U7992 (N_7992,N_7001,N_7214);
nand U7993 (N_7993,N_7425,N_7052);
nand U7994 (N_7994,N_7491,N_7381);
or U7995 (N_7995,N_7212,N_7253);
and U7996 (N_7996,N_7120,N_7314);
and U7997 (N_7997,N_7092,N_7111);
nor U7998 (N_7998,N_7161,N_7268);
xor U7999 (N_7999,N_7227,N_7062);
nor U8000 (N_8000,N_7521,N_7770);
nor U8001 (N_8001,N_7979,N_7848);
and U8002 (N_8002,N_7828,N_7697);
nand U8003 (N_8003,N_7586,N_7615);
and U8004 (N_8004,N_7850,N_7780);
and U8005 (N_8005,N_7565,N_7693);
nor U8006 (N_8006,N_7632,N_7500);
and U8007 (N_8007,N_7569,N_7746);
and U8008 (N_8008,N_7846,N_7610);
nand U8009 (N_8009,N_7662,N_7691);
nand U8010 (N_8010,N_7965,N_7916);
or U8011 (N_8011,N_7687,N_7651);
nand U8012 (N_8012,N_7609,N_7668);
or U8013 (N_8013,N_7556,N_7952);
or U8014 (N_8014,N_7743,N_7690);
nor U8015 (N_8015,N_7958,N_7826);
nor U8016 (N_8016,N_7821,N_7608);
or U8017 (N_8017,N_7625,N_7929);
and U8018 (N_8018,N_7849,N_7857);
nor U8019 (N_8019,N_7841,N_7967);
xor U8020 (N_8020,N_7736,N_7805);
or U8021 (N_8021,N_7833,N_7520);
nor U8022 (N_8022,N_7585,N_7811);
nand U8023 (N_8023,N_7573,N_7781);
and U8024 (N_8024,N_7679,N_7701);
and U8025 (N_8025,N_7506,N_7681);
nor U8026 (N_8026,N_7957,N_7921);
nand U8027 (N_8027,N_7671,N_7657);
nand U8028 (N_8028,N_7791,N_7851);
nand U8029 (N_8029,N_7645,N_7906);
nand U8030 (N_8030,N_7786,N_7815);
and U8031 (N_8031,N_7814,N_7858);
or U8032 (N_8032,N_7750,N_7583);
xor U8033 (N_8033,N_7755,N_7594);
nor U8034 (N_8034,N_7990,N_7935);
or U8035 (N_8035,N_7898,N_7545);
nor U8036 (N_8036,N_7896,N_7882);
nor U8037 (N_8037,N_7852,N_7718);
nor U8038 (N_8038,N_7802,N_7533);
or U8039 (N_8039,N_7526,N_7536);
or U8040 (N_8040,N_7871,N_7963);
nand U8041 (N_8041,N_7669,N_7682);
or U8042 (N_8042,N_7931,N_7689);
nand U8043 (N_8043,N_7540,N_7968);
or U8044 (N_8044,N_7908,N_7999);
nand U8045 (N_8045,N_7670,N_7872);
nor U8046 (N_8046,N_7989,N_7923);
nor U8047 (N_8047,N_7706,N_7897);
nand U8048 (N_8048,N_7991,N_7947);
and U8049 (N_8049,N_7733,N_7862);
and U8050 (N_8050,N_7593,N_7883);
nor U8051 (N_8051,N_7982,N_7723);
nor U8052 (N_8052,N_7887,N_7727);
nand U8053 (N_8053,N_7675,N_7759);
or U8054 (N_8054,N_7638,N_7604);
nor U8055 (N_8055,N_7894,N_7809);
and U8056 (N_8056,N_7808,N_7732);
and U8057 (N_8057,N_7795,N_7839);
nand U8058 (N_8058,N_7823,N_7793);
or U8059 (N_8059,N_7650,N_7762);
and U8060 (N_8060,N_7634,N_7817);
nand U8061 (N_8061,N_7734,N_7885);
nand U8062 (N_8062,N_7960,N_7729);
nor U8063 (N_8063,N_7873,N_7856);
or U8064 (N_8064,N_7877,N_7724);
and U8065 (N_8065,N_7505,N_7768);
nand U8066 (N_8066,N_7584,N_7579);
nand U8067 (N_8067,N_7859,N_7943);
nand U8068 (N_8068,N_7725,N_7562);
nor U8069 (N_8069,N_7629,N_7720);
and U8070 (N_8070,N_7970,N_7806);
and U8071 (N_8071,N_7580,N_7591);
nand U8072 (N_8072,N_7756,N_7938);
nor U8073 (N_8073,N_7603,N_7909);
and U8074 (N_8074,N_7904,N_7782);
nand U8075 (N_8075,N_7899,N_7900);
or U8076 (N_8076,N_7685,N_7757);
nand U8077 (N_8077,N_7698,N_7758);
nor U8078 (N_8078,N_7854,N_7787);
or U8079 (N_8079,N_7560,N_7740);
nand U8080 (N_8080,N_7546,N_7981);
or U8081 (N_8081,N_7978,N_7961);
nor U8082 (N_8082,N_7834,N_7654);
nor U8083 (N_8083,N_7719,N_7576);
or U8084 (N_8084,N_7881,N_7529);
and U8085 (N_8085,N_7715,N_7642);
and U8086 (N_8086,N_7618,N_7575);
xor U8087 (N_8087,N_7702,N_7653);
and U8088 (N_8088,N_7910,N_7503);
or U8089 (N_8089,N_7644,N_7577);
and U8090 (N_8090,N_7507,N_7796);
and U8091 (N_8091,N_7951,N_7964);
or U8092 (N_8092,N_7731,N_7622);
and U8093 (N_8093,N_7527,N_7504);
and U8094 (N_8094,N_7647,N_7643);
nor U8095 (N_8095,N_7518,N_7656);
and U8096 (N_8096,N_7548,N_7774);
or U8097 (N_8097,N_7804,N_7836);
nand U8098 (N_8098,N_7514,N_7624);
nor U8099 (N_8099,N_7599,N_7678);
or U8100 (N_8100,N_7633,N_7926);
or U8101 (N_8101,N_7600,N_7950);
nand U8102 (N_8102,N_7557,N_7879);
nor U8103 (N_8103,N_7892,N_7790);
or U8104 (N_8104,N_7924,N_7801);
and U8105 (N_8105,N_7630,N_7807);
or U8106 (N_8106,N_7710,N_7735);
nor U8107 (N_8107,N_7803,N_7542);
or U8108 (N_8108,N_7972,N_7934);
and U8109 (N_8109,N_7954,N_7554);
nand U8110 (N_8110,N_7700,N_7860);
and U8111 (N_8111,N_7712,N_7832);
or U8112 (N_8112,N_7648,N_7799);
or U8113 (N_8113,N_7831,N_7692);
or U8114 (N_8114,N_7646,N_7601);
or U8115 (N_8115,N_7611,N_7582);
or U8116 (N_8116,N_7661,N_7571);
nand U8117 (N_8117,N_7818,N_7936);
and U8118 (N_8118,N_7984,N_7893);
or U8119 (N_8119,N_7837,N_7513);
or U8120 (N_8120,N_7639,N_7663);
and U8121 (N_8121,N_7528,N_7620);
nor U8122 (N_8122,N_7766,N_7987);
xnor U8123 (N_8123,N_7744,N_7867);
xor U8124 (N_8124,N_7523,N_7707);
nor U8125 (N_8125,N_7855,N_7721);
and U8126 (N_8126,N_7863,N_7544);
or U8127 (N_8127,N_7930,N_7907);
and U8128 (N_8128,N_7946,N_7798);
nor U8129 (N_8129,N_7515,N_7800);
xnor U8130 (N_8130,N_7783,N_7640);
and U8131 (N_8131,N_7709,N_7674);
nand U8132 (N_8132,N_7502,N_7714);
and U8133 (N_8133,N_7775,N_7819);
or U8134 (N_8134,N_7953,N_7959);
xnor U8135 (N_8135,N_7581,N_7613);
xnor U8136 (N_8136,N_7975,N_7912);
and U8137 (N_8137,N_7816,N_7754);
and U8138 (N_8138,N_7568,N_7616);
nor U8139 (N_8139,N_7684,N_7539);
xor U8140 (N_8140,N_7983,N_7997);
or U8141 (N_8141,N_7605,N_7771);
and U8142 (N_8142,N_7917,N_7886);
or U8143 (N_8143,N_7574,N_7920);
or U8144 (N_8144,N_7868,N_7797);
xnor U8145 (N_8145,N_7534,N_7563);
or U8146 (N_8146,N_7884,N_7524);
nand U8147 (N_8147,N_7538,N_7739);
and U8148 (N_8148,N_7680,N_7595);
nor U8149 (N_8149,N_7519,N_7636);
nand U8150 (N_8150,N_7761,N_7728);
or U8151 (N_8151,N_7631,N_7903);
nand U8152 (N_8152,N_7752,N_7876);
nor U8153 (N_8153,N_7748,N_7933);
or U8154 (N_8154,N_7792,N_7665);
and U8155 (N_8155,N_7861,N_7772);
nand U8156 (N_8156,N_7711,N_7925);
or U8157 (N_8157,N_7922,N_7777);
xor U8158 (N_8158,N_7765,N_7673);
and U8159 (N_8159,N_7658,N_7776);
nand U8160 (N_8160,N_7976,N_7511);
or U8161 (N_8161,N_7512,N_7564);
nand U8162 (N_8162,N_7956,N_7626);
nand U8163 (N_8163,N_7566,N_7888);
nand U8164 (N_8164,N_7971,N_7530);
or U8165 (N_8165,N_7649,N_7699);
and U8166 (N_8166,N_7655,N_7590);
nand U8167 (N_8167,N_7704,N_7998);
nor U8168 (N_8168,N_7891,N_7708);
nor U8169 (N_8169,N_7747,N_7703);
and U8170 (N_8170,N_7794,N_7659);
or U8171 (N_8171,N_7785,N_7589);
nor U8172 (N_8172,N_7986,N_7928);
and U8173 (N_8173,N_7870,N_7558);
and U8174 (N_8174,N_7869,N_7901);
nor U8175 (N_8175,N_7864,N_7813);
and U8176 (N_8176,N_7778,N_7945);
xor U8177 (N_8177,N_7614,N_7713);
nand U8178 (N_8178,N_7667,N_7940);
or U8179 (N_8179,N_7623,N_7516);
or U8180 (N_8180,N_7890,N_7764);
nor U8181 (N_8181,N_7822,N_7994);
xnor U8182 (N_8182,N_7779,N_7835);
nor U8183 (N_8183,N_7672,N_7716);
nand U8184 (N_8184,N_7878,N_7843);
and U8185 (N_8185,N_7572,N_7977);
or U8186 (N_8186,N_7722,N_7914);
nor U8187 (N_8187,N_7606,N_7596);
and U8188 (N_8188,N_7559,N_7501);
xnor U8189 (N_8189,N_7829,N_7769);
nand U8190 (N_8190,N_7578,N_7677);
or U8191 (N_8191,N_7866,N_7974);
and U8192 (N_8192,N_7810,N_7830);
or U8193 (N_8193,N_7635,N_7549);
and U8194 (N_8194,N_7607,N_7683);
nand U8195 (N_8195,N_7932,N_7812);
or U8196 (N_8196,N_7918,N_7726);
or U8197 (N_8197,N_7588,N_7717);
or U8198 (N_8198,N_7696,N_7551);
and U8199 (N_8199,N_7510,N_7567);
nand U8200 (N_8200,N_7985,N_7738);
xnor U8201 (N_8201,N_7597,N_7737);
or U8202 (N_8202,N_7955,N_7641);
or U8203 (N_8203,N_7995,N_7637);
nand U8204 (N_8204,N_7784,N_7751);
and U8205 (N_8205,N_7937,N_7525);
xor U8206 (N_8206,N_7973,N_7652);
or U8207 (N_8207,N_7915,N_7842);
and U8208 (N_8208,N_7969,N_7911);
and U8209 (N_8209,N_7587,N_7508);
nand U8210 (N_8210,N_7941,N_7767);
or U8211 (N_8211,N_7944,N_7992);
nor U8212 (N_8212,N_7695,N_7592);
or U8213 (N_8213,N_7621,N_7825);
nand U8214 (N_8214,N_7535,N_7773);
nor U8215 (N_8215,N_7763,N_7942);
nor U8216 (N_8216,N_7745,N_7845);
or U8217 (N_8217,N_7875,N_7996);
xor U8218 (N_8218,N_7628,N_7840);
and U8219 (N_8219,N_7853,N_7820);
and U8220 (N_8220,N_7676,N_7939);
nor U8221 (N_8221,N_7962,N_7619);
or U8222 (N_8222,N_7509,N_7874);
and U8223 (N_8223,N_7532,N_7612);
or U8224 (N_8224,N_7537,N_7570);
and U8225 (N_8225,N_7980,N_7517);
nand U8226 (N_8226,N_7705,N_7760);
or U8227 (N_8227,N_7789,N_7550);
nor U8228 (N_8228,N_7844,N_7686);
xnor U8229 (N_8229,N_7949,N_7543);
or U8230 (N_8230,N_7552,N_7742);
and U8231 (N_8231,N_7666,N_7902);
nand U8232 (N_8232,N_7688,N_7555);
or U8233 (N_8233,N_7865,N_7788);
nand U8234 (N_8234,N_7522,N_7664);
nor U8235 (N_8235,N_7617,N_7847);
and U8236 (N_8236,N_7824,N_7602);
nand U8237 (N_8237,N_7993,N_7895);
or U8238 (N_8238,N_7838,N_7753);
nor U8239 (N_8239,N_7889,N_7827);
or U8240 (N_8240,N_7919,N_7741);
or U8241 (N_8241,N_7927,N_7547);
and U8242 (N_8242,N_7694,N_7553);
nor U8243 (N_8243,N_7913,N_7598);
xor U8244 (N_8244,N_7905,N_7948);
nor U8245 (N_8245,N_7531,N_7966);
xor U8246 (N_8246,N_7880,N_7660);
and U8247 (N_8247,N_7627,N_7749);
nor U8248 (N_8248,N_7988,N_7730);
nor U8249 (N_8249,N_7561,N_7541);
nand U8250 (N_8250,N_7893,N_7606);
xor U8251 (N_8251,N_7581,N_7947);
xnor U8252 (N_8252,N_7540,N_7782);
and U8253 (N_8253,N_7624,N_7694);
and U8254 (N_8254,N_7644,N_7685);
xor U8255 (N_8255,N_7781,N_7761);
nand U8256 (N_8256,N_7509,N_7542);
nand U8257 (N_8257,N_7647,N_7972);
xor U8258 (N_8258,N_7790,N_7909);
xor U8259 (N_8259,N_7945,N_7528);
nand U8260 (N_8260,N_7792,N_7774);
and U8261 (N_8261,N_7813,N_7968);
nand U8262 (N_8262,N_7746,N_7988);
nand U8263 (N_8263,N_7649,N_7852);
nand U8264 (N_8264,N_7747,N_7920);
or U8265 (N_8265,N_7768,N_7798);
or U8266 (N_8266,N_7924,N_7930);
nand U8267 (N_8267,N_7918,N_7704);
or U8268 (N_8268,N_7694,N_7814);
nor U8269 (N_8269,N_7839,N_7660);
or U8270 (N_8270,N_7624,N_7667);
nand U8271 (N_8271,N_7605,N_7975);
and U8272 (N_8272,N_7717,N_7537);
nor U8273 (N_8273,N_7844,N_7799);
and U8274 (N_8274,N_7865,N_7770);
nand U8275 (N_8275,N_7817,N_7990);
nor U8276 (N_8276,N_7608,N_7626);
and U8277 (N_8277,N_7672,N_7846);
and U8278 (N_8278,N_7749,N_7527);
nor U8279 (N_8279,N_7886,N_7563);
or U8280 (N_8280,N_7516,N_7826);
nand U8281 (N_8281,N_7636,N_7560);
xor U8282 (N_8282,N_7634,N_7955);
nor U8283 (N_8283,N_7825,N_7558);
and U8284 (N_8284,N_7926,N_7580);
nor U8285 (N_8285,N_7938,N_7899);
or U8286 (N_8286,N_7881,N_7686);
or U8287 (N_8287,N_7949,N_7864);
nand U8288 (N_8288,N_7945,N_7808);
xnor U8289 (N_8289,N_7558,N_7897);
nor U8290 (N_8290,N_7780,N_7884);
or U8291 (N_8291,N_7858,N_7998);
nand U8292 (N_8292,N_7688,N_7819);
or U8293 (N_8293,N_7666,N_7791);
nor U8294 (N_8294,N_7533,N_7668);
nor U8295 (N_8295,N_7536,N_7901);
nand U8296 (N_8296,N_7735,N_7961);
and U8297 (N_8297,N_7687,N_7894);
nand U8298 (N_8298,N_7815,N_7540);
nand U8299 (N_8299,N_7604,N_7931);
or U8300 (N_8300,N_7683,N_7645);
nand U8301 (N_8301,N_7611,N_7686);
nor U8302 (N_8302,N_7872,N_7646);
nand U8303 (N_8303,N_7876,N_7613);
nand U8304 (N_8304,N_7503,N_7678);
nor U8305 (N_8305,N_7671,N_7632);
xnor U8306 (N_8306,N_7717,N_7907);
or U8307 (N_8307,N_7794,N_7812);
and U8308 (N_8308,N_7503,N_7721);
or U8309 (N_8309,N_7611,N_7831);
or U8310 (N_8310,N_7721,N_7988);
nor U8311 (N_8311,N_7709,N_7942);
nor U8312 (N_8312,N_7844,N_7827);
and U8313 (N_8313,N_7573,N_7504);
or U8314 (N_8314,N_7875,N_7727);
nor U8315 (N_8315,N_7628,N_7787);
or U8316 (N_8316,N_7992,N_7673);
and U8317 (N_8317,N_7896,N_7609);
nand U8318 (N_8318,N_7714,N_7791);
nand U8319 (N_8319,N_7501,N_7533);
or U8320 (N_8320,N_7512,N_7584);
or U8321 (N_8321,N_7584,N_7547);
nand U8322 (N_8322,N_7764,N_7643);
xor U8323 (N_8323,N_7503,N_7632);
and U8324 (N_8324,N_7930,N_7654);
or U8325 (N_8325,N_7937,N_7610);
nor U8326 (N_8326,N_7671,N_7639);
nand U8327 (N_8327,N_7760,N_7633);
nand U8328 (N_8328,N_7774,N_7795);
and U8329 (N_8329,N_7862,N_7610);
and U8330 (N_8330,N_7727,N_7877);
xnor U8331 (N_8331,N_7872,N_7755);
and U8332 (N_8332,N_7606,N_7685);
nor U8333 (N_8333,N_7908,N_7731);
or U8334 (N_8334,N_7691,N_7802);
and U8335 (N_8335,N_7776,N_7585);
or U8336 (N_8336,N_7729,N_7650);
nor U8337 (N_8337,N_7655,N_7812);
and U8338 (N_8338,N_7911,N_7658);
nand U8339 (N_8339,N_7634,N_7858);
or U8340 (N_8340,N_7755,N_7512);
and U8341 (N_8341,N_7724,N_7733);
or U8342 (N_8342,N_7905,N_7659);
nor U8343 (N_8343,N_7522,N_7776);
xnor U8344 (N_8344,N_7725,N_7773);
nor U8345 (N_8345,N_7530,N_7560);
and U8346 (N_8346,N_7874,N_7936);
nor U8347 (N_8347,N_7872,N_7973);
or U8348 (N_8348,N_7787,N_7551);
and U8349 (N_8349,N_7733,N_7686);
nor U8350 (N_8350,N_7892,N_7945);
nand U8351 (N_8351,N_7663,N_7594);
xnor U8352 (N_8352,N_7557,N_7528);
nor U8353 (N_8353,N_7577,N_7529);
nor U8354 (N_8354,N_7732,N_7951);
or U8355 (N_8355,N_7879,N_7713);
nand U8356 (N_8356,N_7892,N_7967);
nor U8357 (N_8357,N_7560,N_7909);
xnor U8358 (N_8358,N_7978,N_7766);
and U8359 (N_8359,N_7622,N_7558);
or U8360 (N_8360,N_7547,N_7585);
and U8361 (N_8361,N_7744,N_7979);
or U8362 (N_8362,N_7745,N_7602);
and U8363 (N_8363,N_7580,N_7842);
and U8364 (N_8364,N_7511,N_7833);
and U8365 (N_8365,N_7855,N_7552);
nand U8366 (N_8366,N_7938,N_7561);
or U8367 (N_8367,N_7846,N_7927);
nand U8368 (N_8368,N_7508,N_7664);
and U8369 (N_8369,N_7663,N_7565);
or U8370 (N_8370,N_7563,N_7511);
and U8371 (N_8371,N_7939,N_7964);
or U8372 (N_8372,N_7550,N_7764);
nor U8373 (N_8373,N_7652,N_7530);
and U8374 (N_8374,N_7657,N_7910);
and U8375 (N_8375,N_7532,N_7695);
and U8376 (N_8376,N_7897,N_7602);
and U8377 (N_8377,N_7662,N_7521);
nor U8378 (N_8378,N_7944,N_7750);
nor U8379 (N_8379,N_7771,N_7916);
or U8380 (N_8380,N_7788,N_7682);
nor U8381 (N_8381,N_7886,N_7719);
nand U8382 (N_8382,N_7559,N_7927);
and U8383 (N_8383,N_7977,N_7930);
or U8384 (N_8384,N_7794,N_7605);
nor U8385 (N_8385,N_7985,N_7597);
nor U8386 (N_8386,N_7798,N_7546);
nor U8387 (N_8387,N_7684,N_7657);
nand U8388 (N_8388,N_7745,N_7916);
and U8389 (N_8389,N_7931,N_7588);
nor U8390 (N_8390,N_7968,N_7742);
nor U8391 (N_8391,N_7999,N_7807);
xnor U8392 (N_8392,N_7536,N_7570);
nand U8393 (N_8393,N_7799,N_7720);
or U8394 (N_8394,N_7910,N_7927);
nand U8395 (N_8395,N_7664,N_7826);
nor U8396 (N_8396,N_7703,N_7501);
nor U8397 (N_8397,N_7556,N_7650);
and U8398 (N_8398,N_7557,N_7751);
or U8399 (N_8399,N_7618,N_7806);
nand U8400 (N_8400,N_7513,N_7771);
nand U8401 (N_8401,N_7651,N_7755);
nand U8402 (N_8402,N_7904,N_7618);
nand U8403 (N_8403,N_7972,N_7825);
or U8404 (N_8404,N_7839,N_7503);
or U8405 (N_8405,N_7784,N_7687);
nand U8406 (N_8406,N_7789,N_7944);
nand U8407 (N_8407,N_7837,N_7698);
or U8408 (N_8408,N_7947,N_7789);
nand U8409 (N_8409,N_7519,N_7647);
and U8410 (N_8410,N_7602,N_7846);
or U8411 (N_8411,N_7644,N_7650);
nor U8412 (N_8412,N_7647,N_7758);
or U8413 (N_8413,N_7819,N_7689);
nand U8414 (N_8414,N_7521,N_7672);
nor U8415 (N_8415,N_7956,N_7986);
or U8416 (N_8416,N_7856,N_7983);
nor U8417 (N_8417,N_7572,N_7812);
nand U8418 (N_8418,N_7775,N_7575);
and U8419 (N_8419,N_7570,N_7883);
or U8420 (N_8420,N_7838,N_7675);
and U8421 (N_8421,N_7554,N_7859);
nand U8422 (N_8422,N_7800,N_7696);
or U8423 (N_8423,N_7545,N_7813);
and U8424 (N_8424,N_7867,N_7692);
and U8425 (N_8425,N_7681,N_7911);
nor U8426 (N_8426,N_7897,N_7658);
nand U8427 (N_8427,N_7860,N_7501);
or U8428 (N_8428,N_7769,N_7959);
nor U8429 (N_8429,N_7897,N_7778);
or U8430 (N_8430,N_7768,N_7568);
or U8431 (N_8431,N_7791,N_7746);
nor U8432 (N_8432,N_7703,N_7617);
nor U8433 (N_8433,N_7870,N_7592);
or U8434 (N_8434,N_7664,N_7696);
or U8435 (N_8435,N_7704,N_7960);
nand U8436 (N_8436,N_7580,N_7679);
nand U8437 (N_8437,N_7548,N_7948);
nand U8438 (N_8438,N_7951,N_7936);
xor U8439 (N_8439,N_7512,N_7605);
xor U8440 (N_8440,N_7596,N_7573);
nor U8441 (N_8441,N_7926,N_7670);
or U8442 (N_8442,N_7958,N_7864);
nor U8443 (N_8443,N_7585,N_7681);
nor U8444 (N_8444,N_7932,N_7745);
nand U8445 (N_8445,N_7861,N_7900);
and U8446 (N_8446,N_7960,N_7854);
nand U8447 (N_8447,N_7594,N_7515);
xnor U8448 (N_8448,N_7571,N_7562);
or U8449 (N_8449,N_7988,N_7940);
nand U8450 (N_8450,N_7821,N_7805);
xnor U8451 (N_8451,N_7608,N_7968);
nor U8452 (N_8452,N_7518,N_7710);
nand U8453 (N_8453,N_7831,N_7892);
nor U8454 (N_8454,N_7964,N_7577);
nand U8455 (N_8455,N_7531,N_7928);
nand U8456 (N_8456,N_7790,N_7523);
nand U8457 (N_8457,N_7901,N_7970);
and U8458 (N_8458,N_7667,N_7970);
or U8459 (N_8459,N_7951,N_7649);
xnor U8460 (N_8460,N_7853,N_7516);
and U8461 (N_8461,N_7958,N_7800);
nor U8462 (N_8462,N_7627,N_7953);
or U8463 (N_8463,N_7607,N_7719);
nand U8464 (N_8464,N_7680,N_7558);
nor U8465 (N_8465,N_7534,N_7725);
nand U8466 (N_8466,N_7886,N_7870);
nor U8467 (N_8467,N_7952,N_7627);
and U8468 (N_8468,N_7983,N_7769);
or U8469 (N_8469,N_7593,N_7971);
or U8470 (N_8470,N_7803,N_7658);
or U8471 (N_8471,N_7977,N_7985);
nand U8472 (N_8472,N_7523,N_7541);
nand U8473 (N_8473,N_7913,N_7800);
and U8474 (N_8474,N_7951,N_7961);
nor U8475 (N_8475,N_7620,N_7775);
nor U8476 (N_8476,N_7909,N_7935);
or U8477 (N_8477,N_7767,N_7679);
or U8478 (N_8478,N_7615,N_7935);
xnor U8479 (N_8479,N_7508,N_7983);
or U8480 (N_8480,N_7694,N_7655);
and U8481 (N_8481,N_7712,N_7991);
nand U8482 (N_8482,N_7556,N_7600);
nor U8483 (N_8483,N_7799,N_7602);
nor U8484 (N_8484,N_7760,N_7603);
or U8485 (N_8485,N_7958,N_7714);
nand U8486 (N_8486,N_7646,N_7622);
nand U8487 (N_8487,N_7756,N_7525);
or U8488 (N_8488,N_7895,N_7648);
or U8489 (N_8489,N_7604,N_7990);
nand U8490 (N_8490,N_7990,N_7770);
and U8491 (N_8491,N_7696,N_7790);
or U8492 (N_8492,N_7711,N_7516);
xor U8493 (N_8493,N_7647,N_7783);
nand U8494 (N_8494,N_7592,N_7717);
or U8495 (N_8495,N_7909,N_7923);
or U8496 (N_8496,N_7566,N_7621);
and U8497 (N_8497,N_7655,N_7849);
nor U8498 (N_8498,N_7767,N_7624);
nand U8499 (N_8499,N_7863,N_7731);
nor U8500 (N_8500,N_8454,N_8440);
or U8501 (N_8501,N_8075,N_8044);
nand U8502 (N_8502,N_8185,N_8322);
nor U8503 (N_8503,N_8333,N_8474);
nor U8504 (N_8504,N_8175,N_8173);
or U8505 (N_8505,N_8152,N_8041);
and U8506 (N_8506,N_8424,N_8006);
and U8507 (N_8507,N_8060,N_8203);
nand U8508 (N_8508,N_8427,N_8222);
nand U8509 (N_8509,N_8218,N_8233);
nand U8510 (N_8510,N_8331,N_8473);
and U8511 (N_8511,N_8104,N_8335);
nand U8512 (N_8512,N_8094,N_8019);
or U8513 (N_8513,N_8141,N_8409);
or U8514 (N_8514,N_8423,N_8392);
nor U8515 (N_8515,N_8193,N_8114);
or U8516 (N_8516,N_8068,N_8268);
and U8517 (N_8517,N_8270,N_8323);
or U8518 (N_8518,N_8192,N_8441);
and U8519 (N_8519,N_8340,N_8237);
xor U8520 (N_8520,N_8299,N_8495);
and U8521 (N_8521,N_8157,N_8490);
xnor U8522 (N_8522,N_8304,N_8425);
xor U8523 (N_8523,N_8083,N_8017);
and U8524 (N_8524,N_8036,N_8384);
nand U8525 (N_8525,N_8415,N_8401);
nand U8526 (N_8526,N_8267,N_8210);
and U8527 (N_8527,N_8007,N_8158);
nor U8528 (N_8528,N_8405,N_8363);
nor U8529 (N_8529,N_8342,N_8265);
xor U8530 (N_8530,N_8232,N_8053);
xor U8531 (N_8531,N_8489,N_8099);
nor U8532 (N_8532,N_8015,N_8277);
and U8533 (N_8533,N_8271,N_8391);
and U8534 (N_8534,N_8123,N_8010);
or U8535 (N_8535,N_8330,N_8071);
xor U8536 (N_8536,N_8397,N_8062);
nand U8537 (N_8537,N_8212,N_8054);
xnor U8538 (N_8538,N_8453,N_8498);
nand U8539 (N_8539,N_8418,N_8096);
xnor U8540 (N_8540,N_8022,N_8181);
and U8541 (N_8541,N_8052,N_8438);
nand U8542 (N_8542,N_8180,N_8122);
nor U8543 (N_8543,N_8219,N_8130);
or U8544 (N_8544,N_8178,N_8263);
and U8545 (N_8545,N_8110,N_8197);
or U8546 (N_8546,N_8244,N_8482);
nor U8547 (N_8547,N_8465,N_8038);
and U8548 (N_8548,N_8201,N_8264);
nand U8549 (N_8549,N_8442,N_8381);
nand U8550 (N_8550,N_8061,N_8162);
nor U8551 (N_8551,N_8356,N_8153);
nor U8552 (N_8552,N_8013,N_8283);
nand U8553 (N_8553,N_8005,N_8382);
nand U8554 (N_8554,N_8393,N_8085);
nand U8555 (N_8555,N_8261,N_8383);
and U8556 (N_8556,N_8084,N_8198);
or U8557 (N_8557,N_8359,N_8477);
and U8558 (N_8558,N_8480,N_8136);
nand U8559 (N_8559,N_8479,N_8009);
nor U8560 (N_8560,N_8021,N_8220);
nor U8561 (N_8561,N_8118,N_8250);
nand U8562 (N_8562,N_8253,N_8371);
and U8563 (N_8563,N_8055,N_8443);
nand U8564 (N_8564,N_8213,N_8476);
nand U8565 (N_8565,N_8460,N_8414);
nor U8566 (N_8566,N_8432,N_8155);
nand U8567 (N_8567,N_8103,N_8372);
and U8568 (N_8568,N_8080,N_8150);
and U8569 (N_8569,N_8360,N_8303);
or U8570 (N_8570,N_8191,N_8296);
nor U8571 (N_8571,N_8182,N_8134);
xnor U8572 (N_8572,N_8279,N_8089);
and U8573 (N_8573,N_8031,N_8127);
nand U8574 (N_8574,N_8327,N_8368);
nor U8575 (N_8575,N_8137,N_8273);
nand U8576 (N_8576,N_8107,N_8126);
nand U8577 (N_8577,N_8163,N_8190);
nor U8578 (N_8578,N_8352,N_8408);
nand U8579 (N_8579,N_8417,N_8001);
nor U8580 (N_8580,N_8289,N_8487);
nor U8581 (N_8581,N_8217,N_8351);
or U8582 (N_8582,N_8170,N_8004);
and U8583 (N_8583,N_8204,N_8147);
and U8584 (N_8584,N_8077,N_8018);
or U8585 (N_8585,N_8366,N_8111);
nor U8586 (N_8586,N_8156,N_8298);
or U8587 (N_8587,N_8098,N_8470);
nand U8588 (N_8588,N_8369,N_8288);
nand U8589 (N_8589,N_8262,N_8025);
or U8590 (N_8590,N_8446,N_8324);
nand U8591 (N_8591,N_8241,N_8499);
nor U8592 (N_8592,N_8135,N_8467);
and U8593 (N_8593,N_8469,N_8164);
nor U8594 (N_8594,N_8257,N_8228);
nand U8595 (N_8595,N_8439,N_8026);
nand U8596 (N_8596,N_8295,N_8419);
nand U8597 (N_8597,N_8399,N_8171);
nor U8598 (N_8598,N_8457,N_8086);
or U8599 (N_8599,N_8205,N_8370);
or U8600 (N_8600,N_8235,N_8145);
nand U8601 (N_8601,N_8406,N_8353);
and U8602 (N_8602,N_8344,N_8373);
nand U8603 (N_8603,N_8362,N_8410);
and U8604 (N_8604,N_8462,N_8389);
and U8605 (N_8605,N_8485,N_8159);
or U8606 (N_8606,N_8374,N_8326);
nand U8607 (N_8607,N_8252,N_8347);
nand U8608 (N_8608,N_8154,N_8112);
or U8609 (N_8609,N_8483,N_8195);
and U8610 (N_8610,N_8073,N_8321);
nand U8611 (N_8611,N_8315,N_8040);
nor U8612 (N_8612,N_8249,N_8272);
or U8613 (N_8613,N_8033,N_8293);
and U8614 (N_8614,N_8269,N_8276);
or U8615 (N_8615,N_8367,N_8000);
nor U8616 (N_8616,N_8102,N_8236);
xor U8617 (N_8617,N_8002,N_8422);
nor U8618 (N_8618,N_8259,N_8176);
nand U8619 (N_8619,N_8196,N_8248);
nand U8620 (N_8620,N_8496,N_8355);
and U8621 (N_8621,N_8493,N_8484);
and U8622 (N_8622,N_8088,N_8200);
xor U8623 (N_8623,N_8497,N_8124);
and U8624 (N_8624,N_8119,N_8003);
nor U8625 (N_8625,N_8254,N_8452);
and U8626 (N_8626,N_8275,N_8278);
nand U8627 (N_8627,N_8229,N_8300);
nor U8628 (N_8628,N_8030,N_8435);
or U8629 (N_8629,N_8357,N_8420);
and U8630 (N_8630,N_8494,N_8144);
or U8631 (N_8631,N_8390,N_8208);
nand U8632 (N_8632,N_8128,N_8207);
and U8633 (N_8633,N_8065,N_8328);
nor U8634 (N_8634,N_8206,N_8108);
and U8635 (N_8635,N_8050,N_8471);
nand U8636 (N_8636,N_8168,N_8142);
nor U8637 (N_8637,N_8459,N_8143);
xor U8638 (N_8638,N_8349,N_8234);
xor U8639 (N_8639,N_8214,N_8202);
nor U8640 (N_8640,N_8069,N_8230);
nor U8641 (N_8641,N_8199,N_8386);
nand U8642 (N_8642,N_8402,N_8165);
nor U8643 (N_8643,N_8140,N_8306);
nand U8644 (N_8644,N_8106,N_8057);
nand U8645 (N_8645,N_8394,N_8121);
or U8646 (N_8646,N_8309,N_8129);
nor U8647 (N_8647,N_8437,N_8243);
xnor U8648 (N_8648,N_8105,N_8255);
and U8649 (N_8649,N_8070,N_8448);
nand U8650 (N_8650,N_8132,N_8297);
xor U8651 (N_8651,N_8285,N_8274);
and U8652 (N_8652,N_8125,N_8308);
nor U8653 (N_8653,N_8395,N_8358);
and U8654 (N_8654,N_8095,N_8133);
and U8655 (N_8655,N_8447,N_8450);
or U8656 (N_8656,N_8318,N_8101);
and U8657 (N_8657,N_8431,N_8047);
xnor U8658 (N_8658,N_8348,N_8231);
and U8659 (N_8659,N_8227,N_8365);
nand U8660 (N_8660,N_8436,N_8314);
xnor U8661 (N_8661,N_8421,N_8043);
nor U8662 (N_8662,N_8354,N_8093);
nor U8663 (N_8663,N_8375,N_8266);
and U8664 (N_8664,N_8037,N_8416);
or U8665 (N_8665,N_8345,N_8247);
nand U8666 (N_8666,N_8238,N_8377);
xor U8667 (N_8667,N_8472,N_8319);
nor U8668 (N_8668,N_8239,N_8316);
and U8669 (N_8669,N_8188,N_8032);
nor U8670 (N_8670,N_8329,N_8117);
and U8671 (N_8671,N_8379,N_8307);
or U8672 (N_8672,N_8341,N_8066);
or U8673 (N_8673,N_8411,N_8429);
nor U8674 (N_8674,N_8292,N_8148);
nand U8675 (N_8675,N_8161,N_8023);
and U8676 (N_8676,N_8337,N_8048);
or U8677 (N_8677,N_8024,N_8310);
nor U8678 (N_8678,N_8014,N_8294);
nor U8679 (N_8679,N_8169,N_8090);
nor U8680 (N_8680,N_8281,N_8475);
nor U8681 (N_8681,N_8412,N_8151);
or U8682 (N_8682,N_8387,N_8413);
nor U8683 (N_8683,N_8100,N_8078);
xor U8684 (N_8684,N_8449,N_8445);
and U8685 (N_8685,N_8146,N_8079);
nand U8686 (N_8686,N_8177,N_8138);
and U8687 (N_8687,N_8035,N_8029);
nand U8688 (N_8688,N_8216,N_8074);
or U8689 (N_8689,N_8388,N_8172);
nand U8690 (N_8690,N_8160,N_8346);
or U8691 (N_8691,N_8183,N_8058);
nor U8692 (N_8692,N_8403,N_8116);
nand U8693 (N_8693,N_8313,N_8317);
nand U8694 (N_8694,N_8028,N_8097);
or U8695 (N_8695,N_8451,N_8067);
or U8696 (N_8696,N_8486,N_8225);
nand U8697 (N_8697,N_8027,N_8492);
nand U8698 (N_8698,N_8221,N_8115);
xor U8699 (N_8699,N_8286,N_8332);
xnor U8700 (N_8700,N_8012,N_8284);
nand U8701 (N_8701,N_8045,N_8302);
nor U8702 (N_8702,N_8082,N_8046);
and U8703 (N_8703,N_8245,N_8456);
and U8704 (N_8704,N_8396,N_8072);
nor U8705 (N_8705,N_8478,N_8224);
nand U8706 (N_8706,N_8139,N_8380);
or U8707 (N_8707,N_8215,N_8209);
nand U8708 (N_8708,N_8184,N_8179);
or U8709 (N_8709,N_8251,N_8282);
nand U8710 (N_8710,N_8056,N_8312);
nand U8711 (N_8711,N_8187,N_8189);
nor U8712 (N_8712,N_8034,N_8076);
nand U8713 (N_8713,N_8051,N_8226);
and U8714 (N_8714,N_8011,N_8320);
nor U8715 (N_8715,N_8194,N_8311);
or U8716 (N_8716,N_8385,N_8338);
xor U8717 (N_8717,N_8301,N_8343);
or U8718 (N_8718,N_8290,N_8378);
or U8719 (N_8719,N_8400,N_8404);
and U8720 (N_8720,N_8081,N_8113);
or U8721 (N_8721,N_8491,N_8242);
or U8722 (N_8722,N_8258,N_8350);
nor U8723 (N_8723,N_8376,N_8287);
or U8724 (N_8724,N_8059,N_8211);
or U8725 (N_8725,N_8223,N_8240);
and U8726 (N_8726,N_8149,N_8120);
nor U8727 (N_8727,N_8186,N_8049);
xor U8728 (N_8728,N_8325,N_8364);
xnor U8729 (N_8729,N_8426,N_8016);
and U8730 (N_8730,N_8458,N_8361);
nand U8731 (N_8731,N_8466,N_8334);
nor U8732 (N_8732,N_8336,N_8131);
or U8733 (N_8733,N_8305,N_8280);
nor U8734 (N_8734,N_8430,N_8339);
and U8735 (N_8735,N_8042,N_8461);
or U8736 (N_8736,N_8291,N_8174);
nand U8737 (N_8737,N_8434,N_8433);
nor U8738 (N_8738,N_8468,N_8260);
nor U8739 (N_8739,N_8488,N_8398);
or U8740 (N_8740,N_8008,N_8481);
and U8741 (N_8741,N_8463,N_8166);
and U8742 (N_8742,N_8039,N_8064);
nor U8743 (N_8743,N_8428,N_8092);
xnor U8744 (N_8744,N_8109,N_8444);
and U8745 (N_8745,N_8455,N_8063);
and U8746 (N_8746,N_8246,N_8407);
and U8747 (N_8747,N_8167,N_8087);
or U8748 (N_8748,N_8020,N_8464);
nor U8749 (N_8749,N_8091,N_8256);
and U8750 (N_8750,N_8162,N_8179);
nor U8751 (N_8751,N_8165,N_8162);
xnor U8752 (N_8752,N_8377,N_8487);
or U8753 (N_8753,N_8126,N_8049);
or U8754 (N_8754,N_8464,N_8424);
and U8755 (N_8755,N_8431,N_8239);
nor U8756 (N_8756,N_8339,N_8435);
and U8757 (N_8757,N_8028,N_8373);
or U8758 (N_8758,N_8323,N_8493);
or U8759 (N_8759,N_8291,N_8069);
nor U8760 (N_8760,N_8143,N_8148);
nand U8761 (N_8761,N_8201,N_8367);
nor U8762 (N_8762,N_8497,N_8307);
nor U8763 (N_8763,N_8398,N_8317);
nand U8764 (N_8764,N_8391,N_8174);
nor U8765 (N_8765,N_8080,N_8193);
and U8766 (N_8766,N_8224,N_8018);
nor U8767 (N_8767,N_8146,N_8459);
or U8768 (N_8768,N_8193,N_8230);
or U8769 (N_8769,N_8139,N_8279);
nor U8770 (N_8770,N_8020,N_8302);
xnor U8771 (N_8771,N_8044,N_8319);
or U8772 (N_8772,N_8378,N_8227);
nor U8773 (N_8773,N_8082,N_8080);
and U8774 (N_8774,N_8187,N_8471);
nor U8775 (N_8775,N_8098,N_8286);
nor U8776 (N_8776,N_8213,N_8042);
nand U8777 (N_8777,N_8390,N_8002);
or U8778 (N_8778,N_8017,N_8391);
nor U8779 (N_8779,N_8385,N_8216);
nor U8780 (N_8780,N_8112,N_8390);
nor U8781 (N_8781,N_8256,N_8353);
nor U8782 (N_8782,N_8342,N_8104);
and U8783 (N_8783,N_8089,N_8184);
nor U8784 (N_8784,N_8078,N_8334);
nor U8785 (N_8785,N_8406,N_8155);
nand U8786 (N_8786,N_8080,N_8352);
nor U8787 (N_8787,N_8323,N_8246);
nand U8788 (N_8788,N_8295,N_8338);
nand U8789 (N_8789,N_8493,N_8452);
xnor U8790 (N_8790,N_8076,N_8130);
xnor U8791 (N_8791,N_8116,N_8224);
or U8792 (N_8792,N_8171,N_8308);
or U8793 (N_8793,N_8298,N_8137);
nor U8794 (N_8794,N_8384,N_8084);
and U8795 (N_8795,N_8479,N_8378);
nand U8796 (N_8796,N_8263,N_8372);
nand U8797 (N_8797,N_8165,N_8049);
or U8798 (N_8798,N_8276,N_8086);
xnor U8799 (N_8799,N_8060,N_8025);
nand U8800 (N_8800,N_8406,N_8018);
xor U8801 (N_8801,N_8377,N_8205);
or U8802 (N_8802,N_8006,N_8211);
or U8803 (N_8803,N_8164,N_8402);
xor U8804 (N_8804,N_8099,N_8326);
nand U8805 (N_8805,N_8142,N_8126);
nor U8806 (N_8806,N_8424,N_8476);
and U8807 (N_8807,N_8444,N_8222);
and U8808 (N_8808,N_8095,N_8138);
and U8809 (N_8809,N_8015,N_8195);
nand U8810 (N_8810,N_8114,N_8125);
or U8811 (N_8811,N_8385,N_8462);
nor U8812 (N_8812,N_8142,N_8097);
nand U8813 (N_8813,N_8322,N_8466);
nor U8814 (N_8814,N_8144,N_8008);
xor U8815 (N_8815,N_8271,N_8172);
or U8816 (N_8816,N_8421,N_8341);
nor U8817 (N_8817,N_8433,N_8094);
nor U8818 (N_8818,N_8263,N_8248);
nor U8819 (N_8819,N_8331,N_8089);
nand U8820 (N_8820,N_8283,N_8343);
nor U8821 (N_8821,N_8195,N_8057);
and U8822 (N_8822,N_8146,N_8175);
or U8823 (N_8823,N_8264,N_8440);
nand U8824 (N_8824,N_8177,N_8497);
or U8825 (N_8825,N_8484,N_8198);
and U8826 (N_8826,N_8171,N_8130);
nand U8827 (N_8827,N_8152,N_8239);
xnor U8828 (N_8828,N_8479,N_8270);
nand U8829 (N_8829,N_8097,N_8180);
or U8830 (N_8830,N_8309,N_8429);
and U8831 (N_8831,N_8349,N_8063);
nor U8832 (N_8832,N_8092,N_8489);
and U8833 (N_8833,N_8425,N_8061);
or U8834 (N_8834,N_8495,N_8176);
and U8835 (N_8835,N_8140,N_8002);
nor U8836 (N_8836,N_8360,N_8409);
nand U8837 (N_8837,N_8321,N_8185);
xnor U8838 (N_8838,N_8332,N_8276);
nand U8839 (N_8839,N_8180,N_8395);
or U8840 (N_8840,N_8463,N_8050);
or U8841 (N_8841,N_8250,N_8165);
and U8842 (N_8842,N_8384,N_8218);
xor U8843 (N_8843,N_8401,N_8440);
or U8844 (N_8844,N_8401,N_8363);
nor U8845 (N_8845,N_8127,N_8340);
nand U8846 (N_8846,N_8263,N_8074);
nor U8847 (N_8847,N_8053,N_8410);
and U8848 (N_8848,N_8213,N_8496);
xor U8849 (N_8849,N_8067,N_8467);
or U8850 (N_8850,N_8026,N_8209);
or U8851 (N_8851,N_8306,N_8472);
nand U8852 (N_8852,N_8097,N_8246);
nor U8853 (N_8853,N_8364,N_8474);
nand U8854 (N_8854,N_8277,N_8178);
or U8855 (N_8855,N_8163,N_8034);
nor U8856 (N_8856,N_8256,N_8089);
and U8857 (N_8857,N_8136,N_8047);
or U8858 (N_8858,N_8137,N_8223);
or U8859 (N_8859,N_8432,N_8467);
or U8860 (N_8860,N_8182,N_8415);
and U8861 (N_8861,N_8058,N_8152);
nor U8862 (N_8862,N_8270,N_8472);
nand U8863 (N_8863,N_8187,N_8076);
nor U8864 (N_8864,N_8252,N_8270);
nand U8865 (N_8865,N_8080,N_8461);
or U8866 (N_8866,N_8335,N_8307);
and U8867 (N_8867,N_8425,N_8436);
nand U8868 (N_8868,N_8076,N_8073);
nor U8869 (N_8869,N_8308,N_8455);
nand U8870 (N_8870,N_8196,N_8203);
nand U8871 (N_8871,N_8172,N_8171);
or U8872 (N_8872,N_8304,N_8295);
and U8873 (N_8873,N_8282,N_8115);
nor U8874 (N_8874,N_8277,N_8247);
nand U8875 (N_8875,N_8397,N_8094);
and U8876 (N_8876,N_8065,N_8228);
xor U8877 (N_8877,N_8237,N_8388);
or U8878 (N_8878,N_8448,N_8079);
and U8879 (N_8879,N_8079,N_8496);
nor U8880 (N_8880,N_8350,N_8460);
nand U8881 (N_8881,N_8210,N_8387);
xor U8882 (N_8882,N_8145,N_8297);
and U8883 (N_8883,N_8102,N_8211);
and U8884 (N_8884,N_8003,N_8250);
nand U8885 (N_8885,N_8436,N_8234);
or U8886 (N_8886,N_8183,N_8410);
nand U8887 (N_8887,N_8194,N_8491);
or U8888 (N_8888,N_8407,N_8457);
xor U8889 (N_8889,N_8271,N_8103);
or U8890 (N_8890,N_8087,N_8117);
nand U8891 (N_8891,N_8122,N_8490);
nand U8892 (N_8892,N_8113,N_8105);
or U8893 (N_8893,N_8350,N_8060);
or U8894 (N_8894,N_8072,N_8189);
nand U8895 (N_8895,N_8116,N_8260);
nand U8896 (N_8896,N_8000,N_8396);
or U8897 (N_8897,N_8351,N_8110);
xnor U8898 (N_8898,N_8337,N_8006);
xnor U8899 (N_8899,N_8007,N_8122);
nor U8900 (N_8900,N_8414,N_8111);
or U8901 (N_8901,N_8174,N_8067);
or U8902 (N_8902,N_8178,N_8068);
and U8903 (N_8903,N_8143,N_8375);
or U8904 (N_8904,N_8065,N_8218);
nand U8905 (N_8905,N_8260,N_8244);
xnor U8906 (N_8906,N_8154,N_8481);
nor U8907 (N_8907,N_8111,N_8323);
or U8908 (N_8908,N_8315,N_8287);
and U8909 (N_8909,N_8382,N_8108);
and U8910 (N_8910,N_8038,N_8250);
nor U8911 (N_8911,N_8150,N_8415);
xnor U8912 (N_8912,N_8338,N_8488);
nor U8913 (N_8913,N_8416,N_8342);
or U8914 (N_8914,N_8194,N_8237);
nand U8915 (N_8915,N_8167,N_8061);
nor U8916 (N_8916,N_8243,N_8236);
nor U8917 (N_8917,N_8025,N_8140);
nand U8918 (N_8918,N_8252,N_8229);
nand U8919 (N_8919,N_8389,N_8425);
nor U8920 (N_8920,N_8396,N_8460);
xor U8921 (N_8921,N_8159,N_8430);
and U8922 (N_8922,N_8258,N_8102);
nand U8923 (N_8923,N_8468,N_8436);
nand U8924 (N_8924,N_8114,N_8366);
nand U8925 (N_8925,N_8464,N_8370);
or U8926 (N_8926,N_8414,N_8328);
or U8927 (N_8927,N_8153,N_8086);
nand U8928 (N_8928,N_8494,N_8319);
and U8929 (N_8929,N_8480,N_8238);
or U8930 (N_8930,N_8291,N_8295);
nor U8931 (N_8931,N_8210,N_8348);
or U8932 (N_8932,N_8051,N_8463);
and U8933 (N_8933,N_8478,N_8359);
and U8934 (N_8934,N_8440,N_8289);
nor U8935 (N_8935,N_8048,N_8290);
and U8936 (N_8936,N_8245,N_8361);
nand U8937 (N_8937,N_8215,N_8250);
or U8938 (N_8938,N_8197,N_8265);
nor U8939 (N_8939,N_8324,N_8329);
nor U8940 (N_8940,N_8018,N_8422);
or U8941 (N_8941,N_8305,N_8155);
or U8942 (N_8942,N_8068,N_8410);
nor U8943 (N_8943,N_8005,N_8192);
nor U8944 (N_8944,N_8044,N_8202);
and U8945 (N_8945,N_8443,N_8248);
nand U8946 (N_8946,N_8252,N_8187);
nor U8947 (N_8947,N_8383,N_8032);
or U8948 (N_8948,N_8101,N_8141);
and U8949 (N_8949,N_8340,N_8083);
or U8950 (N_8950,N_8225,N_8161);
xor U8951 (N_8951,N_8034,N_8289);
nor U8952 (N_8952,N_8091,N_8438);
and U8953 (N_8953,N_8390,N_8343);
nand U8954 (N_8954,N_8186,N_8441);
nand U8955 (N_8955,N_8097,N_8120);
and U8956 (N_8956,N_8017,N_8250);
nand U8957 (N_8957,N_8458,N_8199);
and U8958 (N_8958,N_8372,N_8052);
nor U8959 (N_8959,N_8433,N_8049);
nor U8960 (N_8960,N_8489,N_8369);
or U8961 (N_8961,N_8028,N_8285);
nor U8962 (N_8962,N_8169,N_8481);
or U8963 (N_8963,N_8242,N_8306);
nor U8964 (N_8964,N_8278,N_8273);
and U8965 (N_8965,N_8270,N_8262);
or U8966 (N_8966,N_8201,N_8379);
xnor U8967 (N_8967,N_8107,N_8007);
and U8968 (N_8968,N_8228,N_8135);
nor U8969 (N_8969,N_8469,N_8334);
nand U8970 (N_8970,N_8012,N_8165);
and U8971 (N_8971,N_8070,N_8359);
or U8972 (N_8972,N_8477,N_8061);
nand U8973 (N_8973,N_8082,N_8010);
and U8974 (N_8974,N_8069,N_8449);
or U8975 (N_8975,N_8493,N_8319);
nor U8976 (N_8976,N_8354,N_8044);
nand U8977 (N_8977,N_8325,N_8490);
xnor U8978 (N_8978,N_8190,N_8340);
or U8979 (N_8979,N_8405,N_8022);
nor U8980 (N_8980,N_8356,N_8365);
or U8981 (N_8981,N_8179,N_8045);
nand U8982 (N_8982,N_8107,N_8203);
nor U8983 (N_8983,N_8379,N_8089);
or U8984 (N_8984,N_8248,N_8160);
nor U8985 (N_8985,N_8406,N_8474);
nand U8986 (N_8986,N_8476,N_8092);
nor U8987 (N_8987,N_8448,N_8440);
nor U8988 (N_8988,N_8309,N_8096);
and U8989 (N_8989,N_8178,N_8238);
nand U8990 (N_8990,N_8300,N_8063);
and U8991 (N_8991,N_8037,N_8277);
and U8992 (N_8992,N_8148,N_8080);
or U8993 (N_8993,N_8153,N_8014);
nand U8994 (N_8994,N_8173,N_8287);
or U8995 (N_8995,N_8330,N_8443);
nor U8996 (N_8996,N_8273,N_8064);
xnor U8997 (N_8997,N_8139,N_8474);
nand U8998 (N_8998,N_8281,N_8279);
and U8999 (N_8999,N_8447,N_8300);
nand U9000 (N_9000,N_8676,N_8592);
or U9001 (N_9001,N_8680,N_8994);
nor U9002 (N_9002,N_8836,N_8510);
or U9003 (N_9003,N_8565,N_8528);
nor U9004 (N_9004,N_8767,N_8660);
nor U9005 (N_9005,N_8538,N_8533);
nand U9006 (N_9006,N_8876,N_8991);
or U9007 (N_9007,N_8539,N_8606);
and U9008 (N_9008,N_8916,N_8535);
and U9009 (N_9009,N_8794,N_8973);
and U9010 (N_9010,N_8590,N_8752);
or U9011 (N_9011,N_8632,N_8785);
nand U9012 (N_9012,N_8749,N_8748);
or U9013 (N_9013,N_8883,N_8503);
and U9014 (N_9014,N_8620,N_8781);
nor U9015 (N_9015,N_8512,N_8703);
and U9016 (N_9016,N_8722,N_8837);
nand U9017 (N_9017,N_8677,N_8868);
nor U9018 (N_9018,N_8804,N_8736);
nand U9019 (N_9019,N_8627,N_8926);
nand U9020 (N_9020,N_8754,N_8980);
and U9021 (N_9021,N_8835,N_8936);
xnor U9022 (N_9022,N_8910,N_8981);
and U9023 (N_9023,N_8745,N_8901);
nor U9024 (N_9024,N_8937,N_8576);
and U9025 (N_9025,N_8733,N_8791);
nor U9026 (N_9026,N_8775,N_8738);
nor U9027 (N_9027,N_8704,N_8674);
nand U9028 (N_9028,N_8848,N_8999);
or U9029 (N_9029,N_8502,N_8721);
nor U9030 (N_9030,N_8692,N_8955);
and U9031 (N_9031,N_8633,N_8894);
xnor U9032 (N_9032,N_8905,N_8734);
nand U9033 (N_9033,N_8712,N_8800);
and U9034 (N_9034,N_8558,N_8619);
nand U9035 (N_9035,N_8669,N_8945);
nor U9036 (N_9036,N_8758,N_8623);
nand U9037 (N_9037,N_8621,N_8751);
nor U9038 (N_9038,N_8851,N_8789);
or U9039 (N_9039,N_8922,N_8650);
or U9040 (N_9040,N_8562,N_8971);
and U9041 (N_9041,N_8902,N_8671);
or U9042 (N_9042,N_8543,N_8885);
and U9043 (N_9043,N_8824,N_8879);
nor U9044 (N_9044,N_8717,N_8920);
xor U9045 (N_9045,N_8846,N_8839);
xnor U9046 (N_9046,N_8730,N_8747);
or U9047 (N_9047,N_8770,N_8521);
or U9048 (N_9048,N_8607,N_8665);
nand U9049 (N_9049,N_8988,N_8811);
and U9050 (N_9050,N_8634,N_8954);
nor U9051 (N_9051,N_8656,N_8821);
or U9052 (N_9052,N_8854,N_8556);
nor U9053 (N_9053,N_8643,N_8690);
nand U9054 (N_9054,N_8630,N_8777);
xnor U9055 (N_9055,N_8881,N_8959);
or U9056 (N_9056,N_8915,N_8519);
nor U9057 (N_9057,N_8731,N_8649);
nand U9058 (N_9058,N_8699,N_8688);
nor U9059 (N_9059,N_8501,N_8909);
and U9060 (N_9060,N_8581,N_8628);
or U9061 (N_9061,N_8817,N_8641);
nor U9062 (N_9062,N_8939,N_8983);
or U9063 (N_9063,N_8530,N_8842);
or U9064 (N_9064,N_8525,N_8697);
and U9065 (N_9065,N_8657,N_8853);
xor U9066 (N_9066,N_8829,N_8892);
and U9067 (N_9067,N_8517,N_8993);
nor U9068 (N_9068,N_8838,N_8976);
xor U9069 (N_9069,N_8647,N_8832);
nand U9070 (N_9070,N_8571,N_8640);
or U9071 (N_9071,N_8813,N_8584);
and U9072 (N_9072,N_8707,N_8865);
xor U9073 (N_9073,N_8998,N_8808);
xor U9074 (N_9074,N_8918,N_8589);
nor U9075 (N_9075,N_8977,N_8522);
nor U9076 (N_9076,N_8534,N_8953);
and U9077 (N_9077,N_8867,N_8552);
nand U9078 (N_9078,N_8984,N_8694);
and U9079 (N_9079,N_8756,N_8615);
xor U9080 (N_9080,N_8764,N_8626);
nor U9081 (N_9081,N_8900,N_8588);
and U9082 (N_9082,N_8520,N_8871);
nor U9083 (N_9083,N_8548,N_8689);
and U9084 (N_9084,N_8924,N_8792);
or U9085 (N_9085,N_8812,N_8931);
nand U9086 (N_9086,N_8594,N_8618);
nor U9087 (N_9087,N_8899,N_8595);
and U9088 (N_9088,N_8750,N_8889);
or U9089 (N_9089,N_8516,N_8617);
nand U9090 (N_9090,N_8890,N_8536);
nor U9091 (N_9091,N_8989,N_8573);
and U9092 (N_9092,N_8771,N_8961);
or U9093 (N_9093,N_8996,N_8819);
nand U9094 (N_9094,N_8670,N_8833);
or U9095 (N_9095,N_8695,N_8687);
and U9096 (N_9096,N_8629,N_8965);
nand U9097 (N_9097,N_8579,N_8739);
and U9098 (N_9098,N_8608,N_8672);
nand U9099 (N_9099,N_8952,N_8526);
and U9100 (N_9100,N_8639,N_8978);
xor U9101 (N_9101,N_8511,N_8946);
nor U9102 (N_9102,N_8898,N_8719);
nor U9103 (N_9103,N_8743,N_8822);
or U9104 (N_9104,N_8863,N_8716);
and U9105 (N_9105,N_8951,N_8872);
xor U9106 (N_9106,N_8875,N_8551);
nor U9107 (N_9107,N_8787,N_8841);
or U9108 (N_9108,N_8663,N_8682);
nor U9109 (N_9109,N_8960,N_8807);
and U9110 (N_9110,N_8818,N_8948);
and U9111 (N_9111,N_8500,N_8570);
or U9112 (N_9112,N_8642,N_8801);
and U9113 (N_9113,N_8648,N_8893);
and U9114 (N_9114,N_8995,N_8675);
nand U9115 (N_9115,N_8577,N_8602);
and U9116 (N_9116,N_8788,N_8609);
and U9117 (N_9117,N_8659,N_8917);
nor U9118 (N_9118,N_8840,N_8509);
and U9119 (N_9119,N_8599,N_8987);
nand U9120 (N_9120,N_8715,N_8852);
or U9121 (N_9121,N_8685,N_8887);
and U9122 (N_9122,N_8776,N_8985);
or U9123 (N_9123,N_8843,N_8969);
or U9124 (N_9124,N_8825,N_8966);
or U9125 (N_9125,N_8857,N_8856);
xnor U9126 (N_9126,N_8666,N_8907);
or U9127 (N_9127,N_8698,N_8759);
or U9128 (N_9128,N_8904,N_8944);
or U9129 (N_9129,N_8831,N_8653);
nand U9130 (N_9130,N_8796,N_8933);
xor U9131 (N_9131,N_8683,N_8782);
or U9132 (N_9132,N_8964,N_8555);
or U9133 (N_9133,N_8744,N_8919);
nand U9134 (N_9134,N_8979,N_8932);
and U9135 (N_9135,N_8550,N_8823);
nand U9136 (N_9136,N_8596,N_8622);
or U9137 (N_9137,N_8802,N_8869);
or U9138 (N_9138,N_8566,N_8803);
nor U9139 (N_9139,N_8700,N_8601);
nand U9140 (N_9140,N_8947,N_8508);
nand U9141 (N_9141,N_8827,N_8962);
nor U9142 (N_9142,N_8949,N_8970);
nor U9143 (N_9143,N_8578,N_8805);
and U9144 (N_9144,N_8927,N_8631);
or U9145 (N_9145,N_8661,N_8956);
nor U9146 (N_9146,N_8810,N_8725);
nor U9147 (N_9147,N_8547,N_8652);
nand U9148 (N_9148,N_8798,N_8524);
or U9149 (N_9149,N_8815,N_8681);
nor U9150 (N_9150,N_8740,N_8709);
and U9151 (N_9151,N_8742,N_8720);
or U9152 (N_9152,N_8702,N_8580);
or U9153 (N_9153,N_8678,N_8799);
xnor U9154 (N_9154,N_8943,N_8616);
and U9155 (N_9155,N_8772,N_8705);
and U9156 (N_9156,N_8532,N_8784);
or U9157 (N_9157,N_8968,N_8816);
and U9158 (N_9158,N_8724,N_8963);
or U9159 (N_9159,N_8941,N_8515);
nor U9160 (N_9160,N_8612,N_8549);
or U9161 (N_9161,N_8507,N_8793);
nor U9162 (N_9162,N_8884,N_8760);
or U9163 (N_9163,N_8711,N_8611);
and U9164 (N_9164,N_8940,N_8809);
and U9165 (N_9165,N_8928,N_8790);
and U9166 (N_9166,N_8997,N_8847);
nand U9167 (N_9167,N_8912,N_8934);
and U9168 (N_9168,N_8625,N_8614);
xnor U9169 (N_9169,N_8529,N_8726);
or U9170 (N_9170,N_8882,N_8654);
and U9171 (N_9171,N_8828,N_8982);
and U9172 (N_9172,N_8975,N_8553);
nand U9173 (N_9173,N_8575,N_8950);
nor U9174 (N_9174,N_8561,N_8701);
or U9175 (N_9175,N_8753,N_8765);
nand U9176 (N_9176,N_8582,N_8723);
nor U9177 (N_9177,N_8880,N_8518);
nor U9178 (N_9178,N_8544,N_8768);
and U9179 (N_9179,N_8877,N_8583);
or U9180 (N_9180,N_8870,N_8860);
xor U9181 (N_9181,N_8990,N_8859);
nor U9182 (N_9182,N_8929,N_8773);
nand U9183 (N_9183,N_8598,N_8537);
and U9184 (N_9184,N_8605,N_8651);
nor U9185 (N_9185,N_8906,N_8914);
nand U9186 (N_9186,N_8858,N_8957);
nand U9187 (N_9187,N_8942,N_8911);
xnor U9188 (N_9188,N_8644,N_8673);
xor U9189 (N_9189,N_8779,N_8664);
or U9190 (N_9190,N_8523,N_8729);
nor U9191 (N_9191,N_8714,N_8992);
xnor U9192 (N_9192,N_8826,N_8593);
or U9193 (N_9193,N_8545,N_8585);
nand U9194 (N_9194,N_8541,N_8693);
or U9195 (N_9195,N_8958,N_8527);
nor U9196 (N_9196,N_8667,N_8814);
xor U9197 (N_9197,N_8830,N_8967);
nor U9198 (N_9198,N_8986,N_8774);
nand U9199 (N_9199,N_8591,N_8786);
xor U9200 (N_9200,N_8741,N_8554);
and U9201 (N_9201,N_8886,N_8710);
nor U9202 (N_9202,N_8780,N_8624);
and U9203 (N_9203,N_8713,N_8938);
or U9204 (N_9204,N_8806,N_8797);
xnor U9205 (N_9205,N_8874,N_8557);
or U9206 (N_9206,N_8897,N_8610);
nor U9207 (N_9207,N_8923,N_8896);
nand U9208 (N_9208,N_8604,N_8861);
nor U9209 (N_9209,N_8844,N_8560);
nand U9210 (N_9210,N_8888,N_8567);
or U9211 (N_9211,N_8795,N_8913);
xor U9212 (N_9212,N_8696,N_8762);
nand U9213 (N_9213,N_8864,N_8766);
and U9214 (N_9214,N_8925,N_8646);
nor U9215 (N_9215,N_8757,N_8662);
nand U9216 (N_9216,N_8668,N_8728);
nor U9217 (N_9217,N_8587,N_8542);
nand U9218 (N_9218,N_8635,N_8679);
nor U9219 (N_9219,N_8862,N_8572);
nor U9220 (N_9220,N_8645,N_8873);
nor U9221 (N_9221,N_8531,N_8755);
or U9222 (N_9222,N_8563,N_8658);
nor U9223 (N_9223,N_8866,N_8638);
nor U9224 (N_9224,N_8908,N_8540);
nor U9225 (N_9225,N_8569,N_8735);
nand U9226 (N_9226,N_8513,N_8834);
nand U9227 (N_9227,N_8691,N_8974);
and U9228 (N_9228,N_8769,N_8783);
or U9229 (N_9229,N_8505,N_8600);
or U9230 (N_9230,N_8574,N_8737);
and U9231 (N_9231,N_8546,N_8891);
or U9232 (N_9232,N_8636,N_8506);
or U9233 (N_9233,N_8706,N_8849);
and U9234 (N_9234,N_8686,N_8763);
and U9235 (N_9235,N_8718,N_8514);
nor U9236 (N_9236,N_8586,N_8568);
nand U9237 (N_9237,N_8597,N_8935);
or U9238 (N_9238,N_8850,N_8921);
nand U9239 (N_9239,N_8564,N_8732);
and U9240 (N_9240,N_8820,N_8559);
nand U9241 (N_9241,N_8855,N_8708);
and U9242 (N_9242,N_8504,N_8727);
nand U9243 (N_9243,N_8972,N_8761);
nor U9244 (N_9244,N_8878,N_8930);
nor U9245 (N_9245,N_8613,N_8845);
nand U9246 (N_9246,N_8746,N_8778);
nand U9247 (N_9247,N_8903,N_8603);
and U9248 (N_9248,N_8637,N_8655);
nor U9249 (N_9249,N_8684,N_8895);
nor U9250 (N_9250,N_8595,N_8515);
and U9251 (N_9251,N_8690,N_8627);
nand U9252 (N_9252,N_8636,N_8508);
and U9253 (N_9253,N_8906,N_8883);
xor U9254 (N_9254,N_8714,N_8993);
or U9255 (N_9255,N_8504,N_8679);
or U9256 (N_9256,N_8645,N_8868);
nor U9257 (N_9257,N_8817,N_8992);
nand U9258 (N_9258,N_8653,N_8846);
nand U9259 (N_9259,N_8525,N_8961);
and U9260 (N_9260,N_8841,N_8734);
nand U9261 (N_9261,N_8853,N_8621);
xor U9262 (N_9262,N_8502,N_8999);
nor U9263 (N_9263,N_8946,N_8954);
and U9264 (N_9264,N_8972,N_8828);
xnor U9265 (N_9265,N_8721,N_8910);
and U9266 (N_9266,N_8801,N_8563);
and U9267 (N_9267,N_8670,N_8582);
nand U9268 (N_9268,N_8717,N_8784);
nand U9269 (N_9269,N_8828,N_8913);
or U9270 (N_9270,N_8947,N_8807);
nand U9271 (N_9271,N_8746,N_8863);
xor U9272 (N_9272,N_8767,N_8648);
and U9273 (N_9273,N_8903,N_8676);
nand U9274 (N_9274,N_8941,N_8855);
nand U9275 (N_9275,N_8739,N_8640);
and U9276 (N_9276,N_8646,N_8683);
nand U9277 (N_9277,N_8656,N_8503);
nand U9278 (N_9278,N_8989,N_8784);
or U9279 (N_9279,N_8957,N_8970);
nor U9280 (N_9280,N_8975,N_8755);
xnor U9281 (N_9281,N_8609,N_8703);
or U9282 (N_9282,N_8800,N_8638);
nor U9283 (N_9283,N_8879,N_8974);
or U9284 (N_9284,N_8832,N_8616);
or U9285 (N_9285,N_8851,N_8762);
nor U9286 (N_9286,N_8850,N_8843);
and U9287 (N_9287,N_8517,N_8723);
nor U9288 (N_9288,N_8811,N_8517);
nor U9289 (N_9289,N_8670,N_8935);
nor U9290 (N_9290,N_8631,N_8868);
or U9291 (N_9291,N_8559,N_8743);
or U9292 (N_9292,N_8621,N_8511);
nor U9293 (N_9293,N_8927,N_8655);
xor U9294 (N_9294,N_8994,N_8527);
or U9295 (N_9295,N_8735,N_8653);
or U9296 (N_9296,N_8816,N_8912);
and U9297 (N_9297,N_8648,N_8652);
nand U9298 (N_9298,N_8758,N_8842);
nand U9299 (N_9299,N_8560,N_8715);
and U9300 (N_9300,N_8738,N_8502);
xor U9301 (N_9301,N_8562,N_8779);
nor U9302 (N_9302,N_8860,N_8676);
and U9303 (N_9303,N_8807,N_8661);
and U9304 (N_9304,N_8731,N_8777);
or U9305 (N_9305,N_8848,N_8623);
xnor U9306 (N_9306,N_8505,N_8654);
nand U9307 (N_9307,N_8882,N_8768);
and U9308 (N_9308,N_8526,N_8885);
nand U9309 (N_9309,N_8786,N_8998);
nand U9310 (N_9310,N_8547,N_8561);
nand U9311 (N_9311,N_8711,N_8552);
nand U9312 (N_9312,N_8783,N_8778);
xor U9313 (N_9313,N_8709,N_8704);
xor U9314 (N_9314,N_8636,N_8625);
nand U9315 (N_9315,N_8816,N_8550);
nand U9316 (N_9316,N_8620,N_8550);
nor U9317 (N_9317,N_8936,N_8519);
or U9318 (N_9318,N_8712,N_8582);
or U9319 (N_9319,N_8794,N_8578);
xnor U9320 (N_9320,N_8600,N_8856);
nand U9321 (N_9321,N_8641,N_8917);
nor U9322 (N_9322,N_8974,N_8617);
xnor U9323 (N_9323,N_8519,N_8920);
nand U9324 (N_9324,N_8849,N_8726);
nor U9325 (N_9325,N_8778,N_8700);
and U9326 (N_9326,N_8738,N_8809);
and U9327 (N_9327,N_8677,N_8983);
nand U9328 (N_9328,N_8704,N_8731);
and U9329 (N_9329,N_8775,N_8666);
nand U9330 (N_9330,N_8988,N_8886);
xor U9331 (N_9331,N_8703,N_8810);
nand U9332 (N_9332,N_8898,N_8676);
and U9333 (N_9333,N_8704,N_8857);
nor U9334 (N_9334,N_8889,N_8789);
or U9335 (N_9335,N_8521,N_8563);
nand U9336 (N_9336,N_8969,N_8566);
xnor U9337 (N_9337,N_8852,N_8599);
or U9338 (N_9338,N_8919,N_8932);
xor U9339 (N_9339,N_8506,N_8722);
and U9340 (N_9340,N_8749,N_8956);
nand U9341 (N_9341,N_8979,N_8850);
xnor U9342 (N_9342,N_8977,N_8798);
nand U9343 (N_9343,N_8658,N_8844);
nand U9344 (N_9344,N_8664,N_8851);
nand U9345 (N_9345,N_8719,N_8866);
and U9346 (N_9346,N_8696,N_8516);
nor U9347 (N_9347,N_8570,N_8598);
or U9348 (N_9348,N_8939,N_8649);
nor U9349 (N_9349,N_8612,N_8954);
or U9350 (N_9350,N_8596,N_8666);
nor U9351 (N_9351,N_8711,N_8736);
and U9352 (N_9352,N_8644,N_8757);
nor U9353 (N_9353,N_8827,N_8505);
and U9354 (N_9354,N_8905,N_8644);
and U9355 (N_9355,N_8722,N_8988);
or U9356 (N_9356,N_8760,N_8543);
and U9357 (N_9357,N_8790,N_8541);
nor U9358 (N_9358,N_8930,N_8879);
or U9359 (N_9359,N_8592,N_8718);
and U9360 (N_9360,N_8626,N_8686);
nand U9361 (N_9361,N_8803,N_8898);
nand U9362 (N_9362,N_8790,N_8971);
or U9363 (N_9363,N_8778,N_8589);
xor U9364 (N_9364,N_8691,N_8699);
xnor U9365 (N_9365,N_8829,N_8898);
and U9366 (N_9366,N_8959,N_8625);
nor U9367 (N_9367,N_8827,N_8891);
or U9368 (N_9368,N_8923,N_8965);
and U9369 (N_9369,N_8529,N_8944);
and U9370 (N_9370,N_8716,N_8544);
nand U9371 (N_9371,N_8555,N_8972);
nor U9372 (N_9372,N_8651,N_8589);
and U9373 (N_9373,N_8747,N_8797);
and U9374 (N_9374,N_8995,N_8898);
or U9375 (N_9375,N_8735,N_8860);
and U9376 (N_9376,N_8587,N_8907);
xor U9377 (N_9377,N_8514,N_8756);
nand U9378 (N_9378,N_8547,N_8888);
nor U9379 (N_9379,N_8830,N_8644);
and U9380 (N_9380,N_8807,N_8799);
nand U9381 (N_9381,N_8694,N_8769);
nor U9382 (N_9382,N_8661,N_8853);
or U9383 (N_9383,N_8901,N_8667);
and U9384 (N_9384,N_8586,N_8783);
nand U9385 (N_9385,N_8645,N_8656);
and U9386 (N_9386,N_8908,N_8902);
xnor U9387 (N_9387,N_8839,N_8503);
nand U9388 (N_9388,N_8748,N_8519);
xnor U9389 (N_9389,N_8978,N_8631);
xnor U9390 (N_9390,N_8723,N_8962);
nand U9391 (N_9391,N_8523,N_8904);
and U9392 (N_9392,N_8568,N_8922);
nand U9393 (N_9393,N_8970,N_8959);
nor U9394 (N_9394,N_8915,N_8969);
or U9395 (N_9395,N_8615,N_8858);
and U9396 (N_9396,N_8871,N_8539);
and U9397 (N_9397,N_8543,N_8514);
nor U9398 (N_9398,N_8924,N_8591);
nor U9399 (N_9399,N_8848,N_8945);
or U9400 (N_9400,N_8567,N_8670);
or U9401 (N_9401,N_8957,N_8767);
nand U9402 (N_9402,N_8585,N_8717);
and U9403 (N_9403,N_8908,N_8826);
xor U9404 (N_9404,N_8589,N_8648);
nand U9405 (N_9405,N_8634,N_8643);
or U9406 (N_9406,N_8997,N_8852);
xnor U9407 (N_9407,N_8985,N_8894);
nor U9408 (N_9408,N_8633,N_8582);
nand U9409 (N_9409,N_8635,N_8899);
or U9410 (N_9410,N_8711,N_8526);
nand U9411 (N_9411,N_8581,N_8739);
or U9412 (N_9412,N_8977,N_8674);
and U9413 (N_9413,N_8506,N_8585);
nand U9414 (N_9414,N_8783,N_8963);
nor U9415 (N_9415,N_8625,N_8635);
or U9416 (N_9416,N_8745,N_8968);
and U9417 (N_9417,N_8761,N_8826);
nand U9418 (N_9418,N_8707,N_8902);
nand U9419 (N_9419,N_8824,N_8548);
nor U9420 (N_9420,N_8568,N_8526);
and U9421 (N_9421,N_8559,N_8764);
and U9422 (N_9422,N_8780,N_8626);
or U9423 (N_9423,N_8902,N_8941);
nand U9424 (N_9424,N_8666,N_8737);
or U9425 (N_9425,N_8708,N_8921);
and U9426 (N_9426,N_8717,N_8710);
xnor U9427 (N_9427,N_8942,N_8695);
nor U9428 (N_9428,N_8829,N_8555);
nor U9429 (N_9429,N_8917,N_8999);
and U9430 (N_9430,N_8688,N_8760);
and U9431 (N_9431,N_8784,N_8823);
or U9432 (N_9432,N_8925,N_8723);
nor U9433 (N_9433,N_8523,N_8763);
and U9434 (N_9434,N_8782,N_8857);
xnor U9435 (N_9435,N_8577,N_8786);
nor U9436 (N_9436,N_8772,N_8830);
and U9437 (N_9437,N_8802,N_8537);
xnor U9438 (N_9438,N_8543,N_8907);
nor U9439 (N_9439,N_8693,N_8799);
and U9440 (N_9440,N_8855,N_8673);
nand U9441 (N_9441,N_8738,N_8699);
nor U9442 (N_9442,N_8968,N_8609);
and U9443 (N_9443,N_8509,N_8899);
xnor U9444 (N_9444,N_8990,N_8807);
or U9445 (N_9445,N_8742,N_8643);
or U9446 (N_9446,N_8585,N_8570);
nor U9447 (N_9447,N_8674,N_8884);
nor U9448 (N_9448,N_8641,N_8742);
nor U9449 (N_9449,N_8744,N_8532);
and U9450 (N_9450,N_8959,N_8624);
nor U9451 (N_9451,N_8648,N_8912);
nand U9452 (N_9452,N_8624,N_8639);
and U9453 (N_9453,N_8776,N_8740);
or U9454 (N_9454,N_8534,N_8765);
or U9455 (N_9455,N_8683,N_8698);
nor U9456 (N_9456,N_8617,N_8648);
or U9457 (N_9457,N_8868,N_8555);
nor U9458 (N_9458,N_8504,N_8799);
or U9459 (N_9459,N_8862,N_8767);
and U9460 (N_9460,N_8572,N_8939);
and U9461 (N_9461,N_8752,N_8706);
nand U9462 (N_9462,N_8745,N_8641);
and U9463 (N_9463,N_8665,N_8600);
xnor U9464 (N_9464,N_8983,N_8783);
and U9465 (N_9465,N_8559,N_8966);
xor U9466 (N_9466,N_8572,N_8871);
nor U9467 (N_9467,N_8946,N_8890);
and U9468 (N_9468,N_8530,N_8841);
nor U9469 (N_9469,N_8993,N_8903);
nor U9470 (N_9470,N_8528,N_8858);
nor U9471 (N_9471,N_8851,N_8542);
nor U9472 (N_9472,N_8753,N_8951);
nand U9473 (N_9473,N_8754,N_8886);
xnor U9474 (N_9474,N_8741,N_8634);
and U9475 (N_9475,N_8856,N_8678);
and U9476 (N_9476,N_8582,N_8541);
nand U9477 (N_9477,N_8995,N_8633);
or U9478 (N_9478,N_8906,N_8564);
or U9479 (N_9479,N_8971,N_8816);
nor U9480 (N_9480,N_8805,N_8604);
or U9481 (N_9481,N_8582,N_8584);
nand U9482 (N_9482,N_8574,N_8548);
nor U9483 (N_9483,N_8710,N_8540);
and U9484 (N_9484,N_8522,N_8931);
nor U9485 (N_9485,N_8717,N_8805);
nand U9486 (N_9486,N_8782,N_8952);
nor U9487 (N_9487,N_8762,N_8855);
nand U9488 (N_9488,N_8734,N_8800);
nor U9489 (N_9489,N_8635,N_8882);
xnor U9490 (N_9490,N_8611,N_8686);
nor U9491 (N_9491,N_8854,N_8591);
xor U9492 (N_9492,N_8994,N_8579);
and U9493 (N_9493,N_8673,N_8916);
or U9494 (N_9494,N_8670,N_8715);
nand U9495 (N_9495,N_8944,N_8876);
nor U9496 (N_9496,N_8754,N_8772);
xor U9497 (N_9497,N_8688,N_8531);
xnor U9498 (N_9498,N_8704,N_8978);
nand U9499 (N_9499,N_8742,N_8743);
nand U9500 (N_9500,N_9240,N_9449);
xor U9501 (N_9501,N_9007,N_9006);
nand U9502 (N_9502,N_9104,N_9019);
or U9503 (N_9503,N_9096,N_9044);
or U9504 (N_9504,N_9027,N_9308);
and U9505 (N_9505,N_9169,N_9424);
or U9506 (N_9506,N_9099,N_9213);
xnor U9507 (N_9507,N_9369,N_9325);
nor U9508 (N_9508,N_9060,N_9314);
nand U9509 (N_9509,N_9273,N_9095);
and U9510 (N_9510,N_9335,N_9394);
nand U9511 (N_9511,N_9079,N_9408);
or U9512 (N_9512,N_9397,N_9038);
nor U9513 (N_9513,N_9320,N_9256);
nand U9514 (N_9514,N_9339,N_9439);
or U9515 (N_9515,N_9464,N_9321);
and U9516 (N_9516,N_9187,N_9153);
and U9517 (N_9517,N_9102,N_9221);
nor U9518 (N_9518,N_9289,N_9459);
nor U9519 (N_9519,N_9119,N_9300);
nor U9520 (N_9520,N_9302,N_9171);
and U9521 (N_9521,N_9114,N_9090);
nor U9522 (N_9522,N_9233,N_9245);
nand U9523 (N_9523,N_9117,N_9043);
nand U9524 (N_9524,N_9155,N_9101);
nor U9525 (N_9525,N_9278,N_9107);
nor U9526 (N_9526,N_9462,N_9016);
nand U9527 (N_9527,N_9146,N_9175);
nor U9528 (N_9528,N_9026,N_9342);
nor U9529 (N_9529,N_9264,N_9124);
or U9530 (N_9530,N_9077,N_9242);
xor U9531 (N_9531,N_9253,N_9094);
xor U9532 (N_9532,N_9133,N_9196);
or U9533 (N_9533,N_9160,N_9219);
nor U9534 (N_9534,N_9283,N_9235);
nand U9535 (N_9535,N_9103,N_9398);
nand U9536 (N_9536,N_9429,N_9334);
and U9537 (N_9537,N_9034,N_9435);
nand U9538 (N_9538,N_9154,N_9494);
nand U9539 (N_9539,N_9017,N_9159);
and U9540 (N_9540,N_9474,N_9396);
nand U9541 (N_9541,N_9036,N_9176);
or U9542 (N_9542,N_9121,N_9150);
or U9543 (N_9543,N_9358,N_9493);
and U9544 (N_9544,N_9041,N_9333);
nor U9545 (N_9545,N_9267,N_9002);
xnor U9546 (N_9546,N_9450,N_9265);
and U9547 (N_9547,N_9152,N_9147);
and U9548 (N_9548,N_9414,N_9310);
nor U9549 (N_9549,N_9499,N_9349);
nor U9550 (N_9550,N_9243,N_9456);
nand U9551 (N_9551,N_9033,N_9475);
nor U9552 (N_9552,N_9063,N_9372);
and U9553 (N_9553,N_9151,N_9357);
or U9554 (N_9554,N_9307,N_9177);
or U9555 (N_9555,N_9422,N_9336);
nor U9556 (N_9556,N_9074,N_9049);
and U9557 (N_9557,N_9269,N_9042);
xnor U9558 (N_9558,N_9228,N_9092);
and U9559 (N_9559,N_9488,N_9292);
nor U9560 (N_9560,N_9113,N_9483);
xnor U9561 (N_9561,N_9317,N_9251);
nand U9562 (N_9562,N_9409,N_9427);
nand U9563 (N_9563,N_9337,N_9201);
xnor U9564 (N_9564,N_9197,N_9445);
or U9565 (N_9565,N_9178,N_9039);
nor U9566 (N_9566,N_9384,N_9270);
nand U9567 (N_9567,N_9353,N_9469);
nand U9568 (N_9568,N_9471,N_9305);
xnor U9569 (N_9569,N_9073,N_9188);
or U9570 (N_9570,N_9425,N_9135);
or U9571 (N_9571,N_9365,N_9131);
nor U9572 (N_9572,N_9272,N_9056);
and U9573 (N_9573,N_9089,N_9141);
nor U9574 (N_9574,N_9489,N_9360);
nand U9575 (N_9575,N_9066,N_9401);
xor U9576 (N_9576,N_9008,N_9029);
nor U9577 (N_9577,N_9127,N_9189);
or U9578 (N_9578,N_9013,N_9247);
nor U9579 (N_9579,N_9014,N_9323);
and U9580 (N_9580,N_9004,N_9476);
nand U9581 (N_9581,N_9291,N_9313);
nand U9582 (N_9582,N_9037,N_9279);
and U9583 (N_9583,N_9340,N_9120);
or U9584 (N_9584,N_9125,N_9479);
and U9585 (N_9585,N_9416,N_9181);
or U9586 (N_9586,N_9254,N_9454);
xor U9587 (N_9587,N_9343,N_9156);
or U9588 (N_9588,N_9093,N_9434);
and U9589 (N_9589,N_9136,N_9129);
and U9590 (N_9590,N_9072,N_9182);
nor U9591 (N_9591,N_9405,N_9229);
nor U9592 (N_9592,N_9382,N_9379);
or U9593 (N_9593,N_9438,N_9238);
nand U9594 (N_9594,N_9012,N_9210);
or U9595 (N_9595,N_9170,N_9106);
nor U9596 (N_9596,N_9164,N_9123);
and U9597 (N_9597,N_9330,N_9359);
xor U9598 (N_9598,N_9158,N_9194);
and U9599 (N_9599,N_9259,N_9260);
or U9600 (N_9600,N_9311,N_9443);
and U9601 (N_9601,N_9419,N_9352);
nor U9602 (N_9602,N_9485,N_9491);
or U9603 (N_9603,N_9068,N_9185);
or U9604 (N_9604,N_9395,N_9461);
and U9605 (N_9605,N_9070,N_9148);
and U9606 (N_9606,N_9137,N_9216);
nand U9607 (N_9607,N_9436,N_9391);
nor U9608 (N_9608,N_9015,N_9220);
nand U9609 (N_9609,N_9234,N_9457);
nand U9610 (N_9610,N_9287,N_9071);
nor U9611 (N_9611,N_9028,N_9258);
nand U9612 (N_9612,N_9318,N_9306);
nor U9613 (N_9613,N_9297,N_9458);
nor U9614 (N_9614,N_9275,N_9055);
and U9615 (N_9615,N_9288,N_9341);
and U9616 (N_9616,N_9040,N_9115);
or U9617 (N_9617,N_9277,N_9246);
xnor U9618 (N_9618,N_9091,N_9322);
and U9619 (N_9619,N_9466,N_9385);
nor U9620 (N_9620,N_9280,N_9168);
nor U9621 (N_9621,N_9215,N_9083);
nand U9622 (N_9622,N_9430,N_9067);
nand U9623 (N_9623,N_9142,N_9389);
xnor U9624 (N_9624,N_9338,N_9199);
nor U9625 (N_9625,N_9411,N_9418);
xor U9626 (N_9626,N_9161,N_9285);
nand U9627 (N_9627,N_9186,N_9410);
and U9628 (N_9628,N_9399,N_9440);
nand U9629 (N_9629,N_9467,N_9144);
nand U9630 (N_9630,N_9380,N_9174);
nor U9631 (N_9631,N_9286,N_9203);
nor U9632 (N_9632,N_9162,N_9354);
or U9633 (N_9633,N_9324,N_9362);
xnor U9634 (N_9634,N_9370,N_9390);
or U9635 (N_9635,N_9165,N_9375);
nor U9636 (N_9636,N_9364,N_9080);
and U9637 (N_9637,N_9282,N_9139);
nand U9638 (N_9638,N_9046,N_9437);
nor U9639 (N_9639,N_9172,N_9261);
nand U9640 (N_9640,N_9298,N_9252);
nand U9641 (N_9641,N_9329,N_9209);
nor U9642 (N_9642,N_9415,N_9442);
or U9643 (N_9643,N_9312,N_9350);
nor U9644 (N_9644,N_9271,N_9022);
or U9645 (N_9645,N_9010,N_9400);
or U9646 (N_9646,N_9248,N_9241);
and U9647 (N_9647,N_9250,N_9118);
xor U9648 (N_9648,N_9085,N_9426);
nor U9649 (N_9649,N_9392,N_9447);
and U9650 (N_9650,N_9200,N_9363);
nor U9651 (N_9651,N_9035,N_9208);
nor U9652 (N_9652,N_9472,N_9183);
nor U9653 (N_9653,N_9191,N_9145);
or U9654 (N_9654,N_9140,N_9021);
or U9655 (N_9655,N_9290,N_9361);
nand U9656 (N_9656,N_9226,N_9157);
nand U9657 (N_9657,N_9407,N_9180);
xor U9658 (N_9658,N_9138,N_9374);
and U9659 (N_9659,N_9478,N_9451);
nor U9660 (N_9660,N_9281,N_9296);
and U9661 (N_9661,N_9348,N_9387);
or U9662 (N_9662,N_9403,N_9232);
or U9663 (N_9663,N_9406,N_9227);
nor U9664 (N_9664,N_9061,N_9444);
nand U9665 (N_9665,N_9257,N_9167);
or U9666 (N_9666,N_9223,N_9225);
xnor U9667 (N_9667,N_9381,N_9355);
or U9668 (N_9668,N_9054,N_9284);
and U9669 (N_9669,N_9078,N_9222);
and U9670 (N_9670,N_9003,N_9051);
or U9671 (N_9671,N_9239,N_9423);
and U9672 (N_9672,N_9058,N_9347);
and U9673 (N_9673,N_9274,N_9053);
and U9674 (N_9674,N_9486,N_9386);
nor U9675 (N_9675,N_9214,N_9130);
nand U9676 (N_9676,N_9366,N_9453);
or U9677 (N_9677,N_9332,N_9098);
nor U9678 (N_9678,N_9480,N_9309);
and U9679 (N_9679,N_9446,N_9326);
nand U9680 (N_9680,N_9470,N_9477);
or U9681 (N_9681,N_9076,N_9217);
or U9682 (N_9682,N_9088,N_9207);
nand U9683 (N_9683,N_9075,N_9346);
xnor U9684 (N_9684,N_9082,N_9303);
nand U9685 (N_9685,N_9025,N_9132);
and U9686 (N_9686,N_9448,N_9244);
and U9687 (N_9687,N_9050,N_9059);
nor U9688 (N_9688,N_9441,N_9344);
xor U9689 (N_9689,N_9498,N_9108);
nand U9690 (N_9690,N_9249,N_9378);
or U9691 (N_9691,N_9212,N_9412);
and U9692 (N_9692,N_9484,N_9032);
and U9693 (N_9693,N_9268,N_9084);
or U9694 (N_9694,N_9293,N_9202);
and U9695 (N_9695,N_9388,N_9179);
and U9696 (N_9696,N_9473,N_9134);
and U9697 (N_9697,N_9218,N_9294);
nand U9698 (N_9698,N_9237,N_9081);
nor U9699 (N_9699,N_9356,N_9149);
nor U9700 (N_9700,N_9045,N_9417);
nand U9701 (N_9701,N_9376,N_9373);
nor U9702 (N_9702,N_9111,N_9020);
nand U9703 (N_9703,N_9367,N_9163);
and U9704 (N_9704,N_9345,N_9327);
and U9705 (N_9705,N_9295,N_9110);
xnor U9706 (N_9706,N_9481,N_9126);
nor U9707 (N_9707,N_9112,N_9064);
nand U9708 (N_9708,N_9087,N_9299);
xnor U9709 (N_9709,N_9432,N_9143);
or U9710 (N_9710,N_9351,N_9266);
xnor U9711 (N_9711,N_9404,N_9204);
or U9712 (N_9712,N_9192,N_9371);
nand U9713 (N_9713,N_9497,N_9224);
or U9714 (N_9714,N_9490,N_9231);
and U9715 (N_9715,N_9190,N_9166);
xnor U9716 (N_9716,N_9393,N_9487);
and U9717 (N_9717,N_9496,N_9030);
and U9718 (N_9718,N_9205,N_9048);
nor U9719 (N_9719,N_9184,N_9428);
and U9720 (N_9720,N_9195,N_9105);
or U9721 (N_9721,N_9047,N_9465);
and U9722 (N_9722,N_9368,N_9031);
and U9723 (N_9723,N_9377,N_9463);
or U9724 (N_9724,N_9116,N_9109);
nor U9725 (N_9725,N_9230,N_9468);
nand U9726 (N_9726,N_9263,N_9000);
nor U9727 (N_9727,N_9431,N_9421);
or U9728 (N_9728,N_9319,N_9023);
nor U9729 (N_9729,N_9128,N_9173);
nand U9730 (N_9730,N_9009,N_9276);
nor U9731 (N_9731,N_9100,N_9452);
and U9732 (N_9732,N_9255,N_9420);
nand U9733 (N_9733,N_9211,N_9383);
and U9734 (N_9734,N_9236,N_9011);
nand U9735 (N_9735,N_9328,N_9460);
nor U9736 (N_9736,N_9304,N_9262);
nor U9737 (N_9737,N_9001,N_9122);
xor U9738 (N_9738,N_9086,N_9482);
and U9739 (N_9739,N_9024,N_9315);
or U9740 (N_9740,N_9402,N_9495);
and U9741 (N_9741,N_9316,N_9057);
xnor U9742 (N_9742,N_9455,N_9331);
or U9743 (N_9743,N_9062,N_9198);
and U9744 (N_9744,N_9005,N_9193);
nor U9745 (N_9745,N_9065,N_9052);
and U9746 (N_9746,N_9301,N_9433);
nor U9747 (N_9747,N_9097,N_9206);
nor U9748 (N_9748,N_9492,N_9069);
xnor U9749 (N_9749,N_9018,N_9413);
nand U9750 (N_9750,N_9150,N_9090);
or U9751 (N_9751,N_9497,N_9038);
nand U9752 (N_9752,N_9135,N_9330);
and U9753 (N_9753,N_9200,N_9160);
or U9754 (N_9754,N_9070,N_9259);
and U9755 (N_9755,N_9467,N_9323);
nor U9756 (N_9756,N_9140,N_9450);
xor U9757 (N_9757,N_9463,N_9271);
nand U9758 (N_9758,N_9490,N_9159);
or U9759 (N_9759,N_9010,N_9394);
nand U9760 (N_9760,N_9492,N_9094);
or U9761 (N_9761,N_9217,N_9128);
and U9762 (N_9762,N_9417,N_9143);
or U9763 (N_9763,N_9005,N_9179);
nor U9764 (N_9764,N_9109,N_9053);
or U9765 (N_9765,N_9246,N_9451);
nand U9766 (N_9766,N_9304,N_9245);
and U9767 (N_9767,N_9355,N_9269);
and U9768 (N_9768,N_9354,N_9222);
or U9769 (N_9769,N_9054,N_9317);
nor U9770 (N_9770,N_9474,N_9110);
or U9771 (N_9771,N_9260,N_9411);
and U9772 (N_9772,N_9182,N_9123);
nor U9773 (N_9773,N_9236,N_9404);
or U9774 (N_9774,N_9002,N_9481);
nor U9775 (N_9775,N_9473,N_9162);
nor U9776 (N_9776,N_9136,N_9229);
nand U9777 (N_9777,N_9171,N_9259);
or U9778 (N_9778,N_9418,N_9226);
or U9779 (N_9779,N_9230,N_9320);
or U9780 (N_9780,N_9170,N_9295);
nand U9781 (N_9781,N_9245,N_9048);
nand U9782 (N_9782,N_9474,N_9434);
and U9783 (N_9783,N_9204,N_9022);
and U9784 (N_9784,N_9166,N_9173);
and U9785 (N_9785,N_9003,N_9463);
or U9786 (N_9786,N_9343,N_9204);
and U9787 (N_9787,N_9182,N_9375);
nand U9788 (N_9788,N_9199,N_9010);
nand U9789 (N_9789,N_9472,N_9467);
or U9790 (N_9790,N_9333,N_9326);
or U9791 (N_9791,N_9100,N_9028);
and U9792 (N_9792,N_9213,N_9021);
nor U9793 (N_9793,N_9492,N_9246);
xor U9794 (N_9794,N_9467,N_9006);
xor U9795 (N_9795,N_9379,N_9217);
nand U9796 (N_9796,N_9245,N_9224);
or U9797 (N_9797,N_9421,N_9035);
or U9798 (N_9798,N_9297,N_9191);
xnor U9799 (N_9799,N_9211,N_9331);
nand U9800 (N_9800,N_9287,N_9242);
xnor U9801 (N_9801,N_9106,N_9380);
nand U9802 (N_9802,N_9202,N_9051);
and U9803 (N_9803,N_9041,N_9062);
or U9804 (N_9804,N_9195,N_9097);
xor U9805 (N_9805,N_9019,N_9421);
nor U9806 (N_9806,N_9098,N_9061);
nor U9807 (N_9807,N_9355,N_9047);
or U9808 (N_9808,N_9177,N_9300);
nand U9809 (N_9809,N_9000,N_9006);
or U9810 (N_9810,N_9243,N_9474);
xnor U9811 (N_9811,N_9380,N_9055);
or U9812 (N_9812,N_9162,N_9349);
nor U9813 (N_9813,N_9023,N_9358);
and U9814 (N_9814,N_9024,N_9020);
nand U9815 (N_9815,N_9341,N_9029);
xor U9816 (N_9816,N_9197,N_9497);
and U9817 (N_9817,N_9403,N_9334);
and U9818 (N_9818,N_9276,N_9315);
nor U9819 (N_9819,N_9254,N_9264);
and U9820 (N_9820,N_9049,N_9058);
nand U9821 (N_9821,N_9260,N_9047);
nor U9822 (N_9822,N_9230,N_9186);
xnor U9823 (N_9823,N_9278,N_9403);
and U9824 (N_9824,N_9465,N_9052);
nor U9825 (N_9825,N_9327,N_9171);
or U9826 (N_9826,N_9308,N_9301);
nor U9827 (N_9827,N_9137,N_9264);
nor U9828 (N_9828,N_9161,N_9304);
nand U9829 (N_9829,N_9254,N_9052);
xor U9830 (N_9830,N_9053,N_9330);
nor U9831 (N_9831,N_9084,N_9336);
and U9832 (N_9832,N_9199,N_9297);
nand U9833 (N_9833,N_9495,N_9308);
nand U9834 (N_9834,N_9484,N_9457);
or U9835 (N_9835,N_9372,N_9145);
or U9836 (N_9836,N_9307,N_9425);
nand U9837 (N_9837,N_9334,N_9179);
or U9838 (N_9838,N_9132,N_9147);
and U9839 (N_9839,N_9223,N_9158);
and U9840 (N_9840,N_9379,N_9486);
nand U9841 (N_9841,N_9498,N_9166);
xnor U9842 (N_9842,N_9463,N_9316);
and U9843 (N_9843,N_9203,N_9309);
and U9844 (N_9844,N_9183,N_9335);
nor U9845 (N_9845,N_9453,N_9359);
nor U9846 (N_9846,N_9476,N_9316);
and U9847 (N_9847,N_9194,N_9331);
or U9848 (N_9848,N_9164,N_9189);
and U9849 (N_9849,N_9199,N_9155);
or U9850 (N_9850,N_9301,N_9421);
and U9851 (N_9851,N_9105,N_9113);
nor U9852 (N_9852,N_9239,N_9318);
and U9853 (N_9853,N_9335,N_9273);
xnor U9854 (N_9854,N_9089,N_9105);
xor U9855 (N_9855,N_9199,N_9092);
nor U9856 (N_9856,N_9457,N_9476);
or U9857 (N_9857,N_9399,N_9482);
or U9858 (N_9858,N_9444,N_9103);
nor U9859 (N_9859,N_9380,N_9379);
nor U9860 (N_9860,N_9337,N_9022);
or U9861 (N_9861,N_9454,N_9448);
nor U9862 (N_9862,N_9013,N_9282);
nor U9863 (N_9863,N_9280,N_9143);
or U9864 (N_9864,N_9035,N_9409);
xor U9865 (N_9865,N_9074,N_9308);
and U9866 (N_9866,N_9294,N_9049);
nor U9867 (N_9867,N_9312,N_9408);
nor U9868 (N_9868,N_9423,N_9370);
and U9869 (N_9869,N_9050,N_9222);
or U9870 (N_9870,N_9066,N_9419);
nor U9871 (N_9871,N_9394,N_9011);
xnor U9872 (N_9872,N_9003,N_9045);
or U9873 (N_9873,N_9447,N_9009);
or U9874 (N_9874,N_9316,N_9101);
or U9875 (N_9875,N_9254,N_9332);
and U9876 (N_9876,N_9253,N_9149);
nand U9877 (N_9877,N_9334,N_9402);
and U9878 (N_9878,N_9059,N_9256);
or U9879 (N_9879,N_9297,N_9160);
nor U9880 (N_9880,N_9057,N_9187);
or U9881 (N_9881,N_9023,N_9303);
nor U9882 (N_9882,N_9288,N_9182);
nor U9883 (N_9883,N_9282,N_9337);
nor U9884 (N_9884,N_9154,N_9141);
nor U9885 (N_9885,N_9122,N_9405);
nand U9886 (N_9886,N_9369,N_9211);
and U9887 (N_9887,N_9453,N_9144);
or U9888 (N_9888,N_9205,N_9113);
or U9889 (N_9889,N_9213,N_9080);
nor U9890 (N_9890,N_9083,N_9149);
nor U9891 (N_9891,N_9055,N_9252);
nand U9892 (N_9892,N_9174,N_9113);
nor U9893 (N_9893,N_9370,N_9297);
or U9894 (N_9894,N_9403,N_9250);
nand U9895 (N_9895,N_9249,N_9350);
nor U9896 (N_9896,N_9207,N_9435);
nor U9897 (N_9897,N_9287,N_9327);
or U9898 (N_9898,N_9369,N_9341);
or U9899 (N_9899,N_9000,N_9174);
and U9900 (N_9900,N_9304,N_9042);
xor U9901 (N_9901,N_9402,N_9068);
xnor U9902 (N_9902,N_9318,N_9237);
nor U9903 (N_9903,N_9340,N_9021);
nand U9904 (N_9904,N_9299,N_9361);
and U9905 (N_9905,N_9060,N_9480);
and U9906 (N_9906,N_9479,N_9133);
and U9907 (N_9907,N_9255,N_9457);
or U9908 (N_9908,N_9452,N_9008);
and U9909 (N_9909,N_9499,N_9228);
nand U9910 (N_9910,N_9435,N_9139);
and U9911 (N_9911,N_9055,N_9313);
nor U9912 (N_9912,N_9366,N_9143);
nand U9913 (N_9913,N_9285,N_9281);
or U9914 (N_9914,N_9453,N_9075);
or U9915 (N_9915,N_9244,N_9082);
nor U9916 (N_9916,N_9130,N_9068);
and U9917 (N_9917,N_9209,N_9373);
nor U9918 (N_9918,N_9169,N_9397);
nand U9919 (N_9919,N_9241,N_9406);
nand U9920 (N_9920,N_9460,N_9402);
and U9921 (N_9921,N_9139,N_9259);
nand U9922 (N_9922,N_9298,N_9098);
or U9923 (N_9923,N_9405,N_9419);
nor U9924 (N_9924,N_9440,N_9151);
or U9925 (N_9925,N_9277,N_9190);
nor U9926 (N_9926,N_9357,N_9212);
nor U9927 (N_9927,N_9165,N_9208);
and U9928 (N_9928,N_9184,N_9395);
xnor U9929 (N_9929,N_9392,N_9449);
or U9930 (N_9930,N_9225,N_9198);
or U9931 (N_9931,N_9068,N_9393);
or U9932 (N_9932,N_9417,N_9072);
nand U9933 (N_9933,N_9397,N_9223);
and U9934 (N_9934,N_9140,N_9005);
nand U9935 (N_9935,N_9060,N_9052);
or U9936 (N_9936,N_9452,N_9406);
and U9937 (N_9937,N_9163,N_9358);
or U9938 (N_9938,N_9043,N_9310);
nor U9939 (N_9939,N_9169,N_9371);
nor U9940 (N_9940,N_9293,N_9072);
xnor U9941 (N_9941,N_9398,N_9474);
and U9942 (N_9942,N_9032,N_9062);
and U9943 (N_9943,N_9210,N_9403);
nor U9944 (N_9944,N_9498,N_9424);
nor U9945 (N_9945,N_9051,N_9122);
or U9946 (N_9946,N_9161,N_9315);
nor U9947 (N_9947,N_9222,N_9250);
or U9948 (N_9948,N_9401,N_9272);
nor U9949 (N_9949,N_9174,N_9302);
nor U9950 (N_9950,N_9039,N_9198);
and U9951 (N_9951,N_9288,N_9465);
and U9952 (N_9952,N_9201,N_9252);
nand U9953 (N_9953,N_9474,N_9075);
nand U9954 (N_9954,N_9138,N_9111);
nand U9955 (N_9955,N_9204,N_9005);
and U9956 (N_9956,N_9331,N_9212);
or U9957 (N_9957,N_9473,N_9337);
or U9958 (N_9958,N_9497,N_9132);
and U9959 (N_9959,N_9398,N_9033);
nor U9960 (N_9960,N_9040,N_9387);
and U9961 (N_9961,N_9297,N_9320);
nand U9962 (N_9962,N_9306,N_9128);
nand U9963 (N_9963,N_9272,N_9131);
and U9964 (N_9964,N_9156,N_9405);
nor U9965 (N_9965,N_9313,N_9109);
xor U9966 (N_9966,N_9235,N_9284);
and U9967 (N_9967,N_9309,N_9045);
nand U9968 (N_9968,N_9326,N_9291);
or U9969 (N_9969,N_9252,N_9184);
nand U9970 (N_9970,N_9286,N_9109);
and U9971 (N_9971,N_9250,N_9449);
nand U9972 (N_9972,N_9156,N_9137);
nor U9973 (N_9973,N_9034,N_9431);
nor U9974 (N_9974,N_9247,N_9436);
nand U9975 (N_9975,N_9123,N_9096);
nand U9976 (N_9976,N_9000,N_9337);
xnor U9977 (N_9977,N_9240,N_9061);
or U9978 (N_9978,N_9197,N_9210);
and U9979 (N_9979,N_9055,N_9153);
nor U9980 (N_9980,N_9208,N_9196);
or U9981 (N_9981,N_9269,N_9163);
nor U9982 (N_9982,N_9278,N_9353);
xor U9983 (N_9983,N_9318,N_9460);
nand U9984 (N_9984,N_9032,N_9431);
nand U9985 (N_9985,N_9322,N_9394);
and U9986 (N_9986,N_9496,N_9319);
nor U9987 (N_9987,N_9364,N_9015);
nand U9988 (N_9988,N_9202,N_9346);
and U9989 (N_9989,N_9173,N_9175);
nand U9990 (N_9990,N_9492,N_9269);
nand U9991 (N_9991,N_9084,N_9124);
or U9992 (N_9992,N_9116,N_9441);
nor U9993 (N_9993,N_9408,N_9303);
nand U9994 (N_9994,N_9032,N_9300);
xnor U9995 (N_9995,N_9203,N_9117);
or U9996 (N_9996,N_9215,N_9076);
nand U9997 (N_9997,N_9305,N_9227);
nand U9998 (N_9998,N_9401,N_9293);
and U9999 (N_9999,N_9210,N_9066);
nor U10000 (N_10000,N_9886,N_9580);
or U10001 (N_10001,N_9946,N_9772);
and U10002 (N_10002,N_9988,N_9829);
nand U10003 (N_10003,N_9502,N_9859);
nor U10004 (N_10004,N_9658,N_9897);
nor U10005 (N_10005,N_9895,N_9800);
xor U10006 (N_10006,N_9602,N_9584);
or U10007 (N_10007,N_9742,N_9585);
nand U10008 (N_10008,N_9758,N_9938);
nor U10009 (N_10009,N_9522,N_9728);
and U10010 (N_10010,N_9595,N_9646);
nand U10011 (N_10011,N_9633,N_9773);
xor U10012 (N_10012,N_9509,N_9830);
or U10013 (N_10013,N_9521,N_9757);
nand U10014 (N_10014,N_9930,N_9870);
nor U10015 (N_10015,N_9849,N_9969);
or U10016 (N_10016,N_9611,N_9511);
or U10017 (N_10017,N_9604,N_9724);
or U10018 (N_10018,N_9581,N_9795);
and U10019 (N_10019,N_9572,N_9819);
or U10020 (N_10020,N_9915,N_9810);
nor U10021 (N_10021,N_9891,N_9540);
and U10022 (N_10022,N_9562,N_9873);
nand U10023 (N_10023,N_9642,N_9620);
nor U10024 (N_10024,N_9740,N_9710);
nand U10025 (N_10025,N_9600,N_9679);
nand U10026 (N_10026,N_9889,N_9631);
nor U10027 (N_10027,N_9902,N_9559);
or U10028 (N_10028,N_9677,N_9605);
or U10029 (N_10029,N_9627,N_9689);
and U10030 (N_10030,N_9615,N_9641);
and U10031 (N_10031,N_9623,N_9796);
or U10032 (N_10032,N_9993,N_9541);
and U10033 (N_10033,N_9507,N_9530);
and U10034 (N_10034,N_9578,N_9911);
nor U10035 (N_10035,N_9838,N_9753);
or U10036 (N_10036,N_9945,N_9931);
nor U10037 (N_10037,N_9943,N_9713);
nor U10038 (N_10038,N_9546,N_9591);
or U10039 (N_10039,N_9869,N_9699);
xor U10040 (N_10040,N_9697,N_9548);
and U10041 (N_10041,N_9506,N_9529);
nor U10042 (N_10042,N_9702,N_9929);
and U10043 (N_10043,N_9955,N_9735);
xor U10044 (N_10044,N_9860,N_9711);
and U10045 (N_10045,N_9709,N_9857);
or U10046 (N_10046,N_9893,N_9894);
and U10047 (N_10047,N_9538,N_9885);
and U10048 (N_10048,N_9972,N_9630);
nand U10049 (N_10049,N_9793,N_9835);
or U10050 (N_10050,N_9828,N_9625);
and U10051 (N_10051,N_9613,N_9832);
nor U10052 (N_10052,N_9537,N_9947);
or U10053 (N_10053,N_9996,N_9966);
and U10054 (N_10054,N_9571,N_9610);
or U10055 (N_10055,N_9552,N_9906);
nand U10056 (N_10056,N_9640,N_9590);
and U10057 (N_10057,N_9748,N_9942);
nor U10058 (N_10058,N_9504,N_9834);
nand U10059 (N_10059,N_9618,N_9898);
nor U10060 (N_10060,N_9525,N_9965);
nand U10061 (N_10061,N_9771,N_9567);
xor U10062 (N_10062,N_9779,N_9706);
or U10063 (N_10063,N_9659,N_9953);
or U10064 (N_10064,N_9576,N_9649);
and U10065 (N_10065,N_9652,N_9647);
nor U10066 (N_10066,N_9547,N_9896);
nand U10067 (N_10067,N_9596,N_9928);
or U10068 (N_10068,N_9816,N_9674);
nand U10069 (N_10069,N_9939,N_9801);
nand U10070 (N_10070,N_9990,N_9734);
or U10071 (N_10071,N_9935,N_9936);
or U10072 (N_10072,N_9961,N_9905);
nand U10073 (N_10073,N_9650,N_9629);
nor U10074 (N_10074,N_9846,N_9684);
xor U10075 (N_10075,N_9839,N_9926);
nand U10076 (N_10076,N_9764,N_9937);
nand U10077 (N_10077,N_9863,N_9637);
nor U10078 (N_10078,N_9919,N_9743);
xor U10079 (N_10079,N_9790,N_9954);
xnor U10080 (N_10080,N_9565,N_9617);
and U10081 (N_10081,N_9843,N_9705);
or U10082 (N_10082,N_9768,N_9730);
or U10083 (N_10083,N_9957,N_9660);
and U10084 (N_10084,N_9797,N_9880);
nor U10085 (N_10085,N_9696,N_9675);
and U10086 (N_10086,N_9909,N_9573);
nor U10087 (N_10087,N_9823,N_9974);
or U10088 (N_10088,N_9979,N_9651);
or U10089 (N_10089,N_9967,N_9803);
nor U10090 (N_10090,N_9688,N_9991);
and U10091 (N_10091,N_9874,N_9503);
nand U10092 (N_10092,N_9814,N_9704);
nand U10093 (N_10093,N_9827,N_9738);
and U10094 (N_10094,N_9731,N_9775);
nor U10095 (N_10095,N_9975,N_9887);
or U10096 (N_10096,N_9791,N_9553);
nand U10097 (N_10097,N_9986,N_9933);
nor U10098 (N_10098,N_9608,N_9519);
or U10099 (N_10099,N_9851,N_9820);
xnor U10100 (N_10100,N_9932,N_9720);
nand U10101 (N_10101,N_9760,N_9622);
or U10102 (N_10102,N_9989,N_9815);
xnor U10103 (N_10103,N_9976,N_9516);
or U10104 (N_10104,N_9528,N_9666);
xor U10105 (N_10105,N_9501,N_9575);
nand U10106 (N_10106,N_9635,N_9876);
and U10107 (N_10107,N_9999,N_9862);
xnor U10108 (N_10108,N_9598,N_9907);
and U10109 (N_10109,N_9599,N_9695);
and U10110 (N_10110,N_9958,N_9554);
and U10111 (N_10111,N_9856,N_9681);
or U10112 (N_10112,N_9632,N_9638);
or U10113 (N_10113,N_9985,N_9557);
and U10114 (N_10114,N_9708,N_9747);
nand U10115 (N_10115,N_9781,N_9766);
or U10116 (N_10116,N_9570,N_9566);
nand U10117 (N_10117,N_9736,N_9569);
xor U10118 (N_10118,N_9558,N_9992);
nor U10119 (N_10119,N_9845,N_9531);
xor U10120 (N_10120,N_9754,N_9904);
and U10121 (N_10121,N_9561,N_9987);
and U10122 (N_10122,N_9715,N_9539);
or U10123 (N_10123,N_9648,N_9872);
and U10124 (N_10124,N_9523,N_9916);
nor U10125 (N_10125,N_9712,N_9850);
nor U10126 (N_10126,N_9746,N_9913);
and U10127 (N_10127,N_9749,N_9837);
nand U10128 (N_10128,N_9807,N_9836);
nand U10129 (N_10129,N_9841,N_9668);
nor U10130 (N_10130,N_9950,N_9861);
nand U10131 (N_10131,N_9698,N_9729);
nand U10132 (N_10132,N_9995,N_9783);
nor U10133 (N_10133,N_9587,N_9984);
or U10134 (N_10134,N_9682,N_9717);
nand U10135 (N_10135,N_9513,N_9914);
or U10136 (N_10136,N_9520,N_9788);
xor U10137 (N_10137,N_9890,N_9798);
or U10138 (N_10138,N_9512,N_9669);
and U10139 (N_10139,N_9665,N_9645);
nor U10140 (N_10140,N_9722,N_9899);
or U10141 (N_10141,N_9741,N_9601);
nand U10142 (N_10142,N_9878,N_9733);
nor U10143 (N_10143,N_9639,N_9982);
or U10144 (N_10144,N_9517,N_9643);
nand U10145 (N_10145,N_9616,N_9844);
and U10146 (N_10146,N_9854,N_9903);
or U10147 (N_10147,N_9805,N_9952);
nand U10148 (N_10148,N_9607,N_9968);
xnor U10149 (N_10149,N_9774,N_9694);
and U10150 (N_10150,N_9609,N_9978);
or U10151 (N_10151,N_9744,N_9818);
or U10152 (N_10152,N_9664,N_9817);
nor U10153 (N_10153,N_9917,N_9714);
and U10154 (N_10154,N_9824,N_9685);
and U10155 (N_10155,N_9994,N_9518);
and U10156 (N_10156,N_9535,N_9770);
and U10157 (N_10157,N_9657,N_9515);
nand U10158 (N_10158,N_9971,N_9944);
nor U10159 (N_10159,N_9543,N_9867);
or U10160 (N_10160,N_9808,N_9809);
nor U10161 (N_10161,N_9691,N_9727);
and U10162 (N_10162,N_9802,N_9901);
xnor U10163 (N_10163,N_9787,N_9782);
nand U10164 (N_10164,N_9550,N_9716);
nand U10165 (N_10165,N_9508,N_9551);
and U10166 (N_10166,N_9732,N_9923);
and U10167 (N_10167,N_9606,N_9761);
nor U10168 (N_10168,N_9750,N_9564);
nand U10169 (N_10169,N_9769,N_9621);
nand U10170 (N_10170,N_9737,N_9582);
or U10171 (N_10171,N_9960,N_9866);
nor U10172 (N_10172,N_9505,N_9555);
nand U10173 (N_10173,N_9794,N_9912);
nand U10174 (N_10174,N_9811,N_9686);
and U10175 (N_10175,N_9763,N_9921);
nor U10176 (N_10176,N_9678,N_9888);
nand U10177 (N_10177,N_9981,N_9532);
or U10178 (N_10178,N_9804,N_9977);
or U10179 (N_10179,N_9799,N_9925);
and U10180 (N_10180,N_9594,N_9723);
and U10181 (N_10181,N_9780,N_9778);
and U10182 (N_10182,N_9739,N_9603);
nand U10183 (N_10183,N_9822,N_9980);
and U10184 (N_10184,N_9784,N_9619);
nor U10185 (N_10185,N_9671,N_9514);
nor U10186 (N_10186,N_9959,N_9868);
or U10187 (N_10187,N_9721,N_9776);
or U10188 (N_10188,N_9568,N_9700);
xnor U10189 (N_10189,N_9612,N_9589);
nand U10190 (N_10190,N_9527,N_9725);
nand U10191 (N_10191,N_9833,N_9579);
and U10192 (N_10192,N_9628,N_9910);
nor U10193 (N_10193,N_9583,N_9879);
nor U10194 (N_10194,N_9973,N_9847);
nor U10195 (N_10195,N_9821,N_9526);
nor U10196 (N_10196,N_9786,N_9500);
or U10197 (N_10197,N_9556,N_9892);
or U10198 (N_10198,N_9624,N_9871);
nand U10199 (N_10199,N_9962,N_9577);
nor U10200 (N_10200,N_9670,N_9812);
and U10201 (N_10201,N_9544,N_9908);
and U10202 (N_10202,N_9542,N_9667);
or U10203 (N_10203,N_9881,N_9875);
nand U10204 (N_10204,N_9970,N_9941);
nor U10205 (N_10205,N_9922,N_9653);
nor U10206 (N_10206,N_9842,N_9692);
or U10207 (N_10207,N_9534,N_9656);
or U10208 (N_10208,N_9662,N_9884);
nand U10209 (N_10209,N_9683,N_9680);
nor U10210 (N_10210,N_9672,N_9777);
and U10211 (N_10211,N_9964,N_9673);
nor U10212 (N_10212,N_9983,N_9853);
nor U10213 (N_10213,N_9510,N_9877);
or U10214 (N_10214,N_9592,N_9864);
and U10215 (N_10215,N_9755,N_9762);
and U10216 (N_10216,N_9718,N_9951);
nand U10217 (N_10217,N_9998,N_9536);
nand U10218 (N_10218,N_9586,N_9997);
nor U10219 (N_10219,N_9963,N_9813);
nand U10220 (N_10220,N_9690,N_9719);
nor U10221 (N_10221,N_9940,N_9759);
xor U10222 (N_10222,N_9707,N_9767);
nor U10223 (N_10223,N_9636,N_9745);
or U10224 (N_10224,N_9882,N_9756);
or U10225 (N_10225,N_9524,N_9806);
xor U10226 (N_10226,N_9831,N_9593);
and U10227 (N_10227,N_9792,N_9789);
xnor U10228 (N_10228,N_9865,N_9701);
or U10229 (N_10229,N_9655,N_9597);
xnor U10230 (N_10230,N_9563,N_9924);
xnor U10231 (N_10231,N_9765,N_9858);
nor U10232 (N_10232,N_9533,N_9825);
nand U10233 (N_10233,N_9934,N_9883);
or U10234 (N_10234,N_9693,N_9920);
nand U10235 (N_10235,N_9752,N_9687);
nor U10236 (N_10236,N_9588,N_9634);
and U10237 (N_10237,N_9676,N_9848);
or U10238 (N_10238,N_9663,N_9626);
or U10239 (N_10239,N_9785,N_9918);
and U10240 (N_10240,N_9956,N_9840);
nand U10241 (N_10241,N_9751,N_9927);
xor U10242 (N_10242,N_9855,N_9654);
and U10243 (N_10243,N_9644,N_9726);
nor U10244 (N_10244,N_9900,N_9852);
nand U10245 (N_10245,N_9560,N_9614);
nor U10246 (N_10246,N_9661,N_9826);
and U10247 (N_10247,N_9703,N_9949);
and U10248 (N_10248,N_9948,N_9549);
nand U10249 (N_10249,N_9545,N_9574);
nand U10250 (N_10250,N_9950,N_9955);
nand U10251 (N_10251,N_9647,N_9705);
nand U10252 (N_10252,N_9889,N_9819);
or U10253 (N_10253,N_9823,N_9610);
nand U10254 (N_10254,N_9981,N_9852);
and U10255 (N_10255,N_9534,N_9709);
xnor U10256 (N_10256,N_9745,N_9975);
nand U10257 (N_10257,N_9563,N_9917);
nand U10258 (N_10258,N_9715,N_9615);
xnor U10259 (N_10259,N_9602,N_9790);
or U10260 (N_10260,N_9674,N_9534);
or U10261 (N_10261,N_9705,N_9948);
or U10262 (N_10262,N_9985,N_9512);
nand U10263 (N_10263,N_9987,N_9860);
nor U10264 (N_10264,N_9630,N_9813);
or U10265 (N_10265,N_9840,N_9812);
or U10266 (N_10266,N_9932,N_9569);
and U10267 (N_10267,N_9856,N_9742);
nor U10268 (N_10268,N_9521,N_9609);
and U10269 (N_10269,N_9948,N_9514);
or U10270 (N_10270,N_9594,N_9572);
and U10271 (N_10271,N_9925,N_9623);
nor U10272 (N_10272,N_9800,N_9612);
and U10273 (N_10273,N_9929,N_9666);
or U10274 (N_10274,N_9529,N_9595);
nand U10275 (N_10275,N_9627,N_9581);
or U10276 (N_10276,N_9712,N_9997);
or U10277 (N_10277,N_9807,N_9665);
nand U10278 (N_10278,N_9710,N_9761);
or U10279 (N_10279,N_9518,N_9924);
and U10280 (N_10280,N_9676,N_9885);
nor U10281 (N_10281,N_9854,N_9852);
and U10282 (N_10282,N_9633,N_9886);
nor U10283 (N_10283,N_9924,N_9918);
and U10284 (N_10284,N_9890,N_9557);
or U10285 (N_10285,N_9799,N_9948);
nor U10286 (N_10286,N_9791,N_9776);
nor U10287 (N_10287,N_9938,N_9925);
nand U10288 (N_10288,N_9978,N_9894);
or U10289 (N_10289,N_9693,N_9684);
nand U10290 (N_10290,N_9923,N_9883);
nor U10291 (N_10291,N_9812,N_9579);
nand U10292 (N_10292,N_9767,N_9909);
or U10293 (N_10293,N_9680,N_9939);
and U10294 (N_10294,N_9774,N_9628);
xnor U10295 (N_10295,N_9689,N_9853);
xor U10296 (N_10296,N_9873,N_9566);
or U10297 (N_10297,N_9746,N_9853);
or U10298 (N_10298,N_9502,N_9808);
xnor U10299 (N_10299,N_9951,N_9856);
and U10300 (N_10300,N_9718,N_9783);
nand U10301 (N_10301,N_9784,N_9545);
and U10302 (N_10302,N_9973,N_9952);
xnor U10303 (N_10303,N_9798,N_9771);
and U10304 (N_10304,N_9687,N_9715);
and U10305 (N_10305,N_9900,N_9961);
and U10306 (N_10306,N_9966,N_9561);
nand U10307 (N_10307,N_9666,N_9668);
nor U10308 (N_10308,N_9619,N_9796);
xnor U10309 (N_10309,N_9935,N_9932);
and U10310 (N_10310,N_9604,N_9988);
and U10311 (N_10311,N_9897,N_9594);
nor U10312 (N_10312,N_9889,N_9838);
nand U10313 (N_10313,N_9624,N_9817);
nand U10314 (N_10314,N_9820,N_9514);
xor U10315 (N_10315,N_9578,N_9973);
or U10316 (N_10316,N_9790,N_9752);
or U10317 (N_10317,N_9695,N_9678);
or U10318 (N_10318,N_9675,N_9838);
and U10319 (N_10319,N_9611,N_9618);
or U10320 (N_10320,N_9893,N_9981);
or U10321 (N_10321,N_9963,N_9918);
nand U10322 (N_10322,N_9797,N_9742);
or U10323 (N_10323,N_9796,N_9711);
xnor U10324 (N_10324,N_9728,N_9518);
or U10325 (N_10325,N_9816,N_9762);
xnor U10326 (N_10326,N_9989,N_9677);
nand U10327 (N_10327,N_9930,N_9916);
nor U10328 (N_10328,N_9749,N_9983);
nor U10329 (N_10329,N_9974,N_9761);
nor U10330 (N_10330,N_9869,N_9956);
nand U10331 (N_10331,N_9833,N_9821);
and U10332 (N_10332,N_9913,N_9786);
xor U10333 (N_10333,N_9569,N_9734);
xor U10334 (N_10334,N_9508,N_9992);
and U10335 (N_10335,N_9841,N_9795);
or U10336 (N_10336,N_9509,N_9925);
or U10337 (N_10337,N_9889,N_9743);
or U10338 (N_10338,N_9857,N_9774);
xor U10339 (N_10339,N_9579,N_9815);
nand U10340 (N_10340,N_9598,N_9758);
nand U10341 (N_10341,N_9959,N_9727);
or U10342 (N_10342,N_9533,N_9680);
xor U10343 (N_10343,N_9921,N_9755);
or U10344 (N_10344,N_9632,N_9521);
nand U10345 (N_10345,N_9881,N_9904);
nor U10346 (N_10346,N_9774,N_9543);
or U10347 (N_10347,N_9557,N_9655);
nor U10348 (N_10348,N_9752,N_9748);
xnor U10349 (N_10349,N_9608,N_9947);
nor U10350 (N_10350,N_9641,N_9731);
nand U10351 (N_10351,N_9625,N_9584);
nand U10352 (N_10352,N_9613,N_9547);
and U10353 (N_10353,N_9955,N_9647);
and U10354 (N_10354,N_9727,N_9510);
xnor U10355 (N_10355,N_9571,N_9971);
xor U10356 (N_10356,N_9601,N_9973);
xnor U10357 (N_10357,N_9865,N_9666);
nor U10358 (N_10358,N_9628,N_9996);
and U10359 (N_10359,N_9554,N_9681);
and U10360 (N_10360,N_9564,N_9943);
or U10361 (N_10361,N_9889,N_9590);
nor U10362 (N_10362,N_9777,N_9536);
or U10363 (N_10363,N_9832,N_9567);
and U10364 (N_10364,N_9806,N_9943);
nor U10365 (N_10365,N_9984,N_9798);
nand U10366 (N_10366,N_9888,N_9999);
nor U10367 (N_10367,N_9898,N_9712);
and U10368 (N_10368,N_9676,N_9549);
and U10369 (N_10369,N_9761,N_9507);
or U10370 (N_10370,N_9840,N_9790);
nor U10371 (N_10371,N_9881,N_9787);
and U10372 (N_10372,N_9941,N_9813);
and U10373 (N_10373,N_9936,N_9507);
or U10374 (N_10374,N_9925,N_9965);
nor U10375 (N_10375,N_9715,N_9946);
nor U10376 (N_10376,N_9624,N_9683);
or U10377 (N_10377,N_9869,N_9540);
and U10378 (N_10378,N_9814,N_9818);
nor U10379 (N_10379,N_9817,N_9708);
and U10380 (N_10380,N_9686,N_9930);
nor U10381 (N_10381,N_9600,N_9695);
nand U10382 (N_10382,N_9588,N_9603);
nor U10383 (N_10383,N_9795,N_9978);
nand U10384 (N_10384,N_9731,N_9570);
and U10385 (N_10385,N_9855,N_9854);
nor U10386 (N_10386,N_9796,N_9550);
nor U10387 (N_10387,N_9874,N_9552);
nand U10388 (N_10388,N_9938,N_9631);
xor U10389 (N_10389,N_9829,N_9898);
and U10390 (N_10390,N_9927,N_9741);
and U10391 (N_10391,N_9785,N_9505);
nand U10392 (N_10392,N_9862,N_9601);
nand U10393 (N_10393,N_9998,N_9868);
nor U10394 (N_10394,N_9736,N_9688);
nand U10395 (N_10395,N_9510,N_9863);
nor U10396 (N_10396,N_9638,N_9877);
xnor U10397 (N_10397,N_9572,N_9881);
xnor U10398 (N_10398,N_9965,N_9549);
nand U10399 (N_10399,N_9815,N_9839);
or U10400 (N_10400,N_9704,N_9787);
and U10401 (N_10401,N_9658,N_9751);
nor U10402 (N_10402,N_9886,N_9936);
nand U10403 (N_10403,N_9999,N_9932);
nor U10404 (N_10404,N_9607,N_9953);
or U10405 (N_10405,N_9915,N_9749);
xnor U10406 (N_10406,N_9941,N_9653);
nand U10407 (N_10407,N_9650,N_9862);
nor U10408 (N_10408,N_9975,N_9692);
nand U10409 (N_10409,N_9787,N_9835);
xnor U10410 (N_10410,N_9876,N_9787);
and U10411 (N_10411,N_9967,N_9674);
xor U10412 (N_10412,N_9637,N_9618);
nand U10413 (N_10413,N_9987,N_9806);
nor U10414 (N_10414,N_9552,N_9531);
nand U10415 (N_10415,N_9885,N_9509);
nand U10416 (N_10416,N_9605,N_9737);
and U10417 (N_10417,N_9625,N_9633);
or U10418 (N_10418,N_9816,N_9879);
or U10419 (N_10419,N_9939,N_9917);
or U10420 (N_10420,N_9632,N_9621);
and U10421 (N_10421,N_9786,N_9748);
and U10422 (N_10422,N_9900,N_9614);
nor U10423 (N_10423,N_9698,N_9980);
nor U10424 (N_10424,N_9557,N_9726);
nand U10425 (N_10425,N_9841,N_9503);
nand U10426 (N_10426,N_9521,N_9748);
and U10427 (N_10427,N_9828,N_9906);
xor U10428 (N_10428,N_9599,N_9931);
and U10429 (N_10429,N_9649,N_9993);
and U10430 (N_10430,N_9549,N_9865);
nand U10431 (N_10431,N_9942,N_9913);
xnor U10432 (N_10432,N_9710,N_9811);
nand U10433 (N_10433,N_9745,N_9635);
and U10434 (N_10434,N_9513,N_9957);
nor U10435 (N_10435,N_9732,N_9775);
xnor U10436 (N_10436,N_9764,N_9967);
or U10437 (N_10437,N_9798,N_9925);
nand U10438 (N_10438,N_9894,N_9542);
nor U10439 (N_10439,N_9553,N_9797);
nor U10440 (N_10440,N_9501,N_9826);
xnor U10441 (N_10441,N_9509,N_9869);
or U10442 (N_10442,N_9565,N_9576);
xnor U10443 (N_10443,N_9625,N_9887);
nor U10444 (N_10444,N_9670,N_9578);
and U10445 (N_10445,N_9528,N_9905);
or U10446 (N_10446,N_9712,N_9683);
and U10447 (N_10447,N_9860,N_9986);
nand U10448 (N_10448,N_9676,N_9918);
or U10449 (N_10449,N_9667,N_9892);
or U10450 (N_10450,N_9992,N_9778);
and U10451 (N_10451,N_9512,N_9951);
and U10452 (N_10452,N_9875,N_9751);
nor U10453 (N_10453,N_9643,N_9990);
or U10454 (N_10454,N_9538,N_9884);
and U10455 (N_10455,N_9643,N_9825);
or U10456 (N_10456,N_9614,N_9845);
nor U10457 (N_10457,N_9530,N_9767);
nor U10458 (N_10458,N_9951,N_9982);
nor U10459 (N_10459,N_9807,N_9875);
nand U10460 (N_10460,N_9756,N_9969);
or U10461 (N_10461,N_9701,N_9613);
xnor U10462 (N_10462,N_9911,N_9634);
nand U10463 (N_10463,N_9830,N_9585);
and U10464 (N_10464,N_9675,N_9729);
nand U10465 (N_10465,N_9927,N_9808);
nor U10466 (N_10466,N_9682,N_9595);
nand U10467 (N_10467,N_9557,N_9810);
or U10468 (N_10468,N_9958,N_9980);
xor U10469 (N_10469,N_9624,N_9948);
nor U10470 (N_10470,N_9587,N_9749);
nand U10471 (N_10471,N_9740,N_9806);
or U10472 (N_10472,N_9540,N_9827);
or U10473 (N_10473,N_9782,N_9853);
and U10474 (N_10474,N_9678,N_9810);
nand U10475 (N_10475,N_9630,N_9902);
and U10476 (N_10476,N_9519,N_9727);
or U10477 (N_10477,N_9777,N_9564);
nand U10478 (N_10478,N_9878,N_9952);
or U10479 (N_10479,N_9578,N_9972);
nand U10480 (N_10480,N_9598,N_9562);
or U10481 (N_10481,N_9683,N_9564);
or U10482 (N_10482,N_9644,N_9904);
nor U10483 (N_10483,N_9660,N_9624);
or U10484 (N_10484,N_9957,N_9663);
nor U10485 (N_10485,N_9812,N_9601);
or U10486 (N_10486,N_9743,N_9759);
or U10487 (N_10487,N_9555,N_9508);
nand U10488 (N_10488,N_9666,N_9980);
and U10489 (N_10489,N_9779,N_9920);
nand U10490 (N_10490,N_9611,N_9950);
or U10491 (N_10491,N_9713,N_9614);
nand U10492 (N_10492,N_9944,N_9562);
nor U10493 (N_10493,N_9728,N_9701);
nor U10494 (N_10494,N_9781,N_9765);
and U10495 (N_10495,N_9856,N_9997);
nand U10496 (N_10496,N_9879,N_9779);
or U10497 (N_10497,N_9639,N_9577);
and U10498 (N_10498,N_9655,N_9661);
or U10499 (N_10499,N_9518,N_9522);
nor U10500 (N_10500,N_10324,N_10002);
and U10501 (N_10501,N_10420,N_10379);
or U10502 (N_10502,N_10454,N_10244);
nor U10503 (N_10503,N_10074,N_10446);
nand U10504 (N_10504,N_10090,N_10099);
and U10505 (N_10505,N_10155,N_10092);
nand U10506 (N_10506,N_10243,N_10374);
nor U10507 (N_10507,N_10165,N_10472);
xnor U10508 (N_10508,N_10350,N_10283);
nor U10509 (N_10509,N_10333,N_10176);
or U10510 (N_10510,N_10315,N_10382);
nand U10511 (N_10511,N_10105,N_10117);
or U10512 (N_10512,N_10085,N_10214);
and U10513 (N_10513,N_10273,N_10299);
nand U10514 (N_10514,N_10358,N_10162);
nor U10515 (N_10515,N_10488,N_10292);
or U10516 (N_10516,N_10052,N_10349);
and U10517 (N_10517,N_10175,N_10259);
and U10518 (N_10518,N_10432,N_10112);
and U10519 (N_10519,N_10400,N_10263);
and U10520 (N_10520,N_10410,N_10058);
nor U10521 (N_10521,N_10107,N_10422);
or U10522 (N_10522,N_10027,N_10051);
and U10523 (N_10523,N_10285,N_10178);
and U10524 (N_10524,N_10386,N_10113);
and U10525 (N_10525,N_10414,N_10039);
and U10526 (N_10526,N_10206,N_10030);
nor U10527 (N_10527,N_10218,N_10055);
nand U10528 (N_10528,N_10252,N_10097);
nor U10529 (N_10529,N_10319,N_10373);
or U10530 (N_10530,N_10148,N_10241);
nand U10531 (N_10531,N_10017,N_10317);
nand U10532 (N_10532,N_10024,N_10257);
or U10533 (N_10533,N_10050,N_10225);
or U10534 (N_10534,N_10466,N_10485);
nor U10535 (N_10535,N_10023,N_10106);
or U10536 (N_10536,N_10494,N_10134);
nand U10537 (N_10537,N_10473,N_10355);
nor U10538 (N_10538,N_10098,N_10197);
nand U10539 (N_10539,N_10413,N_10450);
and U10540 (N_10540,N_10075,N_10332);
or U10541 (N_10541,N_10191,N_10347);
or U10542 (N_10542,N_10281,N_10397);
or U10543 (N_10543,N_10093,N_10004);
and U10544 (N_10544,N_10160,N_10471);
nor U10545 (N_10545,N_10448,N_10409);
and U10546 (N_10546,N_10198,N_10069);
nor U10547 (N_10547,N_10268,N_10267);
nand U10548 (N_10548,N_10128,N_10076);
nand U10549 (N_10549,N_10284,N_10111);
xor U10550 (N_10550,N_10266,N_10094);
or U10551 (N_10551,N_10272,N_10036);
nand U10552 (N_10552,N_10102,N_10083);
xnor U10553 (N_10553,N_10343,N_10444);
nand U10554 (N_10554,N_10223,N_10354);
nand U10555 (N_10555,N_10262,N_10322);
nor U10556 (N_10556,N_10337,N_10145);
or U10557 (N_10557,N_10288,N_10101);
nand U10558 (N_10558,N_10242,N_10313);
or U10559 (N_10559,N_10362,N_10059);
or U10560 (N_10560,N_10141,N_10452);
nor U10561 (N_10561,N_10161,N_10378);
nor U10562 (N_10562,N_10224,N_10303);
nand U10563 (N_10563,N_10238,N_10384);
nand U10564 (N_10564,N_10202,N_10486);
or U10565 (N_10565,N_10264,N_10327);
nand U10566 (N_10566,N_10103,N_10309);
and U10567 (N_10567,N_10046,N_10121);
and U10568 (N_10568,N_10330,N_10217);
nor U10569 (N_10569,N_10174,N_10199);
or U10570 (N_10570,N_10290,N_10497);
and U10571 (N_10571,N_10430,N_10153);
or U10572 (N_10572,N_10367,N_10345);
or U10573 (N_10573,N_10431,N_10269);
or U10574 (N_10574,N_10133,N_10037);
nor U10575 (N_10575,N_10169,N_10275);
or U10576 (N_10576,N_10368,N_10192);
nor U10577 (N_10577,N_10163,N_10477);
xnor U10578 (N_10578,N_10171,N_10467);
or U10579 (N_10579,N_10261,N_10212);
or U10580 (N_10580,N_10061,N_10032);
xor U10581 (N_10581,N_10247,N_10395);
xnor U10582 (N_10582,N_10108,N_10479);
nand U10583 (N_10583,N_10219,N_10132);
and U10584 (N_10584,N_10047,N_10120);
nor U10585 (N_10585,N_10063,N_10307);
or U10586 (N_10586,N_10230,N_10271);
and U10587 (N_10587,N_10189,N_10158);
or U10588 (N_10588,N_10054,N_10442);
and U10589 (N_10589,N_10460,N_10240);
xor U10590 (N_10590,N_10087,N_10496);
nor U10591 (N_10591,N_10416,N_10402);
nor U10592 (N_10592,N_10360,N_10072);
and U10593 (N_10593,N_10136,N_10482);
and U10594 (N_10594,N_10455,N_10065);
nand U10595 (N_10595,N_10179,N_10251);
nor U10596 (N_10596,N_10260,N_10321);
xnor U10597 (N_10597,N_10369,N_10270);
nand U10598 (N_10598,N_10351,N_10078);
nor U10599 (N_10599,N_10335,N_10041);
xnor U10600 (N_10600,N_10383,N_10417);
and U10601 (N_10601,N_10449,N_10089);
and U10602 (N_10602,N_10375,N_10484);
or U10603 (N_10603,N_10492,N_10205);
and U10604 (N_10604,N_10186,N_10201);
nor U10605 (N_10605,N_10211,N_10234);
or U10606 (N_10606,N_10091,N_10012);
nor U10607 (N_10607,N_10018,N_10125);
nand U10608 (N_10608,N_10489,N_10237);
and U10609 (N_10609,N_10480,N_10325);
or U10610 (N_10610,N_10487,N_10067);
or U10611 (N_10611,N_10038,N_10437);
nand U10612 (N_10612,N_10329,N_10361);
and U10613 (N_10613,N_10000,N_10468);
nor U10614 (N_10614,N_10068,N_10356);
or U10615 (N_10615,N_10282,N_10221);
and U10616 (N_10616,N_10289,N_10233);
and U10617 (N_10617,N_10157,N_10256);
and U10618 (N_10618,N_10081,N_10139);
or U10619 (N_10619,N_10143,N_10474);
nand U10620 (N_10620,N_10405,N_10295);
or U10621 (N_10621,N_10095,N_10159);
nand U10622 (N_10622,N_10415,N_10291);
and U10623 (N_10623,N_10210,N_10129);
and U10624 (N_10624,N_10394,N_10499);
or U10625 (N_10625,N_10286,N_10183);
nor U10626 (N_10626,N_10249,N_10483);
nand U10627 (N_10627,N_10014,N_10232);
xor U10628 (N_10628,N_10147,N_10478);
and U10629 (N_10629,N_10399,N_10056);
nor U10630 (N_10630,N_10131,N_10433);
and U10631 (N_10631,N_10213,N_10130);
nand U10632 (N_10632,N_10021,N_10293);
and U10633 (N_10633,N_10001,N_10035);
nor U10634 (N_10634,N_10436,N_10306);
nor U10635 (N_10635,N_10184,N_10071);
or U10636 (N_10636,N_10173,N_10421);
and U10637 (N_10637,N_10438,N_10254);
or U10638 (N_10638,N_10138,N_10328);
nor U10639 (N_10639,N_10008,N_10019);
or U10640 (N_10640,N_10190,N_10418);
nor U10641 (N_10641,N_10043,N_10458);
nor U10642 (N_10642,N_10048,N_10045);
nand U10643 (N_10643,N_10152,N_10428);
or U10644 (N_10644,N_10470,N_10044);
nor U10645 (N_10645,N_10073,N_10135);
xor U10646 (N_10646,N_10278,N_10118);
nor U10647 (N_10647,N_10222,N_10311);
nor U10648 (N_10648,N_10334,N_10396);
nor U10649 (N_10649,N_10215,N_10151);
nand U10650 (N_10650,N_10250,N_10235);
and U10651 (N_10651,N_10427,N_10156);
nor U10652 (N_10652,N_10253,N_10393);
xnor U10653 (N_10653,N_10304,N_10364);
xnor U10654 (N_10654,N_10308,N_10344);
or U10655 (N_10655,N_10009,N_10390);
or U10656 (N_10656,N_10167,N_10227);
nor U10657 (N_10657,N_10086,N_10359);
or U10658 (N_10658,N_10022,N_10464);
nor U10659 (N_10659,N_10231,N_10408);
nor U10660 (N_10660,N_10426,N_10406);
or U10661 (N_10661,N_10195,N_10180);
nor U10662 (N_10662,N_10164,N_10419);
and U10663 (N_10663,N_10265,N_10182);
and U10664 (N_10664,N_10387,N_10104);
and U10665 (N_10665,N_10380,N_10392);
nor U10666 (N_10666,N_10126,N_10323);
nor U10667 (N_10667,N_10435,N_10204);
and U10668 (N_10668,N_10287,N_10318);
nand U10669 (N_10669,N_10226,N_10297);
nand U10670 (N_10670,N_10277,N_10025);
and U10671 (N_10671,N_10348,N_10026);
nor U10672 (N_10672,N_10404,N_10080);
nor U10673 (N_10673,N_10124,N_10029);
nor U10674 (N_10674,N_10381,N_10491);
or U10675 (N_10675,N_10209,N_10181);
nor U10676 (N_10676,N_10064,N_10296);
and U10677 (N_10677,N_10049,N_10423);
or U10678 (N_10678,N_10279,N_10403);
or U10679 (N_10679,N_10439,N_10385);
nor U10680 (N_10680,N_10339,N_10248);
nand U10681 (N_10681,N_10185,N_10445);
or U10682 (N_10682,N_10398,N_10168);
nor U10683 (N_10683,N_10336,N_10109);
and U10684 (N_10684,N_10340,N_10114);
or U10685 (N_10685,N_10301,N_10352);
nand U10686 (N_10686,N_10236,N_10376);
nor U10687 (N_10687,N_10388,N_10294);
nand U10688 (N_10688,N_10082,N_10481);
or U10689 (N_10689,N_10434,N_10006);
nor U10690 (N_10690,N_10020,N_10429);
nand U10691 (N_10691,N_10110,N_10365);
or U10692 (N_10692,N_10028,N_10255);
and U10693 (N_10693,N_10057,N_10003);
xor U10694 (N_10694,N_10493,N_10172);
or U10695 (N_10695,N_10137,N_10007);
nand U10696 (N_10696,N_10320,N_10062);
or U10697 (N_10697,N_10475,N_10314);
nor U10698 (N_10698,N_10146,N_10088);
nand U10699 (N_10699,N_10258,N_10342);
and U10700 (N_10700,N_10316,N_10194);
nor U10701 (N_10701,N_10353,N_10401);
and U10702 (N_10702,N_10013,N_10084);
nor U10703 (N_10703,N_10412,N_10011);
and U10704 (N_10704,N_10476,N_10100);
nor U10705 (N_10705,N_10298,N_10469);
nor U10706 (N_10706,N_10363,N_10389);
and U10707 (N_10707,N_10070,N_10440);
and U10708 (N_10708,N_10119,N_10451);
nand U10709 (N_10709,N_10031,N_10077);
and U10710 (N_10710,N_10033,N_10490);
nor U10711 (N_10711,N_10424,N_10443);
xnor U10712 (N_10712,N_10463,N_10425);
nor U10713 (N_10713,N_10203,N_10096);
nand U10714 (N_10714,N_10127,N_10465);
or U10715 (N_10715,N_10193,N_10150);
and U10716 (N_10716,N_10015,N_10276);
and U10717 (N_10717,N_10495,N_10338);
nor U10718 (N_10718,N_10341,N_10461);
nor U10719 (N_10719,N_10229,N_10372);
and U10720 (N_10720,N_10170,N_10122);
nor U10721 (N_10721,N_10177,N_10142);
or U10722 (N_10722,N_10200,N_10371);
or U10723 (N_10723,N_10300,N_10196);
or U10724 (N_10724,N_10040,N_10447);
nor U10725 (N_10725,N_10310,N_10079);
nand U10726 (N_10726,N_10326,N_10274);
and U10727 (N_10727,N_10187,N_10331);
nor U10728 (N_10728,N_10010,N_10280);
nor U10729 (N_10729,N_10391,N_10016);
nor U10730 (N_10730,N_10042,N_10166);
xor U10731 (N_10731,N_10498,N_10245);
xor U10732 (N_10732,N_10228,N_10005);
nor U10733 (N_10733,N_10053,N_10188);
xor U10734 (N_10734,N_10144,N_10060);
and U10735 (N_10735,N_10370,N_10034);
nand U10736 (N_10736,N_10116,N_10302);
and U10737 (N_10737,N_10366,N_10207);
nand U10738 (N_10738,N_10346,N_10154);
nor U10739 (N_10739,N_10407,N_10459);
and U10740 (N_10740,N_10123,N_10140);
and U10741 (N_10741,N_10441,N_10377);
xnor U10742 (N_10742,N_10456,N_10216);
nand U10743 (N_10743,N_10066,N_10357);
or U10744 (N_10744,N_10453,N_10305);
nor U10745 (N_10745,N_10115,N_10208);
or U10746 (N_10746,N_10457,N_10239);
xor U10747 (N_10747,N_10246,N_10220);
and U10748 (N_10748,N_10149,N_10411);
and U10749 (N_10749,N_10312,N_10462);
nor U10750 (N_10750,N_10113,N_10437);
or U10751 (N_10751,N_10053,N_10076);
nor U10752 (N_10752,N_10461,N_10119);
nand U10753 (N_10753,N_10431,N_10126);
nand U10754 (N_10754,N_10302,N_10476);
and U10755 (N_10755,N_10323,N_10184);
nor U10756 (N_10756,N_10324,N_10150);
nand U10757 (N_10757,N_10470,N_10246);
xnor U10758 (N_10758,N_10390,N_10164);
xnor U10759 (N_10759,N_10171,N_10239);
and U10760 (N_10760,N_10337,N_10289);
and U10761 (N_10761,N_10196,N_10331);
nor U10762 (N_10762,N_10391,N_10416);
nand U10763 (N_10763,N_10124,N_10445);
nand U10764 (N_10764,N_10446,N_10253);
and U10765 (N_10765,N_10217,N_10045);
and U10766 (N_10766,N_10275,N_10359);
nand U10767 (N_10767,N_10205,N_10122);
and U10768 (N_10768,N_10406,N_10330);
nor U10769 (N_10769,N_10182,N_10329);
nand U10770 (N_10770,N_10245,N_10106);
and U10771 (N_10771,N_10239,N_10130);
nand U10772 (N_10772,N_10387,N_10484);
xnor U10773 (N_10773,N_10280,N_10116);
and U10774 (N_10774,N_10405,N_10057);
and U10775 (N_10775,N_10316,N_10422);
nor U10776 (N_10776,N_10311,N_10036);
and U10777 (N_10777,N_10202,N_10478);
or U10778 (N_10778,N_10288,N_10062);
or U10779 (N_10779,N_10118,N_10175);
nor U10780 (N_10780,N_10304,N_10104);
nor U10781 (N_10781,N_10201,N_10111);
or U10782 (N_10782,N_10276,N_10136);
or U10783 (N_10783,N_10014,N_10375);
nand U10784 (N_10784,N_10041,N_10076);
xnor U10785 (N_10785,N_10284,N_10377);
nand U10786 (N_10786,N_10203,N_10336);
or U10787 (N_10787,N_10285,N_10116);
xnor U10788 (N_10788,N_10287,N_10042);
and U10789 (N_10789,N_10251,N_10396);
and U10790 (N_10790,N_10086,N_10197);
nand U10791 (N_10791,N_10215,N_10430);
nand U10792 (N_10792,N_10320,N_10049);
nor U10793 (N_10793,N_10445,N_10072);
nor U10794 (N_10794,N_10374,N_10029);
nand U10795 (N_10795,N_10232,N_10292);
and U10796 (N_10796,N_10373,N_10044);
and U10797 (N_10797,N_10350,N_10036);
or U10798 (N_10798,N_10163,N_10438);
nand U10799 (N_10799,N_10244,N_10355);
nand U10800 (N_10800,N_10156,N_10175);
and U10801 (N_10801,N_10346,N_10119);
or U10802 (N_10802,N_10332,N_10499);
xor U10803 (N_10803,N_10415,N_10064);
or U10804 (N_10804,N_10113,N_10470);
nand U10805 (N_10805,N_10070,N_10313);
or U10806 (N_10806,N_10368,N_10050);
nand U10807 (N_10807,N_10098,N_10474);
and U10808 (N_10808,N_10383,N_10468);
xnor U10809 (N_10809,N_10135,N_10268);
and U10810 (N_10810,N_10341,N_10348);
nand U10811 (N_10811,N_10183,N_10418);
and U10812 (N_10812,N_10372,N_10046);
or U10813 (N_10813,N_10092,N_10274);
and U10814 (N_10814,N_10303,N_10256);
nor U10815 (N_10815,N_10007,N_10270);
and U10816 (N_10816,N_10475,N_10462);
or U10817 (N_10817,N_10342,N_10176);
and U10818 (N_10818,N_10308,N_10371);
nand U10819 (N_10819,N_10411,N_10311);
nand U10820 (N_10820,N_10437,N_10412);
nor U10821 (N_10821,N_10167,N_10208);
nand U10822 (N_10822,N_10355,N_10241);
or U10823 (N_10823,N_10461,N_10331);
or U10824 (N_10824,N_10015,N_10411);
nor U10825 (N_10825,N_10402,N_10125);
and U10826 (N_10826,N_10326,N_10485);
or U10827 (N_10827,N_10067,N_10073);
xnor U10828 (N_10828,N_10350,N_10451);
nand U10829 (N_10829,N_10152,N_10236);
or U10830 (N_10830,N_10380,N_10122);
or U10831 (N_10831,N_10177,N_10438);
nand U10832 (N_10832,N_10312,N_10291);
nor U10833 (N_10833,N_10281,N_10081);
or U10834 (N_10834,N_10455,N_10343);
or U10835 (N_10835,N_10446,N_10069);
nand U10836 (N_10836,N_10148,N_10397);
nor U10837 (N_10837,N_10446,N_10245);
and U10838 (N_10838,N_10207,N_10284);
nand U10839 (N_10839,N_10074,N_10014);
nand U10840 (N_10840,N_10410,N_10485);
nor U10841 (N_10841,N_10270,N_10423);
nor U10842 (N_10842,N_10156,N_10399);
and U10843 (N_10843,N_10197,N_10234);
nor U10844 (N_10844,N_10041,N_10345);
or U10845 (N_10845,N_10232,N_10318);
nand U10846 (N_10846,N_10030,N_10212);
nand U10847 (N_10847,N_10235,N_10239);
xor U10848 (N_10848,N_10141,N_10056);
nand U10849 (N_10849,N_10167,N_10321);
xnor U10850 (N_10850,N_10338,N_10126);
and U10851 (N_10851,N_10216,N_10231);
nand U10852 (N_10852,N_10207,N_10198);
or U10853 (N_10853,N_10448,N_10015);
nand U10854 (N_10854,N_10481,N_10149);
and U10855 (N_10855,N_10063,N_10302);
or U10856 (N_10856,N_10337,N_10484);
or U10857 (N_10857,N_10185,N_10231);
nand U10858 (N_10858,N_10280,N_10480);
and U10859 (N_10859,N_10218,N_10033);
or U10860 (N_10860,N_10121,N_10428);
and U10861 (N_10861,N_10173,N_10430);
or U10862 (N_10862,N_10337,N_10020);
and U10863 (N_10863,N_10303,N_10331);
nor U10864 (N_10864,N_10041,N_10268);
nor U10865 (N_10865,N_10051,N_10213);
nand U10866 (N_10866,N_10401,N_10115);
and U10867 (N_10867,N_10162,N_10377);
and U10868 (N_10868,N_10175,N_10440);
or U10869 (N_10869,N_10002,N_10257);
or U10870 (N_10870,N_10097,N_10385);
nand U10871 (N_10871,N_10363,N_10042);
nor U10872 (N_10872,N_10426,N_10388);
nand U10873 (N_10873,N_10122,N_10328);
and U10874 (N_10874,N_10239,N_10113);
nor U10875 (N_10875,N_10333,N_10271);
or U10876 (N_10876,N_10248,N_10289);
or U10877 (N_10877,N_10382,N_10288);
and U10878 (N_10878,N_10005,N_10452);
nor U10879 (N_10879,N_10377,N_10126);
and U10880 (N_10880,N_10233,N_10178);
nand U10881 (N_10881,N_10068,N_10231);
or U10882 (N_10882,N_10423,N_10028);
nor U10883 (N_10883,N_10041,N_10460);
or U10884 (N_10884,N_10499,N_10346);
xnor U10885 (N_10885,N_10338,N_10207);
nand U10886 (N_10886,N_10290,N_10476);
xnor U10887 (N_10887,N_10194,N_10335);
nand U10888 (N_10888,N_10213,N_10091);
or U10889 (N_10889,N_10081,N_10058);
and U10890 (N_10890,N_10454,N_10153);
nor U10891 (N_10891,N_10394,N_10313);
and U10892 (N_10892,N_10016,N_10248);
nor U10893 (N_10893,N_10365,N_10280);
nor U10894 (N_10894,N_10277,N_10243);
or U10895 (N_10895,N_10388,N_10366);
nor U10896 (N_10896,N_10393,N_10065);
nor U10897 (N_10897,N_10387,N_10175);
or U10898 (N_10898,N_10369,N_10468);
and U10899 (N_10899,N_10193,N_10194);
or U10900 (N_10900,N_10123,N_10206);
xor U10901 (N_10901,N_10244,N_10067);
or U10902 (N_10902,N_10068,N_10090);
and U10903 (N_10903,N_10174,N_10077);
and U10904 (N_10904,N_10391,N_10372);
nand U10905 (N_10905,N_10120,N_10377);
nand U10906 (N_10906,N_10434,N_10138);
xor U10907 (N_10907,N_10128,N_10302);
or U10908 (N_10908,N_10391,N_10088);
or U10909 (N_10909,N_10143,N_10492);
nand U10910 (N_10910,N_10304,N_10255);
nand U10911 (N_10911,N_10180,N_10444);
or U10912 (N_10912,N_10279,N_10184);
nand U10913 (N_10913,N_10467,N_10108);
or U10914 (N_10914,N_10058,N_10256);
nor U10915 (N_10915,N_10102,N_10470);
or U10916 (N_10916,N_10395,N_10198);
and U10917 (N_10917,N_10216,N_10237);
or U10918 (N_10918,N_10104,N_10097);
nor U10919 (N_10919,N_10198,N_10414);
nor U10920 (N_10920,N_10424,N_10176);
xor U10921 (N_10921,N_10193,N_10411);
nand U10922 (N_10922,N_10299,N_10353);
and U10923 (N_10923,N_10162,N_10177);
and U10924 (N_10924,N_10439,N_10061);
nand U10925 (N_10925,N_10175,N_10041);
or U10926 (N_10926,N_10130,N_10070);
nor U10927 (N_10927,N_10414,N_10078);
nand U10928 (N_10928,N_10004,N_10258);
and U10929 (N_10929,N_10444,N_10327);
nand U10930 (N_10930,N_10488,N_10138);
and U10931 (N_10931,N_10245,N_10195);
nand U10932 (N_10932,N_10482,N_10133);
or U10933 (N_10933,N_10468,N_10018);
and U10934 (N_10934,N_10136,N_10405);
or U10935 (N_10935,N_10303,N_10382);
xor U10936 (N_10936,N_10143,N_10457);
or U10937 (N_10937,N_10341,N_10304);
and U10938 (N_10938,N_10049,N_10301);
and U10939 (N_10939,N_10316,N_10320);
xnor U10940 (N_10940,N_10447,N_10274);
nand U10941 (N_10941,N_10048,N_10122);
nand U10942 (N_10942,N_10480,N_10202);
and U10943 (N_10943,N_10270,N_10000);
or U10944 (N_10944,N_10355,N_10174);
or U10945 (N_10945,N_10267,N_10475);
or U10946 (N_10946,N_10166,N_10210);
xnor U10947 (N_10947,N_10067,N_10403);
nand U10948 (N_10948,N_10052,N_10129);
and U10949 (N_10949,N_10080,N_10044);
nor U10950 (N_10950,N_10136,N_10361);
and U10951 (N_10951,N_10317,N_10242);
nor U10952 (N_10952,N_10450,N_10184);
nor U10953 (N_10953,N_10456,N_10442);
and U10954 (N_10954,N_10268,N_10152);
and U10955 (N_10955,N_10279,N_10271);
nor U10956 (N_10956,N_10124,N_10409);
and U10957 (N_10957,N_10345,N_10400);
nand U10958 (N_10958,N_10250,N_10154);
nor U10959 (N_10959,N_10464,N_10145);
and U10960 (N_10960,N_10260,N_10252);
and U10961 (N_10961,N_10410,N_10470);
or U10962 (N_10962,N_10444,N_10260);
or U10963 (N_10963,N_10289,N_10161);
nor U10964 (N_10964,N_10048,N_10251);
nand U10965 (N_10965,N_10486,N_10204);
nor U10966 (N_10966,N_10199,N_10127);
nand U10967 (N_10967,N_10200,N_10245);
nor U10968 (N_10968,N_10385,N_10181);
or U10969 (N_10969,N_10117,N_10135);
nand U10970 (N_10970,N_10393,N_10045);
nor U10971 (N_10971,N_10016,N_10326);
nand U10972 (N_10972,N_10255,N_10270);
and U10973 (N_10973,N_10059,N_10485);
nand U10974 (N_10974,N_10319,N_10106);
or U10975 (N_10975,N_10040,N_10226);
xnor U10976 (N_10976,N_10335,N_10251);
nor U10977 (N_10977,N_10454,N_10380);
nor U10978 (N_10978,N_10046,N_10363);
nor U10979 (N_10979,N_10403,N_10014);
or U10980 (N_10980,N_10013,N_10324);
or U10981 (N_10981,N_10232,N_10055);
and U10982 (N_10982,N_10037,N_10262);
or U10983 (N_10983,N_10078,N_10254);
xor U10984 (N_10984,N_10012,N_10433);
and U10985 (N_10985,N_10017,N_10008);
or U10986 (N_10986,N_10017,N_10180);
or U10987 (N_10987,N_10088,N_10476);
and U10988 (N_10988,N_10178,N_10128);
and U10989 (N_10989,N_10097,N_10167);
and U10990 (N_10990,N_10293,N_10277);
or U10991 (N_10991,N_10381,N_10331);
and U10992 (N_10992,N_10144,N_10426);
or U10993 (N_10993,N_10370,N_10301);
and U10994 (N_10994,N_10405,N_10009);
nand U10995 (N_10995,N_10239,N_10132);
xnor U10996 (N_10996,N_10181,N_10381);
nor U10997 (N_10997,N_10138,N_10399);
and U10998 (N_10998,N_10444,N_10069);
and U10999 (N_10999,N_10447,N_10413);
or U11000 (N_11000,N_10870,N_10647);
nor U11001 (N_11001,N_10800,N_10676);
nor U11002 (N_11002,N_10677,N_10701);
nand U11003 (N_11003,N_10743,N_10876);
nor U11004 (N_11004,N_10950,N_10920);
or U11005 (N_11005,N_10696,N_10652);
and U11006 (N_11006,N_10726,N_10672);
and U11007 (N_11007,N_10810,N_10815);
nor U11008 (N_11008,N_10654,N_10767);
or U11009 (N_11009,N_10752,N_10751);
xor U11010 (N_11010,N_10621,N_10711);
and U11011 (N_11011,N_10649,N_10906);
xor U11012 (N_11012,N_10880,N_10771);
and U11013 (N_11013,N_10709,N_10554);
and U11014 (N_11014,N_10718,N_10904);
nor U11015 (N_11015,N_10629,N_10681);
or U11016 (N_11016,N_10566,N_10712);
and U11017 (N_11017,N_10570,N_10531);
or U11018 (N_11018,N_10909,N_10734);
nor U11019 (N_11019,N_10863,N_10731);
or U11020 (N_11020,N_10929,N_10937);
or U11021 (N_11021,N_10979,N_10874);
nor U11022 (N_11022,N_10534,N_10866);
nand U11023 (N_11023,N_10749,N_10998);
nand U11024 (N_11024,N_10759,N_10877);
and U11025 (N_11025,N_10797,N_10873);
and U11026 (N_11026,N_10723,N_10926);
xnor U11027 (N_11027,N_10669,N_10653);
and U11028 (N_11028,N_10804,N_10793);
or U11029 (N_11029,N_10732,N_10747);
and U11030 (N_11030,N_10692,N_10829);
or U11031 (N_11031,N_10957,N_10646);
xor U11032 (N_11032,N_10932,N_10742);
nor U11033 (N_11033,N_10986,N_10820);
nand U11034 (N_11034,N_10883,N_10779);
and U11035 (N_11035,N_10715,N_10660);
and U11036 (N_11036,N_10817,N_10849);
and U11037 (N_11037,N_10781,N_10942);
and U11038 (N_11038,N_10974,N_10834);
or U11039 (N_11039,N_10748,N_10841);
nand U11040 (N_11040,N_10847,N_10875);
nand U11041 (N_11041,N_10643,N_10985);
nand U11042 (N_11042,N_10776,N_10967);
or U11043 (N_11043,N_10869,N_10641);
and U11044 (N_11044,N_10541,N_10801);
nor U11045 (N_11045,N_10609,N_10894);
and U11046 (N_11046,N_10947,N_10903);
nor U11047 (N_11047,N_10954,N_10548);
or U11048 (N_11048,N_10960,N_10618);
xnor U11049 (N_11049,N_10768,N_10547);
and U11050 (N_11050,N_10577,N_10725);
and U11051 (N_11051,N_10746,N_10886);
nand U11052 (N_11052,N_10902,N_10970);
or U11053 (N_11053,N_10520,N_10917);
or U11054 (N_11054,N_10704,N_10995);
or U11055 (N_11055,N_10630,N_10956);
nand U11056 (N_11056,N_10848,N_10750);
xnor U11057 (N_11057,N_10540,N_10586);
nor U11058 (N_11058,N_10924,N_10938);
or U11059 (N_11059,N_10828,N_10941);
nand U11060 (N_11060,N_10864,N_10802);
and U11061 (N_11061,N_10662,N_10513);
and U11062 (N_11062,N_10509,N_10984);
nor U11063 (N_11063,N_10900,N_10683);
nand U11064 (N_11064,N_10708,N_10588);
nor U11065 (N_11065,N_10818,N_10925);
or U11066 (N_11066,N_10843,N_10627);
nand U11067 (N_11067,N_10603,N_10714);
or U11068 (N_11068,N_10699,N_10765);
nor U11069 (N_11069,N_10552,N_10565);
and U11070 (N_11070,N_10961,N_10695);
or U11071 (N_11071,N_10664,N_10506);
nor U11072 (N_11072,N_10582,N_10852);
or U11073 (N_11073,N_10578,N_10790);
and U11074 (N_11074,N_10616,N_10931);
and U11075 (N_11075,N_10968,N_10935);
or U11076 (N_11076,N_10533,N_10576);
nor U11077 (N_11077,N_10831,N_10892);
and U11078 (N_11078,N_10542,N_10997);
and U11079 (N_11079,N_10567,N_10733);
and U11080 (N_11080,N_10936,N_10774);
and U11081 (N_11081,N_10777,N_10607);
nor U11082 (N_11082,N_10637,N_10922);
nor U11083 (N_11083,N_10821,N_10528);
nor U11084 (N_11084,N_10835,N_10933);
nor U11085 (N_11085,N_10888,N_10644);
nand U11086 (N_11086,N_10833,N_10772);
or U11087 (N_11087,N_10661,N_10796);
nand U11088 (N_11088,N_10503,N_10686);
and U11089 (N_11089,N_10898,N_10798);
nand U11090 (N_11090,N_10501,N_10678);
nor U11091 (N_11091,N_10505,N_10812);
and U11092 (N_11092,N_10690,N_10510);
nor U11093 (N_11093,N_10809,N_10901);
nor U11094 (N_11094,N_10530,N_10614);
nand U11095 (N_11095,N_10634,N_10571);
and U11096 (N_11096,N_10885,N_10553);
or U11097 (N_11097,N_10545,N_10787);
xnor U11098 (N_11098,N_10564,N_10899);
nand U11099 (N_11099,N_10978,N_10795);
xnor U11100 (N_11100,N_10601,N_10893);
or U11101 (N_11101,N_10949,N_10700);
nor U11102 (N_11102,N_10626,N_10546);
or U11103 (N_11103,N_10910,N_10816);
or U11104 (N_11104,N_10611,N_10871);
nor U11105 (N_11105,N_10688,N_10955);
nand U11106 (N_11106,N_10918,N_10856);
nor U11107 (N_11107,N_10980,N_10773);
or U11108 (N_11108,N_10791,N_10803);
xor U11109 (N_11109,N_10633,N_10838);
nand U11110 (N_11110,N_10703,N_10551);
or U11111 (N_11111,N_10782,N_10911);
or U11112 (N_11112,N_10517,N_10658);
and U11113 (N_11113,N_10934,N_10550);
or U11114 (N_11114,N_10792,N_10525);
nand U11115 (N_11115,N_10940,N_10555);
nor U11116 (N_11116,N_10764,N_10784);
nor U11117 (N_11117,N_10783,N_10560);
nor U11118 (N_11118,N_10824,N_10504);
nand U11119 (N_11119,N_10663,N_10754);
and U11120 (N_11120,N_10508,N_10832);
or U11121 (N_11121,N_10753,N_10819);
and U11122 (N_11122,N_10854,N_10622);
nor U11123 (N_11123,N_10826,N_10987);
and U11124 (N_11124,N_10994,N_10722);
and U11125 (N_11125,N_10830,N_10656);
and U11126 (N_11126,N_10945,N_10982);
nand U11127 (N_11127,N_10615,N_10671);
nor U11128 (N_11128,N_10972,N_10719);
and U11129 (N_11129,N_10745,N_10666);
nor U11130 (N_11130,N_10685,N_10907);
nor U11131 (N_11131,N_10939,N_10881);
nor U11132 (N_11132,N_10613,N_10868);
and U11133 (N_11133,N_10514,N_10872);
and U11134 (N_11134,N_10697,N_10727);
and U11135 (N_11135,N_10593,N_10993);
nand U11136 (N_11136,N_10916,N_10617);
or U11137 (N_11137,N_10572,N_10558);
nand U11138 (N_11138,N_10515,N_10568);
xor U11139 (N_11139,N_10579,N_10999);
or U11140 (N_11140,N_10963,N_10966);
and U11141 (N_11141,N_10657,N_10535);
nand U11142 (N_11142,N_10702,N_10825);
or U11143 (N_11143,N_10592,N_10665);
and U11144 (N_11144,N_10740,N_10590);
xor U11145 (N_11145,N_10597,N_10775);
and U11146 (N_11146,N_10608,N_10981);
and U11147 (N_11147,N_10707,N_10507);
nor U11148 (N_11148,N_10905,N_10527);
nand U11149 (N_11149,N_10584,N_10575);
nor U11150 (N_11150,N_10602,N_10988);
and U11151 (N_11151,N_10983,N_10595);
nor U11152 (N_11152,N_10735,N_10739);
or U11153 (N_11153,N_10827,N_10573);
or U11154 (N_11154,N_10670,N_10549);
and U11155 (N_11155,N_10591,N_10585);
nor U11156 (N_11156,N_10599,N_10612);
nand U11157 (N_11157,N_10996,N_10887);
nor U11158 (N_11158,N_10822,N_10624);
nor U11159 (N_11159,N_10799,N_10951);
or U11160 (N_11160,N_10655,N_10619);
xnor U11161 (N_11161,N_10919,N_10620);
xor U11162 (N_11162,N_10844,N_10557);
and U11163 (N_11163,N_10559,N_10720);
nand U11164 (N_11164,N_10853,N_10770);
nand U11165 (N_11165,N_10814,N_10605);
nor U11166 (N_11166,N_10758,N_10836);
or U11167 (N_11167,N_10760,N_10561);
nand U11168 (N_11168,N_10895,N_10502);
and U11169 (N_11169,N_10878,N_10581);
nand U11170 (N_11170,N_10842,N_10908);
and U11171 (N_11171,N_10710,N_10857);
nor U11172 (N_11172,N_10921,N_10524);
nor U11173 (N_11173,N_10891,N_10840);
nor U11174 (N_11174,N_10521,N_10964);
or U11175 (N_11175,N_10628,N_10927);
nand U11176 (N_11176,N_10716,N_10511);
nor U11177 (N_11177,N_10958,N_10667);
or U11178 (N_11178,N_10729,N_10890);
or U11179 (N_11179,N_10562,N_10741);
and U11180 (N_11180,N_10589,N_10689);
nor U11181 (N_11181,N_10537,N_10944);
or U11182 (N_11182,N_10896,N_10736);
and U11183 (N_11183,N_10632,N_10539);
or U11184 (N_11184,N_10596,N_10594);
and U11185 (N_11185,N_10807,N_10580);
or U11186 (N_11186,N_10650,N_10912);
or U11187 (N_11187,N_10569,N_10625);
nand U11188 (N_11188,N_10529,N_10992);
xnor U11189 (N_11189,N_10737,N_10691);
nor U11190 (N_11190,N_10543,N_10687);
or U11191 (N_11191,N_10762,N_10674);
nand U11192 (N_11192,N_10648,N_10780);
nand U11193 (N_11193,N_10721,N_10889);
nor U11194 (N_11194,N_10500,N_10860);
nor U11195 (N_11195,N_10913,N_10808);
or U11196 (N_11196,N_10684,N_10522);
and U11197 (N_11197,N_10724,N_10761);
nor U11198 (N_11198,N_10959,N_10642);
and U11199 (N_11199,N_10636,N_10668);
or U11200 (N_11200,N_10813,N_10717);
xor U11201 (N_11201,N_10786,N_10673);
or U11202 (N_11202,N_10823,N_10861);
nor U11203 (N_11203,N_10990,N_10977);
nand U11204 (N_11204,N_10583,N_10518);
xnor U11205 (N_11205,N_10587,N_10846);
nor U11206 (N_11206,N_10850,N_10606);
nor U11207 (N_11207,N_10526,N_10556);
and U11208 (N_11208,N_10788,N_10698);
and U11209 (N_11209,N_10659,N_10989);
and U11210 (N_11210,N_10755,N_10858);
or U11211 (N_11211,N_10682,N_10756);
or U11212 (N_11212,N_10769,N_10794);
and U11213 (N_11213,N_10785,N_10757);
nor U11214 (N_11214,N_10975,N_10705);
or U11215 (N_11215,N_10738,N_10943);
and U11216 (N_11216,N_10915,N_10763);
nand U11217 (N_11217,N_10635,N_10845);
xnor U11218 (N_11218,N_10532,N_10600);
and U11219 (N_11219,N_10694,N_10598);
xor U11220 (N_11220,N_10523,N_10859);
nor U11221 (N_11221,N_10728,N_10930);
nand U11222 (N_11222,N_10512,N_10976);
nand U11223 (N_11223,N_10563,N_10914);
xnor U11224 (N_11224,N_10952,N_10867);
or U11225 (N_11225,N_10882,N_10744);
and U11226 (N_11226,N_10645,N_10638);
nor U11227 (N_11227,N_10706,N_10610);
and U11228 (N_11228,N_10778,N_10538);
nor U11229 (N_11229,N_10675,N_10806);
nand U11230 (N_11230,N_10651,N_10544);
nor U11231 (N_11231,N_10946,N_10884);
or U11232 (N_11232,N_10639,N_10971);
nor U11233 (N_11233,N_10865,N_10805);
nand U11234 (N_11234,N_10897,N_10923);
nand U11235 (N_11235,N_10536,N_10855);
and U11236 (N_11236,N_10693,N_10574);
nor U11237 (N_11237,N_10516,N_10811);
nor U11238 (N_11238,N_10965,N_10680);
or U11239 (N_11239,N_10730,N_10519);
or U11240 (N_11240,N_10928,N_10948);
nor U11241 (N_11241,N_10837,N_10839);
nand U11242 (N_11242,N_10862,N_10851);
and U11243 (N_11243,N_10953,N_10789);
nand U11244 (N_11244,N_10679,N_10973);
xnor U11245 (N_11245,N_10623,N_10713);
nor U11246 (N_11246,N_10969,N_10604);
or U11247 (N_11247,N_10962,N_10631);
or U11248 (N_11248,N_10640,N_10766);
xnor U11249 (N_11249,N_10991,N_10879);
nand U11250 (N_11250,N_10760,N_10916);
nand U11251 (N_11251,N_10954,N_10626);
nand U11252 (N_11252,N_10614,N_10836);
and U11253 (N_11253,N_10917,N_10871);
and U11254 (N_11254,N_10541,N_10710);
and U11255 (N_11255,N_10994,N_10538);
or U11256 (N_11256,N_10550,N_10923);
xor U11257 (N_11257,N_10504,N_10699);
xor U11258 (N_11258,N_10709,N_10782);
xor U11259 (N_11259,N_10510,N_10742);
and U11260 (N_11260,N_10520,N_10616);
and U11261 (N_11261,N_10758,N_10980);
or U11262 (N_11262,N_10870,N_10628);
nor U11263 (N_11263,N_10522,N_10902);
nor U11264 (N_11264,N_10516,N_10727);
and U11265 (N_11265,N_10717,N_10850);
and U11266 (N_11266,N_10818,N_10836);
nor U11267 (N_11267,N_10780,N_10968);
or U11268 (N_11268,N_10760,N_10893);
or U11269 (N_11269,N_10754,N_10559);
or U11270 (N_11270,N_10700,N_10666);
and U11271 (N_11271,N_10840,N_10956);
or U11272 (N_11272,N_10987,N_10951);
nand U11273 (N_11273,N_10876,N_10973);
and U11274 (N_11274,N_10649,N_10544);
and U11275 (N_11275,N_10502,N_10624);
or U11276 (N_11276,N_10964,N_10809);
and U11277 (N_11277,N_10609,N_10711);
nor U11278 (N_11278,N_10840,N_10524);
or U11279 (N_11279,N_10515,N_10556);
or U11280 (N_11280,N_10946,N_10830);
or U11281 (N_11281,N_10567,N_10506);
and U11282 (N_11282,N_10980,N_10986);
and U11283 (N_11283,N_10895,N_10569);
or U11284 (N_11284,N_10785,N_10661);
nor U11285 (N_11285,N_10548,N_10927);
nor U11286 (N_11286,N_10727,N_10974);
nor U11287 (N_11287,N_10781,N_10824);
and U11288 (N_11288,N_10624,N_10672);
and U11289 (N_11289,N_10909,N_10952);
or U11290 (N_11290,N_10831,N_10705);
and U11291 (N_11291,N_10848,N_10776);
or U11292 (N_11292,N_10504,N_10542);
nor U11293 (N_11293,N_10785,N_10885);
or U11294 (N_11294,N_10557,N_10784);
and U11295 (N_11295,N_10772,N_10648);
or U11296 (N_11296,N_10991,N_10579);
nand U11297 (N_11297,N_10874,N_10787);
and U11298 (N_11298,N_10591,N_10668);
and U11299 (N_11299,N_10949,N_10555);
nor U11300 (N_11300,N_10996,N_10610);
and U11301 (N_11301,N_10854,N_10537);
and U11302 (N_11302,N_10554,N_10979);
and U11303 (N_11303,N_10593,N_10535);
nor U11304 (N_11304,N_10936,N_10941);
nor U11305 (N_11305,N_10752,N_10700);
or U11306 (N_11306,N_10701,N_10832);
and U11307 (N_11307,N_10845,N_10509);
nand U11308 (N_11308,N_10789,N_10924);
and U11309 (N_11309,N_10945,N_10618);
and U11310 (N_11310,N_10730,N_10507);
xnor U11311 (N_11311,N_10798,N_10656);
nand U11312 (N_11312,N_10751,N_10932);
nor U11313 (N_11313,N_10664,N_10585);
nor U11314 (N_11314,N_10695,N_10729);
nor U11315 (N_11315,N_10557,N_10798);
or U11316 (N_11316,N_10715,N_10964);
and U11317 (N_11317,N_10518,N_10655);
xor U11318 (N_11318,N_10533,N_10555);
or U11319 (N_11319,N_10909,N_10610);
and U11320 (N_11320,N_10765,N_10925);
nand U11321 (N_11321,N_10771,N_10828);
nor U11322 (N_11322,N_10649,N_10773);
nand U11323 (N_11323,N_10801,N_10704);
nand U11324 (N_11324,N_10667,N_10664);
nor U11325 (N_11325,N_10867,N_10822);
or U11326 (N_11326,N_10777,N_10851);
nand U11327 (N_11327,N_10818,N_10966);
nand U11328 (N_11328,N_10770,N_10687);
nand U11329 (N_11329,N_10686,N_10608);
and U11330 (N_11330,N_10702,N_10669);
xor U11331 (N_11331,N_10589,N_10503);
nor U11332 (N_11332,N_10651,N_10826);
nor U11333 (N_11333,N_10649,N_10577);
nand U11334 (N_11334,N_10739,N_10960);
and U11335 (N_11335,N_10641,N_10862);
nand U11336 (N_11336,N_10990,N_10569);
nand U11337 (N_11337,N_10874,N_10883);
nor U11338 (N_11338,N_10710,N_10571);
xnor U11339 (N_11339,N_10920,N_10982);
or U11340 (N_11340,N_10944,N_10919);
nand U11341 (N_11341,N_10883,N_10621);
nor U11342 (N_11342,N_10828,N_10721);
or U11343 (N_11343,N_10675,N_10937);
and U11344 (N_11344,N_10659,N_10807);
nand U11345 (N_11345,N_10656,N_10542);
or U11346 (N_11346,N_10893,N_10804);
and U11347 (N_11347,N_10612,N_10618);
and U11348 (N_11348,N_10870,N_10676);
nand U11349 (N_11349,N_10612,N_10930);
nand U11350 (N_11350,N_10955,N_10823);
nor U11351 (N_11351,N_10938,N_10705);
and U11352 (N_11352,N_10809,N_10709);
nand U11353 (N_11353,N_10949,N_10556);
nor U11354 (N_11354,N_10574,N_10614);
nand U11355 (N_11355,N_10813,N_10818);
and U11356 (N_11356,N_10716,N_10910);
xnor U11357 (N_11357,N_10828,N_10990);
and U11358 (N_11358,N_10802,N_10909);
nand U11359 (N_11359,N_10868,N_10718);
or U11360 (N_11360,N_10891,N_10950);
or U11361 (N_11361,N_10589,N_10712);
or U11362 (N_11362,N_10734,N_10741);
and U11363 (N_11363,N_10510,N_10592);
nor U11364 (N_11364,N_10582,N_10722);
and U11365 (N_11365,N_10746,N_10740);
or U11366 (N_11366,N_10511,N_10541);
nor U11367 (N_11367,N_10615,N_10759);
or U11368 (N_11368,N_10616,N_10838);
or U11369 (N_11369,N_10744,N_10771);
nand U11370 (N_11370,N_10884,N_10755);
nor U11371 (N_11371,N_10936,N_10522);
or U11372 (N_11372,N_10665,N_10853);
nand U11373 (N_11373,N_10591,N_10584);
and U11374 (N_11374,N_10744,N_10823);
nand U11375 (N_11375,N_10981,N_10898);
nand U11376 (N_11376,N_10642,N_10550);
or U11377 (N_11377,N_10636,N_10792);
or U11378 (N_11378,N_10542,N_10525);
or U11379 (N_11379,N_10922,N_10921);
nor U11380 (N_11380,N_10624,N_10701);
nand U11381 (N_11381,N_10907,N_10766);
nor U11382 (N_11382,N_10966,N_10897);
xnor U11383 (N_11383,N_10698,N_10828);
nor U11384 (N_11384,N_10659,N_10797);
nand U11385 (N_11385,N_10698,N_10580);
and U11386 (N_11386,N_10501,N_10852);
nand U11387 (N_11387,N_10869,N_10566);
nand U11388 (N_11388,N_10698,N_10502);
nand U11389 (N_11389,N_10674,N_10917);
and U11390 (N_11390,N_10793,N_10713);
nand U11391 (N_11391,N_10911,N_10947);
nand U11392 (N_11392,N_10973,N_10862);
xor U11393 (N_11393,N_10755,N_10888);
xnor U11394 (N_11394,N_10640,N_10812);
nor U11395 (N_11395,N_10698,N_10678);
nor U11396 (N_11396,N_10639,N_10551);
nor U11397 (N_11397,N_10632,N_10909);
and U11398 (N_11398,N_10638,N_10683);
xnor U11399 (N_11399,N_10904,N_10589);
or U11400 (N_11400,N_10789,N_10585);
nand U11401 (N_11401,N_10732,N_10766);
nor U11402 (N_11402,N_10868,N_10962);
xor U11403 (N_11403,N_10647,N_10795);
and U11404 (N_11404,N_10660,N_10684);
or U11405 (N_11405,N_10501,N_10849);
or U11406 (N_11406,N_10901,N_10568);
nor U11407 (N_11407,N_10903,N_10635);
or U11408 (N_11408,N_10831,N_10957);
and U11409 (N_11409,N_10555,N_10935);
nand U11410 (N_11410,N_10669,N_10605);
or U11411 (N_11411,N_10636,N_10758);
nand U11412 (N_11412,N_10519,N_10729);
and U11413 (N_11413,N_10790,N_10848);
nand U11414 (N_11414,N_10984,N_10541);
nor U11415 (N_11415,N_10751,N_10540);
xnor U11416 (N_11416,N_10835,N_10752);
nor U11417 (N_11417,N_10522,N_10744);
or U11418 (N_11418,N_10986,N_10728);
nor U11419 (N_11419,N_10572,N_10828);
or U11420 (N_11420,N_10786,N_10808);
and U11421 (N_11421,N_10973,N_10745);
nand U11422 (N_11422,N_10906,N_10653);
or U11423 (N_11423,N_10804,N_10509);
xnor U11424 (N_11424,N_10841,N_10972);
or U11425 (N_11425,N_10913,N_10847);
and U11426 (N_11426,N_10639,N_10534);
nor U11427 (N_11427,N_10719,N_10596);
or U11428 (N_11428,N_10889,N_10779);
nor U11429 (N_11429,N_10563,N_10660);
and U11430 (N_11430,N_10730,N_10857);
nor U11431 (N_11431,N_10783,N_10551);
or U11432 (N_11432,N_10998,N_10718);
nor U11433 (N_11433,N_10777,N_10781);
nor U11434 (N_11434,N_10767,N_10688);
nor U11435 (N_11435,N_10658,N_10765);
or U11436 (N_11436,N_10968,N_10600);
or U11437 (N_11437,N_10585,N_10909);
xor U11438 (N_11438,N_10651,N_10766);
and U11439 (N_11439,N_10615,N_10764);
nand U11440 (N_11440,N_10686,N_10828);
or U11441 (N_11441,N_10530,N_10680);
or U11442 (N_11442,N_10593,N_10983);
nor U11443 (N_11443,N_10994,N_10966);
or U11444 (N_11444,N_10950,N_10928);
nand U11445 (N_11445,N_10973,N_10960);
nand U11446 (N_11446,N_10700,N_10876);
nand U11447 (N_11447,N_10865,N_10961);
nor U11448 (N_11448,N_10560,N_10827);
and U11449 (N_11449,N_10951,N_10586);
xnor U11450 (N_11450,N_10712,N_10569);
nand U11451 (N_11451,N_10743,N_10746);
or U11452 (N_11452,N_10903,N_10610);
or U11453 (N_11453,N_10916,N_10991);
nor U11454 (N_11454,N_10746,N_10791);
and U11455 (N_11455,N_10965,N_10650);
nand U11456 (N_11456,N_10895,N_10884);
nor U11457 (N_11457,N_10799,N_10552);
and U11458 (N_11458,N_10921,N_10798);
and U11459 (N_11459,N_10664,N_10917);
nor U11460 (N_11460,N_10686,N_10577);
xor U11461 (N_11461,N_10512,N_10791);
or U11462 (N_11462,N_10758,N_10719);
and U11463 (N_11463,N_10993,N_10737);
and U11464 (N_11464,N_10702,N_10778);
nor U11465 (N_11465,N_10609,N_10699);
nand U11466 (N_11466,N_10831,N_10950);
nor U11467 (N_11467,N_10921,N_10573);
xnor U11468 (N_11468,N_10916,N_10553);
nor U11469 (N_11469,N_10613,N_10575);
or U11470 (N_11470,N_10579,N_10939);
or U11471 (N_11471,N_10735,N_10774);
nand U11472 (N_11472,N_10759,N_10935);
and U11473 (N_11473,N_10600,N_10502);
xnor U11474 (N_11474,N_10827,N_10514);
and U11475 (N_11475,N_10756,N_10869);
nor U11476 (N_11476,N_10732,N_10814);
or U11477 (N_11477,N_10817,N_10847);
or U11478 (N_11478,N_10952,N_10746);
or U11479 (N_11479,N_10728,N_10914);
nor U11480 (N_11480,N_10500,N_10637);
nand U11481 (N_11481,N_10515,N_10731);
nor U11482 (N_11482,N_10512,N_10671);
and U11483 (N_11483,N_10597,N_10774);
and U11484 (N_11484,N_10584,N_10796);
nand U11485 (N_11485,N_10588,N_10502);
xnor U11486 (N_11486,N_10849,N_10803);
nor U11487 (N_11487,N_10788,N_10656);
or U11488 (N_11488,N_10867,N_10883);
nor U11489 (N_11489,N_10672,N_10538);
nand U11490 (N_11490,N_10828,N_10520);
and U11491 (N_11491,N_10557,N_10863);
nand U11492 (N_11492,N_10775,N_10825);
nor U11493 (N_11493,N_10717,N_10879);
or U11494 (N_11494,N_10638,N_10507);
and U11495 (N_11495,N_10946,N_10688);
nor U11496 (N_11496,N_10914,N_10611);
nor U11497 (N_11497,N_10687,N_10907);
or U11498 (N_11498,N_10691,N_10752);
xnor U11499 (N_11499,N_10557,N_10818);
or U11500 (N_11500,N_11465,N_11145);
nor U11501 (N_11501,N_11264,N_11336);
nor U11502 (N_11502,N_11082,N_11260);
nor U11503 (N_11503,N_11105,N_11249);
nor U11504 (N_11504,N_11030,N_11204);
or U11505 (N_11505,N_11166,N_11431);
nand U11506 (N_11506,N_11257,N_11339);
nor U11507 (N_11507,N_11287,N_11345);
or U11508 (N_11508,N_11319,N_11180);
nand U11509 (N_11509,N_11155,N_11347);
or U11510 (N_11510,N_11410,N_11366);
nor U11511 (N_11511,N_11131,N_11372);
or U11512 (N_11512,N_11058,N_11481);
and U11513 (N_11513,N_11296,N_11151);
or U11514 (N_11514,N_11054,N_11182);
and U11515 (N_11515,N_11087,N_11413);
or U11516 (N_11516,N_11380,N_11268);
nor U11517 (N_11517,N_11171,N_11235);
nor U11518 (N_11518,N_11224,N_11452);
nor U11519 (N_11519,N_11412,N_11229);
nand U11520 (N_11520,N_11346,N_11121);
nor U11521 (N_11521,N_11429,N_11027);
xor U11522 (N_11522,N_11395,N_11497);
nand U11523 (N_11523,N_11302,N_11222);
and U11524 (N_11524,N_11368,N_11373);
nor U11525 (N_11525,N_11169,N_11266);
nor U11526 (N_11526,N_11386,N_11147);
and U11527 (N_11527,N_11250,N_11281);
nand U11528 (N_11528,N_11459,N_11042);
and U11529 (N_11529,N_11137,N_11114);
nor U11530 (N_11530,N_11448,N_11053);
nand U11531 (N_11531,N_11478,N_11305);
nand U11532 (N_11532,N_11450,N_11378);
and U11533 (N_11533,N_11353,N_11449);
and U11534 (N_11534,N_11444,N_11103);
and U11535 (N_11535,N_11462,N_11437);
nor U11536 (N_11536,N_11496,N_11153);
nor U11537 (N_11537,N_11152,N_11390);
xor U11538 (N_11538,N_11328,N_11069);
nand U11539 (N_11539,N_11172,N_11021);
nand U11540 (N_11540,N_11022,N_11217);
nor U11541 (N_11541,N_11117,N_11464);
nand U11542 (N_11542,N_11005,N_11469);
and U11543 (N_11543,N_11015,N_11370);
or U11544 (N_11544,N_11486,N_11348);
nand U11545 (N_11545,N_11074,N_11205);
or U11546 (N_11546,N_11337,N_11426);
nor U11547 (N_11547,N_11394,N_11187);
or U11548 (N_11548,N_11091,N_11483);
nand U11549 (N_11549,N_11482,N_11280);
and U11550 (N_11550,N_11033,N_11416);
and U11551 (N_11551,N_11365,N_11292);
and U11552 (N_11552,N_11270,N_11026);
or U11553 (N_11553,N_11185,N_11445);
or U11554 (N_11554,N_11164,N_11421);
or U11555 (N_11555,N_11234,N_11245);
nor U11556 (N_11556,N_11094,N_11458);
and U11557 (N_11557,N_11442,N_11310);
or U11558 (N_11558,N_11084,N_11119);
or U11559 (N_11559,N_11181,N_11392);
nand U11560 (N_11560,N_11436,N_11133);
and U11561 (N_11561,N_11484,N_11175);
and U11562 (N_11562,N_11001,N_11008);
nand U11563 (N_11563,N_11309,N_11434);
nor U11564 (N_11564,N_11457,N_11326);
and U11565 (N_11565,N_11202,N_11396);
nor U11566 (N_11566,N_11269,N_11025);
and U11567 (N_11567,N_11212,N_11258);
or U11568 (N_11568,N_11439,N_11361);
xnor U11569 (N_11569,N_11067,N_11002);
nor U11570 (N_11570,N_11325,N_11401);
nand U11571 (N_11571,N_11188,N_11013);
xnor U11572 (N_11572,N_11165,N_11453);
nand U11573 (N_11573,N_11277,N_11354);
or U11574 (N_11574,N_11201,N_11350);
or U11575 (N_11575,N_11064,N_11099);
and U11576 (N_11576,N_11290,N_11324);
and U11577 (N_11577,N_11043,N_11112);
and U11578 (N_11578,N_11159,N_11400);
nor U11579 (N_11579,N_11016,N_11340);
and U11580 (N_11580,N_11475,N_11100);
nand U11581 (N_11581,N_11321,N_11037);
nand U11582 (N_11582,N_11075,N_11050);
nand U11583 (N_11583,N_11197,N_11375);
and U11584 (N_11584,N_11108,N_11456);
nand U11585 (N_11585,N_11192,N_11144);
and U11586 (N_11586,N_11077,N_11176);
nand U11587 (N_11587,N_11474,N_11428);
or U11588 (N_11588,N_11048,N_11070);
xor U11589 (N_11589,N_11113,N_11357);
and U11590 (N_11590,N_11190,N_11443);
nand U11591 (N_11591,N_11253,N_11473);
and U11592 (N_11592,N_11355,N_11062);
nor U11593 (N_11593,N_11298,N_11179);
or U11594 (N_11594,N_11383,N_11276);
nor U11595 (N_11595,N_11031,N_11228);
xor U11596 (N_11596,N_11332,N_11300);
nor U11597 (N_11597,N_11135,N_11384);
or U11598 (N_11598,N_11214,N_11402);
xnor U11599 (N_11599,N_11291,N_11265);
xnor U11600 (N_11600,N_11011,N_11338);
xnor U11601 (N_11601,N_11167,N_11284);
nor U11602 (N_11602,N_11476,N_11352);
and U11603 (N_11603,N_11389,N_11393);
nand U11604 (N_11604,N_11415,N_11238);
nand U11605 (N_11605,N_11494,N_11134);
nand U11606 (N_11606,N_11095,N_11498);
nand U11607 (N_11607,N_11195,N_11143);
and U11608 (N_11608,N_11041,N_11407);
nor U11609 (N_11609,N_11161,N_11499);
and U11610 (N_11610,N_11301,N_11023);
xor U11611 (N_11611,N_11071,N_11255);
xnor U11612 (N_11612,N_11262,N_11425);
or U11613 (N_11613,N_11221,N_11460);
nand U11614 (N_11614,N_11010,N_11308);
or U11615 (N_11615,N_11237,N_11492);
and U11616 (N_11616,N_11139,N_11009);
and U11617 (N_11617,N_11274,N_11111);
nand U11618 (N_11618,N_11120,N_11156);
and U11619 (N_11619,N_11468,N_11068);
or U11620 (N_11620,N_11312,N_11126);
and U11621 (N_11621,N_11059,N_11422);
nand U11622 (N_11622,N_11433,N_11404);
and U11623 (N_11623,N_11294,N_11136);
or U11624 (N_11624,N_11200,N_11073);
and U11625 (N_11625,N_11173,N_11186);
or U11626 (N_11626,N_11435,N_11122);
and U11627 (N_11627,N_11351,N_11349);
or U11628 (N_11628,N_11331,N_11055);
nor U11629 (N_11629,N_11007,N_11024);
nand U11630 (N_11630,N_11230,N_11189);
nor U11631 (N_11631,N_11049,N_11261);
nand U11632 (N_11632,N_11226,N_11303);
nor U11633 (N_11633,N_11004,N_11256);
nor U11634 (N_11634,N_11273,N_11223);
nor U11635 (N_11635,N_11216,N_11018);
or U11636 (N_11636,N_11275,N_11382);
and U11637 (N_11637,N_11391,N_11342);
and U11638 (N_11638,N_11109,N_11142);
nor U11639 (N_11639,N_11220,N_11414);
nand U11640 (N_11640,N_11177,N_11304);
nor U11641 (N_11641,N_11129,N_11330);
nand U11642 (N_11642,N_11032,N_11248);
xor U11643 (N_11643,N_11388,N_11405);
or U11644 (N_11644,N_11210,N_11323);
or U11645 (N_11645,N_11282,N_11060);
and U11646 (N_11646,N_11398,N_11063);
and U11647 (N_11647,N_11034,N_11254);
xnor U11648 (N_11648,N_11019,N_11146);
and U11649 (N_11649,N_11000,N_11236);
and U11650 (N_11650,N_11219,N_11397);
and U11651 (N_11651,N_11140,N_11079);
nand U11652 (N_11652,N_11241,N_11012);
or U11653 (N_11653,N_11039,N_11430);
or U11654 (N_11654,N_11411,N_11399);
or U11655 (N_11655,N_11313,N_11097);
nand U11656 (N_11656,N_11006,N_11316);
nand U11657 (N_11657,N_11446,N_11359);
or U11658 (N_11658,N_11240,N_11183);
xor U11659 (N_11659,N_11409,N_11329);
nand U11660 (N_11660,N_11174,N_11490);
and U11661 (N_11661,N_11198,N_11206);
or U11662 (N_11662,N_11440,N_11066);
nor U11663 (N_11663,N_11191,N_11364);
xor U11664 (N_11664,N_11477,N_11061);
nor U11665 (N_11665,N_11267,N_11118);
and U11666 (N_11666,N_11028,N_11045);
or U11667 (N_11667,N_11078,N_11285);
or U11668 (N_11668,N_11093,N_11343);
or U11669 (N_11669,N_11252,N_11488);
or U11670 (N_11670,N_11208,N_11056);
nand U11671 (N_11671,N_11088,N_11227);
nor U11672 (N_11672,N_11115,N_11242);
nor U11673 (N_11673,N_11184,N_11090);
and U11674 (N_11674,N_11320,N_11215);
or U11675 (N_11675,N_11288,N_11318);
or U11676 (N_11676,N_11017,N_11376);
or U11677 (N_11677,N_11387,N_11107);
and U11678 (N_11678,N_11125,N_11403);
and U11679 (N_11679,N_11193,N_11051);
nand U11680 (N_11680,N_11038,N_11480);
nor U11681 (N_11681,N_11160,N_11283);
and U11682 (N_11682,N_11072,N_11209);
or U11683 (N_11683,N_11315,N_11489);
or U11684 (N_11684,N_11154,N_11295);
or U11685 (N_11685,N_11232,N_11096);
nand U11686 (N_11686,N_11035,N_11307);
nor U11687 (N_11687,N_11451,N_11057);
and U11688 (N_11688,N_11196,N_11344);
and U11689 (N_11689,N_11106,N_11044);
nand U11690 (N_11690,N_11132,N_11263);
and U11691 (N_11691,N_11163,N_11385);
nand U11692 (N_11692,N_11279,N_11334);
nor U11693 (N_11693,N_11360,N_11243);
nand U11694 (N_11694,N_11029,N_11149);
and U11695 (N_11695,N_11487,N_11085);
or U11696 (N_11696,N_11363,N_11341);
or U11697 (N_11697,N_11374,N_11116);
xnor U11698 (N_11698,N_11225,N_11046);
or U11699 (N_11699,N_11211,N_11369);
nor U11700 (N_11700,N_11362,N_11239);
nand U11701 (N_11701,N_11485,N_11199);
or U11702 (N_11702,N_11246,N_11178);
xor U11703 (N_11703,N_11278,N_11371);
xor U11704 (N_11704,N_11424,N_11148);
xnor U11705 (N_11705,N_11076,N_11098);
or U11706 (N_11706,N_11020,N_11272);
nand U11707 (N_11707,N_11286,N_11333);
or U11708 (N_11708,N_11317,N_11127);
nand U11709 (N_11709,N_11493,N_11311);
xnor U11710 (N_11710,N_11419,N_11138);
and U11711 (N_11711,N_11259,N_11104);
nor U11712 (N_11712,N_11089,N_11470);
and U11713 (N_11713,N_11438,N_11157);
nand U11714 (N_11714,N_11463,N_11335);
and U11715 (N_11715,N_11101,N_11432);
nor U11716 (N_11716,N_11322,N_11036);
xor U11717 (N_11717,N_11003,N_11420);
nor U11718 (N_11718,N_11377,N_11306);
and U11719 (N_11719,N_11158,N_11454);
nand U11720 (N_11720,N_11231,N_11213);
or U11721 (N_11721,N_11130,N_11297);
nor U11722 (N_11722,N_11110,N_11471);
nor U11723 (N_11723,N_11080,N_11356);
or U11724 (N_11724,N_11251,N_11170);
nand U11725 (N_11725,N_11014,N_11083);
nand U11726 (N_11726,N_11408,N_11207);
nor U11727 (N_11727,N_11367,N_11141);
xor U11728 (N_11728,N_11427,N_11289);
nor U11729 (N_11729,N_11081,N_11461);
nor U11730 (N_11730,N_11293,N_11086);
or U11731 (N_11731,N_11092,N_11065);
and U11732 (N_11732,N_11040,N_11455);
nor U11733 (N_11733,N_11271,N_11467);
nor U11734 (N_11734,N_11491,N_11441);
and U11735 (N_11735,N_11406,N_11203);
nor U11736 (N_11736,N_11327,N_11218);
xnor U11737 (N_11737,N_11123,N_11479);
nand U11738 (N_11738,N_11233,N_11381);
xnor U11739 (N_11739,N_11299,N_11244);
xor U11740 (N_11740,N_11472,N_11194);
or U11741 (N_11741,N_11423,N_11124);
nor U11742 (N_11742,N_11447,N_11314);
nand U11743 (N_11743,N_11358,N_11495);
and U11744 (N_11744,N_11162,N_11102);
or U11745 (N_11745,N_11168,N_11418);
and U11746 (N_11746,N_11128,N_11379);
or U11747 (N_11747,N_11417,N_11150);
nor U11748 (N_11748,N_11466,N_11247);
or U11749 (N_11749,N_11052,N_11047);
nand U11750 (N_11750,N_11167,N_11127);
nand U11751 (N_11751,N_11437,N_11032);
nand U11752 (N_11752,N_11372,N_11094);
nand U11753 (N_11753,N_11028,N_11333);
xor U11754 (N_11754,N_11393,N_11323);
nand U11755 (N_11755,N_11148,N_11328);
nor U11756 (N_11756,N_11319,N_11342);
or U11757 (N_11757,N_11176,N_11119);
nor U11758 (N_11758,N_11105,N_11455);
nand U11759 (N_11759,N_11439,N_11404);
and U11760 (N_11760,N_11118,N_11431);
and U11761 (N_11761,N_11434,N_11181);
or U11762 (N_11762,N_11374,N_11258);
and U11763 (N_11763,N_11365,N_11367);
or U11764 (N_11764,N_11267,N_11484);
nor U11765 (N_11765,N_11366,N_11078);
and U11766 (N_11766,N_11017,N_11246);
nor U11767 (N_11767,N_11228,N_11062);
and U11768 (N_11768,N_11340,N_11316);
and U11769 (N_11769,N_11491,N_11090);
and U11770 (N_11770,N_11177,N_11341);
nor U11771 (N_11771,N_11372,N_11042);
or U11772 (N_11772,N_11132,N_11429);
or U11773 (N_11773,N_11003,N_11263);
nand U11774 (N_11774,N_11204,N_11264);
or U11775 (N_11775,N_11163,N_11390);
nand U11776 (N_11776,N_11468,N_11318);
xor U11777 (N_11777,N_11084,N_11364);
xnor U11778 (N_11778,N_11181,N_11179);
and U11779 (N_11779,N_11107,N_11469);
and U11780 (N_11780,N_11433,N_11320);
xor U11781 (N_11781,N_11188,N_11498);
nor U11782 (N_11782,N_11178,N_11245);
nand U11783 (N_11783,N_11356,N_11339);
xor U11784 (N_11784,N_11493,N_11020);
nor U11785 (N_11785,N_11144,N_11121);
and U11786 (N_11786,N_11331,N_11032);
nor U11787 (N_11787,N_11076,N_11127);
and U11788 (N_11788,N_11309,N_11103);
or U11789 (N_11789,N_11412,N_11398);
xor U11790 (N_11790,N_11448,N_11228);
nor U11791 (N_11791,N_11428,N_11346);
xor U11792 (N_11792,N_11054,N_11417);
and U11793 (N_11793,N_11055,N_11438);
nor U11794 (N_11794,N_11221,N_11361);
and U11795 (N_11795,N_11130,N_11066);
nor U11796 (N_11796,N_11472,N_11070);
and U11797 (N_11797,N_11230,N_11407);
or U11798 (N_11798,N_11479,N_11216);
or U11799 (N_11799,N_11371,N_11091);
nor U11800 (N_11800,N_11356,N_11001);
nor U11801 (N_11801,N_11107,N_11259);
xnor U11802 (N_11802,N_11457,N_11464);
xor U11803 (N_11803,N_11181,N_11166);
or U11804 (N_11804,N_11147,N_11107);
and U11805 (N_11805,N_11471,N_11257);
nor U11806 (N_11806,N_11084,N_11100);
nor U11807 (N_11807,N_11055,N_11132);
and U11808 (N_11808,N_11005,N_11037);
or U11809 (N_11809,N_11191,N_11325);
xor U11810 (N_11810,N_11424,N_11194);
and U11811 (N_11811,N_11386,N_11056);
and U11812 (N_11812,N_11274,N_11344);
nor U11813 (N_11813,N_11032,N_11170);
and U11814 (N_11814,N_11178,N_11370);
or U11815 (N_11815,N_11209,N_11302);
nor U11816 (N_11816,N_11481,N_11290);
or U11817 (N_11817,N_11032,N_11207);
xnor U11818 (N_11818,N_11049,N_11093);
and U11819 (N_11819,N_11382,N_11425);
xor U11820 (N_11820,N_11000,N_11235);
or U11821 (N_11821,N_11359,N_11221);
xnor U11822 (N_11822,N_11141,N_11007);
or U11823 (N_11823,N_11119,N_11232);
nor U11824 (N_11824,N_11408,N_11446);
nor U11825 (N_11825,N_11267,N_11328);
xor U11826 (N_11826,N_11002,N_11056);
nor U11827 (N_11827,N_11230,N_11449);
nand U11828 (N_11828,N_11357,N_11316);
and U11829 (N_11829,N_11441,N_11304);
nand U11830 (N_11830,N_11232,N_11085);
xnor U11831 (N_11831,N_11319,N_11400);
and U11832 (N_11832,N_11029,N_11141);
and U11833 (N_11833,N_11211,N_11379);
or U11834 (N_11834,N_11138,N_11316);
nand U11835 (N_11835,N_11209,N_11417);
xor U11836 (N_11836,N_11458,N_11426);
nand U11837 (N_11837,N_11333,N_11045);
xnor U11838 (N_11838,N_11068,N_11039);
nor U11839 (N_11839,N_11016,N_11258);
nand U11840 (N_11840,N_11344,N_11387);
and U11841 (N_11841,N_11490,N_11164);
or U11842 (N_11842,N_11311,N_11345);
nor U11843 (N_11843,N_11269,N_11427);
or U11844 (N_11844,N_11265,N_11299);
nand U11845 (N_11845,N_11184,N_11401);
or U11846 (N_11846,N_11374,N_11094);
or U11847 (N_11847,N_11053,N_11150);
nand U11848 (N_11848,N_11046,N_11464);
or U11849 (N_11849,N_11034,N_11079);
or U11850 (N_11850,N_11188,N_11248);
nor U11851 (N_11851,N_11470,N_11083);
or U11852 (N_11852,N_11490,N_11446);
nand U11853 (N_11853,N_11423,N_11180);
nor U11854 (N_11854,N_11123,N_11170);
or U11855 (N_11855,N_11012,N_11171);
nor U11856 (N_11856,N_11064,N_11265);
and U11857 (N_11857,N_11041,N_11063);
nor U11858 (N_11858,N_11452,N_11104);
or U11859 (N_11859,N_11322,N_11485);
and U11860 (N_11860,N_11195,N_11260);
nand U11861 (N_11861,N_11070,N_11237);
and U11862 (N_11862,N_11229,N_11463);
or U11863 (N_11863,N_11298,N_11030);
nor U11864 (N_11864,N_11105,N_11234);
nor U11865 (N_11865,N_11194,N_11027);
and U11866 (N_11866,N_11421,N_11301);
xor U11867 (N_11867,N_11414,N_11207);
or U11868 (N_11868,N_11054,N_11343);
or U11869 (N_11869,N_11130,N_11478);
nand U11870 (N_11870,N_11073,N_11002);
nand U11871 (N_11871,N_11060,N_11201);
nand U11872 (N_11872,N_11261,N_11183);
nand U11873 (N_11873,N_11484,N_11034);
or U11874 (N_11874,N_11173,N_11079);
nand U11875 (N_11875,N_11124,N_11492);
nand U11876 (N_11876,N_11011,N_11411);
nand U11877 (N_11877,N_11003,N_11034);
xor U11878 (N_11878,N_11298,N_11290);
xnor U11879 (N_11879,N_11265,N_11219);
xnor U11880 (N_11880,N_11470,N_11367);
and U11881 (N_11881,N_11300,N_11375);
xor U11882 (N_11882,N_11495,N_11410);
nand U11883 (N_11883,N_11468,N_11497);
nand U11884 (N_11884,N_11145,N_11298);
nand U11885 (N_11885,N_11371,N_11050);
or U11886 (N_11886,N_11370,N_11093);
nand U11887 (N_11887,N_11343,N_11291);
and U11888 (N_11888,N_11116,N_11496);
or U11889 (N_11889,N_11070,N_11159);
and U11890 (N_11890,N_11314,N_11308);
nor U11891 (N_11891,N_11327,N_11312);
and U11892 (N_11892,N_11315,N_11497);
or U11893 (N_11893,N_11317,N_11051);
and U11894 (N_11894,N_11254,N_11410);
nor U11895 (N_11895,N_11366,N_11010);
and U11896 (N_11896,N_11415,N_11047);
and U11897 (N_11897,N_11081,N_11360);
nor U11898 (N_11898,N_11295,N_11175);
nand U11899 (N_11899,N_11143,N_11312);
nor U11900 (N_11900,N_11139,N_11062);
or U11901 (N_11901,N_11122,N_11414);
xor U11902 (N_11902,N_11475,N_11081);
and U11903 (N_11903,N_11118,N_11268);
nor U11904 (N_11904,N_11071,N_11070);
nor U11905 (N_11905,N_11330,N_11126);
and U11906 (N_11906,N_11437,N_11029);
nand U11907 (N_11907,N_11109,N_11097);
and U11908 (N_11908,N_11470,N_11469);
nand U11909 (N_11909,N_11421,N_11358);
nor U11910 (N_11910,N_11006,N_11166);
xnor U11911 (N_11911,N_11449,N_11164);
nand U11912 (N_11912,N_11007,N_11405);
and U11913 (N_11913,N_11160,N_11180);
or U11914 (N_11914,N_11159,N_11287);
nor U11915 (N_11915,N_11170,N_11292);
nor U11916 (N_11916,N_11080,N_11284);
and U11917 (N_11917,N_11076,N_11397);
nor U11918 (N_11918,N_11185,N_11230);
nor U11919 (N_11919,N_11079,N_11328);
or U11920 (N_11920,N_11217,N_11184);
nand U11921 (N_11921,N_11342,N_11296);
or U11922 (N_11922,N_11175,N_11050);
or U11923 (N_11923,N_11159,N_11259);
or U11924 (N_11924,N_11429,N_11293);
nor U11925 (N_11925,N_11257,N_11242);
nor U11926 (N_11926,N_11313,N_11480);
nand U11927 (N_11927,N_11219,N_11327);
or U11928 (N_11928,N_11160,N_11247);
or U11929 (N_11929,N_11153,N_11301);
and U11930 (N_11930,N_11244,N_11470);
and U11931 (N_11931,N_11465,N_11055);
nand U11932 (N_11932,N_11162,N_11011);
nor U11933 (N_11933,N_11228,N_11041);
nor U11934 (N_11934,N_11366,N_11287);
nand U11935 (N_11935,N_11026,N_11457);
and U11936 (N_11936,N_11284,N_11289);
and U11937 (N_11937,N_11281,N_11127);
nor U11938 (N_11938,N_11220,N_11224);
or U11939 (N_11939,N_11254,N_11319);
nand U11940 (N_11940,N_11210,N_11296);
and U11941 (N_11941,N_11113,N_11420);
xor U11942 (N_11942,N_11088,N_11167);
or U11943 (N_11943,N_11062,N_11391);
nor U11944 (N_11944,N_11141,N_11300);
or U11945 (N_11945,N_11389,N_11429);
or U11946 (N_11946,N_11043,N_11208);
and U11947 (N_11947,N_11486,N_11492);
and U11948 (N_11948,N_11401,N_11472);
nor U11949 (N_11949,N_11104,N_11456);
nor U11950 (N_11950,N_11469,N_11360);
xor U11951 (N_11951,N_11419,N_11166);
and U11952 (N_11952,N_11238,N_11354);
or U11953 (N_11953,N_11150,N_11147);
or U11954 (N_11954,N_11237,N_11087);
nor U11955 (N_11955,N_11323,N_11013);
or U11956 (N_11956,N_11188,N_11224);
and U11957 (N_11957,N_11246,N_11008);
and U11958 (N_11958,N_11367,N_11455);
and U11959 (N_11959,N_11381,N_11311);
nand U11960 (N_11960,N_11150,N_11208);
nor U11961 (N_11961,N_11076,N_11494);
nor U11962 (N_11962,N_11473,N_11448);
xnor U11963 (N_11963,N_11497,N_11436);
and U11964 (N_11964,N_11069,N_11393);
and U11965 (N_11965,N_11073,N_11334);
xnor U11966 (N_11966,N_11335,N_11282);
nor U11967 (N_11967,N_11052,N_11418);
nor U11968 (N_11968,N_11484,N_11054);
nand U11969 (N_11969,N_11056,N_11026);
and U11970 (N_11970,N_11483,N_11346);
nor U11971 (N_11971,N_11042,N_11184);
nand U11972 (N_11972,N_11472,N_11491);
nand U11973 (N_11973,N_11332,N_11483);
and U11974 (N_11974,N_11125,N_11246);
nand U11975 (N_11975,N_11397,N_11194);
and U11976 (N_11976,N_11383,N_11412);
or U11977 (N_11977,N_11285,N_11124);
nand U11978 (N_11978,N_11018,N_11060);
and U11979 (N_11979,N_11007,N_11014);
nand U11980 (N_11980,N_11216,N_11458);
or U11981 (N_11981,N_11086,N_11230);
nand U11982 (N_11982,N_11313,N_11399);
nor U11983 (N_11983,N_11411,N_11480);
nor U11984 (N_11984,N_11398,N_11097);
and U11985 (N_11985,N_11005,N_11408);
and U11986 (N_11986,N_11132,N_11157);
nand U11987 (N_11987,N_11155,N_11383);
and U11988 (N_11988,N_11344,N_11424);
or U11989 (N_11989,N_11007,N_11482);
nand U11990 (N_11990,N_11222,N_11348);
or U11991 (N_11991,N_11264,N_11458);
nor U11992 (N_11992,N_11108,N_11259);
xnor U11993 (N_11993,N_11186,N_11222);
and U11994 (N_11994,N_11174,N_11229);
or U11995 (N_11995,N_11443,N_11494);
and U11996 (N_11996,N_11120,N_11075);
or U11997 (N_11997,N_11062,N_11101);
and U11998 (N_11998,N_11481,N_11238);
or U11999 (N_11999,N_11111,N_11069);
nand U12000 (N_12000,N_11809,N_11878);
or U12001 (N_12001,N_11978,N_11858);
nor U12002 (N_12002,N_11576,N_11646);
nor U12003 (N_12003,N_11928,N_11921);
nand U12004 (N_12004,N_11746,N_11521);
nand U12005 (N_12005,N_11630,N_11572);
nor U12006 (N_12006,N_11694,N_11654);
xnor U12007 (N_12007,N_11670,N_11527);
xor U12008 (N_12008,N_11591,N_11951);
nand U12009 (N_12009,N_11692,N_11816);
nand U12010 (N_12010,N_11782,N_11536);
nand U12011 (N_12011,N_11737,N_11733);
nor U12012 (N_12012,N_11698,N_11947);
or U12013 (N_12013,N_11941,N_11881);
or U12014 (N_12014,N_11587,N_11803);
nand U12015 (N_12015,N_11865,N_11937);
nand U12016 (N_12016,N_11853,N_11915);
or U12017 (N_12017,N_11934,N_11609);
nor U12018 (N_12018,N_11965,N_11776);
nor U12019 (N_12019,N_11907,N_11815);
or U12020 (N_12020,N_11932,N_11872);
and U12021 (N_12021,N_11952,N_11665);
or U12022 (N_12022,N_11603,N_11671);
and U12023 (N_12023,N_11677,N_11756);
nor U12024 (N_12024,N_11987,N_11807);
nor U12025 (N_12025,N_11675,N_11653);
nand U12026 (N_12026,N_11613,N_11571);
and U12027 (N_12027,N_11574,N_11836);
or U12028 (N_12028,N_11797,N_11908);
and U12029 (N_12029,N_11819,N_11844);
xnor U12030 (N_12030,N_11993,N_11939);
nand U12031 (N_12031,N_11989,N_11940);
xor U12032 (N_12032,N_11863,N_11829);
nor U12033 (N_12033,N_11718,N_11680);
xnor U12034 (N_12034,N_11531,N_11559);
and U12035 (N_12035,N_11754,N_11599);
nand U12036 (N_12036,N_11592,N_11784);
nand U12037 (N_12037,N_11795,N_11641);
nor U12038 (N_12038,N_11847,N_11936);
or U12039 (N_12039,N_11780,N_11873);
nor U12040 (N_12040,N_11808,N_11799);
or U12041 (N_12041,N_11667,N_11787);
and U12042 (N_12042,N_11535,N_11501);
or U12043 (N_12043,N_11734,N_11731);
xnor U12044 (N_12044,N_11639,N_11842);
and U12045 (N_12045,N_11553,N_11607);
nor U12046 (N_12046,N_11906,N_11648);
or U12047 (N_12047,N_11598,N_11973);
nor U12048 (N_12048,N_11685,N_11916);
xor U12049 (N_12049,N_11988,N_11569);
nor U12050 (N_12050,N_11831,N_11511);
nand U12051 (N_12051,N_11625,N_11583);
and U12052 (N_12052,N_11614,N_11699);
or U12053 (N_12053,N_11732,N_11505);
xor U12054 (N_12054,N_11738,N_11683);
nor U12055 (N_12055,N_11517,N_11977);
and U12056 (N_12056,N_11918,N_11870);
nor U12057 (N_12057,N_11768,N_11530);
or U12058 (N_12058,N_11770,N_11860);
nand U12059 (N_12059,N_11550,N_11626);
nor U12060 (N_12060,N_11659,N_11628);
nor U12061 (N_12061,N_11636,N_11538);
xnor U12062 (N_12062,N_11741,N_11929);
nor U12063 (N_12063,N_11760,N_11752);
nor U12064 (N_12064,N_11961,N_11589);
or U12065 (N_12065,N_11769,N_11856);
or U12066 (N_12066,N_11931,N_11975);
nor U12067 (N_12067,N_11946,N_11642);
or U12068 (N_12068,N_11739,N_11850);
nor U12069 (N_12069,N_11689,N_11990);
or U12070 (N_12070,N_11830,N_11657);
nand U12071 (N_12071,N_11875,N_11664);
or U12072 (N_12072,N_11621,N_11820);
xnor U12073 (N_12073,N_11658,N_11834);
nand U12074 (N_12074,N_11637,N_11917);
or U12075 (N_12075,N_11516,N_11673);
xor U12076 (N_12076,N_11982,N_11845);
and U12077 (N_12077,N_11925,N_11660);
nor U12078 (N_12078,N_11611,N_11682);
and U12079 (N_12079,N_11502,N_11790);
nor U12080 (N_12080,N_11676,N_11837);
or U12081 (N_12081,N_11522,N_11943);
xor U12082 (N_12082,N_11500,N_11547);
nor U12083 (N_12083,N_11712,N_11529);
nor U12084 (N_12084,N_11827,N_11761);
nor U12085 (N_12085,N_11736,N_11714);
and U12086 (N_12086,N_11608,N_11744);
and U12087 (N_12087,N_11833,N_11693);
or U12088 (N_12088,N_11801,N_11980);
or U12089 (N_12089,N_11606,N_11713);
nor U12090 (N_12090,N_11528,N_11955);
and U12091 (N_12091,N_11866,N_11730);
nand U12092 (N_12092,N_11696,N_11617);
nor U12093 (N_12093,N_11838,N_11788);
nor U12094 (N_12094,N_11588,N_11579);
or U12095 (N_12095,N_11890,N_11884);
nand U12096 (N_12096,N_11781,N_11892);
or U12097 (N_12097,N_11891,N_11524);
or U12098 (N_12098,N_11767,N_11810);
nand U12099 (N_12099,N_11519,N_11513);
or U12100 (N_12100,N_11706,N_11909);
xnor U12101 (N_12101,N_11817,N_11930);
nor U12102 (N_12102,N_11899,N_11604);
or U12103 (N_12103,N_11554,N_11555);
and U12104 (N_12104,N_11805,N_11632);
nand U12105 (N_12105,N_11794,N_11888);
and U12106 (N_12106,N_11526,N_11627);
or U12107 (N_12107,N_11605,N_11610);
xnor U12108 (N_12108,N_11710,N_11766);
or U12109 (N_12109,N_11887,N_11745);
or U12110 (N_12110,N_11893,N_11723);
and U12111 (N_12111,N_11825,N_11911);
or U12112 (N_12112,N_11813,N_11577);
nand U12113 (N_12113,N_11974,N_11691);
nor U12114 (N_12114,N_11601,N_11668);
nor U12115 (N_12115,N_11945,N_11772);
and U12116 (N_12116,N_11570,N_11966);
and U12117 (N_12117,N_11635,N_11624);
nand U12118 (N_12118,N_11902,N_11775);
nand U12119 (N_12119,N_11968,N_11715);
nor U12120 (N_12120,N_11541,N_11523);
and U12121 (N_12121,N_11962,N_11949);
nand U12122 (N_12122,N_11688,N_11904);
nor U12123 (N_12123,N_11765,N_11789);
or U12124 (N_12124,N_11512,N_11562);
nand U12125 (N_12125,N_11996,N_11542);
and U12126 (N_12126,N_11864,N_11645);
nand U12127 (N_12127,N_11868,N_11901);
nor U12128 (N_12128,N_11859,N_11534);
nand U12129 (N_12129,N_11747,N_11631);
nor U12130 (N_12130,N_11594,N_11634);
nand U12131 (N_12131,N_11964,N_11735);
nand U12132 (N_12132,N_11620,N_11652);
and U12133 (N_12133,N_11832,N_11972);
and U12134 (N_12134,N_11774,N_11567);
or U12135 (N_12135,N_11950,N_11959);
xnor U12136 (N_12136,N_11679,N_11618);
and U12137 (N_12137,N_11509,N_11581);
and U12138 (N_12138,N_11869,N_11725);
nand U12139 (N_12139,N_11672,N_11882);
nor U12140 (N_12140,N_11661,N_11848);
and U12141 (N_12141,N_11721,N_11565);
nor U12142 (N_12142,N_11649,N_11716);
or U12143 (N_12143,N_11508,N_11926);
nor U12144 (N_12144,N_11690,N_11806);
or U12145 (N_12145,N_11897,N_11783);
nor U12146 (N_12146,N_11702,N_11709);
nand U12147 (N_12147,N_11840,N_11584);
and U12148 (N_12148,N_11963,N_11729);
nand U12149 (N_12149,N_11826,N_11503);
and U12150 (N_12150,N_11506,N_11724);
and U12151 (N_12151,N_11976,N_11879);
nand U12152 (N_12152,N_11995,N_11666);
and U12153 (N_12153,N_11900,N_11701);
and U12154 (N_12154,N_11755,N_11678);
nor U12155 (N_12155,N_11898,N_11811);
and U12156 (N_12156,N_11786,N_11719);
or U12157 (N_12157,N_11684,N_11674);
nand U12158 (N_12158,N_11533,N_11944);
and U12159 (N_12159,N_11507,N_11750);
or U12160 (N_12160,N_11985,N_11686);
or U12161 (N_12161,N_11969,N_11851);
or U12162 (N_12162,N_11981,N_11796);
and U12163 (N_12163,N_11753,N_11586);
xnor U12164 (N_12164,N_11785,N_11956);
nor U12165 (N_12165,N_11935,N_11896);
and U12166 (N_12166,N_11854,N_11551);
nor U12167 (N_12167,N_11913,N_11800);
xor U12168 (N_12168,N_11757,N_11862);
nand U12169 (N_12169,N_11532,N_11705);
or U12170 (N_12170,N_11843,N_11759);
xnor U12171 (N_12171,N_11580,N_11793);
nand U12172 (N_12172,N_11556,N_11999);
nand U12173 (N_12173,N_11812,N_11595);
nand U12174 (N_12174,N_11994,N_11984);
xor U12175 (N_12175,N_11504,N_11773);
nand U12176 (N_12176,N_11841,N_11644);
nand U12177 (N_12177,N_11564,N_11633);
or U12178 (N_12178,N_11590,N_11623);
xor U12179 (N_12179,N_11798,N_11728);
nand U12180 (N_12180,N_11711,N_11707);
and U12181 (N_12181,N_11883,N_11905);
or U12182 (N_12182,N_11991,N_11877);
and U12183 (N_12183,N_11933,N_11663);
or U12184 (N_12184,N_11640,N_11600);
or U12185 (N_12185,N_11764,N_11566);
xnor U12186 (N_12186,N_11818,N_11704);
nor U12187 (N_12187,N_11740,N_11669);
nand U12188 (N_12188,N_11717,N_11697);
and U12189 (N_12189,N_11593,N_11920);
or U12190 (N_12190,N_11986,N_11543);
xor U12191 (N_12191,N_11828,N_11681);
or U12192 (N_12192,N_11792,N_11616);
nand U12193 (N_12193,N_11612,N_11839);
or U12194 (N_12194,N_11824,N_11722);
nor U12195 (N_12195,N_11578,N_11849);
and U12196 (N_12196,N_11514,N_11914);
nor U12197 (N_12197,N_11544,N_11938);
nand U12198 (N_12198,N_11763,N_11537);
nor U12199 (N_12199,N_11983,N_11855);
xor U12200 (N_12200,N_11557,N_11703);
nor U12201 (N_12201,N_11742,N_11924);
nand U12202 (N_12202,N_11771,N_11662);
or U12203 (N_12203,N_11561,N_11510);
nand U12204 (N_12204,N_11823,N_11560);
nor U12205 (N_12205,N_11802,N_11971);
nand U12206 (N_12206,N_11727,N_11585);
or U12207 (N_12207,N_11922,N_11814);
nor U12208 (N_12208,N_11546,N_11846);
and U12209 (N_12209,N_11778,N_11643);
nor U12210 (N_12210,N_11549,N_11548);
and U12211 (N_12211,N_11720,N_11582);
or U12212 (N_12212,N_11835,N_11619);
nor U12213 (N_12213,N_11602,N_11762);
nand U12214 (N_12214,N_11857,N_11910);
nor U12215 (N_12215,N_11997,N_11708);
and U12216 (N_12216,N_11948,N_11743);
nand U12217 (N_12217,N_11923,N_11545);
xor U12218 (N_12218,N_11954,N_11960);
nor U12219 (N_12219,N_11876,N_11539);
nand U12220 (N_12220,N_11552,N_11871);
and U12221 (N_12221,N_11779,N_11615);
nand U12222 (N_12222,N_11953,N_11687);
or U12223 (N_12223,N_11656,N_11927);
or U12224 (N_12224,N_11967,N_11970);
or U12225 (N_12225,N_11821,N_11700);
and U12226 (N_12226,N_11726,N_11596);
or U12227 (N_12227,N_11650,N_11748);
xor U12228 (N_12228,N_11758,N_11992);
xor U12229 (N_12229,N_11651,N_11749);
nand U12230 (N_12230,N_11894,N_11568);
or U12231 (N_12231,N_11558,N_11861);
and U12232 (N_12232,N_11880,N_11942);
or U12233 (N_12233,N_11919,N_11518);
or U12234 (N_12234,N_11777,N_11804);
and U12235 (N_12235,N_11515,N_11822);
and U12236 (N_12236,N_11958,N_11573);
or U12237 (N_12237,N_11525,N_11751);
or U12238 (N_12238,N_11695,N_11889);
and U12239 (N_12239,N_11563,N_11575);
and U12240 (N_12240,N_11912,N_11957);
nor U12241 (N_12241,N_11867,N_11540);
nand U12242 (N_12242,N_11979,N_11629);
nand U12243 (N_12243,N_11886,N_11852);
or U12244 (N_12244,N_11647,N_11791);
xor U12245 (N_12245,N_11597,N_11903);
and U12246 (N_12246,N_11655,N_11638);
nor U12247 (N_12247,N_11874,N_11622);
and U12248 (N_12248,N_11520,N_11998);
nand U12249 (N_12249,N_11885,N_11895);
xnor U12250 (N_12250,N_11892,N_11795);
nand U12251 (N_12251,N_11889,N_11758);
nand U12252 (N_12252,N_11800,N_11864);
or U12253 (N_12253,N_11780,N_11638);
xor U12254 (N_12254,N_11550,N_11534);
xor U12255 (N_12255,N_11609,N_11627);
or U12256 (N_12256,N_11824,N_11769);
nor U12257 (N_12257,N_11957,N_11565);
and U12258 (N_12258,N_11773,N_11769);
or U12259 (N_12259,N_11926,N_11815);
or U12260 (N_12260,N_11577,N_11598);
xor U12261 (N_12261,N_11523,N_11933);
nor U12262 (N_12262,N_11574,N_11713);
and U12263 (N_12263,N_11743,N_11914);
or U12264 (N_12264,N_11684,N_11604);
and U12265 (N_12265,N_11793,N_11940);
nor U12266 (N_12266,N_11613,N_11912);
and U12267 (N_12267,N_11616,N_11857);
or U12268 (N_12268,N_11748,N_11743);
nand U12269 (N_12269,N_11698,N_11503);
nor U12270 (N_12270,N_11925,N_11939);
xor U12271 (N_12271,N_11791,N_11825);
xor U12272 (N_12272,N_11601,N_11678);
nor U12273 (N_12273,N_11743,N_11955);
or U12274 (N_12274,N_11675,N_11609);
or U12275 (N_12275,N_11869,N_11831);
xor U12276 (N_12276,N_11688,N_11862);
or U12277 (N_12277,N_11642,N_11602);
or U12278 (N_12278,N_11541,N_11589);
and U12279 (N_12279,N_11550,N_11618);
xnor U12280 (N_12280,N_11534,N_11966);
nor U12281 (N_12281,N_11925,N_11587);
xor U12282 (N_12282,N_11615,N_11512);
nor U12283 (N_12283,N_11507,N_11644);
or U12284 (N_12284,N_11534,N_11817);
nor U12285 (N_12285,N_11629,N_11798);
and U12286 (N_12286,N_11508,N_11835);
nor U12287 (N_12287,N_11753,N_11547);
nand U12288 (N_12288,N_11796,N_11589);
nand U12289 (N_12289,N_11794,N_11788);
nand U12290 (N_12290,N_11670,N_11721);
and U12291 (N_12291,N_11946,N_11799);
or U12292 (N_12292,N_11641,N_11599);
nand U12293 (N_12293,N_11886,N_11933);
or U12294 (N_12294,N_11833,N_11501);
nor U12295 (N_12295,N_11879,N_11618);
and U12296 (N_12296,N_11686,N_11942);
nor U12297 (N_12297,N_11587,N_11576);
nor U12298 (N_12298,N_11585,N_11614);
nor U12299 (N_12299,N_11684,N_11959);
or U12300 (N_12300,N_11909,N_11599);
nand U12301 (N_12301,N_11617,N_11885);
and U12302 (N_12302,N_11911,N_11521);
nand U12303 (N_12303,N_11983,N_11602);
or U12304 (N_12304,N_11922,N_11951);
and U12305 (N_12305,N_11574,N_11680);
xor U12306 (N_12306,N_11850,N_11715);
or U12307 (N_12307,N_11903,N_11702);
and U12308 (N_12308,N_11668,N_11537);
nor U12309 (N_12309,N_11513,N_11917);
and U12310 (N_12310,N_11668,N_11962);
or U12311 (N_12311,N_11624,N_11607);
nand U12312 (N_12312,N_11874,N_11652);
xnor U12313 (N_12313,N_11862,N_11963);
or U12314 (N_12314,N_11647,N_11509);
nor U12315 (N_12315,N_11787,N_11504);
nor U12316 (N_12316,N_11934,N_11555);
or U12317 (N_12317,N_11824,N_11896);
or U12318 (N_12318,N_11641,N_11582);
and U12319 (N_12319,N_11692,N_11731);
and U12320 (N_12320,N_11637,N_11792);
xnor U12321 (N_12321,N_11660,N_11783);
xnor U12322 (N_12322,N_11915,N_11685);
nand U12323 (N_12323,N_11732,N_11582);
xnor U12324 (N_12324,N_11850,N_11735);
and U12325 (N_12325,N_11687,N_11653);
nor U12326 (N_12326,N_11744,N_11549);
xor U12327 (N_12327,N_11547,N_11917);
nand U12328 (N_12328,N_11607,N_11617);
nor U12329 (N_12329,N_11816,N_11946);
and U12330 (N_12330,N_11537,N_11704);
nand U12331 (N_12331,N_11741,N_11753);
nor U12332 (N_12332,N_11646,N_11930);
nor U12333 (N_12333,N_11614,N_11533);
xor U12334 (N_12334,N_11864,N_11675);
and U12335 (N_12335,N_11687,N_11680);
nand U12336 (N_12336,N_11839,N_11965);
nand U12337 (N_12337,N_11748,N_11506);
nor U12338 (N_12338,N_11661,N_11908);
nor U12339 (N_12339,N_11573,N_11966);
or U12340 (N_12340,N_11884,N_11586);
nand U12341 (N_12341,N_11801,N_11620);
and U12342 (N_12342,N_11976,N_11733);
or U12343 (N_12343,N_11899,N_11972);
nand U12344 (N_12344,N_11886,N_11972);
nor U12345 (N_12345,N_11677,N_11577);
or U12346 (N_12346,N_11916,N_11613);
xor U12347 (N_12347,N_11862,N_11503);
nor U12348 (N_12348,N_11898,N_11751);
nand U12349 (N_12349,N_11710,N_11733);
nand U12350 (N_12350,N_11542,N_11518);
xor U12351 (N_12351,N_11861,N_11841);
or U12352 (N_12352,N_11793,N_11930);
nor U12353 (N_12353,N_11669,N_11678);
and U12354 (N_12354,N_11758,N_11689);
nand U12355 (N_12355,N_11934,N_11961);
xor U12356 (N_12356,N_11978,N_11620);
or U12357 (N_12357,N_11886,N_11600);
or U12358 (N_12358,N_11530,N_11637);
nor U12359 (N_12359,N_11975,N_11744);
and U12360 (N_12360,N_11855,N_11572);
nand U12361 (N_12361,N_11649,N_11653);
nand U12362 (N_12362,N_11731,N_11871);
or U12363 (N_12363,N_11677,N_11685);
and U12364 (N_12364,N_11875,N_11770);
xnor U12365 (N_12365,N_11501,N_11887);
xor U12366 (N_12366,N_11589,N_11539);
and U12367 (N_12367,N_11792,N_11910);
or U12368 (N_12368,N_11507,N_11896);
and U12369 (N_12369,N_11604,N_11881);
xor U12370 (N_12370,N_11911,N_11941);
or U12371 (N_12371,N_11779,N_11946);
nand U12372 (N_12372,N_11853,N_11942);
xnor U12373 (N_12373,N_11730,N_11846);
nor U12374 (N_12374,N_11655,N_11823);
nand U12375 (N_12375,N_11704,N_11553);
and U12376 (N_12376,N_11562,N_11729);
nand U12377 (N_12377,N_11973,N_11585);
or U12378 (N_12378,N_11604,N_11836);
nand U12379 (N_12379,N_11533,N_11766);
nand U12380 (N_12380,N_11885,N_11534);
xor U12381 (N_12381,N_11808,N_11659);
and U12382 (N_12382,N_11860,N_11635);
nand U12383 (N_12383,N_11526,N_11556);
nor U12384 (N_12384,N_11670,N_11635);
and U12385 (N_12385,N_11789,N_11714);
nand U12386 (N_12386,N_11578,N_11677);
nand U12387 (N_12387,N_11681,N_11805);
or U12388 (N_12388,N_11534,N_11608);
nor U12389 (N_12389,N_11791,N_11809);
and U12390 (N_12390,N_11737,N_11569);
or U12391 (N_12391,N_11500,N_11985);
xnor U12392 (N_12392,N_11904,N_11650);
or U12393 (N_12393,N_11805,N_11787);
and U12394 (N_12394,N_11629,N_11815);
nor U12395 (N_12395,N_11548,N_11662);
nor U12396 (N_12396,N_11733,N_11944);
and U12397 (N_12397,N_11993,N_11703);
nand U12398 (N_12398,N_11772,N_11996);
and U12399 (N_12399,N_11817,N_11582);
or U12400 (N_12400,N_11768,N_11626);
nand U12401 (N_12401,N_11793,N_11988);
xnor U12402 (N_12402,N_11782,N_11636);
or U12403 (N_12403,N_11888,N_11545);
or U12404 (N_12404,N_11935,N_11809);
xor U12405 (N_12405,N_11860,N_11684);
xnor U12406 (N_12406,N_11898,N_11845);
or U12407 (N_12407,N_11796,N_11574);
or U12408 (N_12408,N_11713,N_11981);
nor U12409 (N_12409,N_11641,N_11734);
nor U12410 (N_12410,N_11655,N_11544);
or U12411 (N_12411,N_11760,N_11917);
nand U12412 (N_12412,N_11989,N_11689);
nand U12413 (N_12413,N_11732,N_11907);
or U12414 (N_12414,N_11645,N_11930);
nand U12415 (N_12415,N_11963,N_11951);
and U12416 (N_12416,N_11989,N_11935);
or U12417 (N_12417,N_11580,N_11569);
nor U12418 (N_12418,N_11643,N_11726);
and U12419 (N_12419,N_11906,N_11749);
nand U12420 (N_12420,N_11674,N_11538);
nor U12421 (N_12421,N_11757,N_11838);
nor U12422 (N_12422,N_11996,N_11500);
and U12423 (N_12423,N_11678,N_11942);
or U12424 (N_12424,N_11942,N_11869);
xor U12425 (N_12425,N_11644,N_11869);
nand U12426 (N_12426,N_11514,N_11894);
and U12427 (N_12427,N_11555,N_11916);
nand U12428 (N_12428,N_11711,N_11986);
and U12429 (N_12429,N_11962,N_11946);
or U12430 (N_12430,N_11909,N_11810);
xor U12431 (N_12431,N_11912,N_11943);
and U12432 (N_12432,N_11711,N_11626);
and U12433 (N_12433,N_11728,N_11653);
xnor U12434 (N_12434,N_11641,N_11538);
or U12435 (N_12435,N_11735,N_11789);
nor U12436 (N_12436,N_11802,N_11733);
and U12437 (N_12437,N_11995,N_11559);
and U12438 (N_12438,N_11726,N_11601);
nor U12439 (N_12439,N_11512,N_11532);
and U12440 (N_12440,N_11675,N_11634);
nand U12441 (N_12441,N_11673,N_11749);
nor U12442 (N_12442,N_11609,N_11625);
and U12443 (N_12443,N_11772,N_11624);
nor U12444 (N_12444,N_11603,N_11879);
nand U12445 (N_12445,N_11706,N_11928);
and U12446 (N_12446,N_11737,N_11686);
and U12447 (N_12447,N_11717,N_11591);
nand U12448 (N_12448,N_11521,N_11601);
xor U12449 (N_12449,N_11721,N_11641);
nand U12450 (N_12450,N_11567,N_11987);
nand U12451 (N_12451,N_11785,N_11945);
and U12452 (N_12452,N_11711,N_11663);
or U12453 (N_12453,N_11788,N_11504);
and U12454 (N_12454,N_11799,N_11890);
xor U12455 (N_12455,N_11645,N_11655);
nor U12456 (N_12456,N_11530,N_11535);
xnor U12457 (N_12457,N_11841,N_11815);
and U12458 (N_12458,N_11987,N_11907);
nand U12459 (N_12459,N_11778,N_11755);
nand U12460 (N_12460,N_11674,N_11581);
and U12461 (N_12461,N_11803,N_11642);
and U12462 (N_12462,N_11731,N_11701);
or U12463 (N_12463,N_11957,N_11558);
xor U12464 (N_12464,N_11626,N_11853);
and U12465 (N_12465,N_11734,N_11544);
nand U12466 (N_12466,N_11987,N_11746);
or U12467 (N_12467,N_11590,N_11540);
nand U12468 (N_12468,N_11569,N_11856);
nor U12469 (N_12469,N_11651,N_11970);
xnor U12470 (N_12470,N_11912,N_11753);
nor U12471 (N_12471,N_11891,N_11993);
or U12472 (N_12472,N_11962,N_11923);
nand U12473 (N_12473,N_11792,N_11882);
nor U12474 (N_12474,N_11673,N_11742);
nand U12475 (N_12475,N_11940,N_11874);
xor U12476 (N_12476,N_11601,N_11967);
and U12477 (N_12477,N_11743,N_11949);
nand U12478 (N_12478,N_11792,N_11900);
or U12479 (N_12479,N_11997,N_11705);
or U12480 (N_12480,N_11721,N_11820);
and U12481 (N_12481,N_11740,N_11915);
nor U12482 (N_12482,N_11852,N_11981);
xnor U12483 (N_12483,N_11607,N_11864);
or U12484 (N_12484,N_11661,N_11727);
and U12485 (N_12485,N_11738,N_11893);
and U12486 (N_12486,N_11509,N_11892);
nor U12487 (N_12487,N_11890,N_11931);
nor U12488 (N_12488,N_11663,N_11681);
nand U12489 (N_12489,N_11517,N_11985);
nor U12490 (N_12490,N_11790,N_11841);
or U12491 (N_12491,N_11630,N_11578);
or U12492 (N_12492,N_11877,N_11626);
or U12493 (N_12493,N_11752,N_11832);
and U12494 (N_12494,N_11748,N_11887);
and U12495 (N_12495,N_11787,N_11722);
or U12496 (N_12496,N_11694,N_11939);
nand U12497 (N_12497,N_11524,N_11620);
and U12498 (N_12498,N_11907,N_11766);
nor U12499 (N_12499,N_11838,N_11860);
and U12500 (N_12500,N_12262,N_12158);
nor U12501 (N_12501,N_12497,N_12277);
or U12502 (N_12502,N_12398,N_12041);
or U12503 (N_12503,N_12233,N_12055);
nand U12504 (N_12504,N_12216,N_12498);
or U12505 (N_12505,N_12074,N_12480);
nand U12506 (N_12506,N_12176,N_12283);
xnor U12507 (N_12507,N_12380,N_12438);
and U12508 (N_12508,N_12125,N_12095);
nor U12509 (N_12509,N_12457,N_12200);
nand U12510 (N_12510,N_12444,N_12291);
or U12511 (N_12511,N_12173,N_12435);
nand U12512 (N_12512,N_12440,N_12460);
nor U12513 (N_12513,N_12169,N_12311);
and U12514 (N_12514,N_12486,N_12228);
xnor U12515 (N_12515,N_12028,N_12107);
or U12516 (N_12516,N_12007,N_12054);
or U12517 (N_12517,N_12255,N_12036);
xnor U12518 (N_12518,N_12297,N_12415);
or U12519 (N_12519,N_12265,N_12001);
and U12520 (N_12520,N_12210,N_12131);
or U12521 (N_12521,N_12057,N_12263);
nand U12522 (N_12522,N_12012,N_12000);
nor U12523 (N_12523,N_12379,N_12324);
nor U12524 (N_12524,N_12052,N_12247);
and U12525 (N_12525,N_12383,N_12185);
and U12526 (N_12526,N_12439,N_12328);
nand U12527 (N_12527,N_12226,N_12071);
nand U12528 (N_12528,N_12410,N_12455);
nor U12529 (N_12529,N_12326,N_12269);
nor U12530 (N_12530,N_12432,N_12144);
or U12531 (N_12531,N_12085,N_12449);
or U12532 (N_12532,N_12307,N_12402);
nor U12533 (N_12533,N_12215,N_12385);
xor U12534 (N_12534,N_12197,N_12374);
nor U12535 (N_12535,N_12043,N_12303);
nor U12536 (N_12536,N_12251,N_12335);
nor U12537 (N_12537,N_12142,N_12353);
or U12538 (N_12538,N_12014,N_12302);
nand U12539 (N_12539,N_12021,N_12378);
xnor U12540 (N_12540,N_12189,N_12414);
nand U12541 (N_12541,N_12063,N_12155);
and U12542 (N_12542,N_12248,N_12177);
and U12543 (N_12543,N_12266,N_12088);
xnor U12544 (N_12544,N_12395,N_12096);
or U12545 (N_12545,N_12179,N_12275);
xnor U12546 (N_12546,N_12428,N_12267);
nand U12547 (N_12547,N_12163,N_12033);
and U12548 (N_12548,N_12219,N_12495);
nor U12549 (N_12549,N_12093,N_12221);
or U12550 (N_12550,N_12412,N_12124);
nand U12551 (N_12551,N_12035,N_12005);
or U12552 (N_12552,N_12331,N_12134);
xor U12553 (N_12553,N_12238,N_12422);
nand U12554 (N_12554,N_12253,N_12334);
nand U12555 (N_12555,N_12019,N_12048);
or U12556 (N_12556,N_12489,N_12069);
xor U12557 (N_12557,N_12076,N_12116);
or U12558 (N_12558,N_12049,N_12109);
or U12559 (N_12559,N_12212,N_12211);
or U12560 (N_12560,N_12154,N_12401);
nor U12561 (N_12561,N_12184,N_12137);
nand U12562 (N_12562,N_12191,N_12301);
nand U12563 (N_12563,N_12332,N_12222);
and U12564 (N_12564,N_12492,N_12360);
and U12565 (N_12565,N_12080,N_12314);
nor U12566 (N_12566,N_12425,N_12465);
or U12567 (N_12567,N_12104,N_12446);
and U12568 (N_12568,N_12464,N_12084);
and U12569 (N_12569,N_12366,N_12135);
and U12570 (N_12570,N_12299,N_12220);
and U12571 (N_12571,N_12298,N_12241);
or U12572 (N_12572,N_12406,N_12394);
nand U12573 (N_12573,N_12227,N_12034);
nand U12574 (N_12574,N_12454,N_12140);
nand U12575 (N_12575,N_12249,N_12382);
xnor U12576 (N_12576,N_12310,N_12290);
or U12577 (N_12577,N_12192,N_12451);
and U12578 (N_12578,N_12106,N_12389);
nor U12579 (N_12579,N_12499,N_12458);
xnor U12580 (N_12580,N_12305,N_12214);
and U12581 (N_12581,N_12348,N_12162);
or U12582 (N_12582,N_12289,N_12487);
nor U12583 (N_12583,N_12045,N_12256);
nand U12584 (N_12584,N_12208,N_12170);
or U12585 (N_12585,N_12025,N_12408);
nand U12586 (N_12586,N_12183,N_12120);
or U12587 (N_12587,N_12419,N_12463);
nor U12588 (N_12588,N_12224,N_12016);
nand U12589 (N_12589,N_12268,N_12296);
and U12590 (N_12590,N_12032,N_12278);
nand U12591 (N_12591,N_12285,N_12145);
and U12592 (N_12592,N_12481,N_12362);
nand U12593 (N_12593,N_12138,N_12011);
nand U12594 (N_12594,N_12100,N_12445);
nand U12595 (N_12595,N_12427,N_12400);
nand U12596 (N_12596,N_12391,N_12168);
nand U12597 (N_12597,N_12437,N_12058);
or U12598 (N_12598,N_12089,N_12318);
nor U12599 (N_12599,N_12196,N_12064);
xor U12600 (N_12600,N_12044,N_12230);
or U12601 (N_12601,N_12418,N_12203);
nand U12602 (N_12602,N_12008,N_12456);
xnor U12603 (N_12603,N_12347,N_12376);
nand U12604 (N_12604,N_12274,N_12209);
nand U12605 (N_12605,N_12494,N_12309);
nor U12606 (N_12606,N_12354,N_12264);
xor U12607 (N_12607,N_12060,N_12308);
nor U12608 (N_12608,N_12204,N_12083);
nand U12609 (N_12609,N_12413,N_12094);
xor U12610 (N_12610,N_12159,N_12370);
or U12611 (N_12611,N_12235,N_12341);
nor U12612 (N_12612,N_12340,N_12294);
nor U12613 (N_12613,N_12450,N_12143);
nand U12614 (N_12614,N_12260,N_12424);
or U12615 (N_12615,N_12153,N_12244);
or U12616 (N_12616,N_12423,N_12270);
and U12617 (N_12617,N_12363,N_12037);
nor U12618 (N_12618,N_12018,N_12122);
or U12619 (N_12619,N_12146,N_12167);
or U12620 (N_12620,N_12442,N_12101);
nand U12621 (N_12621,N_12113,N_12186);
nor U12622 (N_12622,N_12488,N_12316);
nand U12623 (N_12623,N_12062,N_12344);
nand U12624 (N_12624,N_12243,N_12375);
nor U12625 (N_12625,N_12053,N_12188);
nor U12626 (N_12626,N_12276,N_12342);
nand U12627 (N_12627,N_12404,N_12031);
nand U12628 (N_12628,N_12322,N_12436);
nand U12629 (N_12629,N_12369,N_12286);
nor U12630 (N_12630,N_12453,N_12119);
nor U12631 (N_12631,N_12421,N_12156);
nor U12632 (N_12632,N_12115,N_12381);
and U12633 (N_12633,N_12284,N_12172);
nor U12634 (N_12634,N_12242,N_12467);
xnor U12635 (N_12635,N_12462,N_12079);
or U12636 (N_12636,N_12472,N_12367);
nand U12637 (N_12637,N_12246,N_12190);
and U12638 (N_12638,N_12046,N_12013);
xor U12639 (N_12639,N_12337,N_12430);
nand U12640 (N_12640,N_12252,N_12357);
nand U12641 (N_12641,N_12490,N_12194);
nand U12642 (N_12642,N_12452,N_12112);
xnor U12643 (N_12643,N_12443,N_12448);
or U12644 (N_12644,N_12232,N_12090);
nor U12645 (N_12645,N_12359,N_12160);
or U12646 (N_12646,N_12346,N_12384);
nor U12647 (N_12647,N_12121,N_12420);
nor U12648 (N_12648,N_12466,N_12047);
nand U12649 (N_12649,N_12461,N_12387);
nand U12650 (N_12650,N_12441,N_12250);
nand U12651 (N_12651,N_12361,N_12349);
and U12652 (N_12652,N_12358,N_12050);
xnor U12653 (N_12653,N_12181,N_12373);
and U12654 (N_12654,N_12234,N_12202);
and U12655 (N_12655,N_12006,N_12459);
or U12656 (N_12656,N_12206,N_12087);
nor U12657 (N_12657,N_12127,N_12468);
nor U12658 (N_12658,N_12149,N_12067);
nor U12659 (N_12659,N_12287,N_12312);
or U12660 (N_12660,N_12010,N_12485);
and U12661 (N_12661,N_12097,N_12081);
nand U12662 (N_12662,N_12434,N_12431);
nor U12663 (N_12663,N_12026,N_12282);
or U12664 (N_12664,N_12004,N_12279);
xnor U12665 (N_12665,N_12426,N_12039);
xnor U12666 (N_12666,N_12447,N_12023);
and U12667 (N_12667,N_12139,N_12352);
xnor U12668 (N_12668,N_12470,N_12065);
and U12669 (N_12669,N_12273,N_12392);
xor U12670 (N_12670,N_12272,N_12330);
and U12671 (N_12671,N_12180,N_12174);
and U12672 (N_12672,N_12141,N_12491);
nand U12673 (N_12673,N_12479,N_12105);
nand U12674 (N_12674,N_12483,N_12218);
and U12675 (N_12675,N_12077,N_12295);
nor U12676 (N_12676,N_12317,N_12136);
nor U12677 (N_12677,N_12020,N_12029);
and U12678 (N_12678,N_12148,N_12355);
or U12679 (N_12679,N_12325,N_12030);
nand U12680 (N_12680,N_12066,N_12075);
nand U12681 (N_12681,N_12372,N_12365);
nand U12682 (N_12682,N_12198,N_12416);
nand U12683 (N_12683,N_12403,N_12386);
nor U12684 (N_12684,N_12207,N_12166);
nor U12685 (N_12685,N_12390,N_12175);
or U12686 (N_12686,N_12300,N_12072);
or U12687 (N_12687,N_12205,N_12042);
nand U12688 (N_12688,N_12061,N_12009);
nand U12689 (N_12689,N_12223,N_12130);
and U12690 (N_12690,N_12245,N_12399);
or U12691 (N_12691,N_12471,N_12429);
nor U12692 (N_12692,N_12102,N_12108);
nand U12693 (N_12693,N_12474,N_12091);
nor U12694 (N_12694,N_12165,N_12147);
or U12695 (N_12695,N_12329,N_12350);
or U12696 (N_12696,N_12133,N_12099);
nor U12697 (N_12697,N_12339,N_12114);
nand U12698 (N_12698,N_12128,N_12237);
xor U12699 (N_12699,N_12469,N_12259);
or U12700 (N_12700,N_12288,N_12129);
nand U12701 (N_12701,N_12195,N_12068);
or U12702 (N_12702,N_12051,N_12356);
and U12703 (N_12703,N_12003,N_12323);
nand U12704 (N_12704,N_12118,N_12123);
nor U12705 (N_12705,N_12017,N_12473);
nor U12706 (N_12706,N_12336,N_12152);
nor U12707 (N_12707,N_12271,N_12229);
and U12708 (N_12708,N_12280,N_12338);
or U12709 (N_12709,N_12171,N_12092);
xnor U12710 (N_12710,N_12261,N_12405);
nor U12711 (N_12711,N_12407,N_12476);
or U12712 (N_12712,N_12225,N_12126);
nor U12713 (N_12713,N_12477,N_12371);
nand U12714 (N_12714,N_12110,N_12027);
and U12715 (N_12715,N_12151,N_12213);
nand U12716 (N_12716,N_12493,N_12484);
or U12717 (N_12717,N_12368,N_12231);
nor U12718 (N_12718,N_12002,N_12056);
and U12719 (N_12719,N_12478,N_12161);
and U12720 (N_12720,N_12078,N_12150);
nor U12721 (N_12721,N_12364,N_12239);
nand U12722 (N_12722,N_12433,N_12345);
or U12723 (N_12723,N_12073,N_12022);
or U12724 (N_12724,N_12038,N_12321);
and U12725 (N_12725,N_12351,N_12397);
or U12726 (N_12726,N_12396,N_12315);
nor U12727 (N_12727,N_12327,N_12236);
nor U12728 (N_12728,N_12409,N_12199);
nor U12729 (N_12729,N_12178,N_12319);
nand U12730 (N_12730,N_12187,N_12496);
and U12731 (N_12731,N_12193,N_12254);
and U12732 (N_12732,N_12292,N_12164);
nand U12733 (N_12733,N_12024,N_12306);
nand U12734 (N_12734,N_12098,N_12070);
and U12735 (N_12735,N_12015,N_12182);
and U12736 (N_12736,N_12393,N_12304);
or U12737 (N_12737,N_12293,N_12320);
and U12738 (N_12738,N_12217,N_12117);
and U12739 (N_12739,N_12201,N_12240);
and U12740 (N_12740,N_12411,N_12281);
nor U12741 (N_12741,N_12111,N_12059);
and U12742 (N_12742,N_12132,N_12333);
and U12743 (N_12743,N_12103,N_12343);
nand U12744 (N_12744,N_12040,N_12475);
and U12745 (N_12745,N_12417,N_12257);
or U12746 (N_12746,N_12482,N_12377);
or U12747 (N_12747,N_12313,N_12157);
nor U12748 (N_12748,N_12258,N_12082);
nand U12749 (N_12749,N_12086,N_12388);
and U12750 (N_12750,N_12394,N_12179);
and U12751 (N_12751,N_12381,N_12103);
xnor U12752 (N_12752,N_12332,N_12364);
and U12753 (N_12753,N_12485,N_12075);
and U12754 (N_12754,N_12492,N_12472);
and U12755 (N_12755,N_12040,N_12059);
nor U12756 (N_12756,N_12426,N_12229);
and U12757 (N_12757,N_12237,N_12475);
nand U12758 (N_12758,N_12335,N_12312);
or U12759 (N_12759,N_12002,N_12255);
xor U12760 (N_12760,N_12106,N_12009);
nor U12761 (N_12761,N_12259,N_12497);
nand U12762 (N_12762,N_12238,N_12201);
nand U12763 (N_12763,N_12121,N_12475);
nand U12764 (N_12764,N_12036,N_12097);
nor U12765 (N_12765,N_12274,N_12161);
or U12766 (N_12766,N_12267,N_12473);
and U12767 (N_12767,N_12353,N_12335);
nor U12768 (N_12768,N_12357,N_12194);
nor U12769 (N_12769,N_12362,N_12400);
xnor U12770 (N_12770,N_12336,N_12208);
xor U12771 (N_12771,N_12239,N_12053);
and U12772 (N_12772,N_12443,N_12342);
or U12773 (N_12773,N_12168,N_12142);
xor U12774 (N_12774,N_12311,N_12226);
and U12775 (N_12775,N_12332,N_12453);
or U12776 (N_12776,N_12090,N_12129);
nand U12777 (N_12777,N_12239,N_12159);
and U12778 (N_12778,N_12454,N_12414);
or U12779 (N_12779,N_12352,N_12421);
and U12780 (N_12780,N_12238,N_12491);
nor U12781 (N_12781,N_12487,N_12304);
nand U12782 (N_12782,N_12438,N_12463);
or U12783 (N_12783,N_12478,N_12065);
and U12784 (N_12784,N_12083,N_12397);
nor U12785 (N_12785,N_12267,N_12471);
xnor U12786 (N_12786,N_12106,N_12171);
or U12787 (N_12787,N_12012,N_12491);
and U12788 (N_12788,N_12044,N_12299);
or U12789 (N_12789,N_12280,N_12403);
and U12790 (N_12790,N_12085,N_12428);
or U12791 (N_12791,N_12266,N_12126);
nand U12792 (N_12792,N_12157,N_12455);
nand U12793 (N_12793,N_12010,N_12365);
nor U12794 (N_12794,N_12129,N_12482);
and U12795 (N_12795,N_12007,N_12408);
or U12796 (N_12796,N_12254,N_12379);
or U12797 (N_12797,N_12167,N_12112);
and U12798 (N_12798,N_12420,N_12370);
nor U12799 (N_12799,N_12319,N_12338);
nor U12800 (N_12800,N_12395,N_12360);
nor U12801 (N_12801,N_12369,N_12299);
nor U12802 (N_12802,N_12470,N_12015);
or U12803 (N_12803,N_12299,N_12193);
and U12804 (N_12804,N_12309,N_12252);
or U12805 (N_12805,N_12279,N_12011);
nand U12806 (N_12806,N_12276,N_12399);
nor U12807 (N_12807,N_12058,N_12085);
nand U12808 (N_12808,N_12185,N_12054);
or U12809 (N_12809,N_12428,N_12042);
nand U12810 (N_12810,N_12334,N_12188);
nand U12811 (N_12811,N_12356,N_12162);
nor U12812 (N_12812,N_12481,N_12325);
nor U12813 (N_12813,N_12054,N_12407);
nand U12814 (N_12814,N_12471,N_12109);
or U12815 (N_12815,N_12317,N_12051);
xor U12816 (N_12816,N_12437,N_12007);
nand U12817 (N_12817,N_12351,N_12418);
nor U12818 (N_12818,N_12276,N_12112);
xor U12819 (N_12819,N_12018,N_12356);
or U12820 (N_12820,N_12411,N_12065);
nand U12821 (N_12821,N_12365,N_12458);
nor U12822 (N_12822,N_12244,N_12197);
and U12823 (N_12823,N_12274,N_12160);
nand U12824 (N_12824,N_12248,N_12067);
and U12825 (N_12825,N_12206,N_12310);
xnor U12826 (N_12826,N_12261,N_12008);
nor U12827 (N_12827,N_12044,N_12043);
nor U12828 (N_12828,N_12213,N_12129);
nor U12829 (N_12829,N_12473,N_12174);
nor U12830 (N_12830,N_12029,N_12167);
or U12831 (N_12831,N_12017,N_12499);
and U12832 (N_12832,N_12431,N_12265);
and U12833 (N_12833,N_12221,N_12448);
and U12834 (N_12834,N_12314,N_12480);
nand U12835 (N_12835,N_12257,N_12078);
or U12836 (N_12836,N_12180,N_12050);
or U12837 (N_12837,N_12024,N_12257);
nand U12838 (N_12838,N_12272,N_12207);
nor U12839 (N_12839,N_12217,N_12236);
and U12840 (N_12840,N_12311,N_12497);
and U12841 (N_12841,N_12429,N_12030);
and U12842 (N_12842,N_12133,N_12420);
nor U12843 (N_12843,N_12185,N_12317);
and U12844 (N_12844,N_12218,N_12242);
or U12845 (N_12845,N_12146,N_12244);
and U12846 (N_12846,N_12475,N_12186);
nor U12847 (N_12847,N_12194,N_12270);
nand U12848 (N_12848,N_12307,N_12253);
or U12849 (N_12849,N_12183,N_12298);
or U12850 (N_12850,N_12190,N_12285);
or U12851 (N_12851,N_12466,N_12050);
and U12852 (N_12852,N_12019,N_12261);
nand U12853 (N_12853,N_12450,N_12367);
or U12854 (N_12854,N_12372,N_12028);
and U12855 (N_12855,N_12401,N_12453);
nor U12856 (N_12856,N_12483,N_12055);
or U12857 (N_12857,N_12420,N_12407);
and U12858 (N_12858,N_12006,N_12122);
nand U12859 (N_12859,N_12401,N_12462);
or U12860 (N_12860,N_12220,N_12182);
nand U12861 (N_12861,N_12228,N_12276);
nand U12862 (N_12862,N_12010,N_12484);
nor U12863 (N_12863,N_12387,N_12225);
and U12864 (N_12864,N_12328,N_12423);
nor U12865 (N_12865,N_12423,N_12478);
nand U12866 (N_12866,N_12223,N_12099);
or U12867 (N_12867,N_12397,N_12099);
nand U12868 (N_12868,N_12226,N_12446);
or U12869 (N_12869,N_12482,N_12020);
or U12870 (N_12870,N_12002,N_12380);
and U12871 (N_12871,N_12333,N_12449);
and U12872 (N_12872,N_12485,N_12288);
or U12873 (N_12873,N_12051,N_12335);
or U12874 (N_12874,N_12278,N_12274);
or U12875 (N_12875,N_12494,N_12132);
or U12876 (N_12876,N_12432,N_12421);
and U12877 (N_12877,N_12243,N_12164);
nand U12878 (N_12878,N_12175,N_12176);
and U12879 (N_12879,N_12424,N_12410);
or U12880 (N_12880,N_12050,N_12028);
and U12881 (N_12881,N_12364,N_12022);
nor U12882 (N_12882,N_12186,N_12135);
or U12883 (N_12883,N_12205,N_12465);
and U12884 (N_12884,N_12459,N_12339);
and U12885 (N_12885,N_12478,N_12032);
xnor U12886 (N_12886,N_12011,N_12048);
or U12887 (N_12887,N_12459,N_12353);
or U12888 (N_12888,N_12113,N_12297);
and U12889 (N_12889,N_12443,N_12412);
or U12890 (N_12890,N_12235,N_12453);
nand U12891 (N_12891,N_12111,N_12276);
and U12892 (N_12892,N_12237,N_12025);
nand U12893 (N_12893,N_12010,N_12295);
and U12894 (N_12894,N_12323,N_12289);
nor U12895 (N_12895,N_12434,N_12122);
and U12896 (N_12896,N_12164,N_12422);
nor U12897 (N_12897,N_12076,N_12264);
nand U12898 (N_12898,N_12041,N_12361);
or U12899 (N_12899,N_12098,N_12416);
or U12900 (N_12900,N_12444,N_12189);
nand U12901 (N_12901,N_12109,N_12015);
xnor U12902 (N_12902,N_12356,N_12344);
nand U12903 (N_12903,N_12407,N_12278);
or U12904 (N_12904,N_12328,N_12283);
nor U12905 (N_12905,N_12033,N_12323);
or U12906 (N_12906,N_12226,N_12356);
nand U12907 (N_12907,N_12290,N_12325);
nor U12908 (N_12908,N_12185,N_12034);
and U12909 (N_12909,N_12395,N_12020);
nor U12910 (N_12910,N_12465,N_12345);
nor U12911 (N_12911,N_12379,N_12042);
nand U12912 (N_12912,N_12324,N_12258);
nor U12913 (N_12913,N_12124,N_12020);
nand U12914 (N_12914,N_12074,N_12383);
and U12915 (N_12915,N_12285,N_12106);
and U12916 (N_12916,N_12460,N_12008);
nor U12917 (N_12917,N_12161,N_12069);
nand U12918 (N_12918,N_12209,N_12375);
nand U12919 (N_12919,N_12287,N_12248);
and U12920 (N_12920,N_12072,N_12134);
nand U12921 (N_12921,N_12290,N_12335);
nor U12922 (N_12922,N_12077,N_12142);
nand U12923 (N_12923,N_12421,N_12495);
and U12924 (N_12924,N_12205,N_12426);
nor U12925 (N_12925,N_12101,N_12407);
nor U12926 (N_12926,N_12198,N_12112);
or U12927 (N_12927,N_12354,N_12127);
nand U12928 (N_12928,N_12016,N_12078);
nor U12929 (N_12929,N_12170,N_12381);
nand U12930 (N_12930,N_12076,N_12083);
nand U12931 (N_12931,N_12246,N_12282);
nand U12932 (N_12932,N_12448,N_12242);
and U12933 (N_12933,N_12363,N_12337);
nor U12934 (N_12934,N_12201,N_12458);
or U12935 (N_12935,N_12387,N_12175);
nor U12936 (N_12936,N_12030,N_12057);
nor U12937 (N_12937,N_12382,N_12187);
nor U12938 (N_12938,N_12181,N_12286);
nor U12939 (N_12939,N_12367,N_12257);
xor U12940 (N_12940,N_12259,N_12326);
xor U12941 (N_12941,N_12137,N_12289);
and U12942 (N_12942,N_12052,N_12313);
nand U12943 (N_12943,N_12100,N_12391);
and U12944 (N_12944,N_12174,N_12455);
and U12945 (N_12945,N_12043,N_12056);
and U12946 (N_12946,N_12179,N_12429);
nand U12947 (N_12947,N_12465,N_12207);
or U12948 (N_12948,N_12137,N_12096);
nor U12949 (N_12949,N_12070,N_12240);
or U12950 (N_12950,N_12436,N_12121);
nor U12951 (N_12951,N_12415,N_12024);
or U12952 (N_12952,N_12073,N_12216);
and U12953 (N_12953,N_12309,N_12358);
xor U12954 (N_12954,N_12422,N_12432);
and U12955 (N_12955,N_12119,N_12110);
nand U12956 (N_12956,N_12275,N_12080);
nor U12957 (N_12957,N_12400,N_12045);
or U12958 (N_12958,N_12355,N_12070);
nor U12959 (N_12959,N_12013,N_12370);
or U12960 (N_12960,N_12249,N_12123);
and U12961 (N_12961,N_12497,N_12168);
nand U12962 (N_12962,N_12291,N_12288);
nand U12963 (N_12963,N_12236,N_12456);
nand U12964 (N_12964,N_12306,N_12369);
or U12965 (N_12965,N_12114,N_12447);
nor U12966 (N_12966,N_12046,N_12273);
or U12967 (N_12967,N_12479,N_12352);
and U12968 (N_12968,N_12161,N_12253);
nand U12969 (N_12969,N_12142,N_12135);
and U12970 (N_12970,N_12454,N_12246);
and U12971 (N_12971,N_12102,N_12105);
and U12972 (N_12972,N_12352,N_12237);
nand U12973 (N_12973,N_12313,N_12019);
nor U12974 (N_12974,N_12425,N_12191);
nor U12975 (N_12975,N_12112,N_12034);
xor U12976 (N_12976,N_12041,N_12476);
nand U12977 (N_12977,N_12189,N_12411);
xnor U12978 (N_12978,N_12213,N_12344);
and U12979 (N_12979,N_12329,N_12119);
nor U12980 (N_12980,N_12354,N_12243);
or U12981 (N_12981,N_12470,N_12045);
nor U12982 (N_12982,N_12053,N_12464);
nor U12983 (N_12983,N_12149,N_12177);
nor U12984 (N_12984,N_12186,N_12369);
or U12985 (N_12985,N_12280,N_12358);
or U12986 (N_12986,N_12283,N_12224);
xnor U12987 (N_12987,N_12048,N_12350);
nor U12988 (N_12988,N_12287,N_12054);
nand U12989 (N_12989,N_12265,N_12085);
or U12990 (N_12990,N_12355,N_12146);
xnor U12991 (N_12991,N_12315,N_12349);
and U12992 (N_12992,N_12213,N_12235);
nand U12993 (N_12993,N_12041,N_12459);
nand U12994 (N_12994,N_12119,N_12334);
nand U12995 (N_12995,N_12298,N_12278);
nand U12996 (N_12996,N_12143,N_12130);
xnor U12997 (N_12997,N_12440,N_12398);
xor U12998 (N_12998,N_12021,N_12060);
xor U12999 (N_12999,N_12158,N_12136);
nor U13000 (N_13000,N_12860,N_12934);
nand U13001 (N_13001,N_12718,N_12686);
nand U13002 (N_13002,N_12746,N_12960);
nor U13003 (N_13003,N_12891,N_12771);
nand U13004 (N_13004,N_12975,N_12827);
nand U13005 (N_13005,N_12550,N_12561);
nand U13006 (N_13006,N_12678,N_12831);
nor U13007 (N_13007,N_12578,N_12539);
nor U13008 (N_13008,N_12616,N_12872);
nor U13009 (N_13009,N_12669,N_12576);
or U13010 (N_13010,N_12765,N_12835);
xor U13011 (N_13011,N_12999,N_12711);
nand U13012 (N_13012,N_12613,N_12738);
nand U13013 (N_13013,N_12736,N_12627);
nor U13014 (N_13014,N_12668,N_12573);
and U13015 (N_13015,N_12659,N_12972);
or U13016 (N_13016,N_12956,N_12713);
nor U13017 (N_13017,N_12599,N_12569);
nand U13018 (N_13018,N_12877,N_12581);
nor U13019 (N_13019,N_12864,N_12784);
or U13020 (N_13020,N_12935,N_12532);
and U13021 (N_13021,N_12818,N_12901);
or U13022 (N_13022,N_12774,N_12502);
or U13023 (N_13023,N_12551,N_12634);
nand U13024 (N_13024,N_12694,N_12874);
and U13025 (N_13025,N_12828,N_12854);
and U13026 (N_13026,N_12527,N_12662);
and U13027 (N_13027,N_12665,N_12781);
or U13028 (N_13028,N_12504,N_12846);
and U13029 (N_13029,N_12510,N_12714);
xor U13030 (N_13030,N_12692,N_12633);
and U13031 (N_13031,N_12590,N_12756);
xor U13032 (N_13032,N_12884,N_12571);
nand U13033 (N_13033,N_12897,N_12726);
nand U13034 (N_13034,N_12703,N_12788);
nor U13035 (N_13035,N_12710,N_12879);
nand U13036 (N_13036,N_12509,N_12838);
and U13037 (N_13037,N_12801,N_12516);
nor U13038 (N_13038,N_12688,N_12913);
nand U13039 (N_13039,N_12518,N_12648);
and U13040 (N_13040,N_12947,N_12789);
nand U13041 (N_13041,N_12525,N_12990);
nand U13042 (N_13042,N_12521,N_12607);
xor U13043 (N_13043,N_12836,N_12855);
nor U13044 (N_13044,N_12931,N_12605);
nand U13045 (N_13045,N_12790,N_12664);
and U13046 (N_13046,N_12555,N_12973);
nor U13047 (N_13047,N_12825,N_12820);
or U13048 (N_13048,N_12522,N_12957);
and U13049 (N_13049,N_12780,N_12923);
or U13050 (N_13050,N_12841,N_12566);
and U13051 (N_13051,N_12614,N_12565);
xor U13052 (N_13052,N_12908,N_12536);
xnor U13053 (N_13053,N_12865,N_12862);
nor U13054 (N_13054,N_12554,N_12528);
and U13055 (N_13055,N_12829,N_12951);
or U13056 (N_13056,N_12916,N_12684);
or U13057 (N_13057,N_12524,N_12941);
and U13058 (N_13058,N_12940,N_12873);
and U13059 (N_13059,N_12988,N_12823);
xor U13060 (N_13060,N_12986,N_12851);
nor U13061 (N_13061,N_12671,N_12606);
nor U13062 (N_13062,N_12965,N_12690);
or U13063 (N_13063,N_12587,N_12677);
nand U13064 (N_13064,N_12776,N_12600);
xnor U13065 (N_13065,N_12506,N_12579);
nand U13066 (N_13066,N_12775,N_12933);
and U13067 (N_13067,N_12501,N_12712);
nor U13068 (N_13068,N_12515,N_12593);
and U13069 (N_13069,N_12920,N_12803);
or U13070 (N_13070,N_12870,N_12995);
nor U13071 (N_13071,N_12770,N_12572);
nor U13072 (N_13072,N_12924,N_12954);
and U13073 (N_13073,N_12980,N_12882);
nor U13074 (N_13074,N_12859,N_12927);
nand U13075 (N_13075,N_12592,N_12700);
nand U13076 (N_13076,N_12507,N_12716);
xor U13077 (N_13077,N_12702,N_12612);
and U13078 (N_13078,N_12969,N_12608);
nor U13079 (N_13079,N_12643,N_12763);
nor U13080 (N_13080,N_12869,N_12748);
or U13081 (N_13081,N_12867,N_12837);
and U13082 (N_13082,N_12826,N_12833);
nor U13083 (N_13083,N_12666,N_12529);
nor U13084 (N_13084,N_12556,N_12946);
nor U13085 (N_13085,N_12892,N_12812);
nand U13086 (N_13086,N_12844,N_12583);
nand U13087 (N_13087,N_12996,N_12758);
or U13088 (N_13088,N_12834,N_12798);
or U13089 (N_13089,N_12961,N_12866);
and U13090 (N_13090,N_12697,N_12562);
or U13091 (N_13091,N_12992,N_12548);
and U13092 (N_13092,N_12853,N_12785);
or U13093 (N_13093,N_12753,N_12511);
nor U13094 (N_13094,N_12685,N_12595);
or U13095 (N_13095,N_12845,N_12655);
or U13096 (N_13096,N_12977,N_12989);
and U13097 (N_13097,N_12681,N_12647);
or U13098 (N_13098,N_12883,N_12728);
nand U13099 (N_13099,N_12640,N_12707);
nand U13100 (N_13100,N_12537,N_12840);
or U13101 (N_13101,N_12907,N_12638);
xnor U13102 (N_13102,N_12601,N_12952);
or U13103 (N_13103,N_12672,N_12603);
or U13104 (N_13104,N_12793,N_12783);
and U13105 (N_13105,N_12657,N_12904);
nand U13106 (N_13106,N_12729,N_12886);
and U13107 (N_13107,N_12899,N_12651);
nor U13108 (N_13108,N_12821,N_12708);
and U13109 (N_13109,N_12768,N_12810);
or U13110 (N_13110,N_12804,N_12800);
nor U13111 (N_13111,N_12675,N_12778);
xor U13112 (N_13112,N_12949,N_12856);
or U13113 (N_13113,N_12535,N_12722);
nand U13114 (N_13114,N_12584,N_12863);
xor U13115 (N_13115,N_12609,N_12575);
and U13116 (N_13116,N_12628,N_12549);
nand U13117 (N_13117,N_12880,N_12811);
or U13118 (N_13118,N_12586,N_12689);
or U13119 (N_13119,N_12805,N_12623);
or U13120 (N_13120,N_12531,N_12630);
nand U13121 (N_13121,N_12902,N_12849);
or U13122 (N_13122,N_12629,N_12759);
nand U13123 (N_13123,N_12626,N_12791);
or U13124 (N_13124,N_12797,N_12932);
xor U13125 (N_13125,N_12898,N_12721);
xnor U13126 (N_13126,N_12937,N_12842);
and U13127 (N_13127,N_12558,N_12503);
xnor U13128 (N_13128,N_12964,N_12585);
nor U13129 (N_13129,N_12762,N_12676);
nand U13130 (N_13130,N_12679,N_12912);
or U13131 (N_13131,N_12598,N_12602);
and U13132 (N_13132,N_12682,N_12611);
xnor U13133 (N_13133,N_12559,N_12795);
nand U13134 (N_13134,N_12750,N_12887);
or U13135 (N_13135,N_12896,N_12693);
nand U13136 (N_13136,N_12832,N_12513);
nor U13137 (N_13137,N_12918,N_12589);
nor U13138 (N_13138,N_12786,N_12876);
or U13139 (N_13139,N_12661,N_12691);
and U13140 (N_13140,N_12725,N_12921);
and U13141 (N_13141,N_12588,N_12747);
xor U13142 (N_13142,N_12755,N_12983);
and U13143 (N_13143,N_12993,N_12893);
nor U13144 (N_13144,N_12991,N_12761);
nor U13145 (N_13145,N_12766,N_12740);
or U13146 (N_13146,N_12542,N_12695);
nor U13147 (N_13147,N_12981,N_12610);
nand U13148 (N_13148,N_12654,N_12772);
nand U13149 (N_13149,N_12731,N_12839);
or U13150 (N_13150,N_12928,N_12696);
nand U13151 (N_13151,N_12724,N_12512);
or U13152 (N_13152,N_12520,N_12757);
nand U13153 (N_13153,N_12807,N_12948);
nor U13154 (N_13154,N_12802,N_12631);
xnor U13155 (N_13155,N_12717,N_12936);
xnor U13156 (N_13156,N_12580,N_12822);
or U13157 (N_13157,N_12777,N_12751);
nor U13158 (N_13158,N_12929,N_12955);
nor U13159 (N_13159,N_12792,N_12597);
nand U13160 (N_13160,N_12909,N_12922);
xnor U13161 (N_13161,N_12773,N_12744);
or U13162 (N_13162,N_12698,N_12878);
nand U13163 (N_13163,N_12754,N_12741);
and U13164 (N_13164,N_12799,N_12644);
nand U13165 (N_13165,N_12958,N_12656);
nand U13166 (N_13166,N_12560,N_12557);
or U13167 (N_13167,N_12649,N_12653);
nand U13168 (N_13168,N_12641,N_12925);
nor U13169 (N_13169,N_12543,N_12737);
nor U13170 (N_13170,N_12984,N_12687);
nor U13171 (N_13171,N_12540,N_12767);
xnor U13172 (N_13172,N_12815,N_12742);
nand U13173 (N_13173,N_12500,N_12787);
nand U13174 (N_13174,N_12544,N_12619);
nor U13175 (N_13175,N_12782,N_12615);
nor U13176 (N_13176,N_12945,N_12514);
nand U13177 (N_13177,N_12885,N_12505);
or U13178 (N_13178,N_12848,N_12743);
nand U13179 (N_13179,N_12959,N_12914);
nor U13180 (N_13180,N_12541,N_12976);
nor U13181 (N_13181,N_12739,N_12814);
or U13182 (N_13182,N_12979,N_12889);
and U13183 (N_13183,N_12683,N_12674);
and U13184 (N_13184,N_12652,N_12906);
and U13185 (N_13185,N_12594,N_12637);
xor U13186 (N_13186,N_12546,N_12850);
or U13187 (N_13187,N_12817,N_12705);
nand U13188 (N_13188,N_12646,N_12706);
xnor U13189 (N_13189,N_12534,N_12670);
or U13190 (N_13190,N_12888,N_12919);
xor U13191 (N_13191,N_12950,N_12764);
nand U13192 (N_13192,N_12582,N_12660);
xnor U13193 (N_13193,N_12596,N_12806);
nand U13194 (N_13194,N_12568,N_12732);
nand U13195 (N_13195,N_12944,N_12760);
xor U13196 (N_13196,N_12624,N_12938);
xor U13197 (N_13197,N_12733,N_12701);
nor U13198 (N_13198,N_12987,N_12861);
or U13199 (N_13199,N_12830,N_12604);
nand U13200 (N_13200,N_12966,N_12868);
nor U13201 (N_13201,N_12577,N_12719);
nor U13202 (N_13202,N_12658,N_12723);
xnor U13203 (N_13203,N_12858,N_12808);
nor U13204 (N_13204,N_12939,N_12620);
nor U13205 (N_13205,N_12667,N_12997);
xor U13206 (N_13206,N_12813,N_12545);
and U13207 (N_13207,N_12622,N_12915);
or U13208 (N_13208,N_12796,N_12962);
nand U13209 (N_13209,N_12632,N_12968);
nand U13210 (N_13210,N_12971,N_12749);
nor U13211 (N_13211,N_12843,N_12847);
or U13212 (N_13212,N_12564,N_12635);
or U13213 (N_13213,N_12745,N_12663);
or U13214 (N_13214,N_12617,N_12895);
or U13215 (N_13215,N_12517,N_12720);
nor U13216 (N_13216,N_12530,N_12769);
and U13217 (N_13217,N_12890,N_12523);
xnor U13218 (N_13218,N_12680,N_12553);
and U13219 (N_13219,N_12591,N_12943);
nor U13220 (N_13220,N_12639,N_12926);
or U13221 (N_13221,N_12538,N_12978);
nor U13222 (N_13222,N_12752,N_12875);
and U13223 (N_13223,N_12735,N_12519);
nand U13224 (N_13224,N_12852,N_12871);
nor U13225 (N_13225,N_12998,N_12819);
and U13226 (N_13226,N_12816,N_12730);
nand U13227 (N_13227,N_12570,N_12809);
or U13228 (N_13228,N_12894,N_12533);
or U13229 (N_13229,N_12636,N_12552);
and U13230 (N_13230,N_12699,N_12974);
xor U13231 (N_13231,N_12618,N_12625);
xnor U13232 (N_13232,N_12903,N_12905);
nor U13233 (N_13233,N_12645,N_12930);
nor U13234 (N_13234,N_12547,N_12563);
nand U13235 (N_13235,N_12911,N_12567);
and U13236 (N_13236,N_12917,N_12982);
nand U13237 (N_13237,N_12734,N_12704);
or U13238 (N_13238,N_12727,N_12824);
and U13239 (N_13239,N_12985,N_12650);
nor U13240 (N_13240,N_12994,N_12794);
and U13241 (N_13241,N_12715,N_12900);
or U13242 (N_13242,N_12910,N_12574);
and U13243 (N_13243,N_12953,N_12970);
xor U13244 (N_13244,N_12779,N_12967);
and U13245 (N_13245,N_12526,N_12709);
nand U13246 (N_13246,N_12673,N_12857);
nor U13247 (N_13247,N_12621,N_12508);
nand U13248 (N_13248,N_12642,N_12942);
xor U13249 (N_13249,N_12963,N_12881);
and U13250 (N_13250,N_12811,N_12653);
xnor U13251 (N_13251,N_12929,N_12610);
and U13252 (N_13252,N_12723,N_12775);
and U13253 (N_13253,N_12776,N_12573);
or U13254 (N_13254,N_12588,N_12557);
nor U13255 (N_13255,N_12885,N_12772);
or U13256 (N_13256,N_12593,N_12868);
nand U13257 (N_13257,N_12998,N_12610);
nor U13258 (N_13258,N_12797,N_12811);
nor U13259 (N_13259,N_12782,N_12938);
or U13260 (N_13260,N_12733,N_12723);
or U13261 (N_13261,N_12776,N_12760);
nand U13262 (N_13262,N_12544,N_12754);
or U13263 (N_13263,N_12746,N_12952);
nor U13264 (N_13264,N_12905,N_12645);
or U13265 (N_13265,N_12917,N_12540);
and U13266 (N_13266,N_12872,N_12949);
and U13267 (N_13267,N_12528,N_12841);
and U13268 (N_13268,N_12750,N_12840);
nor U13269 (N_13269,N_12926,N_12598);
or U13270 (N_13270,N_12888,N_12769);
nand U13271 (N_13271,N_12967,N_12839);
nor U13272 (N_13272,N_12971,N_12554);
and U13273 (N_13273,N_12537,N_12768);
xor U13274 (N_13274,N_12880,N_12740);
or U13275 (N_13275,N_12650,N_12982);
or U13276 (N_13276,N_12601,N_12801);
or U13277 (N_13277,N_12669,N_12583);
and U13278 (N_13278,N_12592,N_12610);
nor U13279 (N_13279,N_12735,N_12878);
nand U13280 (N_13280,N_12890,N_12506);
nor U13281 (N_13281,N_12748,N_12614);
xor U13282 (N_13282,N_12822,N_12983);
nand U13283 (N_13283,N_12742,N_12669);
and U13284 (N_13284,N_12803,N_12959);
or U13285 (N_13285,N_12868,N_12992);
nor U13286 (N_13286,N_12924,N_12712);
nor U13287 (N_13287,N_12855,N_12777);
or U13288 (N_13288,N_12701,N_12566);
xor U13289 (N_13289,N_12715,N_12663);
and U13290 (N_13290,N_12876,N_12784);
and U13291 (N_13291,N_12974,N_12804);
or U13292 (N_13292,N_12704,N_12502);
nor U13293 (N_13293,N_12809,N_12782);
or U13294 (N_13294,N_12956,N_12780);
nand U13295 (N_13295,N_12537,N_12992);
nand U13296 (N_13296,N_12983,N_12688);
nand U13297 (N_13297,N_12860,N_12513);
or U13298 (N_13298,N_12835,N_12762);
or U13299 (N_13299,N_12757,N_12739);
nor U13300 (N_13300,N_12798,N_12982);
or U13301 (N_13301,N_12829,N_12957);
nand U13302 (N_13302,N_12758,N_12602);
nand U13303 (N_13303,N_12547,N_12653);
nor U13304 (N_13304,N_12643,N_12944);
xor U13305 (N_13305,N_12613,N_12552);
or U13306 (N_13306,N_12649,N_12844);
nand U13307 (N_13307,N_12739,N_12626);
or U13308 (N_13308,N_12510,N_12992);
or U13309 (N_13309,N_12653,N_12810);
nand U13310 (N_13310,N_12989,N_12753);
and U13311 (N_13311,N_12673,N_12828);
nand U13312 (N_13312,N_12859,N_12691);
xor U13313 (N_13313,N_12876,N_12660);
or U13314 (N_13314,N_12896,N_12976);
or U13315 (N_13315,N_12710,N_12857);
nand U13316 (N_13316,N_12867,N_12817);
nor U13317 (N_13317,N_12726,N_12705);
and U13318 (N_13318,N_12837,N_12829);
nand U13319 (N_13319,N_12602,N_12841);
nor U13320 (N_13320,N_12580,N_12775);
nand U13321 (N_13321,N_12586,N_12709);
and U13322 (N_13322,N_12942,N_12514);
nor U13323 (N_13323,N_12929,N_12501);
nor U13324 (N_13324,N_12886,N_12805);
and U13325 (N_13325,N_12574,N_12849);
or U13326 (N_13326,N_12542,N_12661);
and U13327 (N_13327,N_12560,N_12849);
and U13328 (N_13328,N_12580,N_12546);
nor U13329 (N_13329,N_12691,N_12703);
nor U13330 (N_13330,N_12547,N_12875);
or U13331 (N_13331,N_12896,N_12986);
and U13332 (N_13332,N_12757,N_12789);
and U13333 (N_13333,N_12902,N_12642);
nor U13334 (N_13334,N_12727,N_12511);
xor U13335 (N_13335,N_12685,N_12857);
nand U13336 (N_13336,N_12787,N_12837);
nand U13337 (N_13337,N_12663,N_12609);
or U13338 (N_13338,N_12963,N_12944);
and U13339 (N_13339,N_12879,N_12609);
and U13340 (N_13340,N_12985,N_12966);
and U13341 (N_13341,N_12949,N_12597);
nor U13342 (N_13342,N_12678,N_12746);
nor U13343 (N_13343,N_12903,N_12979);
xor U13344 (N_13344,N_12662,N_12826);
nand U13345 (N_13345,N_12735,N_12797);
and U13346 (N_13346,N_12571,N_12674);
nor U13347 (N_13347,N_12786,N_12897);
and U13348 (N_13348,N_12957,N_12614);
xor U13349 (N_13349,N_12958,N_12765);
nor U13350 (N_13350,N_12973,N_12504);
nand U13351 (N_13351,N_12550,N_12695);
and U13352 (N_13352,N_12896,N_12882);
or U13353 (N_13353,N_12577,N_12864);
nand U13354 (N_13354,N_12839,N_12866);
nand U13355 (N_13355,N_12813,N_12916);
nor U13356 (N_13356,N_12742,N_12864);
nand U13357 (N_13357,N_12721,N_12574);
nor U13358 (N_13358,N_12779,N_12793);
or U13359 (N_13359,N_12570,N_12873);
nand U13360 (N_13360,N_12611,N_12860);
nand U13361 (N_13361,N_12565,N_12877);
and U13362 (N_13362,N_12625,N_12701);
or U13363 (N_13363,N_12926,N_12761);
or U13364 (N_13364,N_12914,N_12933);
and U13365 (N_13365,N_12628,N_12885);
and U13366 (N_13366,N_12689,N_12601);
nor U13367 (N_13367,N_12685,N_12942);
and U13368 (N_13368,N_12736,N_12971);
nor U13369 (N_13369,N_12705,N_12805);
and U13370 (N_13370,N_12733,N_12930);
nor U13371 (N_13371,N_12636,N_12995);
and U13372 (N_13372,N_12758,N_12579);
or U13373 (N_13373,N_12607,N_12621);
and U13374 (N_13374,N_12561,N_12742);
xor U13375 (N_13375,N_12809,N_12632);
and U13376 (N_13376,N_12522,N_12787);
nand U13377 (N_13377,N_12727,N_12930);
nand U13378 (N_13378,N_12844,N_12587);
and U13379 (N_13379,N_12837,N_12743);
and U13380 (N_13380,N_12785,N_12562);
nor U13381 (N_13381,N_12863,N_12885);
nor U13382 (N_13382,N_12689,N_12871);
nand U13383 (N_13383,N_12707,N_12892);
nor U13384 (N_13384,N_12823,N_12844);
or U13385 (N_13385,N_12714,N_12737);
or U13386 (N_13386,N_12910,N_12967);
nand U13387 (N_13387,N_12588,N_12807);
nor U13388 (N_13388,N_12672,N_12632);
and U13389 (N_13389,N_12919,N_12565);
nor U13390 (N_13390,N_12892,N_12535);
nor U13391 (N_13391,N_12671,N_12563);
xnor U13392 (N_13392,N_12802,N_12599);
and U13393 (N_13393,N_12809,N_12914);
nand U13394 (N_13394,N_12611,N_12999);
and U13395 (N_13395,N_12856,N_12720);
nor U13396 (N_13396,N_12788,N_12959);
and U13397 (N_13397,N_12519,N_12825);
and U13398 (N_13398,N_12764,N_12868);
nand U13399 (N_13399,N_12690,N_12632);
or U13400 (N_13400,N_12624,N_12977);
nand U13401 (N_13401,N_12690,N_12513);
or U13402 (N_13402,N_12918,N_12508);
nor U13403 (N_13403,N_12533,N_12534);
nor U13404 (N_13404,N_12862,N_12676);
or U13405 (N_13405,N_12616,N_12909);
nor U13406 (N_13406,N_12997,N_12986);
nand U13407 (N_13407,N_12824,N_12661);
xnor U13408 (N_13408,N_12786,N_12862);
and U13409 (N_13409,N_12835,N_12513);
and U13410 (N_13410,N_12553,N_12931);
nand U13411 (N_13411,N_12683,N_12612);
or U13412 (N_13412,N_12594,N_12715);
and U13413 (N_13413,N_12632,N_12732);
nand U13414 (N_13414,N_12762,N_12673);
nor U13415 (N_13415,N_12503,N_12928);
nand U13416 (N_13416,N_12935,N_12602);
nand U13417 (N_13417,N_12720,N_12597);
nand U13418 (N_13418,N_12849,N_12889);
nand U13419 (N_13419,N_12738,N_12526);
nand U13420 (N_13420,N_12801,N_12706);
and U13421 (N_13421,N_12616,N_12742);
and U13422 (N_13422,N_12753,N_12735);
and U13423 (N_13423,N_12656,N_12723);
nor U13424 (N_13424,N_12576,N_12613);
nand U13425 (N_13425,N_12883,N_12666);
and U13426 (N_13426,N_12782,N_12533);
nand U13427 (N_13427,N_12669,N_12594);
nor U13428 (N_13428,N_12642,N_12612);
or U13429 (N_13429,N_12661,N_12626);
nor U13430 (N_13430,N_12674,N_12879);
or U13431 (N_13431,N_12796,N_12710);
and U13432 (N_13432,N_12611,N_12567);
nor U13433 (N_13433,N_12589,N_12508);
and U13434 (N_13434,N_12577,N_12838);
xor U13435 (N_13435,N_12599,N_12916);
and U13436 (N_13436,N_12672,N_12565);
and U13437 (N_13437,N_12737,N_12744);
nor U13438 (N_13438,N_12680,N_12783);
nor U13439 (N_13439,N_12921,N_12602);
xor U13440 (N_13440,N_12756,N_12615);
nand U13441 (N_13441,N_12932,N_12711);
nand U13442 (N_13442,N_12665,N_12716);
nor U13443 (N_13443,N_12542,N_12665);
and U13444 (N_13444,N_12990,N_12802);
or U13445 (N_13445,N_12728,N_12636);
nand U13446 (N_13446,N_12846,N_12815);
or U13447 (N_13447,N_12934,N_12835);
nor U13448 (N_13448,N_12618,N_12891);
and U13449 (N_13449,N_12761,N_12503);
nand U13450 (N_13450,N_12842,N_12700);
nor U13451 (N_13451,N_12549,N_12508);
nor U13452 (N_13452,N_12876,N_12767);
and U13453 (N_13453,N_12594,N_12602);
or U13454 (N_13454,N_12628,N_12785);
nor U13455 (N_13455,N_12861,N_12722);
nand U13456 (N_13456,N_12746,N_12751);
or U13457 (N_13457,N_12711,N_12961);
nor U13458 (N_13458,N_12693,N_12665);
nand U13459 (N_13459,N_12932,N_12844);
nor U13460 (N_13460,N_12634,N_12600);
nor U13461 (N_13461,N_12621,N_12691);
xnor U13462 (N_13462,N_12619,N_12830);
and U13463 (N_13463,N_12666,N_12876);
xor U13464 (N_13464,N_12749,N_12587);
or U13465 (N_13465,N_12964,N_12945);
nor U13466 (N_13466,N_12574,N_12961);
nand U13467 (N_13467,N_12705,N_12590);
nor U13468 (N_13468,N_12980,N_12864);
and U13469 (N_13469,N_12616,N_12976);
nand U13470 (N_13470,N_12640,N_12962);
or U13471 (N_13471,N_12527,N_12725);
or U13472 (N_13472,N_12572,N_12623);
nor U13473 (N_13473,N_12820,N_12920);
and U13474 (N_13474,N_12875,N_12597);
and U13475 (N_13475,N_12850,N_12998);
or U13476 (N_13476,N_12562,N_12680);
or U13477 (N_13477,N_12886,N_12851);
and U13478 (N_13478,N_12674,N_12947);
nand U13479 (N_13479,N_12618,N_12793);
or U13480 (N_13480,N_12822,N_12516);
nand U13481 (N_13481,N_12919,N_12977);
and U13482 (N_13482,N_12968,N_12541);
or U13483 (N_13483,N_12830,N_12720);
xnor U13484 (N_13484,N_12530,N_12785);
nor U13485 (N_13485,N_12507,N_12593);
and U13486 (N_13486,N_12583,N_12831);
and U13487 (N_13487,N_12508,N_12780);
or U13488 (N_13488,N_12754,N_12822);
and U13489 (N_13489,N_12951,N_12593);
nand U13490 (N_13490,N_12563,N_12868);
and U13491 (N_13491,N_12506,N_12733);
nor U13492 (N_13492,N_12993,N_12940);
or U13493 (N_13493,N_12801,N_12932);
or U13494 (N_13494,N_12542,N_12906);
nor U13495 (N_13495,N_12535,N_12807);
or U13496 (N_13496,N_12585,N_12928);
nand U13497 (N_13497,N_12825,N_12550);
or U13498 (N_13498,N_12630,N_12961);
and U13499 (N_13499,N_12550,N_12910);
and U13500 (N_13500,N_13312,N_13092);
xnor U13501 (N_13501,N_13222,N_13063);
nand U13502 (N_13502,N_13045,N_13382);
nand U13503 (N_13503,N_13004,N_13113);
and U13504 (N_13504,N_13325,N_13460);
and U13505 (N_13505,N_13474,N_13193);
xnor U13506 (N_13506,N_13061,N_13131);
and U13507 (N_13507,N_13095,N_13040);
or U13508 (N_13508,N_13455,N_13087);
nand U13509 (N_13509,N_13009,N_13037);
nand U13510 (N_13510,N_13191,N_13082);
nand U13511 (N_13511,N_13297,N_13362);
or U13512 (N_13512,N_13167,N_13052);
nor U13513 (N_13513,N_13072,N_13376);
or U13514 (N_13514,N_13258,N_13392);
xnor U13515 (N_13515,N_13238,N_13085);
nor U13516 (N_13516,N_13070,N_13013);
or U13517 (N_13517,N_13340,N_13133);
or U13518 (N_13518,N_13233,N_13399);
xor U13519 (N_13519,N_13111,N_13398);
and U13520 (N_13520,N_13213,N_13093);
nor U13521 (N_13521,N_13304,N_13026);
or U13522 (N_13522,N_13302,N_13059);
nor U13523 (N_13523,N_13003,N_13378);
or U13524 (N_13524,N_13469,N_13029);
nor U13525 (N_13525,N_13413,N_13465);
xnor U13526 (N_13526,N_13106,N_13114);
nor U13527 (N_13527,N_13220,N_13300);
and U13528 (N_13528,N_13162,N_13475);
or U13529 (N_13529,N_13083,N_13478);
nand U13530 (N_13530,N_13268,N_13492);
nand U13531 (N_13531,N_13326,N_13195);
or U13532 (N_13532,N_13089,N_13159);
and U13533 (N_13533,N_13345,N_13077);
or U13534 (N_13534,N_13034,N_13311);
nand U13535 (N_13535,N_13110,N_13036);
nor U13536 (N_13536,N_13301,N_13410);
or U13537 (N_13537,N_13482,N_13486);
nand U13538 (N_13538,N_13384,N_13174);
and U13539 (N_13539,N_13188,N_13314);
nand U13540 (N_13540,N_13002,N_13256);
and U13541 (N_13541,N_13352,N_13155);
xnor U13542 (N_13542,N_13309,N_13246);
xnor U13543 (N_13543,N_13494,N_13221);
nor U13544 (N_13544,N_13489,N_13338);
nand U13545 (N_13545,N_13138,N_13261);
xor U13546 (N_13546,N_13423,N_13129);
xnor U13547 (N_13547,N_13480,N_13315);
and U13548 (N_13548,N_13028,N_13288);
nand U13549 (N_13549,N_13019,N_13344);
xnor U13550 (N_13550,N_13347,N_13463);
nor U13551 (N_13551,N_13086,N_13144);
nor U13552 (N_13552,N_13435,N_13397);
and U13553 (N_13553,N_13068,N_13183);
xnor U13554 (N_13554,N_13441,N_13043);
or U13555 (N_13555,N_13108,N_13056);
or U13556 (N_13556,N_13281,N_13449);
or U13557 (N_13557,N_13198,N_13065);
and U13558 (N_13558,N_13042,N_13137);
nand U13559 (N_13559,N_13411,N_13454);
nor U13560 (N_13560,N_13151,N_13098);
nor U13561 (N_13561,N_13287,N_13308);
and U13562 (N_13562,N_13296,N_13263);
nand U13563 (N_13563,N_13430,N_13060);
nand U13564 (N_13564,N_13030,N_13130);
nor U13565 (N_13565,N_13270,N_13136);
nor U13566 (N_13566,N_13425,N_13395);
or U13567 (N_13567,N_13359,N_13126);
and U13568 (N_13568,N_13280,N_13484);
and U13569 (N_13569,N_13217,N_13402);
and U13570 (N_13570,N_13283,N_13274);
nor U13571 (N_13571,N_13023,N_13205);
and U13572 (N_13572,N_13374,N_13289);
nand U13573 (N_13573,N_13215,N_13244);
or U13574 (N_13574,N_13496,N_13324);
nand U13575 (N_13575,N_13192,N_13127);
or U13576 (N_13576,N_13462,N_13365);
nor U13577 (N_13577,N_13421,N_13457);
nand U13578 (N_13578,N_13225,N_13190);
nor U13579 (N_13579,N_13400,N_13153);
or U13580 (N_13580,N_13212,N_13169);
nand U13581 (N_13581,N_13208,N_13424);
nand U13582 (N_13582,N_13418,N_13495);
or U13583 (N_13583,N_13154,N_13076);
nand U13584 (N_13584,N_13305,N_13237);
nand U13585 (N_13585,N_13440,N_13267);
or U13586 (N_13586,N_13391,N_13416);
or U13587 (N_13587,N_13331,N_13223);
or U13588 (N_13588,N_13269,N_13016);
nor U13589 (N_13589,N_13409,N_13071);
nand U13590 (N_13590,N_13211,N_13243);
xnor U13591 (N_13591,N_13158,N_13218);
nand U13592 (N_13592,N_13290,N_13118);
nand U13593 (N_13593,N_13363,N_13292);
or U13594 (N_13594,N_13091,N_13079);
nand U13595 (N_13595,N_13354,N_13249);
nor U13596 (N_13596,N_13135,N_13104);
or U13597 (N_13597,N_13172,N_13229);
or U13598 (N_13598,N_13214,N_13149);
nand U13599 (N_13599,N_13011,N_13055);
nor U13600 (N_13600,N_13005,N_13240);
or U13601 (N_13601,N_13075,N_13176);
xor U13602 (N_13602,N_13485,N_13039);
or U13603 (N_13603,N_13447,N_13487);
nor U13604 (N_13604,N_13342,N_13022);
or U13605 (N_13605,N_13181,N_13147);
and U13606 (N_13606,N_13250,N_13184);
nand U13607 (N_13607,N_13069,N_13049);
and U13608 (N_13608,N_13320,N_13027);
nand U13609 (N_13609,N_13241,N_13255);
nor U13610 (N_13610,N_13081,N_13295);
and U13611 (N_13611,N_13146,N_13349);
or U13612 (N_13612,N_13259,N_13335);
nor U13613 (N_13613,N_13206,N_13096);
xnor U13614 (N_13614,N_13128,N_13367);
xnor U13615 (N_13615,N_13000,N_13330);
nand U13616 (N_13616,N_13429,N_13401);
and U13617 (N_13617,N_13178,N_13414);
or U13618 (N_13618,N_13053,N_13119);
nand U13619 (N_13619,N_13168,N_13031);
nor U13620 (N_13620,N_13062,N_13386);
nand U13621 (N_13621,N_13080,N_13007);
and U13622 (N_13622,N_13318,N_13385);
and U13623 (N_13623,N_13124,N_13317);
or U13624 (N_13624,N_13125,N_13235);
and U13625 (N_13625,N_13074,N_13464);
nor U13626 (N_13626,N_13142,N_13064);
and U13627 (N_13627,N_13476,N_13293);
xnor U13628 (N_13628,N_13099,N_13383);
nor U13629 (N_13629,N_13390,N_13008);
or U13630 (N_13630,N_13035,N_13444);
nor U13631 (N_13631,N_13490,N_13373);
nand U13632 (N_13632,N_13251,N_13298);
and U13633 (N_13633,N_13445,N_13497);
and U13634 (N_13634,N_13185,N_13156);
nor U13635 (N_13635,N_13145,N_13471);
nand U13636 (N_13636,N_13182,N_13433);
or U13637 (N_13637,N_13117,N_13219);
xnor U13638 (N_13638,N_13434,N_13406);
and U13639 (N_13639,N_13361,N_13372);
nand U13640 (N_13640,N_13291,N_13199);
xor U13641 (N_13641,N_13278,N_13247);
or U13642 (N_13642,N_13366,N_13179);
nand U13643 (N_13643,N_13470,N_13100);
nand U13644 (N_13644,N_13122,N_13266);
nand U13645 (N_13645,N_13187,N_13341);
nand U13646 (N_13646,N_13321,N_13488);
and U13647 (N_13647,N_13157,N_13186);
nor U13648 (N_13648,N_13033,N_13426);
nor U13649 (N_13649,N_13499,N_13436);
xor U13650 (N_13650,N_13044,N_13346);
and U13651 (N_13651,N_13058,N_13336);
and U13652 (N_13652,N_13403,N_13405);
and U13653 (N_13653,N_13066,N_13306);
xor U13654 (N_13654,N_13407,N_13348);
or U13655 (N_13655,N_13264,N_13275);
nor U13656 (N_13656,N_13163,N_13328);
nor U13657 (N_13657,N_13101,N_13015);
nor U13658 (N_13658,N_13282,N_13006);
nor U13659 (N_13659,N_13166,N_13161);
xor U13660 (N_13660,N_13116,N_13332);
nand U13661 (N_13661,N_13189,N_13364);
nor U13662 (N_13662,N_13160,N_13356);
nor U13663 (N_13663,N_13276,N_13369);
or U13664 (N_13664,N_13201,N_13232);
or U13665 (N_13665,N_13438,N_13084);
nand U13666 (N_13666,N_13360,N_13001);
nor U13667 (N_13667,N_13236,N_13017);
nor U13668 (N_13668,N_13242,N_13253);
and U13669 (N_13669,N_13450,N_13358);
and U13670 (N_13670,N_13210,N_13396);
nor U13671 (N_13671,N_13048,N_13472);
or U13672 (N_13672,N_13097,N_13483);
and U13673 (N_13673,N_13134,N_13196);
xor U13674 (N_13674,N_13123,N_13164);
and U13675 (N_13675,N_13032,N_13299);
xor U13676 (N_13676,N_13073,N_13428);
nand U13677 (N_13677,N_13307,N_13025);
nor U13678 (N_13678,N_13094,N_13226);
nand U13679 (N_13679,N_13047,N_13265);
nor U13680 (N_13680,N_13046,N_13024);
nand U13681 (N_13681,N_13377,N_13173);
and U13682 (N_13682,N_13078,N_13417);
nor U13683 (N_13683,N_13415,N_13197);
nand U13684 (N_13684,N_13313,N_13468);
or U13685 (N_13685,N_13466,N_13432);
xnor U13686 (N_13686,N_13054,N_13143);
and U13687 (N_13687,N_13453,N_13171);
or U13688 (N_13688,N_13140,N_13343);
or U13689 (N_13689,N_13194,N_13148);
and U13690 (N_13690,N_13443,N_13393);
or U13691 (N_13691,N_13209,N_13088);
nor U13692 (N_13692,N_13408,N_13170);
xnor U13693 (N_13693,N_13254,N_13412);
and U13694 (N_13694,N_13310,N_13370);
or U13695 (N_13695,N_13014,N_13458);
and U13696 (N_13696,N_13446,N_13021);
and U13697 (N_13697,N_13090,N_13277);
or U13698 (N_13698,N_13051,N_13448);
or U13699 (N_13699,N_13422,N_13120);
or U13700 (N_13700,N_13351,N_13459);
or U13701 (N_13701,N_13105,N_13067);
nor U13702 (N_13702,N_13319,N_13285);
nor U13703 (N_13703,N_13467,N_13473);
xor U13704 (N_13704,N_13057,N_13177);
and U13705 (N_13705,N_13404,N_13389);
nor U13706 (N_13706,N_13491,N_13286);
and U13707 (N_13707,N_13224,N_13175);
or U13708 (N_13708,N_13150,N_13481);
and U13709 (N_13709,N_13165,N_13050);
or U13710 (N_13710,N_13273,N_13020);
or U13711 (N_13711,N_13252,N_13323);
nor U13712 (N_13712,N_13204,N_13322);
and U13713 (N_13713,N_13334,N_13420);
and U13714 (N_13714,N_13303,N_13394);
nand U13715 (N_13715,N_13234,N_13271);
and U13716 (N_13716,N_13350,N_13333);
or U13717 (N_13717,N_13231,N_13461);
nand U13718 (N_13718,N_13316,N_13442);
or U13719 (N_13719,N_13010,N_13437);
xor U13720 (N_13720,N_13477,N_13257);
or U13721 (N_13721,N_13379,N_13115);
nor U13722 (N_13722,N_13041,N_13498);
and U13723 (N_13723,N_13239,N_13109);
nor U13724 (N_13724,N_13431,N_13357);
or U13725 (N_13725,N_13207,N_13375);
nor U13726 (N_13726,N_13368,N_13112);
nor U13727 (N_13727,N_13227,N_13228);
or U13728 (N_13728,N_13279,N_13132);
xnor U13729 (N_13729,N_13294,N_13107);
and U13730 (N_13730,N_13339,N_13427);
and U13731 (N_13731,N_13419,N_13387);
nor U13732 (N_13732,N_13284,N_13451);
or U13733 (N_13733,N_13038,N_13439);
and U13734 (N_13734,N_13456,N_13381);
xnor U13735 (N_13735,N_13012,N_13180);
nor U13736 (N_13736,N_13141,N_13230);
nand U13737 (N_13737,N_13018,N_13262);
xnor U13738 (N_13738,N_13353,N_13203);
nand U13739 (N_13739,N_13327,N_13380);
or U13740 (N_13740,N_13200,N_13121);
or U13741 (N_13741,N_13329,N_13139);
or U13742 (N_13742,N_13452,N_13245);
xnor U13743 (N_13743,N_13388,N_13202);
or U13744 (N_13744,N_13102,N_13371);
nor U13745 (N_13745,N_13355,N_13272);
nor U13746 (N_13746,N_13216,N_13479);
nor U13747 (N_13747,N_13493,N_13337);
or U13748 (N_13748,N_13152,N_13248);
xor U13749 (N_13749,N_13260,N_13103);
and U13750 (N_13750,N_13227,N_13180);
or U13751 (N_13751,N_13171,N_13491);
and U13752 (N_13752,N_13442,N_13437);
nor U13753 (N_13753,N_13226,N_13494);
and U13754 (N_13754,N_13198,N_13355);
nand U13755 (N_13755,N_13211,N_13061);
and U13756 (N_13756,N_13381,N_13303);
nand U13757 (N_13757,N_13438,N_13279);
or U13758 (N_13758,N_13159,N_13434);
or U13759 (N_13759,N_13401,N_13212);
nor U13760 (N_13760,N_13228,N_13392);
xnor U13761 (N_13761,N_13102,N_13498);
or U13762 (N_13762,N_13114,N_13217);
or U13763 (N_13763,N_13244,N_13178);
or U13764 (N_13764,N_13320,N_13111);
and U13765 (N_13765,N_13156,N_13002);
nor U13766 (N_13766,N_13000,N_13407);
or U13767 (N_13767,N_13061,N_13478);
xnor U13768 (N_13768,N_13014,N_13245);
and U13769 (N_13769,N_13299,N_13487);
and U13770 (N_13770,N_13367,N_13242);
nor U13771 (N_13771,N_13191,N_13282);
xnor U13772 (N_13772,N_13169,N_13221);
xor U13773 (N_13773,N_13011,N_13043);
or U13774 (N_13774,N_13301,N_13379);
nand U13775 (N_13775,N_13092,N_13486);
nor U13776 (N_13776,N_13161,N_13173);
or U13777 (N_13777,N_13231,N_13307);
and U13778 (N_13778,N_13268,N_13348);
nor U13779 (N_13779,N_13421,N_13414);
nand U13780 (N_13780,N_13061,N_13066);
xnor U13781 (N_13781,N_13400,N_13159);
nor U13782 (N_13782,N_13027,N_13236);
nor U13783 (N_13783,N_13440,N_13173);
nor U13784 (N_13784,N_13380,N_13292);
and U13785 (N_13785,N_13044,N_13393);
nand U13786 (N_13786,N_13293,N_13350);
nand U13787 (N_13787,N_13031,N_13346);
nand U13788 (N_13788,N_13063,N_13379);
nand U13789 (N_13789,N_13049,N_13311);
nand U13790 (N_13790,N_13294,N_13218);
and U13791 (N_13791,N_13147,N_13489);
nor U13792 (N_13792,N_13244,N_13428);
and U13793 (N_13793,N_13391,N_13323);
and U13794 (N_13794,N_13490,N_13244);
or U13795 (N_13795,N_13013,N_13066);
nor U13796 (N_13796,N_13266,N_13270);
and U13797 (N_13797,N_13337,N_13043);
or U13798 (N_13798,N_13161,N_13444);
nand U13799 (N_13799,N_13161,N_13391);
nand U13800 (N_13800,N_13064,N_13028);
nand U13801 (N_13801,N_13152,N_13492);
xor U13802 (N_13802,N_13038,N_13054);
nand U13803 (N_13803,N_13344,N_13435);
nand U13804 (N_13804,N_13384,N_13290);
or U13805 (N_13805,N_13353,N_13157);
and U13806 (N_13806,N_13049,N_13355);
nor U13807 (N_13807,N_13054,N_13388);
xor U13808 (N_13808,N_13252,N_13408);
or U13809 (N_13809,N_13259,N_13129);
and U13810 (N_13810,N_13486,N_13119);
or U13811 (N_13811,N_13321,N_13348);
nand U13812 (N_13812,N_13364,N_13477);
nand U13813 (N_13813,N_13267,N_13469);
or U13814 (N_13814,N_13080,N_13115);
nand U13815 (N_13815,N_13307,N_13109);
or U13816 (N_13816,N_13285,N_13186);
nand U13817 (N_13817,N_13371,N_13228);
nor U13818 (N_13818,N_13070,N_13484);
nor U13819 (N_13819,N_13255,N_13063);
or U13820 (N_13820,N_13067,N_13495);
nand U13821 (N_13821,N_13310,N_13223);
or U13822 (N_13822,N_13294,N_13313);
and U13823 (N_13823,N_13173,N_13485);
and U13824 (N_13824,N_13145,N_13384);
xor U13825 (N_13825,N_13196,N_13494);
or U13826 (N_13826,N_13119,N_13172);
and U13827 (N_13827,N_13180,N_13499);
and U13828 (N_13828,N_13308,N_13405);
nor U13829 (N_13829,N_13369,N_13379);
and U13830 (N_13830,N_13455,N_13106);
or U13831 (N_13831,N_13186,N_13027);
and U13832 (N_13832,N_13352,N_13069);
or U13833 (N_13833,N_13265,N_13412);
nand U13834 (N_13834,N_13172,N_13023);
or U13835 (N_13835,N_13359,N_13170);
or U13836 (N_13836,N_13485,N_13432);
nor U13837 (N_13837,N_13090,N_13169);
and U13838 (N_13838,N_13231,N_13415);
nand U13839 (N_13839,N_13087,N_13186);
or U13840 (N_13840,N_13102,N_13025);
and U13841 (N_13841,N_13334,N_13235);
nor U13842 (N_13842,N_13087,N_13273);
or U13843 (N_13843,N_13104,N_13055);
and U13844 (N_13844,N_13025,N_13411);
and U13845 (N_13845,N_13327,N_13173);
nor U13846 (N_13846,N_13158,N_13284);
and U13847 (N_13847,N_13470,N_13131);
nand U13848 (N_13848,N_13145,N_13287);
and U13849 (N_13849,N_13086,N_13057);
nand U13850 (N_13850,N_13213,N_13345);
nor U13851 (N_13851,N_13377,N_13011);
nand U13852 (N_13852,N_13201,N_13197);
and U13853 (N_13853,N_13051,N_13100);
nand U13854 (N_13854,N_13442,N_13172);
nand U13855 (N_13855,N_13464,N_13209);
and U13856 (N_13856,N_13453,N_13021);
nand U13857 (N_13857,N_13367,N_13200);
xor U13858 (N_13858,N_13472,N_13316);
xnor U13859 (N_13859,N_13446,N_13294);
nand U13860 (N_13860,N_13252,N_13444);
and U13861 (N_13861,N_13478,N_13439);
xor U13862 (N_13862,N_13360,N_13363);
and U13863 (N_13863,N_13162,N_13342);
or U13864 (N_13864,N_13180,N_13484);
or U13865 (N_13865,N_13011,N_13044);
or U13866 (N_13866,N_13403,N_13133);
nor U13867 (N_13867,N_13310,N_13147);
nand U13868 (N_13868,N_13406,N_13385);
xnor U13869 (N_13869,N_13065,N_13248);
nor U13870 (N_13870,N_13142,N_13036);
nand U13871 (N_13871,N_13045,N_13007);
or U13872 (N_13872,N_13420,N_13081);
xor U13873 (N_13873,N_13104,N_13288);
nor U13874 (N_13874,N_13202,N_13163);
or U13875 (N_13875,N_13024,N_13094);
xor U13876 (N_13876,N_13016,N_13489);
and U13877 (N_13877,N_13034,N_13108);
nand U13878 (N_13878,N_13499,N_13481);
nand U13879 (N_13879,N_13383,N_13455);
nor U13880 (N_13880,N_13348,N_13185);
nor U13881 (N_13881,N_13436,N_13350);
xor U13882 (N_13882,N_13348,N_13277);
xnor U13883 (N_13883,N_13049,N_13486);
and U13884 (N_13884,N_13052,N_13179);
and U13885 (N_13885,N_13436,N_13351);
or U13886 (N_13886,N_13322,N_13050);
and U13887 (N_13887,N_13038,N_13238);
and U13888 (N_13888,N_13084,N_13057);
and U13889 (N_13889,N_13423,N_13265);
nor U13890 (N_13890,N_13004,N_13114);
or U13891 (N_13891,N_13049,N_13002);
or U13892 (N_13892,N_13023,N_13012);
and U13893 (N_13893,N_13179,N_13008);
nand U13894 (N_13894,N_13325,N_13046);
or U13895 (N_13895,N_13440,N_13363);
nor U13896 (N_13896,N_13481,N_13296);
nor U13897 (N_13897,N_13083,N_13452);
and U13898 (N_13898,N_13162,N_13499);
and U13899 (N_13899,N_13170,N_13045);
nand U13900 (N_13900,N_13260,N_13479);
and U13901 (N_13901,N_13013,N_13306);
nand U13902 (N_13902,N_13057,N_13226);
or U13903 (N_13903,N_13043,N_13476);
or U13904 (N_13904,N_13491,N_13170);
nand U13905 (N_13905,N_13387,N_13341);
and U13906 (N_13906,N_13104,N_13372);
or U13907 (N_13907,N_13149,N_13435);
xnor U13908 (N_13908,N_13178,N_13297);
nor U13909 (N_13909,N_13335,N_13003);
nor U13910 (N_13910,N_13185,N_13124);
nor U13911 (N_13911,N_13084,N_13148);
nor U13912 (N_13912,N_13491,N_13407);
nand U13913 (N_13913,N_13155,N_13328);
nand U13914 (N_13914,N_13176,N_13355);
or U13915 (N_13915,N_13160,N_13163);
and U13916 (N_13916,N_13395,N_13394);
or U13917 (N_13917,N_13120,N_13122);
nand U13918 (N_13918,N_13013,N_13036);
or U13919 (N_13919,N_13136,N_13056);
nor U13920 (N_13920,N_13068,N_13374);
nor U13921 (N_13921,N_13063,N_13484);
nand U13922 (N_13922,N_13303,N_13116);
nand U13923 (N_13923,N_13247,N_13240);
and U13924 (N_13924,N_13183,N_13057);
and U13925 (N_13925,N_13181,N_13082);
or U13926 (N_13926,N_13187,N_13342);
or U13927 (N_13927,N_13460,N_13024);
or U13928 (N_13928,N_13073,N_13188);
nor U13929 (N_13929,N_13451,N_13292);
nand U13930 (N_13930,N_13450,N_13070);
and U13931 (N_13931,N_13001,N_13169);
and U13932 (N_13932,N_13480,N_13305);
xnor U13933 (N_13933,N_13036,N_13240);
nand U13934 (N_13934,N_13332,N_13061);
xnor U13935 (N_13935,N_13475,N_13145);
nand U13936 (N_13936,N_13309,N_13345);
nand U13937 (N_13937,N_13138,N_13495);
and U13938 (N_13938,N_13216,N_13197);
and U13939 (N_13939,N_13072,N_13239);
and U13940 (N_13940,N_13203,N_13069);
nand U13941 (N_13941,N_13484,N_13093);
nor U13942 (N_13942,N_13478,N_13060);
or U13943 (N_13943,N_13204,N_13064);
xor U13944 (N_13944,N_13227,N_13205);
nand U13945 (N_13945,N_13033,N_13364);
or U13946 (N_13946,N_13000,N_13188);
nor U13947 (N_13947,N_13340,N_13267);
or U13948 (N_13948,N_13469,N_13376);
and U13949 (N_13949,N_13369,N_13495);
xor U13950 (N_13950,N_13218,N_13204);
nand U13951 (N_13951,N_13435,N_13452);
or U13952 (N_13952,N_13360,N_13119);
and U13953 (N_13953,N_13318,N_13080);
nand U13954 (N_13954,N_13211,N_13386);
and U13955 (N_13955,N_13352,N_13323);
xor U13956 (N_13956,N_13330,N_13134);
nor U13957 (N_13957,N_13362,N_13285);
or U13958 (N_13958,N_13323,N_13152);
nand U13959 (N_13959,N_13253,N_13316);
or U13960 (N_13960,N_13473,N_13059);
nor U13961 (N_13961,N_13251,N_13436);
xor U13962 (N_13962,N_13041,N_13187);
nand U13963 (N_13963,N_13402,N_13277);
or U13964 (N_13964,N_13468,N_13443);
nand U13965 (N_13965,N_13236,N_13477);
nor U13966 (N_13966,N_13248,N_13123);
nand U13967 (N_13967,N_13279,N_13339);
or U13968 (N_13968,N_13212,N_13248);
nor U13969 (N_13969,N_13371,N_13053);
nor U13970 (N_13970,N_13457,N_13376);
or U13971 (N_13971,N_13171,N_13193);
nor U13972 (N_13972,N_13009,N_13317);
xor U13973 (N_13973,N_13453,N_13064);
xor U13974 (N_13974,N_13028,N_13272);
and U13975 (N_13975,N_13037,N_13150);
nand U13976 (N_13976,N_13390,N_13017);
or U13977 (N_13977,N_13173,N_13105);
nand U13978 (N_13978,N_13291,N_13164);
or U13979 (N_13979,N_13398,N_13193);
xnor U13980 (N_13980,N_13407,N_13183);
or U13981 (N_13981,N_13387,N_13127);
or U13982 (N_13982,N_13247,N_13402);
nor U13983 (N_13983,N_13033,N_13273);
nor U13984 (N_13984,N_13016,N_13057);
nor U13985 (N_13985,N_13449,N_13166);
nor U13986 (N_13986,N_13027,N_13265);
and U13987 (N_13987,N_13234,N_13115);
xor U13988 (N_13988,N_13108,N_13388);
xnor U13989 (N_13989,N_13339,N_13161);
nor U13990 (N_13990,N_13377,N_13441);
and U13991 (N_13991,N_13385,N_13272);
nor U13992 (N_13992,N_13009,N_13271);
nand U13993 (N_13993,N_13078,N_13470);
nand U13994 (N_13994,N_13470,N_13272);
and U13995 (N_13995,N_13134,N_13463);
nor U13996 (N_13996,N_13422,N_13188);
nand U13997 (N_13997,N_13283,N_13154);
xor U13998 (N_13998,N_13169,N_13390);
and U13999 (N_13999,N_13273,N_13145);
or U14000 (N_14000,N_13787,N_13709);
or U14001 (N_14001,N_13953,N_13774);
xor U14002 (N_14002,N_13678,N_13745);
or U14003 (N_14003,N_13917,N_13796);
and U14004 (N_14004,N_13508,N_13880);
or U14005 (N_14005,N_13510,N_13962);
and U14006 (N_14006,N_13506,N_13977);
nand U14007 (N_14007,N_13795,N_13575);
or U14008 (N_14008,N_13927,N_13567);
and U14009 (N_14009,N_13714,N_13680);
nor U14010 (N_14010,N_13667,N_13625);
xor U14011 (N_14011,N_13932,N_13650);
nand U14012 (N_14012,N_13525,N_13549);
nor U14013 (N_14013,N_13729,N_13583);
nor U14014 (N_14014,N_13644,N_13829);
and U14015 (N_14015,N_13949,N_13775);
or U14016 (N_14016,N_13661,N_13719);
nand U14017 (N_14017,N_13532,N_13755);
nand U14018 (N_14018,N_13684,N_13915);
nor U14019 (N_14019,N_13867,N_13564);
nand U14020 (N_14020,N_13903,N_13612);
nor U14021 (N_14021,N_13986,N_13555);
nor U14022 (N_14022,N_13766,N_13842);
nor U14023 (N_14023,N_13582,N_13744);
or U14024 (N_14024,N_13733,N_13788);
xor U14025 (N_14025,N_13891,N_13534);
nand U14026 (N_14026,N_13707,N_13754);
nand U14027 (N_14027,N_13770,N_13780);
xor U14028 (N_14028,N_13634,N_13799);
or U14029 (N_14029,N_13852,N_13598);
and U14030 (N_14030,N_13548,N_13771);
and U14031 (N_14031,N_13964,N_13654);
or U14032 (N_14032,N_13646,N_13621);
xor U14033 (N_14033,N_13991,N_13809);
or U14034 (N_14034,N_13854,N_13984);
or U14035 (N_14035,N_13730,N_13833);
or U14036 (N_14036,N_13703,N_13942);
and U14037 (N_14037,N_13988,N_13820);
nand U14038 (N_14038,N_13956,N_13528);
and U14039 (N_14039,N_13793,N_13571);
nand U14040 (N_14040,N_13702,N_13831);
nand U14041 (N_14041,N_13577,N_13839);
nor U14042 (N_14042,N_13906,N_13562);
nand U14043 (N_14043,N_13605,N_13759);
or U14044 (N_14044,N_13551,N_13732);
and U14045 (N_14045,N_13761,N_13686);
nor U14046 (N_14046,N_13887,N_13655);
nand U14047 (N_14047,N_13731,N_13950);
nand U14048 (N_14048,N_13993,N_13804);
or U14049 (N_14049,N_13519,N_13692);
nand U14050 (N_14050,N_13837,N_13767);
nor U14051 (N_14051,N_13924,N_13568);
nor U14052 (N_14052,N_13936,N_13723);
nor U14053 (N_14053,N_13537,N_13890);
nand U14054 (N_14054,N_13981,N_13581);
nor U14055 (N_14055,N_13710,N_13836);
or U14056 (N_14056,N_13619,N_13700);
nor U14057 (N_14057,N_13560,N_13687);
nor U14058 (N_14058,N_13615,N_13756);
nor U14059 (N_14059,N_13651,N_13800);
nor U14060 (N_14060,N_13789,N_13504);
xor U14061 (N_14061,N_13943,N_13859);
or U14062 (N_14062,N_13827,N_13566);
xor U14063 (N_14063,N_13810,N_13814);
or U14064 (N_14064,N_13670,N_13841);
nand U14065 (N_14065,N_13585,N_13899);
xnor U14066 (N_14066,N_13630,N_13921);
or U14067 (N_14067,N_13706,N_13955);
nand U14068 (N_14068,N_13769,N_13613);
nand U14069 (N_14069,N_13838,N_13864);
or U14070 (N_14070,N_13987,N_13503);
nand U14071 (N_14071,N_13892,N_13524);
and U14072 (N_14072,N_13606,N_13860);
xnor U14073 (N_14073,N_13967,N_13965);
xor U14074 (N_14074,N_13657,N_13970);
or U14075 (N_14075,N_13505,N_13725);
nor U14076 (N_14076,N_13999,N_13747);
and U14077 (N_14077,N_13749,N_13996);
and U14078 (N_14078,N_13816,N_13570);
and U14079 (N_14079,N_13527,N_13523);
nor U14080 (N_14080,N_13883,N_13888);
and U14081 (N_14081,N_13791,N_13643);
and U14082 (N_14082,N_13536,N_13579);
xor U14083 (N_14083,N_13811,N_13632);
and U14084 (N_14084,N_13803,N_13994);
or U14085 (N_14085,N_13812,N_13909);
and U14086 (N_14086,N_13861,N_13783);
or U14087 (N_14087,N_13834,N_13937);
or U14088 (N_14088,N_13507,N_13518);
xnor U14089 (N_14089,N_13699,N_13514);
or U14090 (N_14090,N_13901,N_13845);
xnor U14091 (N_14091,N_13979,N_13750);
nor U14092 (N_14092,N_13900,N_13533);
nor U14093 (N_14093,N_13526,N_13720);
or U14094 (N_14094,N_13957,N_13968);
and U14095 (N_14095,N_13728,N_13858);
or U14096 (N_14096,N_13781,N_13640);
or U14097 (N_14097,N_13576,N_13718);
and U14098 (N_14098,N_13794,N_13825);
or U14099 (N_14099,N_13521,N_13734);
or U14100 (N_14100,N_13776,N_13618);
xor U14101 (N_14101,N_13826,N_13617);
nor U14102 (N_14102,N_13724,N_13552);
and U14103 (N_14103,N_13642,N_13969);
nand U14104 (N_14104,N_13773,N_13871);
or U14105 (N_14105,N_13588,N_13547);
nor U14106 (N_14106,N_13603,N_13772);
and U14107 (N_14107,N_13884,N_13786);
nor U14108 (N_14108,N_13765,N_13609);
or U14109 (N_14109,N_13762,N_13666);
and U14110 (N_14110,N_13778,N_13539);
nand U14111 (N_14111,N_13653,N_13512);
nand U14112 (N_14112,N_13954,N_13975);
and U14113 (N_14113,N_13938,N_13853);
nor U14114 (N_14114,N_13947,N_13601);
and U14115 (N_14115,N_13922,N_13974);
nor U14116 (N_14116,N_13959,N_13662);
nand U14117 (N_14117,N_13631,N_13624);
or U14118 (N_14118,N_13997,N_13983);
nand U14119 (N_14119,N_13722,N_13550);
nand U14120 (N_14120,N_13541,N_13727);
nor U14121 (N_14121,N_13698,N_13961);
nand U14122 (N_14122,N_13701,N_13889);
nor U14123 (N_14123,N_13792,N_13556);
nor U14124 (N_14124,N_13515,N_13513);
or U14125 (N_14125,N_13821,N_13940);
or U14126 (N_14126,N_13849,N_13885);
and U14127 (N_14127,N_13535,N_13501);
or U14128 (N_14128,N_13876,N_13748);
xor U14129 (N_14129,N_13591,N_13530);
nand U14130 (N_14130,N_13584,N_13870);
nor U14131 (N_14131,N_13865,N_13565);
nand U14132 (N_14132,N_13976,N_13593);
or U14133 (N_14133,N_13608,N_13638);
nand U14134 (N_14134,N_13835,N_13679);
xor U14135 (N_14135,N_13573,N_13897);
nor U14136 (N_14136,N_13681,N_13659);
or U14137 (N_14137,N_13531,N_13597);
xnor U14138 (N_14138,N_13875,N_13929);
nand U14139 (N_14139,N_13908,N_13690);
or U14140 (N_14140,N_13801,N_13933);
nor U14141 (N_14141,N_13763,N_13673);
or U14142 (N_14142,N_13878,N_13869);
nor U14143 (N_14143,N_13910,N_13676);
xor U14144 (N_14144,N_13543,N_13726);
xnor U14145 (N_14145,N_13656,N_13946);
and U14146 (N_14146,N_13779,N_13738);
nand U14147 (N_14147,N_13721,N_13939);
nand U14148 (N_14148,N_13607,N_13658);
nor U14149 (N_14149,N_13648,N_13647);
or U14150 (N_14150,N_13682,N_13509);
and U14151 (N_14151,N_13866,N_13637);
nor U14152 (N_14152,N_13604,N_13600);
nand U14153 (N_14153,N_13639,N_13751);
and U14154 (N_14154,N_13911,N_13664);
or U14155 (N_14155,N_13611,N_13960);
and U14156 (N_14156,N_13824,N_13660);
xnor U14157 (N_14157,N_13819,N_13978);
or U14158 (N_14158,N_13741,N_13758);
or U14159 (N_14159,N_13764,N_13623);
nand U14160 (N_14160,N_13898,N_13695);
and U14161 (N_14161,N_13895,N_13952);
and U14162 (N_14162,N_13777,N_13990);
and U14163 (N_14163,N_13563,N_13705);
nand U14164 (N_14164,N_13628,N_13985);
nor U14165 (N_14165,N_13935,N_13830);
and U14166 (N_14166,N_13636,N_13920);
xor U14167 (N_14167,N_13840,N_13522);
and U14168 (N_14168,N_13554,N_13912);
and U14169 (N_14169,N_13879,N_13691);
nor U14170 (N_14170,N_13973,N_13677);
nand U14171 (N_14171,N_13544,N_13737);
nand U14172 (N_14172,N_13822,N_13948);
xor U14173 (N_14173,N_13907,N_13672);
and U14174 (N_14174,N_13784,N_13916);
and U14175 (N_14175,N_13561,N_13872);
and U14176 (N_14176,N_13944,N_13802);
and U14177 (N_14177,N_13704,N_13592);
nand U14178 (N_14178,N_13805,N_13931);
nor U14179 (N_14179,N_13529,N_13500);
or U14180 (N_14180,N_13982,N_13708);
or U14181 (N_14181,N_13992,N_13629);
nand U14182 (N_14182,N_13757,N_13951);
and U14183 (N_14183,N_13596,N_13972);
nor U14184 (N_14184,N_13893,N_13668);
and U14185 (N_14185,N_13590,N_13904);
or U14186 (N_14186,N_13671,N_13941);
nand U14187 (N_14187,N_13716,N_13574);
nand U14188 (N_14188,N_13649,N_13971);
and U14189 (N_14189,N_13928,N_13693);
nor U14190 (N_14190,N_13516,N_13572);
and U14191 (N_14191,N_13553,N_13520);
nand U14192 (N_14192,N_13557,N_13918);
nor U14193 (N_14193,N_13913,N_13886);
xor U14194 (N_14194,N_13877,N_13620);
xor U14195 (N_14195,N_13711,N_13540);
nand U14196 (N_14196,N_13546,N_13815);
xnor U14197 (N_14197,N_13817,N_13742);
nand U14198 (N_14198,N_13569,N_13641);
and U14199 (N_14199,N_13934,N_13782);
nand U14200 (N_14200,N_13848,N_13760);
and U14201 (N_14201,N_13752,N_13635);
nor U14202 (N_14202,N_13851,N_13685);
xnor U14203 (N_14203,N_13545,N_13712);
or U14204 (N_14204,N_13925,N_13602);
nand U14205 (N_14205,N_13882,N_13905);
nor U14206 (N_14206,N_13958,N_13674);
nand U14207 (N_14207,N_13843,N_13914);
nand U14208 (N_14208,N_13578,N_13595);
nor U14209 (N_14209,N_13622,N_13980);
nor U14210 (N_14210,N_13844,N_13808);
and U14211 (N_14211,N_13739,N_13797);
and U14212 (N_14212,N_13896,N_13768);
xor U14213 (N_14213,N_13689,N_13645);
and U14214 (N_14214,N_13926,N_13559);
xnor U14215 (N_14215,N_13517,N_13832);
nor U14216 (N_14216,N_13785,N_13717);
nand U14217 (N_14217,N_13862,N_13989);
and U14218 (N_14218,N_13846,N_13863);
or U14219 (N_14219,N_13683,N_13599);
nor U14220 (N_14220,N_13542,N_13856);
nor U14221 (N_14221,N_13806,N_13873);
xnor U14222 (N_14222,N_13586,N_13902);
xor U14223 (N_14223,N_13696,N_13663);
and U14224 (N_14224,N_13675,N_13616);
or U14225 (N_14225,N_13511,N_13894);
nor U14226 (N_14226,N_13589,N_13594);
nand U14227 (N_14227,N_13813,N_13735);
or U14228 (N_14228,N_13746,N_13963);
xnor U14229 (N_14229,N_13669,N_13652);
nand U14230 (N_14230,N_13627,N_13807);
nor U14231 (N_14231,N_13881,N_13874);
nand U14232 (N_14232,N_13715,N_13694);
nand U14233 (N_14233,N_13740,N_13868);
or U14234 (N_14234,N_13713,N_13798);
xor U14235 (N_14235,N_13665,N_13823);
or U14236 (N_14236,N_13855,N_13587);
or U14237 (N_14237,N_13923,N_13580);
nand U14238 (N_14238,N_13626,N_13828);
or U14239 (N_14239,N_13610,N_13995);
xor U14240 (N_14240,N_13538,N_13743);
or U14241 (N_14241,N_13818,N_13753);
nor U14242 (N_14242,N_13930,N_13614);
nand U14243 (N_14243,N_13857,N_13633);
and U14244 (N_14244,N_13998,N_13919);
nor U14245 (N_14245,N_13850,N_13966);
and U14246 (N_14246,N_13945,N_13688);
and U14247 (N_14247,N_13790,N_13502);
nand U14248 (N_14248,N_13736,N_13558);
and U14249 (N_14249,N_13697,N_13847);
or U14250 (N_14250,N_13823,N_13730);
nor U14251 (N_14251,N_13506,N_13863);
or U14252 (N_14252,N_13586,N_13569);
or U14253 (N_14253,N_13887,N_13559);
nor U14254 (N_14254,N_13522,N_13964);
or U14255 (N_14255,N_13889,N_13594);
and U14256 (N_14256,N_13633,N_13945);
xor U14257 (N_14257,N_13962,N_13698);
and U14258 (N_14258,N_13514,N_13510);
nand U14259 (N_14259,N_13687,N_13748);
or U14260 (N_14260,N_13508,N_13777);
nand U14261 (N_14261,N_13689,N_13615);
nand U14262 (N_14262,N_13866,N_13676);
or U14263 (N_14263,N_13737,N_13724);
and U14264 (N_14264,N_13555,N_13561);
or U14265 (N_14265,N_13890,N_13650);
and U14266 (N_14266,N_13984,N_13695);
xnor U14267 (N_14267,N_13889,N_13685);
nand U14268 (N_14268,N_13858,N_13661);
nand U14269 (N_14269,N_13761,N_13639);
and U14270 (N_14270,N_13501,N_13729);
or U14271 (N_14271,N_13889,N_13525);
nand U14272 (N_14272,N_13941,N_13502);
xor U14273 (N_14273,N_13873,N_13747);
nand U14274 (N_14274,N_13521,N_13777);
nor U14275 (N_14275,N_13605,N_13842);
nor U14276 (N_14276,N_13711,N_13769);
nor U14277 (N_14277,N_13795,N_13554);
nand U14278 (N_14278,N_13857,N_13517);
nor U14279 (N_14279,N_13565,N_13554);
and U14280 (N_14280,N_13523,N_13587);
nor U14281 (N_14281,N_13999,N_13898);
and U14282 (N_14282,N_13591,N_13625);
nand U14283 (N_14283,N_13527,N_13690);
xor U14284 (N_14284,N_13776,N_13553);
and U14285 (N_14285,N_13660,N_13966);
and U14286 (N_14286,N_13520,N_13847);
and U14287 (N_14287,N_13739,N_13719);
nand U14288 (N_14288,N_13597,N_13741);
nand U14289 (N_14289,N_13679,N_13929);
nand U14290 (N_14290,N_13603,N_13791);
nor U14291 (N_14291,N_13529,N_13558);
and U14292 (N_14292,N_13528,N_13680);
nand U14293 (N_14293,N_13586,N_13511);
or U14294 (N_14294,N_13580,N_13823);
and U14295 (N_14295,N_13844,N_13980);
xor U14296 (N_14296,N_13625,N_13812);
nand U14297 (N_14297,N_13869,N_13689);
nor U14298 (N_14298,N_13504,N_13666);
and U14299 (N_14299,N_13884,N_13823);
or U14300 (N_14300,N_13814,N_13584);
nor U14301 (N_14301,N_13708,N_13743);
xnor U14302 (N_14302,N_13971,N_13656);
nor U14303 (N_14303,N_13836,N_13683);
and U14304 (N_14304,N_13764,N_13608);
xnor U14305 (N_14305,N_13878,N_13552);
nand U14306 (N_14306,N_13708,N_13552);
nand U14307 (N_14307,N_13891,N_13786);
and U14308 (N_14308,N_13714,N_13803);
nand U14309 (N_14309,N_13604,N_13776);
or U14310 (N_14310,N_13547,N_13630);
nand U14311 (N_14311,N_13816,N_13864);
nor U14312 (N_14312,N_13537,N_13956);
nand U14313 (N_14313,N_13776,N_13866);
and U14314 (N_14314,N_13704,N_13974);
nor U14315 (N_14315,N_13519,N_13864);
or U14316 (N_14316,N_13828,N_13677);
or U14317 (N_14317,N_13951,N_13654);
and U14318 (N_14318,N_13691,N_13788);
or U14319 (N_14319,N_13610,N_13766);
nor U14320 (N_14320,N_13821,N_13977);
nand U14321 (N_14321,N_13616,N_13591);
nor U14322 (N_14322,N_13750,N_13764);
and U14323 (N_14323,N_13773,N_13599);
nor U14324 (N_14324,N_13705,N_13886);
nand U14325 (N_14325,N_13866,N_13982);
nor U14326 (N_14326,N_13813,N_13907);
xor U14327 (N_14327,N_13603,N_13812);
or U14328 (N_14328,N_13553,N_13819);
nor U14329 (N_14329,N_13557,N_13749);
or U14330 (N_14330,N_13664,N_13728);
nand U14331 (N_14331,N_13557,N_13596);
and U14332 (N_14332,N_13979,N_13510);
or U14333 (N_14333,N_13796,N_13695);
nor U14334 (N_14334,N_13780,N_13894);
xnor U14335 (N_14335,N_13594,N_13803);
nor U14336 (N_14336,N_13989,N_13718);
and U14337 (N_14337,N_13923,N_13507);
and U14338 (N_14338,N_13568,N_13674);
nand U14339 (N_14339,N_13711,N_13762);
xor U14340 (N_14340,N_13658,N_13695);
and U14341 (N_14341,N_13532,N_13613);
and U14342 (N_14342,N_13600,N_13658);
xnor U14343 (N_14343,N_13917,N_13770);
and U14344 (N_14344,N_13782,N_13814);
nor U14345 (N_14345,N_13507,N_13598);
or U14346 (N_14346,N_13584,N_13763);
nand U14347 (N_14347,N_13912,N_13923);
or U14348 (N_14348,N_13542,N_13910);
or U14349 (N_14349,N_13635,N_13565);
or U14350 (N_14350,N_13696,N_13973);
or U14351 (N_14351,N_13897,N_13878);
nand U14352 (N_14352,N_13530,N_13631);
and U14353 (N_14353,N_13759,N_13536);
and U14354 (N_14354,N_13580,N_13742);
or U14355 (N_14355,N_13779,N_13829);
or U14356 (N_14356,N_13758,N_13781);
nor U14357 (N_14357,N_13919,N_13719);
nor U14358 (N_14358,N_13542,N_13888);
or U14359 (N_14359,N_13993,N_13913);
nand U14360 (N_14360,N_13576,N_13748);
or U14361 (N_14361,N_13535,N_13982);
or U14362 (N_14362,N_13912,N_13510);
nor U14363 (N_14363,N_13509,N_13801);
nor U14364 (N_14364,N_13967,N_13888);
or U14365 (N_14365,N_13855,N_13939);
and U14366 (N_14366,N_13940,N_13842);
or U14367 (N_14367,N_13648,N_13563);
xnor U14368 (N_14368,N_13967,N_13935);
and U14369 (N_14369,N_13961,N_13868);
and U14370 (N_14370,N_13884,N_13529);
nand U14371 (N_14371,N_13978,N_13998);
and U14372 (N_14372,N_13508,N_13846);
or U14373 (N_14373,N_13614,N_13873);
nor U14374 (N_14374,N_13588,N_13907);
nand U14375 (N_14375,N_13662,N_13880);
and U14376 (N_14376,N_13803,N_13837);
or U14377 (N_14377,N_13542,N_13595);
and U14378 (N_14378,N_13807,N_13958);
or U14379 (N_14379,N_13753,N_13604);
or U14380 (N_14380,N_13937,N_13607);
or U14381 (N_14381,N_13640,N_13962);
nor U14382 (N_14382,N_13560,N_13719);
or U14383 (N_14383,N_13677,N_13781);
and U14384 (N_14384,N_13735,N_13957);
nand U14385 (N_14385,N_13779,N_13884);
or U14386 (N_14386,N_13706,N_13639);
or U14387 (N_14387,N_13957,N_13612);
or U14388 (N_14388,N_13732,N_13822);
and U14389 (N_14389,N_13536,N_13570);
xor U14390 (N_14390,N_13671,N_13768);
xor U14391 (N_14391,N_13911,N_13636);
nand U14392 (N_14392,N_13845,N_13690);
and U14393 (N_14393,N_13644,N_13699);
and U14394 (N_14394,N_13612,N_13545);
nand U14395 (N_14395,N_13963,N_13553);
nand U14396 (N_14396,N_13892,N_13796);
nor U14397 (N_14397,N_13631,N_13840);
or U14398 (N_14398,N_13577,N_13705);
nand U14399 (N_14399,N_13990,N_13787);
nor U14400 (N_14400,N_13902,N_13814);
and U14401 (N_14401,N_13814,N_13847);
or U14402 (N_14402,N_13808,N_13690);
or U14403 (N_14403,N_13985,N_13521);
and U14404 (N_14404,N_13965,N_13928);
and U14405 (N_14405,N_13810,N_13807);
nand U14406 (N_14406,N_13576,N_13612);
xnor U14407 (N_14407,N_13744,N_13664);
nand U14408 (N_14408,N_13802,N_13801);
or U14409 (N_14409,N_13750,N_13926);
nand U14410 (N_14410,N_13839,N_13914);
nor U14411 (N_14411,N_13929,N_13819);
and U14412 (N_14412,N_13901,N_13809);
or U14413 (N_14413,N_13756,N_13856);
nor U14414 (N_14414,N_13962,N_13882);
or U14415 (N_14415,N_13615,N_13882);
or U14416 (N_14416,N_13542,N_13737);
xnor U14417 (N_14417,N_13575,N_13735);
and U14418 (N_14418,N_13906,N_13648);
or U14419 (N_14419,N_13724,N_13505);
nand U14420 (N_14420,N_13808,N_13698);
nand U14421 (N_14421,N_13870,N_13958);
nor U14422 (N_14422,N_13792,N_13699);
and U14423 (N_14423,N_13765,N_13760);
nand U14424 (N_14424,N_13716,N_13818);
xnor U14425 (N_14425,N_13837,N_13963);
nand U14426 (N_14426,N_13833,N_13974);
nand U14427 (N_14427,N_13819,N_13630);
xor U14428 (N_14428,N_13621,N_13553);
nor U14429 (N_14429,N_13987,N_13870);
nand U14430 (N_14430,N_13632,N_13521);
nand U14431 (N_14431,N_13566,N_13806);
xnor U14432 (N_14432,N_13502,N_13513);
or U14433 (N_14433,N_13758,N_13784);
xnor U14434 (N_14434,N_13640,N_13692);
nand U14435 (N_14435,N_13772,N_13694);
and U14436 (N_14436,N_13952,N_13786);
and U14437 (N_14437,N_13675,N_13690);
xnor U14438 (N_14438,N_13779,N_13530);
nor U14439 (N_14439,N_13881,N_13639);
nor U14440 (N_14440,N_13918,N_13748);
and U14441 (N_14441,N_13857,N_13731);
nor U14442 (N_14442,N_13859,N_13649);
and U14443 (N_14443,N_13918,N_13986);
and U14444 (N_14444,N_13966,N_13811);
nand U14445 (N_14445,N_13968,N_13555);
nand U14446 (N_14446,N_13941,N_13884);
nor U14447 (N_14447,N_13978,N_13632);
or U14448 (N_14448,N_13651,N_13832);
nand U14449 (N_14449,N_13520,N_13973);
nand U14450 (N_14450,N_13509,N_13829);
xnor U14451 (N_14451,N_13577,N_13779);
xnor U14452 (N_14452,N_13521,N_13806);
or U14453 (N_14453,N_13723,N_13783);
nor U14454 (N_14454,N_13951,N_13815);
nor U14455 (N_14455,N_13505,N_13767);
nor U14456 (N_14456,N_13541,N_13540);
or U14457 (N_14457,N_13745,N_13526);
or U14458 (N_14458,N_13623,N_13763);
and U14459 (N_14459,N_13861,N_13651);
nand U14460 (N_14460,N_13520,N_13641);
or U14461 (N_14461,N_13510,N_13580);
xnor U14462 (N_14462,N_13978,N_13788);
nand U14463 (N_14463,N_13761,N_13903);
nor U14464 (N_14464,N_13927,N_13714);
nand U14465 (N_14465,N_13666,N_13657);
xor U14466 (N_14466,N_13908,N_13680);
or U14467 (N_14467,N_13562,N_13823);
xnor U14468 (N_14468,N_13635,N_13507);
xnor U14469 (N_14469,N_13996,N_13549);
and U14470 (N_14470,N_13607,N_13814);
or U14471 (N_14471,N_13967,N_13998);
or U14472 (N_14472,N_13698,N_13958);
or U14473 (N_14473,N_13571,N_13762);
and U14474 (N_14474,N_13938,N_13554);
nor U14475 (N_14475,N_13741,N_13574);
and U14476 (N_14476,N_13886,N_13955);
nor U14477 (N_14477,N_13848,N_13770);
and U14478 (N_14478,N_13808,N_13668);
or U14479 (N_14479,N_13691,N_13750);
nor U14480 (N_14480,N_13981,N_13881);
and U14481 (N_14481,N_13509,N_13727);
nor U14482 (N_14482,N_13793,N_13541);
nand U14483 (N_14483,N_13647,N_13709);
or U14484 (N_14484,N_13855,N_13551);
nand U14485 (N_14485,N_13848,N_13816);
and U14486 (N_14486,N_13851,N_13882);
or U14487 (N_14487,N_13634,N_13866);
or U14488 (N_14488,N_13927,N_13991);
nand U14489 (N_14489,N_13816,N_13817);
nor U14490 (N_14490,N_13592,N_13710);
and U14491 (N_14491,N_13759,N_13867);
nand U14492 (N_14492,N_13736,N_13772);
or U14493 (N_14493,N_13705,N_13755);
nand U14494 (N_14494,N_13876,N_13950);
or U14495 (N_14495,N_13624,N_13873);
or U14496 (N_14496,N_13557,N_13964);
nand U14497 (N_14497,N_13673,N_13788);
nor U14498 (N_14498,N_13664,N_13733);
nand U14499 (N_14499,N_13973,N_13572);
and U14500 (N_14500,N_14494,N_14033);
nand U14501 (N_14501,N_14136,N_14249);
or U14502 (N_14502,N_14004,N_14142);
nor U14503 (N_14503,N_14200,N_14143);
or U14504 (N_14504,N_14066,N_14371);
or U14505 (N_14505,N_14123,N_14068);
xor U14506 (N_14506,N_14338,N_14348);
nor U14507 (N_14507,N_14165,N_14190);
nor U14508 (N_14508,N_14141,N_14070);
and U14509 (N_14509,N_14458,N_14427);
xnor U14510 (N_14510,N_14057,N_14048);
or U14511 (N_14511,N_14281,N_14199);
nand U14512 (N_14512,N_14075,N_14009);
or U14513 (N_14513,N_14417,N_14430);
nor U14514 (N_14514,N_14031,N_14162);
nand U14515 (N_14515,N_14416,N_14337);
xor U14516 (N_14516,N_14381,N_14473);
nand U14517 (N_14517,N_14446,N_14362);
nor U14518 (N_14518,N_14243,N_14469);
nand U14519 (N_14519,N_14299,N_14477);
xnor U14520 (N_14520,N_14399,N_14104);
nand U14521 (N_14521,N_14139,N_14134);
nand U14522 (N_14522,N_14278,N_14043);
or U14523 (N_14523,N_14151,N_14122);
or U14524 (N_14524,N_14431,N_14255);
xnor U14525 (N_14525,N_14270,N_14313);
nand U14526 (N_14526,N_14246,N_14219);
nor U14527 (N_14527,N_14392,N_14476);
xnor U14528 (N_14528,N_14091,N_14160);
nand U14529 (N_14529,N_14305,N_14466);
nand U14530 (N_14530,N_14340,N_14126);
nand U14531 (N_14531,N_14154,N_14051);
or U14532 (N_14532,N_14029,N_14413);
nand U14533 (N_14533,N_14288,N_14342);
xnor U14534 (N_14534,N_14148,N_14410);
or U14535 (N_14535,N_14149,N_14214);
or U14536 (N_14536,N_14412,N_14448);
and U14537 (N_14537,N_14077,N_14235);
and U14538 (N_14538,N_14450,N_14156);
nand U14539 (N_14539,N_14183,N_14307);
nor U14540 (N_14540,N_14047,N_14432);
xor U14541 (N_14541,N_14326,N_14181);
and U14542 (N_14542,N_14359,N_14178);
nand U14543 (N_14543,N_14279,N_14024);
and U14544 (N_14544,N_14087,N_14333);
nor U14545 (N_14545,N_14022,N_14481);
nor U14546 (N_14546,N_14056,N_14407);
and U14547 (N_14547,N_14483,N_14101);
nand U14548 (N_14548,N_14370,N_14394);
and U14549 (N_14549,N_14295,N_14163);
and U14550 (N_14550,N_14130,N_14028);
nor U14551 (N_14551,N_14328,N_14109);
nand U14552 (N_14552,N_14010,N_14213);
nand U14553 (N_14553,N_14236,N_14291);
or U14554 (N_14554,N_14275,N_14310);
or U14555 (N_14555,N_14258,N_14452);
nand U14556 (N_14556,N_14069,N_14019);
and U14557 (N_14557,N_14368,N_14099);
or U14558 (N_14558,N_14485,N_14231);
xnor U14559 (N_14559,N_14088,N_14300);
nor U14560 (N_14560,N_14095,N_14084);
or U14561 (N_14561,N_14355,N_14217);
or U14562 (N_14562,N_14127,N_14499);
or U14563 (N_14563,N_14286,N_14119);
nand U14564 (N_14564,N_14072,N_14212);
nand U14565 (N_14565,N_14405,N_14277);
xnor U14566 (N_14566,N_14497,N_14115);
xor U14567 (N_14567,N_14132,N_14110);
and U14568 (N_14568,N_14321,N_14262);
or U14569 (N_14569,N_14414,N_14331);
xor U14570 (N_14570,N_14191,N_14210);
nor U14571 (N_14571,N_14346,N_14196);
and U14572 (N_14572,N_14011,N_14422);
xor U14573 (N_14573,N_14224,N_14030);
nor U14574 (N_14574,N_14059,N_14350);
xor U14575 (N_14575,N_14389,N_14460);
and U14576 (N_14576,N_14425,N_14013);
nand U14577 (N_14577,N_14456,N_14420);
and U14578 (N_14578,N_14007,N_14027);
or U14579 (N_14579,N_14147,N_14225);
nand U14580 (N_14580,N_14471,N_14146);
and U14581 (N_14581,N_14474,N_14001);
nor U14582 (N_14582,N_14478,N_14040);
and U14583 (N_14583,N_14369,N_14245);
nand U14584 (N_14584,N_14250,N_14000);
or U14585 (N_14585,N_14092,N_14206);
nand U14586 (N_14586,N_14211,N_14254);
or U14587 (N_14587,N_14222,N_14419);
or U14588 (N_14588,N_14021,N_14322);
or U14589 (N_14589,N_14005,N_14131);
nand U14590 (N_14590,N_14232,N_14408);
and U14591 (N_14591,N_14071,N_14363);
nor U14592 (N_14592,N_14145,N_14032);
nor U14593 (N_14593,N_14423,N_14315);
nand U14594 (N_14594,N_14128,N_14185);
nor U14595 (N_14595,N_14108,N_14182);
nor U14596 (N_14596,N_14044,N_14223);
or U14597 (N_14597,N_14402,N_14179);
or U14598 (N_14598,N_14144,N_14496);
nor U14599 (N_14599,N_14100,N_14433);
nand U14600 (N_14600,N_14424,N_14118);
nand U14601 (N_14601,N_14393,N_14140);
nand U14602 (N_14602,N_14221,N_14050);
nor U14603 (N_14603,N_14455,N_14294);
or U14604 (N_14604,N_14352,N_14129);
nor U14605 (N_14605,N_14272,N_14229);
or U14606 (N_14606,N_14449,N_14105);
and U14607 (N_14607,N_14388,N_14240);
and U14608 (N_14608,N_14153,N_14386);
and U14609 (N_14609,N_14360,N_14264);
nor U14610 (N_14610,N_14035,N_14492);
nor U14611 (N_14611,N_14269,N_14319);
nor U14612 (N_14612,N_14170,N_14470);
nand U14613 (N_14613,N_14227,N_14353);
nor U14614 (N_14614,N_14308,N_14230);
nor U14615 (N_14615,N_14008,N_14445);
nand U14616 (N_14616,N_14252,N_14113);
and U14617 (N_14617,N_14261,N_14111);
nor U14618 (N_14618,N_14081,N_14395);
xor U14619 (N_14619,N_14318,N_14304);
or U14620 (N_14620,N_14336,N_14239);
xor U14621 (N_14621,N_14054,N_14094);
and U14622 (N_14622,N_14042,N_14398);
or U14623 (N_14623,N_14330,N_14023);
nor U14624 (N_14624,N_14403,N_14058);
nand U14625 (N_14625,N_14486,N_14133);
nand U14626 (N_14626,N_14265,N_14158);
nor U14627 (N_14627,N_14292,N_14479);
nand U14628 (N_14628,N_14314,N_14285);
xnor U14629 (N_14629,N_14434,N_14465);
and U14630 (N_14630,N_14186,N_14276);
nand U14631 (N_14631,N_14096,N_14303);
or U14632 (N_14632,N_14312,N_14107);
nand U14633 (N_14633,N_14463,N_14203);
nor U14634 (N_14634,N_14037,N_14396);
xnor U14635 (N_14635,N_14406,N_14480);
or U14636 (N_14636,N_14390,N_14184);
and U14637 (N_14637,N_14475,N_14055);
nand U14638 (N_14638,N_14358,N_14038);
and U14639 (N_14639,N_14161,N_14046);
nor U14640 (N_14640,N_14085,N_14493);
nand U14641 (N_14641,N_14124,N_14379);
or U14642 (N_14642,N_14382,N_14006);
nand U14643 (N_14643,N_14188,N_14332);
nand U14644 (N_14644,N_14220,N_14168);
nand U14645 (N_14645,N_14025,N_14065);
or U14646 (N_14646,N_14484,N_14383);
and U14647 (N_14647,N_14063,N_14429);
nor U14648 (N_14648,N_14459,N_14097);
nor U14649 (N_14649,N_14385,N_14339);
or U14650 (N_14650,N_14437,N_14067);
xor U14651 (N_14651,N_14334,N_14045);
or U14652 (N_14652,N_14343,N_14082);
nand U14653 (N_14653,N_14472,N_14026);
or U14654 (N_14654,N_14377,N_14282);
xnor U14655 (N_14655,N_14172,N_14189);
nand U14656 (N_14656,N_14017,N_14194);
and U14657 (N_14657,N_14093,N_14457);
nand U14658 (N_14658,N_14039,N_14137);
nand U14659 (N_14659,N_14159,N_14349);
and U14660 (N_14660,N_14102,N_14441);
or U14661 (N_14661,N_14274,N_14323);
nor U14662 (N_14662,N_14138,N_14444);
and U14663 (N_14663,N_14268,N_14074);
nor U14664 (N_14664,N_14014,N_14073);
nor U14665 (N_14665,N_14438,N_14418);
nor U14666 (N_14666,N_14062,N_14461);
nor U14667 (N_14667,N_14209,N_14283);
or U14668 (N_14668,N_14193,N_14256);
or U14669 (N_14669,N_14378,N_14311);
nor U14670 (N_14670,N_14233,N_14451);
nor U14671 (N_14671,N_14155,N_14324);
nor U14672 (N_14672,N_14290,N_14228);
nand U14673 (N_14673,N_14157,N_14078);
nand U14674 (N_14674,N_14114,N_14079);
or U14675 (N_14675,N_14491,N_14301);
xnor U14676 (N_14676,N_14041,N_14356);
and U14677 (N_14677,N_14380,N_14273);
xnor U14678 (N_14678,N_14176,N_14247);
or U14679 (N_14679,N_14052,N_14173);
nand U14680 (N_14680,N_14207,N_14175);
and U14681 (N_14681,N_14327,N_14267);
nor U14682 (N_14682,N_14482,N_14428);
and U14683 (N_14683,N_14204,N_14192);
or U14684 (N_14684,N_14218,N_14316);
and U14685 (N_14685,N_14121,N_14280);
xor U14686 (N_14686,N_14036,N_14354);
or U14687 (N_14687,N_14366,N_14345);
nand U14688 (N_14688,N_14060,N_14198);
and U14689 (N_14689,N_14177,N_14226);
and U14690 (N_14690,N_14016,N_14384);
nand U14691 (N_14691,N_14495,N_14364);
and U14692 (N_14692,N_14015,N_14376);
or U14693 (N_14693,N_14297,N_14090);
nand U14694 (N_14694,N_14341,N_14329);
nor U14695 (N_14695,N_14248,N_14253);
and U14696 (N_14696,N_14053,N_14464);
nor U14697 (N_14697,N_14309,N_14241);
nor U14698 (N_14698,N_14487,N_14086);
nand U14699 (N_14699,N_14259,N_14488);
or U14700 (N_14700,N_14397,N_14365);
nor U14701 (N_14701,N_14317,N_14490);
and U14702 (N_14702,N_14169,N_14400);
and U14703 (N_14703,N_14298,N_14012);
nor U14704 (N_14704,N_14293,N_14083);
nor U14705 (N_14705,N_14171,N_14462);
nor U14706 (N_14706,N_14103,N_14263);
nor U14707 (N_14707,N_14372,N_14061);
or U14708 (N_14708,N_14447,N_14443);
nor U14709 (N_14709,N_14251,N_14296);
or U14710 (N_14710,N_14034,N_14440);
nand U14711 (N_14711,N_14435,N_14106);
or U14712 (N_14712,N_14208,N_14335);
and U14713 (N_14713,N_14215,N_14266);
and U14714 (N_14714,N_14387,N_14197);
nor U14715 (N_14715,N_14152,N_14174);
xnor U14716 (N_14716,N_14271,N_14367);
and U14717 (N_14717,N_14202,N_14257);
nand U14718 (N_14718,N_14002,N_14467);
and U14719 (N_14719,N_14180,N_14325);
and U14720 (N_14720,N_14421,N_14411);
and U14721 (N_14721,N_14426,N_14409);
nor U14722 (N_14722,N_14351,N_14076);
nand U14723 (N_14723,N_14167,N_14391);
xor U14724 (N_14724,N_14089,N_14344);
nand U14725 (N_14725,N_14195,N_14242);
and U14726 (N_14726,N_14238,N_14453);
and U14727 (N_14727,N_14361,N_14404);
and U14728 (N_14728,N_14375,N_14498);
or U14729 (N_14729,N_14320,N_14187);
and U14730 (N_14730,N_14287,N_14442);
nand U14731 (N_14731,N_14150,N_14436);
or U14732 (N_14732,N_14260,N_14125);
xor U14733 (N_14733,N_14166,N_14357);
and U14734 (N_14734,N_14120,N_14164);
xnor U14735 (N_14735,N_14302,N_14454);
nor U14736 (N_14736,N_14116,N_14374);
and U14737 (N_14737,N_14205,N_14112);
nor U14738 (N_14738,N_14117,N_14098);
xor U14739 (N_14739,N_14003,N_14244);
or U14740 (N_14740,N_14049,N_14080);
and U14741 (N_14741,N_14289,N_14306);
and U14742 (N_14742,N_14234,N_14415);
xor U14743 (N_14743,N_14216,N_14284);
nor U14744 (N_14744,N_14064,N_14489);
nor U14745 (N_14745,N_14020,N_14018);
nand U14746 (N_14746,N_14135,N_14347);
xor U14747 (N_14747,N_14439,N_14468);
and U14748 (N_14748,N_14201,N_14237);
xnor U14749 (N_14749,N_14401,N_14373);
and U14750 (N_14750,N_14366,N_14466);
nor U14751 (N_14751,N_14108,N_14146);
nor U14752 (N_14752,N_14375,N_14424);
xor U14753 (N_14753,N_14292,N_14113);
or U14754 (N_14754,N_14274,N_14289);
nand U14755 (N_14755,N_14258,N_14237);
and U14756 (N_14756,N_14371,N_14178);
nand U14757 (N_14757,N_14300,N_14052);
xor U14758 (N_14758,N_14304,N_14459);
xor U14759 (N_14759,N_14330,N_14409);
and U14760 (N_14760,N_14440,N_14023);
and U14761 (N_14761,N_14315,N_14186);
nand U14762 (N_14762,N_14129,N_14493);
xnor U14763 (N_14763,N_14210,N_14288);
or U14764 (N_14764,N_14039,N_14043);
and U14765 (N_14765,N_14218,N_14082);
xnor U14766 (N_14766,N_14259,N_14320);
nor U14767 (N_14767,N_14482,N_14434);
and U14768 (N_14768,N_14268,N_14409);
nand U14769 (N_14769,N_14405,N_14202);
nand U14770 (N_14770,N_14484,N_14224);
and U14771 (N_14771,N_14310,N_14460);
or U14772 (N_14772,N_14007,N_14373);
xor U14773 (N_14773,N_14177,N_14267);
and U14774 (N_14774,N_14325,N_14054);
nand U14775 (N_14775,N_14100,N_14414);
and U14776 (N_14776,N_14192,N_14355);
nand U14777 (N_14777,N_14101,N_14211);
and U14778 (N_14778,N_14040,N_14492);
nand U14779 (N_14779,N_14165,N_14209);
or U14780 (N_14780,N_14131,N_14067);
nand U14781 (N_14781,N_14152,N_14106);
and U14782 (N_14782,N_14218,N_14055);
and U14783 (N_14783,N_14205,N_14275);
and U14784 (N_14784,N_14342,N_14253);
nand U14785 (N_14785,N_14142,N_14421);
or U14786 (N_14786,N_14107,N_14376);
or U14787 (N_14787,N_14403,N_14112);
nor U14788 (N_14788,N_14096,N_14109);
nand U14789 (N_14789,N_14197,N_14213);
xnor U14790 (N_14790,N_14035,N_14268);
and U14791 (N_14791,N_14017,N_14146);
and U14792 (N_14792,N_14295,N_14199);
nor U14793 (N_14793,N_14407,N_14307);
nand U14794 (N_14794,N_14350,N_14369);
nor U14795 (N_14795,N_14237,N_14015);
nor U14796 (N_14796,N_14117,N_14299);
and U14797 (N_14797,N_14364,N_14163);
or U14798 (N_14798,N_14338,N_14373);
or U14799 (N_14799,N_14393,N_14179);
and U14800 (N_14800,N_14364,N_14290);
nor U14801 (N_14801,N_14464,N_14016);
and U14802 (N_14802,N_14182,N_14401);
nor U14803 (N_14803,N_14120,N_14292);
nor U14804 (N_14804,N_14048,N_14101);
xnor U14805 (N_14805,N_14120,N_14316);
or U14806 (N_14806,N_14386,N_14438);
nand U14807 (N_14807,N_14041,N_14159);
nand U14808 (N_14808,N_14010,N_14056);
nand U14809 (N_14809,N_14265,N_14000);
or U14810 (N_14810,N_14473,N_14295);
nor U14811 (N_14811,N_14468,N_14172);
and U14812 (N_14812,N_14307,N_14085);
xor U14813 (N_14813,N_14037,N_14310);
and U14814 (N_14814,N_14065,N_14151);
or U14815 (N_14815,N_14286,N_14393);
nand U14816 (N_14816,N_14450,N_14181);
or U14817 (N_14817,N_14164,N_14481);
nand U14818 (N_14818,N_14316,N_14462);
or U14819 (N_14819,N_14150,N_14030);
and U14820 (N_14820,N_14100,N_14016);
xnor U14821 (N_14821,N_14198,N_14208);
and U14822 (N_14822,N_14180,N_14260);
and U14823 (N_14823,N_14338,N_14061);
nand U14824 (N_14824,N_14094,N_14346);
nand U14825 (N_14825,N_14472,N_14293);
nor U14826 (N_14826,N_14368,N_14430);
or U14827 (N_14827,N_14315,N_14166);
and U14828 (N_14828,N_14308,N_14127);
nor U14829 (N_14829,N_14387,N_14304);
or U14830 (N_14830,N_14058,N_14331);
nand U14831 (N_14831,N_14149,N_14388);
nand U14832 (N_14832,N_14084,N_14479);
and U14833 (N_14833,N_14485,N_14054);
or U14834 (N_14834,N_14405,N_14418);
or U14835 (N_14835,N_14259,N_14423);
and U14836 (N_14836,N_14284,N_14187);
or U14837 (N_14837,N_14245,N_14035);
and U14838 (N_14838,N_14246,N_14346);
and U14839 (N_14839,N_14399,N_14402);
nor U14840 (N_14840,N_14423,N_14464);
nor U14841 (N_14841,N_14279,N_14302);
and U14842 (N_14842,N_14097,N_14383);
nor U14843 (N_14843,N_14036,N_14029);
nand U14844 (N_14844,N_14129,N_14382);
or U14845 (N_14845,N_14297,N_14055);
or U14846 (N_14846,N_14058,N_14336);
xor U14847 (N_14847,N_14098,N_14165);
and U14848 (N_14848,N_14396,N_14218);
or U14849 (N_14849,N_14240,N_14011);
nor U14850 (N_14850,N_14149,N_14197);
or U14851 (N_14851,N_14225,N_14368);
nand U14852 (N_14852,N_14133,N_14023);
and U14853 (N_14853,N_14323,N_14443);
or U14854 (N_14854,N_14011,N_14437);
nand U14855 (N_14855,N_14155,N_14235);
and U14856 (N_14856,N_14370,N_14255);
and U14857 (N_14857,N_14016,N_14015);
and U14858 (N_14858,N_14403,N_14304);
and U14859 (N_14859,N_14180,N_14442);
xnor U14860 (N_14860,N_14408,N_14129);
or U14861 (N_14861,N_14018,N_14179);
nand U14862 (N_14862,N_14048,N_14063);
xnor U14863 (N_14863,N_14011,N_14051);
or U14864 (N_14864,N_14445,N_14016);
or U14865 (N_14865,N_14112,N_14252);
or U14866 (N_14866,N_14411,N_14066);
xor U14867 (N_14867,N_14289,N_14217);
and U14868 (N_14868,N_14060,N_14054);
xnor U14869 (N_14869,N_14327,N_14388);
nor U14870 (N_14870,N_14447,N_14282);
and U14871 (N_14871,N_14170,N_14078);
or U14872 (N_14872,N_14401,N_14414);
nand U14873 (N_14873,N_14429,N_14170);
and U14874 (N_14874,N_14347,N_14418);
xor U14875 (N_14875,N_14275,N_14405);
or U14876 (N_14876,N_14393,N_14097);
or U14877 (N_14877,N_14385,N_14212);
xor U14878 (N_14878,N_14142,N_14140);
nor U14879 (N_14879,N_14203,N_14493);
or U14880 (N_14880,N_14426,N_14198);
xor U14881 (N_14881,N_14205,N_14058);
and U14882 (N_14882,N_14309,N_14493);
or U14883 (N_14883,N_14052,N_14145);
and U14884 (N_14884,N_14128,N_14227);
and U14885 (N_14885,N_14316,N_14183);
or U14886 (N_14886,N_14107,N_14004);
nand U14887 (N_14887,N_14143,N_14314);
and U14888 (N_14888,N_14382,N_14341);
nand U14889 (N_14889,N_14006,N_14316);
nand U14890 (N_14890,N_14448,N_14332);
or U14891 (N_14891,N_14207,N_14379);
nand U14892 (N_14892,N_14437,N_14028);
or U14893 (N_14893,N_14014,N_14364);
nor U14894 (N_14894,N_14030,N_14060);
or U14895 (N_14895,N_14191,N_14168);
nor U14896 (N_14896,N_14173,N_14366);
and U14897 (N_14897,N_14334,N_14048);
and U14898 (N_14898,N_14455,N_14221);
nand U14899 (N_14899,N_14479,N_14155);
xnor U14900 (N_14900,N_14080,N_14315);
and U14901 (N_14901,N_14065,N_14043);
nand U14902 (N_14902,N_14075,N_14416);
xor U14903 (N_14903,N_14424,N_14014);
and U14904 (N_14904,N_14493,N_14378);
nor U14905 (N_14905,N_14047,N_14488);
nand U14906 (N_14906,N_14321,N_14405);
or U14907 (N_14907,N_14035,N_14078);
nor U14908 (N_14908,N_14277,N_14472);
and U14909 (N_14909,N_14246,N_14469);
nand U14910 (N_14910,N_14273,N_14173);
and U14911 (N_14911,N_14305,N_14338);
and U14912 (N_14912,N_14468,N_14476);
or U14913 (N_14913,N_14268,N_14293);
nor U14914 (N_14914,N_14093,N_14277);
xor U14915 (N_14915,N_14174,N_14104);
and U14916 (N_14916,N_14426,N_14174);
nor U14917 (N_14917,N_14429,N_14360);
nand U14918 (N_14918,N_14438,N_14334);
or U14919 (N_14919,N_14170,N_14156);
nor U14920 (N_14920,N_14397,N_14113);
and U14921 (N_14921,N_14355,N_14376);
nor U14922 (N_14922,N_14460,N_14093);
nand U14923 (N_14923,N_14416,N_14318);
nand U14924 (N_14924,N_14337,N_14159);
nand U14925 (N_14925,N_14161,N_14489);
or U14926 (N_14926,N_14180,N_14221);
xnor U14927 (N_14927,N_14448,N_14489);
nor U14928 (N_14928,N_14300,N_14108);
nand U14929 (N_14929,N_14396,N_14140);
xnor U14930 (N_14930,N_14083,N_14052);
or U14931 (N_14931,N_14246,N_14443);
and U14932 (N_14932,N_14398,N_14053);
and U14933 (N_14933,N_14427,N_14316);
nor U14934 (N_14934,N_14360,N_14073);
nor U14935 (N_14935,N_14077,N_14232);
nor U14936 (N_14936,N_14185,N_14493);
and U14937 (N_14937,N_14467,N_14362);
or U14938 (N_14938,N_14480,N_14000);
and U14939 (N_14939,N_14234,N_14159);
or U14940 (N_14940,N_14196,N_14188);
nor U14941 (N_14941,N_14458,N_14373);
nand U14942 (N_14942,N_14033,N_14286);
and U14943 (N_14943,N_14252,N_14195);
nor U14944 (N_14944,N_14361,N_14058);
and U14945 (N_14945,N_14011,N_14176);
and U14946 (N_14946,N_14216,N_14310);
or U14947 (N_14947,N_14190,N_14076);
nor U14948 (N_14948,N_14298,N_14060);
nand U14949 (N_14949,N_14074,N_14466);
and U14950 (N_14950,N_14340,N_14497);
or U14951 (N_14951,N_14355,N_14374);
xnor U14952 (N_14952,N_14267,N_14297);
or U14953 (N_14953,N_14102,N_14490);
and U14954 (N_14954,N_14312,N_14313);
and U14955 (N_14955,N_14370,N_14101);
nand U14956 (N_14956,N_14188,N_14144);
nand U14957 (N_14957,N_14055,N_14458);
xor U14958 (N_14958,N_14286,N_14292);
and U14959 (N_14959,N_14463,N_14207);
nor U14960 (N_14960,N_14394,N_14016);
and U14961 (N_14961,N_14037,N_14226);
or U14962 (N_14962,N_14485,N_14435);
and U14963 (N_14963,N_14494,N_14066);
and U14964 (N_14964,N_14017,N_14400);
nand U14965 (N_14965,N_14363,N_14437);
and U14966 (N_14966,N_14011,N_14173);
nor U14967 (N_14967,N_14173,N_14068);
nor U14968 (N_14968,N_14155,N_14256);
xnor U14969 (N_14969,N_14173,N_14072);
nand U14970 (N_14970,N_14336,N_14341);
nor U14971 (N_14971,N_14123,N_14342);
or U14972 (N_14972,N_14290,N_14156);
xor U14973 (N_14973,N_14029,N_14143);
nand U14974 (N_14974,N_14483,N_14372);
and U14975 (N_14975,N_14393,N_14266);
nand U14976 (N_14976,N_14233,N_14177);
or U14977 (N_14977,N_14260,N_14208);
and U14978 (N_14978,N_14467,N_14034);
or U14979 (N_14979,N_14177,N_14277);
and U14980 (N_14980,N_14283,N_14168);
nor U14981 (N_14981,N_14283,N_14014);
and U14982 (N_14982,N_14292,N_14352);
and U14983 (N_14983,N_14363,N_14388);
nor U14984 (N_14984,N_14288,N_14152);
or U14985 (N_14985,N_14223,N_14150);
or U14986 (N_14986,N_14461,N_14393);
or U14987 (N_14987,N_14422,N_14060);
and U14988 (N_14988,N_14280,N_14161);
or U14989 (N_14989,N_14093,N_14076);
and U14990 (N_14990,N_14355,N_14023);
or U14991 (N_14991,N_14365,N_14484);
xor U14992 (N_14992,N_14167,N_14433);
nor U14993 (N_14993,N_14210,N_14172);
and U14994 (N_14994,N_14494,N_14136);
and U14995 (N_14995,N_14162,N_14248);
and U14996 (N_14996,N_14223,N_14389);
or U14997 (N_14997,N_14384,N_14374);
and U14998 (N_14998,N_14149,N_14289);
nand U14999 (N_14999,N_14260,N_14052);
and UO_0 (O_0,N_14565,N_14760);
nand UO_1 (O_1,N_14749,N_14780);
nand UO_2 (O_2,N_14828,N_14568);
xor UO_3 (O_3,N_14811,N_14668);
and UO_4 (O_4,N_14580,N_14927);
nor UO_5 (O_5,N_14889,N_14964);
nor UO_6 (O_6,N_14783,N_14516);
and UO_7 (O_7,N_14843,N_14698);
nor UO_8 (O_8,N_14761,N_14982);
nor UO_9 (O_9,N_14710,N_14748);
and UO_10 (O_10,N_14688,N_14706);
or UO_11 (O_11,N_14894,N_14980);
nor UO_12 (O_12,N_14531,N_14941);
nor UO_13 (O_13,N_14664,N_14744);
nor UO_14 (O_14,N_14502,N_14678);
and UO_15 (O_15,N_14902,N_14996);
nand UO_16 (O_16,N_14983,N_14949);
nor UO_17 (O_17,N_14607,N_14563);
nor UO_18 (O_18,N_14882,N_14839);
nor UO_19 (O_19,N_14908,N_14835);
xor UO_20 (O_20,N_14583,N_14567);
nor UO_21 (O_21,N_14998,N_14615);
nand UO_22 (O_22,N_14766,N_14562);
nor UO_23 (O_23,N_14703,N_14801);
and UO_24 (O_24,N_14781,N_14548);
nand UO_25 (O_25,N_14573,N_14545);
xor UO_26 (O_26,N_14827,N_14662);
or UO_27 (O_27,N_14620,N_14955);
nand UO_28 (O_28,N_14920,N_14917);
nor UO_29 (O_29,N_14851,N_14966);
nor UO_30 (O_30,N_14546,N_14916);
nand UO_31 (O_31,N_14750,N_14768);
nand UO_32 (O_32,N_14708,N_14693);
and UO_33 (O_33,N_14576,N_14915);
or UO_34 (O_34,N_14676,N_14547);
and UO_35 (O_35,N_14740,N_14560);
nand UO_36 (O_36,N_14841,N_14844);
nor UO_37 (O_37,N_14868,N_14684);
and UO_38 (O_38,N_14532,N_14985);
or UO_39 (O_39,N_14695,N_14705);
and UO_40 (O_40,N_14850,N_14707);
or UO_41 (O_41,N_14875,N_14924);
nand UO_42 (O_42,N_14819,N_14519);
and UO_43 (O_43,N_14679,N_14711);
nor UO_44 (O_44,N_14566,N_14880);
and UO_45 (O_45,N_14810,N_14747);
xor UO_46 (O_46,N_14727,N_14988);
nand UO_47 (O_47,N_14777,N_14773);
and UO_48 (O_48,N_14993,N_14833);
and UO_49 (O_49,N_14655,N_14696);
or UO_50 (O_50,N_14922,N_14824);
or UO_51 (O_51,N_14571,N_14556);
nor UO_52 (O_52,N_14891,N_14601);
nor UO_53 (O_53,N_14570,N_14623);
nor UO_54 (O_54,N_14956,N_14855);
and UO_55 (O_55,N_14793,N_14522);
and UO_56 (O_56,N_14618,N_14867);
or UO_57 (O_57,N_14815,N_14848);
nand UO_58 (O_58,N_14722,N_14559);
or UO_59 (O_59,N_14860,N_14670);
or UO_60 (O_60,N_14837,N_14730);
or UO_61 (O_61,N_14977,N_14903);
and UO_62 (O_62,N_14899,N_14539);
or UO_63 (O_63,N_14804,N_14614);
or UO_64 (O_64,N_14869,N_14513);
and UO_65 (O_65,N_14973,N_14669);
xnor UO_66 (O_66,N_14770,N_14685);
or UO_67 (O_67,N_14714,N_14856);
nand UO_68 (O_68,N_14659,N_14729);
or UO_69 (O_69,N_14650,N_14818);
nor UO_70 (O_70,N_14501,N_14737);
or UO_71 (O_71,N_14692,N_14881);
nor UO_72 (O_72,N_14665,N_14950);
nor UO_73 (O_73,N_14677,N_14933);
nor UO_74 (O_74,N_14959,N_14912);
nand UO_75 (O_75,N_14581,N_14610);
nand UO_76 (O_76,N_14598,N_14872);
or UO_77 (O_77,N_14552,N_14879);
or UO_78 (O_78,N_14632,N_14716);
or UO_79 (O_79,N_14579,N_14575);
nor UO_80 (O_80,N_14978,N_14757);
and UO_81 (O_81,N_14803,N_14967);
and UO_82 (O_82,N_14800,N_14930);
or UO_83 (O_83,N_14736,N_14914);
and UO_84 (O_84,N_14994,N_14549);
nor UO_85 (O_85,N_14942,N_14555);
and UO_86 (O_86,N_14589,N_14782);
xor UO_87 (O_87,N_14686,N_14754);
or UO_88 (O_88,N_14790,N_14765);
xor UO_89 (O_89,N_14762,N_14822);
nand UO_90 (O_90,N_14619,N_14554);
and UO_91 (O_91,N_14758,N_14640);
or UO_92 (O_92,N_14616,N_14578);
nand UO_93 (O_93,N_14896,N_14667);
nand UO_94 (O_94,N_14734,N_14763);
nand UO_95 (O_95,N_14738,N_14767);
or UO_96 (O_96,N_14723,N_14681);
nor UO_97 (O_97,N_14660,N_14979);
and UO_98 (O_98,N_14853,N_14699);
nand UO_99 (O_99,N_14597,N_14622);
and UO_100 (O_100,N_14820,N_14741);
or UO_101 (O_101,N_14909,N_14874);
nor UO_102 (O_102,N_14671,N_14595);
nor UO_103 (O_103,N_14728,N_14642);
and UO_104 (O_104,N_14588,N_14506);
nor UO_105 (O_105,N_14928,N_14937);
and UO_106 (O_106,N_14943,N_14649);
nor UO_107 (O_107,N_14520,N_14558);
nor UO_108 (O_108,N_14742,N_14582);
and UO_109 (O_109,N_14631,N_14628);
and UO_110 (O_110,N_14764,N_14512);
or UO_111 (O_111,N_14842,N_14687);
nor UO_112 (O_112,N_14641,N_14821);
nand UO_113 (O_113,N_14961,N_14887);
and UO_114 (O_114,N_14858,N_14829);
nor UO_115 (O_115,N_14798,N_14591);
or UO_116 (O_116,N_14600,N_14521);
or UO_117 (O_117,N_14538,N_14795);
and UO_118 (O_118,N_14986,N_14852);
or UO_119 (O_119,N_14523,N_14613);
nand UO_120 (O_120,N_14859,N_14604);
or UO_121 (O_121,N_14854,N_14785);
nor UO_122 (O_122,N_14883,N_14505);
and UO_123 (O_123,N_14931,N_14823);
or UO_124 (O_124,N_14504,N_14787);
nand UO_125 (O_125,N_14605,N_14816);
nor UO_126 (O_126,N_14938,N_14789);
nor UO_127 (O_127,N_14926,N_14774);
and UO_128 (O_128,N_14550,N_14906);
and UO_129 (O_129,N_14694,N_14704);
and UO_130 (O_130,N_14957,N_14630);
and UO_131 (O_131,N_14892,N_14617);
nor UO_132 (O_132,N_14673,N_14680);
xnor UO_133 (O_133,N_14769,N_14870);
or UO_134 (O_134,N_14786,N_14826);
nor UO_135 (O_135,N_14971,N_14886);
nor UO_136 (O_136,N_14796,N_14536);
xnor UO_137 (O_137,N_14947,N_14845);
and UO_138 (O_138,N_14745,N_14861);
nor UO_139 (O_139,N_14974,N_14543);
and UO_140 (O_140,N_14753,N_14759);
and UO_141 (O_141,N_14923,N_14529);
or UO_142 (O_142,N_14683,N_14814);
nor UO_143 (O_143,N_14900,N_14779);
nand UO_144 (O_144,N_14788,N_14514);
xor UO_145 (O_145,N_14807,N_14962);
nor UO_146 (O_146,N_14592,N_14639);
xor UO_147 (O_147,N_14907,N_14661);
nand UO_148 (O_148,N_14603,N_14528);
or UO_149 (O_149,N_14526,N_14645);
nor UO_150 (O_150,N_14954,N_14825);
nand UO_151 (O_151,N_14876,N_14871);
or UO_152 (O_152,N_14999,N_14739);
and UO_153 (O_153,N_14602,N_14846);
or UO_154 (O_154,N_14689,N_14958);
nor UO_155 (O_155,N_14885,N_14893);
nor UO_156 (O_156,N_14690,N_14771);
nand UO_157 (O_157,N_14776,N_14658);
and UO_158 (O_158,N_14792,N_14901);
or UO_159 (O_159,N_14731,N_14976);
and UO_160 (O_160,N_14975,N_14997);
nand UO_161 (O_161,N_14895,N_14525);
nor UO_162 (O_162,N_14633,N_14718);
and UO_163 (O_163,N_14541,N_14500);
nand UO_164 (O_164,N_14542,N_14663);
and UO_165 (O_165,N_14572,N_14577);
and UO_166 (O_166,N_14989,N_14540);
nor UO_167 (O_167,N_14991,N_14561);
and UO_168 (O_168,N_14965,N_14935);
nor UO_169 (O_169,N_14551,N_14960);
or UO_170 (O_170,N_14569,N_14726);
xnor UO_171 (O_171,N_14715,N_14621);
nor UO_172 (O_172,N_14511,N_14653);
or UO_173 (O_173,N_14953,N_14934);
or UO_174 (O_174,N_14878,N_14674);
nand UO_175 (O_175,N_14805,N_14948);
and UO_176 (O_176,N_14877,N_14863);
nand UO_177 (O_177,N_14585,N_14784);
nand UO_178 (O_178,N_14637,N_14553);
and UO_179 (O_179,N_14725,N_14596);
nand UO_180 (O_180,N_14936,N_14697);
and UO_181 (O_181,N_14702,N_14629);
or UO_182 (O_182,N_14939,N_14508);
nor UO_183 (O_183,N_14918,N_14813);
nand UO_184 (O_184,N_14509,N_14831);
nor UO_185 (O_185,N_14862,N_14832);
nor UO_186 (O_186,N_14682,N_14574);
nand UO_187 (O_187,N_14524,N_14636);
nand UO_188 (O_188,N_14712,N_14952);
nand UO_189 (O_189,N_14751,N_14987);
and UO_190 (O_190,N_14656,N_14651);
and UO_191 (O_191,N_14992,N_14535);
nor UO_192 (O_192,N_14691,N_14590);
nor UO_193 (O_193,N_14945,N_14969);
nand UO_194 (O_194,N_14817,N_14534);
or UO_195 (O_195,N_14995,N_14913);
nand UO_196 (O_196,N_14806,N_14984);
and UO_197 (O_197,N_14611,N_14990);
nor UO_198 (O_198,N_14627,N_14772);
nand UO_199 (O_199,N_14724,N_14517);
nor UO_200 (O_200,N_14634,N_14756);
and UO_201 (O_201,N_14544,N_14840);
nor UO_202 (O_202,N_14503,N_14657);
nor UO_203 (O_203,N_14612,N_14733);
nor UO_204 (O_204,N_14701,N_14672);
and UO_205 (O_205,N_14797,N_14646);
nand UO_206 (O_206,N_14932,N_14515);
nand UO_207 (O_207,N_14857,N_14905);
nand UO_208 (O_208,N_14530,N_14865);
and UO_209 (O_209,N_14925,N_14537);
nor UO_210 (O_210,N_14652,N_14970);
nand UO_211 (O_211,N_14735,N_14904);
or UO_212 (O_212,N_14866,N_14951);
and UO_213 (O_213,N_14599,N_14638);
and UO_214 (O_214,N_14752,N_14518);
nand UO_215 (O_215,N_14719,N_14721);
and UO_216 (O_216,N_14775,N_14981);
nand UO_217 (O_217,N_14910,N_14849);
nor UO_218 (O_218,N_14564,N_14890);
or UO_219 (O_219,N_14743,N_14713);
or UO_220 (O_220,N_14587,N_14864);
or UO_221 (O_221,N_14606,N_14709);
nand UO_222 (O_222,N_14608,N_14898);
nor UO_223 (O_223,N_14921,N_14812);
nor UO_224 (O_224,N_14666,N_14897);
and UO_225 (O_225,N_14802,N_14647);
and UO_226 (O_226,N_14584,N_14700);
nor UO_227 (O_227,N_14838,N_14963);
and UO_228 (O_228,N_14873,N_14830);
and UO_229 (O_229,N_14746,N_14648);
nor UO_230 (O_230,N_14809,N_14778);
xor UO_231 (O_231,N_14929,N_14625);
or UO_232 (O_232,N_14884,N_14968);
and UO_233 (O_233,N_14755,N_14834);
nor UO_234 (O_234,N_14533,N_14510);
nor UO_235 (O_235,N_14720,N_14791);
or UO_236 (O_236,N_14717,N_14609);
nor UO_237 (O_237,N_14919,N_14940);
or UO_238 (O_238,N_14593,N_14794);
nor UO_239 (O_239,N_14946,N_14557);
and UO_240 (O_240,N_14644,N_14527);
nor UO_241 (O_241,N_14888,N_14654);
or UO_242 (O_242,N_14586,N_14675);
xor UO_243 (O_243,N_14808,N_14626);
nand UO_244 (O_244,N_14799,N_14944);
nand UO_245 (O_245,N_14732,N_14594);
nor UO_246 (O_246,N_14507,N_14972);
nand UO_247 (O_247,N_14836,N_14847);
or UO_248 (O_248,N_14643,N_14911);
or UO_249 (O_249,N_14635,N_14624);
xnor UO_250 (O_250,N_14947,N_14698);
nand UO_251 (O_251,N_14947,N_14550);
nor UO_252 (O_252,N_14838,N_14613);
and UO_253 (O_253,N_14596,N_14847);
nor UO_254 (O_254,N_14529,N_14525);
or UO_255 (O_255,N_14717,N_14691);
nor UO_256 (O_256,N_14917,N_14562);
nor UO_257 (O_257,N_14591,N_14890);
nand UO_258 (O_258,N_14723,N_14677);
xor UO_259 (O_259,N_14944,N_14933);
nor UO_260 (O_260,N_14526,N_14793);
or UO_261 (O_261,N_14893,N_14693);
nor UO_262 (O_262,N_14689,N_14808);
nand UO_263 (O_263,N_14863,N_14796);
nand UO_264 (O_264,N_14893,N_14939);
nand UO_265 (O_265,N_14790,N_14856);
nand UO_266 (O_266,N_14718,N_14861);
and UO_267 (O_267,N_14560,N_14657);
xnor UO_268 (O_268,N_14850,N_14989);
or UO_269 (O_269,N_14561,N_14565);
or UO_270 (O_270,N_14814,N_14865);
and UO_271 (O_271,N_14545,N_14976);
or UO_272 (O_272,N_14864,N_14688);
nor UO_273 (O_273,N_14570,N_14919);
nand UO_274 (O_274,N_14577,N_14554);
and UO_275 (O_275,N_14943,N_14617);
nor UO_276 (O_276,N_14598,N_14988);
nor UO_277 (O_277,N_14553,N_14985);
nor UO_278 (O_278,N_14758,N_14775);
and UO_279 (O_279,N_14797,N_14867);
and UO_280 (O_280,N_14744,N_14626);
and UO_281 (O_281,N_14705,N_14976);
nand UO_282 (O_282,N_14929,N_14963);
nor UO_283 (O_283,N_14885,N_14537);
and UO_284 (O_284,N_14632,N_14741);
nand UO_285 (O_285,N_14965,N_14882);
or UO_286 (O_286,N_14815,N_14691);
or UO_287 (O_287,N_14911,N_14892);
and UO_288 (O_288,N_14629,N_14875);
or UO_289 (O_289,N_14749,N_14784);
nor UO_290 (O_290,N_14736,N_14526);
xnor UO_291 (O_291,N_14627,N_14653);
xnor UO_292 (O_292,N_14599,N_14569);
nor UO_293 (O_293,N_14696,N_14691);
or UO_294 (O_294,N_14969,N_14527);
xnor UO_295 (O_295,N_14678,N_14789);
and UO_296 (O_296,N_14951,N_14603);
or UO_297 (O_297,N_14726,N_14659);
nand UO_298 (O_298,N_14814,N_14626);
or UO_299 (O_299,N_14963,N_14503);
xnor UO_300 (O_300,N_14947,N_14998);
or UO_301 (O_301,N_14741,N_14960);
and UO_302 (O_302,N_14873,N_14899);
or UO_303 (O_303,N_14542,N_14682);
nor UO_304 (O_304,N_14723,N_14814);
nor UO_305 (O_305,N_14599,N_14830);
and UO_306 (O_306,N_14982,N_14888);
nor UO_307 (O_307,N_14983,N_14508);
or UO_308 (O_308,N_14848,N_14830);
and UO_309 (O_309,N_14555,N_14685);
nand UO_310 (O_310,N_14830,N_14667);
nand UO_311 (O_311,N_14512,N_14509);
xor UO_312 (O_312,N_14628,N_14602);
or UO_313 (O_313,N_14589,N_14728);
and UO_314 (O_314,N_14911,N_14786);
nor UO_315 (O_315,N_14642,N_14754);
and UO_316 (O_316,N_14680,N_14516);
nor UO_317 (O_317,N_14635,N_14752);
nor UO_318 (O_318,N_14981,N_14858);
nand UO_319 (O_319,N_14884,N_14533);
and UO_320 (O_320,N_14898,N_14970);
nand UO_321 (O_321,N_14663,N_14865);
and UO_322 (O_322,N_14968,N_14826);
or UO_323 (O_323,N_14610,N_14957);
or UO_324 (O_324,N_14585,N_14972);
xor UO_325 (O_325,N_14970,N_14768);
and UO_326 (O_326,N_14840,N_14748);
and UO_327 (O_327,N_14696,N_14546);
and UO_328 (O_328,N_14641,N_14675);
or UO_329 (O_329,N_14692,N_14978);
and UO_330 (O_330,N_14584,N_14563);
or UO_331 (O_331,N_14979,N_14807);
and UO_332 (O_332,N_14616,N_14803);
nand UO_333 (O_333,N_14739,N_14633);
nor UO_334 (O_334,N_14987,N_14785);
or UO_335 (O_335,N_14861,N_14855);
and UO_336 (O_336,N_14864,N_14691);
nand UO_337 (O_337,N_14517,N_14613);
or UO_338 (O_338,N_14721,N_14664);
nand UO_339 (O_339,N_14956,N_14870);
or UO_340 (O_340,N_14671,N_14551);
or UO_341 (O_341,N_14879,N_14927);
nor UO_342 (O_342,N_14629,N_14527);
nand UO_343 (O_343,N_14782,N_14772);
nor UO_344 (O_344,N_14710,N_14550);
xor UO_345 (O_345,N_14795,N_14566);
and UO_346 (O_346,N_14734,N_14799);
nand UO_347 (O_347,N_14812,N_14920);
and UO_348 (O_348,N_14888,N_14912);
or UO_349 (O_349,N_14931,N_14506);
nor UO_350 (O_350,N_14752,N_14606);
nor UO_351 (O_351,N_14591,N_14683);
and UO_352 (O_352,N_14993,N_14952);
and UO_353 (O_353,N_14925,N_14988);
and UO_354 (O_354,N_14723,N_14928);
nand UO_355 (O_355,N_14536,N_14912);
or UO_356 (O_356,N_14635,N_14743);
and UO_357 (O_357,N_14516,N_14796);
nor UO_358 (O_358,N_14602,N_14932);
nand UO_359 (O_359,N_14737,N_14691);
nand UO_360 (O_360,N_14616,N_14862);
nor UO_361 (O_361,N_14905,N_14910);
or UO_362 (O_362,N_14609,N_14872);
nor UO_363 (O_363,N_14946,N_14763);
nor UO_364 (O_364,N_14780,N_14635);
xnor UO_365 (O_365,N_14910,N_14940);
or UO_366 (O_366,N_14652,N_14685);
xnor UO_367 (O_367,N_14966,N_14916);
nor UO_368 (O_368,N_14896,N_14849);
nor UO_369 (O_369,N_14740,N_14543);
or UO_370 (O_370,N_14812,N_14967);
and UO_371 (O_371,N_14978,N_14750);
and UO_372 (O_372,N_14684,N_14863);
nor UO_373 (O_373,N_14810,N_14539);
xnor UO_374 (O_374,N_14865,N_14816);
nor UO_375 (O_375,N_14543,N_14832);
xor UO_376 (O_376,N_14738,N_14731);
xnor UO_377 (O_377,N_14787,N_14636);
nor UO_378 (O_378,N_14539,N_14661);
xnor UO_379 (O_379,N_14842,N_14549);
nor UO_380 (O_380,N_14784,N_14591);
nand UO_381 (O_381,N_14960,N_14881);
and UO_382 (O_382,N_14831,N_14525);
nand UO_383 (O_383,N_14773,N_14656);
xor UO_384 (O_384,N_14550,N_14636);
nor UO_385 (O_385,N_14893,N_14841);
nor UO_386 (O_386,N_14585,N_14732);
and UO_387 (O_387,N_14586,N_14744);
nand UO_388 (O_388,N_14714,N_14666);
nor UO_389 (O_389,N_14546,N_14767);
xor UO_390 (O_390,N_14627,N_14996);
nor UO_391 (O_391,N_14771,N_14714);
or UO_392 (O_392,N_14655,N_14952);
nand UO_393 (O_393,N_14505,N_14977);
or UO_394 (O_394,N_14504,N_14958);
or UO_395 (O_395,N_14600,N_14875);
nand UO_396 (O_396,N_14813,N_14936);
nand UO_397 (O_397,N_14938,N_14779);
nor UO_398 (O_398,N_14667,N_14884);
nand UO_399 (O_399,N_14738,N_14770);
or UO_400 (O_400,N_14672,N_14983);
or UO_401 (O_401,N_14957,N_14527);
and UO_402 (O_402,N_14854,N_14866);
and UO_403 (O_403,N_14724,N_14813);
nand UO_404 (O_404,N_14927,N_14902);
nor UO_405 (O_405,N_14673,N_14755);
and UO_406 (O_406,N_14572,N_14837);
nor UO_407 (O_407,N_14686,N_14889);
nor UO_408 (O_408,N_14820,N_14784);
nor UO_409 (O_409,N_14515,N_14501);
nor UO_410 (O_410,N_14621,N_14624);
xnor UO_411 (O_411,N_14666,N_14778);
nor UO_412 (O_412,N_14883,N_14634);
xor UO_413 (O_413,N_14606,N_14579);
and UO_414 (O_414,N_14689,N_14778);
nand UO_415 (O_415,N_14922,N_14672);
nor UO_416 (O_416,N_14711,N_14581);
nor UO_417 (O_417,N_14506,N_14500);
or UO_418 (O_418,N_14862,N_14758);
xnor UO_419 (O_419,N_14737,N_14570);
nand UO_420 (O_420,N_14756,N_14973);
or UO_421 (O_421,N_14567,N_14577);
nand UO_422 (O_422,N_14628,N_14577);
and UO_423 (O_423,N_14966,N_14909);
nand UO_424 (O_424,N_14924,N_14967);
or UO_425 (O_425,N_14801,N_14826);
and UO_426 (O_426,N_14921,N_14809);
nor UO_427 (O_427,N_14948,N_14767);
nand UO_428 (O_428,N_14885,N_14956);
nand UO_429 (O_429,N_14805,N_14696);
xnor UO_430 (O_430,N_14924,N_14688);
and UO_431 (O_431,N_14980,N_14757);
and UO_432 (O_432,N_14705,N_14847);
or UO_433 (O_433,N_14598,N_14622);
nor UO_434 (O_434,N_14894,N_14839);
and UO_435 (O_435,N_14505,N_14979);
and UO_436 (O_436,N_14925,N_14877);
or UO_437 (O_437,N_14520,N_14820);
or UO_438 (O_438,N_14784,N_14661);
nand UO_439 (O_439,N_14805,N_14861);
nand UO_440 (O_440,N_14904,N_14528);
nor UO_441 (O_441,N_14669,N_14572);
nand UO_442 (O_442,N_14804,N_14915);
or UO_443 (O_443,N_14968,N_14923);
nand UO_444 (O_444,N_14847,N_14697);
or UO_445 (O_445,N_14890,N_14942);
nand UO_446 (O_446,N_14881,N_14605);
xor UO_447 (O_447,N_14609,N_14918);
nand UO_448 (O_448,N_14749,N_14625);
nor UO_449 (O_449,N_14891,N_14612);
and UO_450 (O_450,N_14643,N_14709);
nand UO_451 (O_451,N_14548,N_14640);
and UO_452 (O_452,N_14790,N_14989);
nor UO_453 (O_453,N_14785,N_14820);
or UO_454 (O_454,N_14517,N_14684);
xnor UO_455 (O_455,N_14713,N_14924);
nand UO_456 (O_456,N_14953,N_14739);
nor UO_457 (O_457,N_14677,N_14871);
and UO_458 (O_458,N_14992,N_14946);
or UO_459 (O_459,N_14610,N_14662);
xnor UO_460 (O_460,N_14996,N_14571);
nand UO_461 (O_461,N_14585,N_14531);
and UO_462 (O_462,N_14621,N_14583);
xnor UO_463 (O_463,N_14576,N_14789);
nor UO_464 (O_464,N_14983,N_14538);
xor UO_465 (O_465,N_14643,N_14646);
nand UO_466 (O_466,N_14721,N_14691);
and UO_467 (O_467,N_14573,N_14541);
nand UO_468 (O_468,N_14973,N_14994);
nor UO_469 (O_469,N_14953,N_14856);
or UO_470 (O_470,N_14594,N_14772);
nor UO_471 (O_471,N_14508,N_14786);
nor UO_472 (O_472,N_14787,N_14714);
xnor UO_473 (O_473,N_14737,N_14653);
nor UO_474 (O_474,N_14960,N_14603);
nand UO_475 (O_475,N_14980,N_14633);
and UO_476 (O_476,N_14674,N_14759);
or UO_477 (O_477,N_14810,N_14858);
nand UO_478 (O_478,N_14705,N_14898);
or UO_479 (O_479,N_14585,N_14507);
nand UO_480 (O_480,N_14607,N_14809);
nand UO_481 (O_481,N_14970,N_14556);
and UO_482 (O_482,N_14692,N_14669);
nand UO_483 (O_483,N_14597,N_14765);
or UO_484 (O_484,N_14732,N_14871);
and UO_485 (O_485,N_14756,N_14892);
and UO_486 (O_486,N_14972,N_14803);
xnor UO_487 (O_487,N_14984,N_14561);
nand UO_488 (O_488,N_14595,N_14783);
nand UO_489 (O_489,N_14871,N_14583);
nand UO_490 (O_490,N_14514,N_14540);
or UO_491 (O_491,N_14629,N_14880);
or UO_492 (O_492,N_14678,N_14859);
and UO_493 (O_493,N_14646,N_14860);
xor UO_494 (O_494,N_14793,N_14651);
or UO_495 (O_495,N_14828,N_14590);
or UO_496 (O_496,N_14948,N_14947);
or UO_497 (O_497,N_14588,N_14876);
or UO_498 (O_498,N_14670,N_14680);
or UO_499 (O_499,N_14774,N_14767);
nor UO_500 (O_500,N_14743,N_14973);
nand UO_501 (O_501,N_14988,N_14915);
nand UO_502 (O_502,N_14711,N_14685);
nand UO_503 (O_503,N_14702,N_14543);
and UO_504 (O_504,N_14526,N_14533);
nor UO_505 (O_505,N_14541,N_14764);
or UO_506 (O_506,N_14623,N_14599);
nor UO_507 (O_507,N_14884,N_14924);
nand UO_508 (O_508,N_14791,N_14789);
and UO_509 (O_509,N_14928,N_14884);
or UO_510 (O_510,N_14783,N_14964);
xor UO_511 (O_511,N_14891,N_14514);
nand UO_512 (O_512,N_14792,N_14811);
nor UO_513 (O_513,N_14504,N_14598);
and UO_514 (O_514,N_14918,N_14616);
and UO_515 (O_515,N_14668,N_14690);
and UO_516 (O_516,N_14858,N_14507);
nand UO_517 (O_517,N_14524,N_14856);
xnor UO_518 (O_518,N_14573,N_14966);
nor UO_519 (O_519,N_14628,N_14579);
or UO_520 (O_520,N_14638,N_14584);
or UO_521 (O_521,N_14798,N_14599);
nand UO_522 (O_522,N_14767,N_14551);
and UO_523 (O_523,N_14995,N_14789);
and UO_524 (O_524,N_14744,N_14506);
and UO_525 (O_525,N_14920,N_14747);
nor UO_526 (O_526,N_14748,N_14664);
and UO_527 (O_527,N_14764,N_14730);
nand UO_528 (O_528,N_14523,N_14678);
and UO_529 (O_529,N_14550,N_14801);
and UO_530 (O_530,N_14675,N_14553);
nand UO_531 (O_531,N_14802,N_14771);
nor UO_532 (O_532,N_14912,N_14883);
nor UO_533 (O_533,N_14984,N_14930);
nand UO_534 (O_534,N_14725,N_14668);
or UO_535 (O_535,N_14632,N_14743);
or UO_536 (O_536,N_14630,N_14954);
and UO_537 (O_537,N_14715,N_14635);
and UO_538 (O_538,N_14894,N_14717);
xor UO_539 (O_539,N_14578,N_14501);
nand UO_540 (O_540,N_14880,N_14850);
xor UO_541 (O_541,N_14848,N_14521);
or UO_542 (O_542,N_14901,N_14625);
or UO_543 (O_543,N_14688,N_14721);
nor UO_544 (O_544,N_14614,N_14993);
and UO_545 (O_545,N_14934,N_14503);
or UO_546 (O_546,N_14665,N_14663);
and UO_547 (O_547,N_14563,N_14817);
or UO_548 (O_548,N_14510,N_14812);
nor UO_549 (O_549,N_14509,N_14514);
or UO_550 (O_550,N_14929,N_14724);
and UO_551 (O_551,N_14518,N_14780);
and UO_552 (O_552,N_14684,N_14620);
nor UO_553 (O_553,N_14898,N_14888);
and UO_554 (O_554,N_14553,N_14819);
nand UO_555 (O_555,N_14967,N_14706);
nand UO_556 (O_556,N_14757,N_14520);
nand UO_557 (O_557,N_14775,N_14968);
xnor UO_558 (O_558,N_14931,N_14867);
nand UO_559 (O_559,N_14976,N_14606);
nor UO_560 (O_560,N_14599,N_14592);
and UO_561 (O_561,N_14804,N_14648);
nor UO_562 (O_562,N_14860,N_14813);
nand UO_563 (O_563,N_14761,N_14646);
nor UO_564 (O_564,N_14867,N_14704);
and UO_565 (O_565,N_14728,N_14626);
xnor UO_566 (O_566,N_14879,N_14984);
xnor UO_567 (O_567,N_14597,N_14516);
nand UO_568 (O_568,N_14873,N_14569);
and UO_569 (O_569,N_14817,N_14646);
and UO_570 (O_570,N_14610,N_14576);
and UO_571 (O_571,N_14725,N_14953);
nand UO_572 (O_572,N_14971,N_14973);
or UO_573 (O_573,N_14936,N_14927);
nor UO_574 (O_574,N_14741,N_14828);
and UO_575 (O_575,N_14684,N_14965);
nor UO_576 (O_576,N_14827,N_14665);
and UO_577 (O_577,N_14967,N_14966);
nor UO_578 (O_578,N_14910,N_14655);
nand UO_579 (O_579,N_14892,N_14532);
xor UO_580 (O_580,N_14690,N_14635);
nand UO_581 (O_581,N_14802,N_14741);
or UO_582 (O_582,N_14709,N_14585);
or UO_583 (O_583,N_14770,N_14524);
and UO_584 (O_584,N_14937,N_14741);
and UO_585 (O_585,N_14918,N_14967);
xnor UO_586 (O_586,N_14740,N_14503);
nand UO_587 (O_587,N_14556,N_14543);
and UO_588 (O_588,N_14594,N_14937);
nor UO_589 (O_589,N_14895,N_14810);
nor UO_590 (O_590,N_14818,N_14729);
or UO_591 (O_591,N_14735,N_14612);
xnor UO_592 (O_592,N_14675,N_14932);
and UO_593 (O_593,N_14735,N_14618);
xnor UO_594 (O_594,N_14515,N_14968);
or UO_595 (O_595,N_14535,N_14968);
nand UO_596 (O_596,N_14897,N_14781);
nand UO_597 (O_597,N_14689,N_14746);
or UO_598 (O_598,N_14638,N_14539);
nand UO_599 (O_599,N_14956,N_14904);
and UO_600 (O_600,N_14802,N_14503);
nand UO_601 (O_601,N_14917,N_14933);
nor UO_602 (O_602,N_14780,N_14651);
nand UO_603 (O_603,N_14854,N_14971);
xor UO_604 (O_604,N_14922,N_14564);
and UO_605 (O_605,N_14944,N_14804);
and UO_606 (O_606,N_14980,N_14822);
and UO_607 (O_607,N_14863,N_14966);
nand UO_608 (O_608,N_14522,N_14896);
or UO_609 (O_609,N_14937,N_14604);
or UO_610 (O_610,N_14594,N_14556);
xnor UO_611 (O_611,N_14940,N_14741);
or UO_612 (O_612,N_14572,N_14868);
or UO_613 (O_613,N_14777,N_14730);
nand UO_614 (O_614,N_14835,N_14733);
nand UO_615 (O_615,N_14561,N_14968);
nor UO_616 (O_616,N_14688,N_14866);
nor UO_617 (O_617,N_14500,N_14925);
or UO_618 (O_618,N_14740,N_14794);
xor UO_619 (O_619,N_14550,N_14585);
nor UO_620 (O_620,N_14606,N_14820);
and UO_621 (O_621,N_14848,N_14560);
and UO_622 (O_622,N_14636,N_14880);
and UO_623 (O_623,N_14879,N_14748);
nand UO_624 (O_624,N_14942,N_14596);
or UO_625 (O_625,N_14820,N_14564);
nor UO_626 (O_626,N_14845,N_14648);
or UO_627 (O_627,N_14587,N_14618);
nor UO_628 (O_628,N_14908,N_14518);
nand UO_629 (O_629,N_14664,N_14688);
nor UO_630 (O_630,N_14758,N_14813);
or UO_631 (O_631,N_14732,N_14971);
and UO_632 (O_632,N_14933,N_14880);
nor UO_633 (O_633,N_14828,N_14659);
nor UO_634 (O_634,N_14549,N_14672);
xnor UO_635 (O_635,N_14656,N_14706);
or UO_636 (O_636,N_14787,N_14700);
and UO_637 (O_637,N_14537,N_14624);
nand UO_638 (O_638,N_14697,N_14888);
nor UO_639 (O_639,N_14968,N_14602);
nand UO_640 (O_640,N_14617,N_14854);
nor UO_641 (O_641,N_14607,N_14716);
nand UO_642 (O_642,N_14952,N_14521);
or UO_643 (O_643,N_14715,N_14576);
and UO_644 (O_644,N_14866,N_14887);
nor UO_645 (O_645,N_14591,N_14534);
or UO_646 (O_646,N_14811,N_14910);
nand UO_647 (O_647,N_14719,N_14635);
xnor UO_648 (O_648,N_14913,N_14756);
or UO_649 (O_649,N_14764,N_14543);
or UO_650 (O_650,N_14643,N_14781);
xnor UO_651 (O_651,N_14926,N_14510);
and UO_652 (O_652,N_14725,N_14708);
or UO_653 (O_653,N_14664,N_14763);
nand UO_654 (O_654,N_14976,N_14938);
and UO_655 (O_655,N_14893,N_14925);
nor UO_656 (O_656,N_14514,N_14848);
nor UO_657 (O_657,N_14943,N_14865);
nand UO_658 (O_658,N_14843,N_14618);
nor UO_659 (O_659,N_14745,N_14770);
or UO_660 (O_660,N_14860,N_14718);
and UO_661 (O_661,N_14866,N_14585);
xor UO_662 (O_662,N_14551,N_14718);
and UO_663 (O_663,N_14826,N_14994);
nor UO_664 (O_664,N_14870,N_14726);
nor UO_665 (O_665,N_14525,N_14863);
nand UO_666 (O_666,N_14636,N_14777);
or UO_667 (O_667,N_14975,N_14878);
nor UO_668 (O_668,N_14653,N_14644);
or UO_669 (O_669,N_14798,N_14818);
xor UO_670 (O_670,N_14986,N_14959);
nand UO_671 (O_671,N_14509,N_14723);
nor UO_672 (O_672,N_14539,N_14618);
or UO_673 (O_673,N_14672,N_14984);
and UO_674 (O_674,N_14744,N_14937);
or UO_675 (O_675,N_14835,N_14720);
or UO_676 (O_676,N_14755,N_14898);
nand UO_677 (O_677,N_14672,N_14945);
or UO_678 (O_678,N_14804,N_14929);
nor UO_679 (O_679,N_14765,N_14850);
or UO_680 (O_680,N_14574,N_14575);
nand UO_681 (O_681,N_14775,N_14771);
xor UO_682 (O_682,N_14956,N_14821);
nor UO_683 (O_683,N_14888,N_14700);
nand UO_684 (O_684,N_14826,N_14844);
nor UO_685 (O_685,N_14605,N_14825);
nand UO_686 (O_686,N_14927,N_14523);
nand UO_687 (O_687,N_14853,N_14769);
and UO_688 (O_688,N_14715,N_14676);
and UO_689 (O_689,N_14786,N_14925);
or UO_690 (O_690,N_14744,N_14957);
nor UO_691 (O_691,N_14632,N_14729);
nand UO_692 (O_692,N_14776,N_14515);
and UO_693 (O_693,N_14571,N_14879);
and UO_694 (O_694,N_14989,N_14544);
nor UO_695 (O_695,N_14636,N_14986);
nor UO_696 (O_696,N_14859,N_14527);
nor UO_697 (O_697,N_14619,N_14770);
nor UO_698 (O_698,N_14558,N_14909);
xor UO_699 (O_699,N_14545,N_14821);
nand UO_700 (O_700,N_14890,N_14828);
and UO_701 (O_701,N_14705,N_14876);
or UO_702 (O_702,N_14868,N_14902);
nand UO_703 (O_703,N_14923,N_14734);
or UO_704 (O_704,N_14769,N_14886);
nor UO_705 (O_705,N_14765,N_14570);
nand UO_706 (O_706,N_14804,N_14547);
and UO_707 (O_707,N_14505,N_14828);
or UO_708 (O_708,N_14957,N_14574);
nor UO_709 (O_709,N_14943,N_14828);
nor UO_710 (O_710,N_14783,N_14735);
nand UO_711 (O_711,N_14512,N_14576);
nor UO_712 (O_712,N_14600,N_14874);
xnor UO_713 (O_713,N_14853,N_14654);
or UO_714 (O_714,N_14740,N_14940);
or UO_715 (O_715,N_14872,N_14553);
and UO_716 (O_716,N_14955,N_14546);
and UO_717 (O_717,N_14761,N_14724);
and UO_718 (O_718,N_14650,N_14545);
and UO_719 (O_719,N_14547,N_14972);
or UO_720 (O_720,N_14556,N_14777);
xor UO_721 (O_721,N_14889,N_14886);
or UO_722 (O_722,N_14931,N_14915);
nor UO_723 (O_723,N_14598,N_14599);
nand UO_724 (O_724,N_14923,N_14564);
or UO_725 (O_725,N_14830,N_14636);
and UO_726 (O_726,N_14711,N_14871);
or UO_727 (O_727,N_14639,N_14590);
and UO_728 (O_728,N_14645,N_14717);
and UO_729 (O_729,N_14953,N_14517);
nand UO_730 (O_730,N_14578,N_14689);
nand UO_731 (O_731,N_14787,N_14862);
xnor UO_732 (O_732,N_14740,N_14722);
nor UO_733 (O_733,N_14801,N_14877);
or UO_734 (O_734,N_14826,N_14680);
nand UO_735 (O_735,N_14587,N_14506);
and UO_736 (O_736,N_14509,N_14823);
nand UO_737 (O_737,N_14502,N_14523);
or UO_738 (O_738,N_14910,N_14624);
nand UO_739 (O_739,N_14684,N_14767);
or UO_740 (O_740,N_14857,N_14875);
and UO_741 (O_741,N_14947,N_14971);
or UO_742 (O_742,N_14766,N_14783);
or UO_743 (O_743,N_14725,N_14511);
and UO_744 (O_744,N_14551,N_14656);
nand UO_745 (O_745,N_14552,N_14603);
nor UO_746 (O_746,N_14614,N_14726);
nor UO_747 (O_747,N_14599,N_14993);
or UO_748 (O_748,N_14554,N_14719);
and UO_749 (O_749,N_14856,N_14657);
or UO_750 (O_750,N_14797,N_14517);
and UO_751 (O_751,N_14779,N_14530);
nor UO_752 (O_752,N_14666,N_14980);
and UO_753 (O_753,N_14776,N_14513);
or UO_754 (O_754,N_14839,N_14680);
nand UO_755 (O_755,N_14531,N_14619);
and UO_756 (O_756,N_14519,N_14895);
and UO_757 (O_757,N_14740,N_14619);
nand UO_758 (O_758,N_14871,N_14671);
nand UO_759 (O_759,N_14861,N_14948);
or UO_760 (O_760,N_14862,N_14830);
nand UO_761 (O_761,N_14912,N_14508);
nand UO_762 (O_762,N_14639,N_14735);
nor UO_763 (O_763,N_14953,N_14625);
nor UO_764 (O_764,N_14892,N_14916);
nand UO_765 (O_765,N_14599,N_14733);
and UO_766 (O_766,N_14887,N_14545);
nor UO_767 (O_767,N_14594,N_14765);
or UO_768 (O_768,N_14542,N_14501);
or UO_769 (O_769,N_14983,N_14970);
and UO_770 (O_770,N_14578,N_14767);
nand UO_771 (O_771,N_14646,N_14551);
xor UO_772 (O_772,N_14513,N_14982);
or UO_773 (O_773,N_14732,N_14748);
and UO_774 (O_774,N_14853,N_14694);
nor UO_775 (O_775,N_14535,N_14562);
nand UO_776 (O_776,N_14633,N_14630);
and UO_777 (O_777,N_14915,N_14708);
xnor UO_778 (O_778,N_14785,N_14700);
nand UO_779 (O_779,N_14965,N_14983);
and UO_780 (O_780,N_14533,N_14870);
nand UO_781 (O_781,N_14773,N_14920);
and UO_782 (O_782,N_14994,N_14964);
nor UO_783 (O_783,N_14523,N_14797);
nand UO_784 (O_784,N_14842,N_14911);
nor UO_785 (O_785,N_14827,N_14694);
nor UO_786 (O_786,N_14664,N_14896);
nor UO_787 (O_787,N_14681,N_14819);
or UO_788 (O_788,N_14673,N_14999);
xnor UO_789 (O_789,N_14740,N_14554);
or UO_790 (O_790,N_14647,N_14715);
nand UO_791 (O_791,N_14527,N_14576);
or UO_792 (O_792,N_14983,N_14998);
nor UO_793 (O_793,N_14835,N_14566);
nand UO_794 (O_794,N_14995,N_14696);
or UO_795 (O_795,N_14680,N_14960);
nor UO_796 (O_796,N_14643,N_14663);
nand UO_797 (O_797,N_14886,N_14682);
nand UO_798 (O_798,N_14845,N_14782);
nor UO_799 (O_799,N_14828,N_14711);
nor UO_800 (O_800,N_14932,N_14825);
and UO_801 (O_801,N_14683,N_14894);
nand UO_802 (O_802,N_14713,N_14836);
nor UO_803 (O_803,N_14644,N_14990);
nand UO_804 (O_804,N_14773,N_14559);
nand UO_805 (O_805,N_14835,N_14705);
or UO_806 (O_806,N_14776,N_14837);
nand UO_807 (O_807,N_14726,N_14910);
nand UO_808 (O_808,N_14923,N_14708);
nand UO_809 (O_809,N_14737,N_14906);
or UO_810 (O_810,N_14737,N_14614);
or UO_811 (O_811,N_14552,N_14810);
nand UO_812 (O_812,N_14979,N_14608);
nand UO_813 (O_813,N_14539,N_14613);
and UO_814 (O_814,N_14663,N_14828);
or UO_815 (O_815,N_14730,N_14685);
or UO_816 (O_816,N_14742,N_14671);
nor UO_817 (O_817,N_14631,N_14767);
and UO_818 (O_818,N_14789,N_14542);
and UO_819 (O_819,N_14504,N_14748);
xnor UO_820 (O_820,N_14875,N_14957);
and UO_821 (O_821,N_14689,N_14608);
or UO_822 (O_822,N_14711,N_14831);
xor UO_823 (O_823,N_14533,N_14597);
nor UO_824 (O_824,N_14951,N_14696);
and UO_825 (O_825,N_14500,N_14715);
and UO_826 (O_826,N_14976,N_14751);
nand UO_827 (O_827,N_14866,N_14757);
nand UO_828 (O_828,N_14997,N_14784);
or UO_829 (O_829,N_14689,N_14520);
nor UO_830 (O_830,N_14985,N_14747);
xnor UO_831 (O_831,N_14795,N_14509);
and UO_832 (O_832,N_14575,N_14981);
and UO_833 (O_833,N_14865,N_14926);
nand UO_834 (O_834,N_14864,N_14933);
or UO_835 (O_835,N_14584,N_14687);
nand UO_836 (O_836,N_14527,N_14658);
nor UO_837 (O_837,N_14596,N_14644);
xnor UO_838 (O_838,N_14640,N_14769);
nor UO_839 (O_839,N_14787,N_14994);
and UO_840 (O_840,N_14917,N_14802);
nor UO_841 (O_841,N_14995,N_14576);
nor UO_842 (O_842,N_14593,N_14874);
nand UO_843 (O_843,N_14634,N_14816);
or UO_844 (O_844,N_14778,N_14820);
nor UO_845 (O_845,N_14830,N_14606);
nand UO_846 (O_846,N_14975,N_14874);
nand UO_847 (O_847,N_14535,N_14599);
xor UO_848 (O_848,N_14547,N_14991);
or UO_849 (O_849,N_14887,N_14639);
nor UO_850 (O_850,N_14536,N_14938);
or UO_851 (O_851,N_14608,N_14903);
nand UO_852 (O_852,N_14623,N_14843);
and UO_853 (O_853,N_14850,N_14505);
and UO_854 (O_854,N_14991,N_14506);
and UO_855 (O_855,N_14782,N_14885);
nor UO_856 (O_856,N_14620,N_14639);
nor UO_857 (O_857,N_14503,N_14691);
nand UO_858 (O_858,N_14887,N_14680);
nand UO_859 (O_859,N_14849,N_14993);
xor UO_860 (O_860,N_14684,N_14604);
nor UO_861 (O_861,N_14985,N_14679);
nor UO_862 (O_862,N_14570,N_14508);
xnor UO_863 (O_863,N_14957,N_14530);
nand UO_864 (O_864,N_14962,N_14627);
nand UO_865 (O_865,N_14852,N_14747);
nand UO_866 (O_866,N_14906,N_14908);
and UO_867 (O_867,N_14603,N_14946);
nand UO_868 (O_868,N_14684,N_14651);
and UO_869 (O_869,N_14923,N_14558);
nand UO_870 (O_870,N_14614,N_14680);
nand UO_871 (O_871,N_14623,N_14567);
nand UO_872 (O_872,N_14506,N_14852);
or UO_873 (O_873,N_14587,N_14984);
nand UO_874 (O_874,N_14511,N_14932);
or UO_875 (O_875,N_14621,N_14516);
nor UO_876 (O_876,N_14509,N_14678);
nand UO_877 (O_877,N_14743,N_14985);
nand UO_878 (O_878,N_14766,N_14571);
or UO_879 (O_879,N_14547,N_14742);
or UO_880 (O_880,N_14586,N_14942);
or UO_881 (O_881,N_14515,N_14753);
nor UO_882 (O_882,N_14537,N_14875);
nor UO_883 (O_883,N_14533,N_14584);
and UO_884 (O_884,N_14729,N_14912);
nor UO_885 (O_885,N_14522,N_14942);
and UO_886 (O_886,N_14845,N_14678);
and UO_887 (O_887,N_14853,N_14823);
nor UO_888 (O_888,N_14688,N_14838);
nor UO_889 (O_889,N_14703,N_14566);
or UO_890 (O_890,N_14567,N_14692);
and UO_891 (O_891,N_14917,N_14617);
xnor UO_892 (O_892,N_14706,N_14931);
nand UO_893 (O_893,N_14706,N_14969);
and UO_894 (O_894,N_14509,N_14958);
nand UO_895 (O_895,N_14850,N_14594);
and UO_896 (O_896,N_14734,N_14930);
and UO_897 (O_897,N_14991,N_14944);
xnor UO_898 (O_898,N_14859,N_14657);
xor UO_899 (O_899,N_14586,N_14610);
and UO_900 (O_900,N_14814,N_14579);
and UO_901 (O_901,N_14737,N_14759);
nor UO_902 (O_902,N_14780,N_14892);
nand UO_903 (O_903,N_14656,N_14685);
or UO_904 (O_904,N_14602,N_14613);
nor UO_905 (O_905,N_14534,N_14920);
or UO_906 (O_906,N_14584,N_14922);
and UO_907 (O_907,N_14686,N_14899);
nor UO_908 (O_908,N_14857,N_14729);
and UO_909 (O_909,N_14504,N_14821);
and UO_910 (O_910,N_14800,N_14595);
and UO_911 (O_911,N_14545,N_14984);
nand UO_912 (O_912,N_14933,N_14661);
nand UO_913 (O_913,N_14549,N_14889);
or UO_914 (O_914,N_14977,N_14614);
and UO_915 (O_915,N_14546,N_14626);
nand UO_916 (O_916,N_14847,N_14615);
nor UO_917 (O_917,N_14727,N_14791);
nand UO_918 (O_918,N_14610,N_14674);
nand UO_919 (O_919,N_14857,N_14869);
or UO_920 (O_920,N_14743,N_14838);
or UO_921 (O_921,N_14849,N_14989);
nor UO_922 (O_922,N_14801,N_14844);
nor UO_923 (O_923,N_14575,N_14991);
and UO_924 (O_924,N_14854,N_14780);
nand UO_925 (O_925,N_14692,N_14817);
or UO_926 (O_926,N_14978,N_14521);
and UO_927 (O_927,N_14775,N_14570);
or UO_928 (O_928,N_14658,N_14759);
and UO_929 (O_929,N_14962,N_14550);
and UO_930 (O_930,N_14819,N_14736);
nand UO_931 (O_931,N_14906,N_14878);
nand UO_932 (O_932,N_14967,N_14995);
nand UO_933 (O_933,N_14637,N_14845);
and UO_934 (O_934,N_14633,N_14977);
nor UO_935 (O_935,N_14796,N_14616);
nor UO_936 (O_936,N_14917,N_14658);
nand UO_937 (O_937,N_14590,N_14913);
and UO_938 (O_938,N_14745,N_14890);
and UO_939 (O_939,N_14571,N_14686);
nor UO_940 (O_940,N_14555,N_14759);
nor UO_941 (O_941,N_14994,N_14825);
and UO_942 (O_942,N_14856,N_14898);
and UO_943 (O_943,N_14642,N_14561);
and UO_944 (O_944,N_14543,N_14835);
or UO_945 (O_945,N_14884,N_14608);
and UO_946 (O_946,N_14862,N_14922);
or UO_947 (O_947,N_14779,N_14749);
and UO_948 (O_948,N_14913,N_14508);
nor UO_949 (O_949,N_14660,N_14897);
and UO_950 (O_950,N_14695,N_14587);
and UO_951 (O_951,N_14530,N_14878);
nand UO_952 (O_952,N_14660,N_14611);
and UO_953 (O_953,N_14693,N_14968);
or UO_954 (O_954,N_14641,N_14694);
nand UO_955 (O_955,N_14538,N_14588);
and UO_956 (O_956,N_14754,N_14985);
nor UO_957 (O_957,N_14852,N_14737);
nor UO_958 (O_958,N_14629,N_14907);
nor UO_959 (O_959,N_14572,N_14587);
and UO_960 (O_960,N_14539,N_14542);
nand UO_961 (O_961,N_14838,N_14662);
and UO_962 (O_962,N_14510,N_14538);
and UO_963 (O_963,N_14634,N_14832);
nor UO_964 (O_964,N_14799,N_14770);
and UO_965 (O_965,N_14974,N_14801);
and UO_966 (O_966,N_14958,N_14925);
or UO_967 (O_967,N_14612,N_14806);
and UO_968 (O_968,N_14772,N_14643);
and UO_969 (O_969,N_14786,N_14949);
or UO_970 (O_970,N_14646,N_14644);
nor UO_971 (O_971,N_14555,N_14848);
or UO_972 (O_972,N_14553,N_14558);
and UO_973 (O_973,N_14636,N_14923);
nand UO_974 (O_974,N_14966,N_14618);
and UO_975 (O_975,N_14534,N_14882);
nand UO_976 (O_976,N_14868,N_14797);
and UO_977 (O_977,N_14739,N_14881);
or UO_978 (O_978,N_14932,N_14736);
and UO_979 (O_979,N_14994,N_14528);
and UO_980 (O_980,N_14826,N_14858);
nor UO_981 (O_981,N_14563,N_14945);
nor UO_982 (O_982,N_14713,N_14511);
nor UO_983 (O_983,N_14559,N_14949);
xnor UO_984 (O_984,N_14760,N_14821);
nor UO_985 (O_985,N_14750,N_14550);
or UO_986 (O_986,N_14564,N_14957);
nand UO_987 (O_987,N_14639,N_14854);
or UO_988 (O_988,N_14771,N_14794);
and UO_989 (O_989,N_14617,N_14829);
and UO_990 (O_990,N_14576,N_14641);
and UO_991 (O_991,N_14962,N_14969);
or UO_992 (O_992,N_14951,N_14530);
xor UO_993 (O_993,N_14816,N_14970);
nor UO_994 (O_994,N_14579,N_14777);
nand UO_995 (O_995,N_14861,N_14819);
or UO_996 (O_996,N_14573,N_14795);
nand UO_997 (O_997,N_14768,N_14678);
nor UO_998 (O_998,N_14866,N_14710);
nand UO_999 (O_999,N_14717,N_14507);
nor UO_1000 (O_1000,N_14907,N_14624);
nand UO_1001 (O_1001,N_14501,N_14753);
and UO_1002 (O_1002,N_14717,N_14583);
and UO_1003 (O_1003,N_14872,N_14530);
xor UO_1004 (O_1004,N_14881,N_14589);
or UO_1005 (O_1005,N_14824,N_14802);
and UO_1006 (O_1006,N_14981,N_14681);
and UO_1007 (O_1007,N_14803,N_14778);
nor UO_1008 (O_1008,N_14899,N_14844);
nor UO_1009 (O_1009,N_14720,N_14934);
nand UO_1010 (O_1010,N_14894,N_14533);
or UO_1011 (O_1011,N_14833,N_14503);
nor UO_1012 (O_1012,N_14751,N_14916);
nor UO_1013 (O_1013,N_14894,N_14854);
or UO_1014 (O_1014,N_14777,N_14903);
and UO_1015 (O_1015,N_14599,N_14769);
nand UO_1016 (O_1016,N_14711,N_14576);
xnor UO_1017 (O_1017,N_14928,N_14576);
or UO_1018 (O_1018,N_14963,N_14901);
nand UO_1019 (O_1019,N_14735,N_14989);
nand UO_1020 (O_1020,N_14777,N_14580);
and UO_1021 (O_1021,N_14685,N_14653);
and UO_1022 (O_1022,N_14607,N_14980);
xor UO_1023 (O_1023,N_14520,N_14723);
xor UO_1024 (O_1024,N_14739,N_14772);
and UO_1025 (O_1025,N_14801,N_14984);
nor UO_1026 (O_1026,N_14581,N_14882);
nand UO_1027 (O_1027,N_14674,N_14968);
nand UO_1028 (O_1028,N_14653,N_14835);
nor UO_1029 (O_1029,N_14916,N_14538);
and UO_1030 (O_1030,N_14684,N_14687);
xnor UO_1031 (O_1031,N_14524,N_14581);
nor UO_1032 (O_1032,N_14677,N_14973);
or UO_1033 (O_1033,N_14685,N_14689);
xnor UO_1034 (O_1034,N_14748,N_14522);
nand UO_1035 (O_1035,N_14676,N_14967);
nand UO_1036 (O_1036,N_14810,N_14961);
xor UO_1037 (O_1037,N_14617,N_14601);
nand UO_1038 (O_1038,N_14982,N_14529);
nor UO_1039 (O_1039,N_14676,N_14583);
or UO_1040 (O_1040,N_14626,N_14966);
and UO_1041 (O_1041,N_14921,N_14813);
nor UO_1042 (O_1042,N_14587,N_14892);
and UO_1043 (O_1043,N_14992,N_14671);
or UO_1044 (O_1044,N_14728,N_14560);
or UO_1045 (O_1045,N_14727,N_14725);
nor UO_1046 (O_1046,N_14576,N_14639);
or UO_1047 (O_1047,N_14890,N_14767);
nor UO_1048 (O_1048,N_14895,N_14888);
and UO_1049 (O_1049,N_14896,N_14873);
xor UO_1050 (O_1050,N_14733,N_14868);
nand UO_1051 (O_1051,N_14724,N_14908);
xor UO_1052 (O_1052,N_14640,N_14910);
nand UO_1053 (O_1053,N_14875,N_14583);
and UO_1054 (O_1054,N_14629,N_14926);
nand UO_1055 (O_1055,N_14626,N_14629);
and UO_1056 (O_1056,N_14763,N_14573);
nand UO_1057 (O_1057,N_14906,N_14520);
or UO_1058 (O_1058,N_14519,N_14818);
nor UO_1059 (O_1059,N_14513,N_14890);
xnor UO_1060 (O_1060,N_14734,N_14824);
nor UO_1061 (O_1061,N_14699,N_14607);
nor UO_1062 (O_1062,N_14765,N_14720);
xnor UO_1063 (O_1063,N_14830,N_14893);
nor UO_1064 (O_1064,N_14921,N_14565);
and UO_1065 (O_1065,N_14971,N_14797);
nor UO_1066 (O_1066,N_14928,N_14540);
nand UO_1067 (O_1067,N_14665,N_14736);
or UO_1068 (O_1068,N_14924,N_14727);
and UO_1069 (O_1069,N_14606,N_14897);
nor UO_1070 (O_1070,N_14876,N_14614);
or UO_1071 (O_1071,N_14865,N_14883);
nand UO_1072 (O_1072,N_14931,N_14748);
or UO_1073 (O_1073,N_14783,N_14698);
nand UO_1074 (O_1074,N_14754,N_14510);
nand UO_1075 (O_1075,N_14872,N_14915);
nand UO_1076 (O_1076,N_14509,N_14732);
xor UO_1077 (O_1077,N_14500,N_14821);
xor UO_1078 (O_1078,N_14523,N_14922);
nand UO_1079 (O_1079,N_14705,N_14692);
nand UO_1080 (O_1080,N_14562,N_14633);
nor UO_1081 (O_1081,N_14611,N_14763);
nand UO_1082 (O_1082,N_14792,N_14621);
nor UO_1083 (O_1083,N_14562,N_14564);
and UO_1084 (O_1084,N_14988,N_14814);
nand UO_1085 (O_1085,N_14935,N_14643);
or UO_1086 (O_1086,N_14793,N_14934);
and UO_1087 (O_1087,N_14519,N_14988);
or UO_1088 (O_1088,N_14601,N_14696);
nor UO_1089 (O_1089,N_14620,N_14918);
xor UO_1090 (O_1090,N_14696,N_14708);
and UO_1091 (O_1091,N_14839,N_14509);
or UO_1092 (O_1092,N_14672,N_14694);
nand UO_1093 (O_1093,N_14955,N_14621);
and UO_1094 (O_1094,N_14620,N_14953);
nand UO_1095 (O_1095,N_14917,N_14632);
and UO_1096 (O_1096,N_14556,N_14690);
or UO_1097 (O_1097,N_14648,N_14979);
nor UO_1098 (O_1098,N_14825,N_14873);
and UO_1099 (O_1099,N_14812,N_14728);
or UO_1100 (O_1100,N_14942,N_14779);
nand UO_1101 (O_1101,N_14683,N_14606);
or UO_1102 (O_1102,N_14994,N_14770);
and UO_1103 (O_1103,N_14849,N_14708);
and UO_1104 (O_1104,N_14813,N_14555);
nor UO_1105 (O_1105,N_14735,N_14705);
nand UO_1106 (O_1106,N_14728,N_14939);
nor UO_1107 (O_1107,N_14589,N_14947);
and UO_1108 (O_1108,N_14822,N_14896);
nand UO_1109 (O_1109,N_14894,N_14969);
nor UO_1110 (O_1110,N_14975,N_14991);
or UO_1111 (O_1111,N_14970,N_14632);
and UO_1112 (O_1112,N_14705,N_14711);
nor UO_1113 (O_1113,N_14522,N_14533);
and UO_1114 (O_1114,N_14801,N_14576);
nor UO_1115 (O_1115,N_14893,N_14836);
nor UO_1116 (O_1116,N_14797,N_14885);
or UO_1117 (O_1117,N_14847,N_14794);
or UO_1118 (O_1118,N_14913,N_14862);
or UO_1119 (O_1119,N_14938,N_14621);
and UO_1120 (O_1120,N_14850,N_14841);
or UO_1121 (O_1121,N_14850,N_14840);
or UO_1122 (O_1122,N_14602,N_14963);
and UO_1123 (O_1123,N_14741,N_14657);
or UO_1124 (O_1124,N_14512,N_14954);
xor UO_1125 (O_1125,N_14581,N_14787);
and UO_1126 (O_1126,N_14746,N_14576);
xor UO_1127 (O_1127,N_14574,N_14737);
nor UO_1128 (O_1128,N_14818,N_14612);
and UO_1129 (O_1129,N_14796,N_14899);
xor UO_1130 (O_1130,N_14762,N_14660);
nor UO_1131 (O_1131,N_14611,N_14615);
nand UO_1132 (O_1132,N_14757,N_14576);
or UO_1133 (O_1133,N_14523,N_14734);
nand UO_1134 (O_1134,N_14611,N_14988);
nand UO_1135 (O_1135,N_14696,N_14905);
or UO_1136 (O_1136,N_14667,N_14898);
nor UO_1137 (O_1137,N_14957,N_14667);
and UO_1138 (O_1138,N_14815,N_14914);
or UO_1139 (O_1139,N_14562,N_14604);
nand UO_1140 (O_1140,N_14759,N_14910);
xnor UO_1141 (O_1141,N_14528,N_14998);
nand UO_1142 (O_1142,N_14844,N_14854);
nand UO_1143 (O_1143,N_14829,N_14976);
and UO_1144 (O_1144,N_14637,N_14843);
or UO_1145 (O_1145,N_14856,N_14925);
and UO_1146 (O_1146,N_14661,N_14763);
or UO_1147 (O_1147,N_14696,N_14994);
nand UO_1148 (O_1148,N_14838,N_14751);
nand UO_1149 (O_1149,N_14810,N_14706);
xor UO_1150 (O_1150,N_14833,N_14916);
xnor UO_1151 (O_1151,N_14871,N_14756);
nor UO_1152 (O_1152,N_14589,N_14872);
or UO_1153 (O_1153,N_14624,N_14793);
nand UO_1154 (O_1154,N_14852,N_14721);
nor UO_1155 (O_1155,N_14807,N_14744);
nor UO_1156 (O_1156,N_14768,N_14996);
nor UO_1157 (O_1157,N_14855,N_14534);
nand UO_1158 (O_1158,N_14843,N_14813);
and UO_1159 (O_1159,N_14877,N_14816);
or UO_1160 (O_1160,N_14520,N_14593);
nor UO_1161 (O_1161,N_14753,N_14702);
and UO_1162 (O_1162,N_14831,N_14940);
nor UO_1163 (O_1163,N_14774,N_14702);
nor UO_1164 (O_1164,N_14848,N_14863);
nor UO_1165 (O_1165,N_14775,N_14870);
nand UO_1166 (O_1166,N_14502,N_14898);
and UO_1167 (O_1167,N_14540,N_14666);
or UO_1168 (O_1168,N_14731,N_14941);
xor UO_1169 (O_1169,N_14613,N_14753);
nor UO_1170 (O_1170,N_14968,N_14564);
or UO_1171 (O_1171,N_14872,N_14956);
xor UO_1172 (O_1172,N_14703,N_14814);
and UO_1173 (O_1173,N_14648,N_14518);
and UO_1174 (O_1174,N_14895,N_14545);
xnor UO_1175 (O_1175,N_14999,N_14551);
nand UO_1176 (O_1176,N_14760,N_14861);
xor UO_1177 (O_1177,N_14842,N_14595);
and UO_1178 (O_1178,N_14721,N_14573);
or UO_1179 (O_1179,N_14679,N_14887);
nor UO_1180 (O_1180,N_14596,N_14706);
nand UO_1181 (O_1181,N_14526,N_14600);
and UO_1182 (O_1182,N_14611,N_14676);
xnor UO_1183 (O_1183,N_14979,N_14666);
and UO_1184 (O_1184,N_14710,N_14623);
or UO_1185 (O_1185,N_14996,N_14752);
nand UO_1186 (O_1186,N_14942,N_14729);
nor UO_1187 (O_1187,N_14856,N_14833);
nor UO_1188 (O_1188,N_14680,N_14514);
nand UO_1189 (O_1189,N_14692,N_14633);
nor UO_1190 (O_1190,N_14644,N_14684);
xnor UO_1191 (O_1191,N_14501,N_14885);
and UO_1192 (O_1192,N_14512,N_14653);
nand UO_1193 (O_1193,N_14785,N_14680);
xnor UO_1194 (O_1194,N_14916,N_14601);
and UO_1195 (O_1195,N_14572,N_14871);
and UO_1196 (O_1196,N_14749,N_14853);
nor UO_1197 (O_1197,N_14721,N_14557);
nand UO_1198 (O_1198,N_14837,N_14540);
and UO_1199 (O_1199,N_14820,N_14561);
nor UO_1200 (O_1200,N_14544,N_14589);
nand UO_1201 (O_1201,N_14679,N_14872);
or UO_1202 (O_1202,N_14779,N_14962);
and UO_1203 (O_1203,N_14526,N_14558);
nand UO_1204 (O_1204,N_14851,N_14726);
and UO_1205 (O_1205,N_14871,N_14540);
nor UO_1206 (O_1206,N_14849,N_14514);
and UO_1207 (O_1207,N_14835,N_14861);
nor UO_1208 (O_1208,N_14917,N_14657);
nand UO_1209 (O_1209,N_14751,N_14997);
nand UO_1210 (O_1210,N_14542,N_14862);
nor UO_1211 (O_1211,N_14805,N_14500);
nor UO_1212 (O_1212,N_14858,N_14925);
or UO_1213 (O_1213,N_14633,N_14502);
or UO_1214 (O_1214,N_14870,N_14679);
xnor UO_1215 (O_1215,N_14581,N_14505);
nor UO_1216 (O_1216,N_14762,N_14941);
or UO_1217 (O_1217,N_14696,N_14615);
nor UO_1218 (O_1218,N_14888,N_14852);
xnor UO_1219 (O_1219,N_14782,N_14507);
and UO_1220 (O_1220,N_14636,N_14731);
and UO_1221 (O_1221,N_14954,N_14562);
nor UO_1222 (O_1222,N_14668,N_14695);
or UO_1223 (O_1223,N_14864,N_14767);
nor UO_1224 (O_1224,N_14768,N_14538);
or UO_1225 (O_1225,N_14826,N_14542);
nand UO_1226 (O_1226,N_14535,N_14538);
nor UO_1227 (O_1227,N_14697,N_14564);
or UO_1228 (O_1228,N_14824,N_14951);
xnor UO_1229 (O_1229,N_14680,N_14797);
nand UO_1230 (O_1230,N_14893,N_14536);
or UO_1231 (O_1231,N_14835,N_14597);
nand UO_1232 (O_1232,N_14568,N_14800);
nor UO_1233 (O_1233,N_14568,N_14613);
nand UO_1234 (O_1234,N_14643,N_14897);
nor UO_1235 (O_1235,N_14695,N_14744);
nand UO_1236 (O_1236,N_14678,N_14736);
nand UO_1237 (O_1237,N_14575,N_14838);
and UO_1238 (O_1238,N_14865,N_14949);
or UO_1239 (O_1239,N_14618,N_14744);
nor UO_1240 (O_1240,N_14538,N_14516);
or UO_1241 (O_1241,N_14938,N_14710);
nor UO_1242 (O_1242,N_14583,N_14949);
nand UO_1243 (O_1243,N_14845,N_14803);
or UO_1244 (O_1244,N_14651,N_14738);
or UO_1245 (O_1245,N_14617,N_14697);
and UO_1246 (O_1246,N_14838,N_14635);
nand UO_1247 (O_1247,N_14505,N_14752);
nor UO_1248 (O_1248,N_14710,N_14529);
nor UO_1249 (O_1249,N_14997,N_14976);
and UO_1250 (O_1250,N_14904,N_14740);
and UO_1251 (O_1251,N_14795,N_14584);
nor UO_1252 (O_1252,N_14732,N_14713);
nor UO_1253 (O_1253,N_14622,N_14848);
nor UO_1254 (O_1254,N_14955,N_14715);
or UO_1255 (O_1255,N_14799,N_14728);
or UO_1256 (O_1256,N_14672,N_14621);
or UO_1257 (O_1257,N_14709,N_14679);
nand UO_1258 (O_1258,N_14691,N_14903);
nand UO_1259 (O_1259,N_14601,N_14785);
and UO_1260 (O_1260,N_14546,N_14987);
nor UO_1261 (O_1261,N_14780,N_14805);
and UO_1262 (O_1262,N_14607,N_14971);
nor UO_1263 (O_1263,N_14712,N_14768);
nand UO_1264 (O_1264,N_14947,N_14966);
and UO_1265 (O_1265,N_14730,N_14615);
or UO_1266 (O_1266,N_14917,N_14973);
and UO_1267 (O_1267,N_14704,N_14789);
nor UO_1268 (O_1268,N_14909,N_14755);
xnor UO_1269 (O_1269,N_14862,N_14742);
or UO_1270 (O_1270,N_14794,N_14757);
xnor UO_1271 (O_1271,N_14652,N_14839);
and UO_1272 (O_1272,N_14843,N_14750);
and UO_1273 (O_1273,N_14778,N_14690);
and UO_1274 (O_1274,N_14978,N_14788);
nor UO_1275 (O_1275,N_14638,N_14775);
nor UO_1276 (O_1276,N_14599,N_14595);
and UO_1277 (O_1277,N_14568,N_14683);
and UO_1278 (O_1278,N_14626,N_14779);
nor UO_1279 (O_1279,N_14762,N_14949);
or UO_1280 (O_1280,N_14676,N_14520);
nand UO_1281 (O_1281,N_14972,N_14945);
or UO_1282 (O_1282,N_14802,N_14905);
nor UO_1283 (O_1283,N_14896,N_14748);
and UO_1284 (O_1284,N_14500,N_14583);
nor UO_1285 (O_1285,N_14912,N_14697);
nor UO_1286 (O_1286,N_14584,N_14619);
nor UO_1287 (O_1287,N_14546,N_14514);
nand UO_1288 (O_1288,N_14804,N_14997);
or UO_1289 (O_1289,N_14616,N_14748);
nor UO_1290 (O_1290,N_14532,N_14572);
nand UO_1291 (O_1291,N_14597,N_14627);
and UO_1292 (O_1292,N_14810,N_14830);
nand UO_1293 (O_1293,N_14966,N_14572);
or UO_1294 (O_1294,N_14637,N_14776);
and UO_1295 (O_1295,N_14612,N_14533);
nor UO_1296 (O_1296,N_14591,N_14742);
or UO_1297 (O_1297,N_14534,N_14649);
nor UO_1298 (O_1298,N_14529,N_14517);
xnor UO_1299 (O_1299,N_14825,N_14548);
and UO_1300 (O_1300,N_14730,N_14568);
nand UO_1301 (O_1301,N_14746,N_14644);
or UO_1302 (O_1302,N_14968,N_14892);
and UO_1303 (O_1303,N_14693,N_14641);
and UO_1304 (O_1304,N_14644,N_14908);
nor UO_1305 (O_1305,N_14952,N_14969);
xnor UO_1306 (O_1306,N_14847,N_14851);
or UO_1307 (O_1307,N_14724,N_14603);
and UO_1308 (O_1308,N_14713,N_14846);
nor UO_1309 (O_1309,N_14711,N_14678);
nor UO_1310 (O_1310,N_14810,N_14555);
and UO_1311 (O_1311,N_14541,N_14708);
nor UO_1312 (O_1312,N_14693,N_14908);
nand UO_1313 (O_1313,N_14768,N_14950);
or UO_1314 (O_1314,N_14666,N_14707);
xnor UO_1315 (O_1315,N_14622,N_14586);
or UO_1316 (O_1316,N_14683,N_14728);
nor UO_1317 (O_1317,N_14625,N_14631);
and UO_1318 (O_1318,N_14916,N_14697);
nand UO_1319 (O_1319,N_14766,N_14822);
and UO_1320 (O_1320,N_14721,N_14647);
and UO_1321 (O_1321,N_14920,N_14736);
xnor UO_1322 (O_1322,N_14557,N_14547);
or UO_1323 (O_1323,N_14615,N_14596);
and UO_1324 (O_1324,N_14528,N_14928);
nand UO_1325 (O_1325,N_14642,N_14503);
xor UO_1326 (O_1326,N_14576,N_14826);
and UO_1327 (O_1327,N_14905,N_14573);
nor UO_1328 (O_1328,N_14518,N_14631);
xnor UO_1329 (O_1329,N_14780,N_14757);
nand UO_1330 (O_1330,N_14549,N_14811);
xor UO_1331 (O_1331,N_14767,N_14875);
or UO_1332 (O_1332,N_14597,N_14652);
and UO_1333 (O_1333,N_14837,N_14757);
nor UO_1334 (O_1334,N_14882,N_14906);
nand UO_1335 (O_1335,N_14651,N_14629);
nand UO_1336 (O_1336,N_14957,N_14533);
nor UO_1337 (O_1337,N_14500,N_14634);
xor UO_1338 (O_1338,N_14609,N_14757);
nor UO_1339 (O_1339,N_14627,N_14868);
or UO_1340 (O_1340,N_14859,N_14577);
and UO_1341 (O_1341,N_14919,N_14518);
nor UO_1342 (O_1342,N_14835,N_14684);
or UO_1343 (O_1343,N_14597,N_14976);
and UO_1344 (O_1344,N_14696,N_14887);
or UO_1345 (O_1345,N_14608,N_14965);
xnor UO_1346 (O_1346,N_14519,N_14715);
and UO_1347 (O_1347,N_14883,N_14787);
and UO_1348 (O_1348,N_14686,N_14989);
or UO_1349 (O_1349,N_14799,N_14584);
and UO_1350 (O_1350,N_14934,N_14742);
xnor UO_1351 (O_1351,N_14876,N_14755);
and UO_1352 (O_1352,N_14518,N_14670);
or UO_1353 (O_1353,N_14981,N_14770);
nor UO_1354 (O_1354,N_14546,N_14689);
and UO_1355 (O_1355,N_14945,N_14600);
nor UO_1356 (O_1356,N_14641,N_14510);
nand UO_1357 (O_1357,N_14540,N_14744);
nor UO_1358 (O_1358,N_14717,N_14881);
and UO_1359 (O_1359,N_14949,N_14800);
nand UO_1360 (O_1360,N_14540,N_14631);
and UO_1361 (O_1361,N_14852,N_14806);
and UO_1362 (O_1362,N_14547,N_14537);
and UO_1363 (O_1363,N_14958,N_14989);
and UO_1364 (O_1364,N_14884,N_14697);
or UO_1365 (O_1365,N_14881,N_14902);
or UO_1366 (O_1366,N_14624,N_14616);
and UO_1367 (O_1367,N_14658,N_14813);
nand UO_1368 (O_1368,N_14668,N_14526);
and UO_1369 (O_1369,N_14816,N_14687);
nand UO_1370 (O_1370,N_14632,N_14670);
nand UO_1371 (O_1371,N_14910,N_14836);
nor UO_1372 (O_1372,N_14625,N_14932);
nor UO_1373 (O_1373,N_14721,N_14828);
nand UO_1374 (O_1374,N_14978,N_14766);
nor UO_1375 (O_1375,N_14611,N_14686);
and UO_1376 (O_1376,N_14957,N_14679);
nor UO_1377 (O_1377,N_14971,N_14748);
and UO_1378 (O_1378,N_14569,N_14647);
or UO_1379 (O_1379,N_14533,N_14682);
and UO_1380 (O_1380,N_14810,N_14540);
nand UO_1381 (O_1381,N_14990,N_14961);
nand UO_1382 (O_1382,N_14612,N_14986);
or UO_1383 (O_1383,N_14939,N_14814);
nor UO_1384 (O_1384,N_14648,N_14819);
nor UO_1385 (O_1385,N_14546,N_14910);
nor UO_1386 (O_1386,N_14727,N_14797);
xor UO_1387 (O_1387,N_14774,N_14740);
nand UO_1388 (O_1388,N_14822,N_14946);
and UO_1389 (O_1389,N_14528,N_14977);
nor UO_1390 (O_1390,N_14597,N_14697);
nor UO_1391 (O_1391,N_14544,N_14843);
nand UO_1392 (O_1392,N_14807,N_14929);
or UO_1393 (O_1393,N_14546,N_14725);
nor UO_1394 (O_1394,N_14930,N_14651);
and UO_1395 (O_1395,N_14980,N_14878);
nand UO_1396 (O_1396,N_14585,N_14668);
and UO_1397 (O_1397,N_14982,N_14801);
nand UO_1398 (O_1398,N_14716,N_14955);
or UO_1399 (O_1399,N_14893,N_14669);
or UO_1400 (O_1400,N_14774,N_14700);
or UO_1401 (O_1401,N_14722,N_14723);
or UO_1402 (O_1402,N_14990,N_14684);
nor UO_1403 (O_1403,N_14814,N_14864);
xor UO_1404 (O_1404,N_14846,N_14771);
nor UO_1405 (O_1405,N_14984,N_14977);
xor UO_1406 (O_1406,N_14783,N_14934);
nor UO_1407 (O_1407,N_14827,N_14947);
and UO_1408 (O_1408,N_14757,N_14830);
xnor UO_1409 (O_1409,N_14518,N_14748);
nor UO_1410 (O_1410,N_14960,N_14780);
and UO_1411 (O_1411,N_14987,N_14832);
nand UO_1412 (O_1412,N_14819,N_14554);
xor UO_1413 (O_1413,N_14806,N_14559);
or UO_1414 (O_1414,N_14700,N_14954);
nand UO_1415 (O_1415,N_14997,N_14503);
or UO_1416 (O_1416,N_14898,N_14868);
nor UO_1417 (O_1417,N_14913,N_14968);
xor UO_1418 (O_1418,N_14783,N_14997);
nor UO_1419 (O_1419,N_14617,N_14595);
or UO_1420 (O_1420,N_14816,N_14657);
nand UO_1421 (O_1421,N_14801,N_14607);
and UO_1422 (O_1422,N_14800,N_14924);
or UO_1423 (O_1423,N_14751,N_14667);
nand UO_1424 (O_1424,N_14798,N_14917);
or UO_1425 (O_1425,N_14670,N_14602);
nor UO_1426 (O_1426,N_14802,N_14605);
and UO_1427 (O_1427,N_14745,N_14512);
nand UO_1428 (O_1428,N_14847,N_14952);
and UO_1429 (O_1429,N_14928,N_14624);
nor UO_1430 (O_1430,N_14555,N_14548);
nand UO_1431 (O_1431,N_14813,N_14935);
or UO_1432 (O_1432,N_14860,N_14922);
nor UO_1433 (O_1433,N_14642,N_14857);
nand UO_1434 (O_1434,N_14942,N_14907);
nand UO_1435 (O_1435,N_14801,N_14557);
and UO_1436 (O_1436,N_14664,N_14725);
xnor UO_1437 (O_1437,N_14978,N_14646);
or UO_1438 (O_1438,N_14759,N_14878);
or UO_1439 (O_1439,N_14701,N_14580);
nand UO_1440 (O_1440,N_14759,N_14774);
nand UO_1441 (O_1441,N_14668,N_14575);
or UO_1442 (O_1442,N_14983,N_14746);
nand UO_1443 (O_1443,N_14788,N_14814);
nand UO_1444 (O_1444,N_14964,N_14501);
or UO_1445 (O_1445,N_14741,N_14544);
nand UO_1446 (O_1446,N_14817,N_14804);
and UO_1447 (O_1447,N_14971,N_14556);
nor UO_1448 (O_1448,N_14583,N_14668);
nor UO_1449 (O_1449,N_14999,N_14852);
nor UO_1450 (O_1450,N_14749,N_14724);
and UO_1451 (O_1451,N_14881,N_14531);
xor UO_1452 (O_1452,N_14533,N_14585);
and UO_1453 (O_1453,N_14669,N_14696);
and UO_1454 (O_1454,N_14546,N_14844);
or UO_1455 (O_1455,N_14994,N_14823);
and UO_1456 (O_1456,N_14952,N_14766);
and UO_1457 (O_1457,N_14608,N_14810);
nor UO_1458 (O_1458,N_14508,N_14764);
nand UO_1459 (O_1459,N_14758,N_14947);
nor UO_1460 (O_1460,N_14653,N_14748);
or UO_1461 (O_1461,N_14614,N_14660);
nand UO_1462 (O_1462,N_14767,N_14601);
nor UO_1463 (O_1463,N_14763,N_14785);
xor UO_1464 (O_1464,N_14933,N_14768);
or UO_1465 (O_1465,N_14575,N_14712);
nor UO_1466 (O_1466,N_14789,N_14787);
xor UO_1467 (O_1467,N_14885,N_14730);
xnor UO_1468 (O_1468,N_14582,N_14597);
nand UO_1469 (O_1469,N_14541,N_14778);
and UO_1470 (O_1470,N_14674,N_14969);
nand UO_1471 (O_1471,N_14673,N_14689);
nor UO_1472 (O_1472,N_14629,N_14663);
and UO_1473 (O_1473,N_14544,N_14500);
and UO_1474 (O_1474,N_14942,N_14947);
xnor UO_1475 (O_1475,N_14836,N_14699);
or UO_1476 (O_1476,N_14919,N_14541);
and UO_1477 (O_1477,N_14988,N_14926);
or UO_1478 (O_1478,N_14680,N_14840);
or UO_1479 (O_1479,N_14602,N_14923);
and UO_1480 (O_1480,N_14956,N_14852);
or UO_1481 (O_1481,N_14840,N_14990);
and UO_1482 (O_1482,N_14864,N_14761);
nand UO_1483 (O_1483,N_14648,N_14745);
and UO_1484 (O_1484,N_14783,N_14737);
and UO_1485 (O_1485,N_14965,N_14995);
or UO_1486 (O_1486,N_14769,N_14999);
or UO_1487 (O_1487,N_14645,N_14756);
and UO_1488 (O_1488,N_14501,N_14613);
and UO_1489 (O_1489,N_14701,N_14679);
or UO_1490 (O_1490,N_14702,N_14927);
nand UO_1491 (O_1491,N_14953,N_14701);
nor UO_1492 (O_1492,N_14763,N_14621);
nor UO_1493 (O_1493,N_14712,N_14931);
and UO_1494 (O_1494,N_14670,N_14869);
nand UO_1495 (O_1495,N_14847,N_14986);
nor UO_1496 (O_1496,N_14712,N_14922);
and UO_1497 (O_1497,N_14838,N_14558);
and UO_1498 (O_1498,N_14955,N_14974);
nand UO_1499 (O_1499,N_14508,N_14811);
nor UO_1500 (O_1500,N_14595,N_14834);
or UO_1501 (O_1501,N_14705,N_14541);
nor UO_1502 (O_1502,N_14854,N_14615);
nor UO_1503 (O_1503,N_14778,N_14990);
or UO_1504 (O_1504,N_14500,N_14956);
nor UO_1505 (O_1505,N_14831,N_14854);
and UO_1506 (O_1506,N_14845,N_14645);
nand UO_1507 (O_1507,N_14653,N_14725);
nor UO_1508 (O_1508,N_14758,N_14854);
or UO_1509 (O_1509,N_14784,N_14717);
and UO_1510 (O_1510,N_14815,N_14827);
nor UO_1511 (O_1511,N_14871,N_14555);
nor UO_1512 (O_1512,N_14813,N_14561);
xor UO_1513 (O_1513,N_14668,N_14705);
or UO_1514 (O_1514,N_14519,N_14925);
nor UO_1515 (O_1515,N_14519,N_14955);
nor UO_1516 (O_1516,N_14762,N_14899);
nand UO_1517 (O_1517,N_14940,N_14514);
and UO_1518 (O_1518,N_14679,N_14732);
and UO_1519 (O_1519,N_14893,N_14657);
nand UO_1520 (O_1520,N_14998,N_14556);
nand UO_1521 (O_1521,N_14603,N_14660);
nor UO_1522 (O_1522,N_14679,N_14877);
nand UO_1523 (O_1523,N_14514,N_14662);
nor UO_1524 (O_1524,N_14797,N_14577);
xor UO_1525 (O_1525,N_14787,N_14900);
nor UO_1526 (O_1526,N_14518,N_14936);
and UO_1527 (O_1527,N_14827,N_14952);
or UO_1528 (O_1528,N_14632,N_14551);
or UO_1529 (O_1529,N_14610,N_14508);
nor UO_1530 (O_1530,N_14567,N_14798);
nor UO_1531 (O_1531,N_14651,N_14986);
and UO_1532 (O_1532,N_14754,N_14961);
and UO_1533 (O_1533,N_14851,N_14592);
nor UO_1534 (O_1534,N_14537,N_14630);
or UO_1535 (O_1535,N_14533,N_14902);
xor UO_1536 (O_1536,N_14563,N_14941);
or UO_1537 (O_1537,N_14981,N_14528);
nor UO_1538 (O_1538,N_14691,N_14768);
xnor UO_1539 (O_1539,N_14952,N_14646);
or UO_1540 (O_1540,N_14798,N_14812);
and UO_1541 (O_1541,N_14647,N_14990);
nand UO_1542 (O_1542,N_14510,N_14576);
and UO_1543 (O_1543,N_14601,N_14594);
nand UO_1544 (O_1544,N_14700,N_14871);
and UO_1545 (O_1545,N_14735,N_14819);
and UO_1546 (O_1546,N_14897,N_14945);
and UO_1547 (O_1547,N_14857,N_14949);
or UO_1548 (O_1548,N_14610,N_14800);
and UO_1549 (O_1549,N_14748,N_14586);
nand UO_1550 (O_1550,N_14974,N_14645);
or UO_1551 (O_1551,N_14818,N_14530);
nand UO_1552 (O_1552,N_14754,N_14976);
nand UO_1553 (O_1553,N_14597,N_14514);
and UO_1554 (O_1554,N_14553,N_14514);
and UO_1555 (O_1555,N_14841,N_14732);
nand UO_1556 (O_1556,N_14783,N_14883);
nand UO_1557 (O_1557,N_14831,N_14900);
nor UO_1558 (O_1558,N_14611,N_14606);
nand UO_1559 (O_1559,N_14923,N_14514);
and UO_1560 (O_1560,N_14659,N_14835);
and UO_1561 (O_1561,N_14939,N_14805);
or UO_1562 (O_1562,N_14598,N_14602);
nand UO_1563 (O_1563,N_14937,N_14542);
and UO_1564 (O_1564,N_14858,N_14904);
nor UO_1565 (O_1565,N_14519,N_14833);
nor UO_1566 (O_1566,N_14501,N_14512);
or UO_1567 (O_1567,N_14532,N_14615);
or UO_1568 (O_1568,N_14557,N_14810);
nor UO_1569 (O_1569,N_14526,N_14887);
and UO_1570 (O_1570,N_14808,N_14845);
and UO_1571 (O_1571,N_14803,N_14609);
nand UO_1572 (O_1572,N_14740,N_14788);
xor UO_1573 (O_1573,N_14610,N_14697);
nand UO_1574 (O_1574,N_14621,N_14841);
nand UO_1575 (O_1575,N_14953,N_14732);
and UO_1576 (O_1576,N_14951,N_14908);
and UO_1577 (O_1577,N_14536,N_14671);
and UO_1578 (O_1578,N_14939,N_14638);
or UO_1579 (O_1579,N_14539,N_14864);
and UO_1580 (O_1580,N_14549,N_14830);
nor UO_1581 (O_1581,N_14676,N_14927);
and UO_1582 (O_1582,N_14543,N_14512);
and UO_1583 (O_1583,N_14860,N_14861);
or UO_1584 (O_1584,N_14754,N_14540);
and UO_1585 (O_1585,N_14786,N_14731);
and UO_1586 (O_1586,N_14523,N_14699);
nand UO_1587 (O_1587,N_14698,N_14867);
or UO_1588 (O_1588,N_14709,N_14778);
and UO_1589 (O_1589,N_14956,N_14767);
xor UO_1590 (O_1590,N_14502,N_14521);
nor UO_1591 (O_1591,N_14885,N_14930);
nand UO_1592 (O_1592,N_14651,N_14799);
nand UO_1593 (O_1593,N_14885,N_14717);
nor UO_1594 (O_1594,N_14928,N_14729);
nor UO_1595 (O_1595,N_14668,N_14898);
nand UO_1596 (O_1596,N_14553,N_14778);
and UO_1597 (O_1597,N_14528,N_14797);
or UO_1598 (O_1598,N_14977,N_14890);
or UO_1599 (O_1599,N_14695,N_14958);
nor UO_1600 (O_1600,N_14744,N_14711);
xor UO_1601 (O_1601,N_14777,N_14684);
xnor UO_1602 (O_1602,N_14619,N_14816);
nor UO_1603 (O_1603,N_14712,N_14802);
nand UO_1604 (O_1604,N_14974,N_14710);
nand UO_1605 (O_1605,N_14612,N_14617);
and UO_1606 (O_1606,N_14737,N_14978);
nand UO_1607 (O_1607,N_14527,N_14929);
nand UO_1608 (O_1608,N_14928,N_14732);
nor UO_1609 (O_1609,N_14777,N_14576);
nand UO_1610 (O_1610,N_14516,N_14549);
or UO_1611 (O_1611,N_14752,N_14891);
xnor UO_1612 (O_1612,N_14527,N_14750);
nor UO_1613 (O_1613,N_14622,N_14897);
nor UO_1614 (O_1614,N_14996,N_14834);
xor UO_1615 (O_1615,N_14521,N_14781);
xnor UO_1616 (O_1616,N_14922,N_14881);
xor UO_1617 (O_1617,N_14921,N_14801);
nand UO_1618 (O_1618,N_14969,N_14861);
nand UO_1619 (O_1619,N_14758,N_14845);
nor UO_1620 (O_1620,N_14559,N_14719);
nor UO_1621 (O_1621,N_14642,N_14838);
nand UO_1622 (O_1622,N_14951,N_14963);
nor UO_1623 (O_1623,N_14548,N_14620);
nand UO_1624 (O_1624,N_14834,N_14920);
nand UO_1625 (O_1625,N_14631,N_14884);
nand UO_1626 (O_1626,N_14813,N_14585);
or UO_1627 (O_1627,N_14816,N_14638);
xnor UO_1628 (O_1628,N_14823,N_14873);
and UO_1629 (O_1629,N_14602,N_14538);
or UO_1630 (O_1630,N_14950,N_14836);
or UO_1631 (O_1631,N_14553,N_14988);
nand UO_1632 (O_1632,N_14655,N_14647);
or UO_1633 (O_1633,N_14733,N_14559);
nor UO_1634 (O_1634,N_14857,N_14926);
and UO_1635 (O_1635,N_14563,N_14939);
nor UO_1636 (O_1636,N_14980,N_14775);
and UO_1637 (O_1637,N_14888,N_14974);
or UO_1638 (O_1638,N_14573,N_14954);
nand UO_1639 (O_1639,N_14899,N_14760);
xnor UO_1640 (O_1640,N_14762,N_14806);
and UO_1641 (O_1641,N_14961,N_14730);
xor UO_1642 (O_1642,N_14557,N_14700);
and UO_1643 (O_1643,N_14538,N_14771);
nor UO_1644 (O_1644,N_14669,N_14751);
nand UO_1645 (O_1645,N_14634,N_14567);
and UO_1646 (O_1646,N_14689,N_14659);
nand UO_1647 (O_1647,N_14861,N_14588);
or UO_1648 (O_1648,N_14642,N_14609);
nor UO_1649 (O_1649,N_14689,N_14962);
and UO_1650 (O_1650,N_14832,N_14630);
nand UO_1651 (O_1651,N_14655,N_14806);
nand UO_1652 (O_1652,N_14613,N_14646);
xnor UO_1653 (O_1653,N_14636,N_14569);
or UO_1654 (O_1654,N_14876,N_14518);
nand UO_1655 (O_1655,N_14568,N_14838);
or UO_1656 (O_1656,N_14719,N_14706);
nor UO_1657 (O_1657,N_14873,N_14572);
and UO_1658 (O_1658,N_14500,N_14751);
nor UO_1659 (O_1659,N_14769,N_14713);
nand UO_1660 (O_1660,N_14850,N_14564);
nor UO_1661 (O_1661,N_14712,N_14573);
or UO_1662 (O_1662,N_14852,N_14941);
or UO_1663 (O_1663,N_14770,N_14940);
or UO_1664 (O_1664,N_14977,N_14736);
and UO_1665 (O_1665,N_14955,N_14889);
or UO_1666 (O_1666,N_14787,N_14668);
and UO_1667 (O_1667,N_14737,N_14732);
nand UO_1668 (O_1668,N_14793,N_14883);
nor UO_1669 (O_1669,N_14593,N_14531);
and UO_1670 (O_1670,N_14832,N_14705);
nor UO_1671 (O_1671,N_14735,N_14500);
and UO_1672 (O_1672,N_14892,N_14901);
and UO_1673 (O_1673,N_14728,N_14876);
nor UO_1674 (O_1674,N_14906,N_14700);
nand UO_1675 (O_1675,N_14709,N_14590);
nand UO_1676 (O_1676,N_14924,N_14763);
and UO_1677 (O_1677,N_14905,N_14764);
or UO_1678 (O_1678,N_14883,N_14673);
nor UO_1679 (O_1679,N_14687,N_14554);
and UO_1680 (O_1680,N_14810,N_14866);
and UO_1681 (O_1681,N_14863,N_14852);
nor UO_1682 (O_1682,N_14674,N_14711);
nor UO_1683 (O_1683,N_14967,N_14598);
xor UO_1684 (O_1684,N_14975,N_14972);
xor UO_1685 (O_1685,N_14522,N_14827);
and UO_1686 (O_1686,N_14939,N_14531);
xnor UO_1687 (O_1687,N_14904,N_14791);
nand UO_1688 (O_1688,N_14595,N_14968);
nand UO_1689 (O_1689,N_14556,N_14505);
or UO_1690 (O_1690,N_14942,N_14697);
and UO_1691 (O_1691,N_14545,N_14969);
or UO_1692 (O_1692,N_14550,N_14666);
or UO_1693 (O_1693,N_14760,N_14784);
nor UO_1694 (O_1694,N_14596,N_14796);
and UO_1695 (O_1695,N_14500,N_14730);
or UO_1696 (O_1696,N_14833,N_14966);
nor UO_1697 (O_1697,N_14819,N_14701);
or UO_1698 (O_1698,N_14690,N_14897);
or UO_1699 (O_1699,N_14682,N_14885);
nor UO_1700 (O_1700,N_14715,N_14779);
nor UO_1701 (O_1701,N_14798,N_14641);
and UO_1702 (O_1702,N_14849,N_14580);
or UO_1703 (O_1703,N_14906,N_14716);
and UO_1704 (O_1704,N_14667,N_14624);
and UO_1705 (O_1705,N_14725,N_14797);
and UO_1706 (O_1706,N_14554,N_14620);
and UO_1707 (O_1707,N_14679,N_14538);
or UO_1708 (O_1708,N_14938,N_14652);
xnor UO_1709 (O_1709,N_14663,N_14897);
xnor UO_1710 (O_1710,N_14982,N_14785);
and UO_1711 (O_1711,N_14587,N_14748);
nand UO_1712 (O_1712,N_14680,N_14658);
nor UO_1713 (O_1713,N_14932,N_14811);
nor UO_1714 (O_1714,N_14907,N_14704);
nor UO_1715 (O_1715,N_14582,N_14951);
and UO_1716 (O_1716,N_14923,N_14955);
nand UO_1717 (O_1717,N_14736,N_14940);
or UO_1718 (O_1718,N_14931,N_14702);
xor UO_1719 (O_1719,N_14528,N_14651);
or UO_1720 (O_1720,N_14670,N_14551);
nor UO_1721 (O_1721,N_14748,N_14961);
xor UO_1722 (O_1722,N_14577,N_14670);
nand UO_1723 (O_1723,N_14772,N_14650);
or UO_1724 (O_1724,N_14869,N_14506);
and UO_1725 (O_1725,N_14919,N_14558);
nand UO_1726 (O_1726,N_14600,N_14954);
and UO_1727 (O_1727,N_14584,N_14906);
or UO_1728 (O_1728,N_14752,N_14923);
or UO_1729 (O_1729,N_14575,N_14733);
and UO_1730 (O_1730,N_14759,N_14701);
and UO_1731 (O_1731,N_14781,N_14754);
nand UO_1732 (O_1732,N_14660,N_14696);
xor UO_1733 (O_1733,N_14674,N_14667);
nor UO_1734 (O_1734,N_14541,N_14969);
nor UO_1735 (O_1735,N_14972,N_14748);
and UO_1736 (O_1736,N_14628,N_14747);
and UO_1737 (O_1737,N_14652,N_14722);
and UO_1738 (O_1738,N_14721,N_14542);
xnor UO_1739 (O_1739,N_14574,N_14895);
nand UO_1740 (O_1740,N_14591,N_14528);
and UO_1741 (O_1741,N_14860,N_14640);
and UO_1742 (O_1742,N_14519,N_14651);
and UO_1743 (O_1743,N_14800,N_14970);
and UO_1744 (O_1744,N_14666,N_14521);
and UO_1745 (O_1745,N_14528,N_14563);
and UO_1746 (O_1746,N_14879,N_14817);
nand UO_1747 (O_1747,N_14525,N_14634);
or UO_1748 (O_1748,N_14797,N_14936);
or UO_1749 (O_1749,N_14899,N_14707);
nand UO_1750 (O_1750,N_14908,N_14519);
and UO_1751 (O_1751,N_14772,N_14553);
nand UO_1752 (O_1752,N_14950,N_14555);
xor UO_1753 (O_1753,N_14779,N_14586);
nor UO_1754 (O_1754,N_14768,N_14916);
or UO_1755 (O_1755,N_14836,N_14807);
or UO_1756 (O_1756,N_14507,N_14987);
nor UO_1757 (O_1757,N_14685,N_14762);
nand UO_1758 (O_1758,N_14876,N_14665);
nand UO_1759 (O_1759,N_14990,N_14565);
xnor UO_1760 (O_1760,N_14808,N_14557);
nand UO_1761 (O_1761,N_14882,N_14819);
and UO_1762 (O_1762,N_14952,N_14981);
nor UO_1763 (O_1763,N_14824,N_14576);
nand UO_1764 (O_1764,N_14910,N_14694);
nor UO_1765 (O_1765,N_14547,N_14579);
or UO_1766 (O_1766,N_14851,N_14666);
nor UO_1767 (O_1767,N_14877,N_14536);
or UO_1768 (O_1768,N_14654,N_14544);
xor UO_1769 (O_1769,N_14900,N_14854);
and UO_1770 (O_1770,N_14868,N_14545);
and UO_1771 (O_1771,N_14990,N_14595);
and UO_1772 (O_1772,N_14993,N_14795);
or UO_1773 (O_1773,N_14863,N_14566);
or UO_1774 (O_1774,N_14849,N_14788);
and UO_1775 (O_1775,N_14759,N_14594);
or UO_1776 (O_1776,N_14918,N_14959);
nand UO_1777 (O_1777,N_14516,N_14700);
or UO_1778 (O_1778,N_14661,N_14535);
and UO_1779 (O_1779,N_14560,N_14925);
nand UO_1780 (O_1780,N_14698,N_14609);
nor UO_1781 (O_1781,N_14518,N_14720);
nor UO_1782 (O_1782,N_14680,N_14958);
nand UO_1783 (O_1783,N_14665,N_14705);
and UO_1784 (O_1784,N_14837,N_14517);
and UO_1785 (O_1785,N_14827,N_14838);
and UO_1786 (O_1786,N_14930,N_14619);
and UO_1787 (O_1787,N_14714,N_14808);
nor UO_1788 (O_1788,N_14621,N_14979);
nand UO_1789 (O_1789,N_14790,N_14747);
nand UO_1790 (O_1790,N_14776,N_14707);
nand UO_1791 (O_1791,N_14848,N_14613);
or UO_1792 (O_1792,N_14576,N_14834);
or UO_1793 (O_1793,N_14550,N_14720);
xnor UO_1794 (O_1794,N_14618,N_14678);
and UO_1795 (O_1795,N_14860,N_14828);
or UO_1796 (O_1796,N_14542,N_14799);
nand UO_1797 (O_1797,N_14813,N_14881);
or UO_1798 (O_1798,N_14676,N_14892);
nand UO_1799 (O_1799,N_14914,N_14814);
nand UO_1800 (O_1800,N_14736,N_14947);
nor UO_1801 (O_1801,N_14761,N_14917);
xor UO_1802 (O_1802,N_14894,N_14675);
or UO_1803 (O_1803,N_14844,N_14528);
or UO_1804 (O_1804,N_14644,N_14698);
or UO_1805 (O_1805,N_14860,N_14680);
nor UO_1806 (O_1806,N_14829,N_14929);
or UO_1807 (O_1807,N_14881,N_14606);
nor UO_1808 (O_1808,N_14601,N_14709);
nor UO_1809 (O_1809,N_14570,N_14854);
xor UO_1810 (O_1810,N_14974,N_14659);
nor UO_1811 (O_1811,N_14895,N_14793);
xor UO_1812 (O_1812,N_14934,N_14740);
xnor UO_1813 (O_1813,N_14982,N_14926);
nor UO_1814 (O_1814,N_14821,N_14763);
nor UO_1815 (O_1815,N_14677,N_14829);
nand UO_1816 (O_1816,N_14899,N_14698);
or UO_1817 (O_1817,N_14915,N_14767);
and UO_1818 (O_1818,N_14836,N_14663);
and UO_1819 (O_1819,N_14880,N_14672);
or UO_1820 (O_1820,N_14899,N_14818);
and UO_1821 (O_1821,N_14547,N_14684);
and UO_1822 (O_1822,N_14704,N_14829);
nand UO_1823 (O_1823,N_14711,N_14735);
and UO_1824 (O_1824,N_14634,N_14890);
xor UO_1825 (O_1825,N_14601,N_14589);
or UO_1826 (O_1826,N_14650,N_14770);
nor UO_1827 (O_1827,N_14901,N_14898);
xnor UO_1828 (O_1828,N_14707,N_14965);
or UO_1829 (O_1829,N_14791,N_14566);
and UO_1830 (O_1830,N_14690,N_14853);
nor UO_1831 (O_1831,N_14961,N_14673);
or UO_1832 (O_1832,N_14749,N_14988);
nand UO_1833 (O_1833,N_14706,N_14639);
or UO_1834 (O_1834,N_14882,N_14593);
and UO_1835 (O_1835,N_14634,N_14593);
and UO_1836 (O_1836,N_14624,N_14700);
and UO_1837 (O_1837,N_14965,N_14791);
nand UO_1838 (O_1838,N_14712,N_14873);
nor UO_1839 (O_1839,N_14738,N_14695);
or UO_1840 (O_1840,N_14612,N_14994);
nor UO_1841 (O_1841,N_14731,N_14518);
nand UO_1842 (O_1842,N_14514,N_14583);
nand UO_1843 (O_1843,N_14620,N_14831);
and UO_1844 (O_1844,N_14740,N_14916);
nor UO_1845 (O_1845,N_14571,N_14882);
and UO_1846 (O_1846,N_14835,N_14648);
or UO_1847 (O_1847,N_14852,N_14552);
and UO_1848 (O_1848,N_14861,N_14968);
or UO_1849 (O_1849,N_14501,N_14721);
or UO_1850 (O_1850,N_14601,N_14582);
nor UO_1851 (O_1851,N_14624,N_14904);
nor UO_1852 (O_1852,N_14613,N_14708);
xnor UO_1853 (O_1853,N_14815,N_14785);
nand UO_1854 (O_1854,N_14666,N_14671);
or UO_1855 (O_1855,N_14828,N_14836);
and UO_1856 (O_1856,N_14764,N_14691);
nor UO_1857 (O_1857,N_14878,N_14979);
and UO_1858 (O_1858,N_14909,N_14997);
and UO_1859 (O_1859,N_14749,N_14742);
nor UO_1860 (O_1860,N_14522,N_14969);
or UO_1861 (O_1861,N_14724,N_14772);
nand UO_1862 (O_1862,N_14656,N_14547);
and UO_1863 (O_1863,N_14769,N_14749);
nand UO_1864 (O_1864,N_14887,N_14535);
nor UO_1865 (O_1865,N_14837,N_14978);
and UO_1866 (O_1866,N_14542,N_14884);
or UO_1867 (O_1867,N_14909,N_14591);
nor UO_1868 (O_1868,N_14968,N_14589);
nor UO_1869 (O_1869,N_14685,N_14787);
xnor UO_1870 (O_1870,N_14790,N_14678);
and UO_1871 (O_1871,N_14505,N_14559);
nand UO_1872 (O_1872,N_14663,N_14985);
nand UO_1873 (O_1873,N_14743,N_14775);
and UO_1874 (O_1874,N_14928,N_14558);
or UO_1875 (O_1875,N_14937,N_14953);
or UO_1876 (O_1876,N_14841,N_14639);
nand UO_1877 (O_1877,N_14674,N_14877);
or UO_1878 (O_1878,N_14732,N_14523);
nand UO_1879 (O_1879,N_14528,N_14984);
nor UO_1880 (O_1880,N_14677,N_14818);
and UO_1881 (O_1881,N_14580,N_14973);
nand UO_1882 (O_1882,N_14664,N_14686);
xor UO_1883 (O_1883,N_14732,N_14817);
nand UO_1884 (O_1884,N_14813,N_14805);
xnor UO_1885 (O_1885,N_14990,N_14983);
nor UO_1886 (O_1886,N_14753,N_14662);
nor UO_1887 (O_1887,N_14827,N_14569);
nor UO_1888 (O_1888,N_14667,N_14999);
or UO_1889 (O_1889,N_14890,N_14965);
nand UO_1890 (O_1890,N_14838,N_14610);
nand UO_1891 (O_1891,N_14597,N_14663);
and UO_1892 (O_1892,N_14895,N_14837);
or UO_1893 (O_1893,N_14960,N_14975);
nand UO_1894 (O_1894,N_14536,N_14883);
nand UO_1895 (O_1895,N_14991,N_14930);
and UO_1896 (O_1896,N_14812,N_14617);
nor UO_1897 (O_1897,N_14613,N_14507);
nand UO_1898 (O_1898,N_14688,N_14593);
nor UO_1899 (O_1899,N_14970,N_14538);
nand UO_1900 (O_1900,N_14942,N_14679);
nor UO_1901 (O_1901,N_14724,N_14853);
or UO_1902 (O_1902,N_14931,N_14885);
nand UO_1903 (O_1903,N_14888,N_14905);
and UO_1904 (O_1904,N_14510,N_14965);
or UO_1905 (O_1905,N_14633,N_14723);
xor UO_1906 (O_1906,N_14678,N_14624);
nand UO_1907 (O_1907,N_14539,N_14978);
nor UO_1908 (O_1908,N_14529,N_14613);
xor UO_1909 (O_1909,N_14640,N_14848);
nor UO_1910 (O_1910,N_14816,N_14951);
nand UO_1911 (O_1911,N_14522,N_14652);
nor UO_1912 (O_1912,N_14579,N_14816);
nand UO_1913 (O_1913,N_14839,N_14979);
and UO_1914 (O_1914,N_14915,N_14569);
or UO_1915 (O_1915,N_14874,N_14785);
or UO_1916 (O_1916,N_14792,N_14706);
nand UO_1917 (O_1917,N_14778,N_14670);
nor UO_1918 (O_1918,N_14792,N_14927);
and UO_1919 (O_1919,N_14598,N_14914);
and UO_1920 (O_1920,N_14523,N_14961);
and UO_1921 (O_1921,N_14975,N_14736);
or UO_1922 (O_1922,N_14646,N_14741);
nor UO_1923 (O_1923,N_14998,N_14610);
and UO_1924 (O_1924,N_14883,N_14570);
nor UO_1925 (O_1925,N_14760,N_14935);
nand UO_1926 (O_1926,N_14835,N_14685);
nor UO_1927 (O_1927,N_14928,N_14508);
xnor UO_1928 (O_1928,N_14682,N_14750);
and UO_1929 (O_1929,N_14772,N_14597);
nand UO_1930 (O_1930,N_14501,N_14968);
nand UO_1931 (O_1931,N_14634,N_14844);
xor UO_1932 (O_1932,N_14911,N_14646);
or UO_1933 (O_1933,N_14954,N_14534);
nor UO_1934 (O_1934,N_14715,N_14657);
and UO_1935 (O_1935,N_14588,N_14877);
nor UO_1936 (O_1936,N_14999,N_14545);
or UO_1937 (O_1937,N_14784,N_14947);
xnor UO_1938 (O_1938,N_14628,N_14558);
nand UO_1939 (O_1939,N_14655,N_14948);
and UO_1940 (O_1940,N_14881,N_14634);
nor UO_1941 (O_1941,N_14661,N_14815);
and UO_1942 (O_1942,N_14622,N_14711);
or UO_1943 (O_1943,N_14721,N_14997);
nor UO_1944 (O_1944,N_14973,N_14536);
xor UO_1945 (O_1945,N_14649,N_14846);
nand UO_1946 (O_1946,N_14536,N_14966);
and UO_1947 (O_1947,N_14592,N_14742);
and UO_1948 (O_1948,N_14629,N_14822);
and UO_1949 (O_1949,N_14516,N_14725);
xnor UO_1950 (O_1950,N_14602,N_14586);
and UO_1951 (O_1951,N_14944,N_14518);
and UO_1952 (O_1952,N_14643,N_14703);
xor UO_1953 (O_1953,N_14723,N_14762);
nor UO_1954 (O_1954,N_14976,N_14870);
or UO_1955 (O_1955,N_14502,N_14976);
nor UO_1956 (O_1956,N_14697,N_14797);
and UO_1957 (O_1957,N_14869,N_14847);
or UO_1958 (O_1958,N_14619,N_14712);
nor UO_1959 (O_1959,N_14938,N_14666);
nor UO_1960 (O_1960,N_14957,N_14868);
and UO_1961 (O_1961,N_14625,N_14867);
or UO_1962 (O_1962,N_14751,N_14517);
nor UO_1963 (O_1963,N_14680,N_14671);
and UO_1964 (O_1964,N_14949,N_14930);
nand UO_1965 (O_1965,N_14747,N_14545);
and UO_1966 (O_1966,N_14935,N_14904);
nor UO_1967 (O_1967,N_14981,N_14609);
and UO_1968 (O_1968,N_14914,N_14778);
or UO_1969 (O_1969,N_14805,N_14831);
nor UO_1970 (O_1970,N_14869,N_14550);
or UO_1971 (O_1971,N_14718,N_14849);
and UO_1972 (O_1972,N_14857,N_14807);
and UO_1973 (O_1973,N_14700,N_14770);
and UO_1974 (O_1974,N_14583,N_14862);
or UO_1975 (O_1975,N_14874,N_14755);
or UO_1976 (O_1976,N_14817,N_14744);
and UO_1977 (O_1977,N_14709,N_14802);
nand UO_1978 (O_1978,N_14594,N_14684);
nand UO_1979 (O_1979,N_14979,N_14547);
nor UO_1980 (O_1980,N_14956,N_14657);
nand UO_1981 (O_1981,N_14729,N_14714);
and UO_1982 (O_1982,N_14595,N_14774);
or UO_1983 (O_1983,N_14782,N_14725);
nor UO_1984 (O_1984,N_14516,N_14534);
nor UO_1985 (O_1985,N_14815,N_14776);
xor UO_1986 (O_1986,N_14746,N_14565);
or UO_1987 (O_1987,N_14822,N_14956);
nor UO_1988 (O_1988,N_14912,N_14889);
nand UO_1989 (O_1989,N_14667,N_14585);
and UO_1990 (O_1990,N_14934,N_14944);
nand UO_1991 (O_1991,N_14807,N_14801);
nand UO_1992 (O_1992,N_14529,N_14553);
nand UO_1993 (O_1993,N_14746,N_14845);
or UO_1994 (O_1994,N_14517,N_14831);
or UO_1995 (O_1995,N_14907,N_14993);
xor UO_1996 (O_1996,N_14515,N_14517);
xnor UO_1997 (O_1997,N_14787,N_14724);
nand UO_1998 (O_1998,N_14612,N_14851);
and UO_1999 (O_1999,N_14896,N_14893);
endmodule