module basic_500_3000_500_4_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xor U0 (N_0,In_172,In_264);
nor U1 (N_1,In_150,In_140);
nand U2 (N_2,In_194,In_201);
and U3 (N_3,In_432,In_22);
nor U4 (N_4,In_281,In_436);
nand U5 (N_5,In_0,In_441);
and U6 (N_6,In_202,In_420);
nor U7 (N_7,In_303,In_120);
or U8 (N_8,In_402,In_474);
nand U9 (N_9,In_372,In_380);
nand U10 (N_10,In_57,In_289);
nand U11 (N_11,In_349,In_215);
and U12 (N_12,In_255,In_62);
or U13 (N_13,In_142,In_195);
nor U14 (N_14,In_182,In_30);
and U15 (N_15,In_374,In_112);
nand U16 (N_16,In_111,In_222);
or U17 (N_17,In_337,In_45);
nand U18 (N_18,In_400,In_173);
nor U19 (N_19,In_406,In_200);
or U20 (N_20,In_344,In_229);
nor U21 (N_21,In_26,In_351);
nor U22 (N_22,In_302,In_253);
nor U23 (N_23,In_453,In_309);
or U24 (N_24,In_65,In_88);
or U25 (N_25,In_292,In_188);
or U26 (N_26,In_216,In_262);
or U27 (N_27,In_211,In_440);
nor U28 (N_28,In_25,In_178);
and U29 (N_29,In_297,In_390);
and U30 (N_30,In_245,In_270);
nor U31 (N_31,In_166,In_80);
nor U32 (N_32,In_44,In_312);
and U33 (N_33,In_284,In_471);
nor U34 (N_34,In_118,In_332);
or U35 (N_35,In_359,In_385);
or U36 (N_36,In_386,In_59);
and U37 (N_37,In_268,In_75);
or U38 (N_38,In_14,In_473);
nor U39 (N_39,In_313,In_336);
and U40 (N_40,In_83,In_35);
nand U41 (N_41,In_449,In_477);
or U42 (N_42,In_176,In_50);
nand U43 (N_43,In_73,In_6);
and U44 (N_44,In_261,In_158);
and U45 (N_45,In_405,In_493);
and U46 (N_46,In_242,In_148);
and U47 (N_47,In_227,In_422);
or U48 (N_48,In_445,In_177);
or U49 (N_49,In_362,In_114);
or U50 (N_50,In_295,In_237);
nor U51 (N_51,In_240,In_437);
or U52 (N_52,In_410,In_156);
and U53 (N_53,In_171,In_11);
nand U54 (N_54,In_190,In_481);
and U55 (N_55,In_326,In_259);
nand U56 (N_56,In_257,In_18);
nor U57 (N_57,In_451,In_373);
or U58 (N_58,In_2,In_91);
nand U59 (N_59,In_151,In_498);
nor U60 (N_60,In_276,In_363);
nand U61 (N_61,In_52,In_497);
nand U62 (N_62,In_354,In_483);
or U63 (N_63,In_10,In_224);
and U64 (N_64,In_321,In_263);
xnor U65 (N_65,In_128,In_423);
or U66 (N_66,In_494,In_484);
nand U67 (N_67,In_170,In_67);
nand U68 (N_68,In_51,In_149);
nand U69 (N_69,In_357,In_461);
and U70 (N_70,In_465,In_1);
nor U71 (N_71,In_191,In_104);
or U72 (N_72,In_464,In_492);
and U73 (N_73,In_282,In_443);
or U74 (N_74,In_298,In_233);
or U75 (N_75,In_347,In_430);
nor U76 (N_76,In_327,In_243);
nand U77 (N_77,In_379,In_322);
nor U78 (N_78,In_294,In_343);
nand U79 (N_79,In_248,In_458);
or U80 (N_80,In_399,In_89);
nand U81 (N_81,In_205,In_370);
nand U82 (N_82,In_192,In_418);
and U83 (N_83,In_116,In_274);
and U84 (N_84,In_232,In_95);
nor U85 (N_85,In_266,In_117);
nand U86 (N_86,In_7,In_183);
and U87 (N_87,In_241,In_345);
and U88 (N_88,In_180,In_371);
and U89 (N_89,In_376,In_393);
or U90 (N_90,In_283,In_33);
nand U91 (N_91,In_132,In_16);
and U92 (N_92,In_115,In_291);
or U93 (N_93,In_37,In_275);
or U94 (N_94,In_186,In_5);
or U95 (N_95,In_324,In_444);
nor U96 (N_96,In_375,In_81);
or U97 (N_97,In_395,In_439);
nor U98 (N_98,In_61,In_323);
and U99 (N_99,In_185,In_31);
and U100 (N_100,In_366,In_278);
nand U101 (N_101,In_365,In_467);
or U102 (N_102,In_13,In_92);
or U103 (N_103,In_109,In_234);
nand U104 (N_104,In_250,In_404);
or U105 (N_105,In_213,In_38);
and U106 (N_106,In_384,In_134);
nand U107 (N_107,In_113,In_207);
nand U108 (N_108,In_3,In_198);
nor U109 (N_109,In_15,In_175);
and U110 (N_110,In_133,In_47);
nor U111 (N_111,In_17,In_448);
nor U112 (N_112,In_346,In_455);
and U113 (N_113,In_368,In_361);
and U114 (N_114,In_446,In_165);
nor U115 (N_115,In_119,In_144);
or U116 (N_116,In_29,In_101);
and U117 (N_117,In_267,In_66);
nor U118 (N_118,In_478,In_77);
xor U119 (N_119,In_247,In_157);
nand U120 (N_120,In_228,In_482);
nand U121 (N_121,In_391,In_181);
nand U122 (N_122,In_208,In_490);
nand U123 (N_123,In_93,In_367);
or U124 (N_124,In_315,In_163);
xor U125 (N_125,In_339,In_90);
nor U126 (N_126,In_426,In_433);
nor U127 (N_127,In_454,In_381);
and U128 (N_128,In_335,In_293);
nor U129 (N_129,In_476,In_486);
or U130 (N_130,In_273,In_318);
and U131 (N_131,In_417,In_197);
nand U132 (N_132,In_21,In_121);
and U133 (N_133,In_56,In_20);
nor U134 (N_134,In_287,In_43);
and U135 (N_135,In_383,In_314);
nor U136 (N_136,In_308,In_491);
nand U137 (N_137,In_470,In_152);
nor U138 (N_138,In_131,In_325);
or U139 (N_139,In_489,In_41);
or U140 (N_140,In_27,In_69);
or U141 (N_141,In_311,In_398);
or U142 (N_142,In_435,In_272);
nand U143 (N_143,In_169,In_457);
and U144 (N_144,In_179,In_206);
or U145 (N_145,In_277,In_204);
nor U146 (N_146,In_244,In_103);
nor U147 (N_147,In_280,In_64);
and U148 (N_148,In_258,In_388);
nor U149 (N_149,In_136,In_416);
nor U150 (N_150,In_427,In_209);
nand U151 (N_151,In_286,In_341);
nor U152 (N_152,In_352,In_251);
or U153 (N_153,In_333,In_71);
xor U154 (N_154,In_23,In_184);
or U155 (N_155,In_24,In_218);
and U156 (N_156,In_424,In_468);
and U157 (N_157,In_496,In_231);
nor U158 (N_158,In_130,In_86);
and U159 (N_159,In_348,In_394);
nand U160 (N_160,In_60,In_409);
nand U161 (N_161,In_137,In_28);
nor U162 (N_162,In_48,In_76);
or U163 (N_163,In_110,In_32);
xnor U164 (N_164,In_53,In_431);
nor U165 (N_165,In_279,In_403);
or U166 (N_166,In_189,In_40);
nor U167 (N_167,In_220,In_269);
xnor U168 (N_168,In_290,In_145);
nor U169 (N_169,In_12,In_155);
or U170 (N_170,In_305,In_296);
or U171 (N_171,In_256,In_138);
or U172 (N_172,In_306,In_329);
or U173 (N_173,In_221,In_238);
xnor U174 (N_174,In_19,In_55);
or U175 (N_175,In_78,In_42);
and U176 (N_176,In_97,In_320);
nor U177 (N_177,In_58,In_252);
and U178 (N_178,In_174,In_217);
nor U179 (N_179,In_122,In_107);
and U180 (N_180,In_450,In_301);
and U181 (N_181,In_411,In_36);
or U182 (N_182,In_389,In_360);
nor U183 (N_183,In_469,In_330);
and U184 (N_184,In_230,In_419);
nand U185 (N_185,In_235,In_63);
nor U186 (N_186,In_340,In_350);
or U187 (N_187,In_68,In_254);
and U188 (N_188,In_94,In_162);
nand U189 (N_189,In_84,In_414);
and U190 (N_190,In_147,In_225);
and U191 (N_191,In_167,In_462);
nand U192 (N_192,In_39,In_187);
nor U193 (N_193,In_463,In_105);
and U194 (N_194,In_485,In_214);
and U195 (N_195,In_358,In_299);
nor U196 (N_196,In_396,In_203);
nand U197 (N_197,In_98,In_108);
nor U198 (N_198,In_34,In_271);
nand U199 (N_199,In_168,In_401);
and U200 (N_200,In_219,In_425);
and U201 (N_201,In_265,In_126);
and U202 (N_202,In_317,In_364);
nand U203 (N_203,In_100,In_472);
nand U204 (N_204,In_499,In_387);
or U205 (N_205,In_434,In_407);
xnor U206 (N_206,In_377,In_139);
nand U207 (N_207,In_85,In_310);
nor U208 (N_208,In_164,In_428);
nand U209 (N_209,In_452,In_196);
and U210 (N_210,In_438,In_70);
or U211 (N_211,In_54,In_307);
and U212 (N_212,In_79,In_480);
or U213 (N_213,In_421,In_459);
and U214 (N_214,In_153,In_460);
or U215 (N_215,In_304,In_127);
or U216 (N_216,In_338,In_334);
nor U217 (N_217,In_331,In_125);
xor U218 (N_218,In_49,In_4);
or U219 (N_219,In_260,In_475);
and U220 (N_220,In_8,In_300);
nor U221 (N_221,In_397,In_226);
nand U222 (N_222,In_356,In_246);
and U223 (N_223,In_74,In_141);
or U224 (N_224,In_124,In_413);
and U225 (N_225,In_479,In_369);
nand U226 (N_226,In_82,In_87);
and U227 (N_227,In_288,In_382);
nand U228 (N_228,In_212,In_316);
xor U229 (N_229,In_159,In_488);
nand U230 (N_230,In_429,In_285);
or U231 (N_231,In_328,In_442);
or U232 (N_232,In_342,In_447);
nor U233 (N_233,In_102,In_106);
or U234 (N_234,In_161,In_160);
nor U235 (N_235,In_199,In_392);
nand U236 (N_236,In_72,In_456);
nand U237 (N_237,In_415,In_353);
and U238 (N_238,In_146,In_9);
or U239 (N_239,In_239,In_123);
nor U240 (N_240,In_487,In_236);
nand U241 (N_241,In_210,In_408);
nor U242 (N_242,In_129,In_99);
nor U243 (N_243,In_143,In_223);
nand U244 (N_244,In_355,In_495);
and U245 (N_245,In_378,In_135);
or U246 (N_246,In_193,In_96);
and U247 (N_247,In_154,In_46);
xnor U248 (N_248,In_466,In_319);
nor U249 (N_249,In_412,In_249);
or U250 (N_250,In_131,In_463);
nor U251 (N_251,In_191,In_121);
nor U252 (N_252,In_467,In_413);
nor U253 (N_253,In_23,In_55);
and U254 (N_254,In_200,In_497);
nand U255 (N_255,In_98,In_455);
nor U256 (N_256,In_185,In_112);
nand U257 (N_257,In_268,In_175);
nand U258 (N_258,In_246,In_240);
nor U259 (N_259,In_267,In_327);
nor U260 (N_260,In_409,In_154);
nor U261 (N_261,In_129,In_161);
and U262 (N_262,In_80,In_467);
and U263 (N_263,In_47,In_139);
or U264 (N_264,In_181,In_319);
and U265 (N_265,In_349,In_460);
or U266 (N_266,In_457,In_449);
nand U267 (N_267,In_425,In_21);
nor U268 (N_268,In_496,In_209);
nand U269 (N_269,In_491,In_30);
nor U270 (N_270,In_266,In_326);
nand U271 (N_271,In_141,In_208);
and U272 (N_272,In_417,In_331);
or U273 (N_273,In_101,In_417);
nand U274 (N_274,In_130,In_467);
nor U275 (N_275,In_6,In_317);
or U276 (N_276,In_323,In_49);
and U277 (N_277,In_12,In_460);
or U278 (N_278,In_87,In_247);
nand U279 (N_279,In_157,In_376);
xnor U280 (N_280,In_132,In_294);
or U281 (N_281,In_454,In_189);
xor U282 (N_282,In_340,In_442);
xor U283 (N_283,In_469,In_388);
or U284 (N_284,In_317,In_264);
nor U285 (N_285,In_418,In_19);
xnor U286 (N_286,In_400,In_392);
and U287 (N_287,In_313,In_159);
and U288 (N_288,In_492,In_121);
nand U289 (N_289,In_67,In_2);
nor U290 (N_290,In_127,In_208);
or U291 (N_291,In_289,In_302);
nand U292 (N_292,In_103,In_92);
or U293 (N_293,In_372,In_68);
nor U294 (N_294,In_398,In_374);
and U295 (N_295,In_110,In_275);
nor U296 (N_296,In_124,In_315);
nand U297 (N_297,In_57,In_59);
nor U298 (N_298,In_3,In_228);
nor U299 (N_299,In_200,In_172);
nor U300 (N_300,In_355,In_441);
and U301 (N_301,In_360,In_247);
nand U302 (N_302,In_154,In_471);
and U303 (N_303,In_146,In_276);
or U304 (N_304,In_497,In_459);
or U305 (N_305,In_498,In_384);
nand U306 (N_306,In_42,In_271);
nand U307 (N_307,In_379,In_406);
nor U308 (N_308,In_226,In_144);
nand U309 (N_309,In_217,In_489);
xnor U310 (N_310,In_406,In_245);
or U311 (N_311,In_393,In_131);
or U312 (N_312,In_144,In_343);
and U313 (N_313,In_102,In_379);
or U314 (N_314,In_299,In_396);
nand U315 (N_315,In_86,In_136);
or U316 (N_316,In_235,In_142);
and U317 (N_317,In_337,In_63);
nor U318 (N_318,In_494,In_103);
nand U319 (N_319,In_111,In_380);
nand U320 (N_320,In_102,In_197);
nand U321 (N_321,In_234,In_104);
nand U322 (N_322,In_449,In_55);
nor U323 (N_323,In_283,In_197);
and U324 (N_324,In_83,In_433);
nor U325 (N_325,In_438,In_73);
nand U326 (N_326,In_205,In_355);
or U327 (N_327,In_84,In_296);
or U328 (N_328,In_134,In_421);
or U329 (N_329,In_385,In_266);
nor U330 (N_330,In_425,In_265);
and U331 (N_331,In_62,In_465);
nor U332 (N_332,In_162,In_229);
nand U333 (N_333,In_376,In_284);
or U334 (N_334,In_48,In_127);
nor U335 (N_335,In_198,In_362);
nand U336 (N_336,In_33,In_165);
and U337 (N_337,In_153,In_357);
or U338 (N_338,In_378,In_437);
or U339 (N_339,In_465,In_389);
nor U340 (N_340,In_470,In_408);
or U341 (N_341,In_226,In_145);
nand U342 (N_342,In_123,In_492);
and U343 (N_343,In_454,In_247);
nor U344 (N_344,In_11,In_294);
nor U345 (N_345,In_7,In_397);
nand U346 (N_346,In_370,In_441);
nand U347 (N_347,In_93,In_173);
and U348 (N_348,In_307,In_126);
or U349 (N_349,In_206,In_223);
nor U350 (N_350,In_437,In_477);
or U351 (N_351,In_337,In_157);
or U352 (N_352,In_408,In_136);
nor U353 (N_353,In_324,In_389);
or U354 (N_354,In_163,In_277);
or U355 (N_355,In_264,In_41);
nand U356 (N_356,In_238,In_333);
and U357 (N_357,In_30,In_492);
nand U358 (N_358,In_166,In_152);
xnor U359 (N_359,In_410,In_21);
nand U360 (N_360,In_197,In_302);
nor U361 (N_361,In_15,In_198);
nor U362 (N_362,In_219,In_315);
or U363 (N_363,In_355,In_7);
nand U364 (N_364,In_284,In_145);
nor U365 (N_365,In_43,In_390);
and U366 (N_366,In_452,In_308);
nand U367 (N_367,In_129,In_97);
nand U368 (N_368,In_103,In_108);
or U369 (N_369,In_159,In_310);
or U370 (N_370,In_374,In_461);
nor U371 (N_371,In_283,In_127);
nand U372 (N_372,In_32,In_281);
and U373 (N_373,In_14,In_249);
nor U374 (N_374,In_199,In_13);
and U375 (N_375,In_484,In_374);
nand U376 (N_376,In_348,In_156);
nor U377 (N_377,In_318,In_204);
and U378 (N_378,In_243,In_497);
or U379 (N_379,In_342,In_268);
or U380 (N_380,In_307,In_11);
nand U381 (N_381,In_60,In_270);
nor U382 (N_382,In_254,In_95);
or U383 (N_383,In_194,In_91);
nand U384 (N_384,In_121,In_426);
or U385 (N_385,In_466,In_403);
nand U386 (N_386,In_74,In_68);
nor U387 (N_387,In_139,In_9);
xor U388 (N_388,In_209,In_308);
nand U389 (N_389,In_314,In_469);
and U390 (N_390,In_469,In_369);
or U391 (N_391,In_353,In_352);
or U392 (N_392,In_350,In_459);
and U393 (N_393,In_40,In_116);
nand U394 (N_394,In_119,In_260);
nand U395 (N_395,In_187,In_235);
nand U396 (N_396,In_328,In_353);
nand U397 (N_397,In_258,In_405);
and U398 (N_398,In_431,In_407);
and U399 (N_399,In_365,In_343);
and U400 (N_400,In_85,In_484);
nand U401 (N_401,In_459,In_461);
and U402 (N_402,In_235,In_426);
xor U403 (N_403,In_161,In_132);
nor U404 (N_404,In_92,In_184);
nand U405 (N_405,In_239,In_82);
nor U406 (N_406,In_430,In_380);
or U407 (N_407,In_180,In_141);
nor U408 (N_408,In_352,In_182);
and U409 (N_409,In_396,In_231);
and U410 (N_410,In_244,In_310);
nor U411 (N_411,In_399,In_107);
and U412 (N_412,In_296,In_444);
nand U413 (N_413,In_282,In_46);
or U414 (N_414,In_278,In_148);
and U415 (N_415,In_142,In_346);
or U416 (N_416,In_155,In_366);
nand U417 (N_417,In_341,In_399);
and U418 (N_418,In_25,In_235);
nor U419 (N_419,In_280,In_39);
nor U420 (N_420,In_81,In_64);
nor U421 (N_421,In_358,In_131);
xor U422 (N_422,In_481,In_97);
nor U423 (N_423,In_156,In_483);
and U424 (N_424,In_420,In_274);
nand U425 (N_425,In_194,In_61);
or U426 (N_426,In_0,In_191);
nand U427 (N_427,In_459,In_167);
or U428 (N_428,In_376,In_228);
or U429 (N_429,In_212,In_33);
nand U430 (N_430,In_193,In_62);
nand U431 (N_431,In_348,In_283);
and U432 (N_432,In_72,In_348);
or U433 (N_433,In_380,In_58);
nand U434 (N_434,In_53,In_486);
and U435 (N_435,In_450,In_477);
nor U436 (N_436,In_357,In_224);
or U437 (N_437,In_14,In_204);
nor U438 (N_438,In_99,In_33);
nand U439 (N_439,In_23,In_410);
nand U440 (N_440,In_345,In_76);
nor U441 (N_441,In_388,In_392);
and U442 (N_442,In_34,In_0);
and U443 (N_443,In_280,In_485);
and U444 (N_444,In_382,In_319);
or U445 (N_445,In_324,In_434);
or U446 (N_446,In_439,In_254);
xor U447 (N_447,In_499,In_95);
nand U448 (N_448,In_286,In_208);
or U449 (N_449,In_391,In_113);
nor U450 (N_450,In_206,In_225);
nand U451 (N_451,In_303,In_296);
nor U452 (N_452,In_370,In_262);
nor U453 (N_453,In_278,In_29);
nand U454 (N_454,In_212,In_420);
nand U455 (N_455,In_459,In_72);
xnor U456 (N_456,In_383,In_77);
or U457 (N_457,In_187,In_317);
nor U458 (N_458,In_206,In_156);
xnor U459 (N_459,In_91,In_359);
nor U460 (N_460,In_393,In_98);
nand U461 (N_461,In_33,In_8);
nand U462 (N_462,In_422,In_117);
nor U463 (N_463,In_106,In_346);
or U464 (N_464,In_439,In_215);
and U465 (N_465,In_255,In_23);
or U466 (N_466,In_389,In_352);
nand U467 (N_467,In_231,In_154);
or U468 (N_468,In_269,In_169);
and U469 (N_469,In_270,In_255);
and U470 (N_470,In_81,In_213);
and U471 (N_471,In_157,In_330);
nor U472 (N_472,In_497,In_452);
nor U473 (N_473,In_324,In_479);
or U474 (N_474,In_122,In_45);
nor U475 (N_475,In_272,In_355);
and U476 (N_476,In_441,In_257);
nor U477 (N_477,In_256,In_283);
nand U478 (N_478,In_61,In_279);
or U479 (N_479,In_353,In_43);
nand U480 (N_480,In_47,In_430);
nand U481 (N_481,In_338,In_487);
and U482 (N_482,In_190,In_343);
nor U483 (N_483,In_431,In_397);
and U484 (N_484,In_118,In_130);
nand U485 (N_485,In_394,In_134);
or U486 (N_486,In_3,In_10);
and U487 (N_487,In_225,In_482);
and U488 (N_488,In_318,In_322);
nand U489 (N_489,In_51,In_230);
nand U490 (N_490,In_51,In_87);
and U491 (N_491,In_347,In_329);
and U492 (N_492,In_11,In_215);
nand U493 (N_493,In_390,In_303);
or U494 (N_494,In_472,In_74);
nand U495 (N_495,In_72,In_416);
nand U496 (N_496,In_171,In_32);
or U497 (N_497,In_350,In_14);
nor U498 (N_498,In_404,In_286);
or U499 (N_499,In_115,In_283);
and U500 (N_500,In_45,In_368);
nor U501 (N_501,In_12,In_33);
xor U502 (N_502,In_338,In_335);
nand U503 (N_503,In_166,In_457);
or U504 (N_504,In_460,In_475);
nor U505 (N_505,In_41,In_278);
and U506 (N_506,In_347,In_325);
or U507 (N_507,In_329,In_163);
nand U508 (N_508,In_263,In_51);
and U509 (N_509,In_255,In_60);
or U510 (N_510,In_359,In_409);
nor U511 (N_511,In_136,In_125);
or U512 (N_512,In_70,In_2);
or U513 (N_513,In_57,In_251);
nor U514 (N_514,In_394,In_333);
or U515 (N_515,In_56,In_350);
or U516 (N_516,In_427,In_318);
and U517 (N_517,In_167,In_384);
nor U518 (N_518,In_213,In_462);
and U519 (N_519,In_41,In_89);
nand U520 (N_520,In_314,In_233);
xor U521 (N_521,In_55,In_49);
or U522 (N_522,In_73,In_427);
nor U523 (N_523,In_115,In_233);
nor U524 (N_524,In_7,In_256);
and U525 (N_525,In_11,In_275);
nor U526 (N_526,In_361,In_466);
and U527 (N_527,In_261,In_126);
nand U528 (N_528,In_188,In_303);
or U529 (N_529,In_83,In_72);
and U530 (N_530,In_165,In_322);
nor U531 (N_531,In_169,In_345);
nor U532 (N_532,In_13,In_252);
or U533 (N_533,In_79,In_337);
and U534 (N_534,In_285,In_396);
nand U535 (N_535,In_46,In_288);
nand U536 (N_536,In_22,In_450);
nor U537 (N_537,In_275,In_124);
nand U538 (N_538,In_443,In_384);
and U539 (N_539,In_313,In_226);
or U540 (N_540,In_220,In_475);
and U541 (N_541,In_165,In_107);
or U542 (N_542,In_114,In_452);
nor U543 (N_543,In_232,In_332);
and U544 (N_544,In_244,In_433);
or U545 (N_545,In_18,In_275);
nand U546 (N_546,In_479,In_417);
nand U547 (N_547,In_414,In_383);
or U548 (N_548,In_495,In_97);
nor U549 (N_549,In_231,In_290);
or U550 (N_550,In_384,In_102);
nor U551 (N_551,In_149,In_334);
or U552 (N_552,In_478,In_405);
nand U553 (N_553,In_474,In_437);
nor U554 (N_554,In_382,In_436);
or U555 (N_555,In_221,In_38);
nor U556 (N_556,In_101,In_336);
or U557 (N_557,In_89,In_390);
nand U558 (N_558,In_487,In_365);
nor U559 (N_559,In_104,In_59);
nor U560 (N_560,In_383,In_20);
nand U561 (N_561,In_331,In_455);
and U562 (N_562,In_235,In_18);
nand U563 (N_563,In_496,In_69);
nand U564 (N_564,In_424,In_130);
nand U565 (N_565,In_23,In_316);
nor U566 (N_566,In_89,In_285);
xnor U567 (N_567,In_1,In_387);
nand U568 (N_568,In_291,In_445);
nand U569 (N_569,In_444,In_307);
nor U570 (N_570,In_358,In_114);
or U571 (N_571,In_5,In_405);
nand U572 (N_572,In_191,In_468);
nor U573 (N_573,In_453,In_406);
nand U574 (N_574,In_129,In_177);
xnor U575 (N_575,In_121,In_462);
nor U576 (N_576,In_138,In_335);
or U577 (N_577,In_45,In_364);
and U578 (N_578,In_303,In_25);
nor U579 (N_579,In_97,In_85);
or U580 (N_580,In_316,In_240);
or U581 (N_581,In_379,In_109);
and U582 (N_582,In_308,In_67);
and U583 (N_583,In_427,In_31);
or U584 (N_584,In_343,In_137);
or U585 (N_585,In_391,In_25);
nor U586 (N_586,In_267,In_134);
nor U587 (N_587,In_45,In_279);
xnor U588 (N_588,In_115,In_386);
nand U589 (N_589,In_482,In_190);
and U590 (N_590,In_55,In_180);
nor U591 (N_591,In_361,In_2);
nand U592 (N_592,In_91,In_78);
or U593 (N_593,In_494,In_386);
nand U594 (N_594,In_298,In_147);
nor U595 (N_595,In_334,In_248);
nor U596 (N_596,In_366,In_177);
or U597 (N_597,In_462,In_413);
nand U598 (N_598,In_260,In_305);
nand U599 (N_599,In_370,In_485);
nor U600 (N_600,In_101,In_273);
or U601 (N_601,In_238,In_194);
or U602 (N_602,In_294,In_429);
and U603 (N_603,In_277,In_223);
or U604 (N_604,In_487,In_479);
or U605 (N_605,In_414,In_176);
or U606 (N_606,In_300,In_113);
nor U607 (N_607,In_426,In_59);
and U608 (N_608,In_188,In_1);
and U609 (N_609,In_26,In_489);
or U610 (N_610,In_385,In_225);
and U611 (N_611,In_477,In_291);
nor U612 (N_612,In_377,In_136);
nor U613 (N_613,In_56,In_364);
or U614 (N_614,In_230,In_31);
or U615 (N_615,In_466,In_472);
nor U616 (N_616,In_12,In_107);
nor U617 (N_617,In_235,In_76);
nand U618 (N_618,In_237,In_274);
nand U619 (N_619,In_174,In_98);
nand U620 (N_620,In_349,In_428);
or U621 (N_621,In_441,In_139);
or U622 (N_622,In_58,In_27);
or U623 (N_623,In_110,In_366);
and U624 (N_624,In_209,In_411);
nand U625 (N_625,In_139,In_172);
and U626 (N_626,In_77,In_323);
and U627 (N_627,In_252,In_16);
and U628 (N_628,In_96,In_333);
or U629 (N_629,In_92,In_234);
nor U630 (N_630,In_322,In_341);
and U631 (N_631,In_150,In_73);
nor U632 (N_632,In_238,In_215);
or U633 (N_633,In_208,In_45);
or U634 (N_634,In_374,In_142);
xnor U635 (N_635,In_415,In_381);
xor U636 (N_636,In_137,In_189);
nor U637 (N_637,In_294,In_138);
nor U638 (N_638,In_59,In_308);
or U639 (N_639,In_61,In_373);
nand U640 (N_640,In_398,In_460);
or U641 (N_641,In_289,In_293);
and U642 (N_642,In_288,In_138);
xor U643 (N_643,In_163,In_54);
and U644 (N_644,In_305,In_306);
and U645 (N_645,In_373,In_8);
nand U646 (N_646,In_27,In_420);
nor U647 (N_647,In_489,In_478);
or U648 (N_648,In_29,In_229);
or U649 (N_649,In_336,In_178);
or U650 (N_650,In_186,In_327);
and U651 (N_651,In_357,In_356);
nand U652 (N_652,In_485,In_450);
or U653 (N_653,In_87,In_88);
nand U654 (N_654,In_2,In_300);
or U655 (N_655,In_167,In_140);
nor U656 (N_656,In_80,In_314);
and U657 (N_657,In_394,In_425);
nand U658 (N_658,In_365,In_207);
nor U659 (N_659,In_399,In_309);
nand U660 (N_660,In_316,In_58);
or U661 (N_661,In_153,In_318);
or U662 (N_662,In_436,In_343);
nor U663 (N_663,In_162,In_189);
nand U664 (N_664,In_257,In_161);
nand U665 (N_665,In_229,In_95);
nor U666 (N_666,In_212,In_77);
and U667 (N_667,In_109,In_270);
nor U668 (N_668,In_169,In_476);
or U669 (N_669,In_276,In_481);
nand U670 (N_670,In_161,In_442);
nor U671 (N_671,In_301,In_148);
nand U672 (N_672,In_86,In_173);
or U673 (N_673,In_243,In_400);
nand U674 (N_674,In_229,In_142);
nand U675 (N_675,In_107,In_484);
nand U676 (N_676,In_31,In_108);
nand U677 (N_677,In_43,In_436);
nor U678 (N_678,In_73,In_68);
nor U679 (N_679,In_15,In_278);
or U680 (N_680,In_456,In_297);
and U681 (N_681,In_242,In_201);
and U682 (N_682,In_73,In_142);
and U683 (N_683,In_75,In_81);
nor U684 (N_684,In_88,In_236);
or U685 (N_685,In_366,In_97);
nand U686 (N_686,In_183,In_476);
xor U687 (N_687,In_258,In_185);
nand U688 (N_688,In_341,In_390);
or U689 (N_689,In_217,In_198);
nand U690 (N_690,In_164,In_479);
nand U691 (N_691,In_466,In_108);
nand U692 (N_692,In_384,In_375);
nor U693 (N_693,In_238,In_355);
nand U694 (N_694,In_144,In_23);
or U695 (N_695,In_444,In_93);
or U696 (N_696,In_264,In_169);
or U697 (N_697,In_493,In_67);
and U698 (N_698,In_142,In_67);
nand U699 (N_699,In_290,In_474);
nand U700 (N_700,In_230,In_3);
and U701 (N_701,In_22,In_460);
nor U702 (N_702,In_193,In_268);
nand U703 (N_703,In_172,In_487);
and U704 (N_704,In_196,In_111);
and U705 (N_705,In_350,In_364);
nor U706 (N_706,In_346,In_497);
or U707 (N_707,In_102,In_251);
or U708 (N_708,In_260,In_281);
nor U709 (N_709,In_374,In_286);
nor U710 (N_710,In_24,In_94);
xor U711 (N_711,In_211,In_97);
or U712 (N_712,In_355,In_386);
and U713 (N_713,In_238,In_442);
and U714 (N_714,In_388,In_279);
and U715 (N_715,In_312,In_164);
and U716 (N_716,In_79,In_242);
nand U717 (N_717,In_144,In_460);
or U718 (N_718,In_212,In_337);
xnor U719 (N_719,In_35,In_300);
nand U720 (N_720,In_268,In_79);
nor U721 (N_721,In_120,In_232);
nor U722 (N_722,In_86,In_281);
or U723 (N_723,In_339,In_210);
nand U724 (N_724,In_301,In_481);
and U725 (N_725,In_130,In_98);
and U726 (N_726,In_340,In_406);
nor U727 (N_727,In_334,In_374);
and U728 (N_728,In_207,In_171);
and U729 (N_729,In_359,In_300);
nor U730 (N_730,In_260,In_299);
or U731 (N_731,In_342,In_307);
nor U732 (N_732,In_246,In_427);
or U733 (N_733,In_118,In_288);
xnor U734 (N_734,In_213,In_46);
or U735 (N_735,In_69,In_448);
nand U736 (N_736,In_90,In_134);
nand U737 (N_737,In_19,In_24);
nor U738 (N_738,In_89,In_370);
and U739 (N_739,In_92,In_122);
nor U740 (N_740,In_272,In_29);
and U741 (N_741,In_38,In_131);
and U742 (N_742,In_15,In_261);
nor U743 (N_743,In_193,In_405);
or U744 (N_744,In_178,In_24);
and U745 (N_745,In_277,In_259);
nor U746 (N_746,In_80,In_187);
and U747 (N_747,In_407,In_84);
or U748 (N_748,In_0,In_132);
nor U749 (N_749,In_127,In_403);
nand U750 (N_750,N_626,N_342);
and U751 (N_751,N_41,N_484);
nor U752 (N_752,N_599,N_482);
and U753 (N_753,N_493,N_258);
nand U754 (N_754,N_522,N_634);
nand U755 (N_755,N_26,N_704);
nand U756 (N_756,N_180,N_43);
nor U757 (N_757,N_461,N_149);
nor U758 (N_758,N_458,N_111);
nor U759 (N_759,N_492,N_297);
and U760 (N_760,N_479,N_202);
nor U761 (N_761,N_621,N_344);
nor U762 (N_762,N_619,N_370);
or U763 (N_763,N_734,N_347);
and U764 (N_764,N_93,N_594);
nand U765 (N_765,N_345,N_361);
and U766 (N_766,N_495,N_302);
nor U767 (N_767,N_282,N_736);
and U768 (N_768,N_604,N_505);
and U769 (N_769,N_469,N_655);
and U770 (N_770,N_336,N_680);
and U771 (N_771,N_511,N_671);
nor U772 (N_772,N_133,N_348);
xor U773 (N_773,N_176,N_86);
and U774 (N_774,N_389,N_657);
or U775 (N_775,N_579,N_618);
nand U776 (N_776,N_448,N_230);
or U777 (N_777,N_527,N_506);
and U778 (N_778,N_724,N_94);
and U779 (N_779,N_502,N_318);
and U780 (N_780,N_474,N_185);
nor U781 (N_781,N_18,N_317);
or U782 (N_782,N_309,N_686);
and U783 (N_783,N_32,N_584);
or U784 (N_784,N_20,N_320);
nor U785 (N_785,N_512,N_379);
nor U786 (N_786,N_677,N_683);
and U787 (N_787,N_196,N_614);
nand U788 (N_788,N_744,N_443);
nor U789 (N_789,N_366,N_84);
and U790 (N_790,N_166,N_374);
nand U791 (N_791,N_650,N_627);
nand U792 (N_792,N_652,N_706);
nor U793 (N_793,N_423,N_210);
nand U794 (N_794,N_37,N_333);
nor U795 (N_795,N_556,N_30);
or U796 (N_796,N_748,N_158);
and U797 (N_797,N_433,N_47);
nor U798 (N_798,N_412,N_77);
nor U799 (N_799,N_477,N_384);
or U800 (N_800,N_659,N_606);
nor U801 (N_801,N_431,N_733);
or U802 (N_802,N_540,N_179);
nand U803 (N_803,N_171,N_549);
and U804 (N_804,N_514,N_731);
or U805 (N_805,N_146,N_281);
nor U806 (N_806,N_656,N_268);
nand U807 (N_807,N_689,N_603);
nor U808 (N_808,N_69,N_102);
nor U809 (N_809,N_719,N_82);
and U810 (N_810,N_112,N_548);
and U811 (N_811,N_58,N_245);
or U812 (N_812,N_714,N_265);
and U813 (N_813,N_78,N_647);
or U814 (N_814,N_295,N_516);
nor U815 (N_815,N_216,N_88);
nor U816 (N_816,N_29,N_145);
and U817 (N_817,N_645,N_118);
and U818 (N_818,N_131,N_580);
nand U819 (N_819,N_228,N_184);
nand U820 (N_820,N_161,N_83);
or U821 (N_821,N_221,N_75);
or U822 (N_822,N_546,N_193);
nand U823 (N_823,N_498,N_306);
nor U824 (N_824,N_411,N_515);
nand U825 (N_825,N_497,N_590);
and U826 (N_826,N_369,N_142);
and U827 (N_827,N_526,N_682);
nor U828 (N_828,N_392,N_715);
and U829 (N_829,N_509,N_653);
or U830 (N_830,N_568,N_508);
xor U831 (N_831,N_726,N_292);
xnor U832 (N_832,N_528,N_17);
nor U833 (N_833,N_613,N_698);
and U834 (N_834,N_223,N_643);
xnor U835 (N_835,N_324,N_312);
nor U836 (N_836,N_39,N_141);
nor U837 (N_837,N_359,N_288);
nor U838 (N_838,N_425,N_353);
or U839 (N_839,N_541,N_672);
and U840 (N_840,N_503,N_346);
xnor U841 (N_841,N_91,N_33);
or U842 (N_842,N_194,N_181);
or U843 (N_843,N_625,N_103);
or U844 (N_844,N_520,N_351);
nor U845 (N_845,N_665,N_729);
nand U846 (N_846,N_128,N_319);
nor U847 (N_847,N_406,N_337);
xnor U848 (N_848,N_271,N_561);
or U849 (N_849,N_19,N_373);
or U850 (N_850,N_670,N_447);
nand U851 (N_851,N_340,N_457);
nor U852 (N_852,N_175,N_487);
or U853 (N_853,N_450,N_620);
and U854 (N_854,N_405,N_617);
nor U855 (N_855,N_410,N_674);
or U856 (N_856,N_67,N_50);
or U857 (N_857,N_628,N_428);
nor U858 (N_858,N_415,N_55);
or U859 (N_859,N_162,N_227);
nor U860 (N_860,N_262,N_385);
nor U861 (N_861,N_261,N_441);
xnor U862 (N_862,N_28,N_130);
nor U863 (N_863,N_636,N_700);
xnor U864 (N_864,N_126,N_290);
nand U865 (N_865,N_48,N_298);
nor U866 (N_866,N_589,N_436);
xor U867 (N_867,N_658,N_259);
or U868 (N_868,N_247,N_608);
nand U869 (N_869,N_710,N_3);
nor U870 (N_870,N_574,N_220);
nor U871 (N_871,N_140,N_397);
nor U872 (N_872,N_135,N_115);
nand U873 (N_873,N_570,N_387);
or U874 (N_874,N_473,N_692);
nor U875 (N_875,N_462,N_11);
nor U876 (N_876,N_684,N_496);
and U877 (N_877,N_558,N_195);
and U878 (N_878,N_399,N_721);
xnor U879 (N_879,N_615,N_712);
nor U880 (N_880,N_697,N_99);
and U881 (N_881,N_197,N_738);
and U882 (N_882,N_534,N_163);
or U883 (N_883,N_651,N_96);
nand U884 (N_884,N_113,N_286);
nand U885 (N_885,N_501,N_407);
and U886 (N_886,N_246,N_287);
and U887 (N_887,N_311,N_676);
or U888 (N_888,N_155,N_349);
and U889 (N_889,N_539,N_660);
or U890 (N_890,N_390,N_357);
and U891 (N_891,N_421,N_630);
or U892 (N_892,N_74,N_600);
or U893 (N_893,N_231,N_269);
or U894 (N_894,N_424,N_681);
nand U895 (N_895,N_310,N_23);
nand U896 (N_896,N_530,N_510);
nand U897 (N_897,N_521,N_642);
nand U898 (N_898,N_483,N_709);
nand U899 (N_899,N_485,N_241);
nand U900 (N_900,N_254,N_352);
nand U901 (N_901,N_609,N_275);
nand U902 (N_902,N_679,N_637);
or U903 (N_903,N_593,N_631);
or U904 (N_904,N_662,N_730);
nor U905 (N_905,N_741,N_439);
or U906 (N_906,N_13,N_213);
or U907 (N_907,N_468,N_5);
nand U908 (N_908,N_124,N_622);
nor U909 (N_909,N_576,N_742);
nor U910 (N_910,N_654,N_61);
nand U911 (N_911,N_335,N_240);
nand U912 (N_912,N_648,N_270);
nor U913 (N_913,N_266,N_343);
and U914 (N_914,N_418,N_455);
nor U915 (N_915,N_147,N_587);
nor U916 (N_916,N_56,N_276);
and U917 (N_917,N_170,N_430);
or U918 (N_918,N_393,N_263);
nor U919 (N_919,N_695,N_699);
and U920 (N_920,N_253,N_542);
or U921 (N_921,N_372,N_581);
nor U922 (N_922,N_408,N_460);
nand U923 (N_923,N_136,N_475);
nand U924 (N_924,N_192,N_257);
nand U925 (N_925,N_173,N_577);
and U926 (N_926,N_107,N_693);
nand U927 (N_927,N_138,N_517);
nor U928 (N_928,N_732,N_422);
nand U929 (N_929,N_172,N_416);
xor U930 (N_930,N_440,N_480);
or U931 (N_931,N_190,N_116);
and U932 (N_932,N_85,N_76);
nand U933 (N_933,N_169,N_144);
or U934 (N_934,N_35,N_446);
nor U935 (N_935,N_117,N_187);
nand U936 (N_936,N_545,N_365);
nand U937 (N_937,N_233,N_16);
nor U938 (N_938,N_225,N_217);
nand U939 (N_939,N_567,N_203);
nand U940 (N_940,N_36,N_394);
nand U941 (N_941,N_191,N_442);
and U942 (N_942,N_537,N_623);
or U943 (N_943,N_206,N_396);
or U944 (N_944,N_4,N_350);
nor U945 (N_945,N_745,N_426);
or U946 (N_946,N_316,N_451);
or U947 (N_947,N_7,N_1);
nor U948 (N_948,N_563,N_92);
xor U949 (N_949,N_504,N_691);
nand U950 (N_950,N_331,N_168);
nand U951 (N_951,N_188,N_702);
nand U952 (N_952,N_685,N_236);
or U953 (N_953,N_728,N_582);
and U954 (N_954,N_229,N_696);
and U955 (N_955,N_129,N_400);
nand U956 (N_956,N_256,N_174);
nor U957 (N_957,N_214,N_607);
nand U958 (N_958,N_204,N_720);
or U959 (N_959,N_10,N_363);
nor U960 (N_960,N_419,N_277);
or U961 (N_961,N_201,N_14);
and U962 (N_962,N_68,N_165);
and U963 (N_963,N_597,N_569);
nor U964 (N_964,N_705,N_101);
or U965 (N_965,N_62,N_494);
nand U966 (N_966,N_326,N_747);
nand U967 (N_967,N_553,N_543);
and U968 (N_968,N_137,N_152);
nand U969 (N_969,N_401,N_575);
or U970 (N_970,N_471,N_452);
or U971 (N_971,N_727,N_454);
or U972 (N_972,N_417,N_322);
and U973 (N_973,N_739,N_740);
or U974 (N_974,N_641,N_100);
nand U975 (N_975,N_602,N_313);
or U976 (N_976,N_383,N_81);
nor U977 (N_977,N_669,N_291);
or U978 (N_978,N_27,N_445);
nor U979 (N_979,N_420,N_464);
nand U980 (N_980,N_612,N_703);
nor U981 (N_981,N_182,N_219);
nand U982 (N_982,N_402,N_71);
nor U983 (N_983,N_325,N_189);
or U984 (N_984,N_122,N_592);
and U985 (N_985,N_127,N_255);
nand U986 (N_986,N_252,N_632);
and U987 (N_987,N_591,N_321);
nand U988 (N_988,N_198,N_746);
and U989 (N_989,N_330,N_588);
nand U990 (N_990,N_666,N_434);
nor U991 (N_991,N_2,N_362);
and U992 (N_992,N_376,N_367);
nor U993 (N_993,N_303,N_513);
nand U994 (N_994,N_24,N_109);
or U995 (N_995,N_722,N_123);
and U996 (N_996,N_108,N_339);
or U997 (N_997,N_358,N_60);
or U998 (N_998,N_64,N_6);
or U999 (N_999,N_437,N_209);
or U1000 (N_1000,N_633,N_488);
or U1001 (N_1001,N_8,N_119);
nand U1002 (N_1002,N_157,N_72);
or U1003 (N_1003,N_667,N_150);
nor U1004 (N_1004,N_465,N_486);
nand U1005 (N_1005,N_79,N_578);
nor U1006 (N_1006,N_525,N_564);
or U1007 (N_1007,N_238,N_65);
nand U1008 (N_1008,N_294,N_151);
or U1009 (N_1009,N_183,N_329);
nand U1010 (N_1010,N_249,N_156);
xor U1011 (N_1011,N_300,N_121);
nand U1012 (N_1012,N_713,N_63);
and U1013 (N_1013,N_315,N_284);
nand U1014 (N_1014,N_0,N_524);
nor U1015 (N_1015,N_596,N_559);
nor U1016 (N_1016,N_46,N_435);
or U1017 (N_1017,N_341,N_360);
and U1018 (N_1018,N_519,N_279);
or U1019 (N_1019,N_749,N_31);
nor U1020 (N_1020,N_375,N_668);
or U1021 (N_1021,N_476,N_42);
or U1022 (N_1022,N_551,N_283);
or U1023 (N_1023,N_293,N_199);
or U1024 (N_1024,N_57,N_610);
or U1025 (N_1025,N_605,N_583);
nor U1026 (N_1026,N_177,N_499);
nand U1027 (N_1027,N_489,N_301);
nor U1028 (N_1028,N_586,N_678);
and U1029 (N_1029,N_160,N_646);
nand U1030 (N_1030,N_97,N_212);
nand U1031 (N_1031,N_364,N_244);
nand U1032 (N_1032,N_38,N_148);
or U1033 (N_1033,N_386,N_114);
nand U1034 (N_1034,N_87,N_132);
and U1035 (N_1035,N_500,N_207);
nor U1036 (N_1036,N_226,N_566);
and U1037 (N_1037,N_332,N_388);
nand U1038 (N_1038,N_304,N_444);
nand U1039 (N_1039,N_242,N_98);
nand U1040 (N_1040,N_110,N_66);
and U1041 (N_1041,N_701,N_380);
and U1042 (N_1042,N_711,N_164);
and U1043 (N_1043,N_40,N_694);
or U1044 (N_1044,N_371,N_529);
nor U1045 (N_1045,N_381,N_562);
nor U1046 (N_1046,N_554,N_305);
nor U1047 (N_1047,N_143,N_273);
nor U1048 (N_1048,N_354,N_449);
or U1049 (N_1049,N_251,N_557);
nor U1050 (N_1050,N_552,N_595);
nand U1051 (N_1051,N_218,N_167);
and U1052 (N_1052,N_232,N_153);
nand U1053 (N_1053,N_154,N_565);
nor U1054 (N_1054,N_544,N_456);
or U1055 (N_1055,N_459,N_687);
and U1056 (N_1056,N_378,N_629);
nor U1057 (N_1057,N_743,N_598);
and U1058 (N_1058,N_572,N_125);
nand U1059 (N_1059,N_708,N_250);
and U1060 (N_1060,N_560,N_395);
nor U1061 (N_1061,N_70,N_21);
nor U1062 (N_1062,N_355,N_15);
nor U1063 (N_1063,N_52,N_9);
and U1064 (N_1064,N_601,N_296);
and U1065 (N_1065,N_267,N_314);
or U1066 (N_1066,N_725,N_299);
xnor U1067 (N_1067,N_690,N_611);
or U1068 (N_1068,N_73,N_334);
or U1069 (N_1069,N_532,N_536);
nand U1070 (N_1070,N_640,N_49);
nor U1071 (N_1071,N_272,N_463);
or U1072 (N_1072,N_644,N_573);
nor U1073 (N_1073,N_34,N_531);
nor U1074 (N_1074,N_432,N_90);
nor U1075 (N_1075,N_518,N_438);
or U1076 (N_1076,N_260,N_413);
nand U1077 (N_1077,N_22,N_639);
or U1078 (N_1078,N_186,N_327);
and U1079 (N_1079,N_661,N_718);
nor U1080 (N_1080,N_472,N_550);
or U1081 (N_1081,N_507,N_427);
and U1082 (N_1082,N_45,N_248);
and U1083 (N_1083,N_538,N_274);
nand U1084 (N_1084,N_224,N_547);
and U1085 (N_1085,N_523,N_707);
or U1086 (N_1086,N_264,N_716);
nor U1087 (N_1087,N_105,N_429);
nand U1088 (N_1088,N_571,N_649);
nor U1089 (N_1089,N_139,N_490);
xnor U1090 (N_1090,N_239,N_737);
or U1091 (N_1091,N_382,N_200);
or U1092 (N_1092,N_453,N_89);
nor U1093 (N_1093,N_134,N_673);
nor U1094 (N_1094,N_688,N_289);
nand U1095 (N_1095,N_80,N_470);
nand U1096 (N_1096,N_208,N_663);
nand U1097 (N_1097,N_491,N_178);
and U1098 (N_1098,N_44,N_215);
and U1099 (N_1099,N_403,N_356);
or U1100 (N_1100,N_717,N_106);
and U1101 (N_1101,N_280,N_338);
or U1102 (N_1102,N_243,N_95);
nor U1103 (N_1103,N_723,N_323);
and U1104 (N_1104,N_675,N_409);
or U1105 (N_1105,N_414,N_391);
nand U1106 (N_1106,N_285,N_377);
nor U1107 (N_1107,N_404,N_104);
nand U1108 (N_1108,N_624,N_616);
nand U1109 (N_1109,N_555,N_25);
nor U1110 (N_1110,N_585,N_59);
or U1111 (N_1111,N_120,N_12);
nand U1112 (N_1112,N_481,N_635);
or U1113 (N_1113,N_234,N_54);
nand U1114 (N_1114,N_398,N_535);
nand U1115 (N_1115,N_328,N_478);
and U1116 (N_1116,N_278,N_307);
nand U1117 (N_1117,N_235,N_53);
and U1118 (N_1118,N_159,N_211);
nor U1119 (N_1119,N_222,N_735);
or U1120 (N_1120,N_51,N_205);
nand U1121 (N_1121,N_664,N_237);
nand U1122 (N_1122,N_467,N_368);
or U1123 (N_1123,N_308,N_533);
nand U1124 (N_1124,N_466,N_638);
nor U1125 (N_1125,N_571,N_695);
nor U1126 (N_1126,N_186,N_109);
nand U1127 (N_1127,N_81,N_239);
nor U1128 (N_1128,N_564,N_647);
nor U1129 (N_1129,N_262,N_548);
or U1130 (N_1130,N_533,N_732);
nor U1131 (N_1131,N_335,N_381);
and U1132 (N_1132,N_166,N_124);
or U1133 (N_1133,N_553,N_238);
nor U1134 (N_1134,N_466,N_714);
and U1135 (N_1135,N_474,N_227);
or U1136 (N_1136,N_712,N_174);
nand U1137 (N_1137,N_669,N_278);
nand U1138 (N_1138,N_282,N_682);
nand U1139 (N_1139,N_237,N_178);
and U1140 (N_1140,N_35,N_637);
or U1141 (N_1141,N_392,N_546);
nor U1142 (N_1142,N_721,N_290);
and U1143 (N_1143,N_390,N_47);
or U1144 (N_1144,N_539,N_528);
nand U1145 (N_1145,N_529,N_649);
and U1146 (N_1146,N_378,N_40);
and U1147 (N_1147,N_663,N_571);
and U1148 (N_1148,N_123,N_526);
nor U1149 (N_1149,N_511,N_43);
and U1150 (N_1150,N_179,N_11);
nand U1151 (N_1151,N_23,N_639);
nor U1152 (N_1152,N_442,N_417);
nor U1153 (N_1153,N_8,N_716);
nor U1154 (N_1154,N_676,N_416);
nand U1155 (N_1155,N_337,N_739);
nand U1156 (N_1156,N_268,N_590);
nand U1157 (N_1157,N_601,N_415);
nand U1158 (N_1158,N_619,N_61);
and U1159 (N_1159,N_553,N_314);
or U1160 (N_1160,N_48,N_328);
and U1161 (N_1161,N_612,N_714);
or U1162 (N_1162,N_183,N_473);
nor U1163 (N_1163,N_405,N_267);
or U1164 (N_1164,N_157,N_744);
and U1165 (N_1165,N_465,N_297);
nor U1166 (N_1166,N_192,N_102);
and U1167 (N_1167,N_490,N_303);
nand U1168 (N_1168,N_578,N_473);
nor U1169 (N_1169,N_724,N_469);
nand U1170 (N_1170,N_426,N_261);
nor U1171 (N_1171,N_441,N_3);
nor U1172 (N_1172,N_11,N_210);
nand U1173 (N_1173,N_386,N_562);
or U1174 (N_1174,N_609,N_492);
nor U1175 (N_1175,N_316,N_535);
nand U1176 (N_1176,N_420,N_15);
and U1177 (N_1177,N_378,N_728);
and U1178 (N_1178,N_245,N_220);
and U1179 (N_1179,N_526,N_365);
nand U1180 (N_1180,N_119,N_17);
nor U1181 (N_1181,N_366,N_682);
and U1182 (N_1182,N_152,N_16);
or U1183 (N_1183,N_713,N_499);
or U1184 (N_1184,N_421,N_550);
or U1185 (N_1185,N_262,N_507);
nor U1186 (N_1186,N_163,N_173);
and U1187 (N_1187,N_331,N_201);
nand U1188 (N_1188,N_199,N_306);
or U1189 (N_1189,N_431,N_736);
nor U1190 (N_1190,N_702,N_150);
nor U1191 (N_1191,N_17,N_187);
or U1192 (N_1192,N_58,N_59);
xor U1193 (N_1193,N_59,N_83);
nand U1194 (N_1194,N_452,N_93);
nand U1195 (N_1195,N_31,N_433);
and U1196 (N_1196,N_410,N_100);
nor U1197 (N_1197,N_183,N_47);
nand U1198 (N_1198,N_75,N_155);
or U1199 (N_1199,N_684,N_495);
nand U1200 (N_1200,N_714,N_364);
nand U1201 (N_1201,N_603,N_667);
and U1202 (N_1202,N_289,N_330);
nand U1203 (N_1203,N_258,N_541);
and U1204 (N_1204,N_490,N_744);
nor U1205 (N_1205,N_384,N_126);
nor U1206 (N_1206,N_494,N_1);
nor U1207 (N_1207,N_300,N_541);
nand U1208 (N_1208,N_377,N_380);
and U1209 (N_1209,N_294,N_476);
nor U1210 (N_1210,N_290,N_12);
or U1211 (N_1211,N_527,N_148);
or U1212 (N_1212,N_389,N_656);
or U1213 (N_1213,N_378,N_307);
nor U1214 (N_1214,N_553,N_324);
and U1215 (N_1215,N_162,N_695);
and U1216 (N_1216,N_235,N_237);
nand U1217 (N_1217,N_218,N_677);
or U1218 (N_1218,N_71,N_103);
nand U1219 (N_1219,N_275,N_473);
nand U1220 (N_1220,N_43,N_238);
and U1221 (N_1221,N_477,N_349);
or U1222 (N_1222,N_157,N_8);
nand U1223 (N_1223,N_616,N_552);
and U1224 (N_1224,N_379,N_189);
and U1225 (N_1225,N_382,N_590);
nand U1226 (N_1226,N_606,N_398);
and U1227 (N_1227,N_490,N_673);
and U1228 (N_1228,N_59,N_484);
nor U1229 (N_1229,N_163,N_574);
nor U1230 (N_1230,N_293,N_647);
nor U1231 (N_1231,N_249,N_688);
or U1232 (N_1232,N_696,N_429);
xor U1233 (N_1233,N_295,N_416);
nand U1234 (N_1234,N_433,N_75);
nor U1235 (N_1235,N_366,N_235);
nor U1236 (N_1236,N_660,N_579);
nor U1237 (N_1237,N_223,N_386);
or U1238 (N_1238,N_123,N_426);
nor U1239 (N_1239,N_743,N_131);
or U1240 (N_1240,N_607,N_20);
nand U1241 (N_1241,N_22,N_449);
and U1242 (N_1242,N_712,N_196);
nand U1243 (N_1243,N_192,N_191);
or U1244 (N_1244,N_662,N_698);
and U1245 (N_1245,N_563,N_130);
nor U1246 (N_1246,N_110,N_454);
nand U1247 (N_1247,N_476,N_117);
or U1248 (N_1248,N_482,N_175);
or U1249 (N_1249,N_68,N_118);
nor U1250 (N_1250,N_480,N_570);
nor U1251 (N_1251,N_379,N_577);
or U1252 (N_1252,N_58,N_711);
nor U1253 (N_1253,N_635,N_201);
or U1254 (N_1254,N_336,N_32);
or U1255 (N_1255,N_674,N_68);
or U1256 (N_1256,N_537,N_610);
nor U1257 (N_1257,N_171,N_464);
or U1258 (N_1258,N_626,N_4);
nand U1259 (N_1259,N_252,N_255);
and U1260 (N_1260,N_236,N_163);
nor U1261 (N_1261,N_404,N_235);
nand U1262 (N_1262,N_641,N_735);
or U1263 (N_1263,N_484,N_692);
and U1264 (N_1264,N_529,N_742);
nand U1265 (N_1265,N_440,N_720);
nand U1266 (N_1266,N_314,N_352);
or U1267 (N_1267,N_433,N_543);
nand U1268 (N_1268,N_568,N_567);
and U1269 (N_1269,N_28,N_354);
and U1270 (N_1270,N_179,N_518);
nor U1271 (N_1271,N_36,N_457);
and U1272 (N_1272,N_250,N_329);
or U1273 (N_1273,N_386,N_266);
nand U1274 (N_1274,N_551,N_498);
or U1275 (N_1275,N_430,N_239);
or U1276 (N_1276,N_452,N_657);
nand U1277 (N_1277,N_524,N_620);
nand U1278 (N_1278,N_255,N_6);
or U1279 (N_1279,N_217,N_317);
nor U1280 (N_1280,N_512,N_642);
or U1281 (N_1281,N_154,N_130);
nor U1282 (N_1282,N_537,N_211);
nand U1283 (N_1283,N_628,N_506);
nor U1284 (N_1284,N_595,N_418);
and U1285 (N_1285,N_664,N_37);
or U1286 (N_1286,N_363,N_396);
nand U1287 (N_1287,N_430,N_742);
nor U1288 (N_1288,N_460,N_159);
or U1289 (N_1289,N_519,N_305);
and U1290 (N_1290,N_340,N_625);
nand U1291 (N_1291,N_551,N_572);
nor U1292 (N_1292,N_575,N_374);
or U1293 (N_1293,N_14,N_523);
and U1294 (N_1294,N_745,N_506);
nand U1295 (N_1295,N_500,N_555);
or U1296 (N_1296,N_492,N_151);
and U1297 (N_1297,N_171,N_51);
nand U1298 (N_1298,N_110,N_96);
nor U1299 (N_1299,N_390,N_337);
and U1300 (N_1300,N_378,N_123);
or U1301 (N_1301,N_462,N_13);
nand U1302 (N_1302,N_241,N_486);
or U1303 (N_1303,N_422,N_40);
nand U1304 (N_1304,N_390,N_694);
nor U1305 (N_1305,N_468,N_519);
and U1306 (N_1306,N_478,N_595);
and U1307 (N_1307,N_126,N_449);
or U1308 (N_1308,N_58,N_141);
nor U1309 (N_1309,N_452,N_32);
nand U1310 (N_1310,N_188,N_535);
nor U1311 (N_1311,N_533,N_655);
nor U1312 (N_1312,N_131,N_174);
nand U1313 (N_1313,N_735,N_480);
nor U1314 (N_1314,N_333,N_64);
xor U1315 (N_1315,N_556,N_568);
nand U1316 (N_1316,N_96,N_594);
and U1317 (N_1317,N_258,N_169);
or U1318 (N_1318,N_584,N_392);
xnor U1319 (N_1319,N_318,N_177);
nor U1320 (N_1320,N_292,N_472);
or U1321 (N_1321,N_546,N_23);
or U1322 (N_1322,N_713,N_477);
nand U1323 (N_1323,N_396,N_637);
and U1324 (N_1324,N_319,N_360);
and U1325 (N_1325,N_200,N_742);
and U1326 (N_1326,N_499,N_257);
and U1327 (N_1327,N_298,N_30);
and U1328 (N_1328,N_226,N_499);
nand U1329 (N_1329,N_384,N_67);
xor U1330 (N_1330,N_194,N_698);
and U1331 (N_1331,N_127,N_145);
nand U1332 (N_1332,N_622,N_31);
or U1333 (N_1333,N_610,N_49);
xnor U1334 (N_1334,N_180,N_237);
nand U1335 (N_1335,N_600,N_212);
nand U1336 (N_1336,N_572,N_389);
nor U1337 (N_1337,N_696,N_304);
nand U1338 (N_1338,N_652,N_72);
nor U1339 (N_1339,N_97,N_553);
or U1340 (N_1340,N_94,N_527);
nand U1341 (N_1341,N_252,N_746);
and U1342 (N_1342,N_229,N_413);
and U1343 (N_1343,N_375,N_190);
xor U1344 (N_1344,N_377,N_114);
nand U1345 (N_1345,N_5,N_456);
nor U1346 (N_1346,N_439,N_312);
and U1347 (N_1347,N_307,N_305);
or U1348 (N_1348,N_398,N_457);
and U1349 (N_1349,N_440,N_54);
nor U1350 (N_1350,N_310,N_747);
and U1351 (N_1351,N_654,N_562);
or U1352 (N_1352,N_190,N_161);
nand U1353 (N_1353,N_656,N_460);
or U1354 (N_1354,N_155,N_198);
nor U1355 (N_1355,N_401,N_379);
nor U1356 (N_1356,N_474,N_297);
and U1357 (N_1357,N_239,N_300);
nor U1358 (N_1358,N_343,N_140);
or U1359 (N_1359,N_35,N_327);
or U1360 (N_1360,N_385,N_370);
nor U1361 (N_1361,N_540,N_623);
or U1362 (N_1362,N_85,N_180);
xor U1363 (N_1363,N_531,N_218);
or U1364 (N_1364,N_579,N_38);
nor U1365 (N_1365,N_726,N_144);
nor U1366 (N_1366,N_183,N_155);
nand U1367 (N_1367,N_104,N_246);
nor U1368 (N_1368,N_206,N_261);
and U1369 (N_1369,N_592,N_693);
nor U1370 (N_1370,N_744,N_638);
nor U1371 (N_1371,N_624,N_422);
nor U1372 (N_1372,N_280,N_703);
nand U1373 (N_1373,N_264,N_116);
nor U1374 (N_1374,N_133,N_440);
nand U1375 (N_1375,N_2,N_678);
or U1376 (N_1376,N_120,N_240);
or U1377 (N_1377,N_297,N_57);
nand U1378 (N_1378,N_402,N_508);
and U1379 (N_1379,N_606,N_254);
and U1380 (N_1380,N_141,N_226);
nand U1381 (N_1381,N_446,N_703);
nand U1382 (N_1382,N_711,N_698);
or U1383 (N_1383,N_678,N_635);
nand U1384 (N_1384,N_202,N_481);
nor U1385 (N_1385,N_662,N_599);
or U1386 (N_1386,N_316,N_559);
and U1387 (N_1387,N_377,N_454);
or U1388 (N_1388,N_357,N_642);
nor U1389 (N_1389,N_412,N_308);
nor U1390 (N_1390,N_375,N_10);
nor U1391 (N_1391,N_518,N_267);
nand U1392 (N_1392,N_635,N_590);
nor U1393 (N_1393,N_723,N_187);
and U1394 (N_1394,N_509,N_54);
and U1395 (N_1395,N_159,N_88);
and U1396 (N_1396,N_112,N_66);
and U1397 (N_1397,N_466,N_494);
and U1398 (N_1398,N_258,N_746);
or U1399 (N_1399,N_173,N_625);
and U1400 (N_1400,N_453,N_690);
nor U1401 (N_1401,N_636,N_264);
nor U1402 (N_1402,N_516,N_157);
or U1403 (N_1403,N_528,N_47);
nand U1404 (N_1404,N_278,N_543);
and U1405 (N_1405,N_391,N_142);
nor U1406 (N_1406,N_212,N_34);
and U1407 (N_1407,N_360,N_439);
nor U1408 (N_1408,N_598,N_564);
or U1409 (N_1409,N_125,N_726);
nand U1410 (N_1410,N_372,N_331);
nand U1411 (N_1411,N_575,N_17);
nand U1412 (N_1412,N_319,N_559);
nor U1413 (N_1413,N_498,N_224);
and U1414 (N_1414,N_687,N_350);
nor U1415 (N_1415,N_575,N_172);
and U1416 (N_1416,N_382,N_0);
nor U1417 (N_1417,N_88,N_123);
and U1418 (N_1418,N_450,N_685);
nor U1419 (N_1419,N_326,N_569);
or U1420 (N_1420,N_433,N_404);
nor U1421 (N_1421,N_108,N_280);
or U1422 (N_1422,N_369,N_522);
and U1423 (N_1423,N_731,N_438);
or U1424 (N_1424,N_613,N_189);
and U1425 (N_1425,N_513,N_655);
or U1426 (N_1426,N_736,N_527);
or U1427 (N_1427,N_483,N_330);
and U1428 (N_1428,N_98,N_247);
or U1429 (N_1429,N_86,N_579);
or U1430 (N_1430,N_737,N_521);
or U1431 (N_1431,N_162,N_310);
and U1432 (N_1432,N_290,N_748);
nor U1433 (N_1433,N_97,N_399);
nor U1434 (N_1434,N_15,N_603);
nand U1435 (N_1435,N_445,N_127);
or U1436 (N_1436,N_43,N_201);
and U1437 (N_1437,N_394,N_450);
and U1438 (N_1438,N_106,N_449);
nand U1439 (N_1439,N_692,N_424);
or U1440 (N_1440,N_239,N_147);
nand U1441 (N_1441,N_635,N_570);
nor U1442 (N_1442,N_326,N_386);
or U1443 (N_1443,N_536,N_278);
nand U1444 (N_1444,N_674,N_607);
xnor U1445 (N_1445,N_562,N_406);
xnor U1446 (N_1446,N_398,N_373);
nor U1447 (N_1447,N_164,N_627);
and U1448 (N_1448,N_391,N_15);
nor U1449 (N_1449,N_110,N_602);
nand U1450 (N_1450,N_320,N_61);
nor U1451 (N_1451,N_666,N_691);
or U1452 (N_1452,N_431,N_84);
nor U1453 (N_1453,N_9,N_19);
nand U1454 (N_1454,N_671,N_586);
or U1455 (N_1455,N_646,N_573);
nor U1456 (N_1456,N_226,N_228);
nor U1457 (N_1457,N_541,N_5);
nor U1458 (N_1458,N_192,N_142);
nand U1459 (N_1459,N_503,N_360);
nor U1460 (N_1460,N_347,N_613);
nand U1461 (N_1461,N_541,N_281);
or U1462 (N_1462,N_16,N_610);
nor U1463 (N_1463,N_15,N_739);
nand U1464 (N_1464,N_312,N_69);
and U1465 (N_1465,N_468,N_625);
and U1466 (N_1466,N_538,N_533);
nor U1467 (N_1467,N_460,N_545);
nand U1468 (N_1468,N_102,N_520);
nor U1469 (N_1469,N_6,N_67);
and U1470 (N_1470,N_712,N_277);
nand U1471 (N_1471,N_427,N_599);
or U1472 (N_1472,N_82,N_532);
nor U1473 (N_1473,N_576,N_55);
nor U1474 (N_1474,N_637,N_583);
nand U1475 (N_1475,N_35,N_440);
nand U1476 (N_1476,N_136,N_266);
nor U1477 (N_1477,N_55,N_473);
nand U1478 (N_1478,N_336,N_352);
nor U1479 (N_1479,N_609,N_625);
or U1480 (N_1480,N_631,N_146);
nand U1481 (N_1481,N_747,N_482);
nand U1482 (N_1482,N_171,N_200);
and U1483 (N_1483,N_257,N_575);
and U1484 (N_1484,N_469,N_190);
or U1485 (N_1485,N_76,N_250);
or U1486 (N_1486,N_45,N_470);
nor U1487 (N_1487,N_49,N_449);
or U1488 (N_1488,N_286,N_0);
nor U1489 (N_1489,N_156,N_569);
or U1490 (N_1490,N_193,N_268);
nor U1491 (N_1491,N_539,N_566);
nand U1492 (N_1492,N_281,N_74);
nand U1493 (N_1493,N_36,N_141);
nor U1494 (N_1494,N_555,N_306);
nor U1495 (N_1495,N_346,N_720);
and U1496 (N_1496,N_553,N_520);
nand U1497 (N_1497,N_485,N_172);
or U1498 (N_1498,N_289,N_463);
nand U1499 (N_1499,N_323,N_377);
and U1500 (N_1500,N_1027,N_1482);
nand U1501 (N_1501,N_860,N_1367);
or U1502 (N_1502,N_1360,N_1095);
or U1503 (N_1503,N_1480,N_1340);
or U1504 (N_1504,N_801,N_1311);
nor U1505 (N_1505,N_777,N_789);
and U1506 (N_1506,N_1299,N_1026);
and U1507 (N_1507,N_1384,N_1054);
nor U1508 (N_1508,N_804,N_1020);
or U1509 (N_1509,N_1289,N_1465);
nor U1510 (N_1510,N_918,N_1010);
and U1511 (N_1511,N_969,N_1405);
or U1512 (N_1512,N_1427,N_1454);
nor U1513 (N_1513,N_1025,N_1323);
nand U1514 (N_1514,N_822,N_1392);
or U1515 (N_1515,N_1217,N_1463);
nand U1516 (N_1516,N_1260,N_857);
or U1517 (N_1517,N_1479,N_922);
or U1518 (N_1518,N_1279,N_799);
or U1519 (N_1519,N_1182,N_869);
xnor U1520 (N_1520,N_1146,N_941);
and U1521 (N_1521,N_940,N_1346);
and U1522 (N_1522,N_1021,N_1317);
nand U1523 (N_1523,N_1046,N_768);
nor U1524 (N_1524,N_1339,N_1113);
and U1525 (N_1525,N_946,N_1361);
nand U1526 (N_1526,N_817,N_1183);
or U1527 (N_1527,N_1188,N_1321);
nor U1528 (N_1528,N_938,N_1449);
and U1529 (N_1529,N_805,N_1036);
nand U1530 (N_1530,N_1483,N_1137);
nor U1531 (N_1531,N_1160,N_1022);
nand U1532 (N_1532,N_1013,N_928);
nand U1533 (N_1533,N_1038,N_919);
nor U1534 (N_1534,N_1017,N_1214);
and U1535 (N_1535,N_1060,N_1162);
or U1536 (N_1536,N_1322,N_1108);
and U1537 (N_1537,N_1207,N_1399);
nor U1538 (N_1538,N_983,N_1152);
nand U1539 (N_1539,N_1167,N_1104);
nor U1540 (N_1540,N_1276,N_1144);
nor U1541 (N_1541,N_926,N_1381);
and U1542 (N_1542,N_925,N_1460);
nand U1543 (N_1543,N_1375,N_942);
nand U1544 (N_1544,N_826,N_1351);
and U1545 (N_1545,N_1268,N_1073);
and U1546 (N_1546,N_1007,N_836);
or U1547 (N_1547,N_1139,N_828);
and U1548 (N_1548,N_782,N_855);
and U1549 (N_1549,N_1109,N_1030);
or U1550 (N_1550,N_1261,N_1034);
and U1551 (N_1551,N_1206,N_1239);
or U1552 (N_1552,N_1065,N_1135);
and U1553 (N_1553,N_1028,N_1131);
or U1554 (N_1554,N_820,N_787);
and U1555 (N_1555,N_1213,N_1082);
nand U1556 (N_1556,N_1049,N_997);
nor U1557 (N_1557,N_1499,N_1096);
nor U1558 (N_1558,N_1481,N_792);
and U1559 (N_1559,N_1349,N_793);
or U1560 (N_1560,N_1259,N_1331);
or U1561 (N_1561,N_770,N_963);
and U1562 (N_1562,N_1438,N_1343);
nand U1563 (N_1563,N_1488,N_1379);
and U1564 (N_1564,N_883,N_877);
nor U1565 (N_1565,N_1337,N_1016);
nand U1566 (N_1566,N_923,N_952);
nand U1567 (N_1567,N_1423,N_1411);
and U1568 (N_1568,N_1408,N_1232);
and U1569 (N_1569,N_1040,N_1055);
nor U1570 (N_1570,N_1413,N_1225);
and U1571 (N_1571,N_1426,N_1295);
or U1572 (N_1572,N_1448,N_1453);
and U1573 (N_1573,N_962,N_1132);
xor U1574 (N_1574,N_1332,N_898);
nor U1575 (N_1575,N_866,N_1456);
and U1576 (N_1576,N_846,N_996);
and U1577 (N_1577,N_1461,N_1292);
or U1578 (N_1578,N_861,N_813);
xor U1579 (N_1579,N_1378,N_1068);
nand U1580 (N_1580,N_998,N_1478);
nand U1581 (N_1581,N_1236,N_1165);
or U1582 (N_1582,N_859,N_1249);
and U1583 (N_1583,N_1111,N_1296);
nor U1584 (N_1584,N_1352,N_825);
or U1585 (N_1585,N_881,N_934);
and U1586 (N_1586,N_1059,N_1126);
nor U1587 (N_1587,N_1310,N_1372);
or U1588 (N_1588,N_1210,N_958);
nor U1589 (N_1589,N_1254,N_988);
or U1590 (N_1590,N_901,N_1127);
or U1591 (N_1591,N_1269,N_1284);
and U1592 (N_1592,N_882,N_1312);
and U1593 (N_1593,N_790,N_823);
nand U1594 (N_1594,N_1324,N_1297);
nand U1595 (N_1595,N_975,N_1195);
nor U1596 (N_1596,N_762,N_1286);
or U1597 (N_1597,N_1386,N_1318);
and U1598 (N_1598,N_989,N_896);
nor U1599 (N_1599,N_1475,N_1134);
nor U1600 (N_1600,N_786,N_798);
and U1601 (N_1601,N_1319,N_1198);
nor U1602 (N_1602,N_1099,N_999);
and U1603 (N_1603,N_1485,N_1425);
nor U1604 (N_1604,N_917,N_1204);
nor U1605 (N_1605,N_900,N_1490);
or U1606 (N_1606,N_1177,N_1442);
nor U1607 (N_1607,N_1042,N_1450);
nor U1608 (N_1608,N_1181,N_1000);
or U1609 (N_1609,N_1409,N_890);
nand U1610 (N_1610,N_756,N_1285);
and U1611 (N_1611,N_1302,N_1117);
nand U1612 (N_1612,N_842,N_1307);
nor U1613 (N_1613,N_839,N_1470);
xnor U1614 (N_1614,N_1124,N_1262);
or U1615 (N_1615,N_815,N_1180);
nor U1616 (N_1616,N_1061,N_1084);
nor U1617 (N_1617,N_929,N_864);
nor U1618 (N_1618,N_1057,N_1193);
nor U1619 (N_1619,N_819,N_1230);
or U1620 (N_1620,N_806,N_1265);
or U1621 (N_1621,N_897,N_1176);
nor U1622 (N_1622,N_784,N_1178);
and U1623 (N_1623,N_1467,N_1257);
or U1624 (N_1624,N_879,N_847);
and U1625 (N_1625,N_1190,N_1489);
and U1626 (N_1626,N_1150,N_916);
nor U1627 (N_1627,N_830,N_763);
nor U1628 (N_1628,N_1451,N_1304);
nor U1629 (N_1629,N_1251,N_1224);
nor U1630 (N_1630,N_1002,N_1086);
or U1631 (N_1631,N_755,N_1044);
nor U1632 (N_1632,N_1138,N_1412);
nand U1633 (N_1633,N_1171,N_892);
nand U1634 (N_1634,N_1258,N_921);
or U1635 (N_1635,N_1174,N_886);
nor U1636 (N_1636,N_1415,N_850);
and U1637 (N_1637,N_1334,N_1282);
nand U1638 (N_1638,N_785,N_1091);
or U1639 (N_1639,N_1147,N_1356);
nand U1640 (N_1640,N_1353,N_1402);
nor U1641 (N_1641,N_1266,N_1389);
nor U1642 (N_1642,N_1358,N_1443);
nor U1643 (N_1643,N_987,N_1371);
or U1644 (N_1644,N_1446,N_1458);
nor U1645 (N_1645,N_1306,N_1393);
nand U1646 (N_1646,N_788,N_1434);
and U1647 (N_1647,N_1233,N_1281);
nand U1648 (N_1648,N_1058,N_1106);
or U1649 (N_1649,N_870,N_875);
and U1650 (N_1650,N_1047,N_829);
nor U1651 (N_1651,N_761,N_1118);
nand U1652 (N_1652,N_1243,N_1220);
and U1653 (N_1653,N_1078,N_1001);
and U1654 (N_1654,N_1394,N_1368);
or U1655 (N_1655,N_1255,N_978);
nand U1656 (N_1656,N_769,N_1094);
xor U1657 (N_1657,N_1202,N_956);
nand U1658 (N_1658,N_1487,N_947);
nand U1659 (N_1659,N_994,N_1102);
or U1660 (N_1660,N_1336,N_802);
or U1661 (N_1661,N_1264,N_764);
or U1662 (N_1662,N_1459,N_849);
nand U1663 (N_1663,N_1492,N_1064);
nand U1664 (N_1664,N_796,N_1246);
and U1665 (N_1665,N_1287,N_1215);
nand U1666 (N_1666,N_1237,N_1031);
and U1667 (N_1667,N_1397,N_1452);
or U1668 (N_1668,N_1056,N_863);
or U1669 (N_1669,N_1313,N_1221);
or U1670 (N_1670,N_1029,N_818);
nor U1671 (N_1671,N_1329,N_1196);
nand U1672 (N_1672,N_903,N_1283);
nor U1673 (N_1673,N_1330,N_1420);
and U1674 (N_1674,N_930,N_1345);
and U1675 (N_1675,N_1477,N_1218);
nor U1676 (N_1676,N_1473,N_1173);
nand U1677 (N_1677,N_972,N_1199);
nand U1678 (N_1678,N_1179,N_884);
nor U1679 (N_1679,N_1129,N_1350);
or U1680 (N_1680,N_1417,N_1149);
and U1681 (N_1681,N_812,N_1348);
or U1682 (N_1682,N_1377,N_1400);
and U1683 (N_1683,N_1308,N_1163);
nor U1684 (N_1684,N_1153,N_911);
and U1685 (N_1685,N_1075,N_772);
nand U1686 (N_1686,N_1018,N_867);
and U1687 (N_1687,N_1497,N_1275);
or U1688 (N_1688,N_1341,N_774);
nand U1689 (N_1689,N_1403,N_835);
nand U1690 (N_1690,N_1303,N_979);
nand U1691 (N_1691,N_1320,N_1226);
and U1692 (N_1692,N_780,N_1364);
nor U1693 (N_1693,N_1316,N_1491);
nor U1694 (N_1694,N_1326,N_1291);
nor U1695 (N_1695,N_1376,N_1229);
nor U1696 (N_1696,N_943,N_1192);
nor U1697 (N_1697,N_1051,N_845);
and U1698 (N_1698,N_1374,N_1436);
and U1699 (N_1699,N_1290,N_853);
nor U1700 (N_1700,N_871,N_1164);
and U1701 (N_1701,N_808,N_1333);
and U1702 (N_1702,N_1114,N_807);
nor U1703 (N_1703,N_937,N_1033);
xor U1704 (N_1704,N_1032,N_1466);
and U1705 (N_1705,N_1133,N_971);
nand U1706 (N_1706,N_1252,N_779);
or U1707 (N_1707,N_1216,N_1205);
nor U1708 (N_1708,N_862,N_1039);
nor U1709 (N_1709,N_1315,N_1327);
nor U1710 (N_1710,N_1245,N_776);
or U1711 (N_1711,N_876,N_1136);
nor U1712 (N_1712,N_1247,N_1370);
nand U1713 (N_1713,N_980,N_904);
nand U1714 (N_1714,N_873,N_1219);
nand U1715 (N_1715,N_909,N_1043);
nand U1716 (N_1716,N_984,N_1369);
nand U1717 (N_1717,N_1242,N_887);
nor U1718 (N_1718,N_1066,N_1309);
xnor U1719 (N_1719,N_1140,N_991);
or U1720 (N_1720,N_1416,N_1401);
or U1721 (N_1721,N_1231,N_844);
and U1722 (N_1722,N_1170,N_1083);
or U1723 (N_1723,N_810,N_1168);
nand U1724 (N_1724,N_1090,N_1155);
nor U1725 (N_1725,N_1298,N_955);
and U1726 (N_1726,N_1169,N_995);
nand U1727 (N_1727,N_1186,N_843);
nor U1728 (N_1728,N_1484,N_1263);
nor U1729 (N_1729,N_791,N_1410);
and U1730 (N_1730,N_1203,N_905);
nand U1731 (N_1731,N_1277,N_1390);
and U1732 (N_1732,N_1241,N_990);
or U1733 (N_1733,N_949,N_1305);
nor U1734 (N_1734,N_1363,N_1457);
nand U1735 (N_1735,N_977,N_753);
nor U1736 (N_1736,N_1278,N_1359);
and U1737 (N_1737,N_1079,N_950);
nand U1738 (N_1738,N_854,N_982);
or U1739 (N_1739,N_1256,N_1175);
and U1740 (N_1740,N_765,N_1209);
nor U1741 (N_1741,N_773,N_771);
nor U1742 (N_1742,N_1081,N_1151);
nor U1743 (N_1743,N_1354,N_1435);
and U1744 (N_1744,N_1159,N_874);
nand U1745 (N_1745,N_1471,N_976);
nor U1746 (N_1746,N_920,N_1077);
and U1747 (N_1747,N_1430,N_1223);
and U1748 (N_1748,N_1328,N_910);
or U1749 (N_1749,N_1142,N_915);
and U1750 (N_1750,N_833,N_851);
nand U1751 (N_1751,N_852,N_1143);
nand U1752 (N_1752,N_1469,N_1112);
nor U1753 (N_1753,N_766,N_841);
nand U1754 (N_1754,N_993,N_757);
nor U1755 (N_1755,N_1468,N_1357);
xor U1756 (N_1756,N_1105,N_775);
or U1757 (N_1757,N_1432,N_778);
nand U1758 (N_1758,N_1080,N_1464);
and U1759 (N_1759,N_1293,N_1158);
nor U1760 (N_1760,N_1383,N_1071);
nor U1761 (N_1761,N_1200,N_1005);
nand U1762 (N_1762,N_960,N_927);
or U1763 (N_1763,N_935,N_1062);
nand U1764 (N_1764,N_1141,N_1366);
nor U1765 (N_1765,N_1493,N_795);
or U1766 (N_1766,N_809,N_1355);
nor U1767 (N_1767,N_1486,N_1053);
nor U1768 (N_1768,N_1387,N_961);
nor U1769 (N_1769,N_1006,N_1280);
xnor U1770 (N_1770,N_1414,N_974);
nand U1771 (N_1771,N_1398,N_939);
nand U1772 (N_1772,N_959,N_1385);
and U1773 (N_1773,N_895,N_1267);
and U1774 (N_1774,N_936,N_1063);
or U1775 (N_1775,N_1373,N_781);
and U1776 (N_1776,N_824,N_1388);
and U1777 (N_1777,N_1212,N_1498);
or U1778 (N_1778,N_889,N_783);
and U1779 (N_1779,N_1098,N_1120);
and U1780 (N_1780,N_894,N_1428);
xor U1781 (N_1781,N_1197,N_1072);
nand U1782 (N_1782,N_1093,N_1211);
or U1783 (N_1783,N_1494,N_1050);
and U1784 (N_1784,N_1271,N_1122);
and U1785 (N_1785,N_1208,N_1148);
or U1786 (N_1786,N_908,N_957);
or U1787 (N_1787,N_1130,N_1110);
and U1788 (N_1788,N_1391,N_1100);
nor U1789 (N_1789,N_1496,N_803);
nor U1790 (N_1790,N_1070,N_902);
nand U1791 (N_1791,N_1194,N_992);
or U1792 (N_1792,N_931,N_1419);
or U1793 (N_1793,N_953,N_891);
or U1794 (N_1794,N_924,N_1441);
nor U1795 (N_1795,N_885,N_1092);
nor U1796 (N_1796,N_933,N_1250);
nand U1797 (N_1797,N_1003,N_1455);
or U1798 (N_1798,N_1019,N_868);
and U1799 (N_1799,N_794,N_1116);
nand U1800 (N_1800,N_821,N_985);
nand U1801 (N_1801,N_1395,N_1396);
and U1802 (N_1802,N_1088,N_1037);
and U1803 (N_1803,N_1288,N_1014);
and U1804 (N_1804,N_750,N_1362);
or U1805 (N_1805,N_1103,N_964);
or U1806 (N_1806,N_1445,N_913);
or U1807 (N_1807,N_951,N_751);
and U1808 (N_1808,N_759,N_1009);
nor U1809 (N_1809,N_1069,N_1495);
nor U1810 (N_1810,N_797,N_948);
nor U1811 (N_1811,N_1234,N_1472);
nor U1812 (N_1812,N_1052,N_1347);
nand U1813 (N_1813,N_1335,N_1023);
nor U1814 (N_1814,N_1128,N_1429);
or U1815 (N_1815,N_1041,N_1067);
nor U1816 (N_1816,N_1097,N_1365);
or U1817 (N_1817,N_837,N_970);
nor U1818 (N_1818,N_1300,N_832);
nand U1819 (N_1819,N_1240,N_834);
and U1820 (N_1820,N_893,N_1440);
or U1821 (N_1821,N_1166,N_752);
nor U1822 (N_1822,N_838,N_1107);
nor U1823 (N_1823,N_1074,N_1338);
nor U1824 (N_1824,N_856,N_814);
and U1825 (N_1825,N_932,N_1121);
nor U1826 (N_1826,N_1462,N_912);
nor U1827 (N_1827,N_1184,N_1314);
or U1828 (N_1828,N_1228,N_827);
nand U1829 (N_1829,N_965,N_1406);
nor U1830 (N_1830,N_1185,N_1447);
nor U1831 (N_1831,N_1422,N_1476);
and U1832 (N_1832,N_1087,N_865);
and U1833 (N_1833,N_872,N_1235);
or U1834 (N_1834,N_858,N_1344);
nor U1835 (N_1835,N_1156,N_981);
nor U1836 (N_1836,N_754,N_1101);
or U1837 (N_1837,N_1011,N_1189);
and U1838 (N_1838,N_1172,N_1418);
and U1839 (N_1839,N_1125,N_1008);
nand U1840 (N_1840,N_1145,N_1238);
or U1841 (N_1841,N_1301,N_1407);
or U1842 (N_1842,N_914,N_1187);
nand U1843 (N_1843,N_1444,N_1157);
nand U1844 (N_1844,N_758,N_1274);
and U1845 (N_1845,N_1474,N_1439);
and U1846 (N_1846,N_1045,N_1272);
and U1847 (N_1847,N_1015,N_1342);
and U1848 (N_1848,N_878,N_1201);
nor U1849 (N_1849,N_1123,N_907);
or U1850 (N_1850,N_880,N_1012);
or U1851 (N_1851,N_1085,N_1076);
and U1852 (N_1852,N_1431,N_899);
or U1853 (N_1853,N_840,N_906);
or U1854 (N_1854,N_1433,N_1089);
and U1855 (N_1855,N_1253,N_1244);
nor U1856 (N_1856,N_1024,N_1248);
xnor U1857 (N_1857,N_1048,N_1404);
xnor U1858 (N_1858,N_1380,N_1154);
nor U1859 (N_1859,N_1161,N_1382);
and U1860 (N_1860,N_1115,N_954);
nor U1861 (N_1861,N_1325,N_816);
and U1862 (N_1862,N_767,N_1294);
xnor U1863 (N_1863,N_1191,N_848);
and U1864 (N_1864,N_811,N_968);
xnor U1865 (N_1865,N_1119,N_800);
nor U1866 (N_1866,N_966,N_973);
and U1867 (N_1867,N_888,N_760);
nand U1868 (N_1868,N_1035,N_1004);
and U1869 (N_1869,N_945,N_1437);
nand U1870 (N_1870,N_1222,N_1424);
and U1871 (N_1871,N_1227,N_986);
and U1872 (N_1872,N_1270,N_1421);
nand U1873 (N_1873,N_1273,N_967);
or U1874 (N_1874,N_944,N_831);
nand U1875 (N_1875,N_1121,N_1458);
nor U1876 (N_1876,N_1344,N_807);
nand U1877 (N_1877,N_750,N_921);
or U1878 (N_1878,N_1436,N_789);
nor U1879 (N_1879,N_1437,N_1185);
and U1880 (N_1880,N_862,N_815);
nor U1881 (N_1881,N_1198,N_1160);
nor U1882 (N_1882,N_763,N_950);
nor U1883 (N_1883,N_1182,N_899);
nand U1884 (N_1884,N_1421,N_764);
and U1885 (N_1885,N_1247,N_752);
nor U1886 (N_1886,N_962,N_1444);
or U1887 (N_1887,N_765,N_1060);
and U1888 (N_1888,N_1271,N_961);
and U1889 (N_1889,N_1024,N_1098);
or U1890 (N_1890,N_1220,N_1232);
nor U1891 (N_1891,N_831,N_799);
nor U1892 (N_1892,N_978,N_926);
nand U1893 (N_1893,N_1424,N_1042);
and U1894 (N_1894,N_1316,N_1485);
nor U1895 (N_1895,N_852,N_1120);
or U1896 (N_1896,N_892,N_1132);
and U1897 (N_1897,N_1006,N_828);
or U1898 (N_1898,N_1029,N_1292);
or U1899 (N_1899,N_1370,N_1381);
or U1900 (N_1900,N_1156,N_1340);
and U1901 (N_1901,N_1480,N_1408);
nand U1902 (N_1902,N_833,N_832);
or U1903 (N_1903,N_830,N_1086);
and U1904 (N_1904,N_1151,N_1083);
nand U1905 (N_1905,N_1347,N_1292);
nand U1906 (N_1906,N_1215,N_1460);
or U1907 (N_1907,N_1111,N_1309);
and U1908 (N_1908,N_1034,N_1409);
or U1909 (N_1909,N_870,N_1488);
nor U1910 (N_1910,N_1057,N_1103);
and U1911 (N_1911,N_1005,N_1160);
and U1912 (N_1912,N_849,N_909);
and U1913 (N_1913,N_849,N_843);
nor U1914 (N_1914,N_838,N_936);
nand U1915 (N_1915,N_752,N_1474);
and U1916 (N_1916,N_970,N_833);
nor U1917 (N_1917,N_1431,N_1301);
and U1918 (N_1918,N_1294,N_1207);
or U1919 (N_1919,N_1450,N_905);
nand U1920 (N_1920,N_1194,N_1481);
and U1921 (N_1921,N_1132,N_1152);
or U1922 (N_1922,N_1449,N_821);
and U1923 (N_1923,N_1300,N_1048);
nor U1924 (N_1924,N_1498,N_1390);
nand U1925 (N_1925,N_1074,N_1182);
nand U1926 (N_1926,N_1040,N_1431);
and U1927 (N_1927,N_1353,N_878);
nand U1928 (N_1928,N_1153,N_915);
nor U1929 (N_1929,N_960,N_1459);
and U1930 (N_1930,N_949,N_1286);
and U1931 (N_1931,N_1125,N_1129);
nand U1932 (N_1932,N_1398,N_923);
or U1933 (N_1933,N_1288,N_1320);
or U1934 (N_1934,N_1340,N_1453);
or U1935 (N_1935,N_1182,N_1471);
or U1936 (N_1936,N_1447,N_965);
nand U1937 (N_1937,N_1347,N_847);
nor U1938 (N_1938,N_768,N_1493);
or U1939 (N_1939,N_1117,N_1371);
or U1940 (N_1940,N_1034,N_999);
nand U1941 (N_1941,N_816,N_1085);
nand U1942 (N_1942,N_985,N_1342);
or U1943 (N_1943,N_1142,N_1290);
or U1944 (N_1944,N_929,N_1169);
or U1945 (N_1945,N_1369,N_1339);
nand U1946 (N_1946,N_1342,N_848);
or U1947 (N_1947,N_1128,N_1301);
or U1948 (N_1948,N_1029,N_1108);
nor U1949 (N_1949,N_1089,N_804);
nor U1950 (N_1950,N_1479,N_1166);
nor U1951 (N_1951,N_997,N_1316);
nor U1952 (N_1952,N_1019,N_1224);
and U1953 (N_1953,N_1076,N_1308);
or U1954 (N_1954,N_1243,N_1207);
or U1955 (N_1955,N_786,N_941);
and U1956 (N_1956,N_965,N_1193);
or U1957 (N_1957,N_1112,N_767);
nor U1958 (N_1958,N_1425,N_903);
or U1959 (N_1959,N_1334,N_887);
or U1960 (N_1960,N_1433,N_933);
nor U1961 (N_1961,N_852,N_1423);
nand U1962 (N_1962,N_1048,N_1041);
or U1963 (N_1963,N_967,N_1111);
nor U1964 (N_1964,N_972,N_1321);
and U1965 (N_1965,N_1051,N_1078);
or U1966 (N_1966,N_774,N_1234);
or U1967 (N_1967,N_1142,N_960);
and U1968 (N_1968,N_1209,N_1119);
and U1969 (N_1969,N_1266,N_758);
and U1970 (N_1970,N_1340,N_1394);
nor U1971 (N_1971,N_1071,N_1456);
nand U1972 (N_1972,N_1387,N_1460);
or U1973 (N_1973,N_841,N_1009);
nor U1974 (N_1974,N_807,N_1036);
or U1975 (N_1975,N_1442,N_953);
nor U1976 (N_1976,N_809,N_1388);
nor U1977 (N_1977,N_1014,N_1320);
or U1978 (N_1978,N_1262,N_976);
nand U1979 (N_1979,N_1424,N_898);
nand U1980 (N_1980,N_765,N_1251);
nor U1981 (N_1981,N_956,N_1445);
nor U1982 (N_1982,N_1485,N_836);
and U1983 (N_1983,N_836,N_1118);
nor U1984 (N_1984,N_814,N_1399);
nand U1985 (N_1985,N_1094,N_1057);
nand U1986 (N_1986,N_1245,N_1223);
nor U1987 (N_1987,N_1490,N_1448);
nor U1988 (N_1988,N_1053,N_1165);
nor U1989 (N_1989,N_972,N_1011);
nand U1990 (N_1990,N_1060,N_1359);
nand U1991 (N_1991,N_1368,N_777);
or U1992 (N_1992,N_1374,N_1130);
and U1993 (N_1993,N_893,N_826);
and U1994 (N_1994,N_961,N_1275);
nand U1995 (N_1995,N_1288,N_1433);
and U1996 (N_1996,N_805,N_814);
nor U1997 (N_1997,N_858,N_873);
nand U1998 (N_1998,N_1292,N_968);
nand U1999 (N_1999,N_789,N_910);
nor U2000 (N_2000,N_1126,N_813);
nand U2001 (N_2001,N_1066,N_1091);
or U2002 (N_2002,N_1164,N_854);
nand U2003 (N_2003,N_1057,N_1382);
or U2004 (N_2004,N_986,N_798);
or U2005 (N_2005,N_1138,N_1207);
and U2006 (N_2006,N_1381,N_881);
and U2007 (N_2007,N_1148,N_1338);
or U2008 (N_2008,N_1076,N_1205);
or U2009 (N_2009,N_1261,N_1230);
nor U2010 (N_2010,N_1012,N_876);
and U2011 (N_2011,N_1070,N_1198);
xnor U2012 (N_2012,N_1201,N_1447);
or U2013 (N_2013,N_902,N_1027);
nor U2014 (N_2014,N_1296,N_1468);
nor U2015 (N_2015,N_1069,N_1447);
nor U2016 (N_2016,N_816,N_1072);
xnor U2017 (N_2017,N_795,N_1165);
nand U2018 (N_2018,N_1025,N_999);
and U2019 (N_2019,N_847,N_1058);
and U2020 (N_2020,N_1309,N_856);
nand U2021 (N_2021,N_1018,N_1071);
nor U2022 (N_2022,N_1398,N_886);
and U2023 (N_2023,N_1146,N_1462);
and U2024 (N_2024,N_755,N_1495);
nand U2025 (N_2025,N_1475,N_846);
nor U2026 (N_2026,N_1283,N_1461);
nor U2027 (N_2027,N_1170,N_1001);
or U2028 (N_2028,N_947,N_817);
or U2029 (N_2029,N_1433,N_1055);
or U2030 (N_2030,N_1004,N_1342);
or U2031 (N_2031,N_1273,N_1470);
nand U2032 (N_2032,N_1002,N_1307);
or U2033 (N_2033,N_970,N_1402);
or U2034 (N_2034,N_802,N_811);
or U2035 (N_2035,N_1218,N_1489);
and U2036 (N_2036,N_1224,N_1134);
nor U2037 (N_2037,N_1104,N_1070);
xor U2038 (N_2038,N_1089,N_1251);
and U2039 (N_2039,N_1000,N_1265);
or U2040 (N_2040,N_1037,N_1383);
or U2041 (N_2041,N_885,N_1334);
nor U2042 (N_2042,N_1266,N_1247);
nor U2043 (N_2043,N_940,N_935);
or U2044 (N_2044,N_871,N_1320);
and U2045 (N_2045,N_1159,N_1450);
and U2046 (N_2046,N_1148,N_1235);
and U2047 (N_2047,N_914,N_878);
and U2048 (N_2048,N_1185,N_881);
and U2049 (N_2049,N_970,N_947);
or U2050 (N_2050,N_1100,N_1211);
or U2051 (N_2051,N_1250,N_1095);
nand U2052 (N_2052,N_1000,N_1418);
nor U2053 (N_2053,N_1212,N_1053);
and U2054 (N_2054,N_1034,N_1447);
nand U2055 (N_2055,N_1076,N_825);
and U2056 (N_2056,N_1029,N_1443);
or U2057 (N_2057,N_1477,N_1445);
or U2058 (N_2058,N_1074,N_1230);
nor U2059 (N_2059,N_1471,N_794);
nand U2060 (N_2060,N_1140,N_1177);
nor U2061 (N_2061,N_1118,N_1396);
or U2062 (N_2062,N_1046,N_1495);
nor U2063 (N_2063,N_1264,N_1245);
nor U2064 (N_2064,N_1291,N_750);
nand U2065 (N_2065,N_1347,N_1001);
nand U2066 (N_2066,N_983,N_1332);
nand U2067 (N_2067,N_1025,N_1253);
or U2068 (N_2068,N_756,N_1035);
or U2069 (N_2069,N_1174,N_1153);
or U2070 (N_2070,N_1105,N_1189);
nand U2071 (N_2071,N_815,N_1372);
xnor U2072 (N_2072,N_1338,N_1050);
nand U2073 (N_2073,N_836,N_1082);
nand U2074 (N_2074,N_1292,N_1380);
and U2075 (N_2075,N_1122,N_802);
nand U2076 (N_2076,N_818,N_1040);
nand U2077 (N_2077,N_1360,N_1126);
nand U2078 (N_2078,N_1140,N_1369);
and U2079 (N_2079,N_807,N_854);
xor U2080 (N_2080,N_1358,N_1160);
and U2081 (N_2081,N_868,N_818);
or U2082 (N_2082,N_1042,N_1046);
and U2083 (N_2083,N_1174,N_776);
xor U2084 (N_2084,N_1084,N_1494);
nand U2085 (N_2085,N_1102,N_771);
and U2086 (N_2086,N_901,N_1364);
nor U2087 (N_2087,N_775,N_1058);
or U2088 (N_2088,N_828,N_1223);
nand U2089 (N_2089,N_1243,N_1478);
and U2090 (N_2090,N_1288,N_1248);
nand U2091 (N_2091,N_837,N_923);
nor U2092 (N_2092,N_1425,N_762);
nor U2093 (N_2093,N_1134,N_756);
nand U2094 (N_2094,N_1078,N_1268);
nor U2095 (N_2095,N_1326,N_817);
or U2096 (N_2096,N_1309,N_1391);
and U2097 (N_2097,N_1132,N_1064);
or U2098 (N_2098,N_1283,N_944);
or U2099 (N_2099,N_962,N_1035);
or U2100 (N_2100,N_1045,N_788);
and U2101 (N_2101,N_1111,N_1280);
nor U2102 (N_2102,N_1192,N_991);
nor U2103 (N_2103,N_1279,N_876);
and U2104 (N_2104,N_830,N_1238);
nand U2105 (N_2105,N_875,N_1269);
and U2106 (N_2106,N_873,N_956);
xor U2107 (N_2107,N_1432,N_1311);
xor U2108 (N_2108,N_816,N_836);
nand U2109 (N_2109,N_1035,N_985);
and U2110 (N_2110,N_1283,N_1275);
or U2111 (N_2111,N_1041,N_826);
nand U2112 (N_2112,N_1187,N_1306);
or U2113 (N_2113,N_1214,N_1316);
nand U2114 (N_2114,N_840,N_1326);
xnor U2115 (N_2115,N_1046,N_1217);
and U2116 (N_2116,N_1317,N_1143);
nand U2117 (N_2117,N_783,N_1150);
nand U2118 (N_2118,N_1236,N_857);
or U2119 (N_2119,N_1419,N_1157);
nand U2120 (N_2120,N_1297,N_1304);
or U2121 (N_2121,N_874,N_847);
and U2122 (N_2122,N_1012,N_1019);
and U2123 (N_2123,N_937,N_1237);
nand U2124 (N_2124,N_1126,N_1380);
or U2125 (N_2125,N_1386,N_919);
or U2126 (N_2126,N_1219,N_1489);
nand U2127 (N_2127,N_856,N_910);
or U2128 (N_2128,N_879,N_941);
and U2129 (N_2129,N_815,N_1113);
or U2130 (N_2130,N_942,N_978);
nor U2131 (N_2131,N_1371,N_972);
and U2132 (N_2132,N_840,N_1433);
nor U2133 (N_2133,N_1064,N_864);
or U2134 (N_2134,N_834,N_1267);
or U2135 (N_2135,N_824,N_1041);
or U2136 (N_2136,N_1097,N_1451);
nor U2137 (N_2137,N_995,N_872);
nand U2138 (N_2138,N_1365,N_1141);
nand U2139 (N_2139,N_1261,N_1297);
nand U2140 (N_2140,N_1263,N_789);
and U2141 (N_2141,N_1071,N_1186);
and U2142 (N_2142,N_1004,N_750);
nor U2143 (N_2143,N_882,N_1034);
nor U2144 (N_2144,N_1110,N_1492);
and U2145 (N_2145,N_945,N_1122);
nor U2146 (N_2146,N_779,N_753);
or U2147 (N_2147,N_1018,N_805);
nand U2148 (N_2148,N_1105,N_1061);
and U2149 (N_2149,N_1473,N_777);
nor U2150 (N_2150,N_852,N_1325);
nand U2151 (N_2151,N_834,N_884);
nand U2152 (N_2152,N_1279,N_1202);
or U2153 (N_2153,N_1179,N_797);
and U2154 (N_2154,N_947,N_1395);
and U2155 (N_2155,N_1079,N_876);
and U2156 (N_2156,N_1152,N_1275);
nor U2157 (N_2157,N_952,N_1028);
and U2158 (N_2158,N_882,N_1149);
or U2159 (N_2159,N_1214,N_1332);
or U2160 (N_2160,N_1441,N_849);
or U2161 (N_2161,N_1167,N_1182);
nor U2162 (N_2162,N_889,N_1260);
nand U2163 (N_2163,N_1179,N_779);
nor U2164 (N_2164,N_994,N_1045);
and U2165 (N_2165,N_1408,N_1161);
and U2166 (N_2166,N_875,N_1426);
nor U2167 (N_2167,N_1458,N_1076);
and U2168 (N_2168,N_941,N_1093);
nand U2169 (N_2169,N_1372,N_887);
and U2170 (N_2170,N_912,N_1318);
or U2171 (N_2171,N_984,N_1422);
nand U2172 (N_2172,N_899,N_823);
nand U2173 (N_2173,N_1350,N_1278);
xor U2174 (N_2174,N_1475,N_1466);
and U2175 (N_2175,N_1443,N_954);
nand U2176 (N_2176,N_1321,N_1029);
and U2177 (N_2177,N_1170,N_955);
or U2178 (N_2178,N_1451,N_1350);
nand U2179 (N_2179,N_1033,N_1243);
or U2180 (N_2180,N_1193,N_878);
nor U2181 (N_2181,N_1040,N_972);
and U2182 (N_2182,N_1144,N_1325);
nor U2183 (N_2183,N_1004,N_1241);
nor U2184 (N_2184,N_1176,N_1080);
xor U2185 (N_2185,N_814,N_1127);
nand U2186 (N_2186,N_1229,N_1404);
nor U2187 (N_2187,N_1239,N_1332);
and U2188 (N_2188,N_1283,N_865);
nor U2189 (N_2189,N_1254,N_1285);
nor U2190 (N_2190,N_1179,N_1271);
or U2191 (N_2191,N_890,N_1428);
xor U2192 (N_2192,N_924,N_993);
xor U2193 (N_2193,N_943,N_962);
nor U2194 (N_2194,N_1134,N_831);
nor U2195 (N_2195,N_928,N_1215);
nand U2196 (N_2196,N_1015,N_979);
and U2197 (N_2197,N_1454,N_1312);
and U2198 (N_2198,N_1191,N_1231);
nor U2199 (N_2199,N_1244,N_993);
nand U2200 (N_2200,N_784,N_1452);
nand U2201 (N_2201,N_1028,N_1126);
nand U2202 (N_2202,N_785,N_1329);
nor U2203 (N_2203,N_1092,N_937);
nand U2204 (N_2204,N_1223,N_1088);
nor U2205 (N_2205,N_1081,N_1038);
nor U2206 (N_2206,N_1376,N_1020);
nor U2207 (N_2207,N_943,N_1114);
nor U2208 (N_2208,N_1103,N_980);
nor U2209 (N_2209,N_977,N_1180);
and U2210 (N_2210,N_1275,N_1201);
nor U2211 (N_2211,N_1471,N_1490);
nand U2212 (N_2212,N_1157,N_1306);
nor U2213 (N_2213,N_886,N_947);
nor U2214 (N_2214,N_830,N_1161);
nand U2215 (N_2215,N_754,N_1067);
or U2216 (N_2216,N_909,N_848);
and U2217 (N_2217,N_908,N_1441);
nor U2218 (N_2218,N_975,N_937);
nor U2219 (N_2219,N_1113,N_1007);
xnor U2220 (N_2220,N_803,N_909);
nand U2221 (N_2221,N_1002,N_758);
and U2222 (N_2222,N_1488,N_1337);
xnor U2223 (N_2223,N_1457,N_760);
or U2224 (N_2224,N_1099,N_953);
nand U2225 (N_2225,N_1328,N_791);
and U2226 (N_2226,N_1091,N_1013);
nor U2227 (N_2227,N_1121,N_808);
nand U2228 (N_2228,N_883,N_1158);
and U2229 (N_2229,N_973,N_974);
nor U2230 (N_2230,N_1298,N_878);
nand U2231 (N_2231,N_991,N_1045);
nand U2232 (N_2232,N_1257,N_1062);
and U2233 (N_2233,N_1205,N_932);
nand U2234 (N_2234,N_760,N_839);
and U2235 (N_2235,N_849,N_1197);
xor U2236 (N_2236,N_1343,N_1159);
and U2237 (N_2237,N_769,N_905);
or U2238 (N_2238,N_774,N_1437);
or U2239 (N_2239,N_874,N_1483);
or U2240 (N_2240,N_1238,N_828);
and U2241 (N_2241,N_798,N_1311);
nand U2242 (N_2242,N_944,N_899);
and U2243 (N_2243,N_1264,N_1133);
or U2244 (N_2244,N_876,N_1426);
or U2245 (N_2245,N_863,N_1429);
or U2246 (N_2246,N_846,N_1406);
nand U2247 (N_2247,N_801,N_1308);
and U2248 (N_2248,N_1204,N_1085);
nand U2249 (N_2249,N_826,N_1168);
nor U2250 (N_2250,N_2141,N_2095);
nor U2251 (N_2251,N_1878,N_2075);
nor U2252 (N_2252,N_1528,N_1960);
nor U2253 (N_2253,N_1891,N_1885);
nand U2254 (N_2254,N_1974,N_1625);
and U2255 (N_2255,N_1590,N_1916);
nor U2256 (N_2256,N_2093,N_1649);
xnor U2257 (N_2257,N_1808,N_1876);
and U2258 (N_2258,N_1520,N_2115);
and U2259 (N_2259,N_2008,N_2204);
nand U2260 (N_2260,N_1718,N_1970);
nor U2261 (N_2261,N_1881,N_2221);
and U2262 (N_2262,N_1711,N_2122);
or U2263 (N_2263,N_2230,N_1574);
nor U2264 (N_2264,N_2153,N_1848);
nor U2265 (N_2265,N_2031,N_1683);
or U2266 (N_2266,N_1860,N_1621);
and U2267 (N_2267,N_1775,N_1518);
and U2268 (N_2268,N_1912,N_2051);
nor U2269 (N_2269,N_1715,N_1644);
or U2270 (N_2270,N_1672,N_1598);
or U2271 (N_2271,N_1851,N_1819);
nand U2272 (N_2272,N_2155,N_2111);
or U2273 (N_2273,N_1604,N_1633);
nor U2274 (N_2274,N_1985,N_2034);
or U2275 (N_2275,N_1741,N_1664);
nand U2276 (N_2276,N_1943,N_1762);
xnor U2277 (N_2277,N_1716,N_1822);
and U2278 (N_2278,N_1654,N_2148);
nand U2279 (N_2279,N_1863,N_2218);
nor U2280 (N_2280,N_2028,N_2109);
or U2281 (N_2281,N_1911,N_1591);
and U2282 (N_2282,N_1721,N_2209);
nand U2283 (N_2283,N_1534,N_1723);
or U2284 (N_2284,N_1594,N_1700);
nor U2285 (N_2285,N_2129,N_1844);
nor U2286 (N_2286,N_1769,N_1545);
nand U2287 (N_2287,N_2108,N_1740);
xnor U2288 (N_2288,N_1837,N_1796);
nand U2289 (N_2289,N_2188,N_1557);
or U2290 (N_2290,N_2013,N_1934);
nand U2291 (N_2291,N_1880,N_1870);
nand U2292 (N_2292,N_1527,N_1952);
nor U2293 (N_2293,N_1969,N_1994);
or U2294 (N_2294,N_1615,N_1991);
nor U2295 (N_2295,N_2242,N_2102);
or U2296 (N_2296,N_1751,N_1903);
and U2297 (N_2297,N_1776,N_2107);
and U2298 (N_2298,N_1537,N_2037);
or U2299 (N_2299,N_1632,N_1733);
nand U2300 (N_2300,N_1575,N_2197);
nand U2301 (N_2301,N_1656,N_1768);
nand U2302 (N_2302,N_1995,N_2213);
and U2303 (N_2303,N_1951,N_2241);
and U2304 (N_2304,N_1993,N_2217);
or U2305 (N_2305,N_1523,N_1525);
nor U2306 (N_2306,N_2225,N_2152);
nor U2307 (N_2307,N_2061,N_1629);
nor U2308 (N_2308,N_2165,N_1948);
and U2309 (N_2309,N_1764,N_1918);
or U2310 (N_2310,N_1605,N_1685);
nor U2311 (N_2311,N_2098,N_1820);
and U2312 (N_2312,N_2189,N_2140);
and U2313 (N_2313,N_2058,N_1670);
nand U2314 (N_2314,N_1550,N_2077);
and U2315 (N_2315,N_1555,N_2143);
nand U2316 (N_2316,N_1688,N_1668);
and U2317 (N_2317,N_2159,N_1601);
nand U2318 (N_2318,N_1701,N_2121);
and U2319 (N_2319,N_2179,N_1779);
or U2320 (N_2320,N_1743,N_1818);
nand U2321 (N_2321,N_2081,N_1704);
or U2322 (N_2322,N_2002,N_1785);
nor U2323 (N_2323,N_1758,N_2125);
or U2324 (N_2324,N_1953,N_1850);
or U2325 (N_2325,N_2158,N_1753);
and U2326 (N_2326,N_1856,N_1674);
nor U2327 (N_2327,N_2135,N_1667);
nand U2328 (N_2328,N_1871,N_1532);
and U2329 (N_2329,N_2201,N_1802);
or U2330 (N_2330,N_1515,N_1907);
nand U2331 (N_2331,N_1650,N_2088);
or U2332 (N_2332,N_2147,N_1755);
and U2333 (N_2333,N_1967,N_2178);
nand U2334 (N_2334,N_1500,N_2096);
nand U2335 (N_2335,N_2222,N_1803);
nor U2336 (N_2336,N_1908,N_1724);
or U2337 (N_2337,N_1765,N_2145);
nor U2338 (N_2338,N_2030,N_1902);
or U2339 (N_2339,N_2101,N_2079);
and U2340 (N_2340,N_2022,N_2056);
nor U2341 (N_2341,N_2085,N_2047);
and U2342 (N_2342,N_2005,N_1921);
nor U2343 (N_2343,N_2127,N_1852);
nor U2344 (N_2344,N_2231,N_1507);
nand U2345 (N_2345,N_2083,N_2033);
or U2346 (N_2346,N_2214,N_1983);
or U2347 (N_2347,N_1562,N_1909);
nor U2348 (N_2348,N_1963,N_1989);
and U2349 (N_2349,N_1742,N_2200);
nand U2350 (N_2350,N_1813,N_1593);
nand U2351 (N_2351,N_1547,N_1634);
nand U2352 (N_2352,N_1987,N_1836);
or U2353 (N_2353,N_1945,N_1834);
and U2354 (N_2354,N_1928,N_1665);
or U2355 (N_2355,N_2130,N_2036);
and U2356 (N_2356,N_1693,N_1767);
nor U2357 (N_2357,N_2059,N_2212);
nand U2358 (N_2358,N_2011,N_1760);
nand U2359 (N_2359,N_2126,N_2180);
nand U2360 (N_2360,N_1869,N_1728);
or U2361 (N_2361,N_2166,N_1659);
nand U2362 (N_2362,N_1872,N_1867);
and U2363 (N_2363,N_1774,N_1595);
nand U2364 (N_2364,N_2190,N_2169);
nor U2365 (N_2365,N_1599,N_2114);
and U2366 (N_2366,N_1877,N_2012);
nand U2367 (N_2367,N_1807,N_1787);
xor U2368 (N_2368,N_2078,N_1554);
nor U2369 (N_2369,N_2208,N_1812);
and U2370 (N_2370,N_2228,N_2050);
nor U2371 (N_2371,N_1730,N_1978);
nand U2372 (N_2372,N_1933,N_1623);
and U2373 (N_2373,N_1592,N_2116);
nor U2374 (N_2374,N_2106,N_1564);
or U2375 (N_2375,N_1823,N_2039);
xor U2376 (N_2376,N_1973,N_1661);
nor U2377 (N_2377,N_1505,N_1901);
nand U2378 (N_2378,N_2049,N_2134);
nor U2379 (N_2379,N_1999,N_2035);
nand U2380 (N_2380,N_1846,N_1511);
nand U2381 (N_2381,N_2144,N_1955);
nand U2382 (N_2382,N_1568,N_1913);
and U2383 (N_2383,N_2067,N_1984);
nor U2384 (N_2384,N_2018,N_1900);
nor U2385 (N_2385,N_1620,N_1647);
nand U2386 (N_2386,N_1585,N_2154);
nand U2387 (N_2387,N_2001,N_1666);
or U2388 (N_2388,N_2157,N_1671);
and U2389 (N_2389,N_1795,N_1687);
nand U2390 (N_2390,N_1809,N_1965);
and U2391 (N_2391,N_2080,N_2173);
and U2392 (N_2392,N_2167,N_2027);
and U2393 (N_2393,N_1565,N_1731);
nand U2394 (N_2394,N_1607,N_2063);
and U2395 (N_2395,N_1893,N_1847);
nand U2396 (N_2396,N_1582,N_2046);
or U2397 (N_2397,N_1747,N_2128);
nor U2398 (N_2398,N_1990,N_1662);
nor U2399 (N_2399,N_1636,N_1986);
or U2400 (N_2400,N_1560,N_1502);
nor U2401 (N_2401,N_1691,N_1673);
xnor U2402 (N_2402,N_1556,N_2240);
nand U2403 (N_2403,N_2052,N_1979);
nor U2404 (N_2404,N_1517,N_1992);
nor U2405 (N_2405,N_1791,N_1864);
and U2406 (N_2406,N_1782,N_1503);
or U2407 (N_2407,N_1879,N_2124);
nand U2408 (N_2408,N_1680,N_1857);
nand U2409 (N_2409,N_1538,N_1608);
or U2410 (N_2410,N_1734,N_1602);
nand U2411 (N_2411,N_1966,N_1652);
or U2412 (N_2412,N_1522,N_1640);
xnor U2413 (N_2413,N_2211,N_1759);
and U2414 (N_2414,N_1941,N_1800);
or U2415 (N_2415,N_1577,N_2232);
nand U2416 (N_2416,N_1853,N_2216);
and U2417 (N_2417,N_2246,N_1618);
nor U2418 (N_2418,N_1663,N_2117);
nand U2419 (N_2419,N_1686,N_1890);
nand U2420 (N_2420,N_2105,N_2103);
nor U2421 (N_2421,N_2066,N_2084);
nand U2422 (N_2422,N_1542,N_1959);
and U2423 (N_2423,N_2175,N_2120);
nor U2424 (N_2424,N_1657,N_1587);
nand U2425 (N_2425,N_2029,N_1609);
nand U2426 (N_2426,N_2017,N_1946);
nand U2427 (N_2427,N_1729,N_1514);
or U2428 (N_2428,N_1790,N_2215);
nor U2429 (N_2429,N_2007,N_1923);
or U2430 (N_2430,N_1773,N_1610);
nand U2431 (N_2431,N_2239,N_1676);
and U2432 (N_2432,N_1914,N_2177);
nor U2433 (N_2433,N_1684,N_1692);
and U2434 (N_2434,N_1588,N_2119);
or U2435 (N_2435,N_2151,N_2186);
or U2436 (N_2436,N_1543,N_2170);
xor U2437 (N_2437,N_1763,N_1535);
or U2438 (N_2438,N_2090,N_1801);
nor U2439 (N_2439,N_2192,N_1551);
nand U2440 (N_2440,N_1613,N_2161);
and U2441 (N_2441,N_1971,N_2198);
or U2442 (N_2442,N_1540,N_2131);
nand U2443 (N_2443,N_1996,N_1982);
nor U2444 (N_2444,N_1799,N_1784);
nor U2445 (N_2445,N_1919,N_2025);
and U2446 (N_2446,N_1793,N_1957);
nor U2447 (N_2447,N_1641,N_1578);
nor U2448 (N_2448,N_1754,N_2042);
nor U2449 (N_2449,N_1709,N_1904);
and U2450 (N_2450,N_1868,N_1824);
and U2451 (N_2451,N_2237,N_1703);
nor U2452 (N_2452,N_1521,N_1873);
and U2453 (N_2453,N_1930,N_2062);
nand U2454 (N_2454,N_1761,N_1513);
nor U2455 (N_2455,N_2194,N_1717);
or U2456 (N_2456,N_1645,N_2207);
xnor U2457 (N_2457,N_1858,N_1544);
and U2458 (N_2458,N_2210,N_1886);
nand U2459 (N_2459,N_1713,N_1512);
and U2460 (N_2460,N_1744,N_1694);
nor U2461 (N_2461,N_1596,N_2026);
nor U2462 (N_2462,N_1727,N_1905);
and U2463 (N_2463,N_2181,N_2118);
or U2464 (N_2464,N_1707,N_1695);
and U2465 (N_2465,N_1771,N_2227);
and U2466 (N_2466,N_2057,N_1825);
and U2467 (N_2467,N_1936,N_1975);
nand U2468 (N_2468,N_2183,N_1888);
nor U2469 (N_2469,N_1842,N_1887);
nor U2470 (N_2470,N_1816,N_1726);
and U2471 (N_2471,N_2023,N_1745);
or U2472 (N_2472,N_1789,N_1706);
nand U2473 (N_2473,N_1679,N_1646);
nand U2474 (N_2474,N_1805,N_1536);
or U2475 (N_2475,N_1906,N_1998);
and U2476 (N_2476,N_2195,N_2138);
xnor U2477 (N_2477,N_1546,N_1533);
and U2478 (N_2478,N_2092,N_1506);
nor U2479 (N_2479,N_1897,N_2203);
or U2480 (N_2480,N_2146,N_2206);
nand U2481 (N_2481,N_1637,N_1712);
nor U2482 (N_2482,N_1814,N_2015);
or U2483 (N_2483,N_1746,N_2249);
or U2484 (N_2484,N_2089,N_1932);
or U2485 (N_2485,N_1792,N_1917);
nand U2486 (N_2486,N_1862,N_1770);
and U2487 (N_2487,N_1655,N_2168);
and U2488 (N_2488,N_1861,N_1682);
or U2489 (N_2489,N_2176,N_2219);
xnor U2490 (N_2490,N_1797,N_1708);
nor U2491 (N_2491,N_1579,N_1939);
and U2492 (N_2492,N_1570,N_1892);
or U2493 (N_2493,N_1839,N_1882);
and U2494 (N_2494,N_2236,N_2087);
or U2495 (N_2495,N_2224,N_1958);
nand U2496 (N_2496,N_1580,N_1931);
or U2497 (N_2497,N_2021,N_1735);
xor U2498 (N_2498,N_1828,N_1927);
nor U2499 (N_2499,N_1508,N_1584);
nand U2500 (N_2500,N_2226,N_1516);
nor U2501 (N_2501,N_1614,N_2032);
nand U2502 (N_2502,N_1635,N_2104);
nand U2503 (N_2503,N_2076,N_2038);
and U2504 (N_2504,N_1549,N_1899);
or U2505 (N_2505,N_1558,N_1981);
and U2506 (N_2506,N_2150,N_1722);
or U2507 (N_2507,N_1894,N_2040);
nand U2508 (N_2508,N_1843,N_1781);
nor U2509 (N_2509,N_1772,N_1531);
nand U2510 (N_2510,N_2185,N_1925);
nor U2511 (N_2511,N_1597,N_2229);
or U2512 (N_2512,N_1815,N_1949);
and U2513 (N_2513,N_1849,N_1576);
nor U2514 (N_2514,N_1783,N_1616);
nand U2515 (N_2515,N_2174,N_1895);
nor U2516 (N_2516,N_1651,N_2248);
or U2517 (N_2517,N_1719,N_1737);
nand U2518 (N_2518,N_1938,N_1915);
or U2519 (N_2519,N_1720,N_2070);
and U2520 (N_2520,N_1874,N_1643);
and U2521 (N_2521,N_1950,N_1530);
nor U2522 (N_2522,N_1896,N_1976);
nor U2523 (N_2523,N_1806,N_1732);
nor U2524 (N_2524,N_1826,N_2097);
or U2525 (N_2525,N_1541,N_2163);
and U2526 (N_2526,N_2060,N_1689);
nand U2527 (N_2527,N_2043,N_1788);
nand U2528 (N_2528,N_1980,N_2243);
and U2529 (N_2529,N_1922,N_2123);
nor U2530 (N_2530,N_1841,N_1710);
or U2531 (N_2531,N_2054,N_2072);
nand U2532 (N_2532,N_1942,N_2064);
and U2533 (N_2533,N_1855,N_2162);
or U2534 (N_2534,N_1572,N_1794);
or U2535 (N_2535,N_1875,N_1569);
nor U2536 (N_2536,N_1833,N_2205);
nor U2537 (N_2537,N_2069,N_1845);
nor U2538 (N_2538,N_1961,N_1660);
nand U2539 (N_2539,N_1866,N_1940);
nor U2540 (N_2540,N_2099,N_2041);
nor U2541 (N_2541,N_1519,N_1638);
and U2542 (N_2542,N_2136,N_1944);
or U2543 (N_2543,N_1639,N_1697);
and U2544 (N_2544,N_2048,N_1786);
nor U2545 (N_2545,N_1859,N_1750);
and U2546 (N_2546,N_1628,N_1924);
or U2547 (N_2547,N_1714,N_1977);
or U2548 (N_2548,N_1504,N_2202);
nor U2549 (N_2549,N_2187,N_2074);
nand U2550 (N_2550,N_1736,N_1810);
or U2551 (N_2551,N_2160,N_1889);
and U2552 (N_2552,N_2247,N_1830);
nor U2553 (N_2553,N_1619,N_1835);
nor U2554 (N_2554,N_2220,N_1937);
or U2555 (N_2555,N_1559,N_2010);
nand U2556 (N_2556,N_1630,N_1702);
nand U2557 (N_2557,N_1968,N_1964);
and U2558 (N_2558,N_1669,N_1956);
nor U2559 (N_2559,N_2000,N_1738);
nand U2560 (N_2560,N_2053,N_1972);
nand U2561 (N_2561,N_1696,N_1780);
and U2562 (N_2562,N_1827,N_1524);
or U2563 (N_2563,N_2244,N_2171);
nand U2564 (N_2564,N_1756,N_1501);
nand U2565 (N_2565,N_1606,N_2199);
nor U2566 (N_2566,N_2113,N_2142);
or U2567 (N_2567,N_1811,N_1725);
and U2568 (N_2568,N_2071,N_2014);
nand U2569 (N_2569,N_1757,N_1910);
and U2570 (N_2570,N_1690,N_2132);
or U2571 (N_2571,N_1529,N_1617);
or U2572 (N_2572,N_1539,N_1581);
or U2573 (N_2573,N_2100,N_2196);
or U2574 (N_2574,N_1571,N_2112);
nor U2575 (N_2575,N_1748,N_1988);
or U2576 (N_2576,N_1777,N_2020);
nor U2577 (N_2577,N_1698,N_1658);
or U2578 (N_2578,N_2193,N_1829);
nor U2579 (N_2579,N_1563,N_2235);
or U2580 (N_2580,N_2055,N_2139);
nand U2581 (N_2581,N_2223,N_1926);
and U2582 (N_2582,N_2044,N_2191);
nor U2583 (N_2583,N_1954,N_1962);
xor U2584 (N_2584,N_1935,N_2006);
nor U2585 (N_2585,N_1552,N_1648);
nor U2586 (N_2586,N_1947,N_2133);
nand U2587 (N_2587,N_2172,N_1612);
and U2588 (N_2588,N_1626,N_1553);
nand U2589 (N_2589,N_1883,N_1884);
or U2590 (N_2590,N_2182,N_1600);
and U2591 (N_2591,N_1675,N_1681);
nand U2592 (N_2592,N_2245,N_1817);
and U2593 (N_2593,N_1589,N_1510);
nand U2594 (N_2594,N_2073,N_1798);
nor U2595 (N_2595,N_2184,N_1705);
nor U2596 (N_2596,N_1627,N_1611);
or U2597 (N_2597,N_1622,N_2094);
and U2598 (N_2598,N_2164,N_1778);
nor U2599 (N_2599,N_1865,N_2238);
or U2600 (N_2600,N_2156,N_1561);
or U2601 (N_2601,N_1653,N_1898);
nand U2602 (N_2602,N_1699,N_2091);
or U2603 (N_2603,N_1624,N_1840);
nand U2604 (N_2604,N_2016,N_2045);
xor U2605 (N_2605,N_1821,N_1509);
and U2606 (N_2606,N_2065,N_1854);
or U2607 (N_2607,N_1526,N_1838);
or U2608 (N_2608,N_1749,N_1548);
nand U2609 (N_2609,N_1804,N_2019);
and U2610 (N_2610,N_2149,N_1631);
and U2611 (N_2611,N_1567,N_1831);
and U2612 (N_2612,N_2024,N_1678);
or U2613 (N_2613,N_2003,N_1642);
and U2614 (N_2614,N_2004,N_1583);
and U2615 (N_2615,N_2233,N_2082);
or U2616 (N_2616,N_1929,N_1677);
nand U2617 (N_2617,N_1573,N_1739);
nand U2618 (N_2618,N_1566,N_1832);
nand U2619 (N_2619,N_2086,N_1586);
and U2620 (N_2620,N_1752,N_2137);
xnor U2621 (N_2621,N_1920,N_2009);
and U2622 (N_2622,N_1766,N_1997);
nand U2623 (N_2623,N_1603,N_2110);
or U2624 (N_2624,N_2068,N_2234);
nand U2625 (N_2625,N_1896,N_1796);
and U2626 (N_2626,N_1731,N_1645);
nand U2627 (N_2627,N_1626,N_2029);
or U2628 (N_2628,N_2013,N_1605);
or U2629 (N_2629,N_2025,N_1979);
and U2630 (N_2630,N_1682,N_1873);
nand U2631 (N_2631,N_1533,N_1973);
nand U2632 (N_2632,N_1897,N_1719);
nand U2633 (N_2633,N_2092,N_2169);
and U2634 (N_2634,N_1583,N_1999);
or U2635 (N_2635,N_2014,N_1796);
or U2636 (N_2636,N_1595,N_2067);
or U2637 (N_2637,N_1685,N_1866);
or U2638 (N_2638,N_1925,N_2069);
nand U2639 (N_2639,N_1657,N_2159);
or U2640 (N_2640,N_1875,N_2074);
or U2641 (N_2641,N_1603,N_1614);
nand U2642 (N_2642,N_1845,N_1771);
or U2643 (N_2643,N_2210,N_2055);
nand U2644 (N_2644,N_1569,N_2164);
nor U2645 (N_2645,N_1732,N_1876);
nand U2646 (N_2646,N_1928,N_1888);
and U2647 (N_2647,N_2189,N_1794);
nand U2648 (N_2648,N_1693,N_1647);
nand U2649 (N_2649,N_2136,N_1635);
nand U2650 (N_2650,N_2211,N_1860);
nand U2651 (N_2651,N_2176,N_2009);
and U2652 (N_2652,N_1641,N_1862);
nand U2653 (N_2653,N_1857,N_1974);
and U2654 (N_2654,N_1850,N_1753);
or U2655 (N_2655,N_1856,N_1798);
nor U2656 (N_2656,N_1978,N_1678);
nor U2657 (N_2657,N_2142,N_2000);
xor U2658 (N_2658,N_2041,N_1574);
nand U2659 (N_2659,N_2014,N_1592);
nor U2660 (N_2660,N_2127,N_1887);
nor U2661 (N_2661,N_2200,N_1500);
nor U2662 (N_2662,N_2161,N_2074);
nand U2663 (N_2663,N_1707,N_2117);
nor U2664 (N_2664,N_1726,N_1917);
and U2665 (N_2665,N_2249,N_1722);
or U2666 (N_2666,N_1653,N_1850);
nand U2667 (N_2667,N_1723,N_2073);
nor U2668 (N_2668,N_2217,N_1610);
nor U2669 (N_2669,N_2078,N_2087);
nor U2670 (N_2670,N_1864,N_2116);
nor U2671 (N_2671,N_2127,N_1959);
nor U2672 (N_2672,N_2216,N_1522);
nand U2673 (N_2673,N_1879,N_1557);
and U2674 (N_2674,N_2148,N_1658);
nand U2675 (N_2675,N_2120,N_1758);
nor U2676 (N_2676,N_1552,N_1577);
or U2677 (N_2677,N_1800,N_2216);
or U2678 (N_2678,N_2084,N_1987);
or U2679 (N_2679,N_1620,N_2239);
and U2680 (N_2680,N_2085,N_2154);
xor U2681 (N_2681,N_1545,N_1949);
and U2682 (N_2682,N_1571,N_2248);
nand U2683 (N_2683,N_1644,N_1691);
nand U2684 (N_2684,N_1599,N_1942);
and U2685 (N_2685,N_1833,N_1830);
nor U2686 (N_2686,N_2034,N_2170);
and U2687 (N_2687,N_1788,N_1725);
and U2688 (N_2688,N_2050,N_2188);
or U2689 (N_2689,N_1563,N_2093);
nand U2690 (N_2690,N_1628,N_1906);
nor U2691 (N_2691,N_1578,N_2062);
nand U2692 (N_2692,N_2182,N_1769);
nand U2693 (N_2693,N_2162,N_2081);
or U2694 (N_2694,N_1907,N_1554);
and U2695 (N_2695,N_1601,N_1930);
nand U2696 (N_2696,N_1700,N_1533);
and U2697 (N_2697,N_1956,N_1906);
nand U2698 (N_2698,N_2220,N_1714);
and U2699 (N_2699,N_2210,N_2002);
nand U2700 (N_2700,N_1822,N_1877);
nor U2701 (N_2701,N_2151,N_2242);
or U2702 (N_2702,N_1841,N_2205);
nor U2703 (N_2703,N_2054,N_1980);
and U2704 (N_2704,N_1750,N_1598);
or U2705 (N_2705,N_1631,N_1666);
nand U2706 (N_2706,N_1822,N_1964);
xnor U2707 (N_2707,N_1544,N_1637);
nand U2708 (N_2708,N_1880,N_1563);
or U2709 (N_2709,N_2114,N_1903);
nand U2710 (N_2710,N_2089,N_1737);
nor U2711 (N_2711,N_2176,N_1595);
nor U2712 (N_2712,N_2056,N_2102);
nor U2713 (N_2713,N_2042,N_1600);
nand U2714 (N_2714,N_1878,N_1753);
or U2715 (N_2715,N_2194,N_1595);
and U2716 (N_2716,N_1666,N_1662);
xnor U2717 (N_2717,N_2001,N_2180);
and U2718 (N_2718,N_2138,N_1803);
nor U2719 (N_2719,N_2190,N_1921);
or U2720 (N_2720,N_1803,N_1918);
nor U2721 (N_2721,N_1750,N_1907);
nor U2722 (N_2722,N_2149,N_1596);
or U2723 (N_2723,N_2086,N_2051);
or U2724 (N_2724,N_1737,N_1965);
nor U2725 (N_2725,N_1873,N_2034);
or U2726 (N_2726,N_1993,N_1833);
nor U2727 (N_2727,N_1586,N_2057);
nor U2728 (N_2728,N_1797,N_1921);
nor U2729 (N_2729,N_2042,N_1982);
nor U2730 (N_2730,N_1840,N_1515);
nor U2731 (N_2731,N_1863,N_2234);
nand U2732 (N_2732,N_1546,N_1504);
and U2733 (N_2733,N_1924,N_1799);
xor U2734 (N_2734,N_1625,N_1946);
nand U2735 (N_2735,N_2208,N_1891);
and U2736 (N_2736,N_1850,N_2076);
nor U2737 (N_2737,N_2007,N_1554);
and U2738 (N_2738,N_1668,N_1670);
nand U2739 (N_2739,N_1701,N_2128);
or U2740 (N_2740,N_1944,N_2243);
nand U2741 (N_2741,N_2069,N_1669);
nand U2742 (N_2742,N_1577,N_1753);
nor U2743 (N_2743,N_1687,N_2163);
or U2744 (N_2744,N_2169,N_1852);
or U2745 (N_2745,N_2009,N_1584);
nand U2746 (N_2746,N_1773,N_2089);
nand U2747 (N_2747,N_2223,N_1878);
xnor U2748 (N_2748,N_1689,N_1984);
or U2749 (N_2749,N_1722,N_2123);
nand U2750 (N_2750,N_1719,N_2150);
nor U2751 (N_2751,N_2190,N_1869);
or U2752 (N_2752,N_1994,N_1764);
and U2753 (N_2753,N_1726,N_1745);
nor U2754 (N_2754,N_1724,N_1892);
or U2755 (N_2755,N_1510,N_1704);
and U2756 (N_2756,N_1954,N_2010);
or U2757 (N_2757,N_1824,N_2026);
nand U2758 (N_2758,N_2093,N_1517);
nor U2759 (N_2759,N_1865,N_2149);
and U2760 (N_2760,N_2056,N_1750);
or U2761 (N_2761,N_2095,N_1918);
or U2762 (N_2762,N_1900,N_1958);
nor U2763 (N_2763,N_1524,N_1800);
or U2764 (N_2764,N_1645,N_2153);
or U2765 (N_2765,N_1710,N_1529);
and U2766 (N_2766,N_1594,N_2222);
nor U2767 (N_2767,N_2163,N_1632);
nand U2768 (N_2768,N_1608,N_1990);
or U2769 (N_2769,N_2228,N_1540);
or U2770 (N_2770,N_2151,N_2024);
and U2771 (N_2771,N_1918,N_1745);
nor U2772 (N_2772,N_1725,N_2122);
nand U2773 (N_2773,N_1701,N_2115);
or U2774 (N_2774,N_1995,N_1922);
or U2775 (N_2775,N_1990,N_1808);
nor U2776 (N_2776,N_2196,N_1828);
nor U2777 (N_2777,N_2213,N_2148);
nor U2778 (N_2778,N_1957,N_2247);
nand U2779 (N_2779,N_1589,N_2031);
nor U2780 (N_2780,N_2175,N_2065);
or U2781 (N_2781,N_1919,N_1630);
nand U2782 (N_2782,N_2041,N_2148);
or U2783 (N_2783,N_1945,N_1754);
nand U2784 (N_2784,N_1959,N_2198);
or U2785 (N_2785,N_1622,N_1516);
and U2786 (N_2786,N_1572,N_1640);
nand U2787 (N_2787,N_2246,N_1909);
nor U2788 (N_2788,N_1543,N_1807);
nand U2789 (N_2789,N_1643,N_2202);
or U2790 (N_2790,N_1812,N_1950);
or U2791 (N_2791,N_1554,N_1561);
and U2792 (N_2792,N_1616,N_1812);
and U2793 (N_2793,N_1984,N_1839);
nor U2794 (N_2794,N_1547,N_2066);
or U2795 (N_2795,N_1546,N_2084);
or U2796 (N_2796,N_1941,N_1993);
nand U2797 (N_2797,N_1911,N_1864);
and U2798 (N_2798,N_1526,N_1607);
nand U2799 (N_2799,N_1700,N_1711);
or U2800 (N_2800,N_1757,N_1788);
nand U2801 (N_2801,N_2153,N_1557);
and U2802 (N_2802,N_1607,N_2110);
or U2803 (N_2803,N_1621,N_2067);
or U2804 (N_2804,N_2214,N_1952);
and U2805 (N_2805,N_1855,N_1896);
nand U2806 (N_2806,N_1766,N_1709);
nand U2807 (N_2807,N_1810,N_2165);
nand U2808 (N_2808,N_1626,N_1872);
or U2809 (N_2809,N_1910,N_2115);
nor U2810 (N_2810,N_1896,N_1930);
and U2811 (N_2811,N_2204,N_1808);
nor U2812 (N_2812,N_2183,N_1979);
xnor U2813 (N_2813,N_1546,N_2248);
and U2814 (N_2814,N_2006,N_2088);
nor U2815 (N_2815,N_2052,N_1879);
and U2816 (N_2816,N_2003,N_1952);
nand U2817 (N_2817,N_1793,N_2148);
or U2818 (N_2818,N_2245,N_2168);
or U2819 (N_2819,N_1802,N_1534);
nor U2820 (N_2820,N_2006,N_1575);
nor U2821 (N_2821,N_1861,N_2109);
and U2822 (N_2822,N_1525,N_2079);
nor U2823 (N_2823,N_1646,N_1647);
and U2824 (N_2824,N_1650,N_1626);
or U2825 (N_2825,N_1743,N_1529);
and U2826 (N_2826,N_1635,N_2141);
nor U2827 (N_2827,N_1997,N_2068);
and U2828 (N_2828,N_1733,N_1686);
and U2829 (N_2829,N_1774,N_2065);
nand U2830 (N_2830,N_1647,N_1745);
and U2831 (N_2831,N_2030,N_1795);
or U2832 (N_2832,N_1939,N_1713);
or U2833 (N_2833,N_1717,N_2081);
nor U2834 (N_2834,N_2138,N_1749);
nor U2835 (N_2835,N_1543,N_2017);
or U2836 (N_2836,N_1743,N_2168);
and U2837 (N_2837,N_2223,N_1691);
nand U2838 (N_2838,N_1677,N_1653);
nand U2839 (N_2839,N_1712,N_1549);
nor U2840 (N_2840,N_1501,N_2119);
or U2841 (N_2841,N_2092,N_1819);
nand U2842 (N_2842,N_1808,N_1557);
nand U2843 (N_2843,N_1532,N_1874);
or U2844 (N_2844,N_1823,N_2020);
or U2845 (N_2845,N_1718,N_1910);
nand U2846 (N_2846,N_1682,N_1538);
nand U2847 (N_2847,N_1699,N_1540);
or U2848 (N_2848,N_1889,N_2131);
and U2849 (N_2849,N_2229,N_1664);
nand U2850 (N_2850,N_1947,N_2129);
nor U2851 (N_2851,N_1911,N_1842);
nand U2852 (N_2852,N_1742,N_1839);
or U2853 (N_2853,N_1553,N_1776);
and U2854 (N_2854,N_1970,N_1931);
xor U2855 (N_2855,N_1873,N_2223);
or U2856 (N_2856,N_1991,N_1938);
and U2857 (N_2857,N_2172,N_1877);
nor U2858 (N_2858,N_2197,N_1724);
and U2859 (N_2859,N_1500,N_1699);
nand U2860 (N_2860,N_1677,N_1815);
or U2861 (N_2861,N_1646,N_1668);
and U2862 (N_2862,N_1771,N_2199);
nand U2863 (N_2863,N_2047,N_1730);
nand U2864 (N_2864,N_2101,N_1980);
and U2865 (N_2865,N_1994,N_1565);
nand U2866 (N_2866,N_1970,N_2053);
and U2867 (N_2867,N_1706,N_2160);
and U2868 (N_2868,N_1865,N_2135);
or U2869 (N_2869,N_1665,N_1841);
nand U2870 (N_2870,N_1823,N_2073);
and U2871 (N_2871,N_2129,N_1728);
nand U2872 (N_2872,N_1555,N_2222);
nor U2873 (N_2873,N_1601,N_1999);
xnor U2874 (N_2874,N_2059,N_1675);
nand U2875 (N_2875,N_1787,N_1785);
and U2876 (N_2876,N_2004,N_2029);
xor U2877 (N_2877,N_1822,N_2066);
nand U2878 (N_2878,N_1889,N_1970);
xor U2879 (N_2879,N_1946,N_2205);
or U2880 (N_2880,N_2165,N_1997);
nand U2881 (N_2881,N_1822,N_1827);
nor U2882 (N_2882,N_1833,N_1998);
or U2883 (N_2883,N_1774,N_2177);
and U2884 (N_2884,N_2212,N_2233);
nand U2885 (N_2885,N_1592,N_1756);
nand U2886 (N_2886,N_2152,N_1996);
xnor U2887 (N_2887,N_1863,N_1845);
or U2888 (N_2888,N_1733,N_1704);
and U2889 (N_2889,N_1979,N_1643);
or U2890 (N_2890,N_2148,N_2081);
and U2891 (N_2891,N_2241,N_2207);
and U2892 (N_2892,N_2180,N_1706);
nor U2893 (N_2893,N_2232,N_2223);
nand U2894 (N_2894,N_1587,N_1619);
or U2895 (N_2895,N_1510,N_1731);
nor U2896 (N_2896,N_2167,N_2243);
and U2897 (N_2897,N_1845,N_1795);
or U2898 (N_2898,N_2050,N_1597);
nand U2899 (N_2899,N_1904,N_1576);
and U2900 (N_2900,N_2015,N_1697);
or U2901 (N_2901,N_1781,N_2076);
and U2902 (N_2902,N_1665,N_1722);
and U2903 (N_2903,N_1746,N_2076);
and U2904 (N_2904,N_2047,N_1530);
or U2905 (N_2905,N_1767,N_1970);
nand U2906 (N_2906,N_2215,N_2222);
or U2907 (N_2907,N_1656,N_2200);
nor U2908 (N_2908,N_1770,N_1999);
nand U2909 (N_2909,N_2051,N_1579);
or U2910 (N_2910,N_2225,N_1512);
and U2911 (N_2911,N_1735,N_2007);
or U2912 (N_2912,N_1987,N_2065);
nor U2913 (N_2913,N_2026,N_2082);
nor U2914 (N_2914,N_1795,N_1547);
nand U2915 (N_2915,N_1903,N_1585);
nand U2916 (N_2916,N_2196,N_1693);
nor U2917 (N_2917,N_1508,N_2226);
nor U2918 (N_2918,N_1763,N_1671);
and U2919 (N_2919,N_2150,N_1820);
nand U2920 (N_2920,N_1881,N_2172);
or U2921 (N_2921,N_1736,N_1617);
nand U2922 (N_2922,N_2195,N_1673);
nand U2923 (N_2923,N_1681,N_2144);
or U2924 (N_2924,N_2010,N_1740);
and U2925 (N_2925,N_1758,N_2202);
nand U2926 (N_2926,N_1585,N_1536);
nand U2927 (N_2927,N_2208,N_1716);
or U2928 (N_2928,N_1597,N_1880);
nor U2929 (N_2929,N_1523,N_1975);
and U2930 (N_2930,N_2182,N_1508);
nor U2931 (N_2931,N_1719,N_2113);
nand U2932 (N_2932,N_2201,N_2181);
nor U2933 (N_2933,N_1842,N_2209);
xor U2934 (N_2934,N_1963,N_1659);
nor U2935 (N_2935,N_1915,N_1770);
and U2936 (N_2936,N_1594,N_2137);
and U2937 (N_2937,N_2080,N_2149);
nand U2938 (N_2938,N_1807,N_1984);
nand U2939 (N_2939,N_1646,N_1519);
or U2940 (N_2940,N_1946,N_1672);
or U2941 (N_2941,N_2084,N_1711);
nor U2942 (N_2942,N_1571,N_2151);
or U2943 (N_2943,N_1905,N_1978);
and U2944 (N_2944,N_1831,N_1843);
nand U2945 (N_2945,N_2059,N_1962);
or U2946 (N_2946,N_2177,N_2073);
or U2947 (N_2947,N_1537,N_2124);
nand U2948 (N_2948,N_2036,N_2026);
or U2949 (N_2949,N_2009,N_1719);
and U2950 (N_2950,N_1916,N_2022);
and U2951 (N_2951,N_2218,N_1940);
nor U2952 (N_2952,N_1800,N_1889);
and U2953 (N_2953,N_1769,N_1723);
or U2954 (N_2954,N_2058,N_1768);
nor U2955 (N_2955,N_1537,N_1737);
nand U2956 (N_2956,N_1621,N_1685);
nand U2957 (N_2957,N_1981,N_2096);
nand U2958 (N_2958,N_1994,N_2227);
and U2959 (N_2959,N_1802,N_2134);
and U2960 (N_2960,N_1692,N_1554);
nand U2961 (N_2961,N_2249,N_1613);
and U2962 (N_2962,N_2083,N_1852);
or U2963 (N_2963,N_1865,N_1509);
nor U2964 (N_2964,N_2202,N_2068);
nor U2965 (N_2965,N_1647,N_1981);
or U2966 (N_2966,N_1510,N_2173);
or U2967 (N_2967,N_1661,N_1642);
nand U2968 (N_2968,N_1502,N_1729);
nand U2969 (N_2969,N_1898,N_1864);
or U2970 (N_2970,N_2243,N_1842);
xor U2971 (N_2971,N_2088,N_2132);
or U2972 (N_2972,N_1525,N_2071);
nor U2973 (N_2973,N_1983,N_1670);
nor U2974 (N_2974,N_1891,N_1922);
nand U2975 (N_2975,N_1717,N_2218);
nor U2976 (N_2976,N_1674,N_1783);
nor U2977 (N_2977,N_1595,N_1989);
nand U2978 (N_2978,N_1564,N_1724);
and U2979 (N_2979,N_2206,N_1967);
nor U2980 (N_2980,N_1791,N_2054);
and U2981 (N_2981,N_1904,N_1656);
or U2982 (N_2982,N_1864,N_1690);
or U2983 (N_2983,N_1944,N_1941);
nand U2984 (N_2984,N_2034,N_2184);
and U2985 (N_2985,N_2045,N_1645);
nor U2986 (N_2986,N_1697,N_1559);
and U2987 (N_2987,N_2088,N_2015);
and U2988 (N_2988,N_1903,N_1851);
or U2989 (N_2989,N_2105,N_2137);
nor U2990 (N_2990,N_1556,N_1963);
xnor U2991 (N_2991,N_2064,N_1754);
or U2992 (N_2992,N_1940,N_1760);
nor U2993 (N_2993,N_2085,N_1531);
or U2994 (N_2994,N_1989,N_1611);
nor U2995 (N_2995,N_2245,N_1662);
nand U2996 (N_2996,N_1906,N_1574);
and U2997 (N_2997,N_1639,N_2039);
nand U2998 (N_2998,N_2004,N_2003);
or U2999 (N_2999,N_1620,N_2022);
or UO_0 (O_0,N_2801,N_2738);
and UO_1 (O_1,N_2818,N_2286);
nand UO_2 (O_2,N_2814,N_2646);
and UO_3 (O_3,N_2629,N_2493);
nor UO_4 (O_4,N_2513,N_2532);
or UO_5 (O_5,N_2984,N_2347);
or UO_6 (O_6,N_2500,N_2613);
nand UO_7 (O_7,N_2653,N_2705);
nand UO_8 (O_8,N_2729,N_2438);
or UO_9 (O_9,N_2279,N_2267);
nor UO_10 (O_10,N_2440,N_2293);
and UO_11 (O_11,N_2952,N_2254);
nand UO_12 (O_12,N_2737,N_2869);
nand UO_13 (O_13,N_2605,N_2755);
and UO_14 (O_14,N_2821,N_2315);
or UO_15 (O_15,N_2358,N_2551);
and UO_16 (O_16,N_2461,N_2402);
or UO_17 (O_17,N_2916,N_2921);
or UO_18 (O_18,N_2638,N_2652);
nand UO_19 (O_19,N_2678,N_2446);
xnor UO_20 (O_20,N_2807,N_2606);
nand UO_21 (O_21,N_2560,N_2320);
nand UO_22 (O_22,N_2787,N_2710);
nand UO_23 (O_23,N_2409,N_2651);
xor UO_24 (O_24,N_2890,N_2901);
nand UO_25 (O_25,N_2723,N_2791);
nand UO_26 (O_26,N_2876,N_2837);
nor UO_27 (O_27,N_2879,N_2258);
or UO_28 (O_28,N_2670,N_2745);
nand UO_29 (O_29,N_2387,N_2683);
or UO_30 (O_30,N_2999,N_2675);
nor UO_31 (O_31,N_2484,N_2593);
nand UO_32 (O_32,N_2400,N_2454);
nand UO_33 (O_33,N_2946,N_2371);
nor UO_34 (O_34,N_2832,N_2974);
or UO_35 (O_35,N_2873,N_2650);
nand UO_36 (O_36,N_2968,N_2452);
nand UO_37 (O_37,N_2739,N_2566);
nand UO_38 (O_38,N_2733,N_2702);
and UO_39 (O_39,N_2508,N_2528);
and UO_40 (O_40,N_2956,N_2514);
and UO_41 (O_41,N_2270,N_2852);
and UO_42 (O_42,N_2935,N_2337);
and UO_43 (O_43,N_2796,N_2326);
nor UO_44 (O_44,N_2340,N_2475);
nor UO_45 (O_45,N_2681,N_2268);
and UO_46 (O_46,N_2259,N_2995);
nor UO_47 (O_47,N_2778,N_2771);
and UO_48 (O_48,N_2991,N_2565);
nand UO_49 (O_49,N_2687,N_2630);
nand UO_50 (O_50,N_2838,N_2709);
and UO_51 (O_51,N_2856,N_2392);
nand UO_52 (O_52,N_2717,N_2281);
or UO_53 (O_53,N_2497,N_2919);
and UO_54 (O_54,N_2913,N_2352);
and UO_55 (O_55,N_2834,N_2718);
nor UO_56 (O_56,N_2987,N_2450);
or UO_57 (O_57,N_2313,N_2503);
nor UO_58 (O_58,N_2881,N_2250);
nand UO_59 (O_59,N_2458,N_2261);
or UO_60 (O_60,N_2877,N_2850);
and UO_61 (O_61,N_2769,N_2696);
nand UO_62 (O_62,N_2465,N_2257);
nand UO_63 (O_63,N_2793,N_2483);
nand UO_64 (O_64,N_2707,N_2616);
or UO_65 (O_65,N_2647,N_2361);
and UO_66 (O_66,N_2753,N_2994);
and UO_67 (O_67,N_2453,N_2682);
or UO_68 (O_68,N_2920,N_2841);
and UO_69 (O_69,N_2760,N_2990);
nand UO_70 (O_70,N_2624,N_2586);
or UO_71 (O_71,N_2393,N_2824);
nor UO_72 (O_72,N_2489,N_2482);
and UO_73 (O_73,N_2590,N_2357);
nor UO_74 (O_74,N_2859,N_2468);
or UO_75 (O_75,N_2563,N_2695);
or UO_76 (O_76,N_2985,N_2506);
and UO_77 (O_77,N_2810,N_2800);
nor UO_78 (O_78,N_2966,N_2923);
nor UO_79 (O_79,N_2549,N_2963);
or UO_80 (O_80,N_2958,N_2735);
nor UO_81 (O_81,N_2550,N_2910);
and UO_82 (O_82,N_2444,N_2721);
and UO_83 (O_83,N_2294,N_2636);
nand UO_84 (O_84,N_2331,N_2535);
or UO_85 (O_85,N_2997,N_2897);
and UO_86 (O_86,N_2734,N_2730);
nand UO_87 (O_87,N_2866,N_2385);
nor UO_88 (O_88,N_2295,N_2441);
nand UO_89 (O_89,N_2714,N_2662);
nand UO_90 (O_90,N_2900,N_2490);
or UO_91 (O_91,N_2547,N_2902);
or UO_92 (O_92,N_2266,N_2596);
or UO_93 (O_93,N_2562,N_2936);
nand UO_94 (O_94,N_2414,N_2372);
or UO_95 (O_95,N_2828,N_2580);
or UO_96 (O_96,N_2891,N_2359);
and UO_97 (O_97,N_2456,N_2983);
nand UO_98 (O_98,N_2494,N_2296);
and UO_99 (O_99,N_2280,N_2855);
or UO_100 (O_100,N_2311,N_2748);
nand UO_101 (O_101,N_2561,N_2543);
nand UO_102 (O_102,N_2469,N_2504);
and UO_103 (O_103,N_2459,N_2627);
or UO_104 (O_104,N_2542,N_2564);
nor UO_105 (O_105,N_2533,N_2511);
nor UO_106 (O_106,N_2338,N_2978);
nand UO_107 (O_107,N_2860,N_2570);
nor UO_108 (O_108,N_2263,N_2909);
and UO_109 (O_109,N_2269,N_2623);
nor UO_110 (O_110,N_2307,N_2608);
nor UO_111 (O_111,N_2977,N_2957);
or UO_112 (O_112,N_2439,N_2299);
or UO_113 (O_113,N_2728,N_2431);
nor UO_114 (O_114,N_2278,N_2525);
nor UO_115 (O_115,N_2747,N_2323);
nand UO_116 (O_116,N_2868,N_2430);
nand UO_117 (O_117,N_2880,N_2954);
nand UO_118 (O_118,N_2846,N_2480);
or UO_119 (O_119,N_2945,N_2667);
or UO_120 (O_120,N_2658,N_2727);
nor UO_121 (O_121,N_2905,N_2581);
nand UO_122 (O_122,N_2335,N_2448);
or UO_123 (O_123,N_2621,N_2965);
xor UO_124 (O_124,N_2819,N_2282);
nand UO_125 (O_125,N_2589,N_2460);
and UO_126 (O_126,N_2640,N_2848);
nor UO_127 (O_127,N_2287,N_2631);
or UO_128 (O_128,N_2744,N_2314);
nand UO_129 (O_129,N_2507,N_2327);
nor UO_130 (O_130,N_2384,N_2464);
and UO_131 (O_131,N_2726,N_2492);
nor UO_132 (O_132,N_2350,N_2654);
and UO_133 (O_133,N_2967,N_2376);
nand UO_134 (O_134,N_2959,N_2316);
nor UO_135 (O_135,N_2619,N_2644);
or UO_136 (O_136,N_2424,N_2896);
or UO_137 (O_137,N_2746,N_2688);
and UO_138 (O_138,N_2324,N_2708);
or UO_139 (O_139,N_2693,N_2411);
nand UO_140 (O_140,N_2799,N_2395);
nor UO_141 (O_141,N_2904,N_2495);
and UO_142 (O_142,N_2641,N_2970);
nand UO_143 (O_143,N_2285,N_2540);
or UO_144 (O_144,N_2568,N_2501);
and UO_145 (O_145,N_2782,N_2379);
and UO_146 (O_146,N_2784,N_2704);
xor UO_147 (O_147,N_2764,N_2382);
and UO_148 (O_148,N_2322,N_2413);
and UO_149 (O_149,N_2779,N_2649);
or UO_150 (O_150,N_2854,N_2304);
nand UO_151 (O_151,N_2617,N_2813);
or UO_152 (O_152,N_2825,N_2642);
and UO_153 (O_153,N_2255,N_2584);
nand UO_154 (O_154,N_2447,N_2757);
nor UO_155 (O_155,N_2585,N_2569);
and UO_156 (O_156,N_2491,N_2434);
nor UO_157 (O_157,N_2812,N_2817);
or UO_158 (O_158,N_2772,N_2396);
nand UO_159 (O_159,N_2334,N_2740);
nor UO_160 (O_160,N_2895,N_2575);
and UO_161 (O_161,N_2686,N_2445);
and UO_162 (O_162,N_2763,N_2419);
nand UO_163 (O_163,N_2872,N_2657);
and UO_164 (O_164,N_2499,N_2843);
or UO_165 (O_165,N_2516,N_2684);
or UO_166 (O_166,N_2582,N_2428);
or UO_167 (O_167,N_2878,N_2993);
nor UO_168 (O_168,N_2284,N_2732);
nand UO_169 (O_169,N_2317,N_2773);
and UO_170 (O_170,N_2407,N_2422);
nor UO_171 (O_171,N_2949,N_2780);
and UO_172 (O_172,N_2442,N_2583);
nor UO_173 (O_173,N_2515,N_2816);
or UO_174 (O_174,N_2842,N_2524);
or UO_175 (O_175,N_2716,N_2505);
and UO_176 (O_176,N_2743,N_2853);
and UO_177 (O_177,N_2998,N_2463);
and UO_178 (O_178,N_2473,N_2665);
or UO_179 (O_179,N_2759,N_2598);
nand UO_180 (O_180,N_2942,N_2345);
and UO_181 (O_181,N_2425,N_2899);
nand UO_182 (O_182,N_2436,N_2969);
nand UO_183 (O_183,N_2415,N_2830);
or UO_184 (O_184,N_2941,N_2634);
nand UO_185 (O_185,N_2668,N_2477);
nand UO_186 (O_186,N_2711,N_2487);
nor UO_187 (O_187,N_2697,N_2292);
or UO_188 (O_188,N_2626,N_2907);
and UO_189 (O_189,N_2509,N_2786);
or UO_190 (O_190,N_2822,N_2604);
or UO_191 (O_191,N_2378,N_2301);
or UO_192 (O_192,N_2973,N_2986);
nor UO_193 (O_193,N_2291,N_2521);
or UO_194 (O_194,N_2609,N_2903);
or UO_195 (O_195,N_2297,N_2979);
nand UO_196 (O_196,N_2761,N_2768);
and UO_197 (O_197,N_2546,N_2756);
or UO_198 (O_198,N_2610,N_2394);
and UO_199 (O_199,N_2595,N_2510);
nand UO_200 (O_200,N_2433,N_2274);
nor UO_201 (O_201,N_2368,N_2374);
nand UO_202 (O_202,N_2847,N_2518);
nand UO_203 (O_203,N_2474,N_2861);
and UO_204 (O_204,N_2363,N_2576);
nand UO_205 (O_205,N_2981,N_2423);
or UO_206 (O_206,N_2988,N_2364);
and UO_207 (O_207,N_2399,N_2618);
nand UO_208 (O_208,N_2312,N_2591);
nand UO_209 (O_209,N_2870,N_2758);
nor UO_210 (O_210,N_2719,N_2845);
nor UO_211 (O_211,N_2309,N_2397);
nand UO_212 (O_212,N_2770,N_2792);
nand UO_213 (O_213,N_2289,N_2777);
and UO_214 (O_214,N_2893,N_2804);
or UO_215 (O_215,N_2427,N_2488);
and UO_216 (O_216,N_2332,N_2554);
nor UO_217 (O_217,N_2391,N_2275);
and UO_218 (O_218,N_2599,N_2715);
or UO_219 (O_219,N_2362,N_2950);
and UO_220 (O_220,N_2925,N_2674);
and UO_221 (O_221,N_2579,N_2602);
and UO_222 (O_222,N_2673,N_2265);
or UO_223 (O_223,N_2271,N_2625);
nor UO_224 (O_224,N_2451,N_2534);
and UO_225 (O_225,N_2470,N_2989);
or UO_226 (O_226,N_2346,N_2481);
nand UO_227 (O_227,N_2926,N_2672);
or UO_228 (O_228,N_2976,N_2406);
nand UO_229 (O_229,N_2558,N_2953);
and UO_230 (O_230,N_2614,N_2351);
and UO_231 (O_231,N_2961,N_2948);
nor UO_232 (O_232,N_2403,N_2588);
nor UO_233 (O_233,N_2689,N_2836);
nand UO_234 (O_234,N_2794,N_2632);
and UO_235 (O_235,N_2835,N_2685);
and UO_236 (O_236,N_2522,N_2661);
or UO_237 (O_237,N_2706,N_2930);
and UO_238 (O_238,N_2964,N_2938);
nor UO_239 (O_239,N_2887,N_2932);
nor UO_240 (O_240,N_2405,N_2908);
and UO_241 (O_241,N_2260,N_2703);
or UO_242 (O_242,N_2611,N_2587);
xnor UO_243 (O_243,N_2655,N_2389);
nor UO_244 (O_244,N_2871,N_2353);
or UO_245 (O_245,N_2694,N_2472);
nand UO_246 (O_246,N_2556,N_2573);
nor UO_247 (O_247,N_2398,N_2545);
nor UO_248 (O_248,N_2574,N_2656);
nand UO_249 (O_249,N_2290,N_2882);
or UO_250 (O_250,N_2677,N_2857);
nand UO_251 (O_251,N_2833,N_2552);
nand UO_252 (O_252,N_2512,N_2302);
nand UO_253 (O_253,N_2972,N_2417);
or UO_254 (O_254,N_2319,N_2955);
xnor UO_255 (O_255,N_2633,N_2937);
or UO_256 (O_256,N_2940,N_2671);
nand UO_257 (O_257,N_2333,N_2951);
or UO_258 (O_258,N_2788,N_2874);
or UO_259 (O_259,N_2840,N_2762);
nand UO_260 (O_260,N_2305,N_2783);
or UO_261 (O_261,N_2479,N_2698);
nand UO_262 (O_262,N_2971,N_2601);
nor UO_263 (O_263,N_2865,N_2690);
or UO_264 (O_264,N_2622,N_2437);
nor UO_265 (O_265,N_2498,N_2536);
or UO_266 (O_266,N_2578,N_2555);
or UO_267 (O_267,N_2523,N_2502);
nor UO_268 (O_268,N_2712,N_2380);
nor UO_269 (O_269,N_2262,N_2669);
nor UO_270 (O_270,N_2918,N_2615);
or UO_271 (O_271,N_2659,N_2750);
nand UO_272 (O_272,N_2858,N_2252);
nor UO_273 (O_273,N_2342,N_2639);
and UO_274 (O_274,N_2527,N_2412);
nor UO_275 (O_275,N_2917,N_2520);
nand UO_276 (O_276,N_2366,N_2699);
or UO_277 (O_277,N_2478,N_2823);
or UO_278 (O_278,N_2775,N_2336);
nand UO_279 (O_279,N_2892,N_2864);
and UO_280 (O_280,N_2449,N_2517);
and UO_281 (O_281,N_2785,N_2914);
nor UO_282 (O_282,N_2929,N_2467);
or UO_283 (O_283,N_2386,N_2421);
xor UO_284 (O_284,N_2912,N_2645);
nand UO_285 (O_285,N_2666,N_2557);
nor UO_286 (O_286,N_2339,N_2924);
or UO_287 (O_287,N_2637,N_2519);
or UO_288 (O_288,N_2251,N_2603);
or UO_289 (O_289,N_2466,N_2975);
or UO_290 (O_290,N_2808,N_2643);
or UO_291 (O_291,N_2344,N_2306);
nor UO_292 (O_292,N_2894,N_2538);
or UO_293 (O_293,N_2310,N_2915);
and UO_294 (O_294,N_2594,N_2476);
or UO_295 (O_295,N_2471,N_2933);
nand UO_296 (O_296,N_2485,N_2883);
nand UO_297 (O_297,N_2328,N_2820);
or UO_298 (O_298,N_2612,N_2898);
nand UO_299 (O_299,N_2321,N_2798);
or UO_300 (O_300,N_2815,N_2544);
nor UO_301 (O_301,N_2329,N_2432);
and UO_302 (O_302,N_2531,N_2537);
or UO_303 (O_303,N_2947,N_2369);
nand UO_304 (O_304,N_2373,N_2607);
and UO_305 (O_305,N_2802,N_2939);
nand UO_306 (O_306,N_2889,N_2660);
nand UO_307 (O_307,N_2435,N_2867);
nor UO_308 (O_308,N_2789,N_2680);
nand UO_309 (O_309,N_2298,N_2455);
nand UO_310 (O_310,N_2911,N_2700);
nor UO_311 (O_311,N_2803,N_2388);
or UO_312 (O_312,N_2960,N_2303);
nor UO_313 (O_313,N_2356,N_2805);
and UO_314 (O_314,N_2713,N_2962);
or UO_315 (O_315,N_2343,N_2648);
nand UO_316 (O_316,N_2367,N_2741);
nand UO_317 (O_317,N_2420,N_2539);
and UO_318 (O_318,N_2736,N_2766);
nand UO_319 (O_319,N_2486,N_2992);
nand UO_320 (O_320,N_2462,N_2982);
nor UO_321 (O_321,N_2724,N_2375);
or UO_322 (O_322,N_2354,N_2811);
or UO_323 (O_323,N_2355,N_2370);
nor UO_324 (O_324,N_2457,N_2390);
and UO_325 (O_325,N_2752,N_2862);
nand UO_326 (O_326,N_2429,N_2572);
nand UO_327 (O_327,N_2559,N_2264);
nor UO_328 (O_328,N_2722,N_2571);
and UO_329 (O_329,N_2751,N_2360);
nor UO_330 (O_330,N_2365,N_2906);
and UO_331 (O_331,N_2283,N_2526);
nand UO_332 (O_332,N_2426,N_2664);
nand UO_333 (O_333,N_2790,N_2851);
nand UO_334 (O_334,N_2404,N_2288);
nand UO_335 (O_335,N_2996,N_2774);
nand UO_336 (O_336,N_2795,N_2797);
nand UO_337 (O_337,N_2875,N_2826);
nand UO_338 (O_338,N_2300,N_2831);
or UO_339 (O_339,N_2806,N_2496);
nand UO_340 (O_340,N_2691,N_2341);
or UO_341 (O_341,N_2827,N_2943);
or UO_342 (O_342,N_2928,N_2888);
and UO_343 (O_343,N_2885,N_2980);
nand UO_344 (O_344,N_2749,N_2325);
and UO_345 (O_345,N_2731,N_2276);
and UO_346 (O_346,N_2809,N_2754);
nand UO_347 (O_347,N_2541,N_2577);
nor UO_348 (O_348,N_2253,N_2720);
nand UO_349 (O_349,N_2272,N_2922);
nand UO_350 (O_350,N_2635,N_2273);
nor UO_351 (O_351,N_2725,N_2676);
nor UO_352 (O_352,N_2600,N_2844);
and UO_353 (O_353,N_2530,N_2592);
nand UO_354 (O_354,N_2349,N_2628);
nor UO_355 (O_355,N_2701,N_2548);
or UO_356 (O_356,N_2256,N_2401);
nor UO_357 (O_357,N_2884,N_2863);
and UO_358 (O_358,N_2781,N_2348);
nand UO_359 (O_359,N_2829,N_2663);
or UO_360 (O_360,N_2765,N_2277);
or UO_361 (O_361,N_2839,N_2553);
and UO_362 (O_362,N_2408,N_2377);
and UO_363 (O_363,N_2330,N_2381);
or UO_364 (O_364,N_2934,N_2849);
or UO_365 (O_365,N_2443,N_2620);
nor UO_366 (O_366,N_2567,N_2308);
nand UO_367 (O_367,N_2944,N_2529);
nand UO_368 (O_368,N_2931,N_2767);
nor UO_369 (O_369,N_2886,N_2927);
and UO_370 (O_370,N_2776,N_2742);
nor UO_371 (O_371,N_2410,N_2692);
or UO_372 (O_372,N_2416,N_2318);
nand UO_373 (O_373,N_2383,N_2418);
nor UO_374 (O_374,N_2597,N_2679);
and UO_375 (O_375,N_2690,N_2385);
and UO_376 (O_376,N_2360,N_2260);
and UO_377 (O_377,N_2728,N_2262);
nand UO_378 (O_378,N_2929,N_2804);
nand UO_379 (O_379,N_2938,N_2707);
nand UO_380 (O_380,N_2349,N_2769);
nor UO_381 (O_381,N_2802,N_2600);
and UO_382 (O_382,N_2258,N_2922);
nor UO_383 (O_383,N_2292,N_2706);
nor UO_384 (O_384,N_2988,N_2765);
or UO_385 (O_385,N_2429,N_2534);
or UO_386 (O_386,N_2341,N_2688);
or UO_387 (O_387,N_2965,N_2488);
nand UO_388 (O_388,N_2629,N_2657);
nor UO_389 (O_389,N_2551,N_2755);
or UO_390 (O_390,N_2584,N_2368);
xor UO_391 (O_391,N_2648,N_2916);
or UO_392 (O_392,N_2812,N_2840);
or UO_393 (O_393,N_2653,N_2335);
nor UO_394 (O_394,N_2473,N_2909);
and UO_395 (O_395,N_2714,N_2726);
nand UO_396 (O_396,N_2288,N_2484);
and UO_397 (O_397,N_2713,N_2691);
nor UO_398 (O_398,N_2287,N_2671);
and UO_399 (O_399,N_2989,N_2841);
nand UO_400 (O_400,N_2864,N_2346);
nand UO_401 (O_401,N_2476,N_2471);
or UO_402 (O_402,N_2890,N_2864);
or UO_403 (O_403,N_2364,N_2953);
or UO_404 (O_404,N_2823,N_2675);
and UO_405 (O_405,N_2634,N_2486);
and UO_406 (O_406,N_2913,N_2624);
nor UO_407 (O_407,N_2421,N_2677);
or UO_408 (O_408,N_2885,N_2636);
or UO_409 (O_409,N_2373,N_2897);
nor UO_410 (O_410,N_2548,N_2852);
or UO_411 (O_411,N_2436,N_2649);
and UO_412 (O_412,N_2473,N_2779);
nor UO_413 (O_413,N_2398,N_2395);
and UO_414 (O_414,N_2708,N_2990);
and UO_415 (O_415,N_2318,N_2915);
and UO_416 (O_416,N_2439,N_2513);
or UO_417 (O_417,N_2683,N_2456);
nor UO_418 (O_418,N_2425,N_2572);
or UO_419 (O_419,N_2370,N_2834);
nor UO_420 (O_420,N_2727,N_2269);
nand UO_421 (O_421,N_2844,N_2949);
and UO_422 (O_422,N_2377,N_2343);
nor UO_423 (O_423,N_2769,N_2387);
xnor UO_424 (O_424,N_2256,N_2957);
or UO_425 (O_425,N_2476,N_2752);
nand UO_426 (O_426,N_2685,N_2628);
or UO_427 (O_427,N_2753,N_2378);
and UO_428 (O_428,N_2851,N_2267);
nand UO_429 (O_429,N_2638,N_2735);
or UO_430 (O_430,N_2988,N_2645);
nand UO_431 (O_431,N_2769,N_2904);
nand UO_432 (O_432,N_2857,N_2830);
nor UO_433 (O_433,N_2898,N_2599);
and UO_434 (O_434,N_2519,N_2983);
nor UO_435 (O_435,N_2316,N_2443);
or UO_436 (O_436,N_2587,N_2987);
and UO_437 (O_437,N_2816,N_2850);
nand UO_438 (O_438,N_2617,N_2555);
and UO_439 (O_439,N_2987,N_2767);
nand UO_440 (O_440,N_2957,N_2407);
and UO_441 (O_441,N_2829,N_2912);
nand UO_442 (O_442,N_2299,N_2490);
or UO_443 (O_443,N_2903,N_2497);
and UO_444 (O_444,N_2689,N_2568);
or UO_445 (O_445,N_2524,N_2858);
nor UO_446 (O_446,N_2782,N_2897);
nand UO_447 (O_447,N_2365,N_2976);
and UO_448 (O_448,N_2882,N_2898);
nand UO_449 (O_449,N_2492,N_2403);
nand UO_450 (O_450,N_2275,N_2685);
nand UO_451 (O_451,N_2620,N_2377);
nor UO_452 (O_452,N_2509,N_2929);
nor UO_453 (O_453,N_2467,N_2422);
nor UO_454 (O_454,N_2338,N_2928);
and UO_455 (O_455,N_2477,N_2590);
and UO_456 (O_456,N_2872,N_2581);
and UO_457 (O_457,N_2908,N_2476);
and UO_458 (O_458,N_2294,N_2621);
xor UO_459 (O_459,N_2640,N_2328);
nor UO_460 (O_460,N_2436,N_2809);
nor UO_461 (O_461,N_2323,N_2879);
and UO_462 (O_462,N_2363,N_2984);
nor UO_463 (O_463,N_2910,N_2931);
nor UO_464 (O_464,N_2364,N_2831);
or UO_465 (O_465,N_2801,N_2789);
nor UO_466 (O_466,N_2953,N_2471);
and UO_467 (O_467,N_2720,N_2310);
nand UO_468 (O_468,N_2961,N_2547);
or UO_469 (O_469,N_2457,N_2318);
and UO_470 (O_470,N_2616,N_2272);
nand UO_471 (O_471,N_2492,N_2676);
nand UO_472 (O_472,N_2902,N_2379);
or UO_473 (O_473,N_2375,N_2641);
nor UO_474 (O_474,N_2931,N_2343);
nor UO_475 (O_475,N_2905,N_2962);
nand UO_476 (O_476,N_2677,N_2353);
and UO_477 (O_477,N_2529,N_2384);
nor UO_478 (O_478,N_2615,N_2644);
xnor UO_479 (O_479,N_2563,N_2705);
and UO_480 (O_480,N_2453,N_2340);
nor UO_481 (O_481,N_2868,N_2735);
or UO_482 (O_482,N_2701,N_2471);
nor UO_483 (O_483,N_2674,N_2436);
and UO_484 (O_484,N_2585,N_2416);
or UO_485 (O_485,N_2879,N_2790);
or UO_486 (O_486,N_2351,N_2944);
nand UO_487 (O_487,N_2745,N_2506);
or UO_488 (O_488,N_2360,N_2872);
xor UO_489 (O_489,N_2726,N_2443);
nand UO_490 (O_490,N_2597,N_2636);
or UO_491 (O_491,N_2632,N_2253);
and UO_492 (O_492,N_2665,N_2319);
and UO_493 (O_493,N_2272,N_2872);
nand UO_494 (O_494,N_2551,N_2387);
and UO_495 (O_495,N_2593,N_2263);
or UO_496 (O_496,N_2653,N_2689);
xor UO_497 (O_497,N_2579,N_2293);
nand UO_498 (O_498,N_2749,N_2466);
nand UO_499 (O_499,N_2334,N_2961);
endmodule