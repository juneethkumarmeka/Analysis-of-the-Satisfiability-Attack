module basic_2500_25000_3000_4_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18760,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18985,N_18986,N_18987,N_18988,N_18989,N_18991,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19203,N_19204,N_19205,N_19207,N_19208,N_19209,N_19210,N_19211,N_19213,N_19214,N_19215,N_19216,N_19217,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19344,N_19345,N_19346,N_19347,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19624,N_19625,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19651,N_19652,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19813,N_19814,N_19815,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19921,N_19922,N_19923,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20003,N_20004,N_20005,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20023,N_20024,N_20025,N_20026,N_20027,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20118,N_20119,N_20120,N_20121,N_20122,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20131,N_20132,N_20133,N_20134,N_20135,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20482,N_20483,N_20484,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20587,N_20588,N_20589,N_20591,N_20592,N_20593,N_20594,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20957,N_20958,N_20959,N_20961,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21129,N_21130,N_21131,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21155,N_21157,N_21158,N_21159,N_21160,N_21161,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21309,N_21310,N_21311,N_21312,N_21313,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21615,N_21616,N_21617,N_21618,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21712,N_21713,N_21714,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21817,N_21818,N_21819,N_21820,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21879,N_21881,N_21882,N_21884,N_21885,N_21886,N_21887,N_21888,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22254,N_22255,N_22256,N_22257,N_22258,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22268,N_22269,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22307,N_22308,N_22310,N_22311,N_22312,N_22314,N_22315,N_22317,N_22318,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23628,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23658,N_23659,N_23660,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24165,N_24167,N_24168,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24417,N_24418,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24539,N_24540,N_24541,N_24542,N_24544,N_24545,N_24546,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24708,N_24709,N_24710,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24865,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_51,In_1705);
nor U1 (N_1,In_1886,In_762);
nor U2 (N_2,In_2291,In_1);
nand U3 (N_3,In_1463,In_895);
and U4 (N_4,In_512,In_2095);
or U5 (N_5,In_885,In_1655);
or U6 (N_6,In_2390,In_2104);
or U7 (N_7,In_1126,In_1958);
or U8 (N_8,In_296,In_476);
xor U9 (N_9,In_1283,In_938);
and U10 (N_10,In_1119,In_2468);
and U11 (N_11,In_2364,In_289);
and U12 (N_12,In_2230,In_708);
or U13 (N_13,In_1406,In_1263);
and U14 (N_14,In_2347,In_1538);
nand U15 (N_15,In_112,In_1598);
xnor U16 (N_16,In_1134,In_893);
nor U17 (N_17,In_385,In_1060);
nor U18 (N_18,In_341,In_76);
nand U19 (N_19,In_1569,In_1218);
nand U20 (N_20,In_625,In_688);
xnor U21 (N_21,In_1585,In_1334);
nand U22 (N_22,In_2422,In_1017);
and U23 (N_23,In_1164,In_851);
nor U24 (N_24,In_1482,In_1480);
nand U25 (N_25,In_1107,In_1782);
nand U26 (N_26,In_546,In_751);
xnor U27 (N_27,In_9,In_2020);
nand U28 (N_28,In_2063,In_1548);
nor U29 (N_29,In_1076,In_701);
and U30 (N_30,In_1194,In_1042);
nand U31 (N_31,In_807,In_2457);
or U32 (N_32,In_332,In_1913);
nand U33 (N_33,In_2082,In_493);
nand U34 (N_34,In_866,In_834);
nand U35 (N_35,In_122,In_2265);
nor U36 (N_36,In_1949,In_1328);
or U37 (N_37,In_1120,In_278);
nor U38 (N_38,In_850,In_401);
nand U39 (N_39,In_1847,In_2452);
nand U40 (N_40,In_118,In_982);
and U41 (N_41,In_1362,In_241);
or U42 (N_42,In_845,In_711);
or U43 (N_43,In_1097,In_2184);
and U44 (N_44,In_442,In_1508);
nor U45 (N_45,In_2229,In_1836);
nor U46 (N_46,In_1959,In_317);
nand U47 (N_47,In_964,In_500);
nand U48 (N_48,In_2272,In_2471);
nor U49 (N_49,In_1402,In_1123);
nor U50 (N_50,In_1685,In_227);
and U51 (N_51,In_559,In_435);
xor U52 (N_52,In_1476,In_1141);
or U53 (N_53,In_336,In_117);
xnor U54 (N_54,In_1891,In_2326);
nand U55 (N_55,In_2110,In_2172);
nand U56 (N_56,In_2162,In_91);
and U57 (N_57,In_1666,In_1311);
or U58 (N_58,In_735,In_718);
nor U59 (N_59,In_1525,In_1863);
nand U60 (N_60,In_2085,In_1924);
nor U61 (N_61,In_1781,In_1409);
or U62 (N_62,In_1758,In_1001);
nand U63 (N_63,In_1503,In_962);
and U64 (N_64,In_828,In_495);
xor U65 (N_65,In_2041,In_1618);
nand U66 (N_66,In_1158,In_399);
xor U67 (N_67,In_1893,In_2005);
and U68 (N_68,In_1037,In_277);
or U69 (N_69,In_1006,In_1567);
nand U70 (N_70,In_473,In_2032);
and U71 (N_71,In_248,In_2411);
nor U72 (N_72,In_2330,In_1337);
nor U73 (N_73,In_340,In_108);
and U74 (N_74,In_1136,In_1454);
nand U75 (N_75,In_477,In_1229);
or U76 (N_76,In_69,In_1297);
xnor U77 (N_77,In_328,In_1773);
nor U78 (N_78,In_1388,In_2059);
nand U79 (N_79,In_2339,In_2243);
nand U80 (N_80,In_1797,In_1570);
nand U81 (N_81,In_2431,In_525);
or U82 (N_82,In_420,In_746);
and U83 (N_83,In_1214,In_2123);
or U84 (N_84,In_1361,In_2368);
or U85 (N_85,In_889,In_1807);
nor U86 (N_86,In_183,In_2185);
nand U87 (N_87,In_2001,In_402);
xor U88 (N_88,In_1708,In_2458);
xnor U89 (N_89,In_990,In_1143);
nor U90 (N_90,In_1063,In_2417);
xnor U91 (N_91,In_571,In_970);
and U92 (N_92,In_1360,In_1562);
nand U93 (N_93,In_2008,In_1602);
nand U94 (N_94,In_1871,In_322);
nand U95 (N_95,In_598,In_43);
nor U96 (N_96,In_1803,In_1763);
nor U97 (N_97,In_1951,In_712);
and U98 (N_98,In_873,In_67);
xor U99 (N_99,In_1867,In_809);
and U100 (N_100,In_1207,In_1660);
nand U101 (N_101,In_867,In_2386);
or U102 (N_102,In_413,In_1972);
nand U103 (N_103,In_1246,In_196);
nor U104 (N_104,In_1885,In_1600);
nand U105 (N_105,In_1162,In_698);
nand U106 (N_106,In_738,In_1831);
or U107 (N_107,In_1258,In_526);
or U108 (N_108,In_547,In_1517);
nor U109 (N_109,In_682,In_2017);
xnor U110 (N_110,In_795,In_388);
nor U111 (N_111,In_1298,In_914);
nand U112 (N_112,In_1736,In_1678);
nor U113 (N_113,In_347,In_563);
nor U114 (N_114,In_17,In_556);
nand U115 (N_115,In_301,In_1299);
nor U116 (N_116,In_2264,In_1447);
xnor U117 (N_117,In_165,In_2231);
nand U118 (N_118,In_1918,In_1681);
nand U119 (N_119,In_2072,In_1739);
xnor U120 (N_120,In_1093,In_99);
xor U121 (N_121,In_407,In_1745);
and U122 (N_122,In_2488,In_2052);
or U123 (N_123,In_1855,In_1274);
xor U124 (N_124,In_945,In_2331);
or U125 (N_125,In_1278,In_648);
nand U126 (N_126,In_1295,In_1414);
nor U127 (N_127,In_2371,In_1877);
nor U128 (N_128,In_19,In_740);
and U129 (N_129,In_438,In_449);
or U130 (N_130,In_1520,In_2102);
or U131 (N_131,In_2204,In_1864);
nand U132 (N_132,In_1830,In_34);
and U133 (N_133,In_2199,In_2307);
or U134 (N_134,In_1970,In_63);
and U135 (N_135,In_1316,In_1646);
nor U136 (N_136,In_765,In_2334);
and U137 (N_137,In_2442,In_1024);
nand U138 (N_138,In_932,In_2290);
or U139 (N_139,In_2252,In_218);
nor U140 (N_140,In_323,In_1742);
nor U141 (N_141,In_2496,In_1180);
xnor U142 (N_142,In_406,In_1941);
nor U143 (N_143,In_1057,In_973);
and U144 (N_144,In_142,In_1082);
nor U145 (N_145,In_706,In_209);
or U146 (N_146,In_2257,In_2078);
and U147 (N_147,In_2460,In_2163);
and U148 (N_148,In_1248,In_1765);
nor U149 (N_149,In_594,In_2040);
nor U150 (N_150,In_207,In_775);
nor U151 (N_151,In_1801,In_778);
and U152 (N_152,In_833,In_1080);
nor U153 (N_153,In_1509,In_232);
nor U154 (N_154,In_2152,In_1534);
nand U155 (N_155,In_1704,In_853);
xnor U156 (N_156,In_2293,In_194);
or U157 (N_157,In_904,In_1943);
nand U158 (N_158,In_624,In_806);
nand U159 (N_159,In_768,In_351);
nor U160 (N_160,In_1583,In_414);
and U161 (N_161,In_1731,In_2240);
xnor U162 (N_162,In_1649,In_2277);
nor U163 (N_163,In_1254,In_2481);
nor U164 (N_164,In_1135,In_1329);
xor U165 (N_165,In_1793,In_73);
nor U166 (N_166,In_2129,In_1418);
and U167 (N_167,In_8,In_2299);
xnor U168 (N_168,In_2171,In_1198);
or U169 (N_169,In_59,In_1543);
nand U170 (N_170,In_1215,In_1531);
and U171 (N_171,In_1774,In_1677);
nand U172 (N_172,In_2018,In_1990);
or U173 (N_173,In_287,In_236);
and U174 (N_174,In_1630,In_12);
xnor U175 (N_175,In_1698,In_299);
and U176 (N_176,In_676,In_185);
nand U177 (N_177,In_1167,In_2295);
and U178 (N_178,In_1749,In_1225);
nor U179 (N_179,In_1366,In_1500);
nor U180 (N_180,In_1665,In_1713);
nand U181 (N_181,In_2166,In_274);
nand U182 (N_182,In_632,In_842);
nor U183 (N_183,In_583,In_358);
xor U184 (N_184,In_2055,In_1410);
nor U185 (N_185,In_2215,In_1236);
nor U186 (N_186,In_1485,In_1387);
nor U187 (N_187,In_334,In_2088);
and U188 (N_188,In_573,In_2135);
and U189 (N_189,In_1645,In_2443);
or U190 (N_190,In_1714,In_1268);
nand U191 (N_191,In_392,In_604);
and U192 (N_192,In_1945,In_2077);
or U193 (N_193,In_484,In_1494);
and U194 (N_194,In_2356,In_678);
and U195 (N_195,In_265,In_1232);
and U196 (N_196,In_461,In_285);
nor U197 (N_197,In_1292,In_677);
and U198 (N_198,In_1930,In_629);
or U199 (N_199,In_1746,In_151);
or U200 (N_200,In_864,In_2146);
nor U201 (N_201,In_383,In_1211);
nand U202 (N_202,In_1737,In_2434);
nand U203 (N_203,In_742,In_370);
or U204 (N_204,In_44,In_1858);
or U205 (N_205,In_1721,In_1005);
or U206 (N_206,In_247,In_2190);
nand U207 (N_207,In_1072,In_797);
and U208 (N_208,In_408,In_1286);
nor U209 (N_209,In_298,In_2107);
xnor U210 (N_210,In_2387,In_704);
nand U211 (N_211,In_1000,In_149);
or U212 (N_212,In_1445,In_120);
xor U213 (N_213,In_2062,In_1386);
nor U214 (N_214,In_1908,In_1116);
xor U215 (N_215,In_1213,In_2239);
xnor U216 (N_216,In_899,In_346);
or U217 (N_217,In_1786,In_2051);
nand U218 (N_218,In_309,In_164);
nor U219 (N_219,In_1235,In_1091);
xnor U220 (N_220,In_2357,In_799);
and U221 (N_221,In_1291,In_2416);
and U222 (N_222,In_2149,In_4);
nor U223 (N_223,In_773,In_1623);
and U224 (N_224,In_1224,In_814);
and U225 (N_225,In_577,In_2408);
nor U226 (N_226,In_2377,In_969);
nand U227 (N_227,In_830,In_1809);
or U228 (N_228,In_1344,In_1069);
xor U229 (N_229,In_258,In_444);
xnor U230 (N_230,In_1393,In_1521);
nor U231 (N_231,In_2280,In_515);
or U232 (N_232,In_1439,In_308);
nand U233 (N_233,In_1703,In_1022);
nand U234 (N_234,In_1185,In_1629);
or U235 (N_235,In_1969,In_1619);
and U236 (N_236,In_1039,In_922);
nor U237 (N_237,In_2453,In_804);
nand U238 (N_238,In_61,In_649);
nand U239 (N_239,In_1984,In_1635);
or U240 (N_240,In_1866,In_1154);
and U241 (N_241,In_1377,In_936);
nand U242 (N_242,In_617,In_736);
nor U243 (N_243,In_2116,In_45);
nand U244 (N_244,In_269,In_555);
nor U245 (N_245,In_305,In_1150);
and U246 (N_246,In_652,In_716);
or U247 (N_247,In_696,In_747);
or U248 (N_248,In_968,In_2183);
nand U249 (N_249,In_256,In_2499);
and U250 (N_250,In_1892,In_2208);
and U251 (N_251,In_719,In_2424);
nor U252 (N_252,In_1738,In_2091);
or U253 (N_253,In_168,In_64);
xor U254 (N_254,In_585,In_1834);
or U255 (N_255,In_2134,In_1696);
xnor U256 (N_256,In_60,In_1417);
or U257 (N_257,In_2227,In_1284);
or U258 (N_258,In_2254,In_1820);
xor U259 (N_259,In_455,In_633);
nor U260 (N_260,In_2444,In_57);
nor U261 (N_261,In_350,In_1149);
and U262 (N_262,In_523,In_381);
xnor U263 (N_263,In_1617,In_2130);
and U264 (N_264,In_1083,In_319);
and U265 (N_265,In_2459,In_1579);
xor U266 (N_266,In_1455,In_2474);
nand U267 (N_267,In_543,In_874);
nand U268 (N_268,In_1633,In_933);
or U269 (N_269,In_290,In_602);
and U270 (N_270,In_2470,In_90);
nor U271 (N_271,In_1873,In_1962);
nand U272 (N_272,In_213,In_1441);
nand U273 (N_273,In_1428,In_1385);
and U274 (N_274,In_131,In_2451);
and U275 (N_275,In_2292,In_2436);
xnor U276 (N_276,In_1822,In_1747);
nand U277 (N_277,In_1513,In_235);
or U278 (N_278,In_1935,In_1296);
and U279 (N_279,In_518,In_1347);
and U280 (N_280,In_129,In_786);
nor U281 (N_281,In_1796,In_2296);
and U282 (N_282,In_462,In_2031);
nor U283 (N_283,In_2317,In_86);
and U284 (N_284,In_879,In_1159);
or U285 (N_285,In_1456,In_805);
nand U286 (N_286,In_172,In_592);
or U287 (N_287,In_609,In_2385);
nor U288 (N_288,In_894,In_211);
or U289 (N_289,In_915,In_1272);
and U290 (N_290,In_1353,In_2203);
and U291 (N_291,In_116,In_389);
and U292 (N_292,In_2237,In_204);
xor U293 (N_293,In_2406,In_1186);
and U294 (N_294,In_1880,In_1301);
or U295 (N_295,In_2214,In_1563);
nor U296 (N_296,In_1359,In_2284);
nand U297 (N_297,In_1744,In_753);
and U298 (N_298,In_2177,In_785);
nor U299 (N_299,In_844,In_1785);
nor U300 (N_300,In_450,In_1373);
and U301 (N_301,In_2122,In_1419);
and U302 (N_302,In_841,In_1533);
and U303 (N_303,In_1166,In_910);
nand U304 (N_304,In_2491,In_1589);
or U305 (N_305,In_2044,In_33);
nor U306 (N_306,In_1089,In_789);
nand U307 (N_307,In_987,In_854);
and U308 (N_308,In_1495,In_18);
and U309 (N_309,In_513,In_934);
nand U310 (N_310,In_2086,In_2038);
xnor U311 (N_311,In_254,In_2150);
or U312 (N_312,In_79,In_1070);
and U313 (N_313,In_1112,In_2103);
or U314 (N_314,In_2300,In_1333);
and U315 (N_315,In_2173,In_201);
nand U316 (N_316,In_955,In_2260);
nor U317 (N_317,In_1730,In_1059);
and U318 (N_318,In_2447,In_745);
nand U319 (N_319,In_699,In_2034);
and U320 (N_320,In_1113,In_1733);
or U321 (N_321,In_627,In_1046);
nor U322 (N_322,In_1884,In_1768);
or U323 (N_323,In_1265,In_2169);
or U324 (N_324,In_901,In_2362);
nand U325 (N_325,In_2267,In_1233);
and U326 (N_326,In_1647,In_2024);
nor U327 (N_327,In_2490,In_1461);
and U328 (N_328,In_1147,In_1405);
and U329 (N_329,In_887,In_35);
nand U330 (N_330,In_1110,In_1537);
and U331 (N_331,In_2346,In_2242);
nand U332 (N_332,In_1102,In_663);
or U333 (N_333,In_1887,In_2303);
and U334 (N_334,In_1661,In_2108);
or U335 (N_335,In_466,In_1912);
or U336 (N_336,In_1427,In_2432);
and U337 (N_337,In_863,In_13);
or U338 (N_338,In_2164,In_958);
or U339 (N_339,In_1605,In_2430);
and U340 (N_340,In_1436,In_242);
or U341 (N_341,In_1302,In_1132);
or U342 (N_342,In_950,In_1400);
nor U343 (N_343,In_2333,In_1818);
and U344 (N_344,In_1870,In_997);
and U345 (N_345,In_162,In_292);
xnor U346 (N_346,In_1028,In_318);
and U347 (N_347,In_324,In_212);
nor U348 (N_348,In_1999,In_2094);
nand U349 (N_349,In_1595,In_1364);
or U350 (N_350,In_2493,In_2461);
or U351 (N_351,In_2355,In_1261);
and U352 (N_352,In_584,In_2275);
and U353 (N_353,In_638,In_1289);
and U354 (N_354,In_2492,In_1980);
and U355 (N_355,In_1052,In_1073);
or U356 (N_356,In_1408,In_2429);
or U357 (N_357,In_641,In_1313);
nor U358 (N_358,In_1025,In_41);
or U359 (N_359,In_2392,In_1897);
or U360 (N_360,In_664,In_101);
nand U361 (N_361,In_1068,In_1540);
and U362 (N_362,In_1078,In_672);
or U363 (N_363,In_2439,In_725);
or U364 (N_364,In_1305,In_2101);
xor U365 (N_365,In_1416,In_2067);
or U366 (N_366,In_1222,In_2318);
nor U367 (N_367,In_1691,In_132);
and U368 (N_368,In_104,In_333);
nor U369 (N_369,In_2092,In_1907);
nor U370 (N_370,In_2251,In_1909);
nand U371 (N_371,In_1869,In_1269);
and U372 (N_372,In_1391,In_2035);
xor U373 (N_373,In_2263,In_727);
nand U374 (N_374,In_1824,In_1694);
nor U375 (N_375,In_1477,In_1356);
nand U376 (N_376,In_608,In_974);
and U377 (N_377,In_1620,In_1875);
xor U378 (N_378,In_2310,In_280);
and U379 (N_379,In_2370,In_100);
and U380 (N_380,In_1852,In_426);
and U381 (N_381,In_390,In_417);
or U382 (N_382,In_1199,In_669);
nand U383 (N_383,In_829,In_1055);
nand U384 (N_384,In_1053,In_1898);
nor U385 (N_385,In_1004,In_2202);
or U386 (N_386,In_1491,In_1242);
nand U387 (N_387,In_1420,In_1833);
nor U388 (N_388,In_1290,In_233);
xnor U389 (N_389,In_176,In_1011);
or U390 (N_390,In_1507,In_1524);
nor U391 (N_391,In_1241,In_345);
or U392 (N_392,In_2405,In_2332);
and U393 (N_393,In_1003,In_1812);
and U394 (N_394,In_1710,In_1064);
nor U395 (N_395,In_2142,In_1451);
nor U396 (N_396,In_2403,In_2191);
nand U397 (N_397,In_1784,In_2137);
nand U398 (N_398,In_565,In_1486);
nand U399 (N_399,In_70,In_84);
and U400 (N_400,In_249,In_102);
nor U401 (N_401,In_520,In_1146);
nand U402 (N_402,In_145,In_1839);
nor U403 (N_403,In_1608,In_1558);
nand U404 (N_404,In_0,In_83);
nor U405 (N_405,In_1253,In_593);
and U406 (N_406,In_801,In_705);
nand U407 (N_407,In_423,In_467);
nand U408 (N_408,In_222,In_1170);
or U409 (N_409,In_686,In_1819);
or U410 (N_410,In_822,In_927);
nor U411 (N_411,In_2075,In_198);
and U412 (N_412,In_475,In_1624);
nor U413 (N_413,In_1559,In_2194);
and U414 (N_414,In_511,In_1474);
xnor U415 (N_415,In_238,In_219);
xnor U416 (N_416,In_1842,In_1363);
nand U417 (N_417,In_2445,In_25);
or U418 (N_418,In_2147,In_1823);
and U419 (N_419,In_1648,In_38);
nor U420 (N_420,In_1560,In_816);
nand U421 (N_421,In_549,In_1306);
nor U422 (N_422,In_1860,In_2157);
nor U423 (N_423,In_739,In_337);
and U424 (N_424,In_395,In_1121);
nor U425 (N_425,In_749,In_681);
xnor U426 (N_426,In_1769,In_1881);
or U427 (N_427,In_535,In_2383);
nor U428 (N_428,In_1105,In_1518);
or U429 (N_429,In_1740,In_1156);
xnor U430 (N_430,In_10,In_2158);
or U431 (N_431,In_1148,In_1653);
or U432 (N_432,In_994,In_540);
xnor U433 (N_433,In_271,In_1020);
or U434 (N_434,In_2329,In_155);
xnor U435 (N_435,In_276,In_1826);
and U436 (N_436,In_1716,In_1953);
nand U437 (N_437,In_991,In_1045);
and U438 (N_438,In_2369,In_1526);
nor U439 (N_439,In_2197,In_1392);
xor U440 (N_440,In_1644,In_1549);
nor U441 (N_441,In_1902,In_1193);
and U442 (N_442,In_957,In_1806);
or U443 (N_443,In_3,In_396);
nand U444 (N_444,In_897,In_1168);
nor U445 (N_445,In_926,In_1536);
or U446 (N_446,In_2466,In_1100);
and U447 (N_447,In_675,In_321);
and U448 (N_448,In_2084,In_748);
nand U449 (N_449,In_1075,In_903);
nor U450 (N_450,In_2455,In_42);
or U451 (N_451,In_234,In_642);
nand U452 (N_452,In_1249,In_1937);
or U453 (N_453,In_2047,In_1354);
or U454 (N_454,In_623,In_530);
nand U455 (N_455,In_1270,In_1457);
and U456 (N_456,In_1956,In_1844);
or U457 (N_457,In_2396,In_846);
and U458 (N_458,In_1725,In_1695);
xor U459 (N_459,In_1779,In_39);
and U460 (N_460,In_2249,In_2012);
nor U461 (N_461,In_2168,In_707);
and U462 (N_462,In_421,In_143);
xor U463 (N_463,In_838,In_1030);
nor U464 (N_464,In_921,In_1637);
or U465 (N_465,In_2019,In_569);
and U466 (N_466,In_427,In_1625);
or U467 (N_467,In_2037,In_491);
xor U468 (N_468,In_658,In_110);
or U469 (N_469,In_1950,In_2328);
xnor U470 (N_470,In_597,In_2033);
xnor U471 (N_471,In_1122,In_1621);
nand U472 (N_472,In_1652,In_868);
xor U473 (N_473,In_800,In_2124);
or U474 (N_474,In_875,In_349);
nor U475 (N_475,In_432,In_1169);
nand U476 (N_476,In_224,In_107);
nor U477 (N_477,In_2216,In_405);
and U478 (N_478,In_1805,In_870);
nor U479 (N_479,In_1111,In_810);
or U480 (N_480,In_37,In_2278);
and U481 (N_481,In_11,In_1231);
xnor U482 (N_482,In_48,In_1800);
and U483 (N_483,In_743,In_772);
nor U484 (N_484,In_1978,In_787);
nor U485 (N_485,In_1411,In_2321);
xor U486 (N_486,In_1255,In_1815);
and U487 (N_487,In_2193,In_791);
or U488 (N_488,In_1865,In_1547);
xor U489 (N_489,In_2117,In_480);
xnor U490 (N_490,In_848,In_159);
nand U491 (N_491,In_802,In_158);
and U492 (N_492,In_148,In_521);
nor U493 (N_493,In_1551,In_440);
or U494 (N_494,In_1425,In_2325);
or U495 (N_495,In_542,In_1942);
nor U496 (N_496,In_2112,In_722);
nor U497 (N_497,In_1153,In_517);
xor U498 (N_498,In_275,In_1964);
nand U499 (N_499,In_630,In_1051);
xor U500 (N_500,In_732,In_919);
or U501 (N_501,In_2352,In_1048);
or U502 (N_502,In_1667,In_925);
or U503 (N_503,In_2495,In_948);
xnor U504 (N_504,In_2388,In_1240);
and U505 (N_505,In_2446,In_2427);
nand U506 (N_506,In_516,In_1191);
or U507 (N_507,In_1182,In_20);
and U508 (N_508,In_2138,In_1986);
or U509 (N_509,In_1849,In_1175);
nor U510 (N_510,In_920,In_181);
or U511 (N_511,In_684,In_1614);
xnor U512 (N_512,In_510,In_1103);
nor U513 (N_513,In_246,In_1294);
nor U514 (N_514,In_1933,In_1944);
and U515 (N_515,In_1584,In_2175);
nand U516 (N_516,In_2483,In_1041);
or U517 (N_517,In_214,In_1401);
nand U518 (N_518,In_783,In_1751);
or U519 (N_519,In_1352,In_1783);
or U520 (N_520,In_55,In_56);
nand U521 (N_521,In_1099,In_1165);
or U522 (N_522,In_1394,In_1840);
or U523 (N_523,In_659,In_1587);
xor U524 (N_524,In_362,In_1923);
or U525 (N_525,In_1376,In_2376);
or U526 (N_526,In_776,In_2007);
or U527 (N_527,In_434,In_1047);
xor U528 (N_528,In_2353,In_673);
or U529 (N_529,In_503,In_1217);
nand U530 (N_530,In_645,In_1899);
or U531 (N_531,In_771,In_286);
or U532 (N_532,In_817,In_566);
and U533 (N_533,In_46,In_1903);
xnor U534 (N_534,In_228,In_2367);
and U535 (N_535,In_335,In_1511);
and U536 (N_536,In_2351,In_930);
and U537 (N_537,In_1281,In_1967);
nor U538 (N_538,In_1672,In_2201);
nand U539 (N_539,In_628,In_2494);
nor U540 (N_540,In_1640,In_557);
or U541 (N_541,In_1239,In_2010);
nor U542 (N_542,In_32,In_1501);
or U543 (N_543,In_2176,In_124);
or U544 (N_544,In_2391,In_1267);
and U545 (N_545,In_266,In_1770);
nand U546 (N_546,In_1998,In_1342);
nand U547 (N_547,In_1811,In_325);
nand U548 (N_548,In_796,In_562);
nand U549 (N_549,In_1139,In_524);
nand U550 (N_550,In_1993,In_2304);
xor U551 (N_551,In_2354,In_1780);
and U552 (N_552,In_352,In_1960);
or U553 (N_553,In_996,In_1921);
xor U554 (N_554,In_357,In_2097);
xnor U555 (N_555,In_1914,In_121);
nor U556 (N_556,In_267,In_1176);
nand U557 (N_557,In_1606,In_1627);
nand U558 (N_558,In_693,In_1828);
nor U559 (N_559,In_827,In_1412);
nor U560 (N_560,In_529,In_199);
nor U561 (N_561,In_2400,In_469);
xor U562 (N_562,In_2311,In_1309);
or U563 (N_563,In_506,In_1443);
or U564 (N_564,In_2115,In_1615);
nand U565 (N_565,In_956,In_2143);
nor U566 (N_566,In_544,In_2066);
or U567 (N_567,In_1424,In_1415);
and U568 (N_568,In_2128,In_1516);
or U569 (N_569,In_1756,In_1670);
nand U570 (N_570,In_1426,In_1219);
nor U571 (N_571,In_509,In_878);
nand U572 (N_572,In_813,In_180);
or U573 (N_573,In_574,In_811);
nand U574 (N_574,In_620,In_1192);
or U575 (N_575,In_2132,In_784);
xor U576 (N_576,In_1915,In_250);
or U577 (N_577,In_2437,In_788);
nand U578 (N_578,In_1350,In_448);
nand U579 (N_579,In_7,In_622);
nor U580 (N_580,In_1038,In_891);
nor U581 (N_581,In_626,In_1544);
nand U582 (N_582,In_1395,In_1916);
or U583 (N_583,In_452,In_939);
and U584 (N_584,In_1611,In_2382);
xor U585 (N_585,In_2273,In_1396);
or U586 (N_586,In_1300,In_1378);
xor U587 (N_587,In_1221,In_1118);
and U588 (N_588,In_2454,In_582);
nor U589 (N_589,In_558,In_1755);
xnor U590 (N_590,In_1275,In_2380);
xor U591 (N_591,In_1015,In_690);
and U592 (N_592,In_1040,In_1279);
and U593 (N_593,In_66,In_741);
and U594 (N_594,In_1900,In_689);
xnor U595 (N_595,In_1271,In_1687);
nor U596 (N_596,In_2029,In_182);
or U597 (N_597,In_998,In_1724);
xnor U598 (N_598,In_353,In_1701);
or U599 (N_599,In_186,In_928);
nor U600 (N_600,In_1204,In_312);
and U601 (N_601,In_1137,In_1683);
xnor U602 (N_602,In_2359,In_203);
xnor U603 (N_603,In_587,In_15);
nor U604 (N_604,In_1789,In_1230);
nor U605 (N_605,In_393,In_415);
xor U606 (N_606,In_1821,In_615);
nand U607 (N_607,In_419,In_572);
nand U608 (N_608,In_1307,In_5);
and U609 (N_609,In_1712,In_1981);
or U610 (N_610,In_1195,In_487);
nand U611 (N_611,In_2006,In_29);
nand U612 (N_612,In_152,In_1010);
nand U613 (N_613,In_946,In_2218);
nand U614 (N_614,In_1827,In_1023);
nor U615 (N_615,In_2151,In_2180);
and U616 (N_616,In_1607,In_825);
nand U617 (N_617,In_770,In_709);
and U618 (N_618,In_1722,In_146);
nand U619 (N_619,In_545,In_163);
xnor U620 (N_620,In_902,In_631);
and U621 (N_621,In_1861,In_1926);
nor U622 (N_622,In_522,In_1310);
or U623 (N_623,In_1929,In_847);
nor U624 (N_624,In_2046,In_1228);
nor U625 (N_625,In_1735,In_2256);
nand U626 (N_626,In_1223,In_2200);
or U627 (N_627,In_720,In_137);
nand U628 (N_628,In_2363,In_2297);
or U629 (N_629,In_1762,In_293);
nor U630 (N_630,In_723,In_714);
nand U631 (N_631,In_2011,In_803);
and U632 (N_632,In_1838,In_1804);
and U633 (N_633,In_935,In_2258);
nor U634 (N_634,In_812,In_2410);
and U635 (N_635,In_931,In_1775);
nand U636 (N_636,In_1662,In_941);
and U637 (N_637,In_532,In_754);
nor U638 (N_638,In_2395,In_852);
and U639 (N_639,In_331,In_1188);
and U640 (N_640,In_942,In_1338);
and U641 (N_641,In_77,In_2287);
or U642 (N_642,In_1452,In_655);
or U643 (N_643,In_514,In_1058);
xnor U644 (N_644,In_2282,In_443);
nand U645 (N_645,In_605,In_1398);
nand U646 (N_646,In_193,In_157);
nand U647 (N_647,In_1065,In_1974);
nor U648 (N_648,In_1671,In_504);
nand U649 (N_649,In_1987,In_2366);
nand U650 (N_650,In_273,In_943);
and U651 (N_651,In_1012,In_2423);
or U652 (N_652,In_1019,In_1682);
nor U653 (N_653,In_195,In_832);
or U654 (N_654,In_1613,In_2478);
nand U655 (N_655,In_1965,In_1952);
xnor U656 (N_656,In_1654,In_1889);
or U657 (N_657,In_1505,In_906);
and U658 (N_658,In_2428,In_1568);
nand U659 (N_659,In_855,In_1673);
and U660 (N_660,In_662,In_1098);
or U661 (N_661,In_1971,In_361);
and U662 (N_662,In_750,In_95);
nor U663 (N_663,In_244,In_1920);
nor U664 (N_664,In_486,In_1067);
or U665 (N_665,In_1319,In_2219);
nand U666 (N_666,In_1574,In_179);
and U667 (N_667,In_161,In_1375);
and U668 (N_668,In_369,In_72);
nand U669 (N_669,In_2105,In_428);
and U670 (N_670,In_2337,In_1034);
nor U671 (N_671,In_2327,In_71);
or U672 (N_672,In_1802,In_1471);
or U673 (N_673,In_1129,In_49);
nor U674 (N_674,In_2271,In_951);
nand U675 (N_675,In_1857,In_1133);
and U676 (N_676,In_710,In_1992);
xnor U677 (N_677,In_2222,In_995);
or U678 (N_678,In_454,In_918);
nor U679 (N_679,In_36,In_1383);
and U680 (N_680,In_314,In_1304);
or U681 (N_681,In_1979,In_226);
nand U682 (N_682,In_2279,In_31);
nor U683 (N_683,In_190,In_446);
nand U684 (N_684,In_2479,In_2475);
nor U685 (N_685,In_2213,In_790);
nor U686 (N_686,In_1994,In_611);
nor U687 (N_687,In_1079,In_618);
and U688 (N_688,In_88,In_888);
and U689 (N_689,In_456,In_130);
or U690 (N_690,In_1390,In_1659);
nor U691 (N_691,In_306,In_1925);
or U692 (N_692,In_1026,In_264);
and U693 (N_693,In_191,In_221);
xor U694 (N_694,In_890,In_2407);
nor U695 (N_695,In_1706,In_54);
nand U696 (N_696,In_2114,In_2139);
or U697 (N_697,In_65,In_1458);
or U698 (N_698,In_2090,In_661);
and U699 (N_699,In_575,In_1502);
nor U700 (N_700,In_2312,In_1656);
and U701 (N_701,In_2021,In_437);
nand U702 (N_702,In_1448,In_924);
or U703 (N_703,In_75,In_1315);
xnor U704 (N_704,In_1095,In_940);
nand U705 (N_705,In_189,In_1764);
and U706 (N_706,In_1318,In_1901);
nand U707 (N_707,In_1798,In_1552);
nor U708 (N_708,In_231,In_2083);
and U709 (N_709,In_937,In_1252);
and U710 (N_710,In_429,In_1475);
nand U711 (N_711,In_1966,In_1071);
nand U712 (N_712,In_1514,In_433);
xnor U713 (N_713,In_327,In_2476);
nand U714 (N_714,In_2050,In_560);
nor U715 (N_715,In_2268,In_1326);
or U716 (N_716,In_1905,In_202);
nand U717 (N_717,In_619,In_595);
xor U718 (N_718,In_2415,In_2226);
and U719 (N_719,In_1931,In_1989);
nand U720 (N_720,In_1203,In_366);
and U721 (N_721,In_568,In_757);
and U722 (N_722,In_650,In_237);
nor U723 (N_723,In_1109,In_2087);
and U724 (N_724,In_551,In_113);
and U725 (N_725,In_1497,In_1843);
and U726 (N_726,In_1470,In_2014);
or U727 (N_727,In_798,In_668);
or U728 (N_728,In_715,In_1841);
nor U729 (N_729,In_1968,In_621);
nand U730 (N_730,In_1689,In_1963);
nor U731 (N_731,In_294,In_646);
and U732 (N_732,In_880,In_979);
and U733 (N_733,In_1370,In_965);
or U734 (N_734,In_338,In_653);
and U735 (N_735,In_1173,In_1572);
nor U736 (N_736,In_1324,In_1663);
or U737 (N_737,In_119,In_539);
nor U738 (N_738,In_2418,In_695);
or U739 (N_739,In_774,In_307);
nor U740 (N_740,In_326,In_1565);
xnor U741 (N_741,In_154,In_1530);
or U742 (N_742,In_737,In_1961);
nor U743 (N_743,In_1450,In_2141);
or U744 (N_744,In_1947,In_2360);
nand U745 (N_745,In_2441,In_1700);
and U746 (N_746,In_1566,In_1753);
nor U747 (N_747,In_1594,In_485);
nand U748 (N_748,In_471,In_1504);
and U749 (N_749,In_2261,In_1939);
or U750 (N_750,In_2238,In_1750);
nor U751 (N_751,In_2140,In_2489);
nor U752 (N_752,In_2420,In_2350);
nand U753 (N_753,In_2131,In_382);
nand U754 (N_754,In_2127,In_139);
nand U755 (N_755,In_94,In_177);
nand U756 (N_756,In_1054,In_2419);
nor U757 (N_757,In_1596,In_412);
and U758 (N_758,In_229,In_781);
nand U759 (N_759,In_1056,In_1590);
xnor U760 (N_760,In_637,In_634);
xor U761 (N_761,In_376,In_856);
or U762 (N_762,In_1578,In_2049);
nand U763 (N_763,In_394,In_1546);
or U764 (N_764,In_680,In_793);
or U765 (N_765,In_599,In_1380);
or U766 (N_766,In_1467,In_2378);
nand U767 (N_767,In_683,In_2160);
nand U768 (N_768,In_1260,In_459);
or U769 (N_769,In_2438,In_2119);
or U770 (N_770,In_2281,In_877);
nor U771 (N_771,In_136,In_1179);
and U772 (N_772,In_1718,In_1066);
and U773 (N_773,In_343,In_1856);
xnor U774 (N_774,In_230,In_1106);
and U775 (N_775,In_756,In_2155);
nand U776 (N_776,In_2013,In_860);
or U777 (N_777,In_697,In_1711);
or U778 (N_778,In_14,In_2209);
or U779 (N_779,In_665,In_1727);
nor U780 (N_780,In_1876,In_993);
or U781 (N_781,In_2245,In_1124);
and U782 (N_782,In_378,In_144);
nand U783 (N_783,In_1085,In_2253);
nor U784 (N_784,In_881,In_464);
nand U785 (N_785,In_1832,In_215);
nand U786 (N_786,In_1493,In_766);
nand U787 (N_787,In_1772,In_538);
nand U788 (N_788,In_978,In_150);
xnor U789 (N_789,In_2379,In_169);
nand U790 (N_790,In_1013,In_2309);
and U791 (N_791,In_581,In_425);
or U792 (N_792,In_492,In_197);
nand U793 (N_793,In_330,In_541);
nor U794 (N_794,In_1609,In_2348);
nand U795 (N_795,In_2136,In_553);
nand U796 (N_796,In_508,In_898);
nand U797 (N_797,In_1332,In_1825);
and U798 (N_798,In_304,In_2394);
or U799 (N_799,In_916,In_2004);
or U800 (N_800,In_818,In_734);
or U801 (N_801,In_1808,In_865);
nand U802 (N_802,In_1904,In_839);
or U803 (N_803,In_580,In_1101);
nand U804 (N_804,In_2322,In_913);
and U805 (N_805,In_2182,In_2196);
or U806 (N_806,In_1431,In_2054);
nand U807 (N_807,In_909,In_2285);
and U808 (N_808,In_1948,In_1976);
nand U809 (N_809,In_687,In_667);
nor U810 (N_810,In_125,In_377);
nand U811 (N_811,In_2393,In_138);
nor U812 (N_812,In_1778,In_1752);
or U813 (N_813,In_2413,In_379);
or U814 (N_814,In_2125,In_2221);
nand U815 (N_815,In_1799,In_1460);
nor U816 (N_816,In_208,In_1487);
or U817 (N_817,In_823,In_171);
nand U818 (N_818,In_1435,In_2153);
nor U819 (N_819,In_1145,In_2220);
or U820 (N_820,In_329,In_1610);
nor U821 (N_821,In_1490,In_519);
or U822 (N_822,In_1466,In_1792);
xnor U823 (N_823,In_1357,In_1657);
nand U824 (N_824,In_1688,In_1453);
nand U825 (N_825,In_1946,In_2414);
or U826 (N_826,In_360,In_2302);
or U827 (N_827,In_483,In_1190);
nor U828 (N_828,In_1312,In_2025);
nand U829 (N_829,In_1720,In_606);
nand U830 (N_830,In_1553,In_1152);
nand U831 (N_831,In_253,In_1896);
and U832 (N_832,In_840,In_2343);
nand U833 (N_833,In_1616,In_1340);
nor U834 (N_834,In_1919,In_1601);
and U835 (N_835,In_1519,In_1754);
xnor U836 (N_836,In_578,In_82);
nand U837 (N_837,In_223,In_1335);
nor U838 (N_838,In_1339,In_2324);
nand U839 (N_839,In_170,In_1174);
nor U840 (N_840,In_111,In_1197);
and U841 (N_841,In_2250,In_1557);
and U842 (N_842,In_1092,In_1564);
and U843 (N_843,In_2498,In_2099);
nand U844 (N_844,In_380,In_1591);
nand U845 (N_845,In_2345,In_479);
and U846 (N_846,In_884,In_1636);
xor U847 (N_847,In_2060,In_30);
nand U848 (N_848,In_502,In_1227);
nand U849 (N_849,In_2056,In_1599);
or U850 (N_850,In_188,In_2465);
and U851 (N_851,In_1201,In_2000);
and U852 (N_852,In_1853,In_2093);
and U853 (N_853,In_2323,In_730);
xnor U854 (N_854,In_760,In_1664);
nor U855 (N_855,In_81,In_192);
and U856 (N_856,In_1459,In_463);
nand U857 (N_857,In_1729,In_78);
or U858 (N_858,In_1358,In_2217);
nor U859 (N_859,In_724,In_1555);
nand U860 (N_860,In_929,In_1906);
nand U861 (N_861,In_175,In_2262);
nor U862 (N_862,In_490,In_6);
or U863 (N_863,In_458,In_896);
and U864 (N_864,In_1668,In_1355);
nand U865 (N_865,In_2126,In_567);
and U866 (N_866,In_908,In_187);
xor U867 (N_867,In_1033,In_1846);
or U868 (N_868,In_1128,In_2016);
or U869 (N_869,In_16,In_729);
nor U870 (N_870,In_1707,In_1632);
nand U871 (N_871,In_1556,In_1488);
or U872 (N_872,In_386,In_1317);
nand U873 (N_873,In_651,In_971);
or U874 (N_874,In_410,In_1651);
or U875 (N_875,In_1131,In_507);
nand U876 (N_876,In_2336,In_763);
and U877 (N_877,In_431,In_1975);
nor U878 (N_878,In_1597,In_2120);
nand U879 (N_879,In_1539,In_1226);
or U880 (N_880,In_1257,In_1202);
nand U881 (N_881,In_92,In_1266);
and U882 (N_882,In_2179,In_564);
or U883 (N_883,In_1977,In_2365);
or U884 (N_884,In_1469,In_892);
or U885 (N_885,In_612,In_976);
nand U886 (N_886,In_1715,In_1554);
and U887 (N_887,In_1161,In_1138);
and U888 (N_888,In_536,In_418);
and U889 (N_889,In_534,In_374);
nand U890 (N_890,In_1094,In_279);
nor U891 (N_891,In_1982,In_2036);
nand U892 (N_892,In_1973,In_178);
nor U893 (N_893,In_992,In_1741);
xor U894 (N_894,In_364,In_240);
nand U895 (N_895,In_685,In_2421);
nand U896 (N_896,In_2079,In_2486);
nand U897 (N_897,In_2338,In_1638);
or U898 (N_898,In_1178,In_2096);
and U899 (N_899,In_590,In_216);
and U900 (N_900,In_1086,In_2064);
nand U901 (N_901,In_1287,In_27);
nand U902 (N_902,In_527,In_2022);
and U903 (N_903,In_1837,In_2074);
or U904 (N_904,In_2118,In_1788);
nor U905 (N_905,In_1492,In_2315);
nand U906 (N_906,In_1007,In_1125);
or U907 (N_907,In_596,In_2080);
nand U908 (N_908,In_436,In_656);
nor U909 (N_909,In_1626,In_96);
nor U910 (N_910,In_1814,In_952);
nor U911 (N_911,In_1676,In_591);
xnor U912 (N_912,In_694,In_2440);
xnor U913 (N_913,In_1845,In_2289);
and U914 (N_914,In_2341,In_561);
and U915 (N_915,In_1911,In_251);
and U916 (N_916,In_1872,In_303);
or U917 (N_917,In_21,In_999);
nand U918 (N_918,In_2,In_453);
or U919 (N_919,In_282,In_2070);
nor U920 (N_920,In_601,In_713);
nor U921 (N_921,In_1234,In_1642);
nor U922 (N_922,In_1669,In_1468);
nor U923 (N_923,In_1985,In_1795);
and U924 (N_924,In_1346,In_2167);
and U925 (N_925,In_384,In_1108);
nand U926 (N_926,In_2148,In_210);
or U927 (N_927,In_849,In_1498);
and U928 (N_928,In_1096,In_1140);
or U929 (N_929,In_1422,In_2081);
and U930 (N_930,In_2426,In_1479);
or U931 (N_931,In_2048,In_717);
xnor U932 (N_932,In_2113,In_239);
nand U933 (N_933,In_1934,In_478);
nand U934 (N_934,In_166,In_831);
or U935 (N_935,In_398,In_1432);
nand U936 (N_936,In_2043,In_1895);
and U937 (N_937,In_2224,In_972);
and U938 (N_938,In_1288,In_905);
and U939 (N_939,In_531,In_550);
nor U940 (N_940,In_310,In_2372);
or U941 (N_941,In_283,In_726);
nor U942 (N_942,In_794,In_1612);
nor U943 (N_943,In_1327,In_2174);
and U944 (N_944,In_1686,In_614);
nor U945 (N_945,In_1588,In_445);
nor U946 (N_946,In_2145,In_923);
xnor U947 (N_947,In_983,In_1181);
nor U948 (N_948,In_1160,In_2404);
nor U949 (N_949,In_576,In_1573);
xor U950 (N_950,In_782,In_105);
xor U951 (N_951,In_134,In_1690);
or U952 (N_952,In_959,In_1280);
nand U953 (N_953,In_603,In_2236);
or U954 (N_954,In_2189,In_2401);
nand U955 (N_955,In_2373,In_1894);
nor U956 (N_956,In_2109,In_769);
or U957 (N_957,In_430,In_824);
and U958 (N_958,In_1522,In_2023);
nand U959 (N_959,In_1541,In_949);
nor U960 (N_960,In_1882,In_821);
or U961 (N_961,In_2384,In_1444);
xor U962 (N_962,In_98,In_1776);
or U963 (N_963,In_1791,In_1499);
nor U964 (N_964,In_311,In_1890);
or U965 (N_965,In_2286,In_1367);
nor U966 (N_966,In_610,In_2042);
nor U967 (N_967,In_291,In_62);
xnor U968 (N_968,In_640,In_1478);
and U969 (N_969,In_22,In_1680);
nor U970 (N_970,In_1465,In_1983);
and U971 (N_971,In_1586,In_1384);
nand U972 (N_972,In_548,In_963);
or U973 (N_973,In_1430,In_639);
or U974 (N_974,In_270,In_302);
or U975 (N_975,In_411,In_2206);
xnor U976 (N_976,In_759,In_2283);
xor U977 (N_977,In_1940,In_2485);
and U978 (N_978,In_1813,In_2448);
nor U979 (N_979,In_206,In_1238);
nor U980 (N_980,In_156,In_1308);
and U981 (N_981,In_1527,In_819);
and U982 (N_982,In_1151,In_1777);
nand U983 (N_983,In_954,In_764);
or U984 (N_984,In_1761,In_1592);
nor U985 (N_985,In_1200,In_1349);
or U986 (N_986,In_1404,In_657);
or U987 (N_987,In_220,In_1081);
nor U988 (N_988,In_160,In_416);
xor U989 (N_989,In_1351,In_1008);
xnor U990 (N_990,In_2165,In_2433);
nand U991 (N_991,In_1580,In_2425);
and U992 (N_992,In_2320,In_1561);
nand U993 (N_993,In_700,In_2234);
and U994 (N_994,In_28,In_1675);
and U995 (N_995,In_2071,In_554);
or U996 (N_996,In_1496,In_1910);
or U997 (N_997,In_1879,In_1245);
and U998 (N_998,In_767,In_869);
nor U999 (N_999,In_1262,In_2244);
or U1000 (N_1000,In_1854,In_1336);
or U1001 (N_1001,In_1061,In_2045);
and U1002 (N_1002,In_691,In_2207);
nand U1003 (N_1003,In_2068,In_147);
nor U1004 (N_1004,In_666,In_272);
nand U1005 (N_1005,In_1446,In_1743);
xor U1006 (N_1006,In_498,In_900);
or U1007 (N_1007,In_1787,In_1550);
xor U1008 (N_1008,In_1379,In_1922);
and U1009 (N_1009,In_1874,In_858);
and U1010 (N_1010,In_372,In_947);
nand U1011 (N_1011,In_2003,In_268);
nor U1012 (N_1012,In_2456,In_552);
xor U1013 (N_1013,In_2487,In_115);
nor U1014 (N_1014,In_2298,In_1196);
or U1015 (N_1015,In_1371,In_671);
nor U1016 (N_1016,In_1734,In_2015);
or U1017 (N_1017,In_85,In_780);
and U1018 (N_1018,In_1434,In_2274);
or U1019 (N_1019,In_184,In_988);
and U1020 (N_1020,In_1515,In_2027);
nor U1021 (N_1021,In_1571,In_1382);
and U1022 (N_1022,In_1277,In_579);
or U1023 (N_1023,In_883,In_1077);
and U1024 (N_1024,In_2248,In_1684);
nand U1025 (N_1025,In_1341,In_2450);
nor U1026 (N_1026,In_2225,In_1369);
and U1027 (N_1027,In_1205,In_344);
nand U1028 (N_1028,In_123,In_2195);
and U1029 (N_1029,In_2301,In_2381);
and U1030 (N_1030,In_1473,In_1183);
nor U1031 (N_1031,In_1429,In_1062);
or U1032 (N_1032,In_1603,In_2255);
or U1033 (N_1033,In_1413,In_1650);
nor U1034 (N_1034,In_2154,In_1658);
and U1035 (N_1035,In_460,In_1760);
nor U1036 (N_1036,In_1142,In_2412);
nand U1037 (N_1037,In_2210,In_1050);
or U1038 (N_1038,In_1529,In_859);
nand U1039 (N_1039,In_505,In_1483);
nor U1040 (N_1040,In_1285,In_2276);
nand U1041 (N_1041,In_2306,In_1631);
nand U1042 (N_1042,In_133,In_2198);
nand U1043 (N_1043,In_404,In_2058);
nor U1044 (N_1044,In_497,In_2462);
and U1045 (N_1045,In_2009,In_320);
and U1046 (N_1046,In_2246,In_1757);
nand U1047 (N_1047,In_174,In_613);
nand U1048 (N_1048,In_2361,In_1928);
nand U1049 (N_1049,In_1259,In_1848);
nor U1050 (N_1050,In_2467,In_2188);
or U1051 (N_1051,In_2076,In_1545);
nor U1052 (N_1052,In_2111,In_2098);
or U1053 (N_1053,In_1049,In_1117);
nor U1054 (N_1054,In_47,In_1321);
and U1055 (N_1055,In_288,In_1489);
nor U1056 (N_1056,In_375,In_1325);
and U1057 (N_1057,In_1697,In_1323);
nor U1058 (N_1058,In_1088,In_1927);
nor U1059 (N_1059,In_40,In_1542);
nor U1060 (N_1060,In_636,In_2358);
and U1061 (N_1061,In_2156,In_1593);
nand U1062 (N_1062,In_1184,In_501);
nand U1063 (N_1063,In_2389,In_2073);
nand U1064 (N_1064,In_2335,In_588);
nand U1065 (N_1065,In_1581,In_313);
nand U1066 (N_1066,In_1835,In_257);
or U1067 (N_1067,In_1210,In_1206);
and U1068 (N_1068,In_2375,In_703);
nor U1069 (N_1069,In_876,In_944);
or U1070 (N_1070,In_1251,In_674);
nand U1071 (N_1071,In_1293,In_1130);
and U1072 (N_1072,In_2178,In_2399);
or U1073 (N_1073,In_422,In_1208);
and U1074 (N_1074,In_1693,In_126);
and U1075 (N_1075,In_1481,In_387);
and U1076 (N_1076,In_1421,In_1699);
nor U1077 (N_1077,In_1859,In_1381);
nand U1078 (N_1078,In_1679,In_1403);
and U1079 (N_1079,In_1726,In_808);
or U1080 (N_1080,In_1634,In_1604);
or U1081 (N_1081,In_2100,In_1368);
and U1082 (N_1082,In_1810,In_356);
or U1083 (N_1083,In_1817,In_1029);
or U1084 (N_1084,In_1348,In_2482);
nand U1085 (N_1085,In_339,In_836);
nand U1086 (N_1086,In_777,In_961);
xor U1087 (N_1087,In_758,In_2288);
nand U1088 (N_1088,In_365,In_2270);
or U1089 (N_1089,In_1932,In_1991);
nand U1090 (N_1090,In_2212,In_315);
nor U1091 (N_1091,In_1018,In_1247);
nand U1092 (N_1092,In_1330,In_2463);
and U1093 (N_1093,In_2314,In_843);
or U1094 (N_1094,In_468,In_363);
nor U1095 (N_1095,In_2398,In_1767);
or U1096 (N_1096,In_1957,In_1365);
or U1097 (N_1097,In_589,In_281);
nand U1098 (N_1098,In_1643,In_470);
xor U1099 (N_1099,In_1883,In_1374);
or U1100 (N_1100,In_1273,In_1220);
nor U1101 (N_1101,In_975,In_474);
nand U1102 (N_1102,In_2480,In_917);
xor U1103 (N_1103,In_2133,In_761);
nor U1104 (N_1104,In_1868,In_1264);
nand U1105 (N_1105,In_1759,In_1087);
xor U1106 (N_1106,In_1035,In_348);
and U1107 (N_1107,In_2069,In_217);
xor U1108 (N_1108,In_1021,In_1399);
and U1109 (N_1109,In_1484,In_1009);
nor U1110 (N_1110,In_2247,In_173);
nor U1111 (N_1111,In_114,In_1862);
nand U1112 (N_1112,In_1187,In_871);
nor U1113 (N_1113,In_1276,In_1622);
and U1114 (N_1114,In_74,In_316);
nor U1115 (N_1115,In_989,In_1127);
nor U1116 (N_1116,In_1794,In_779);
or U1117 (N_1117,In_2374,In_835);
or U1118 (N_1118,In_1955,In_200);
and U1119 (N_1119,In_52,In_986);
or U1120 (N_1120,In_50,In_243);
xor U1121 (N_1121,In_2397,In_68);
or U1122 (N_1122,In_439,In_635);
and U1123 (N_1123,In_1709,In_1032);
and U1124 (N_1124,In_2065,In_861);
nor U1125 (N_1125,In_1719,In_2294);
xnor U1126 (N_1126,In_262,In_953);
or U1127 (N_1127,In_1995,In_2089);
or U1128 (N_1128,In_2061,In_1074);
nor U1129 (N_1129,In_2002,In_1766);
xnor U1130 (N_1130,In_907,In_1397);
nor U1131 (N_1131,In_1878,In_1244);
nor U1132 (N_1132,In_2223,In_1717);
or U1133 (N_1133,In_1243,In_1322);
or U1134 (N_1134,In_1027,In_2259);
nor U1135 (N_1135,In_1523,In_1771);
or U1136 (N_1136,In_496,In_472);
and U1137 (N_1137,In_1114,In_1177);
or U1138 (N_1138,In_2187,In_494);
or U1139 (N_1139,In_2186,In_670);
nand U1140 (N_1140,In_1728,In_368);
and U1141 (N_1141,In_342,In_1209);
or U1142 (N_1142,In_259,In_1250);
nor U1143 (N_1143,In_872,In_1014);
nor U1144 (N_1144,In_1155,In_2106);
nand U1145 (N_1145,In_721,In_2266);
nand U1146 (N_1146,In_87,In_1212);
nor U1147 (N_1147,In_1472,In_1104);
nand U1148 (N_1148,In_1343,In_1936);
and U1149 (N_1149,In_255,In_692);
and U1150 (N_1150,In_2449,In_755);
and U1151 (N_1151,In_1576,In_702);
xnor U1152 (N_1152,In_300,In_109);
xnor U1153 (N_1153,In_2342,In_1816);
nand U1154 (N_1154,In_153,In_2409);
nand U1155 (N_1155,In_355,In_261);
or U1156 (N_1156,In_1090,In_981);
nand U1157 (N_1157,In_1996,In_731);
nand U1158 (N_1158,In_586,In_1157);
nand U1159 (N_1159,In_607,In_263);
nand U1160 (N_1160,In_647,In_284);
nand U1161 (N_1161,In_967,In_400);
or U1162 (N_1162,In_295,In_1216);
or U1163 (N_1163,In_1171,In_127);
nand U1164 (N_1164,In_128,In_1535);
or U1165 (N_1165,In_2170,In_654);
nand U1166 (N_1166,In_752,In_1189);
and U1167 (N_1167,In_447,In_465);
or U1168 (N_1168,In_977,In_1954);
and U1169 (N_1169,In_1084,In_533);
nand U1170 (N_1170,In_1829,In_24);
nand U1171 (N_1171,In_93,In_1674);
nand U1172 (N_1172,In_2161,In_2159);
nand U1173 (N_1173,In_882,In_2305);
and U1174 (N_1174,In_1442,In_1016);
or U1175 (N_1175,In_600,In_1528);
nor U1176 (N_1176,In_826,In_424);
or U1177 (N_1177,In_53,In_1850);
nand U1178 (N_1178,In_2477,In_1331);
nand U1179 (N_1179,In_2349,In_857);
and U1180 (N_1180,In_2344,In_728);
and U1181 (N_1181,In_397,In_1639);
or U1182 (N_1182,In_1438,In_1723);
and U1183 (N_1183,In_1988,In_457);
or U1184 (N_1184,In_2026,In_1407);
nand U1185 (N_1185,In_1314,In_2205);
or U1186 (N_1186,In_616,In_245);
or U1187 (N_1187,In_1172,In_2316);
nor U1188 (N_1188,In_528,In_1163);
nand U1189 (N_1189,In_26,In_820);
or U1190 (N_1190,In_1577,In_1115);
and U1191 (N_1191,In_1702,In_1449);
nor U1192 (N_1192,In_140,In_2469);
and U1193 (N_1193,In_1748,In_403);
xnor U1194 (N_1194,In_1002,In_660);
xnor U1195 (N_1195,In_141,In_2228);
and U1196 (N_1196,In_1320,In_2039);
nor U1197 (N_1197,In_2192,In_482);
nand U1198 (N_1198,In_837,In_2435);
and U1199 (N_1199,In_2340,In_1282);
or U1200 (N_1200,In_2028,In_1851);
xnor U1201 (N_1201,In_2211,In_2241);
nand U1202 (N_1202,In_391,In_1532);
or U1203 (N_1203,In_792,In_135);
nor U1204 (N_1204,In_2313,In_2057);
nor U1205 (N_1205,In_297,In_499);
nor U1206 (N_1206,In_570,In_966);
xnor U1207 (N_1207,In_886,In_644);
nor U1208 (N_1208,In_1641,In_1043);
or U1209 (N_1209,In_1433,In_1303);
and U1210 (N_1210,In_2473,In_409);
and U1211 (N_1211,In_1692,In_373);
or U1212 (N_1212,In_252,In_2053);
or U1213 (N_1213,In_488,In_1036);
and U1214 (N_1214,In_1582,In_1628);
or U1215 (N_1215,In_1031,In_1938);
or U1216 (N_1216,In_2269,In_537);
nand U1217 (N_1217,In_167,In_1437);
nand U1218 (N_1218,In_2308,In_1237);
and U1219 (N_1219,In_371,In_451);
nor U1220 (N_1220,In_260,In_2232);
nor U1221 (N_1221,In_205,In_89);
and U1222 (N_1222,In_441,In_744);
and U1223 (N_1223,In_911,In_2121);
nor U1224 (N_1224,In_2484,In_1510);
and U1225 (N_1225,In_1389,In_2233);
nand U1226 (N_1226,In_2464,In_2319);
nor U1227 (N_1227,In_733,In_481);
nor U1228 (N_1228,In_985,In_1440);
nand U1229 (N_1229,In_23,In_1423);
nand U1230 (N_1230,In_1256,In_984);
nor U1231 (N_1231,In_1506,In_1464);
nor U1232 (N_1232,In_643,In_980);
nor U1233 (N_1233,In_1512,In_1888);
nand U1234 (N_1234,In_2402,In_1997);
and U1235 (N_1235,In_1462,In_679);
and U1236 (N_1236,In_2472,In_97);
nand U1237 (N_1237,In_2497,In_1144);
xnor U1238 (N_1238,In_489,In_2235);
nor U1239 (N_1239,In_1917,In_2181);
or U1240 (N_1240,In_1372,In_58);
nor U1241 (N_1241,In_80,In_912);
nor U1242 (N_1242,In_960,In_862);
nor U1243 (N_1243,In_359,In_2144);
or U1244 (N_1244,In_815,In_106);
nor U1245 (N_1245,In_367,In_103);
xor U1246 (N_1246,In_2030,In_225);
nor U1247 (N_1247,In_1575,In_1732);
xor U1248 (N_1248,In_354,In_1790);
nand U1249 (N_1249,In_1345,In_1044);
nor U1250 (N_1250,In_273,In_820);
nor U1251 (N_1251,In_1145,In_812);
or U1252 (N_1252,In_1301,In_1302);
nand U1253 (N_1253,In_1513,In_2343);
and U1254 (N_1254,In_1699,In_2105);
nand U1255 (N_1255,In_281,In_2287);
and U1256 (N_1256,In_2219,In_1514);
nand U1257 (N_1257,In_1693,In_648);
or U1258 (N_1258,In_83,In_2177);
and U1259 (N_1259,In_117,In_524);
or U1260 (N_1260,In_1262,In_1781);
and U1261 (N_1261,In_867,In_1796);
and U1262 (N_1262,In_19,In_1626);
or U1263 (N_1263,In_1012,In_1329);
and U1264 (N_1264,In_1092,In_360);
nor U1265 (N_1265,In_856,In_2488);
and U1266 (N_1266,In_810,In_2124);
and U1267 (N_1267,In_2006,In_1093);
and U1268 (N_1268,In_2424,In_1875);
nand U1269 (N_1269,In_885,In_907);
nor U1270 (N_1270,In_1632,In_543);
xor U1271 (N_1271,In_730,In_839);
nor U1272 (N_1272,In_1291,In_622);
and U1273 (N_1273,In_477,In_1394);
nor U1274 (N_1274,In_868,In_2056);
nand U1275 (N_1275,In_705,In_732);
and U1276 (N_1276,In_1718,In_538);
or U1277 (N_1277,In_486,In_1132);
or U1278 (N_1278,In_499,In_508);
or U1279 (N_1279,In_240,In_1003);
nand U1280 (N_1280,In_1172,In_2400);
nand U1281 (N_1281,In_232,In_1669);
nand U1282 (N_1282,In_1527,In_958);
xor U1283 (N_1283,In_1692,In_636);
nand U1284 (N_1284,In_1201,In_421);
and U1285 (N_1285,In_2126,In_923);
and U1286 (N_1286,In_1487,In_235);
nand U1287 (N_1287,In_242,In_198);
or U1288 (N_1288,In_2433,In_1812);
and U1289 (N_1289,In_1304,In_1754);
or U1290 (N_1290,In_2200,In_862);
and U1291 (N_1291,In_519,In_1830);
xor U1292 (N_1292,In_1751,In_1251);
nand U1293 (N_1293,In_2239,In_1628);
nand U1294 (N_1294,In_1363,In_1280);
nor U1295 (N_1295,In_958,In_2334);
nand U1296 (N_1296,In_1861,In_1198);
nand U1297 (N_1297,In_1248,In_199);
and U1298 (N_1298,In_1072,In_2071);
nor U1299 (N_1299,In_1643,In_500);
nor U1300 (N_1300,In_804,In_254);
and U1301 (N_1301,In_1823,In_1025);
xor U1302 (N_1302,In_191,In_2079);
nor U1303 (N_1303,In_299,In_77);
and U1304 (N_1304,In_171,In_1954);
or U1305 (N_1305,In_1736,In_74);
nand U1306 (N_1306,In_131,In_796);
or U1307 (N_1307,In_1968,In_98);
nand U1308 (N_1308,In_1930,In_2064);
nor U1309 (N_1309,In_1255,In_1390);
or U1310 (N_1310,In_2270,In_800);
nor U1311 (N_1311,In_476,In_2273);
or U1312 (N_1312,In_708,In_3);
nand U1313 (N_1313,In_1539,In_2109);
nand U1314 (N_1314,In_775,In_1307);
or U1315 (N_1315,In_708,In_1589);
nand U1316 (N_1316,In_2128,In_2302);
and U1317 (N_1317,In_75,In_701);
nor U1318 (N_1318,In_347,In_482);
and U1319 (N_1319,In_1438,In_1133);
nand U1320 (N_1320,In_594,In_2445);
nand U1321 (N_1321,In_553,In_1869);
nor U1322 (N_1322,In_47,In_1);
or U1323 (N_1323,In_1812,In_2291);
xor U1324 (N_1324,In_2342,In_1573);
nor U1325 (N_1325,In_2159,In_1428);
and U1326 (N_1326,In_314,In_955);
nand U1327 (N_1327,In_1336,In_824);
and U1328 (N_1328,In_1236,In_2177);
or U1329 (N_1329,In_802,In_1100);
or U1330 (N_1330,In_1875,In_834);
and U1331 (N_1331,In_64,In_2276);
or U1332 (N_1332,In_722,In_439);
nand U1333 (N_1333,In_1840,In_1339);
and U1334 (N_1334,In_192,In_2160);
or U1335 (N_1335,In_78,In_420);
nor U1336 (N_1336,In_168,In_2223);
nor U1337 (N_1337,In_1733,In_1597);
nor U1338 (N_1338,In_802,In_2369);
or U1339 (N_1339,In_1008,In_1731);
nand U1340 (N_1340,In_2250,In_647);
xnor U1341 (N_1341,In_647,In_694);
and U1342 (N_1342,In_852,In_2362);
and U1343 (N_1343,In_57,In_423);
nand U1344 (N_1344,In_686,In_746);
nor U1345 (N_1345,In_1217,In_1230);
nor U1346 (N_1346,In_370,In_1403);
nand U1347 (N_1347,In_1753,In_1311);
or U1348 (N_1348,In_1494,In_695);
nor U1349 (N_1349,In_1711,In_1567);
or U1350 (N_1350,In_39,In_2014);
nand U1351 (N_1351,In_1527,In_2315);
or U1352 (N_1352,In_291,In_2468);
nor U1353 (N_1353,In_1711,In_2322);
and U1354 (N_1354,In_79,In_1921);
nand U1355 (N_1355,In_1638,In_656);
or U1356 (N_1356,In_1518,In_752);
and U1357 (N_1357,In_771,In_1399);
and U1358 (N_1358,In_1588,In_1845);
or U1359 (N_1359,In_1047,In_2135);
nor U1360 (N_1360,In_989,In_1255);
and U1361 (N_1361,In_93,In_1860);
or U1362 (N_1362,In_1363,In_798);
nand U1363 (N_1363,In_774,In_1165);
and U1364 (N_1364,In_1484,In_2481);
nand U1365 (N_1365,In_227,In_550);
nor U1366 (N_1366,In_1012,In_488);
xor U1367 (N_1367,In_1973,In_1122);
nor U1368 (N_1368,In_273,In_6);
or U1369 (N_1369,In_1092,In_1492);
or U1370 (N_1370,In_307,In_1374);
nand U1371 (N_1371,In_1097,In_1791);
and U1372 (N_1372,In_674,In_1609);
nand U1373 (N_1373,In_1516,In_1435);
nor U1374 (N_1374,In_930,In_2218);
and U1375 (N_1375,In_1314,In_2380);
or U1376 (N_1376,In_1038,In_1315);
xor U1377 (N_1377,In_746,In_839);
xnor U1378 (N_1378,In_857,In_2218);
and U1379 (N_1379,In_501,In_745);
and U1380 (N_1380,In_812,In_689);
nand U1381 (N_1381,In_2035,In_2140);
nand U1382 (N_1382,In_1867,In_790);
nor U1383 (N_1383,In_1783,In_551);
and U1384 (N_1384,In_2240,In_693);
and U1385 (N_1385,In_1541,In_1315);
or U1386 (N_1386,In_754,In_179);
and U1387 (N_1387,In_918,In_651);
xor U1388 (N_1388,In_1830,In_267);
xnor U1389 (N_1389,In_1102,In_1286);
nand U1390 (N_1390,In_1293,In_469);
and U1391 (N_1391,In_628,In_1788);
xnor U1392 (N_1392,In_501,In_682);
nor U1393 (N_1393,In_1929,In_418);
and U1394 (N_1394,In_1666,In_1773);
or U1395 (N_1395,In_2008,In_1107);
or U1396 (N_1396,In_1722,In_2463);
nand U1397 (N_1397,In_524,In_1531);
nand U1398 (N_1398,In_1248,In_2220);
xor U1399 (N_1399,In_1819,In_516);
and U1400 (N_1400,In_1548,In_1915);
nor U1401 (N_1401,In_2222,In_1929);
nand U1402 (N_1402,In_2135,In_2242);
nor U1403 (N_1403,In_1292,In_348);
nand U1404 (N_1404,In_2188,In_1960);
and U1405 (N_1405,In_1827,In_1913);
and U1406 (N_1406,In_1592,In_2238);
nand U1407 (N_1407,In_1093,In_854);
nor U1408 (N_1408,In_321,In_1582);
or U1409 (N_1409,In_1793,In_1696);
nand U1410 (N_1410,In_2294,In_86);
and U1411 (N_1411,In_1486,In_1731);
xnor U1412 (N_1412,In_528,In_508);
or U1413 (N_1413,In_787,In_938);
nor U1414 (N_1414,In_1551,In_2157);
or U1415 (N_1415,In_2433,In_1050);
and U1416 (N_1416,In_2318,In_1458);
nor U1417 (N_1417,In_2369,In_2187);
nor U1418 (N_1418,In_313,In_185);
nor U1419 (N_1419,In_1968,In_1852);
nand U1420 (N_1420,In_599,In_807);
nor U1421 (N_1421,In_1233,In_409);
or U1422 (N_1422,In_1516,In_309);
or U1423 (N_1423,In_17,In_1458);
and U1424 (N_1424,In_707,In_825);
nor U1425 (N_1425,In_539,In_2367);
nor U1426 (N_1426,In_228,In_2314);
nor U1427 (N_1427,In_342,In_1245);
nand U1428 (N_1428,In_1329,In_2418);
or U1429 (N_1429,In_1109,In_860);
and U1430 (N_1430,In_189,In_930);
nor U1431 (N_1431,In_948,In_1147);
or U1432 (N_1432,In_1372,In_2478);
or U1433 (N_1433,In_1528,In_859);
and U1434 (N_1434,In_188,In_450);
or U1435 (N_1435,In_1365,In_2301);
or U1436 (N_1436,In_200,In_784);
and U1437 (N_1437,In_2246,In_1322);
nand U1438 (N_1438,In_1770,In_2065);
nand U1439 (N_1439,In_293,In_1079);
nor U1440 (N_1440,In_1978,In_208);
and U1441 (N_1441,In_2419,In_1539);
and U1442 (N_1442,In_1392,In_39);
and U1443 (N_1443,In_982,In_2136);
or U1444 (N_1444,In_828,In_33);
xnor U1445 (N_1445,In_103,In_79);
and U1446 (N_1446,In_1966,In_1300);
nor U1447 (N_1447,In_2225,In_1833);
nor U1448 (N_1448,In_2239,In_618);
xor U1449 (N_1449,In_2423,In_17);
nand U1450 (N_1450,In_34,In_1171);
xnor U1451 (N_1451,In_2122,In_1095);
nor U1452 (N_1452,In_2239,In_2336);
xnor U1453 (N_1453,In_90,In_785);
nand U1454 (N_1454,In_175,In_2193);
nand U1455 (N_1455,In_339,In_484);
nand U1456 (N_1456,In_822,In_150);
or U1457 (N_1457,In_1802,In_396);
xnor U1458 (N_1458,In_2310,In_1827);
and U1459 (N_1459,In_1173,In_730);
and U1460 (N_1460,In_1405,In_420);
and U1461 (N_1461,In_748,In_808);
and U1462 (N_1462,In_1221,In_1198);
nor U1463 (N_1463,In_1513,In_379);
nor U1464 (N_1464,In_516,In_56);
nand U1465 (N_1465,In_1880,In_483);
nor U1466 (N_1466,In_646,In_1052);
nor U1467 (N_1467,In_1875,In_807);
xnor U1468 (N_1468,In_2426,In_1708);
nor U1469 (N_1469,In_851,In_748);
or U1470 (N_1470,In_203,In_463);
or U1471 (N_1471,In_1621,In_2427);
nor U1472 (N_1472,In_195,In_82);
and U1473 (N_1473,In_2276,In_746);
and U1474 (N_1474,In_1097,In_588);
or U1475 (N_1475,In_284,In_1520);
and U1476 (N_1476,In_482,In_1210);
and U1477 (N_1477,In_276,In_12);
nor U1478 (N_1478,In_792,In_1708);
nand U1479 (N_1479,In_2054,In_2185);
nor U1480 (N_1480,In_2148,In_1373);
and U1481 (N_1481,In_7,In_1496);
nand U1482 (N_1482,In_1846,In_1383);
nand U1483 (N_1483,In_1286,In_1033);
and U1484 (N_1484,In_1942,In_1088);
nand U1485 (N_1485,In_1734,In_1598);
and U1486 (N_1486,In_1847,In_314);
and U1487 (N_1487,In_1004,In_1479);
and U1488 (N_1488,In_1064,In_630);
and U1489 (N_1489,In_796,In_1355);
nor U1490 (N_1490,In_2097,In_1359);
or U1491 (N_1491,In_1295,In_1700);
or U1492 (N_1492,In_2441,In_736);
nand U1493 (N_1493,In_65,In_1689);
and U1494 (N_1494,In_621,In_51);
or U1495 (N_1495,In_460,In_1975);
nor U1496 (N_1496,In_172,In_1495);
and U1497 (N_1497,In_779,In_2147);
or U1498 (N_1498,In_707,In_130);
nand U1499 (N_1499,In_870,In_540);
or U1500 (N_1500,In_459,In_1271);
and U1501 (N_1501,In_1634,In_1325);
xnor U1502 (N_1502,In_772,In_2052);
and U1503 (N_1503,In_1923,In_127);
or U1504 (N_1504,In_614,In_900);
or U1505 (N_1505,In_359,In_1047);
xnor U1506 (N_1506,In_2339,In_586);
xor U1507 (N_1507,In_1393,In_312);
nand U1508 (N_1508,In_1054,In_2268);
and U1509 (N_1509,In_988,In_1360);
and U1510 (N_1510,In_2247,In_2059);
or U1511 (N_1511,In_240,In_136);
nand U1512 (N_1512,In_160,In_1064);
and U1513 (N_1513,In_1707,In_1391);
nand U1514 (N_1514,In_2310,In_284);
or U1515 (N_1515,In_1121,In_591);
or U1516 (N_1516,In_470,In_1431);
or U1517 (N_1517,In_53,In_1939);
and U1518 (N_1518,In_233,In_501);
nor U1519 (N_1519,In_172,In_758);
nor U1520 (N_1520,In_644,In_384);
nor U1521 (N_1521,In_989,In_357);
nor U1522 (N_1522,In_2036,In_1511);
or U1523 (N_1523,In_801,In_890);
or U1524 (N_1524,In_448,In_1133);
and U1525 (N_1525,In_2276,In_358);
nor U1526 (N_1526,In_889,In_1110);
xnor U1527 (N_1527,In_1927,In_2008);
nor U1528 (N_1528,In_252,In_708);
and U1529 (N_1529,In_1273,In_643);
nand U1530 (N_1530,In_2324,In_406);
nor U1531 (N_1531,In_1159,In_1053);
nor U1532 (N_1532,In_1987,In_379);
or U1533 (N_1533,In_532,In_860);
nand U1534 (N_1534,In_401,In_116);
and U1535 (N_1535,In_712,In_1515);
xnor U1536 (N_1536,In_1684,In_1088);
or U1537 (N_1537,In_1231,In_1927);
nand U1538 (N_1538,In_381,In_463);
or U1539 (N_1539,In_1759,In_215);
and U1540 (N_1540,In_1861,In_1786);
nand U1541 (N_1541,In_1964,In_224);
or U1542 (N_1542,In_264,In_344);
nand U1543 (N_1543,In_388,In_1199);
nand U1544 (N_1544,In_2131,In_2346);
xnor U1545 (N_1545,In_653,In_847);
nand U1546 (N_1546,In_700,In_1275);
xnor U1547 (N_1547,In_1714,In_2361);
or U1548 (N_1548,In_967,In_683);
and U1549 (N_1549,In_1665,In_446);
nor U1550 (N_1550,In_496,In_701);
xor U1551 (N_1551,In_2147,In_121);
nand U1552 (N_1552,In_940,In_761);
nor U1553 (N_1553,In_1725,In_1330);
nor U1554 (N_1554,In_2154,In_368);
nand U1555 (N_1555,In_2292,In_1856);
nor U1556 (N_1556,In_769,In_225);
or U1557 (N_1557,In_985,In_2071);
and U1558 (N_1558,In_1187,In_229);
nand U1559 (N_1559,In_456,In_446);
xnor U1560 (N_1560,In_520,In_1931);
nor U1561 (N_1561,In_1103,In_2116);
nor U1562 (N_1562,In_2168,In_733);
nor U1563 (N_1563,In_1205,In_1458);
nand U1564 (N_1564,In_2333,In_1014);
nand U1565 (N_1565,In_1597,In_1627);
or U1566 (N_1566,In_2413,In_841);
nor U1567 (N_1567,In_1746,In_1902);
or U1568 (N_1568,In_1530,In_2326);
or U1569 (N_1569,In_651,In_1624);
nor U1570 (N_1570,In_800,In_2283);
xor U1571 (N_1571,In_1576,In_217);
nor U1572 (N_1572,In_454,In_121);
nand U1573 (N_1573,In_329,In_477);
and U1574 (N_1574,In_2292,In_732);
and U1575 (N_1575,In_816,In_2094);
nand U1576 (N_1576,In_1882,In_1215);
and U1577 (N_1577,In_1769,In_1068);
xnor U1578 (N_1578,In_1725,In_2450);
nor U1579 (N_1579,In_370,In_1669);
xor U1580 (N_1580,In_1253,In_708);
nor U1581 (N_1581,In_787,In_1717);
or U1582 (N_1582,In_566,In_1451);
nand U1583 (N_1583,In_1207,In_353);
and U1584 (N_1584,In_250,In_1370);
nand U1585 (N_1585,In_479,In_301);
nand U1586 (N_1586,In_991,In_592);
xnor U1587 (N_1587,In_1875,In_1197);
nor U1588 (N_1588,In_2239,In_2219);
and U1589 (N_1589,In_68,In_1766);
or U1590 (N_1590,In_924,In_1705);
nor U1591 (N_1591,In_1038,In_875);
nand U1592 (N_1592,In_1634,In_2061);
nor U1593 (N_1593,In_2047,In_1432);
nand U1594 (N_1594,In_930,In_76);
nand U1595 (N_1595,In_1759,In_2156);
nor U1596 (N_1596,In_1324,In_1138);
nor U1597 (N_1597,In_1708,In_396);
and U1598 (N_1598,In_1236,In_2082);
and U1599 (N_1599,In_65,In_1549);
or U1600 (N_1600,In_1559,In_737);
or U1601 (N_1601,In_665,In_1879);
and U1602 (N_1602,In_1531,In_966);
nand U1603 (N_1603,In_828,In_856);
nand U1604 (N_1604,In_665,In_1981);
xnor U1605 (N_1605,In_1104,In_469);
nand U1606 (N_1606,In_864,In_881);
and U1607 (N_1607,In_837,In_1061);
and U1608 (N_1608,In_2253,In_2367);
nor U1609 (N_1609,In_2339,In_589);
or U1610 (N_1610,In_239,In_695);
or U1611 (N_1611,In_1999,In_1369);
and U1612 (N_1612,In_2201,In_849);
and U1613 (N_1613,In_90,In_915);
nor U1614 (N_1614,In_2457,In_731);
or U1615 (N_1615,In_2257,In_2419);
nor U1616 (N_1616,In_1926,In_203);
nor U1617 (N_1617,In_1747,In_1938);
and U1618 (N_1618,In_1628,In_1253);
and U1619 (N_1619,In_1434,In_1530);
and U1620 (N_1620,In_2063,In_143);
and U1621 (N_1621,In_1508,In_2099);
nand U1622 (N_1622,In_2160,In_586);
nand U1623 (N_1623,In_1453,In_328);
nor U1624 (N_1624,In_2154,In_2063);
xnor U1625 (N_1625,In_2077,In_1311);
nor U1626 (N_1626,In_364,In_1277);
nand U1627 (N_1627,In_1569,In_960);
nor U1628 (N_1628,In_2041,In_991);
and U1629 (N_1629,In_1953,In_43);
nand U1630 (N_1630,In_1826,In_407);
nand U1631 (N_1631,In_1301,In_2039);
or U1632 (N_1632,In_2357,In_1195);
or U1633 (N_1633,In_1578,In_1043);
nor U1634 (N_1634,In_1247,In_291);
and U1635 (N_1635,In_1743,In_523);
xnor U1636 (N_1636,In_1445,In_1196);
xor U1637 (N_1637,In_1491,In_1920);
nor U1638 (N_1638,In_1335,In_2324);
and U1639 (N_1639,In_851,In_2119);
or U1640 (N_1640,In_332,In_1575);
or U1641 (N_1641,In_1553,In_293);
or U1642 (N_1642,In_1676,In_949);
xor U1643 (N_1643,In_2388,In_1924);
nor U1644 (N_1644,In_779,In_503);
nor U1645 (N_1645,In_512,In_1666);
nand U1646 (N_1646,In_1933,In_1759);
or U1647 (N_1647,In_854,In_1044);
nor U1648 (N_1648,In_1193,In_1835);
and U1649 (N_1649,In_1224,In_1504);
nor U1650 (N_1650,In_2484,In_2181);
or U1651 (N_1651,In_1285,In_1789);
nand U1652 (N_1652,In_2149,In_1255);
and U1653 (N_1653,In_1451,In_1842);
or U1654 (N_1654,In_694,In_250);
nor U1655 (N_1655,In_223,In_2401);
nor U1656 (N_1656,In_1080,In_2469);
nor U1657 (N_1657,In_231,In_1226);
and U1658 (N_1658,In_2112,In_2200);
and U1659 (N_1659,In_1428,In_1648);
or U1660 (N_1660,In_2065,In_1399);
nand U1661 (N_1661,In_1467,In_1135);
xor U1662 (N_1662,In_140,In_1293);
and U1663 (N_1663,In_1681,In_1447);
nor U1664 (N_1664,In_1176,In_114);
or U1665 (N_1665,In_222,In_1905);
and U1666 (N_1666,In_2,In_1214);
and U1667 (N_1667,In_2127,In_290);
and U1668 (N_1668,In_1150,In_1441);
nor U1669 (N_1669,In_1842,In_1058);
or U1670 (N_1670,In_787,In_1230);
nand U1671 (N_1671,In_286,In_1472);
and U1672 (N_1672,In_525,In_1468);
nand U1673 (N_1673,In_1758,In_2433);
and U1674 (N_1674,In_566,In_1041);
or U1675 (N_1675,In_496,In_290);
nand U1676 (N_1676,In_2483,In_690);
or U1677 (N_1677,In_2263,In_1863);
or U1678 (N_1678,In_2151,In_967);
nand U1679 (N_1679,In_561,In_1401);
and U1680 (N_1680,In_531,In_207);
or U1681 (N_1681,In_2165,In_224);
or U1682 (N_1682,In_169,In_1204);
and U1683 (N_1683,In_98,In_1460);
nor U1684 (N_1684,In_1894,In_71);
and U1685 (N_1685,In_2249,In_330);
and U1686 (N_1686,In_1304,In_457);
or U1687 (N_1687,In_811,In_1297);
nand U1688 (N_1688,In_785,In_1526);
nand U1689 (N_1689,In_94,In_1409);
nor U1690 (N_1690,In_326,In_2488);
nand U1691 (N_1691,In_2474,In_1655);
nor U1692 (N_1692,In_873,In_2214);
or U1693 (N_1693,In_2285,In_1929);
or U1694 (N_1694,In_1348,In_32);
or U1695 (N_1695,In_60,In_540);
or U1696 (N_1696,In_1078,In_53);
and U1697 (N_1697,In_1119,In_957);
and U1698 (N_1698,In_328,In_1520);
and U1699 (N_1699,In_1685,In_659);
and U1700 (N_1700,In_383,In_2451);
nor U1701 (N_1701,In_1123,In_747);
and U1702 (N_1702,In_396,In_2217);
nor U1703 (N_1703,In_1202,In_1410);
nor U1704 (N_1704,In_1553,In_1246);
nor U1705 (N_1705,In_2485,In_268);
nor U1706 (N_1706,In_2357,In_1546);
nor U1707 (N_1707,In_198,In_2254);
and U1708 (N_1708,In_1823,In_2090);
nor U1709 (N_1709,In_2123,In_1048);
xnor U1710 (N_1710,In_1075,In_1009);
and U1711 (N_1711,In_1850,In_2229);
nor U1712 (N_1712,In_588,In_176);
or U1713 (N_1713,In_1970,In_1623);
or U1714 (N_1714,In_2173,In_1176);
nor U1715 (N_1715,In_1943,In_1066);
and U1716 (N_1716,In_1746,In_906);
and U1717 (N_1717,In_2320,In_509);
and U1718 (N_1718,In_617,In_1535);
or U1719 (N_1719,In_1306,In_340);
or U1720 (N_1720,In_1300,In_2336);
nor U1721 (N_1721,In_2399,In_229);
and U1722 (N_1722,In_403,In_1124);
or U1723 (N_1723,In_926,In_768);
or U1724 (N_1724,In_1293,In_1347);
nor U1725 (N_1725,In_665,In_1674);
and U1726 (N_1726,In_185,In_2074);
and U1727 (N_1727,In_2356,In_945);
and U1728 (N_1728,In_220,In_687);
xor U1729 (N_1729,In_2028,In_1460);
nor U1730 (N_1730,In_692,In_2403);
nand U1731 (N_1731,In_1996,In_2083);
and U1732 (N_1732,In_686,In_1258);
nand U1733 (N_1733,In_302,In_1163);
and U1734 (N_1734,In_2110,In_875);
xor U1735 (N_1735,In_1126,In_1988);
nor U1736 (N_1736,In_1293,In_1860);
and U1737 (N_1737,In_1953,In_1505);
nor U1738 (N_1738,In_1201,In_1810);
nand U1739 (N_1739,In_635,In_1375);
and U1740 (N_1740,In_2252,In_861);
nor U1741 (N_1741,In_2036,In_223);
xor U1742 (N_1742,In_1831,In_2326);
and U1743 (N_1743,In_2035,In_551);
nand U1744 (N_1744,In_631,In_432);
nand U1745 (N_1745,In_2170,In_646);
xnor U1746 (N_1746,In_2431,In_2181);
nand U1747 (N_1747,In_2167,In_333);
nand U1748 (N_1748,In_1010,In_1011);
nand U1749 (N_1749,In_79,In_662);
and U1750 (N_1750,In_826,In_1811);
or U1751 (N_1751,In_1211,In_1946);
or U1752 (N_1752,In_1010,In_451);
nor U1753 (N_1753,In_192,In_1803);
and U1754 (N_1754,In_362,In_2339);
or U1755 (N_1755,In_1849,In_51);
or U1756 (N_1756,In_557,In_1462);
and U1757 (N_1757,In_2414,In_1172);
and U1758 (N_1758,In_1132,In_323);
and U1759 (N_1759,In_520,In_2401);
nand U1760 (N_1760,In_2431,In_461);
nand U1761 (N_1761,In_1002,In_1835);
or U1762 (N_1762,In_2273,In_556);
and U1763 (N_1763,In_2423,In_2225);
or U1764 (N_1764,In_2408,In_170);
or U1765 (N_1765,In_1664,In_229);
nor U1766 (N_1766,In_391,In_418);
nand U1767 (N_1767,In_1400,In_1784);
and U1768 (N_1768,In_1965,In_2203);
or U1769 (N_1769,In_590,In_1440);
nand U1770 (N_1770,In_1061,In_2366);
and U1771 (N_1771,In_2246,In_426);
and U1772 (N_1772,In_1321,In_171);
or U1773 (N_1773,In_1400,In_1310);
nand U1774 (N_1774,In_778,In_1117);
nand U1775 (N_1775,In_66,In_968);
or U1776 (N_1776,In_2003,In_1414);
nor U1777 (N_1777,In_1920,In_1532);
and U1778 (N_1778,In_1637,In_2383);
nand U1779 (N_1779,In_893,In_1145);
or U1780 (N_1780,In_1547,In_2492);
and U1781 (N_1781,In_2130,In_347);
xnor U1782 (N_1782,In_2178,In_921);
nand U1783 (N_1783,In_1956,In_2369);
and U1784 (N_1784,In_636,In_502);
nand U1785 (N_1785,In_2144,In_2376);
or U1786 (N_1786,In_2280,In_1439);
or U1787 (N_1787,In_229,In_2372);
nor U1788 (N_1788,In_693,In_821);
nand U1789 (N_1789,In_2360,In_1025);
or U1790 (N_1790,In_263,In_1649);
nand U1791 (N_1791,In_1748,In_1991);
nand U1792 (N_1792,In_2298,In_1282);
or U1793 (N_1793,In_722,In_409);
nor U1794 (N_1794,In_1129,In_681);
nand U1795 (N_1795,In_556,In_645);
or U1796 (N_1796,In_1664,In_2193);
and U1797 (N_1797,In_1142,In_2197);
nand U1798 (N_1798,In_1268,In_2253);
nand U1799 (N_1799,In_753,In_374);
or U1800 (N_1800,In_2269,In_644);
nand U1801 (N_1801,In_2043,In_740);
xor U1802 (N_1802,In_2409,In_1819);
and U1803 (N_1803,In_1000,In_980);
or U1804 (N_1804,In_2476,In_564);
nand U1805 (N_1805,In_2175,In_791);
or U1806 (N_1806,In_864,In_260);
or U1807 (N_1807,In_625,In_1167);
xnor U1808 (N_1808,In_2330,In_1728);
and U1809 (N_1809,In_1696,In_61);
and U1810 (N_1810,In_447,In_1070);
nor U1811 (N_1811,In_1383,In_2499);
nand U1812 (N_1812,In_1047,In_165);
and U1813 (N_1813,In_1625,In_1450);
nor U1814 (N_1814,In_1193,In_320);
nor U1815 (N_1815,In_419,In_1643);
nor U1816 (N_1816,In_759,In_2272);
nand U1817 (N_1817,In_1370,In_962);
and U1818 (N_1818,In_479,In_2261);
or U1819 (N_1819,In_1291,In_9);
or U1820 (N_1820,In_769,In_2148);
nor U1821 (N_1821,In_1009,In_1277);
nand U1822 (N_1822,In_1232,In_21);
xnor U1823 (N_1823,In_565,In_1807);
nor U1824 (N_1824,In_2477,In_1089);
nor U1825 (N_1825,In_1653,In_504);
nor U1826 (N_1826,In_2496,In_172);
and U1827 (N_1827,In_392,In_70);
nor U1828 (N_1828,In_1285,In_1185);
and U1829 (N_1829,In_1127,In_642);
nand U1830 (N_1830,In_304,In_2433);
nor U1831 (N_1831,In_39,In_1065);
nand U1832 (N_1832,In_825,In_1227);
xor U1833 (N_1833,In_2222,In_760);
or U1834 (N_1834,In_1581,In_1304);
xnor U1835 (N_1835,In_242,In_1597);
or U1836 (N_1836,In_2035,In_1166);
and U1837 (N_1837,In_872,In_1586);
xor U1838 (N_1838,In_1498,In_440);
nand U1839 (N_1839,In_905,In_369);
nor U1840 (N_1840,In_716,In_601);
nor U1841 (N_1841,In_402,In_2361);
nor U1842 (N_1842,In_1557,In_2097);
xnor U1843 (N_1843,In_704,In_1003);
nand U1844 (N_1844,In_1680,In_999);
and U1845 (N_1845,In_105,In_17);
nor U1846 (N_1846,In_1719,In_1486);
and U1847 (N_1847,In_658,In_239);
xor U1848 (N_1848,In_84,In_1168);
and U1849 (N_1849,In_883,In_1662);
or U1850 (N_1850,In_729,In_1337);
and U1851 (N_1851,In_2396,In_179);
or U1852 (N_1852,In_2227,In_1103);
or U1853 (N_1853,In_47,In_25);
nor U1854 (N_1854,In_1651,In_338);
or U1855 (N_1855,In_2030,In_1516);
or U1856 (N_1856,In_1677,In_1321);
nor U1857 (N_1857,In_1584,In_2482);
nand U1858 (N_1858,In_35,In_2171);
nand U1859 (N_1859,In_493,In_134);
or U1860 (N_1860,In_884,In_1266);
nor U1861 (N_1861,In_149,In_940);
nand U1862 (N_1862,In_117,In_422);
and U1863 (N_1863,In_1501,In_1678);
and U1864 (N_1864,In_1634,In_1842);
nand U1865 (N_1865,In_692,In_1675);
nand U1866 (N_1866,In_1173,In_443);
nand U1867 (N_1867,In_113,In_2352);
or U1868 (N_1868,In_808,In_1314);
and U1869 (N_1869,In_1556,In_121);
nor U1870 (N_1870,In_1732,In_1679);
and U1871 (N_1871,In_459,In_651);
xor U1872 (N_1872,In_2326,In_363);
nor U1873 (N_1873,In_1195,In_450);
nor U1874 (N_1874,In_1214,In_975);
and U1875 (N_1875,In_1014,In_1835);
and U1876 (N_1876,In_374,In_2236);
nand U1877 (N_1877,In_1571,In_576);
or U1878 (N_1878,In_359,In_2469);
or U1879 (N_1879,In_1453,In_988);
or U1880 (N_1880,In_1177,In_2063);
or U1881 (N_1881,In_408,In_1811);
or U1882 (N_1882,In_728,In_1916);
and U1883 (N_1883,In_431,In_2335);
or U1884 (N_1884,In_2029,In_1174);
and U1885 (N_1885,In_1537,In_1575);
nand U1886 (N_1886,In_1004,In_1733);
nor U1887 (N_1887,In_565,In_1028);
nand U1888 (N_1888,In_2232,In_984);
or U1889 (N_1889,In_955,In_1757);
or U1890 (N_1890,In_85,In_2419);
nand U1891 (N_1891,In_1679,In_1468);
or U1892 (N_1892,In_888,In_2230);
nand U1893 (N_1893,In_111,In_2029);
and U1894 (N_1894,In_1278,In_679);
or U1895 (N_1895,In_958,In_782);
nand U1896 (N_1896,In_1699,In_221);
nor U1897 (N_1897,In_2368,In_267);
xnor U1898 (N_1898,In_229,In_505);
or U1899 (N_1899,In_213,In_1688);
nor U1900 (N_1900,In_163,In_211);
xor U1901 (N_1901,In_2084,In_2224);
or U1902 (N_1902,In_900,In_2210);
nand U1903 (N_1903,In_1356,In_610);
nand U1904 (N_1904,In_2481,In_1634);
nor U1905 (N_1905,In_1726,In_2263);
nand U1906 (N_1906,In_1540,In_544);
xnor U1907 (N_1907,In_1743,In_1456);
nor U1908 (N_1908,In_1786,In_42);
nor U1909 (N_1909,In_2143,In_938);
xor U1910 (N_1910,In_2430,In_477);
and U1911 (N_1911,In_1446,In_1514);
or U1912 (N_1912,In_461,In_2194);
nand U1913 (N_1913,In_1591,In_786);
and U1914 (N_1914,In_465,In_1631);
nor U1915 (N_1915,In_1670,In_1330);
or U1916 (N_1916,In_30,In_742);
nor U1917 (N_1917,In_576,In_1730);
or U1918 (N_1918,In_707,In_2376);
or U1919 (N_1919,In_1762,In_1538);
nand U1920 (N_1920,In_1062,In_1158);
nand U1921 (N_1921,In_2328,In_1612);
nand U1922 (N_1922,In_789,In_1348);
nand U1923 (N_1923,In_986,In_1468);
and U1924 (N_1924,In_2045,In_2440);
or U1925 (N_1925,In_1871,In_1229);
and U1926 (N_1926,In_1143,In_664);
and U1927 (N_1927,In_1521,In_995);
or U1928 (N_1928,In_1289,In_370);
or U1929 (N_1929,In_2066,In_1835);
nor U1930 (N_1930,In_556,In_1890);
nor U1931 (N_1931,In_2269,In_1725);
and U1932 (N_1932,In_111,In_473);
xor U1933 (N_1933,In_854,In_1269);
or U1934 (N_1934,In_74,In_2054);
and U1935 (N_1935,In_1363,In_882);
or U1936 (N_1936,In_565,In_103);
nor U1937 (N_1937,In_1595,In_409);
or U1938 (N_1938,In_1711,In_1827);
or U1939 (N_1939,In_348,In_1414);
or U1940 (N_1940,In_946,In_990);
nand U1941 (N_1941,In_631,In_105);
and U1942 (N_1942,In_1670,In_1497);
nor U1943 (N_1943,In_35,In_1247);
and U1944 (N_1944,In_2132,In_2158);
or U1945 (N_1945,In_1645,In_1008);
or U1946 (N_1946,In_2473,In_1724);
xnor U1947 (N_1947,In_1831,In_829);
nand U1948 (N_1948,In_2202,In_2229);
or U1949 (N_1949,In_1566,In_2460);
nand U1950 (N_1950,In_717,In_226);
and U1951 (N_1951,In_1552,In_1586);
nor U1952 (N_1952,In_496,In_2215);
and U1953 (N_1953,In_352,In_2428);
or U1954 (N_1954,In_1547,In_1495);
and U1955 (N_1955,In_1953,In_51);
nor U1956 (N_1956,In_1715,In_1640);
or U1957 (N_1957,In_2049,In_1877);
nand U1958 (N_1958,In_1445,In_1457);
xnor U1959 (N_1959,In_876,In_46);
and U1960 (N_1960,In_407,In_1868);
nand U1961 (N_1961,In_1358,In_1776);
and U1962 (N_1962,In_2290,In_1703);
nor U1963 (N_1963,In_2001,In_658);
or U1964 (N_1964,In_2333,In_1861);
nand U1965 (N_1965,In_2490,In_1081);
and U1966 (N_1966,In_830,In_2014);
or U1967 (N_1967,In_1529,In_2403);
or U1968 (N_1968,In_1889,In_1400);
nand U1969 (N_1969,In_1443,In_1902);
or U1970 (N_1970,In_475,In_555);
and U1971 (N_1971,In_1761,In_2238);
nor U1972 (N_1972,In_1470,In_784);
or U1973 (N_1973,In_2442,In_349);
or U1974 (N_1974,In_872,In_921);
nand U1975 (N_1975,In_28,In_1876);
nor U1976 (N_1976,In_374,In_939);
and U1977 (N_1977,In_1970,In_1261);
xor U1978 (N_1978,In_820,In_1507);
nand U1979 (N_1979,In_681,In_236);
and U1980 (N_1980,In_793,In_1740);
and U1981 (N_1981,In_909,In_539);
and U1982 (N_1982,In_657,In_1976);
xor U1983 (N_1983,In_2387,In_937);
nor U1984 (N_1984,In_2294,In_1753);
nand U1985 (N_1985,In_2040,In_893);
and U1986 (N_1986,In_310,In_393);
nand U1987 (N_1987,In_1587,In_2098);
nor U1988 (N_1988,In_2091,In_1390);
and U1989 (N_1989,In_1107,In_1435);
nor U1990 (N_1990,In_776,In_429);
nor U1991 (N_1991,In_662,In_2128);
and U1992 (N_1992,In_1287,In_2351);
nor U1993 (N_1993,In_954,In_668);
nor U1994 (N_1994,In_1660,In_1311);
and U1995 (N_1995,In_2292,In_327);
xor U1996 (N_1996,In_997,In_926);
nor U1997 (N_1997,In_2309,In_289);
nor U1998 (N_1998,In_1697,In_1039);
nand U1999 (N_1999,In_463,In_834);
nand U2000 (N_2000,In_815,In_1057);
or U2001 (N_2001,In_559,In_142);
nor U2002 (N_2002,In_1785,In_792);
and U2003 (N_2003,In_1583,In_303);
and U2004 (N_2004,In_2117,In_875);
and U2005 (N_2005,In_2211,In_1653);
nor U2006 (N_2006,In_130,In_2122);
xor U2007 (N_2007,In_2254,In_1292);
xor U2008 (N_2008,In_342,In_1229);
and U2009 (N_2009,In_469,In_740);
nor U2010 (N_2010,In_231,In_1705);
nor U2011 (N_2011,In_476,In_279);
and U2012 (N_2012,In_1942,In_918);
nand U2013 (N_2013,In_2178,In_926);
nor U2014 (N_2014,In_2322,In_1933);
nand U2015 (N_2015,In_981,In_190);
and U2016 (N_2016,In_976,In_1183);
or U2017 (N_2017,In_1555,In_2081);
or U2018 (N_2018,In_65,In_1493);
nor U2019 (N_2019,In_521,In_848);
nor U2020 (N_2020,In_1121,In_1749);
xnor U2021 (N_2021,In_666,In_551);
nand U2022 (N_2022,In_34,In_1580);
or U2023 (N_2023,In_567,In_2325);
or U2024 (N_2024,In_1031,In_851);
nor U2025 (N_2025,In_869,In_541);
or U2026 (N_2026,In_1078,In_1018);
or U2027 (N_2027,In_678,In_1243);
nor U2028 (N_2028,In_1498,In_998);
or U2029 (N_2029,In_1994,In_619);
nor U2030 (N_2030,In_1482,In_48);
nor U2031 (N_2031,In_2329,In_846);
nor U2032 (N_2032,In_1992,In_2186);
nand U2033 (N_2033,In_1277,In_1791);
or U2034 (N_2034,In_2416,In_1585);
or U2035 (N_2035,In_2150,In_631);
nand U2036 (N_2036,In_2050,In_2015);
and U2037 (N_2037,In_2165,In_1874);
or U2038 (N_2038,In_1527,In_1200);
or U2039 (N_2039,In_159,In_338);
nor U2040 (N_2040,In_669,In_2066);
nor U2041 (N_2041,In_857,In_1883);
and U2042 (N_2042,In_2377,In_755);
and U2043 (N_2043,In_1323,In_293);
or U2044 (N_2044,In_685,In_1900);
nand U2045 (N_2045,In_1761,In_389);
nor U2046 (N_2046,In_2199,In_1163);
and U2047 (N_2047,In_1960,In_1725);
nor U2048 (N_2048,In_1173,In_2320);
or U2049 (N_2049,In_1348,In_110);
and U2050 (N_2050,In_2354,In_674);
and U2051 (N_2051,In_1697,In_1551);
and U2052 (N_2052,In_2061,In_1048);
nor U2053 (N_2053,In_1291,In_2044);
nor U2054 (N_2054,In_23,In_892);
nor U2055 (N_2055,In_2401,In_831);
or U2056 (N_2056,In_1409,In_776);
and U2057 (N_2057,In_1216,In_533);
xnor U2058 (N_2058,In_1877,In_1084);
or U2059 (N_2059,In_1462,In_852);
or U2060 (N_2060,In_811,In_2242);
and U2061 (N_2061,In_128,In_2127);
nand U2062 (N_2062,In_1688,In_775);
nor U2063 (N_2063,In_2348,In_1089);
nand U2064 (N_2064,In_1908,In_1028);
and U2065 (N_2065,In_1721,In_1260);
nor U2066 (N_2066,In_1324,In_1417);
and U2067 (N_2067,In_315,In_2220);
or U2068 (N_2068,In_2344,In_1046);
and U2069 (N_2069,In_521,In_580);
nand U2070 (N_2070,In_505,In_2140);
nor U2071 (N_2071,In_1033,In_2223);
or U2072 (N_2072,In_1333,In_1486);
xnor U2073 (N_2073,In_1316,In_938);
and U2074 (N_2074,In_1659,In_2027);
and U2075 (N_2075,In_94,In_2369);
and U2076 (N_2076,In_859,In_462);
xor U2077 (N_2077,In_2297,In_678);
and U2078 (N_2078,In_1517,In_2314);
xor U2079 (N_2079,In_2433,In_2346);
and U2080 (N_2080,In_54,In_1959);
nand U2081 (N_2081,In_1262,In_1359);
nand U2082 (N_2082,In_557,In_498);
or U2083 (N_2083,In_881,In_1572);
nand U2084 (N_2084,In_1257,In_7);
and U2085 (N_2085,In_1945,In_2146);
nor U2086 (N_2086,In_1859,In_520);
nor U2087 (N_2087,In_1435,In_1978);
and U2088 (N_2088,In_1007,In_1702);
nand U2089 (N_2089,In_2153,In_1280);
nor U2090 (N_2090,In_2117,In_105);
nor U2091 (N_2091,In_1849,In_357);
xnor U2092 (N_2092,In_471,In_959);
and U2093 (N_2093,In_2141,In_1651);
xor U2094 (N_2094,In_2054,In_882);
and U2095 (N_2095,In_1376,In_1830);
or U2096 (N_2096,In_1492,In_2089);
or U2097 (N_2097,In_2474,In_1306);
and U2098 (N_2098,In_19,In_625);
and U2099 (N_2099,In_1523,In_1915);
nor U2100 (N_2100,In_2152,In_1657);
nand U2101 (N_2101,In_2104,In_1728);
xnor U2102 (N_2102,In_1125,In_1526);
or U2103 (N_2103,In_1658,In_412);
and U2104 (N_2104,In_1937,In_2412);
nand U2105 (N_2105,In_365,In_1604);
and U2106 (N_2106,In_1485,In_1152);
or U2107 (N_2107,In_1587,In_837);
or U2108 (N_2108,In_2068,In_1988);
and U2109 (N_2109,In_837,In_1715);
nor U2110 (N_2110,In_2016,In_1139);
nand U2111 (N_2111,In_802,In_935);
nor U2112 (N_2112,In_306,In_1927);
and U2113 (N_2113,In_2280,In_1793);
nor U2114 (N_2114,In_2499,In_2401);
and U2115 (N_2115,In_714,In_1199);
or U2116 (N_2116,In_1078,In_503);
nand U2117 (N_2117,In_2363,In_144);
nand U2118 (N_2118,In_359,In_1941);
nand U2119 (N_2119,In_2346,In_309);
or U2120 (N_2120,In_1499,In_236);
nand U2121 (N_2121,In_552,In_1490);
and U2122 (N_2122,In_149,In_447);
nand U2123 (N_2123,In_1294,In_1222);
nand U2124 (N_2124,In_1080,In_1572);
or U2125 (N_2125,In_16,In_2290);
xor U2126 (N_2126,In_566,In_1491);
nand U2127 (N_2127,In_1279,In_1515);
and U2128 (N_2128,In_425,In_1233);
or U2129 (N_2129,In_1544,In_896);
nand U2130 (N_2130,In_1172,In_2004);
or U2131 (N_2131,In_792,In_1838);
nand U2132 (N_2132,In_479,In_1375);
xor U2133 (N_2133,In_2475,In_1898);
and U2134 (N_2134,In_679,In_355);
or U2135 (N_2135,In_405,In_846);
and U2136 (N_2136,In_923,In_1486);
nand U2137 (N_2137,In_2065,In_174);
nor U2138 (N_2138,In_340,In_1949);
xnor U2139 (N_2139,In_142,In_2116);
or U2140 (N_2140,In_1446,In_1458);
nor U2141 (N_2141,In_2179,In_637);
nor U2142 (N_2142,In_1687,In_931);
xnor U2143 (N_2143,In_96,In_486);
and U2144 (N_2144,In_2132,In_370);
nand U2145 (N_2145,In_927,In_1595);
and U2146 (N_2146,In_1243,In_2314);
and U2147 (N_2147,In_594,In_2102);
and U2148 (N_2148,In_43,In_1454);
or U2149 (N_2149,In_819,In_728);
or U2150 (N_2150,In_1249,In_632);
or U2151 (N_2151,In_1660,In_2489);
and U2152 (N_2152,In_1250,In_1692);
nor U2153 (N_2153,In_1696,In_149);
or U2154 (N_2154,In_46,In_1421);
xnor U2155 (N_2155,In_2350,In_1604);
or U2156 (N_2156,In_682,In_367);
xnor U2157 (N_2157,In_471,In_1541);
nand U2158 (N_2158,In_1487,In_2354);
and U2159 (N_2159,In_325,In_2289);
nor U2160 (N_2160,In_535,In_2173);
nor U2161 (N_2161,In_2205,In_190);
and U2162 (N_2162,In_1250,In_226);
and U2163 (N_2163,In_220,In_2363);
or U2164 (N_2164,In_960,In_1526);
or U2165 (N_2165,In_2312,In_2083);
and U2166 (N_2166,In_1232,In_1224);
and U2167 (N_2167,In_1807,In_377);
and U2168 (N_2168,In_1908,In_1751);
nor U2169 (N_2169,In_2259,In_1694);
xor U2170 (N_2170,In_465,In_918);
nand U2171 (N_2171,In_787,In_1795);
nor U2172 (N_2172,In_1132,In_1879);
or U2173 (N_2173,In_2052,In_1441);
or U2174 (N_2174,In_2049,In_1351);
or U2175 (N_2175,In_343,In_1210);
and U2176 (N_2176,In_1240,In_1413);
and U2177 (N_2177,In_597,In_756);
and U2178 (N_2178,In_588,In_1493);
or U2179 (N_2179,In_1330,In_1601);
nor U2180 (N_2180,In_1675,In_1796);
xor U2181 (N_2181,In_217,In_2433);
nand U2182 (N_2182,In_1360,In_1442);
or U2183 (N_2183,In_2116,In_1696);
or U2184 (N_2184,In_2045,In_1644);
nand U2185 (N_2185,In_606,In_940);
and U2186 (N_2186,In_2432,In_394);
or U2187 (N_2187,In_1717,In_131);
nand U2188 (N_2188,In_2418,In_2400);
or U2189 (N_2189,In_2024,In_1783);
nor U2190 (N_2190,In_1100,In_99);
or U2191 (N_2191,In_2454,In_1675);
nand U2192 (N_2192,In_540,In_1727);
or U2193 (N_2193,In_2268,In_1152);
and U2194 (N_2194,In_1187,In_1399);
or U2195 (N_2195,In_2190,In_815);
or U2196 (N_2196,In_416,In_2128);
nor U2197 (N_2197,In_77,In_1665);
and U2198 (N_2198,In_2178,In_909);
or U2199 (N_2199,In_541,In_341);
and U2200 (N_2200,In_2221,In_1410);
nor U2201 (N_2201,In_2318,In_1775);
and U2202 (N_2202,In_824,In_2292);
and U2203 (N_2203,In_274,In_2464);
nor U2204 (N_2204,In_730,In_988);
xnor U2205 (N_2205,In_2264,In_1373);
nor U2206 (N_2206,In_1074,In_2181);
nor U2207 (N_2207,In_1901,In_1496);
nand U2208 (N_2208,In_740,In_2292);
or U2209 (N_2209,In_1977,In_1679);
nand U2210 (N_2210,In_2289,In_2206);
nor U2211 (N_2211,In_793,In_2027);
nor U2212 (N_2212,In_1669,In_1238);
or U2213 (N_2213,In_768,In_194);
xor U2214 (N_2214,In_377,In_805);
nand U2215 (N_2215,In_129,In_1560);
nor U2216 (N_2216,In_874,In_2030);
nor U2217 (N_2217,In_194,In_1633);
nor U2218 (N_2218,In_643,In_149);
and U2219 (N_2219,In_954,In_1721);
nand U2220 (N_2220,In_846,In_2270);
xnor U2221 (N_2221,In_2113,In_504);
nand U2222 (N_2222,In_1619,In_569);
and U2223 (N_2223,In_2196,In_2386);
and U2224 (N_2224,In_1383,In_876);
and U2225 (N_2225,In_1378,In_488);
or U2226 (N_2226,In_807,In_1519);
or U2227 (N_2227,In_1499,In_332);
xnor U2228 (N_2228,In_192,In_143);
or U2229 (N_2229,In_1245,In_223);
or U2230 (N_2230,In_358,In_2209);
and U2231 (N_2231,In_1475,In_946);
and U2232 (N_2232,In_1065,In_585);
nor U2233 (N_2233,In_837,In_1417);
nand U2234 (N_2234,In_1433,In_1203);
or U2235 (N_2235,In_1466,In_2080);
nand U2236 (N_2236,In_1261,In_872);
nor U2237 (N_2237,In_343,In_485);
nand U2238 (N_2238,In_1956,In_2198);
nand U2239 (N_2239,In_2042,In_1893);
and U2240 (N_2240,In_383,In_706);
nor U2241 (N_2241,In_41,In_117);
xnor U2242 (N_2242,In_1706,In_642);
and U2243 (N_2243,In_1938,In_1903);
nand U2244 (N_2244,In_890,In_856);
nor U2245 (N_2245,In_644,In_974);
xor U2246 (N_2246,In_1038,In_2453);
nand U2247 (N_2247,In_644,In_953);
xnor U2248 (N_2248,In_445,In_1301);
xnor U2249 (N_2249,In_105,In_196);
and U2250 (N_2250,In_97,In_279);
nor U2251 (N_2251,In_690,In_2419);
nand U2252 (N_2252,In_789,In_1214);
or U2253 (N_2253,In_1476,In_2464);
nand U2254 (N_2254,In_135,In_93);
and U2255 (N_2255,In_389,In_68);
or U2256 (N_2256,In_1598,In_1526);
and U2257 (N_2257,In_2250,In_1854);
or U2258 (N_2258,In_2172,In_1276);
xor U2259 (N_2259,In_766,In_124);
or U2260 (N_2260,In_2297,In_315);
nor U2261 (N_2261,In_2003,In_2480);
or U2262 (N_2262,In_1934,In_1441);
and U2263 (N_2263,In_2405,In_734);
nand U2264 (N_2264,In_1539,In_2038);
or U2265 (N_2265,In_655,In_94);
and U2266 (N_2266,In_2239,In_1681);
nand U2267 (N_2267,In_1775,In_1403);
nand U2268 (N_2268,In_1587,In_1393);
or U2269 (N_2269,In_1985,In_365);
nand U2270 (N_2270,In_459,In_1480);
and U2271 (N_2271,In_2140,In_1818);
nor U2272 (N_2272,In_466,In_1591);
and U2273 (N_2273,In_1075,In_1663);
and U2274 (N_2274,In_204,In_2105);
nor U2275 (N_2275,In_660,In_1448);
nand U2276 (N_2276,In_145,In_1493);
and U2277 (N_2277,In_258,In_1043);
nand U2278 (N_2278,In_933,In_1262);
nand U2279 (N_2279,In_849,In_899);
nand U2280 (N_2280,In_1647,In_1056);
and U2281 (N_2281,In_1256,In_1576);
xor U2282 (N_2282,In_1692,In_1776);
nor U2283 (N_2283,In_318,In_47);
nand U2284 (N_2284,In_1319,In_386);
and U2285 (N_2285,In_423,In_1365);
nor U2286 (N_2286,In_1286,In_1653);
and U2287 (N_2287,In_836,In_1420);
nand U2288 (N_2288,In_2240,In_2475);
nand U2289 (N_2289,In_1660,In_2325);
nand U2290 (N_2290,In_617,In_370);
and U2291 (N_2291,In_194,In_1572);
nor U2292 (N_2292,In_1124,In_212);
or U2293 (N_2293,In_953,In_256);
nor U2294 (N_2294,In_1140,In_291);
nand U2295 (N_2295,In_9,In_108);
and U2296 (N_2296,In_689,In_335);
xor U2297 (N_2297,In_2206,In_428);
or U2298 (N_2298,In_202,In_2194);
nor U2299 (N_2299,In_2310,In_1106);
nand U2300 (N_2300,In_1638,In_1593);
and U2301 (N_2301,In_1891,In_50);
nor U2302 (N_2302,In_1652,In_978);
nor U2303 (N_2303,In_1711,In_575);
nor U2304 (N_2304,In_1439,In_804);
or U2305 (N_2305,In_1454,In_2416);
or U2306 (N_2306,In_413,In_279);
and U2307 (N_2307,In_831,In_48);
nand U2308 (N_2308,In_752,In_896);
and U2309 (N_2309,In_13,In_1659);
or U2310 (N_2310,In_2195,In_820);
xnor U2311 (N_2311,In_589,In_1801);
or U2312 (N_2312,In_554,In_471);
xnor U2313 (N_2313,In_1127,In_1578);
xor U2314 (N_2314,In_439,In_807);
and U2315 (N_2315,In_1875,In_2107);
or U2316 (N_2316,In_1879,In_386);
and U2317 (N_2317,In_1641,In_534);
and U2318 (N_2318,In_1060,In_2061);
nand U2319 (N_2319,In_198,In_2135);
nor U2320 (N_2320,In_1914,In_125);
nor U2321 (N_2321,In_316,In_155);
nor U2322 (N_2322,In_1827,In_1787);
xnor U2323 (N_2323,In_2495,In_892);
and U2324 (N_2324,In_2201,In_512);
nor U2325 (N_2325,In_148,In_833);
or U2326 (N_2326,In_1386,In_1536);
nor U2327 (N_2327,In_1463,In_79);
or U2328 (N_2328,In_579,In_531);
or U2329 (N_2329,In_1545,In_167);
nor U2330 (N_2330,In_1992,In_1906);
nor U2331 (N_2331,In_1826,In_1841);
nor U2332 (N_2332,In_1196,In_681);
and U2333 (N_2333,In_2392,In_1460);
or U2334 (N_2334,In_161,In_1608);
nand U2335 (N_2335,In_1320,In_1747);
xor U2336 (N_2336,In_1770,In_846);
or U2337 (N_2337,In_2237,In_372);
xor U2338 (N_2338,In_50,In_1641);
nor U2339 (N_2339,In_1561,In_2338);
and U2340 (N_2340,In_2441,In_221);
nor U2341 (N_2341,In_2480,In_1641);
nand U2342 (N_2342,In_2112,In_370);
and U2343 (N_2343,In_1894,In_2149);
or U2344 (N_2344,In_1064,In_1954);
nand U2345 (N_2345,In_1316,In_696);
nand U2346 (N_2346,In_1490,In_1342);
and U2347 (N_2347,In_1856,In_1649);
and U2348 (N_2348,In_2124,In_2217);
and U2349 (N_2349,In_525,In_2174);
and U2350 (N_2350,In_2499,In_2387);
nand U2351 (N_2351,In_1692,In_2385);
and U2352 (N_2352,In_2188,In_939);
nand U2353 (N_2353,In_1490,In_614);
nand U2354 (N_2354,In_1566,In_1068);
or U2355 (N_2355,In_1072,In_1792);
and U2356 (N_2356,In_43,In_2167);
nor U2357 (N_2357,In_459,In_1388);
xnor U2358 (N_2358,In_2337,In_1451);
or U2359 (N_2359,In_1159,In_1905);
nand U2360 (N_2360,In_827,In_518);
nand U2361 (N_2361,In_1931,In_1956);
nor U2362 (N_2362,In_602,In_2466);
nor U2363 (N_2363,In_2014,In_2358);
nand U2364 (N_2364,In_93,In_1211);
and U2365 (N_2365,In_1143,In_1784);
or U2366 (N_2366,In_272,In_627);
or U2367 (N_2367,In_2268,In_461);
nand U2368 (N_2368,In_1771,In_1722);
and U2369 (N_2369,In_701,In_402);
or U2370 (N_2370,In_380,In_620);
and U2371 (N_2371,In_929,In_285);
and U2372 (N_2372,In_1467,In_248);
or U2373 (N_2373,In_1424,In_1212);
xnor U2374 (N_2374,In_646,In_2471);
nor U2375 (N_2375,In_1455,In_1226);
or U2376 (N_2376,In_2107,In_186);
nand U2377 (N_2377,In_1261,In_1599);
or U2378 (N_2378,In_2499,In_1732);
and U2379 (N_2379,In_204,In_2287);
and U2380 (N_2380,In_2189,In_484);
nand U2381 (N_2381,In_2006,In_2150);
nand U2382 (N_2382,In_709,In_185);
nand U2383 (N_2383,In_2308,In_1574);
nor U2384 (N_2384,In_392,In_1574);
xor U2385 (N_2385,In_1259,In_1667);
nor U2386 (N_2386,In_1839,In_2150);
nand U2387 (N_2387,In_186,In_2483);
or U2388 (N_2388,In_2134,In_820);
nand U2389 (N_2389,In_2203,In_2442);
xor U2390 (N_2390,In_380,In_1866);
nand U2391 (N_2391,In_1871,In_1926);
nor U2392 (N_2392,In_1306,In_1425);
and U2393 (N_2393,In_2400,In_2037);
nand U2394 (N_2394,In_580,In_1335);
nand U2395 (N_2395,In_46,In_1281);
nor U2396 (N_2396,In_2331,In_479);
nand U2397 (N_2397,In_2431,In_1856);
or U2398 (N_2398,In_1465,In_8);
nand U2399 (N_2399,In_1665,In_2328);
and U2400 (N_2400,In_867,In_1784);
nand U2401 (N_2401,In_1959,In_2410);
nor U2402 (N_2402,In_723,In_557);
nand U2403 (N_2403,In_1554,In_2399);
or U2404 (N_2404,In_2334,In_1106);
nor U2405 (N_2405,In_37,In_2131);
nand U2406 (N_2406,In_1322,In_887);
nor U2407 (N_2407,In_324,In_2144);
nor U2408 (N_2408,In_1276,In_849);
and U2409 (N_2409,In_2205,In_2484);
nand U2410 (N_2410,In_430,In_1404);
nor U2411 (N_2411,In_2023,In_147);
xnor U2412 (N_2412,In_2130,In_1181);
or U2413 (N_2413,In_1471,In_306);
xor U2414 (N_2414,In_895,In_2311);
nand U2415 (N_2415,In_1817,In_626);
nand U2416 (N_2416,In_2020,In_1989);
nor U2417 (N_2417,In_1053,In_2392);
xnor U2418 (N_2418,In_876,In_594);
and U2419 (N_2419,In_944,In_1072);
nand U2420 (N_2420,In_1249,In_886);
xnor U2421 (N_2421,In_2401,In_1144);
nand U2422 (N_2422,In_214,In_860);
nand U2423 (N_2423,In_730,In_2434);
and U2424 (N_2424,In_2436,In_292);
and U2425 (N_2425,In_275,In_2342);
and U2426 (N_2426,In_694,In_1541);
and U2427 (N_2427,In_1392,In_2220);
and U2428 (N_2428,In_530,In_312);
nand U2429 (N_2429,In_2412,In_17);
or U2430 (N_2430,In_302,In_349);
nand U2431 (N_2431,In_746,In_19);
nand U2432 (N_2432,In_2092,In_1289);
and U2433 (N_2433,In_320,In_406);
nand U2434 (N_2434,In_1027,In_1842);
nor U2435 (N_2435,In_1408,In_734);
or U2436 (N_2436,In_724,In_122);
or U2437 (N_2437,In_1206,In_1765);
nand U2438 (N_2438,In_1086,In_802);
and U2439 (N_2439,In_2035,In_1215);
or U2440 (N_2440,In_1986,In_72);
nor U2441 (N_2441,In_149,In_533);
nor U2442 (N_2442,In_2211,In_2306);
or U2443 (N_2443,In_2000,In_1884);
nand U2444 (N_2444,In_1352,In_1567);
and U2445 (N_2445,In_2421,In_27);
or U2446 (N_2446,In_337,In_651);
nor U2447 (N_2447,In_2281,In_564);
nor U2448 (N_2448,In_2301,In_1591);
nor U2449 (N_2449,In_109,In_243);
xor U2450 (N_2450,In_2157,In_923);
and U2451 (N_2451,In_933,In_2040);
nand U2452 (N_2452,In_2102,In_1205);
nand U2453 (N_2453,In_1977,In_417);
or U2454 (N_2454,In_446,In_1826);
and U2455 (N_2455,In_2120,In_698);
nor U2456 (N_2456,In_1772,In_788);
nor U2457 (N_2457,In_1310,In_1319);
nor U2458 (N_2458,In_893,In_1643);
nor U2459 (N_2459,In_1044,In_1626);
nand U2460 (N_2460,In_1431,In_1712);
or U2461 (N_2461,In_764,In_99);
or U2462 (N_2462,In_429,In_1505);
and U2463 (N_2463,In_1253,In_1394);
xor U2464 (N_2464,In_410,In_1819);
nand U2465 (N_2465,In_530,In_421);
nor U2466 (N_2466,In_975,In_1136);
nand U2467 (N_2467,In_1985,In_695);
nor U2468 (N_2468,In_1644,In_2314);
nor U2469 (N_2469,In_2222,In_834);
or U2470 (N_2470,In_261,In_1814);
nor U2471 (N_2471,In_1888,In_2414);
and U2472 (N_2472,In_840,In_555);
and U2473 (N_2473,In_257,In_2328);
or U2474 (N_2474,In_1547,In_363);
and U2475 (N_2475,In_516,In_2151);
nor U2476 (N_2476,In_466,In_2283);
and U2477 (N_2477,In_1682,In_1282);
and U2478 (N_2478,In_88,In_1432);
and U2479 (N_2479,In_885,In_2383);
or U2480 (N_2480,In_440,In_104);
nor U2481 (N_2481,In_1568,In_73);
and U2482 (N_2482,In_1974,In_857);
nor U2483 (N_2483,In_1102,In_475);
nand U2484 (N_2484,In_1328,In_201);
nor U2485 (N_2485,In_1750,In_481);
nor U2486 (N_2486,In_879,In_1054);
nand U2487 (N_2487,In_2394,In_475);
and U2488 (N_2488,In_2225,In_1260);
xnor U2489 (N_2489,In_2005,In_172);
nand U2490 (N_2490,In_1383,In_1472);
nor U2491 (N_2491,In_775,In_1095);
nand U2492 (N_2492,In_554,In_341);
nor U2493 (N_2493,In_426,In_132);
and U2494 (N_2494,In_1754,In_1558);
nor U2495 (N_2495,In_183,In_2260);
xor U2496 (N_2496,In_1826,In_143);
or U2497 (N_2497,In_981,In_256);
xor U2498 (N_2498,In_1858,In_1012);
and U2499 (N_2499,In_1781,In_471);
nor U2500 (N_2500,In_1481,In_1795);
xor U2501 (N_2501,In_1138,In_901);
or U2502 (N_2502,In_1403,In_2414);
and U2503 (N_2503,In_2147,In_1870);
or U2504 (N_2504,In_1455,In_896);
nor U2505 (N_2505,In_809,In_805);
and U2506 (N_2506,In_1007,In_691);
or U2507 (N_2507,In_1097,In_135);
or U2508 (N_2508,In_800,In_2006);
or U2509 (N_2509,In_1651,In_2426);
nor U2510 (N_2510,In_2224,In_67);
nor U2511 (N_2511,In_1017,In_2012);
nor U2512 (N_2512,In_629,In_809);
or U2513 (N_2513,In_1868,In_268);
nor U2514 (N_2514,In_747,In_390);
nor U2515 (N_2515,In_2413,In_1317);
or U2516 (N_2516,In_1928,In_25);
and U2517 (N_2517,In_1285,In_1797);
nand U2518 (N_2518,In_2402,In_1240);
nand U2519 (N_2519,In_1819,In_1460);
nand U2520 (N_2520,In_305,In_696);
or U2521 (N_2521,In_858,In_876);
or U2522 (N_2522,In_222,In_2278);
xnor U2523 (N_2523,In_270,In_906);
or U2524 (N_2524,In_43,In_1705);
or U2525 (N_2525,In_1312,In_1644);
or U2526 (N_2526,In_2006,In_1750);
xor U2527 (N_2527,In_1443,In_2453);
xor U2528 (N_2528,In_1300,In_140);
nand U2529 (N_2529,In_2085,In_1214);
nor U2530 (N_2530,In_610,In_202);
and U2531 (N_2531,In_682,In_2231);
xor U2532 (N_2532,In_905,In_1042);
nor U2533 (N_2533,In_2287,In_305);
nor U2534 (N_2534,In_2087,In_804);
nand U2535 (N_2535,In_1772,In_1834);
nor U2536 (N_2536,In_1629,In_1049);
or U2537 (N_2537,In_185,In_1019);
or U2538 (N_2538,In_978,In_1907);
nand U2539 (N_2539,In_734,In_1268);
nand U2540 (N_2540,In_1252,In_705);
and U2541 (N_2541,In_1672,In_1231);
nor U2542 (N_2542,In_70,In_1080);
nor U2543 (N_2543,In_836,In_1648);
xor U2544 (N_2544,In_1133,In_2331);
nand U2545 (N_2545,In_512,In_660);
and U2546 (N_2546,In_96,In_636);
and U2547 (N_2547,In_1961,In_409);
and U2548 (N_2548,In_1665,In_2167);
nor U2549 (N_2549,In_171,In_639);
nor U2550 (N_2550,In_1281,In_1914);
and U2551 (N_2551,In_658,In_1951);
xor U2552 (N_2552,In_1152,In_1596);
nor U2553 (N_2553,In_1355,In_2226);
nor U2554 (N_2554,In_2159,In_1103);
nand U2555 (N_2555,In_2253,In_1034);
xnor U2556 (N_2556,In_745,In_72);
nand U2557 (N_2557,In_1991,In_1518);
nand U2558 (N_2558,In_754,In_1431);
and U2559 (N_2559,In_2300,In_944);
nand U2560 (N_2560,In_1582,In_463);
xor U2561 (N_2561,In_1019,In_1945);
xor U2562 (N_2562,In_1600,In_827);
nor U2563 (N_2563,In_235,In_1176);
nand U2564 (N_2564,In_2231,In_1640);
and U2565 (N_2565,In_1975,In_1429);
nor U2566 (N_2566,In_2032,In_2049);
or U2567 (N_2567,In_2468,In_1381);
and U2568 (N_2568,In_448,In_923);
and U2569 (N_2569,In_783,In_1387);
nand U2570 (N_2570,In_422,In_1498);
nor U2571 (N_2571,In_2334,In_777);
and U2572 (N_2572,In_1402,In_1356);
nor U2573 (N_2573,In_269,In_1862);
nand U2574 (N_2574,In_1586,In_706);
xnor U2575 (N_2575,In_545,In_1962);
nor U2576 (N_2576,In_1218,In_1252);
or U2577 (N_2577,In_866,In_1564);
xor U2578 (N_2578,In_1172,In_2268);
nand U2579 (N_2579,In_1969,In_1566);
nand U2580 (N_2580,In_1575,In_1337);
or U2581 (N_2581,In_1151,In_1463);
and U2582 (N_2582,In_1241,In_194);
nor U2583 (N_2583,In_2275,In_2269);
xor U2584 (N_2584,In_2169,In_2487);
nand U2585 (N_2585,In_1554,In_21);
xor U2586 (N_2586,In_1124,In_1398);
xnor U2587 (N_2587,In_2260,In_383);
nand U2588 (N_2588,In_1396,In_1448);
and U2589 (N_2589,In_406,In_507);
xnor U2590 (N_2590,In_2346,In_78);
nor U2591 (N_2591,In_1356,In_1493);
or U2592 (N_2592,In_695,In_2260);
xnor U2593 (N_2593,In_803,In_18);
nor U2594 (N_2594,In_1327,In_574);
or U2595 (N_2595,In_859,In_2086);
xor U2596 (N_2596,In_702,In_1099);
and U2597 (N_2597,In_2357,In_1227);
nor U2598 (N_2598,In_2309,In_169);
or U2599 (N_2599,In_213,In_1227);
nor U2600 (N_2600,In_2039,In_1757);
and U2601 (N_2601,In_1891,In_663);
nor U2602 (N_2602,In_560,In_20);
nor U2603 (N_2603,In_830,In_2314);
xnor U2604 (N_2604,In_2051,In_1934);
and U2605 (N_2605,In_2013,In_2273);
nand U2606 (N_2606,In_1262,In_871);
nand U2607 (N_2607,In_1528,In_41);
nor U2608 (N_2608,In_1349,In_2369);
nand U2609 (N_2609,In_456,In_478);
nor U2610 (N_2610,In_573,In_1978);
nand U2611 (N_2611,In_2204,In_1781);
nor U2612 (N_2612,In_2331,In_711);
nand U2613 (N_2613,In_1354,In_1675);
xor U2614 (N_2614,In_1099,In_178);
nand U2615 (N_2615,In_1560,In_304);
or U2616 (N_2616,In_604,In_2290);
nor U2617 (N_2617,In_746,In_915);
or U2618 (N_2618,In_2314,In_1244);
or U2619 (N_2619,In_1140,In_2492);
or U2620 (N_2620,In_1538,In_313);
or U2621 (N_2621,In_406,In_409);
and U2622 (N_2622,In_672,In_1189);
xnor U2623 (N_2623,In_1500,In_77);
nor U2624 (N_2624,In_1645,In_2428);
and U2625 (N_2625,In_2432,In_2226);
or U2626 (N_2626,In_1942,In_1916);
nor U2627 (N_2627,In_1037,In_892);
nor U2628 (N_2628,In_1368,In_122);
nand U2629 (N_2629,In_221,In_147);
xor U2630 (N_2630,In_693,In_1556);
or U2631 (N_2631,In_1582,In_2182);
and U2632 (N_2632,In_1646,In_1868);
nand U2633 (N_2633,In_1542,In_1216);
nor U2634 (N_2634,In_43,In_632);
xor U2635 (N_2635,In_1651,In_1255);
nor U2636 (N_2636,In_10,In_614);
nor U2637 (N_2637,In_1906,In_2450);
and U2638 (N_2638,In_2476,In_1673);
nor U2639 (N_2639,In_1631,In_1109);
xor U2640 (N_2640,In_1776,In_1641);
xnor U2641 (N_2641,In_807,In_985);
nand U2642 (N_2642,In_2206,In_696);
xor U2643 (N_2643,In_1900,In_2339);
nand U2644 (N_2644,In_301,In_447);
nand U2645 (N_2645,In_2101,In_1117);
nor U2646 (N_2646,In_1100,In_2159);
or U2647 (N_2647,In_1098,In_1577);
or U2648 (N_2648,In_2487,In_709);
nand U2649 (N_2649,In_1004,In_1590);
nand U2650 (N_2650,In_1952,In_1886);
and U2651 (N_2651,In_1164,In_1497);
and U2652 (N_2652,In_1205,In_2167);
nor U2653 (N_2653,In_1517,In_535);
or U2654 (N_2654,In_2111,In_2009);
or U2655 (N_2655,In_2398,In_1914);
and U2656 (N_2656,In_913,In_1129);
and U2657 (N_2657,In_2216,In_469);
xor U2658 (N_2658,In_1497,In_1897);
and U2659 (N_2659,In_999,In_1862);
or U2660 (N_2660,In_1105,In_903);
and U2661 (N_2661,In_2030,In_1888);
nor U2662 (N_2662,In_1020,In_1781);
or U2663 (N_2663,In_2144,In_383);
xor U2664 (N_2664,In_1294,In_199);
and U2665 (N_2665,In_1020,In_1140);
nor U2666 (N_2666,In_2234,In_1673);
nand U2667 (N_2667,In_2170,In_153);
nand U2668 (N_2668,In_1099,In_2110);
and U2669 (N_2669,In_120,In_1274);
nand U2670 (N_2670,In_1935,In_2068);
nor U2671 (N_2671,In_852,In_745);
or U2672 (N_2672,In_1820,In_2069);
nor U2673 (N_2673,In_2017,In_213);
nor U2674 (N_2674,In_1660,In_383);
nor U2675 (N_2675,In_1630,In_1800);
nor U2676 (N_2676,In_79,In_1006);
or U2677 (N_2677,In_837,In_1409);
or U2678 (N_2678,In_108,In_261);
nor U2679 (N_2679,In_773,In_501);
and U2680 (N_2680,In_823,In_713);
and U2681 (N_2681,In_1866,In_1412);
nor U2682 (N_2682,In_1832,In_2483);
and U2683 (N_2683,In_2303,In_2120);
nor U2684 (N_2684,In_2180,In_1434);
and U2685 (N_2685,In_2047,In_734);
and U2686 (N_2686,In_491,In_1541);
nand U2687 (N_2687,In_598,In_1850);
and U2688 (N_2688,In_2275,In_88);
xnor U2689 (N_2689,In_1043,In_460);
or U2690 (N_2690,In_2262,In_1116);
nor U2691 (N_2691,In_184,In_1984);
and U2692 (N_2692,In_1300,In_61);
nand U2693 (N_2693,In_960,In_1004);
xor U2694 (N_2694,In_282,In_1936);
xor U2695 (N_2695,In_498,In_2001);
or U2696 (N_2696,In_1435,In_1013);
nand U2697 (N_2697,In_104,In_769);
nor U2698 (N_2698,In_336,In_1825);
xnor U2699 (N_2699,In_2236,In_611);
nand U2700 (N_2700,In_1692,In_915);
and U2701 (N_2701,In_393,In_1286);
nand U2702 (N_2702,In_1042,In_1333);
and U2703 (N_2703,In_1814,In_93);
nor U2704 (N_2704,In_1523,In_543);
nor U2705 (N_2705,In_1431,In_1340);
and U2706 (N_2706,In_283,In_970);
nor U2707 (N_2707,In_1901,In_2394);
and U2708 (N_2708,In_2473,In_2278);
and U2709 (N_2709,In_695,In_915);
nand U2710 (N_2710,In_293,In_1410);
or U2711 (N_2711,In_2328,In_38);
or U2712 (N_2712,In_2336,In_245);
or U2713 (N_2713,In_736,In_2418);
or U2714 (N_2714,In_850,In_1709);
and U2715 (N_2715,In_1185,In_1575);
nor U2716 (N_2716,In_2322,In_318);
nand U2717 (N_2717,In_1488,In_1750);
or U2718 (N_2718,In_1971,In_13);
nand U2719 (N_2719,In_939,In_455);
xnor U2720 (N_2720,In_713,In_264);
xor U2721 (N_2721,In_2106,In_419);
xor U2722 (N_2722,In_152,In_550);
nand U2723 (N_2723,In_1869,In_631);
and U2724 (N_2724,In_2387,In_1574);
xnor U2725 (N_2725,In_788,In_731);
nor U2726 (N_2726,In_1744,In_876);
nor U2727 (N_2727,In_2444,In_502);
and U2728 (N_2728,In_1585,In_717);
and U2729 (N_2729,In_2157,In_350);
nor U2730 (N_2730,In_1006,In_1198);
nor U2731 (N_2731,In_438,In_465);
nor U2732 (N_2732,In_920,In_1340);
nor U2733 (N_2733,In_1107,In_90);
and U2734 (N_2734,In_928,In_1143);
or U2735 (N_2735,In_1639,In_2047);
nor U2736 (N_2736,In_412,In_133);
nor U2737 (N_2737,In_2434,In_1838);
or U2738 (N_2738,In_1506,In_210);
nand U2739 (N_2739,In_916,In_2155);
nor U2740 (N_2740,In_1610,In_1307);
nor U2741 (N_2741,In_1442,In_1808);
and U2742 (N_2742,In_909,In_2184);
nor U2743 (N_2743,In_1638,In_2423);
nand U2744 (N_2744,In_2223,In_1997);
xor U2745 (N_2745,In_2416,In_90);
nor U2746 (N_2746,In_2328,In_283);
and U2747 (N_2747,In_248,In_1219);
or U2748 (N_2748,In_2420,In_1402);
nor U2749 (N_2749,In_2161,In_1586);
nand U2750 (N_2750,In_1757,In_1991);
xor U2751 (N_2751,In_1151,In_1607);
and U2752 (N_2752,In_79,In_1794);
or U2753 (N_2753,In_1037,In_2376);
nor U2754 (N_2754,In_1060,In_791);
xor U2755 (N_2755,In_1455,In_124);
xnor U2756 (N_2756,In_2353,In_215);
nor U2757 (N_2757,In_544,In_2056);
or U2758 (N_2758,In_333,In_718);
nand U2759 (N_2759,In_659,In_54);
xor U2760 (N_2760,In_52,In_1801);
nor U2761 (N_2761,In_1771,In_1790);
and U2762 (N_2762,In_1571,In_504);
and U2763 (N_2763,In_1082,In_1742);
nor U2764 (N_2764,In_180,In_1391);
nor U2765 (N_2765,In_1352,In_386);
nor U2766 (N_2766,In_2184,In_1332);
and U2767 (N_2767,In_2457,In_571);
and U2768 (N_2768,In_91,In_2036);
nor U2769 (N_2769,In_2181,In_2328);
and U2770 (N_2770,In_2168,In_689);
or U2771 (N_2771,In_607,In_1591);
and U2772 (N_2772,In_545,In_2404);
nand U2773 (N_2773,In_1965,In_1649);
nand U2774 (N_2774,In_1331,In_1759);
and U2775 (N_2775,In_1647,In_26);
nand U2776 (N_2776,In_312,In_2142);
or U2777 (N_2777,In_265,In_2373);
nand U2778 (N_2778,In_221,In_291);
or U2779 (N_2779,In_410,In_241);
nand U2780 (N_2780,In_1341,In_2357);
or U2781 (N_2781,In_475,In_2451);
and U2782 (N_2782,In_567,In_385);
and U2783 (N_2783,In_1273,In_2065);
nor U2784 (N_2784,In_1421,In_2160);
nand U2785 (N_2785,In_1560,In_599);
or U2786 (N_2786,In_1886,In_610);
xnor U2787 (N_2787,In_551,In_211);
and U2788 (N_2788,In_702,In_520);
or U2789 (N_2789,In_1933,In_2362);
nand U2790 (N_2790,In_1260,In_1647);
xor U2791 (N_2791,In_783,In_2068);
or U2792 (N_2792,In_1509,In_2372);
nand U2793 (N_2793,In_227,In_1662);
and U2794 (N_2794,In_1152,In_128);
or U2795 (N_2795,In_2221,In_1603);
nand U2796 (N_2796,In_2385,In_1236);
xnor U2797 (N_2797,In_1802,In_1478);
or U2798 (N_2798,In_2002,In_188);
and U2799 (N_2799,In_2176,In_1608);
nand U2800 (N_2800,In_515,In_2040);
and U2801 (N_2801,In_430,In_20);
or U2802 (N_2802,In_398,In_138);
or U2803 (N_2803,In_733,In_1517);
nor U2804 (N_2804,In_2405,In_270);
nor U2805 (N_2805,In_81,In_886);
or U2806 (N_2806,In_774,In_1649);
or U2807 (N_2807,In_1540,In_1105);
nor U2808 (N_2808,In_898,In_1720);
nor U2809 (N_2809,In_549,In_14);
and U2810 (N_2810,In_1881,In_1393);
and U2811 (N_2811,In_1292,In_987);
nor U2812 (N_2812,In_367,In_1884);
and U2813 (N_2813,In_1355,In_349);
or U2814 (N_2814,In_1866,In_1254);
and U2815 (N_2815,In_1121,In_125);
or U2816 (N_2816,In_332,In_2172);
and U2817 (N_2817,In_63,In_1375);
nand U2818 (N_2818,In_1374,In_1260);
nor U2819 (N_2819,In_495,In_1888);
nand U2820 (N_2820,In_1050,In_2196);
xnor U2821 (N_2821,In_648,In_1072);
nand U2822 (N_2822,In_1895,In_1248);
or U2823 (N_2823,In_553,In_1032);
and U2824 (N_2824,In_944,In_1011);
or U2825 (N_2825,In_2447,In_810);
nor U2826 (N_2826,In_1155,In_1364);
and U2827 (N_2827,In_957,In_199);
nand U2828 (N_2828,In_1936,In_1518);
nand U2829 (N_2829,In_1449,In_2429);
xnor U2830 (N_2830,In_330,In_2384);
and U2831 (N_2831,In_861,In_2072);
xor U2832 (N_2832,In_805,In_1583);
or U2833 (N_2833,In_1459,In_288);
and U2834 (N_2834,In_1399,In_253);
and U2835 (N_2835,In_639,In_1874);
nor U2836 (N_2836,In_1268,In_38);
or U2837 (N_2837,In_713,In_2155);
or U2838 (N_2838,In_1521,In_2041);
and U2839 (N_2839,In_2473,In_1195);
or U2840 (N_2840,In_2160,In_1053);
nand U2841 (N_2841,In_2396,In_1838);
and U2842 (N_2842,In_1362,In_680);
nand U2843 (N_2843,In_2043,In_2489);
and U2844 (N_2844,In_1442,In_1680);
xnor U2845 (N_2845,In_999,In_394);
or U2846 (N_2846,In_2272,In_1973);
nor U2847 (N_2847,In_142,In_2082);
and U2848 (N_2848,In_1830,In_543);
nor U2849 (N_2849,In_2208,In_655);
or U2850 (N_2850,In_2016,In_23);
nand U2851 (N_2851,In_431,In_490);
and U2852 (N_2852,In_1797,In_1097);
nor U2853 (N_2853,In_350,In_1834);
or U2854 (N_2854,In_2261,In_2286);
nor U2855 (N_2855,In_1241,In_86);
nand U2856 (N_2856,In_1217,In_2352);
and U2857 (N_2857,In_1441,In_2077);
or U2858 (N_2858,In_1559,In_1054);
or U2859 (N_2859,In_385,In_456);
nor U2860 (N_2860,In_83,In_954);
nor U2861 (N_2861,In_2081,In_1959);
and U2862 (N_2862,In_161,In_2421);
nand U2863 (N_2863,In_455,In_362);
nor U2864 (N_2864,In_1668,In_339);
and U2865 (N_2865,In_1617,In_1990);
nor U2866 (N_2866,In_666,In_1634);
and U2867 (N_2867,In_916,In_2369);
and U2868 (N_2868,In_2305,In_2316);
nand U2869 (N_2869,In_2325,In_2317);
xor U2870 (N_2870,In_1858,In_2339);
and U2871 (N_2871,In_483,In_122);
xnor U2872 (N_2872,In_2239,In_1494);
and U2873 (N_2873,In_433,In_1645);
and U2874 (N_2874,In_2283,In_1366);
or U2875 (N_2875,In_1236,In_1438);
or U2876 (N_2876,In_822,In_1292);
or U2877 (N_2877,In_2022,In_117);
nor U2878 (N_2878,In_1822,In_541);
nand U2879 (N_2879,In_1665,In_335);
nor U2880 (N_2880,In_397,In_377);
nand U2881 (N_2881,In_1007,In_1924);
nor U2882 (N_2882,In_964,In_304);
and U2883 (N_2883,In_396,In_1568);
and U2884 (N_2884,In_794,In_2178);
or U2885 (N_2885,In_1804,In_2031);
nor U2886 (N_2886,In_1373,In_2046);
nand U2887 (N_2887,In_1384,In_2117);
or U2888 (N_2888,In_2154,In_1791);
nand U2889 (N_2889,In_2069,In_364);
nor U2890 (N_2890,In_1498,In_2179);
or U2891 (N_2891,In_1377,In_1060);
or U2892 (N_2892,In_1217,In_1875);
and U2893 (N_2893,In_2100,In_1923);
nand U2894 (N_2894,In_1605,In_1202);
nor U2895 (N_2895,In_1087,In_843);
nor U2896 (N_2896,In_1840,In_1090);
and U2897 (N_2897,In_1223,In_904);
and U2898 (N_2898,In_1443,In_736);
and U2899 (N_2899,In_1707,In_727);
and U2900 (N_2900,In_1704,In_412);
xnor U2901 (N_2901,In_503,In_1102);
nand U2902 (N_2902,In_1505,In_1520);
nor U2903 (N_2903,In_971,In_2181);
nand U2904 (N_2904,In_588,In_2201);
and U2905 (N_2905,In_1753,In_2047);
nand U2906 (N_2906,In_1987,In_1614);
and U2907 (N_2907,In_149,In_587);
or U2908 (N_2908,In_1100,In_1059);
nor U2909 (N_2909,In_530,In_1304);
and U2910 (N_2910,In_924,In_671);
nand U2911 (N_2911,In_953,In_1024);
xor U2912 (N_2912,In_906,In_1917);
or U2913 (N_2913,In_758,In_2476);
nand U2914 (N_2914,In_1449,In_2185);
nor U2915 (N_2915,In_545,In_1035);
or U2916 (N_2916,In_523,In_1348);
and U2917 (N_2917,In_2381,In_1502);
nor U2918 (N_2918,In_1177,In_1196);
nor U2919 (N_2919,In_2048,In_1805);
or U2920 (N_2920,In_1743,In_2491);
nand U2921 (N_2921,In_1401,In_1879);
or U2922 (N_2922,In_2401,In_2379);
and U2923 (N_2923,In_2024,In_1089);
nand U2924 (N_2924,In_1845,In_2204);
xor U2925 (N_2925,In_1104,In_506);
or U2926 (N_2926,In_1819,In_2135);
nand U2927 (N_2927,In_54,In_2376);
xor U2928 (N_2928,In_1478,In_1423);
or U2929 (N_2929,In_336,In_2081);
or U2930 (N_2930,In_1272,In_747);
and U2931 (N_2931,In_8,In_1111);
nand U2932 (N_2932,In_1261,In_2111);
xor U2933 (N_2933,In_1854,In_866);
nand U2934 (N_2934,In_1184,In_1778);
or U2935 (N_2935,In_1553,In_1310);
and U2936 (N_2936,In_1936,In_2156);
and U2937 (N_2937,In_14,In_1532);
nand U2938 (N_2938,In_618,In_567);
xnor U2939 (N_2939,In_1296,In_1565);
or U2940 (N_2940,In_2260,In_391);
and U2941 (N_2941,In_60,In_2302);
xnor U2942 (N_2942,In_1023,In_1859);
nor U2943 (N_2943,In_978,In_518);
or U2944 (N_2944,In_1229,In_2106);
nor U2945 (N_2945,In_2454,In_1987);
nor U2946 (N_2946,In_261,In_1843);
and U2947 (N_2947,In_1521,In_615);
nor U2948 (N_2948,In_1123,In_1755);
or U2949 (N_2949,In_1465,In_163);
and U2950 (N_2950,In_594,In_766);
and U2951 (N_2951,In_1044,In_293);
and U2952 (N_2952,In_1406,In_1011);
and U2953 (N_2953,In_1580,In_2248);
xor U2954 (N_2954,In_331,In_470);
and U2955 (N_2955,In_1302,In_1330);
or U2956 (N_2956,In_335,In_1098);
xor U2957 (N_2957,In_1005,In_2195);
and U2958 (N_2958,In_700,In_2091);
and U2959 (N_2959,In_45,In_93);
nor U2960 (N_2960,In_849,In_538);
and U2961 (N_2961,In_2499,In_305);
and U2962 (N_2962,In_1858,In_1930);
nor U2963 (N_2963,In_1915,In_1237);
and U2964 (N_2964,In_689,In_1648);
and U2965 (N_2965,In_2213,In_2265);
and U2966 (N_2966,In_1873,In_1542);
or U2967 (N_2967,In_873,In_135);
nor U2968 (N_2968,In_53,In_1139);
nor U2969 (N_2969,In_2082,In_2);
or U2970 (N_2970,In_698,In_1208);
or U2971 (N_2971,In_505,In_2019);
or U2972 (N_2972,In_2234,In_1728);
nand U2973 (N_2973,In_94,In_121);
nand U2974 (N_2974,In_934,In_1737);
xor U2975 (N_2975,In_995,In_1740);
xnor U2976 (N_2976,In_132,In_315);
and U2977 (N_2977,In_2022,In_775);
and U2978 (N_2978,In_211,In_1718);
nand U2979 (N_2979,In_1196,In_984);
nor U2980 (N_2980,In_872,In_1552);
or U2981 (N_2981,In_985,In_1245);
and U2982 (N_2982,In_1759,In_35);
nand U2983 (N_2983,In_1844,In_461);
nor U2984 (N_2984,In_171,In_1962);
or U2985 (N_2985,In_949,In_1113);
and U2986 (N_2986,In_2155,In_1175);
and U2987 (N_2987,In_652,In_1441);
and U2988 (N_2988,In_671,In_459);
and U2989 (N_2989,In_2061,In_1516);
nand U2990 (N_2990,In_2287,In_921);
xor U2991 (N_2991,In_1279,In_122);
nor U2992 (N_2992,In_1216,In_2191);
nand U2993 (N_2993,In_248,In_2256);
nand U2994 (N_2994,In_1949,In_417);
or U2995 (N_2995,In_2246,In_542);
or U2996 (N_2996,In_1300,In_2102);
or U2997 (N_2997,In_1133,In_1205);
or U2998 (N_2998,In_1492,In_1216);
nand U2999 (N_2999,In_1765,In_1839);
and U3000 (N_3000,In_2219,In_1576);
or U3001 (N_3001,In_560,In_207);
xor U3002 (N_3002,In_1837,In_1527);
nor U3003 (N_3003,In_1286,In_59);
nor U3004 (N_3004,In_1149,In_291);
xor U3005 (N_3005,In_50,In_1226);
nor U3006 (N_3006,In_1446,In_578);
nand U3007 (N_3007,In_2447,In_2332);
xnor U3008 (N_3008,In_2383,In_1644);
or U3009 (N_3009,In_361,In_647);
or U3010 (N_3010,In_1816,In_852);
and U3011 (N_3011,In_548,In_238);
or U3012 (N_3012,In_1429,In_1017);
and U3013 (N_3013,In_2325,In_1693);
nand U3014 (N_3014,In_1151,In_1084);
or U3015 (N_3015,In_1114,In_875);
or U3016 (N_3016,In_521,In_1184);
and U3017 (N_3017,In_1806,In_1897);
nand U3018 (N_3018,In_848,In_2065);
nor U3019 (N_3019,In_1878,In_2413);
nand U3020 (N_3020,In_758,In_77);
nand U3021 (N_3021,In_507,In_2405);
nor U3022 (N_3022,In_89,In_1834);
nor U3023 (N_3023,In_1209,In_2080);
and U3024 (N_3024,In_1506,In_872);
xnor U3025 (N_3025,In_830,In_2309);
and U3026 (N_3026,In_1960,In_153);
nor U3027 (N_3027,In_1775,In_2168);
xnor U3028 (N_3028,In_2121,In_2300);
nand U3029 (N_3029,In_703,In_393);
nand U3030 (N_3030,In_967,In_1277);
or U3031 (N_3031,In_1938,In_1871);
nor U3032 (N_3032,In_1264,In_476);
or U3033 (N_3033,In_1411,In_1958);
or U3034 (N_3034,In_494,In_1190);
nor U3035 (N_3035,In_2233,In_1541);
nand U3036 (N_3036,In_2386,In_1821);
or U3037 (N_3037,In_22,In_1695);
and U3038 (N_3038,In_1874,In_2384);
and U3039 (N_3039,In_2184,In_859);
nor U3040 (N_3040,In_1366,In_2165);
xnor U3041 (N_3041,In_209,In_1363);
nor U3042 (N_3042,In_1503,In_1476);
nand U3043 (N_3043,In_893,In_1582);
nor U3044 (N_3044,In_1109,In_374);
nand U3045 (N_3045,In_82,In_2062);
and U3046 (N_3046,In_822,In_1316);
or U3047 (N_3047,In_1613,In_1717);
xnor U3048 (N_3048,In_1813,In_962);
or U3049 (N_3049,In_1604,In_453);
xnor U3050 (N_3050,In_610,In_1717);
nand U3051 (N_3051,In_862,In_579);
nor U3052 (N_3052,In_1906,In_1966);
or U3053 (N_3053,In_1311,In_1707);
nor U3054 (N_3054,In_1692,In_1815);
and U3055 (N_3055,In_1434,In_1469);
xnor U3056 (N_3056,In_2152,In_1225);
or U3057 (N_3057,In_1711,In_1511);
and U3058 (N_3058,In_506,In_942);
xor U3059 (N_3059,In_2064,In_52);
or U3060 (N_3060,In_1392,In_155);
nand U3061 (N_3061,In_1201,In_768);
and U3062 (N_3062,In_1635,In_1474);
nand U3063 (N_3063,In_478,In_1008);
nor U3064 (N_3064,In_305,In_1102);
or U3065 (N_3065,In_1097,In_585);
or U3066 (N_3066,In_2442,In_711);
and U3067 (N_3067,In_1688,In_969);
nor U3068 (N_3068,In_1097,In_1105);
nand U3069 (N_3069,In_2104,In_577);
nand U3070 (N_3070,In_1153,In_1463);
xnor U3071 (N_3071,In_1867,In_1252);
nor U3072 (N_3072,In_0,In_928);
xnor U3073 (N_3073,In_1462,In_2094);
or U3074 (N_3074,In_9,In_684);
or U3075 (N_3075,In_2094,In_1342);
nand U3076 (N_3076,In_2054,In_394);
nand U3077 (N_3077,In_2027,In_48);
xor U3078 (N_3078,In_1689,In_2080);
or U3079 (N_3079,In_2103,In_2464);
or U3080 (N_3080,In_685,In_1872);
nor U3081 (N_3081,In_274,In_172);
nor U3082 (N_3082,In_1020,In_1946);
nand U3083 (N_3083,In_261,In_1865);
and U3084 (N_3084,In_685,In_840);
nor U3085 (N_3085,In_2063,In_155);
nand U3086 (N_3086,In_1483,In_1003);
nor U3087 (N_3087,In_1606,In_1584);
nor U3088 (N_3088,In_503,In_2351);
nand U3089 (N_3089,In_542,In_1988);
nor U3090 (N_3090,In_1738,In_2402);
nand U3091 (N_3091,In_663,In_2220);
xnor U3092 (N_3092,In_2237,In_1540);
and U3093 (N_3093,In_994,In_1125);
and U3094 (N_3094,In_307,In_1000);
nor U3095 (N_3095,In_2170,In_546);
and U3096 (N_3096,In_2444,In_1790);
nor U3097 (N_3097,In_1449,In_1537);
or U3098 (N_3098,In_683,In_2155);
nand U3099 (N_3099,In_906,In_343);
xnor U3100 (N_3100,In_2297,In_61);
nor U3101 (N_3101,In_1568,In_2041);
nand U3102 (N_3102,In_2419,In_2352);
nand U3103 (N_3103,In_355,In_1993);
or U3104 (N_3104,In_1547,In_837);
or U3105 (N_3105,In_1538,In_672);
nor U3106 (N_3106,In_610,In_1809);
or U3107 (N_3107,In_2456,In_2324);
nand U3108 (N_3108,In_1445,In_1996);
xnor U3109 (N_3109,In_2005,In_1528);
and U3110 (N_3110,In_20,In_69);
and U3111 (N_3111,In_10,In_2171);
nand U3112 (N_3112,In_1969,In_2444);
nor U3113 (N_3113,In_1133,In_2378);
nor U3114 (N_3114,In_1718,In_480);
and U3115 (N_3115,In_2376,In_939);
nand U3116 (N_3116,In_1856,In_2406);
nand U3117 (N_3117,In_27,In_944);
nand U3118 (N_3118,In_820,In_2143);
or U3119 (N_3119,In_1510,In_584);
nand U3120 (N_3120,In_1694,In_155);
and U3121 (N_3121,In_242,In_1737);
nor U3122 (N_3122,In_434,In_1421);
nor U3123 (N_3123,In_320,In_782);
nor U3124 (N_3124,In_172,In_2234);
nand U3125 (N_3125,In_481,In_77);
nor U3126 (N_3126,In_1239,In_1215);
or U3127 (N_3127,In_2164,In_2277);
nor U3128 (N_3128,In_67,In_584);
nor U3129 (N_3129,In_800,In_571);
and U3130 (N_3130,In_588,In_198);
nand U3131 (N_3131,In_764,In_207);
and U3132 (N_3132,In_60,In_1498);
and U3133 (N_3133,In_200,In_1857);
nor U3134 (N_3134,In_286,In_1895);
or U3135 (N_3135,In_2366,In_261);
nand U3136 (N_3136,In_1345,In_1823);
and U3137 (N_3137,In_546,In_1370);
or U3138 (N_3138,In_904,In_1139);
nor U3139 (N_3139,In_1705,In_11);
nand U3140 (N_3140,In_1903,In_1334);
or U3141 (N_3141,In_481,In_824);
nor U3142 (N_3142,In_1234,In_1179);
nor U3143 (N_3143,In_1888,In_516);
and U3144 (N_3144,In_1123,In_2273);
or U3145 (N_3145,In_1590,In_2078);
nor U3146 (N_3146,In_2305,In_838);
nand U3147 (N_3147,In_99,In_2049);
nor U3148 (N_3148,In_1639,In_2120);
xnor U3149 (N_3149,In_368,In_1537);
or U3150 (N_3150,In_1039,In_425);
or U3151 (N_3151,In_482,In_2416);
and U3152 (N_3152,In_1179,In_1656);
nand U3153 (N_3153,In_909,In_23);
xor U3154 (N_3154,In_1032,In_2154);
or U3155 (N_3155,In_457,In_891);
or U3156 (N_3156,In_259,In_657);
or U3157 (N_3157,In_1134,In_722);
and U3158 (N_3158,In_1834,In_838);
nor U3159 (N_3159,In_912,In_1505);
nand U3160 (N_3160,In_2060,In_370);
nor U3161 (N_3161,In_2288,In_1927);
nand U3162 (N_3162,In_2082,In_1362);
nor U3163 (N_3163,In_365,In_1774);
nor U3164 (N_3164,In_1970,In_1425);
xnor U3165 (N_3165,In_2354,In_2343);
nor U3166 (N_3166,In_659,In_1014);
nand U3167 (N_3167,In_1277,In_1505);
and U3168 (N_3168,In_1339,In_1298);
and U3169 (N_3169,In_129,In_1949);
nand U3170 (N_3170,In_1783,In_830);
nand U3171 (N_3171,In_2340,In_1058);
nand U3172 (N_3172,In_93,In_1713);
nor U3173 (N_3173,In_2283,In_307);
or U3174 (N_3174,In_1952,In_1116);
nor U3175 (N_3175,In_2135,In_1006);
nor U3176 (N_3176,In_153,In_906);
or U3177 (N_3177,In_1188,In_218);
and U3178 (N_3178,In_1448,In_2121);
and U3179 (N_3179,In_2177,In_974);
or U3180 (N_3180,In_2466,In_433);
or U3181 (N_3181,In_1046,In_2369);
nor U3182 (N_3182,In_880,In_2340);
or U3183 (N_3183,In_685,In_1753);
and U3184 (N_3184,In_2336,In_80);
nor U3185 (N_3185,In_408,In_1119);
or U3186 (N_3186,In_1209,In_852);
nand U3187 (N_3187,In_1619,In_1061);
xnor U3188 (N_3188,In_1731,In_2025);
nor U3189 (N_3189,In_2377,In_329);
or U3190 (N_3190,In_1508,In_1044);
nand U3191 (N_3191,In_2022,In_1362);
nand U3192 (N_3192,In_1736,In_1282);
and U3193 (N_3193,In_1612,In_614);
and U3194 (N_3194,In_2134,In_1463);
nand U3195 (N_3195,In_2077,In_2383);
or U3196 (N_3196,In_2402,In_791);
nor U3197 (N_3197,In_277,In_2281);
nand U3198 (N_3198,In_2289,In_541);
nor U3199 (N_3199,In_2317,In_2239);
or U3200 (N_3200,In_732,In_1503);
xor U3201 (N_3201,In_2333,In_2417);
nor U3202 (N_3202,In_669,In_685);
nand U3203 (N_3203,In_470,In_682);
nor U3204 (N_3204,In_905,In_701);
xor U3205 (N_3205,In_1934,In_2010);
nor U3206 (N_3206,In_694,In_1381);
or U3207 (N_3207,In_1976,In_2093);
or U3208 (N_3208,In_480,In_2219);
nand U3209 (N_3209,In_98,In_1593);
and U3210 (N_3210,In_1775,In_1128);
nand U3211 (N_3211,In_1197,In_18);
nand U3212 (N_3212,In_385,In_2416);
nor U3213 (N_3213,In_2185,In_593);
and U3214 (N_3214,In_1339,In_1445);
xnor U3215 (N_3215,In_1085,In_1555);
and U3216 (N_3216,In_627,In_722);
nand U3217 (N_3217,In_1987,In_1996);
or U3218 (N_3218,In_1867,In_190);
nand U3219 (N_3219,In_2011,In_2197);
or U3220 (N_3220,In_1949,In_775);
nor U3221 (N_3221,In_1759,In_1286);
nor U3222 (N_3222,In_1368,In_1879);
nand U3223 (N_3223,In_1727,In_2032);
nand U3224 (N_3224,In_1153,In_609);
and U3225 (N_3225,In_292,In_2342);
nand U3226 (N_3226,In_1725,In_2454);
xor U3227 (N_3227,In_341,In_463);
xnor U3228 (N_3228,In_1368,In_1581);
nor U3229 (N_3229,In_1819,In_1975);
nor U3230 (N_3230,In_1247,In_753);
nor U3231 (N_3231,In_2423,In_498);
nor U3232 (N_3232,In_1550,In_671);
or U3233 (N_3233,In_449,In_413);
nand U3234 (N_3234,In_1233,In_1084);
nand U3235 (N_3235,In_1217,In_1322);
and U3236 (N_3236,In_1126,In_2497);
or U3237 (N_3237,In_1903,In_2133);
or U3238 (N_3238,In_396,In_440);
nand U3239 (N_3239,In_898,In_1239);
or U3240 (N_3240,In_2080,In_2451);
and U3241 (N_3241,In_449,In_1366);
nand U3242 (N_3242,In_111,In_1220);
or U3243 (N_3243,In_1791,In_1947);
and U3244 (N_3244,In_952,In_1893);
nand U3245 (N_3245,In_1861,In_1674);
and U3246 (N_3246,In_589,In_1519);
nand U3247 (N_3247,In_253,In_32);
and U3248 (N_3248,In_2100,In_505);
and U3249 (N_3249,In_792,In_1226);
or U3250 (N_3250,In_1770,In_2005);
nand U3251 (N_3251,In_2419,In_2005);
nor U3252 (N_3252,In_1876,In_1307);
and U3253 (N_3253,In_1015,In_573);
nor U3254 (N_3254,In_971,In_728);
nand U3255 (N_3255,In_2087,In_582);
nand U3256 (N_3256,In_2190,In_1383);
nor U3257 (N_3257,In_1267,In_2299);
nor U3258 (N_3258,In_1464,In_2455);
and U3259 (N_3259,In_1418,In_358);
or U3260 (N_3260,In_2436,In_1735);
or U3261 (N_3261,In_1393,In_605);
nor U3262 (N_3262,In_2423,In_1676);
or U3263 (N_3263,In_2125,In_1043);
nor U3264 (N_3264,In_379,In_757);
xor U3265 (N_3265,In_376,In_1980);
nor U3266 (N_3266,In_884,In_2126);
and U3267 (N_3267,In_197,In_193);
and U3268 (N_3268,In_1192,In_709);
xor U3269 (N_3269,In_10,In_1150);
and U3270 (N_3270,In_1168,In_655);
nand U3271 (N_3271,In_721,In_1241);
or U3272 (N_3272,In_574,In_1969);
and U3273 (N_3273,In_961,In_980);
and U3274 (N_3274,In_1722,In_1458);
xnor U3275 (N_3275,In_2228,In_1323);
nor U3276 (N_3276,In_1320,In_173);
xor U3277 (N_3277,In_261,In_1326);
nand U3278 (N_3278,In_259,In_2025);
xnor U3279 (N_3279,In_25,In_1704);
nor U3280 (N_3280,In_966,In_863);
nor U3281 (N_3281,In_881,In_1579);
xnor U3282 (N_3282,In_244,In_1847);
nand U3283 (N_3283,In_1789,In_1853);
nand U3284 (N_3284,In_1675,In_1469);
or U3285 (N_3285,In_2205,In_131);
and U3286 (N_3286,In_2244,In_2396);
and U3287 (N_3287,In_1007,In_1264);
and U3288 (N_3288,In_2094,In_2482);
and U3289 (N_3289,In_1804,In_856);
and U3290 (N_3290,In_434,In_802);
nor U3291 (N_3291,In_1506,In_1959);
and U3292 (N_3292,In_293,In_1638);
xnor U3293 (N_3293,In_807,In_324);
or U3294 (N_3294,In_1469,In_1501);
or U3295 (N_3295,In_479,In_388);
nor U3296 (N_3296,In_1115,In_1781);
and U3297 (N_3297,In_512,In_98);
or U3298 (N_3298,In_2040,In_1695);
xnor U3299 (N_3299,In_1640,In_861);
and U3300 (N_3300,In_2301,In_32);
and U3301 (N_3301,In_2204,In_847);
and U3302 (N_3302,In_370,In_1364);
nor U3303 (N_3303,In_8,In_846);
xnor U3304 (N_3304,In_2288,In_1532);
xnor U3305 (N_3305,In_2416,In_372);
or U3306 (N_3306,In_735,In_292);
nor U3307 (N_3307,In_2410,In_811);
nor U3308 (N_3308,In_2200,In_1718);
nor U3309 (N_3309,In_2024,In_2279);
nand U3310 (N_3310,In_1792,In_2462);
nand U3311 (N_3311,In_1413,In_1782);
and U3312 (N_3312,In_2069,In_1934);
xnor U3313 (N_3313,In_1701,In_789);
nor U3314 (N_3314,In_17,In_2066);
or U3315 (N_3315,In_613,In_776);
or U3316 (N_3316,In_1829,In_790);
nand U3317 (N_3317,In_183,In_2392);
or U3318 (N_3318,In_2284,In_1851);
nor U3319 (N_3319,In_321,In_705);
nor U3320 (N_3320,In_734,In_1300);
or U3321 (N_3321,In_564,In_2414);
nand U3322 (N_3322,In_1199,In_372);
nand U3323 (N_3323,In_1024,In_123);
or U3324 (N_3324,In_906,In_991);
or U3325 (N_3325,In_1791,In_749);
or U3326 (N_3326,In_1879,In_1228);
nor U3327 (N_3327,In_641,In_2342);
nor U3328 (N_3328,In_1411,In_1550);
and U3329 (N_3329,In_1302,In_39);
nor U3330 (N_3330,In_1909,In_2176);
and U3331 (N_3331,In_242,In_1312);
nand U3332 (N_3332,In_540,In_1006);
or U3333 (N_3333,In_1605,In_114);
nor U3334 (N_3334,In_1439,In_1520);
xnor U3335 (N_3335,In_1316,In_669);
or U3336 (N_3336,In_2162,In_1422);
nand U3337 (N_3337,In_974,In_617);
nor U3338 (N_3338,In_325,In_2071);
nor U3339 (N_3339,In_1836,In_1763);
nor U3340 (N_3340,In_642,In_496);
nor U3341 (N_3341,In_1105,In_2103);
nor U3342 (N_3342,In_256,In_668);
or U3343 (N_3343,In_2414,In_1291);
and U3344 (N_3344,In_207,In_2341);
nor U3345 (N_3345,In_2256,In_445);
or U3346 (N_3346,In_347,In_1308);
and U3347 (N_3347,In_1173,In_1105);
or U3348 (N_3348,In_1805,In_2107);
xor U3349 (N_3349,In_257,In_781);
or U3350 (N_3350,In_1691,In_604);
nor U3351 (N_3351,In_2181,In_986);
nand U3352 (N_3352,In_209,In_1961);
and U3353 (N_3353,In_154,In_2280);
nor U3354 (N_3354,In_47,In_180);
nand U3355 (N_3355,In_575,In_1625);
or U3356 (N_3356,In_330,In_2168);
nor U3357 (N_3357,In_128,In_2351);
and U3358 (N_3358,In_783,In_316);
nand U3359 (N_3359,In_1257,In_121);
nand U3360 (N_3360,In_777,In_2234);
xor U3361 (N_3361,In_99,In_2062);
xor U3362 (N_3362,In_2310,In_2080);
or U3363 (N_3363,In_2351,In_1823);
nor U3364 (N_3364,In_1233,In_111);
or U3365 (N_3365,In_590,In_2239);
nor U3366 (N_3366,In_2217,In_1357);
or U3367 (N_3367,In_1717,In_1168);
and U3368 (N_3368,In_2214,In_2336);
xor U3369 (N_3369,In_1721,In_1249);
xnor U3370 (N_3370,In_1470,In_1047);
or U3371 (N_3371,In_2197,In_378);
nand U3372 (N_3372,In_1685,In_1079);
nor U3373 (N_3373,In_1161,In_1249);
or U3374 (N_3374,In_1370,In_462);
and U3375 (N_3375,In_2212,In_491);
nor U3376 (N_3376,In_1635,In_1997);
or U3377 (N_3377,In_681,In_29);
nand U3378 (N_3378,In_93,In_2439);
and U3379 (N_3379,In_237,In_1174);
nand U3380 (N_3380,In_2319,In_102);
or U3381 (N_3381,In_616,In_1576);
nand U3382 (N_3382,In_64,In_2000);
nand U3383 (N_3383,In_708,In_1869);
nand U3384 (N_3384,In_77,In_1803);
nand U3385 (N_3385,In_2223,In_2413);
or U3386 (N_3386,In_1427,In_166);
nand U3387 (N_3387,In_2250,In_1059);
xnor U3388 (N_3388,In_349,In_676);
and U3389 (N_3389,In_2210,In_793);
nor U3390 (N_3390,In_452,In_772);
and U3391 (N_3391,In_2105,In_855);
or U3392 (N_3392,In_1151,In_793);
xnor U3393 (N_3393,In_330,In_1357);
or U3394 (N_3394,In_1279,In_1611);
and U3395 (N_3395,In_1971,In_1309);
and U3396 (N_3396,In_1825,In_1693);
nor U3397 (N_3397,In_841,In_1210);
and U3398 (N_3398,In_2366,In_586);
nand U3399 (N_3399,In_1367,In_600);
nand U3400 (N_3400,In_977,In_1868);
xnor U3401 (N_3401,In_183,In_2464);
or U3402 (N_3402,In_805,In_1777);
or U3403 (N_3403,In_1274,In_715);
xor U3404 (N_3404,In_2181,In_1590);
nand U3405 (N_3405,In_89,In_1121);
or U3406 (N_3406,In_2342,In_537);
and U3407 (N_3407,In_1334,In_2089);
and U3408 (N_3408,In_2296,In_1349);
or U3409 (N_3409,In_1361,In_1221);
and U3410 (N_3410,In_2464,In_1392);
and U3411 (N_3411,In_228,In_401);
or U3412 (N_3412,In_1423,In_2095);
nor U3413 (N_3413,In_698,In_270);
nand U3414 (N_3414,In_1750,In_2231);
or U3415 (N_3415,In_780,In_884);
or U3416 (N_3416,In_2368,In_1727);
nand U3417 (N_3417,In_427,In_1427);
nand U3418 (N_3418,In_2148,In_951);
nor U3419 (N_3419,In_1158,In_1809);
xnor U3420 (N_3420,In_1464,In_2373);
nand U3421 (N_3421,In_2158,In_592);
nor U3422 (N_3422,In_1091,In_1850);
nand U3423 (N_3423,In_810,In_2261);
and U3424 (N_3424,In_952,In_1310);
or U3425 (N_3425,In_2212,In_570);
nand U3426 (N_3426,In_1791,In_1100);
and U3427 (N_3427,In_2029,In_19);
or U3428 (N_3428,In_671,In_2402);
xor U3429 (N_3429,In_12,In_1820);
or U3430 (N_3430,In_1453,In_363);
nand U3431 (N_3431,In_705,In_1551);
xnor U3432 (N_3432,In_516,In_885);
xor U3433 (N_3433,In_717,In_2379);
and U3434 (N_3434,In_2203,In_411);
nor U3435 (N_3435,In_347,In_677);
or U3436 (N_3436,In_204,In_751);
xnor U3437 (N_3437,In_1034,In_239);
nand U3438 (N_3438,In_1768,In_1653);
nand U3439 (N_3439,In_559,In_1365);
or U3440 (N_3440,In_1448,In_838);
nor U3441 (N_3441,In_107,In_2148);
nand U3442 (N_3442,In_62,In_2359);
xnor U3443 (N_3443,In_1124,In_974);
nand U3444 (N_3444,In_355,In_998);
nor U3445 (N_3445,In_410,In_1583);
nor U3446 (N_3446,In_816,In_1008);
and U3447 (N_3447,In_497,In_1521);
nand U3448 (N_3448,In_1282,In_64);
nor U3449 (N_3449,In_1618,In_703);
xnor U3450 (N_3450,In_26,In_333);
xor U3451 (N_3451,In_648,In_764);
xnor U3452 (N_3452,In_1011,In_653);
or U3453 (N_3453,In_1796,In_791);
nand U3454 (N_3454,In_239,In_1871);
or U3455 (N_3455,In_2053,In_1141);
and U3456 (N_3456,In_2192,In_1300);
and U3457 (N_3457,In_2170,In_1372);
nand U3458 (N_3458,In_2096,In_1291);
nor U3459 (N_3459,In_1508,In_1573);
nor U3460 (N_3460,In_1531,In_1952);
nand U3461 (N_3461,In_2313,In_1280);
nor U3462 (N_3462,In_1344,In_1898);
nand U3463 (N_3463,In_2189,In_1884);
nand U3464 (N_3464,In_21,In_575);
nor U3465 (N_3465,In_1381,In_1823);
nand U3466 (N_3466,In_1814,In_1233);
and U3467 (N_3467,In_2128,In_1501);
nor U3468 (N_3468,In_679,In_113);
xnor U3469 (N_3469,In_331,In_643);
nand U3470 (N_3470,In_720,In_1163);
nand U3471 (N_3471,In_346,In_368);
and U3472 (N_3472,In_1970,In_599);
or U3473 (N_3473,In_527,In_1022);
xor U3474 (N_3474,In_726,In_344);
nor U3475 (N_3475,In_1116,In_1795);
nand U3476 (N_3476,In_614,In_1057);
nor U3477 (N_3477,In_574,In_255);
and U3478 (N_3478,In_1450,In_106);
and U3479 (N_3479,In_899,In_2421);
nand U3480 (N_3480,In_1316,In_419);
and U3481 (N_3481,In_1355,In_1405);
nand U3482 (N_3482,In_1675,In_1634);
nand U3483 (N_3483,In_303,In_993);
or U3484 (N_3484,In_1564,In_2412);
or U3485 (N_3485,In_1356,In_2362);
or U3486 (N_3486,In_1818,In_382);
nor U3487 (N_3487,In_2329,In_1095);
or U3488 (N_3488,In_1673,In_12);
nand U3489 (N_3489,In_1360,In_1402);
xnor U3490 (N_3490,In_243,In_1647);
nand U3491 (N_3491,In_386,In_1363);
and U3492 (N_3492,In_1945,In_1813);
and U3493 (N_3493,In_1388,In_2243);
and U3494 (N_3494,In_1570,In_1433);
or U3495 (N_3495,In_1507,In_94);
and U3496 (N_3496,In_2397,In_1051);
nor U3497 (N_3497,In_2477,In_1328);
and U3498 (N_3498,In_2368,In_2466);
nand U3499 (N_3499,In_72,In_385);
or U3500 (N_3500,In_1594,In_2246);
or U3501 (N_3501,In_2344,In_1476);
nor U3502 (N_3502,In_2489,In_1891);
nand U3503 (N_3503,In_2139,In_413);
nor U3504 (N_3504,In_2156,In_1856);
or U3505 (N_3505,In_1030,In_1693);
nor U3506 (N_3506,In_351,In_1004);
nor U3507 (N_3507,In_956,In_2468);
nand U3508 (N_3508,In_2265,In_1530);
nor U3509 (N_3509,In_2337,In_735);
xor U3510 (N_3510,In_1344,In_904);
nand U3511 (N_3511,In_763,In_816);
nor U3512 (N_3512,In_551,In_2022);
nand U3513 (N_3513,In_187,In_884);
nor U3514 (N_3514,In_2245,In_36);
or U3515 (N_3515,In_66,In_2030);
or U3516 (N_3516,In_1064,In_2123);
or U3517 (N_3517,In_2192,In_879);
xor U3518 (N_3518,In_1844,In_1124);
nand U3519 (N_3519,In_103,In_2219);
or U3520 (N_3520,In_913,In_2048);
nand U3521 (N_3521,In_1199,In_710);
xnor U3522 (N_3522,In_2466,In_1944);
and U3523 (N_3523,In_263,In_612);
nor U3524 (N_3524,In_1488,In_1819);
nor U3525 (N_3525,In_1461,In_262);
or U3526 (N_3526,In_767,In_2342);
and U3527 (N_3527,In_987,In_137);
nand U3528 (N_3528,In_1050,In_473);
or U3529 (N_3529,In_1874,In_286);
xor U3530 (N_3530,In_68,In_2094);
and U3531 (N_3531,In_2191,In_1896);
nand U3532 (N_3532,In_2312,In_1740);
or U3533 (N_3533,In_628,In_1838);
nor U3534 (N_3534,In_1003,In_1146);
and U3535 (N_3535,In_1474,In_1154);
nand U3536 (N_3536,In_1799,In_371);
or U3537 (N_3537,In_1489,In_2007);
or U3538 (N_3538,In_1765,In_371);
nor U3539 (N_3539,In_673,In_1058);
or U3540 (N_3540,In_853,In_90);
nand U3541 (N_3541,In_1488,In_592);
nand U3542 (N_3542,In_1839,In_327);
nand U3543 (N_3543,In_207,In_1502);
and U3544 (N_3544,In_1439,In_784);
nand U3545 (N_3545,In_2235,In_430);
nor U3546 (N_3546,In_2435,In_1796);
or U3547 (N_3547,In_1951,In_1486);
nand U3548 (N_3548,In_2223,In_1792);
and U3549 (N_3549,In_164,In_2496);
nand U3550 (N_3550,In_2157,In_2392);
nand U3551 (N_3551,In_2222,In_1004);
or U3552 (N_3552,In_1355,In_2280);
nand U3553 (N_3553,In_2220,In_64);
nand U3554 (N_3554,In_1638,In_965);
nor U3555 (N_3555,In_902,In_882);
and U3556 (N_3556,In_1506,In_597);
or U3557 (N_3557,In_1231,In_1551);
nor U3558 (N_3558,In_1942,In_1416);
or U3559 (N_3559,In_2495,In_836);
or U3560 (N_3560,In_1101,In_2025);
and U3561 (N_3561,In_1802,In_31);
or U3562 (N_3562,In_1096,In_1412);
and U3563 (N_3563,In_1244,In_1580);
nor U3564 (N_3564,In_1599,In_954);
or U3565 (N_3565,In_2183,In_2313);
xor U3566 (N_3566,In_2077,In_365);
and U3567 (N_3567,In_1510,In_1672);
and U3568 (N_3568,In_690,In_799);
nand U3569 (N_3569,In_2331,In_1713);
or U3570 (N_3570,In_312,In_2153);
nor U3571 (N_3571,In_2025,In_2097);
nand U3572 (N_3572,In_1324,In_975);
or U3573 (N_3573,In_1725,In_362);
nand U3574 (N_3574,In_275,In_2227);
or U3575 (N_3575,In_1825,In_1101);
nand U3576 (N_3576,In_894,In_1230);
xnor U3577 (N_3577,In_2181,In_31);
nand U3578 (N_3578,In_1689,In_780);
xor U3579 (N_3579,In_1303,In_1267);
and U3580 (N_3580,In_1373,In_1489);
nand U3581 (N_3581,In_1508,In_274);
nand U3582 (N_3582,In_2401,In_1384);
and U3583 (N_3583,In_2230,In_2158);
xnor U3584 (N_3584,In_289,In_475);
nor U3585 (N_3585,In_618,In_2421);
or U3586 (N_3586,In_2193,In_588);
nand U3587 (N_3587,In_1840,In_0);
nand U3588 (N_3588,In_293,In_1569);
xnor U3589 (N_3589,In_1668,In_828);
xor U3590 (N_3590,In_1734,In_948);
xnor U3591 (N_3591,In_1213,In_1385);
xnor U3592 (N_3592,In_2456,In_111);
or U3593 (N_3593,In_2412,In_149);
nand U3594 (N_3594,In_491,In_423);
nor U3595 (N_3595,In_1117,In_2049);
nand U3596 (N_3596,In_902,In_1502);
nand U3597 (N_3597,In_445,In_1221);
and U3598 (N_3598,In_944,In_1820);
and U3599 (N_3599,In_2159,In_183);
nand U3600 (N_3600,In_1042,In_2088);
nor U3601 (N_3601,In_1620,In_974);
xnor U3602 (N_3602,In_2136,In_2005);
xnor U3603 (N_3603,In_1818,In_1590);
nand U3604 (N_3604,In_1743,In_1856);
nor U3605 (N_3605,In_214,In_1691);
nand U3606 (N_3606,In_1036,In_1153);
or U3607 (N_3607,In_1149,In_25);
nand U3608 (N_3608,In_1847,In_1263);
and U3609 (N_3609,In_494,In_2423);
and U3610 (N_3610,In_1508,In_1829);
nor U3611 (N_3611,In_14,In_1122);
nor U3612 (N_3612,In_740,In_696);
nand U3613 (N_3613,In_1932,In_1023);
nor U3614 (N_3614,In_1430,In_2055);
nor U3615 (N_3615,In_2079,In_1104);
nor U3616 (N_3616,In_764,In_2161);
nand U3617 (N_3617,In_642,In_608);
and U3618 (N_3618,In_542,In_937);
nand U3619 (N_3619,In_399,In_1696);
and U3620 (N_3620,In_2127,In_300);
nand U3621 (N_3621,In_1155,In_978);
or U3622 (N_3622,In_1572,In_2247);
or U3623 (N_3623,In_389,In_1251);
nand U3624 (N_3624,In_1820,In_1967);
nor U3625 (N_3625,In_1383,In_1388);
xor U3626 (N_3626,In_1790,In_1623);
nor U3627 (N_3627,In_1463,In_2077);
xor U3628 (N_3628,In_620,In_308);
nor U3629 (N_3629,In_1440,In_1567);
and U3630 (N_3630,In_1539,In_1793);
or U3631 (N_3631,In_402,In_1159);
nor U3632 (N_3632,In_248,In_2374);
and U3633 (N_3633,In_1779,In_839);
nor U3634 (N_3634,In_131,In_1975);
nand U3635 (N_3635,In_2299,In_1114);
or U3636 (N_3636,In_185,In_1479);
nand U3637 (N_3637,In_1281,In_1383);
nor U3638 (N_3638,In_737,In_812);
or U3639 (N_3639,In_503,In_1096);
or U3640 (N_3640,In_1217,In_1590);
nand U3641 (N_3641,In_1414,In_29);
nand U3642 (N_3642,In_487,In_1182);
nand U3643 (N_3643,In_933,In_1346);
nor U3644 (N_3644,In_2303,In_434);
or U3645 (N_3645,In_631,In_1788);
and U3646 (N_3646,In_1452,In_2106);
nand U3647 (N_3647,In_715,In_2491);
nor U3648 (N_3648,In_1995,In_2249);
or U3649 (N_3649,In_95,In_1354);
and U3650 (N_3650,In_151,In_1234);
nor U3651 (N_3651,In_1390,In_2041);
and U3652 (N_3652,In_479,In_580);
or U3653 (N_3653,In_778,In_80);
or U3654 (N_3654,In_1885,In_2462);
or U3655 (N_3655,In_2057,In_1435);
nor U3656 (N_3656,In_1782,In_1327);
xnor U3657 (N_3657,In_909,In_1637);
and U3658 (N_3658,In_1408,In_1029);
or U3659 (N_3659,In_1299,In_758);
nand U3660 (N_3660,In_2472,In_2257);
and U3661 (N_3661,In_195,In_1460);
and U3662 (N_3662,In_1161,In_192);
and U3663 (N_3663,In_870,In_232);
nor U3664 (N_3664,In_1213,In_2119);
xnor U3665 (N_3665,In_767,In_2147);
nand U3666 (N_3666,In_1475,In_1303);
nand U3667 (N_3667,In_1937,In_2447);
xor U3668 (N_3668,In_9,In_177);
or U3669 (N_3669,In_287,In_1877);
nand U3670 (N_3670,In_169,In_424);
and U3671 (N_3671,In_1097,In_2188);
xor U3672 (N_3672,In_1824,In_1266);
nand U3673 (N_3673,In_7,In_624);
or U3674 (N_3674,In_301,In_1488);
and U3675 (N_3675,In_1112,In_1533);
nor U3676 (N_3676,In_46,In_634);
nand U3677 (N_3677,In_880,In_609);
and U3678 (N_3678,In_1783,In_1850);
and U3679 (N_3679,In_275,In_1736);
or U3680 (N_3680,In_2265,In_437);
or U3681 (N_3681,In_1069,In_1266);
nor U3682 (N_3682,In_2410,In_349);
and U3683 (N_3683,In_968,In_1730);
nand U3684 (N_3684,In_1222,In_1376);
and U3685 (N_3685,In_2327,In_361);
xor U3686 (N_3686,In_167,In_843);
nor U3687 (N_3687,In_2409,In_1181);
nor U3688 (N_3688,In_81,In_1949);
nor U3689 (N_3689,In_2040,In_1401);
or U3690 (N_3690,In_2447,In_2242);
or U3691 (N_3691,In_2278,In_933);
nand U3692 (N_3692,In_783,In_1485);
nand U3693 (N_3693,In_889,In_142);
and U3694 (N_3694,In_1967,In_2060);
and U3695 (N_3695,In_579,In_2131);
nand U3696 (N_3696,In_1290,In_731);
and U3697 (N_3697,In_103,In_123);
or U3698 (N_3698,In_367,In_218);
or U3699 (N_3699,In_887,In_2272);
or U3700 (N_3700,In_1365,In_749);
nand U3701 (N_3701,In_918,In_2027);
nor U3702 (N_3702,In_2348,In_2326);
or U3703 (N_3703,In_1867,In_1349);
nor U3704 (N_3704,In_2273,In_512);
and U3705 (N_3705,In_258,In_1076);
and U3706 (N_3706,In_510,In_1777);
nand U3707 (N_3707,In_1424,In_1106);
nor U3708 (N_3708,In_2389,In_1418);
or U3709 (N_3709,In_2327,In_564);
nor U3710 (N_3710,In_590,In_1414);
nor U3711 (N_3711,In_145,In_2167);
and U3712 (N_3712,In_272,In_1329);
and U3713 (N_3713,In_2190,In_1083);
nand U3714 (N_3714,In_694,In_742);
xnor U3715 (N_3715,In_1672,In_1732);
or U3716 (N_3716,In_2075,In_2016);
nor U3717 (N_3717,In_948,In_338);
and U3718 (N_3718,In_957,In_637);
or U3719 (N_3719,In_1353,In_491);
xnor U3720 (N_3720,In_1272,In_1074);
or U3721 (N_3721,In_2013,In_277);
nand U3722 (N_3722,In_2226,In_1508);
nand U3723 (N_3723,In_1049,In_251);
nor U3724 (N_3724,In_11,In_2022);
nand U3725 (N_3725,In_1549,In_2083);
or U3726 (N_3726,In_2405,In_1283);
nor U3727 (N_3727,In_2081,In_192);
nand U3728 (N_3728,In_90,In_1055);
nor U3729 (N_3729,In_2369,In_871);
and U3730 (N_3730,In_1011,In_505);
or U3731 (N_3731,In_1253,In_1327);
nand U3732 (N_3732,In_2436,In_1801);
or U3733 (N_3733,In_238,In_1988);
nand U3734 (N_3734,In_2357,In_1552);
or U3735 (N_3735,In_491,In_1229);
nand U3736 (N_3736,In_2161,In_2299);
nor U3737 (N_3737,In_1522,In_1477);
or U3738 (N_3738,In_1913,In_1557);
and U3739 (N_3739,In_2007,In_779);
and U3740 (N_3740,In_1878,In_959);
and U3741 (N_3741,In_1169,In_1464);
nor U3742 (N_3742,In_2262,In_185);
xor U3743 (N_3743,In_890,In_2150);
nand U3744 (N_3744,In_2441,In_289);
nand U3745 (N_3745,In_716,In_1930);
nor U3746 (N_3746,In_1588,In_1638);
and U3747 (N_3747,In_1158,In_1573);
nor U3748 (N_3748,In_1274,In_1198);
nor U3749 (N_3749,In_725,In_634);
and U3750 (N_3750,In_796,In_1901);
nor U3751 (N_3751,In_2379,In_1679);
and U3752 (N_3752,In_2420,In_1282);
nand U3753 (N_3753,In_2190,In_1869);
xor U3754 (N_3754,In_722,In_516);
or U3755 (N_3755,In_1476,In_1882);
xnor U3756 (N_3756,In_1620,In_2498);
and U3757 (N_3757,In_2161,In_1983);
and U3758 (N_3758,In_1464,In_281);
or U3759 (N_3759,In_1753,In_882);
xnor U3760 (N_3760,In_2317,In_1391);
xnor U3761 (N_3761,In_1193,In_2303);
nor U3762 (N_3762,In_274,In_365);
nand U3763 (N_3763,In_777,In_1327);
or U3764 (N_3764,In_1373,In_2227);
nand U3765 (N_3765,In_1236,In_1356);
and U3766 (N_3766,In_1798,In_1682);
or U3767 (N_3767,In_902,In_2231);
or U3768 (N_3768,In_2054,In_148);
nor U3769 (N_3769,In_2103,In_1697);
or U3770 (N_3770,In_300,In_1987);
nor U3771 (N_3771,In_761,In_1057);
and U3772 (N_3772,In_1607,In_1073);
or U3773 (N_3773,In_891,In_2356);
and U3774 (N_3774,In_2391,In_1098);
nor U3775 (N_3775,In_2214,In_1831);
xnor U3776 (N_3776,In_1152,In_367);
xnor U3777 (N_3777,In_1209,In_2178);
nand U3778 (N_3778,In_524,In_268);
nand U3779 (N_3779,In_2209,In_211);
and U3780 (N_3780,In_1226,In_2286);
nor U3781 (N_3781,In_2430,In_1276);
and U3782 (N_3782,In_2329,In_2433);
nor U3783 (N_3783,In_97,In_1228);
or U3784 (N_3784,In_2424,In_200);
or U3785 (N_3785,In_2342,In_2426);
nand U3786 (N_3786,In_1807,In_184);
nand U3787 (N_3787,In_363,In_1014);
and U3788 (N_3788,In_77,In_2342);
nor U3789 (N_3789,In_786,In_2174);
and U3790 (N_3790,In_1256,In_1478);
or U3791 (N_3791,In_1686,In_213);
nand U3792 (N_3792,In_588,In_1663);
or U3793 (N_3793,In_1574,In_2064);
and U3794 (N_3794,In_692,In_1265);
xor U3795 (N_3795,In_2260,In_228);
xnor U3796 (N_3796,In_1127,In_2304);
nor U3797 (N_3797,In_1262,In_576);
nand U3798 (N_3798,In_1918,In_960);
nand U3799 (N_3799,In_1208,In_2182);
nor U3800 (N_3800,In_2002,In_2162);
nand U3801 (N_3801,In_914,In_665);
nor U3802 (N_3802,In_1736,In_1134);
nor U3803 (N_3803,In_1328,In_425);
and U3804 (N_3804,In_375,In_671);
or U3805 (N_3805,In_2074,In_625);
xor U3806 (N_3806,In_117,In_1619);
or U3807 (N_3807,In_2033,In_996);
and U3808 (N_3808,In_1468,In_1618);
nand U3809 (N_3809,In_537,In_490);
nor U3810 (N_3810,In_1252,In_1370);
or U3811 (N_3811,In_2456,In_1930);
nor U3812 (N_3812,In_2069,In_1387);
and U3813 (N_3813,In_1271,In_210);
nand U3814 (N_3814,In_319,In_1012);
nand U3815 (N_3815,In_601,In_471);
and U3816 (N_3816,In_2388,In_144);
and U3817 (N_3817,In_526,In_894);
or U3818 (N_3818,In_1216,In_1878);
or U3819 (N_3819,In_2049,In_271);
or U3820 (N_3820,In_2014,In_1490);
nor U3821 (N_3821,In_1866,In_587);
nand U3822 (N_3822,In_2219,In_757);
and U3823 (N_3823,In_1145,In_2453);
nand U3824 (N_3824,In_761,In_1443);
and U3825 (N_3825,In_1020,In_1614);
nor U3826 (N_3826,In_2329,In_1922);
and U3827 (N_3827,In_17,In_81);
or U3828 (N_3828,In_12,In_1132);
or U3829 (N_3829,In_1850,In_1947);
nand U3830 (N_3830,In_569,In_1389);
nor U3831 (N_3831,In_888,In_1112);
nand U3832 (N_3832,In_1899,In_112);
and U3833 (N_3833,In_212,In_1114);
nand U3834 (N_3834,In_2177,In_128);
and U3835 (N_3835,In_1209,In_1015);
or U3836 (N_3836,In_803,In_1415);
and U3837 (N_3837,In_2415,In_1197);
or U3838 (N_3838,In_1438,In_2392);
or U3839 (N_3839,In_155,In_1730);
and U3840 (N_3840,In_2143,In_2485);
or U3841 (N_3841,In_535,In_1626);
nand U3842 (N_3842,In_2451,In_1233);
nor U3843 (N_3843,In_1561,In_995);
and U3844 (N_3844,In_401,In_210);
nor U3845 (N_3845,In_2169,In_1876);
xnor U3846 (N_3846,In_1588,In_2431);
nand U3847 (N_3847,In_1297,In_1947);
nand U3848 (N_3848,In_890,In_530);
and U3849 (N_3849,In_157,In_502);
and U3850 (N_3850,In_875,In_1814);
nor U3851 (N_3851,In_1138,In_850);
or U3852 (N_3852,In_1413,In_1235);
nand U3853 (N_3853,In_2487,In_2351);
nand U3854 (N_3854,In_1855,In_1539);
nor U3855 (N_3855,In_2240,In_1839);
nor U3856 (N_3856,In_1214,In_479);
nor U3857 (N_3857,In_949,In_1046);
or U3858 (N_3858,In_1496,In_1314);
xnor U3859 (N_3859,In_157,In_897);
and U3860 (N_3860,In_47,In_1707);
nor U3861 (N_3861,In_6,In_2233);
or U3862 (N_3862,In_532,In_778);
nor U3863 (N_3863,In_1175,In_1562);
and U3864 (N_3864,In_707,In_1147);
nor U3865 (N_3865,In_505,In_169);
or U3866 (N_3866,In_736,In_2068);
nor U3867 (N_3867,In_835,In_1507);
or U3868 (N_3868,In_281,In_1513);
or U3869 (N_3869,In_521,In_2196);
or U3870 (N_3870,In_2217,In_132);
nand U3871 (N_3871,In_1163,In_1428);
or U3872 (N_3872,In_1396,In_1043);
or U3873 (N_3873,In_872,In_1673);
and U3874 (N_3874,In_1213,In_81);
nor U3875 (N_3875,In_258,In_2385);
nor U3876 (N_3876,In_1920,In_2479);
nor U3877 (N_3877,In_828,In_799);
and U3878 (N_3878,In_468,In_2361);
and U3879 (N_3879,In_210,In_2394);
nand U3880 (N_3880,In_1513,In_2425);
or U3881 (N_3881,In_685,In_777);
nor U3882 (N_3882,In_355,In_1656);
nor U3883 (N_3883,In_1944,In_2047);
xor U3884 (N_3884,In_2458,In_276);
nor U3885 (N_3885,In_892,In_1867);
and U3886 (N_3886,In_1139,In_2286);
or U3887 (N_3887,In_502,In_2162);
nand U3888 (N_3888,In_1212,In_345);
or U3889 (N_3889,In_1066,In_1439);
nor U3890 (N_3890,In_360,In_2323);
and U3891 (N_3891,In_1250,In_1095);
and U3892 (N_3892,In_216,In_1115);
xor U3893 (N_3893,In_1897,In_1113);
nand U3894 (N_3894,In_174,In_2357);
nor U3895 (N_3895,In_1642,In_1962);
or U3896 (N_3896,In_1601,In_1342);
or U3897 (N_3897,In_1765,In_1255);
nor U3898 (N_3898,In_1985,In_2315);
and U3899 (N_3899,In_2262,In_702);
or U3900 (N_3900,In_279,In_1863);
nand U3901 (N_3901,In_2173,In_1260);
and U3902 (N_3902,In_570,In_1318);
nor U3903 (N_3903,In_1719,In_1238);
nand U3904 (N_3904,In_551,In_1472);
or U3905 (N_3905,In_2212,In_2258);
nor U3906 (N_3906,In_1373,In_234);
nor U3907 (N_3907,In_556,In_1661);
nand U3908 (N_3908,In_2382,In_807);
and U3909 (N_3909,In_1502,In_838);
or U3910 (N_3910,In_99,In_1768);
or U3911 (N_3911,In_741,In_2258);
or U3912 (N_3912,In_1096,In_144);
xor U3913 (N_3913,In_2093,In_1380);
nand U3914 (N_3914,In_311,In_1871);
or U3915 (N_3915,In_1665,In_1098);
nor U3916 (N_3916,In_1816,In_2391);
nor U3917 (N_3917,In_1047,In_1852);
nand U3918 (N_3918,In_669,In_1200);
xnor U3919 (N_3919,In_531,In_1454);
or U3920 (N_3920,In_1831,In_280);
nor U3921 (N_3921,In_300,In_1308);
or U3922 (N_3922,In_2060,In_269);
and U3923 (N_3923,In_2063,In_2260);
or U3924 (N_3924,In_193,In_823);
nand U3925 (N_3925,In_2090,In_1364);
or U3926 (N_3926,In_2378,In_1333);
and U3927 (N_3927,In_730,In_330);
nand U3928 (N_3928,In_184,In_2130);
or U3929 (N_3929,In_1818,In_1087);
or U3930 (N_3930,In_65,In_2414);
or U3931 (N_3931,In_539,In_997);
or U3932 (N_3932,In_1137,In_1100);
nor U3933 (N_3933,In_1059,In_1851);
nand U3934 (N_3934,In_1917,In_2343);
nor U3935 (N_3935,In_1614,In_268);
nand U3936 (N_3936,In_2492,In_446);
or U3937 (N_3937,In_1900,In_1893);
nor U3938 (N_3938,In_2473,In_516);
and U3939 (N_3939,In_1207,In_1140);
or U3940 (N_3940,In_257,In_777);
and U3941 (N_3941,In_2450,In_2306);
nor U3942 (N_3942,In_1292,In_1763);
nand U3943 (N_3943,In_1676,In_18);
xor U3944 (N_3944,In_1693,In_261);
and U3945 (N_3945,In_1605,In_1571);
nor U3946 (N_3946,In_2347,In_1236);
nand U3947 (N_3947,In_574,In_902);
nor U3948 (N_3948,In_1918,In_754);
nor U3949 (N_3949,In_2008,In_2389);
and U3950 (N_3950,In_1243,In_1122);
nand U3951 (N_3951,In_347,In_495);
nand U3952 (N_3952,In_1619,In_2272);
or U3953 (N_3953,In_1388,In_1958);
nand U3954 (N_3954,In_1434,In_78);
nor U3955 (N_3955,In_55,In_1073);
or U3956 (N_3956,In_377,In_1154);
nor U3957 (N_3957,In_308,In_1389);
and U3958 (N_3958,In_529,In_1528);
nor U3959 (N_3959,In_1975,In_862);
xnor U3960 (N_3960,In_597,In_415);
or U3961 (N_3961,In_487,In_1725);
and U3962 (N_3962,In_1230,In_197);
xnor U3963 (N_3963,In_1741,In_371);
and U3964 (N_3964,In_1076,In_2308);
and U3965 (N_3965,In_597,In_490);
nor U3966 (N_3966,In_1442,In_88);
and U3967 (N_3967,In_670,In_1004);
or U3968 (N_3968,In_2341,In_1104);
and U3969 (N_3969,In_183,In_2009);
xor U3970 (N_3970,In_131,In_220);
and U3971 (N_3971,In_86,In_668);
nor U3972 (N_3972,In_911,In_2151);
or U3973 (N_3973,In_1573,In_2049);
nand U3974 (N_3974,In_1496,In_1082);
nand U3975 (N_3975,In_91,In_1047);
nand U3976 (N_3976,In_122,In_2369);
nand U3977 (N_3977,In_1502,In_1171);
nand U3978 (N_3978,In_1589,In_1874);
and U3979 (N_3979,In_1054,In_1644);
and U3980 (N_3980,In_2157,In_1875);
nor U3981 (N_3981,In_1011,In_2085);
and U3982 (N_3982,In_87,In_1733);
nand U3983 (N_3983,In_2108,In_599);
or U3984 (N_3984,In_223,In_345);
and U3985 (N_3985,In_783,In_1892);
and U3986 (N_3986,In_296,In_767);
or U3987 (N_3987,In_2312,In_1793);
nand U3988 (N_3988,In_1808,In_305);
xnor U3989 (N_3989,In_790,In_843);
or U3990 (N_3990,In_899,In_1534);
nor U3991 (N_3991,In_2225,In_439);
and U3992 (N_3992,In_347,In_592);
and U3993 (N_3993,In_1185,In_2401);
or U3994 (N_3994,In_514,In_345);
or U3995 (N_3995,In_1635,In_495);
xnor U3996 (N_3996,In_1174,In_1138);
nand U3997 (N_3997,In_208,In_46);
and U3998 (N_3998,In_2079,In_2495);
and U3999 (N_3999,In_2321,In_2244);
and U4000 (N_4000,In_632,In_1030);
or U4001 (N_4001,In_705,In_1200);
and U4002 (N_4002,In_854,In_65);
xnor U4003 (N_4003,In_875,In_768);
xnor U4004 (N_4004,In_849,In_423);
xnor U4005 (N_4005,In_1735,In_1914);
or U4006 (N_4006,In_1396,In_1859);
nor U4007 (N_4007,In_216,In_963);
and U4008 (N_4008,In_981,In_332);
and U4009 (N_4009,In_238,In_739);
or U4010 (N_4010,In_1365,In_2438);
nor U4011 (N_4011,In_2115,In_2277);
nand U4012 (N_4012,In_2349,In_1855);
or U4013 (N_4013,In_2444,In_1557);
or U4014 (N_4014,In_1999,In_1542);
nand U4015 (N_4015,In_1315,In_1574);
or U4016 (N_4016,In_636,In_357);
nor U4017 (N_4017,In_586,In_961);
xnor U4018 (N_4018,In_82,In_2096);
nor U4019 (N_4019,In_1013,In_1980);
xor U4020 (N_4020,In_2400,In_1299);
nor U4021 (N_4021,In_1324,In_1597);
and U4022 (N_4022,In_714,In_1824);
xnor U4023 (N_4023,In_1132,In_1711);
or U4024 (N_4024,In_1781,In_153);
nor U4025 (N_4025,In_1310,In_2033);
or U4026 (N_4026,In_69,In_837);
and U4027 (N_4027,In_305,In_1086);
nand U4028 (N_4028,In_1967,In_808);
nand U4029 (N_4029,In_784,In_1808);
or U4030 (N_4030,In_2013,In_317);
nor U4031 (N_4031,In_2249,In_1869);
or U4032 (N_4032,In_901,In_145);
nor U4033 (N_4033,In_2438,In_924);
and U4034 (N_4034,In_993,In_940);
or U4035 (N_4035,In_2429,In_1082);
and U4036 (N_4036,In_2085,In_453);
nand U4037 (N_4037,In_1393,In_486);
and U4038 (N_4038,In_2424,In_2186);
and U4039 (N_4039,In_2140,In_847);
nor U4040 (N_4040,In_1839,In_310);
or U4041 (N_4041,In_2303,In_1050);
or U4042 (N_4042,In_2154,In_1121);
nor U4043 (N_4043,In_488,In_655);
nor U4044 (N_4044,In_200,In_204);
xnor U4045 (N_4045,In_1554,In_1634);
and U4046 (N_4046,In_1620,In_1365);
or U4047 (N_4047,In_1322,In_2364);
and U4048 (N_4048,In_359,In_1909);
and U4049 (N_4049,In_2455,In_1250);
and U4050 (N_4050,In_2387,In_1100);
or U4051 (N_4051,In_869,In_1737);
nor U4052 (N_4052,In_2452,In_1742);
and U4053 (N_4053,In_2104,In_329);
nand U4054 (N_4054,In_911,In_1108);
xor U4055 (N_4055,In_1182,In_2148);
or U4056 (N_4056,In_948,In_2267);
nor U4057 (N_4057,In_1735,In_2470);
and U4058 (N_4058,In_2202,In_1056);
or U4059 (N_4059,In_1263,In_1264);
nand U4060 (N_4060,In_70,In_2478);
or U4061 (N_4061,In_2194,In_1071);
and U4062 (N_4062,In_371,In_306);
nor U4063 (N_4063,In_2085,In_1082);
xnor U4064 (N_4064,In_425,In_1586);
xnor U4065 (N_4065,In_2190,In_691);
and U4066 (N_4066,In_1169,In_1625);
nand U4067 (N_4067,In_1479,In_1348);
xor U4068 (N_4068,In_565,In_1489);
or U4069 (N_4069,In_99,In_1266);
xnor U4070 (N_4070,In_1618,In_752);
nor U4071 (N_4071,In_469,In_2100);
xor U4072 (N_4072,In_656,In_176);
nand U4073 (N_4073,In_858,In_1626);
nand U4074 (N_4074,In_2095,In_127);
nor U4075 (N_4075,In_1368,In_1571);
nand U4076 (N_4076,In_2166,In_1975);
nand U4077 (N_4077,In_2119,In_1580);
and U4078 (N_4078,In_1595,In_741);
xnor U4079 (N_4079,In_1955,In_847);
and U4080 (N_4080,In_533,In_2427);
or U4081 (N_4081,In_250,In_1189);
and U4082 (N_4082,In_59,In_1454);
nor U4083 (N_4083,In_1533,In_1382);
and U4084 (N_4084,In_29,In_1242);
or U4085 (N_4085,In_1971,In_585);
xnor U4086 (N_4086,In_945,In_881);
nor U4087 (N_4087,In_1539,In_1909);
nor U4088 (N_4088,In_30,In_1245);
and U4089 (N_4089,In_2352,In_1675);
nand U4090 (N_4090,In_2277,In_408);
nor U4091 (N_4091,In_2155,In_117);
xor U4092 (N_4092,In_1295,In_1015);
or U4093 (N_4093,In_1091,In_453);
and U4094 (N_4094,In_197,In_1279);
nand U4095 (N_4095,In_1889,In_161);
nand U4096 (N_4096,In_484,In_621);
xnor U4097 (N_4097,In_2463,In_1639);
nand U4098 (N_4098,In_1910,In_146);
and U4099 (N_4099,In_2460,In_1995);
nand U4100 (N_4100,In_71,In_1092);
or U4101 (N_4101,In_1460,In_635);
nand U4102 (N_4102,In_2273,In_520);
nand U4103 (N_4103,In_1130,In_956);
and U4104 (N_4104,In_537,In_660);
xor U4105 (N_4105,In_804,In_1814);
and U4106 (N_4106,In_472,In_1588);
nand U4107 (N_4107,In_698,In_277);
nand U4108 (N_4108,In_779,In_1032);
and U4109 (N_4109,In_2347,In_1107);
and U4110 (N_4110,In_1429,In_328);
nand U4111 (N_4111,In_2454,In_256);
nor U4112 (N_4112,In_316,In_247);
nor U4113 (N_4113,In_1586,In_548);
nor U4114 (N_4114,In_732,In_1932);
nand U4115 (N_4115,In_1066,In_2194);
nor U4116 (N_4116,In_2216,In_1849);
xor U4117 (N_4117,In_409,In_864);
nor U4118 (N_4118,In_242,In_2316);
nor U4119 (N_4119,In_1215,In_1381);
nand U4120 (N_4120,In_917,In_2056);
nand U4121 (N_4121,In_2078,In_127);
and U4122 (N_4122,In_572,In_2256);
nand U4123 (N_4123,In_143,In_1846);
nand U4124 (N_4124,In_1055,In_371);
or U4125 (N_4125,In_2284,In_1753);
xor U4126 (N_4126,In_2058,In_840);
xnor U4127 (N_4127,In_1848,In_1112);
or U4128 (N_4128,In_2452,In_1142);
or U4129 (N_4129,In_1811,In_463);
nand U4130 (N_4130,In_2202,In_36);
nor U4131 (N_4131,In_707,In_1330);
and U4132 (N_4132,In_1095,In_723);
or U4133 (N_4133,In_559,In_1176);
and U4134 (N_4134,In_2023,In_337);
nand U4135 (N_4135,In_1186,In_910);
and U4136 (N_4136,In_449,In_1365);
and U4137 (N_4137,In_102,In_324);
and U4138 (N_4138,In_1557,In_442);
nor U4139 (N_4139,In_2113,In_1291);
and U4140 (N_4140,In_753,In_1356);
or U4141 (N_4141,In_666,In_670);
and U4142 (N_4142,In_394,In_2103);
and U4143 (N_4143,In_2094,In_2277);
nor U4144 (N_4144,In_412,In_1723);
or U4145 (N_4145,In_770,In_2029);
or U4146 (N_4146,In_2244,In_56);
xnor U4147 (N_4147,In_1141,In_2216);
or U4148 (N_4148,In_1158,In_307);
xnor U4149 (N_4149,In_701,In_1890);
or U4150 (N_4150,In_1790,In_651);
and U4151 (N_4151,In_837,In_1677);
and U4152 (N_4152,In_2187,In_1576);
nand U4153 (N_4153,In_2161,In_388);
and U4154 (N_4154,In_2451,In_75);
nand U4155 (N_4155,In_2497,In_2245);
nand U4156 (N_4156,In_2380,In_664);
and U4157 (N_4157,In_1202,In_2249);
or U4158 (N_4158,In_2240,In_1523);
nand U4159 (N_4159,In_1439,In_1179);
nand U4160 (N_4160,In_1528,In_85);
and U4161 (N_4161,In_2446,In_1956);
and U4162 (N_4162,In_2046,In_1426);
and U4163 (N_4163,In_972,In_36);
and U4164 (N_4164,In_1204,In_2226);
or U4165 (N_4165,In_1826,In_2299);
nor U4166 (N_4166,In_1919,In_1717);
xor U4167 (N_4167,In_1318,In_1194);
nand U4168 (N_4168,In_437,In_1297);
nor U4169 (N_4169,In_730,In_1586);
xor U4170 (N_4170,In_107,In_1787);
or U4171 (N_4171,In_1819,In_2310);
or U4172 (N_4172,In_2376,In_148);
xor U4173 (N_4173,In_1589,In_325);
and U4174 (N_4174,In_1629,In_1581);
nand U4175 (N_4175,In_285,In_474);
or U4176 (N_4176,In_1097,In_225);
and U4177 (N_4177,In_992,In_1542);
or U4178 (N_4178,In_1484,In_68);
or U4179 (N_4179,In_39,In_2070);
and U4180 (N_4180,In_275,In_936);
nor U4181 (N_4181,In_589,In_1629);
nand U4182 (N_4182,In_2305,In_2086);
nor U4183 (N_4183,In_2244,In_54);
or U4184 (N_4184,In_793,In_301);
or U4185 (N_4185,In_1710,In_1497);
and U4186 (N_4186,In_954,In_560);
nand U4187 (N_4187,In_289,In_1824);
or U4188 (N_4188,In_1724,In_1960);
nor U4189 (N_4189,In_778,In_1883);
and U4190 (N_4190,In_1145,In_1551);
and U4191 (N_4191,In_486,In_2011);
or U4192 (N_4192,In_2216,In_130);
nand U4193 (N_4193,In_1795,In_994);
nand U4194 (N_4194,In_1228,In_1592);
or U4195 (N_4195,In_1977,In_1082);
or U4196 (N_4196,In_1800,In_1568);
xor U4197 (N_4197,In_1710,In_137);
and U4198 (N_4198,In_1017,In_1307);
and U4199 (N_4199,In_1109,In_605);
nor U4200 (N_4200,In_380,In_1521);
or U4201 (N_4201,In_1101,In_886);
nand U4202 (N_4202,In_1698,In_1960);
nor U4203 (N_4203,In_257,In_517);
and U4204 (N_4204,In_237,In_1383);
and U4205 (N_4205,In_2063,In_634);
xnor U4206 (N_4206,In_1129,In_2052);
nand U4207 (N_4207,In_879,In_2432);
and U4208 (N_4208,In_1163,In_963);
nor U4209 (N_4209,In_2400,In_1371);
and U4210 (N_4210,In_2058,In_1141);
and U4211 (N_4211,In_1812,In_1424);
and U4212 (N_4212,In_1433,In_1049);
and U4213 (N_4213,In_2102,In_909);
nor U4214 (N_4214,In_1180,In_1260);
xnor U4215 (N_4215,In_62,In_881);
or U4216 (N_4216,In_335,In_2388);
or U4217 (N_4217,In_1338,In_2347);
nand U4218 (N_4218,In_243,In_2404);
nand U4219 (N_4219,In_82,In_2115);
xor U4220 (N_4220,In_642,In_363);
nor U4221 (N_4221,In_391,In_2347);
nand U4222 (N_4222,In_1996,In_1753);
and U4223 (N_4223,In_809,In_2248);
nor U4224 (N_4224,In_1226,In_1332);
and U4225 (N_4225,In_650,In_1967);
nor U4226 (N_4226,In_877,In_2073);
and U4227 (N_4227,In_651,In_381);
and U4228 (N_4228,In_1931,In_1632);
and U4229 (N_4229,In_1847,In_2253);
nor U4230 (N_4230,In_1899,In_1241);
nor U4231 (N_4231,In_2493,In_1316);
nand U4232 (N_4232,In_1390,In_2000);
nor U4233 (N_4233,In_120,In_1172);
nor U4234 (N_4234,In_489,In_2431);
or U4235 (N_4235,In_650,In_455);
and U4236 (N_4236,In_130,In_2395);
or U4237 (N_4237,In_302,In_1496);
nand U4238 (N_4238,In_1068,In_1827);
nand U4239 (N_4239,In_1951,In_1332);
nand U4240 (N_4240,In_1403,In_618);
or U4241 (N_4241,In_1828,In_858);
or U4242 (N_4242,In_409,In_522);
nor U4243 (N_4243,In_1628,In_1507);
and U4244 (N_4244,In_2069,In_1293);
nor U4245 (N_4245,In_2036,In_9);
or U4246 (N_4246,In_2442,In_516);
xor U4247 (N_4247,In_1833,In_308);
nor U4248 (N_4248,In_6,In_1477);
or U4249 (N_4249,In_2127,In_2029);
and U4250 (N_4250,In_815,In_1832);
and U4251 (N_4251,In_557,In_325);
nand U4252 (N_4252,In_634,In_745);
nand U4253 (N_4253,In_448,In_981);
and U4254 (N_4254,In_1427,In_146);
nor U4255 (N_4255,In_1568,In_389);
nand U4256 (N_4256,In_480,In_2);
or U4257 (N_4257,In_1253,In_1796);
nand U4258 (N_4258,In_704,In_1686);
nor U4259 (N_4259,In_2154,In_2279);
nor U4260 (N_4260,In_743,In_148);
xor U4261 (N_4261,In_2468,In_2219);
nand U4262 (N_4262,In_230,In_2480);
nand U4263 (N_4263,In_706,In_217);
nor U4264 (N_4264,In_2318,In_15);
and U4265 (N_4265,In_924,In_282);
nor U4266 (N_4266,In_589,In_677);
nand U4267 (N_4267,In_1119,In_2344);
or U4268 (N_4268,In_617,In_1364);
and U4269 (N_4269,In_726,In_901);
and U4270 (N_4270,In_25,In_2456);
or U4271 (N_4271,In_462,In_7);
nand U4272 (N_4272,In_1757,In_2439);
xor U4273 (N_4273,In_750,In_2116);
nand U4274 (N_4274,In_2123,In_2307);
xor U4275 (N_4275,In_2497,In_1593);
nand U4276 (N_4276,In_1998,In_319);
nor U4277 (N_4277,In_1798,In_1663);
nand U4278 (N_4278,In_1142,In_1348);
and U4279 (N_4279,In_830,In_649);
xnor U4280 (N_4280,In_2183,In_1124);
xnor U4281 (N_4281,In_1552,In_236);
or U4282 (N_4282,In_676,In_1139);
nor U4283 (N_4283,In_502,In_15);
nand U4284 (N_4284,In_426,In_1799);
nor U4285 (N_4285,In_2087,In_1798);
and U4286 (N_4286,In_1726,In_1641);
or U4287 (N_4287,In_1428,In_1513);
or U4288 (N_4288,In_284,In_2297);
nand U4289 (N_4289,In_1108,In_643);
and U4290 (N_4290,In_160,In_956);
nand U4291 (N_4291,In_2240,In_263);
nor U4292 (N_4292,In_1062,In_1224);
or U4293 (N_4293,In_1210,In_1548);
nor U4294 (N_4294,In_2201,In_1104);
or U4295 (N_4295,In_1358,In_2433);
and U4296 (N_4296,In_464,In_1013);
nor U4297 (N_4297,In_2076,In_1919);
or U4298 (N_4298,In_2101,In_85);
nor U4299 (N_4299,In_105,In_2261);
and U4300 (N_4300,In_1252,In_1729);
or U4301 (N_4301,In_1770,In_1280);
nor U4302 (N_4302,In_792,In_581);
or U4303 (N_4303,In_1886,In_1482);
nand U4304 (N_4304,In_965,In_864);
nand U4305 (N_4305,In_1363,In_2197);
nand U4306 (N_4306,In_2027,In_2319);
nor U4307 (N_4307,In_70,In_1477);
nor U4308 (N_4308,In_270,In_1063);
and U4309 (N_4309,In_734,In_2360);
nor U4310 (N_4310,In_1694,In_2212);
or U4311 (N_4311,In_1757,In_393);
or U4312 (N_4312,In_1182,In_2224);
and U4313 (N_4313,In_2321,In_114);
or U4314 (N_4314,In_153,In_1922);
nor U4315 (N_4315,In_312,In_2017);
or U4316 (N_4316,In_1633,In_1233);
nand U4317 (N_4317,In_340,In_717);
nor U4318 (N_4318,In_2366,In_2259);
nand U4319 (N_4319,In_2166,In_2446);
xor U4320 (N_4320,In_1956,In_6);
xor U4321 (N_4321,In_2262,In_747);
nor U4322 (N_4322,In_1625,In_1050);
or U4323 (N_4323,In_2127,In_1802);
and U4324 (N_4324,In_1439,In_1414);
or U4325 (N_4325,In_464,In_1719);
nor U4326 (N_4326,In_1456,In_193);
xor U4327 (N_4327,In_2052,In_925);
nor U4328 (N_4328,In_2314,In_2093);
or U4329 (N_4329,In_1356,In_939);
and U4330 (N_4330,In_545,In_2213);
nand U4331 (N_4331,In_1155,In_975);
nand U4332 (N_4332,In_544,In_1985);
and U4333 (N_4333,In_1857,In_1406);
nor U4334 (N_4334,In_1954,In_2244);
nor U4335 (N_4335,In_1449,In_2099);
and U4336 (N_4336,In_1008,In_1874);
nor U4337 (N_4337,In_801,In_1063);
xnor U4338 (N_4338,In_2017,In_860);
or U4339 (N_4339,In_25,In_220);
or U4340 (N_4340,In_381,In_2325);
or U4341 (N_4341,In_2432,In_1534);
nand U4342 (N_4342,In_391,In_779);
or U4343 (N_4343,In_2354,In_640);
nand U4344 (N_4344,In_2138,In_1815);
nor U4345 (N_4345,In_799,In_497);
nor U4346 (N_4346,In_2456,In_1673);
or U4347 (N_4347,In_712,In_2325);
xnor U4348 (N_4348,In_266,In_2062);
nor U4349 (N_4349,In_1892,In_1915);
or U4350 (N_4350,In_1466,In_1139);
xnor U4351 (N_4351,In_1911,In_809);
nor U4352 (N_4352,In_1802,In_2492);
or U4353 (N_4353,In_1505,In_1311);
or U4354 (N_4354,In_1491,In_2115);
xor U4355 (N_4355,In_2044,In_2088);
xnor U4356 (N_4356,In_1449,In_991);
and U4357 (N_4357,In_474,In_1982);
or U4358 (N_4358,In_611,In_1475);
and U4359 (N_4359,In_287,In_864);
nand U4360 (N_4360,In_1301,In_1705);
or U4361 (N_4361,In_1557,In_492);
nand U4362 (N_4362,In_2098,In_1802);
or U4363 (N_4363,In_1525,In_1775);
or U4364 (N_4364,In_1757,In_1364);
nand U4365 (N_4365,In_326,In_491);
nand U4366 (N_4366,In_2369,In_1814);
or U4367 (N_4367,In_1275,In_1692);
or U4368 (N_4368,In_252,In_2315);
nor U4369 (N_4369,In_1663,In_982);
nand U4370 (N_4370,In_1778,In_462);
or U4371 (N_4371,In_635,In_1130);
or U4372 (N_4372,In_1635,In_116);
and U4373 (N_4373,In_1194,In_2201);
or U4374 (N_4374,In_182,In_2317);
nor U4375 (N_4375,In_2212,In_485);
nand U4376 (N_4376,In_1195,In_1032);
or U4377 (N_4377,In_2079,In_961);
or U4378 (N_4378,In_1746,In_136);
and U4379 (N_4379,In_2105,In_159);
and U4380 (N_4380,In_1916,In_2259);
or U4381 (N_4381,In_386,In_2200);
and U4382 (N_4382,In_1995,In_579);
and U4383 (N_4383,In_2438,In_721);
or U4384 (N_4384,In_164,In_1918);
nand U4385 (N_4385,In_917,In_1693);
and U4386 (N_4386,In_123,In_1453);
nand U4387 (N_4387,In_2142,In_1459);
nor U4388 (N_4388,In_782,In_1101);
and U4389 (N_4389,In_2083,In_354);
nor U4390 (N_4390,In_2286,In_949);
nor U4391 (N_4391,In_2239,In_1670);
and U4392 (N_4392,In_1606,In_128);
and U4393 (N_4393,In_2453,In_2147);
nand U4394 (N_4394,In_2169,In_21);
nand U4395 (N_4395,In_2295,In_471);
and U4396 (N_4396,In_1027,In_1580);
or U4397 (N_4397,In_495,In_1090);
and U4398 (N_4398,In_510,In_1245);
nand U4399 (N_4399,In_2084,In_1885);
and U4400 (N_4400,In_443,In_299);
nand U4401 (N_4401,In_1076,In_1409);
or U4402 (N_4402,In_212,In_1285);
and U4403 (N_4403,In_2121,In_2223);
nor U4404 (N_4404,In_1113,In_372);
or U4405 (N_4405,In_693,In_81);
and U4406 (N_4406,In_2355,In_1668);
or U4407 (N_4407,In_623,In_1460);
nand U4408 (N_4408,In_444,In_329);
nor U4409 (N_4409,In_1242,In_2131);
or U4410 (N_4410,In_1854,In_2125);
nor U4411 (N_4411,In_614,In_793);
or U4412 (N_4412,In_893,In_721);
xor U4413 (N_4413,In_2358,In_1440);
and U4414 (N_4414,In_1377,In_1086);
and U4415 (N_4415,In_1567,In_1875);
or U4416 (N_4416,In_1950,In_1323);
nor U4417 (N_4417,In_377,In_91);
xnor U4418 (N_4418,In_1261,In_2396);
nand U4419 (N_4419,In_1935,In_881);
or U4420 (N_4420,In_2317,In_782);
xnor U4421 (N_4421,In_1262,In_365);
nand U4422 (N_4422,In_1221,In_1085);
or U4423 (N_4423,In_1727,In_289);
nand U4424 (N_4424,In_1523,In_1725);
nor U4425 (N_4425,In_46,In_1950);
xnor U4426 (N_4426,In_989,In_1072);
xnor U4427 (N_4427,In_479,In_2126);
or U4428 (N_4428,In_1384,In_1171);
or U4429 (N_4429,In_2343,In_2308);
or U4430 (N_4430,In_1378,In_1419);
or U4431 (N_4431,In_2391,In_1800);
nor U4432 (N_4432,In_1538,In_2470);
nor U4433 (N_4433,In_1903,In_1579);
and U4434 (N_4434,In_266,In_983);
nor U4435 (N_4435,In_1391,In_1733);
and U4436 (N_4436,In_1358,In_1974);
xor U4437 (N_4437,In_634,In_350);
nor U4438 (N_4438,In_1787,In_1137);
nor U4439 (N_4439,In_1521,In_1660);
nand U4440 (N_4440,In_2405,In_103);
nor U4441 (N_4441,In_195,In_723);
nand U4442 (N_4442,In_445,In_1215);
xor U4443 (N_4443,In_1967,In_1800);
nor U4444 (N_4444,In_1943,In_1748);
or U4445 (N_4445,In_1004,In_579);
or U4446 (N_4446,In_2027,In_2349);
xnor U4447 (N_4447,In_917,In_2329);
and U4448 (N_4448,In_641,In_253);
xor U4449 (N_4449,In_1886,In_2406);
nand U4450 (N_4450,In_881,In_814);
or U4451 (N_4451,In_245,In_482);
nor U4452 (N_4452,In_982,In_398);
nand U4453 (N_4453,In_591,In_1415);
or U4454 (N_4454,In_825,In_297);
nor U4455 (N_4455,In_1858,In_691);
nor U4456 (N_4456,In_1387,In_922);
or U4457 (N_4457,In_767,In_2000);
or U4458 (N_4458,In_208,In_970);
nor U4459 (N_4459,In_446,In_2382);
and U4460 (N_4460,In_676,In_1489);
and U4461 (N_4461,In_1017,In_1584);
nand U4462 (N_4462,In_2246,In_1853);
nand U4463 (N_4463,In_364,In_1603);
or U4464 (N_4464,In_2038,In_1331);
nor U4465 (N_4465,In_441,In_700);
nand U4466 (N_4466,In_477,In_1792);
and U4467 (N_4467,In_2494,In_1650);
nand U4468 (N_4468,In_116,In_2467);
nor U4469 (N_4469,In_1988,In_717);
nor U4470 (N_4470,In_2112,In_1849);
and U4471 (N_4471,In_2459,In_1140);
or U4472 (N_4472,In_1179,In_691);
nand U4473 (N_4473,In_402,In_448);
nor U4474 (N_4474,In_944,In_1469);
xor U4475 (N_4475,In_1133,In_1080);
or U4476 (N_4476,In_1290,In_1453);
or U4477 (N_4477,In_483,In_1070);
nand U4478 (N_4478,In_1843,In_1655);
or U4479 (N_4479,In_34,In_1581);
nor U4480 (N_4480,In_1927,In_2004);
nand U4481 (N_4481,In_1948,In_1926);
and U4482 (N_4482,In_1340,In_572);
and U4483 (N_4483,In_2414,In_2007);
and U4484 (N_4484,In_1062,In_633);
and U4485 (N_4485,In_1374,In_2347);
nand U4486 (N_4486,In_2304,In_860);
nand U4487 (N_4487,In_1298,In_2317);
or U4488 (N_4488,In_1835,In_2137);
or U4489 (N_4489,In_1407,In_615);
and U4490 (N_4490,In_1517,In_156);
or U4491 (N_4491,In_488,In_1481);
nor U4492 (N_4492,In_957,In_1357);
or U4493 (N_4493,In_1102,In_1668);
and U4494 (N_4494,In_219,In_1500);
xor U4495 (N_4495,In_1542,In_711);
or U4496 (N_4496,In_1760,In_598);
xnor U4497 (N_4497,In_2300,In_2489);
or U4498 (N_4498,In_1699,In_599);
xnor U4499 (N_4499,In_2270,In_96);
and U4500 (N_4500,In_1660,In_906);
nand U4501 (N_4501,In_1320,In_2099);
nor U4502 (N_4502,In_2064,In_1591);
nor U4503 (N_4503,In_1584,In_1072);
nand U4504 (N_4504,In_145,In_501);
nand U4505 (N_4505,In_654,In_2407);
nor U4506 (N_4506,In_1397,In_2024);
nor U4507 (N_4507,In_1752,In_392);
nand U4508 (N_4508,In_288,In_2141);
nor U4509 (N_4509,In_874,In_588);
nor U4510 (N_4510,In_1866,In_1923);
xnor U4511 (N_4511,In_2299,In_16);
or U4512 (N_4512,In_763,In_2240);
and U4513 (N_4513,In_14,In_1424);
and U4514 (N_4514,In_754,In_2079);
nor U4515 (N_4515,In_1009,In_350);
xor U4516 (N_4516,In_421,In_1871);
nand U4517 (N_4517,In_233,In_2365);
or U4518 (N_4518,In_269,In_60);
xnor U4519 (N_4519,In_624,In_841);
or U4520 (N_4520,In_2231,In_2345);
and U4521 (N_4521,In_432,In_1404);
nor U4522 (N_4522,In_1141,In_1919);
xnor U4523 (N_4523,In_1373,In_133);
and U4524 (N_4524,In_2162,In_1693);
or U4525 (N_4525,In_1831,In_752);
nor U4526 (N_4526,In_396,In_2087);
and U4527 (N_4527,In_1714,In_2429);
nor U4528 (N_4528,In_42,In_1096);
and U4529 (N_4529,In_765,In_1157);
and U4530 (N_4530,In_1253,In_2403);
and U4531 (N_4531,In_1415,In_2246);
and U4532 (N_4532,In_1899,In_2484);
nand U4533 (N_4533,In_391,In_257);
nor U4534 (N_4534,In_2064,In_594);
and U4535 (N_4535,In_2251,In_2071);
xor U4536 (N_4536,In_1009,In_2497);
or U4537 (N_4537,In_2005,In_694);
and U4538 (N_4538,In_347,In_1424);
xnor U4539 (N_4539,In_4,In_1155);
or U4540 (N_4540,In_2102,In_777);
xor U4541 (N_4541,In_831,In_1288);
xor U4542 (N_4542,In_2251,In_1159);
or U4543 (N_4543,In_1187,In_1837);
nor U4544 (N_4544,In_1331,In_215);
and U4545 (N_4545,In_127,In_175);
nand U4546 (N_4546,In_177,In_968);
and U4547 (N_4547,In_1956,In_1061);
or U4548 (N_4548,In_1323,In_269);
nand U4549 (N_4549,In_282,In_2005);
or U4550 (N_4550,In_314,In_2018);
and U4551 (N_4551,In_1020,In_2189);
and U4552 (N_4552,In_519,In_59);
nand U4553 (N_4553,In_127,In_563);
and U4554 (N_4554,In_1424,In_349);
nor U4555 (N_4555,In_353,In_1881);
nor U4556 (N_4556,In_1962,In_1762);
or U4557 (N_4557,In_1987,In_1796);
nand U4558 (N_4558,In_2478,In_2234);
nor U4559 (N_4559,In_1603,In_1721);
nand U4560 (N_4560,In_2374,In_2491);
or U4561 (N_4561,In_145,In_768);
or U4562 (N_4562,In_1718,In_836);
nand U4563 (N_4563,In_1333,In_1307);
and U4564 (N_4564,In_956,In_421);
or U4565 (N_4565,In_479,In_2493);
or U4566 (N_4566,In_314,In_63);
and U4567 (N_4567,In_1665,In_2115);
nor U4568 (N_4568,In_2016,In_1570);
nand U4569 (N_4569,In_1414,In_2185);
or U4570 (N_4570,In_495,In_1179);
and U4571 (N_4571,In_1622,In_755);
and U4572 (N_4572,In_1113,In_2176);
or U4573 (N_4573,In_2264,In_2007);
or U4574 (N_4574,In_1014,In_2274);
or U4575 (N_4575,In_1336,In_956);
or U4576 (N_4576,In_1892,In_931);
or U4577 (N_4577,In_1615,In_530);
xor U4578 (N_4578,In_313,In_649);
nor U4579 (N_4579,In_1511,In_1238);
xor U4580 (N_4580,In_1956,In_615);
xnor U4581 (N_4581,In_1457,In_889);
or U4582 (N_4582,In_2274,In_1992);
nand U4583 (N_4583,In_1613,In_192);
nor U4584 (N_4584,In_1539,In_1746);
xnor U4585 (N_4585,In_1204,In_648);
and U4586 (N_4586,In_841,In_2069);
nor U4587 (N_4587,In_1639,In_1953);
or U4588 (N_4588,In_247,In_227);
nand U4589 (N_4589,In_1923,In_688);
and U4590 (N_4590,In_2346,In_549);
and U4591 (N_4591,In_955,In_2489);
nor U4592 (N_4592,In_1992,In_290);
and U4593 (N_4593,In_1267,In_1198);
and U4594 (N_4594,In_911,In_1803);
or U4595 (N_4595,In_1852,In_1843);
nor U4596 (N_4596,In_1843,In_1143);
nor U4597 (N_4597,In_1006,In_1061);
nand U4598 (N_4598,In_806,In_765);
nor U4599 (N_4599,In_2114,In_253);
or U4600 (N_4600,In_1823,In_1072);
xnor U4601 (N_4601,In_1699,In_1639);
or U4602 (N_4602,In_381,In_1031);
or U4603 (N_4603,In_191,In_908);
or U4604 (N_4604,In_285,In_1114);
nor U4605 (N_4605,In_1019,In_1411);
or U4606 (N_4606,In_1671,In_1135);
nor U4607 (N_4607,In_175,In_2171);
or U4608 (N_4608,In_294,In_655);
nand U4609 (N_4609,In_855,In_1089);
nor U4610 (N_4610,In_481,In_20);
nand U4611 (N_4611,In_1187,In_205);
nor U4612 (N_4612,In_2251,In_1059);
nand U4613 (N_4613,In_470,In_1587);
and U4614 (N_4614,In_2250,In_98);
and U4615 (N_4615,In_855,In_2118);
nand U4616 (N_4616,In_2027,In_2217);
or U4617 (N_4617,In_1032,In_2417);
nand U4618 (N_4618,In_511,In_1071);
xnor U4619 (N_4619,In_1329,In_1759);
or U4620 (N_4620,In_1666,In_1914);
or U4621 (N_4621,In_2139,In_2010);
nor U4622 (N_4622,In_371,In_2109);
nand U4623 (N_4623,In_920,In_1156);
nor U4624 (N_4624,In_1318,In_554);
nand U4625 (N_4625,In_1875,In_980);
or U4626 (N_4626,In_1989,In_66);
nor U4627 (N_4627,In_842,In_2151);
nor U4628 (N_4628,In_1669,In_2396);
or U4629 (N_4629,In_443,In_781);
nand U4630 (N_4630,In_2327,In_677);
nand U4631 (N_4631,In_439,In_619);
nor U4632 (N_4632,In_1651,In_610);
or U4633 (N_4633,In_1634,In_189);
nor U4634 (N_4634,In_2286,In_2356);
nand U4635 (N_4635,In_486,In_2459);
nand U4636 (N_4636,In_2257,In_977);
nand U4637 (N_4637,In_1093,In_28);
and U4638 (N_4638,In_1896,In_1484);
nand U4639 (N_4639,In_598,In_289);
nand U4640 (N_4640,In_1378,In_1274);
or U4641 (N_4641,In_646,In_1108);
and U4642 (N_4642,In_1058,In_1536);
nor U4643 (N_4643,In_1023,In_2082);
nand U4644 (N_4644,In_73,In_801);
and U4645 (N_4645,In_1525,In_1149);
nand U4646 (N_4646,In_2154,In_1223);
nand U4647 (N_4647,In_450,In_1062);
nor U4648 (N_4648,In_248,In_1645);
or U4649 (N_4649,In_1743,In_1067);
or U4650 (N_4650,In_2006,In_2176);
nand U4651 (N_4651,In_205,In_82);
or U4652 (N_4652,In_1090,In_898);
nor U4653 (N_4653,In_2375,In_1206);
nor U4654 (N_4654,In_1465,In_663);
nand U4655 (N_4655,In_2388,In_1758);
or U4656 (N_4656,In_925,In_2145);
nand U4657 (N_4657,In_1589,In_201);
and U4658 (N_4658,In_2450,In_1985);
and U4659 (N_4659,In_598,In_609);
and U4660 (N_4660,In_1711,In_1620);
and U4661 (N_4661,In_1354,In_584);
nand U4662 (N_4662,In_1873,In_647);
and U4663 (N_4663,In_2169,In_688);
xnor U4664 (N_4664,In_52,In_2245);
or U4665 (N_4665,In_751,In_195);
nor U4666 (N_4666,In_1637,In_2285);
nor U4667 (N_4667,In_1703,In_1221);
nor U4668 (N_4668,In_1972,In_744);
or U4669 (N_4669,In_1148,In_491);
nand U4670 (N_4670,In_2110,In_546);
nand U4671 (N_4671,In_2216,In_1535);
and U4672 (N_4672,In_1173,In_509);
or U4673 (N_4673,In_1322,In_1889);
and U4674 (N_4674,In_1928,In_629);
and U4675 (N_4675,In_2321,In_1128);
or U4676 (N_4676,In_1307,In_2096);
and U4677 (N_4677,In_1896,In_1007);
and U4678 (N_4678,In_317,In_1478);
nand U4679 (N_4679,In_2238,In_1153);
nor U4680 (N_4680,In_771,In_2131);
nand U4681 (N_4681,In_429,In_1142);
and U4682 (N_4682,In_2476,In_1157);
or U4683 (N_4683,In_1779,In_274);
nor U4684 (N_4684,In_697,In_45);
nor U4685 (N_4685,In_2152,In_1781);
or U4686 (N_4686,In_1011,In_2279);
nor U4687 (N_4687,In_1500,In_1487);
or U4688 (N_4688,In_728,In_103);
and U4689 (N_4689,In_1239,In_2008);
nor U4690 (N_4690,In_1261,In_1334);
xor U4691 (N_4691,In_2412,In_256);
nor U4692 (N_4692,In_1642,In_1300);
nor U4693 (N_4693,In_471,In_171);
or U4694 (N_4694,In_2027,In_2102);
nor U4695 (N_4695,In_807,In_2118);
xor U4696 (N_4696,In_193,In_561);
or U4697 (N_4697,In_444,In_1092);
or U4698 (N_4698,In_1392,In_748);
nor U4699 (N_4699,In_1779,In_1135);
nand U4700 (N_4700,In_1745,In_1467);
nor U4701 (N_4701,In_2062,In_408);
and U4702 (N_4702,In_2093,In_514);
xnor U4703 (N_4703,In_2403,In_1174);
or U4704 (N_4704,In_810,In_1811);
nand U4705 (N_4705,In_2395,In_1478);
nor U4706 (N_4706,In_406,In_1489);
xor U4707 (N_4707,In_1223,In_1710);
nor U4708 (N_4708,In_444,In_420);
and U4709 (N_4709,In_1113,In_1178);
nor U4710 (N_4710,In_490,In_227);
nor U4711 (N_4711,In_1067,In_652);
nand U4712 (N_4712,In_2060,In_2198);
or U4713 (N_4713,In_1370,In_1376);
and U4714 (N_4714,In_1960,In_515);
nor U4715 (N_4715,In_229,In_2411);
nor U4716 (N_4716,In_1719,In_409);
or U4717 (N_4717,In_1892,In_2038);
nor U4718 (N_4718,In_1520,In_1070);
or U4719 (N_4719,In_1184,In_2190);
and U4720 (N_4720,In_790,In_1921);
nand U4721 (N_4721,In_1113,In_469);
nand U4722 (N_4722,In_608,In_544);
and U4723 (N_4723,In_1560,In_590);
or U4724 (N_4724,In_964,In_517);
or U4725 (N_4725,In_545,In_1555);
or U4726 (N_4726,In_2379,In_1901);
nor U4727 (N_4727,In_2162,In_644);
or U4728 (N_4728,In_85,In_1215);
nor U4729 (N_4729,In_136,In_1021);
nor U4730 (N_4730,In_1530,In_778);
xor U4731 (N_4731,In_757,In_3);
nor U4732 (N_4732,In_1979,In_1154);
and U4733 (N_4733,In_2169,In_1891);
nand U4734 (N_4734,In_1217,In_1494);
nand U4735 (N_4735,In_1741,In_745);
xor U4736 (N_4736,In_1753,In_114);
and U4737 (N_4737,In_2036,In_1797);
xor U4738 (N_4738,In_128,In_954);
nand U4739 (N_4739,In_586,In_389);
and U4740 (N_4740,In_1604,In_1117);
and U4741 (N_4741,In_719,In_411);
nand U4742 (N_4742,In_2042,In_614);
and U4743 (N_4743,In_114,In_485);
nor U4744 (N_4744,In_1543,In_1981);
xor U4745 (N_4745,In_692,In_2498);
nor U4746 (N_4746,In_496,In_1840);
or U4747 (N_4747,In_243,In_2345);
xor U4748 (N_4748,In_896,In_695);
and U4749 (N_4749,In_691,In_728);
and U4750 (N_4750,In_761,In_1596);
and U4751 (N_4751,In_1163,In_2140);
nor U4752 (N_4752,In_963,In_51);
and U4753 (N_4753,In_1812,In_51);
or U4754 (N_4754,In_246,In_1452);
and U4755 (N_4755,In_596,In_1303);
nor U4756 (N_4756,In_794,In_664);
nand U4757 (N_4757,In_1716,In_437);
nor U4758 (N_4758,In_76,In_237);
nor U4759 (N_4759,In_1865,In_95);
nor U4760 (N_4760,In_2282,In_1856);
nand U4761 (N_4761,In_1291,In_35);
and U4762 (N_4762,In_778,In_355);
and U4763 (N_4763,In_268,In_121);
xnor U4764 (N_4764,In_1830,In_1622);
nor U4765 (N_4765,In_852,In_1361);
or U4766 (N_4766,In_1108,In_2035);
xnor U4767 (N_4767,In_1510,In_1500);
xnor U4768 (N_4768,In_429,In_1451);
nand U4769 (N_4769,In_1586,In_2328);
and U4770 (N_4770,In_1147,In_2188);
nor U4771 (N_4771,In_892,In_2016);
nor U4772 (N_4772,In_2073,In_1979);
nor U4773 (N_4773,In_112,In_2151);
and U4774 (N_4774,In_2056,In_403);
or U4775 (N_4775,In_772,In_2019);
xnor U4776 (N_4776,In_385,In_1867);
and U4777 (N_4777,In_1315,In_988);
and U4778 (N_4778,In_841,In_846);
nor U4779 (N_4779,In_44,In_2050);
and U4780 (N_4780,In_805,In_1609);
and U4781 (N_4781,In_2215,In_424);
and U4782 (N_4782,In_1796,In_788);
nor U4783 (N_4783,In_2121,In_1708);
nand U4784 (N_4784,In_289,In_898);
nor U4785 (N_4785,In_507,In_1554);
and U4786 (N_4786,In_1147,In_1049);
xnor U4787 (N_4787,In_712,In_2055);
nor U4788 (N_4788,In_757,In_1105);
or U4789 (N_4789,In_1792,In_2041);
and U4790 (N_4790,In_987,In_1590);
xnor U4791 (N_4791,In_2116,In_1386);
nor U4792 (N_4792,In_1672,In_1607);
xnor U4793 (N_4793,In_263,In_1244);
nand U4794 (N_4794,In_740,In_2398);
and U4795 (N_4795,In_542,In_999);
nand U4796 (N_4796,In_507,In_2441);
and U4797 (N_4797,In_102,In_732);
nand U4798 (N_4798,In_497,In_594);
nand U4799 (N_4799,In_1614,In_618);
or U4800 (N_4800,In_417,In_2309);
nand U4801 (N_4801,In_998,In_573);
or U4802 (N_4802,In_2007,In_521);
nand U4803 (N_4803,In_471,In_2360);
nor U4804 (N_4804,In_403,In_1583);
or U4805 (N_4805,In_1521,In_1077);
or U4806 (N_4806,In_2076,In_2080);
and U4807 (N_4807,In_489,In_948);
and U4808 (N_4808,In_1623,In_2257);
nor U4809 (N_4809,In_260,In_731);
nand U4810 (N_4810,In_83,In_685);
nor U4811 (N_4811,In_2201,In_1424);
and U4812 (N_4812,In_2405,In_133);
and U4813 (N_4813,In_2299,In_2215);
or U4814 (N_4814,In_1983,In_150);
nand U4815 (N_4815,In_174,In_486);
or U4816 (N_4816,In_1548,In_68);
and U4817 (N_4817,In_2385,In_778);
nand U4818 (N_4818,In_2334,In_467);
or U4819 (N_4819,In_1248,In_1923);
nand U4820 (N_4820,In_926,In_2235);
nor U4821 (N_4821,In_1615,In_498);
or U4822 (N_4822,In_1795,In_1475);
nand U4823 (N_4823,In_1688,In_464);
nor U4824 (N_4824,In_447,In_59);
and U4825 (N_4825,In_241,In_1972);
nor U4826 (N_4826,In_1458,In_832);
nand U4827 (N_4827,In_5,In_2485);
or U4828 (N_4828,In_1209,In_1757);
nand U4829 (N_4829,In_1158,In_2061);
nand U4830 (N_4830,In_1433,In_2441);
or U4831 (N_4831,In_427,In_264);
nor U4832 (N_4832,In_2396,In_2217);
nand U4833 (N_4833,In_2376,In_2180);
xnor U4834 (N_4834,In_343,In_460);
nor U4835 (N_4835,In_520,In_2495);
nor U4836 (N_4836,In_1629,In_1171);
and U4837 (N_4837,In_2255,In_913);
or U4838 (N_4838,In_41,In_2258);
nand U4839 (N_4839,In_907,In_2021);
nand U4840 (N_4840,In_2366,In_1651);
or U4841 (N_4841,In_1194,In_1331);
or U4842 (N_4842,In_978,In_2260);
and U4843 (N_4843,In_303,In_2123);
nand U4844 (N_4844,In_2242,In_591);
or U4845 (N_4845,In_455,In_404);
or U4846 (N_4846,In_2167,In_982);
or U4847 (N_4847,In_2419,In_920);
nand U4848 (N_4848,In_2477,In_1568);
and U4849 (N_4849,In_766,In_1711);
nor U4850 (N_4850,In_1428,In_1225);
or U4851 (N_4851,In_1004,In_820);
or U4852 (N_4852,In_1714,In_95);
nand U4853 (N_4853,In_2157,In_1328);
or U4854 (N_4854,In_117,In_161);
xnor U4855 (N_4855,In_1442,In_640);
nor U4856 (N_4856,In_1310,In_2489);
nand U4857 (N_4857,In_1689,In_1377);
and U4858 (N_4858,In_496,In_1117);
nor U4859 (N_4859,In_1113,In_152);
or U4860 (N_4860,In_1397,In_1949);
nor U4861 (N_4861,In_470,In_1775);
or U4862 (N_4862,In_1825,In_2413);
nor U4863 (N_4863,In_1696,In_2439);
and U4864 (N_4864,In_2437,In_1666);
nor U4865 (N_4865,In_1594,In_1416);
and U4866 (N_4866,In_516,In_183);
nand U4867 (N_4867,In_209,In_1839);
and U4868 (N_4868,In_354,In_1642);
or U4869 (N_4869,In_48,In_1027);
nor U4870 (N_4870,In_1668,In_1136);
nor U4871 (N_4871,In_1867,In_2439);
or U4872 (N_4872,In_1490,In_1030);
nand U4873 (N_4873,In_151,In_1347);
and U4874 (N_4874,In_1683,In_2379);
nand U4875 (N_4875,In_229,In_1463);
xnor U4876 (N_4876,In_1546,In_701);
xnor U4877 (N_4877,In_1465,In_1539);
or U4878 (N_4878,In_1015,In_623);
and U4879 (N_4879,In_1533,In_1348);
or U4880 (N_4880,In_261,In_2262);
nor U4881 (N_4881,In_2144,In_2029);
or U4882 (N_4882,In_579,In_2433);
and U4883 (N_4883,In_2347,In_383);
or U4884 (N_4884,In_757,In_378);
or U4885 (N_4885,In_684,In_595);
and U4886 (N_4886,In_2089,In_1617);
or U4887 (N_4887,In_92,In_429);
nand U4888 (N_4888,In_609,In_1029);
nand U4889 (N_4889,In_635,In_2251);
nor U4890 (N_4890,In_1740,In_984);
nand U4891 (N_4891,In_630,In_167);
nor U4892 (N_4892,In_1940,In_686);
xor U4893 (N_4893,In_1649,In_178);
and U4894 (N_4894,In_1177,In_1460);
nand U4895 (N_4895,In_1130,In_2404);
nor U4896 (N_4896,In_1106,In_1734);
nand U4897 (N_4897,In_2451,In_1847);
or U4898 (N_4898,In_1574,In_1850);
xnor U4899 (N_4899,In_789,In_457);
nand U4900 (N_4900,In_1103,In_2158);
nor U4901 (N_4901,In_1880,In_819);
or U4902 (N_4902,In_1974,In_84);
nand U4903 (N_4903,In_2425,In_907);
nor U4904 (N_4904,In_1547,In_839);
xnor U4905 (N_4905,In_1197,In_701);
nand U4906 (N_4906,In_1683,In_1201);
xnor U4907 (N_4907,In_2301,In_835);
xor U4908 (N_4908,In_1715,In_34);
nand U4909 (N_4909,In_1736,In_2352);
xnor U4910 (N_4910,In_2271,In_852);
xor U4911 (N_4911,In_538,In_2290);
nand U4912 (N_4912,In_1792,In_1054);
and U4913 (N_4913,In_1279,In_344);
nand U4914 (N_4914,In_139,In_1518);
nand U4915 (N_4915,In_2438,In_302);
nand U4916 (N_4916,In_1739,In_540);
and U4917 (N_4917,In_181,In_2089);
and U4918 (N_4918,In_1522,In_2344);
and U4919 (N_4919,In_460,In_1843);
and U4920 (N_4920,In_2354,In_698);
or U4921 (N_4921,In_2153,In_2225);
and U4922 (N_4922,In_2488,In_801);
or U4923 (N_4923,In_1531,In_338);
and U4924 (N_4924,In_1598,In_1938);
nor U4925 (N_4925,In_2131,In_1943);
nand U4926 (N_4926,In_238,In_2471);
or U4927 (N_4927,In_2408,In_2108);
nand U4928 (N_4928,In_2465,In_1996);
or U4929 (N_4929,In_427,In_761);
nand U4930 (N_4930,In_32,In_1799);
nor U4931 (N_4931,In_1777,In_1482);
nand U4932 (N_4932,In_2490,In_1615);
or U4933 (N_4933,In_486,In_994);
and U4934 (N_4934,In_716,In_82);
or U4935 (N_4935,In_1545,In_1535);
nor U4936 (N_4936,In_689,In_225);
or U4937 (N_4937,In_1219,In_1711);
and U4938 (N_4938,In_1921,In_2208);
or U4939 (N_4939,In_1739,In_247);
or U4940 (N_4940,In_2198,In_182);
xnor U4941 (N_4941,In_1154,In_22);
nand U4942 (N_4942,In_1061,In_1871);
nor U4943 (N_4943,In_1506,In_1743);
nor U4944 (N_4944,In_1861,In_636);
xor U4945 (N_4945,In_1552,In_113);
and U4946 (N_4946,In_494,In_978);
or U4947 (N_4947,In_1662,In_1235);
nor U4948 (N_4948,In_1492,In_1329);
nor U4949 (N_4949,In_1333,In_1099);
or U4950 (N_4950,In_2188,In_741);
xnor U4951 (N_4951,In_1344,In_315);
nand U4952 (N_4952,In_713,In_665);
xor U4953 (N_4953,In_372,In_1507);
or U4954 (N_4954,In_1764,In_2085);
and U4955 (N_4955,In_310,In_805);
nor U4956 (N_4956,In_2257,In_296);
xor U4957 (N_4957,In_2302,In_1449);
or U4958 (N_4958,In_2140,In_471);
nor U4959 (N_4959,In_1516,In_220);
and U4960 (N_4960,In_808,In_1103);
and U4961 (N_4961,In_1955,In_1759);
nand U4962 (N_4962,In_2222,In_1120);
or U4963 (N_4963,In_2225,In_2239);
nor U4964 (N_4964,In_1301,In_2135);
or U4965 (N_4965,In_59,In_1796);
and U4966 (N_4966,In_676,In_650);
and U4967 (N_4967,In_1263,In_995);
or U4968 (N_4968,In_950,In_2308);
nor U4969 (N_4969,In_276,In_2367);
nor U4970 (N_4970,In_1535,In_1386);
nor U4971 (N_4971,In_989,In_1260);
nor U4972 (N_4972,In_1403,In_882);
or U4973 (N_4973,In_1459,In_202);
or U4974 (N_4974,In_2343,In_803);
xor U4975 (N_4975,In_1514,In_1737);
and U4976 (N_4976,In_353,In_1932);
nor U4977 (N_4977,In_592,In_1940);
xnor U4978 (N_4978,In_556,In_690);
or U4979 (N_4979,In_1041,In_1319);
nor U4980 (N_4980,In_829,In_159);
nor U4981 (N_4981,In_2326,In_2398);
nand U4982 (N_4982,In_718,In_2068);
nand U4983 (N_4983,In_599,In_2242);
or U4984 (N_4984,In_1023,In_1578);
xnor U4985 (N_4985,In_1353,In_1600);
and U4986 (N_4986,In_1728,In_899);
nor U4987 (N_4987,In_992,In_1347);
or U4988 (N_4988,In_1306,In_79);
xor U4989 (N_4989,In_2076,In_1870);
nor U4990 (N_4990,In_903,In_259);
nor U4991 (N_4991,In_228,In_1582);
and U4992 (N_4992,In_1207,In_664);
nor U4993 (N_4993,In_1299,In_2016);
nor U4994 (N_4994,In_120,In_1454);
and U4995 (N_4995,In_1692,In_394);
nor U4996 (N_4996,In_1877,In_2367);
nand U4997 (N_4997,In_2061,In_884);
or U4998 (N_4998,In_1443,In_1218);
and U4999 (N_4999,In_950,In_2394);
xor U5000 (N_5000,In_1994,In_638);
nor U5001 (N_5001,In_2115,In_481);
nor U5002 (N_5002,In_1807,In_2108);
nand U5003 (N_5003,In_191,In_2475);
nand U5004 (N_5004,In_1440,In_181);
and U5005 (N_5005,In_1804,In_1915);
nand U5006 (N_5006,In_1330,In_2064);
xnor U5007 (N_5007,In_1926,In_814);
nand U5008 (N_5008,In_2176,In_46);
xor U5009 (N_5009,In_43,In_724);
nand U5010 (N_5010,In_140,In_43);
or U5011 (N_5011,In_1615,In_176);
and U5012 (N_5012,In_1910,In_1850);
nor U5013 (N_5013,In_2189,In_150);
or U5014 (N_5014,In_1213,In_1319);
nor U5015 (N_5015,In_2233,In_753);
nor U5016 (N_5016,In_205,In_1027);
and U5017 (N_5017,In_737,In_1679);
nand U5018 (N_5018,In_1589,In_1532);
and U5019 (N_5019,In_64,In_1209);
nor U5020 (N_5020,In_1352,In_2347);
and U5021 (N_5021,In_983,In_544);
or U5022 (N_5022,In_712,In_1010);
xnor U5023 (N_5023,In_1740,In_1092);
nand U5024 (N_5024,In_41,In_769);
nand U5025 (N_5025,In_391,In_2043);
or U5026 (N_5026,In_2412,In_1867);
and U5027 (N_5027,In_169,In_1638);
and U5028 (N_5028,In_1002,In_1142);
nor U5029 (N_5029,In_1277,In_2199);
or U5030 (N_5030,In_1772,In_930);
nand U5031 (N_5031,In_591,In_710);
nand U5032 (N_5032,In_1601,In_1142);
and U5033 (N_5033,In_1874,In_1155);
nand U5034 (N_5034,In_1635,In_1723);
and U5035 (N_5035,In_421,In_571);
or U5036 (N_5036,In_1501,In_1692);
nand U5037 (N_5037,In_713,In_901);
nor U5038 (N_5038,In_1017,In_149);
xnor U5039 (N_5039,In_1936,In_164);
nand U5040 (N_5040,In_637,In_2300);
nor U5041 (N_5041,In_1874,In_759);
and U5042 (N_5042,In_2027,In_188);
and U5043 (N_5043,In_88,In_40);
nand U5044 (N_5044,In_2370,In_1911);
nor U5045 (N_5045,In_640,In_832);
nor U5046 (N_5046,In_884,In_1623);
or U5047 (N_5047,In_635,In_1409);
and U5048 (N_5048,In_389,In_693);
and U5049 (N_5049,In_807,In_469);
xnor U5050 (N_5050,In_1946,In_508);
xnor U5051 (N_5051,In_647,In_2478);
and U5052 (N_5052,In_917,In_1083);
or U5053 (N_5053,In_2452,In_324);
and U5054 (N_5054,In_906,In_1037);
or U5055 (N_5055,In_1176,In_64);
nor U5056 (N_5056,In_1014,In_2037);
nand U5057 (N_5057,In_1513,In_2138);
nand U5058 (N_5058,In_2268,In_770);
nor U5059 (N_5059,In_457,In_2294);
and U5060 (N_5060,In_2495,In_720);
nor U5061 (N_5061,In_1454,In_333);
nand U5062 (N_5062,In_1049,In_2215);
and U5063 (N_5063,In_514,In_874);
or U5064 (N_5064,In_987,In_2452);
nand U5065 (N_5065,In_130,In_2289);
and U5066 (N_5066,In_1086,In_2289);
nand U5067 (N_5067,In_2228,In_1753);
nor U5068 (N_5068,In_878,In_1963);
nand U5069 (N_5069,In_640,In_1646);
xor U5070 (N_5070,In_814,In_2180);
and U5071 (N_5071,In_1827,In_57);
nand U5072 (N_5072,In_21,In_2164);
xor U5073 (N_5073,In_1262,In_1774);
and U5074 (N_5074,In_940,In_712);
xnor U5075 (N_5075,In_1115,In_568);
nand U5076 (N_5076,In_240,In_2323);
or U5077 (N_5077,In_2382,In_2320);
or U5078 (N_5078,In_572,In_1029);
and U5079 (N_5079,In_2250,In_204);
or U5080 (N_5080,In_2363,In_1301);
and U5081 (N_5081,In_719,In_522);
nor U5082 (N_5082,In_2032,In_1861);
xor U5083 (N_5083,In_2425,In_187);
and U5084 (N_5084,In_1834,In_2387);
and U5085 (N_5085,In_1381,In_2411);
or U5086 (N_5086,In_2372,In_1042);
nand U5087 (N_5087,In_1174,In_1953);
or U5088 (N_5088,In_2160,In_1386);
or U5089 (N_5089,In_494,In_2254);
nand U5090 (N_5090,In_962,In_1117);
nand U5091 (N_5091,In_1896,In_1826);
nor U5092 (N_5092,In_32,In_1001);
nand U5093 (N_5093,In_1407,In_2318);
nor U5094 (N_5094,In_2182,In_2057);
nor U5095 (N_5095,In_1554,In_1517);
and U5096 (N_5096,In_598,In_1353);
nand U5097 (N_5097,In_2123,In_181);
and U5098 (N_5098,In_1853,In_2383);
or U5099 (N_5099,In_1134,In_1878);
and U5100 (N_5100,In_2464,In_1342);
xor U5101 (N_5101,In_1234,In_2398);
xor U5102 (N_5102,In_1457,In_452);
nand U5103 (N_5103,In_1192,In_1615);
xor U5104 (N_5104,In_1171,In_811);
nor U5105 (N_5105,In_645,In_1268);
nand U5106 (N_5106,In_2472,In_785);
and U5107 (N_5107,In_733,In_1202);
nor U5108 (N_5108,In_1588,In_1366);
or U5109 (N_5109,In_1090,In_2319);
or U5110 (N_5110,In_1172,In_1743);
nor U5111 (N_5111,In_1965,In_1961);
nand U5112 (N_5112,In_678,In_1240);
nand U5113 (N_5113,In_1299,In_1179);
and U5114 (N_5114,In_1548,In_1724);
nor U5115 (N_5115,In_643,In_202);
and U5116 (N_5116,In_952,In_1110);
or U5117 (N_5117,In_1968,In_1057);
xor U5118 (N_5118,In_408,In_848);
or U5119 (N_5119,In_1814,In_338);
xnor U5120 (N_5120,In_1620,In_2207);
xor U5121 (N_5121,In_938,In_1729);
nand U5122 (N_5122,In_749,In_540);
or U5123 (N_5123,In_447,In_193);
or U5124 (N_5124,In_959,In_1094);
nand U5125 (N_5125,In_2061,In_1084);
and U5126 (N_5126,In_1192,In_373);
nand U5127 (N_5127,In_116,In_1328);
nand U5128 (N_5128,In_842,In_859);
and U5129 (N_5129,In_719,In_1742);
or U5130 (N_5130,In_2190,In_1933);
and U5131 (N_5131,In_711,In_0);
nand U5132 (N_5132,In_219,In_480);
xor U5133 (N_5133,In_567,In_1257);
nand U5134 (N_5134,In_2182,In_2289);
xor U5135 (N_5135,In_412,In_711);
and U5136 (N_5136,In_1236,In_1122);
or U5137 (N_5137,In_2436,In_1263);
nand U5138 (N_5138,In_1774,In_1349);
xor U5139 (N_5139,In_2185,In_1072);
xnor U5140 (N_5140,In_1077,In_1595);
or U5141 (N_5141,In_1042,In_164);
and U5142 (N_5142,In_790,In_2265);
and U5143 (N_5143,In_843,In_374);
and U5144 (N_5144,In_1651,In_1748);
or U5145 (N_5145,In_1886,In_766);
xnor U5146 (N_5146,In_1733,In_804);
and U5147 (N_5147,In_487,In_1141);
or U5148 (N_5148,In_1793,In_707);
or U5149 (N_5149,In_168,In_422);
nor U5150 (N_5150,In_558,In_1837);
and U5151 (N_5151,In_1208,In_98);
nor U5152 (N_5152,In_1189,In_53);
nor U5153 (N_5153,In_1284,In_719);
xor U5154 (N_5154,In_1580,In_2240);
nand U5155 (N_5155,In_1269,In_1079);
nand U5156 (N_5156,In_801,In_308);
nand U5157 (N_5157,In_2217,In_1763);
or U5158 (N_5158,In_1790,In_1134);
or U5159 (N_5159,In_2380,In_782);
or U5160 (N_5160,In_1252,In_740);
nor U5161 (N_5161,In_106,In_310);
and U5162 (N_5162,In_816,In_446);
or U5163 (N_5163,In_975,In_2355);
or U5164 (N_5164,In_691,In_1287);
nor U5165 (N_5165,In_1013,In_1331);
nor U5166 (N_5166,In_33,In_448);
xor U5167 (N_5167,In_126,In_255);
and U5168 (N_5168,In_320,In_1705);
nand U5169 (N_5169,In_1548,In_2117);
nand U5170 (N_5170,In_1924,In_79);
and U5171 (N_5171,In_1305,In_2431);
or U5172 (N_5172,In_370,In_165);
nor U5173 (N_5173,In_2072,In_2470);
nor U5174 (N_5174,In_1719,In_1516);
or U5175 (N_5175,In_1552,In_115);
nor U5176 (N_5176,In_1496,In_1773);
nor U5177 (N_5177,In_2027,In_2361);
or U5178 (N_5178,In_1090,In_149);
and U5179 (N_5179,In_1179,In_540);
or U5180 (N_5180,In_1633,In_308);
nand U5181 (N_5181,In_2100,In_944);
nor U5182 (N_5182,In_2357,In_1095);
nor U5183 (N_5183,In_1820,In_1638);
or U5184 (N_5184,In_411,In_918);
and U5185 (N_5185,In_1921,In_2477);
or U5186 (N_5186,In_516,In_494);
or U5187 (N_5187,In_1876,In_2479);
or U5188 (N_5188,In_573,In_2114);
nor U5189 (N_5189,In_1077,In_823);
nor U5190 (N_5190,In_1797,In_1266);
xnor U5191 (N_5191,In_245,In_365);
nor U5192 (N_5192,In_1675,In_1726);
and U5193 (N_5193,In_921,In_846);
or U5194 (N_5194,In_383,In_586);
nor U5195 (N_5195,In_1815,In_1169);
and U5196 (N_5196,In_2295,In_1733);
xnor U5197 (N_5197,In_1676,In_959);
nor U5198 (N_5198,In_2173,In_1744);
and U5199 (N_5199,In_1103,In_1920);
nor U5200 (N_5200,In_1138,In_2101);
nand U5201 (N_5201,In_2122,In_1533);
nor U5202 (N_5202,In_95,In_580);
xnor U5203 (N_5203,In_1630,In_1113);
or U5204 (N_5204,In_781,In_2008);
or U5205 (N_5205,In_242,In_463);
nor U5206 (N_5206,In_1358,In_1455);
nand U5207 (N_5207,In_1589,In_1647);
nand U5208 (N_5208,In_2126,In_846);
or U5209 (N_5209,In_309,In_119);
and U5210 (N_5210,In_1771,In_1357);
or U5211 (N_5211,In_408,In_1978);
or U5212 (N_5212,In_2100,In_1077);
or U5213 (N_5213,In_598,In_1600);
nand U5214 (N_5214,In_1459,In_1795);
nor U5215 (N_5215,In_1685,In_498);
nor U5216 (N_5216,In_1355,In_1554);
and U5217 (N_5217,In_1364,In_2158);
nor U5218 (N_5218,In_1841,In_1384);
or U5219 (N_5219,In_808,In_763);
and U5220 (N_5220,In_2127,In_1148);
nand U5221 (N_5221,In_1298,In_2060);
nand U5222 (N_5222,In_917,In_1038);
and U5223 (N_5223,In_352,In_75);
nor U5224 (N_5224,In_710,In_1883);
and U5225 (N_5225,In_1133,In_1176);
nor U5226 (N_5226,In_511,In_1158);
and U5227 (N_5227,In_403,In_610);
nor U5228 (N_5228,In_1959,In_2452);
nand U5229 (N_5229,In_572,In_1977);
or U5230 (N_5230,In_2267,In_1737);
nor U5231 (N_5231,In_1129,In_1966);
or U5232 (N_5232,In_2150,In_935);
or U5233 (N_5233,In_1008,In_952);
xnor U5234 (N_5234,In_109,In_2230);
nor U5235 (N_5235,In_2473,In_1201);
nand U5236 (N_5236,In_1126,In_1368);
nand U5237 (N_5237,In_1853,In_1596);
nand U5238 (N_5238,In_2284,In_105);
nor U5239 (N_5239,In_605,In_1239);
xnor U5240 (N_5240,In_2299,In_56);
nor U5241 (N_5241,In_1870,In_710);
nor U5242 (N_5242,In_1814,In_2160);
xnor U5243 (N_5243,In_82,In_154);
or U5244 (N_5244,In_1452,In_398);
nor U5245 (N_5245,In_1200,In_2381);
xnor U5246 (N_5246,In_817,In_732);
and U5247 (N_5247,In_100,In_146);
xnor U5248 (N_5248,In_270,In_512);
or U5249 (N_5249,In_1935,In_22);
nand U5250 (N_5250,In_1253,In_2376);
or U5251 (N_5251,In_1497,In_1311);
nor U5252 (N_5252,In_1550,In_1458);
nor U5253 (N_5253,In_809,In_1698);
and U5254 (N_5254,In_1552,In_1952);
xor U5255 (N_5255,In_1086,In_676);
nand U5256 (N_5256,In_2377,In_921);
nand U5257 (N_5257,In_1735,In_2352);
nor U5258 (N_5258,In_1869,In_494);
nand U5259 (N_5259,In_868,In_2342);
xor U5260 (N_5260,In_1093,In_723);
nor U5261 (N_5261,In_2259,In_1273);
nor U5262 (N_5262,In_2485,In_596);
nand U5263 (N_5263,In_1345,In_17);
nand U5264 (N_5264,In_2240,In_713);
nor U5265 (N_5265,In_2105,In_561);
xnor U5266 (N_5266,In_1493,In_704);
nand U5267 (N_5267,In_1077,In_713);
nand U5268 (N_5268,In_1312,In_606);
or U5269 (N_5269,In_2477,In_445);
and U5270 (N_5270,In_308,In_1639);
or U5271 (N_5271,In_822,In_1980);
or U5272 (N_5272,In_506,In_1829);
nand U5273 (N_5273,In_734,In_2221);
nand U5274 (N_5274,In_2248,In_1433);
or U5275 (N_5275,In_1865,In_846);
and U5276 (N_5276,In_1197,In_281);
nand U5277 (N_5277,In_1568,In_1233);
and U5278 (N_5278,In_743,In_1851);
nor U5279 (N_5279,In_2445,In_760);
or U5280 (N_5280,In_1793,In_2401);
nor U5281 (N_5281,In_2218,In_429);
nand U5282 (N_5282,In_1905,In_2139);
nor U5283 (N_5283,In_1698,In_561);
xor U5284 (N_5284,In_334,In_1760);
or U5285 (N_5285,In_277,In_1786);
nor U5286 (N_5286,In_5,In_1414);
or U5287 (N_5287,In_967,In_1439);
and U5288 (N_5288,In_1436,In_827);
or U5289 (N_5289,In_320,In_1854);
nor U5290 (N_5290,In_1012,In_1420);
or U5291 (N_5291,In_1514,In_1080);
and U5292 (N_5292,In_1999,In_795);
and U5293 (N_5293,In_2094,In_1614);
nor U5294 (N_5294,In_286,In_53);
nand U5295 (N_5295,In_1328,In_231);
nand U5296 (N_5296,In_2002,In_170);
nand U5297 (N_5297,In_704,In_978);
nand U5298 (N_5298,In_1266,In_1404);
nor U5299 (N_5299,In_56,In_2090);
nor U5300 (N_5300,In_1776,In_522);
nor U5301 (N_5301,In_584,In_739);
nand U5302 (N_5302,In_1225,In_2369);
or U5303 (N_5303,In_650,In_184);
nor U5304 (N_5304,In_681,In_469);
xnor U5305 (N_5305,In_596,In_2115);
nor U5306 (N_5306,In_82,In_221);
or U5307 (N_5307,In_2480,In_311);
nand U5308 (N_5308,In_1426,In_1068);
or U5309 (N_5309,In_2422,In_1470);
or U5310 (N_5310,In_1005,In_1994);
xor U5311 (N_5311,In_605,In_479);
nor U5312 (N_5312,In_718,In_1068);
and U5313 (N_5313,In_683,In_724);
or U5314 (N_5314,In_1596,In_374);
xnor U5315 (N_5315,In_1735,In_1832);
and U5316 (N_5316,In_1956,In_1738);
or U5317 (N_5317,In_2321,In_2008);
xnor U5318 (N_5318,In_1862,In_91);
or U5319 (N_5319,In_2228,In_1689);
nor U5320 (N_5320,In_278,In_1117);
xor U5321 (N_5321,In_1475,In_939);
and U5322 (N_5322,In_440,In_2462);
nor U5323 (N_5323,In_2480,In_1302);
nor U5324 (N_5324,In_2263,In_1696);
or U5325 (N_5325,In_1845,In_1859);
and U5326 (N_5326,In_547,In_930);
nor U5327 (N_5327,In_2349,In_2387);
and U5328 (N_5328,In_1096,In_2318);
or U5329 (N_5329,In_1531,In_1837);
or U5330 (N_5330,In_2359,In_373);
nand U5331 (N_5331,In_2012,In_344);
and U5332 (N_5332,In_1983,In_1823);
and U5333 (N_5333,In_2475,In_1865);
nor U5334 (N_5334,In_945,In_310);
and U5335 (N_5335,In_700,In_129);
or U5336 (N_5336,In_1476,In_436);
nand U5337 (N_5337,In_702,In_1055);
xnor U5338 (N_5338,In_2297,In_1510);
and U5339 (N_5339,In_1684,In_454);
or U5340 (N_5340,In_623,In_1644);
and U5341 (N_5341,In_1781,In_1588);
or U5342 (N_5342,In_818,In_174);
xnor U5343 (N_5343,In_733,In_2459);
nand U5344 (N_5344,In_270,In_105);
and U5345 (N_5345,In_625,In_1772);
or U5346 (N_5346,In_2197,In_1355);
and U5347 (N_5347,In_1318,In_1710);
nor U5348 (N_5348,In_1404,In_2240);
and U5349 (N_5349,In_416,In_89);
nor U5350 (N_5350,In_1362,In_1619);
or U5351 (N_5351,In_2199,In_2019);
or U5352 (N_5352,In_336,In_1570);
or U5353 (N_5353,In_515,In_706);
xor U5354 (N_5354,In_2125,In_1497);
or U5355 (N_5355,In_961,In_1818);
or U5356 (N_5356,In_728,In_512);
nor U5357 (N_5357,In_461,In_1518);
nor U5358 (N_5358,In_1777,In_2078);
or U5359 (N_5359,In_415,In_442);
nand U5360 (N_5360,In_2229,In_1309);
nand U5361 (N_5361,In_755,In_1266);
nand U5362 (N_5362,In_42,In_1706);
nand U5363 (N_5363,In_192,In_2018);
and U5364 (N_5364,In_830,In_1703);
nor U5365 (N_5365,In_1353,In_1635);
or U5366 (N_5366,In_705,In_1137);
xor U5367 (N_5367,In_108,In_2478);
or U5368 (N_5368,In_1164,In_2043);
or U5369 (N_5369,In_2479,In_1932);
xnor U5370 (N_5370,In_1132,In_1186);
xor U5371 (N_5371,In_726,In_163);
or U5372 (N_5372,In_569,In_588);
and U5373 (N_5373,In_1831,In_1628);
nand U5374 (N_5374,In_1067,In_1736);
xnor U5375 (N_5375,In_2128,In_1465);
nand U5376 (N_5376,In_1120,In_2275);
or U5377 (N_5377,In_1227,In_1189);
and U5378 (N_5378,In_1368,In_531);
and U5379 (N_5379,In_885,In_228);
and U5380 (N_5380,In_753,In_39);
nor U5381 (N_5381,In_104,In_343);
or U5382 (N_5382,In_1319,In_1631);
and U5383 (N_5383,In_1253,In_411);
and U5384 (N_5384,In_988,In_1684);
and U5385 (N_5385,In_1012,In_2416);
nand U5386 (N_5386,In_1439,In_1156);
nand U5387 (N_5387,In_2367,In_2091);
nor U5388 (N_5388,In_1762,In_1031);
and U5389 (N_5389,In_183,In_1127);
or U5390 (N_5390,In_1933,In_1442);
or U5391 (N_5391,In_1731,In_2182);
nor U5392 (N_5392,In_385,In_138);
or U5393 (N_5393,In_1080,In_2107);
and U5394 (N_5394,In_1814,In_1068);
xnor U5395 (N_5395,In_902,In_541);
nand U5396 (N_5396,In_1973,In_2274);
or U5397 (N_5397,In_1478,In_1887);
nor U5398 (N_5398,In_861,In_479);
nand U5399 (N_5399,In_684,In_1923);
xnor U5400 (N_5400,In_2185,In_2498);
or U5401 (N_5401,In_1779,In_1346);
and U5402 (N_5402,In_1073,In_2192);
nor U5403 (N_5403,In_1735,In_2498);
nor U5404 (N_5404,In_2438,In_168);
nor U5405 (N_5405,In_1962,In_21);
or U5406 (N_5406,In_2119,In_1603);
or U5407 (N_5407,In_166,In_1331);
nor U5408 (N_5408,In_2139,In_1057);
nand U5409 (N_5409,In_2349,In_1058);
nor U5410 (N_5410,In_450,In_872);
and U5411 (N_5411,In_271,In_544);
nand U5412 (N_5412,In_2405,In_889);
nor U5413 (N_5413,In_963,In_1775);
nor U5414 (N_5414,In_1942,In_493);
and U5415 (N_5415,In_2439,In_598);
nand U5416 (N_5416,In_1161,In_1618);
nand U5417 (N_5417,In_412,In_1513);
nand U5418 (N_5418,In_708,In_2130);
or U5419 (N_5419,In_2070,In_1926);
or U5420 (N_5420,In_244,In_989);
and U5421 (N_5421,In_2253,In_603);
and U5422 (N_5422,In_2298,In_1618);
or U5423 (N_5423,In_1819,In_1246);
nand U5424 (N_5424,In_2425,In_1171);
and U5425 (N_5425,In_2319,In_1032);
or U5426 (N_5426,In_1227,In_319);
nor U5427 (N_5427,In_902,In_1101);
or U5428 (N_5428,In_1728,In_107);
nand U5429 (N_5429,In_486,In_341);
nand U5430 (N_5430,In_2156,In_1320);
and U5431 (N_5431,In_1542,In_575);
and U5432 (N_5432,In_919,In_2344);
and U5433 (N_5433,In_151,In_388);
and U5434 (N_5434,In_1135,In_647);
or U5435 (N_5435,In_925,In_2467);
nand U5436 (N_5436,In_2426,In_2146);
nand U5437 (N_5437,In_1143,In_733);
nor U5438 (N_5438,In_1041,In_279);
nand U5439 (N_5439,In_990,In_1658);
nor U5440 (N_5440,In_2159,In_62);
and U5441 (N_5441,In_19,In_1380);
xnor U5442 (N_5442,In_1889,In_149);
or U5443 (N_5443,In_2283,In_489);
and U5444 (N_5444,In_1257,In_2267);
and U5445 (N_5445,In_2456,In_313);
or U5446 (N_5446,In_1970,In_2001);
nand U5447 (N_5447,In_1042,In_531);
nor U5448 (N_5448,In_2439,In_1386);
or U5449 (N_5449,In_1704,In_134);
xnor U5450 (N_5450,In_2233,In_2109);
or U5451 (N_5451,In_1795,In_1695);
nor U5452 (N_5452,In_1054,In_1944);
or U5453 (N_5453,In_412,In_1321);
xnor U5454 (N_5454,In_764,In_666);
and U5455 (N_5455,In_2416,In_552);
or U5456 (N_5456,In_856,In_772);
and U5457 (N_5457,In_940,In_2444);
and U5458 (N_5458,In_855,In_2346);
xor U5459 (N_5459,In_1974,In_1035);
nor U5460 (N_5460,In_240,In_1761);
or U5461 (N_5461,In_447,In_227);
xor U5462 (N_5462,In_1749,In_1517);
nor U5463 (N_5463,In_180,In_2080);
and U5464 (N_5464,In_1263,In_1046);
nor U5465 (N_5465,In_821,In_1902);
nand U5466 (N_5466,In_619,In_1574);
and U5467 (N_5467,In_1662,In_455);
and U5468 (N_5468,In_2388,In_1446);
and U5469 (N_5469,In_342,In_1889);
nor U5470 (N_5470,In_1651,In_333);
xor U5471 (N_5471,In_1441,In_32);
xnor U5472 (N_5472,In_2159,In_1819);
and U5473 (N_5473,In_1435,In_1313);
or U5474 (N_5474,In_1640,In_774);
or U5475 (N_5475,In_1751,In_2314);
and U5476 (N_5476,In_504,In_925);
and U5477 (N_5477,In_942,In_2469);
nor U5478 (N_5478,In_1449,In_1049);
nor U5479 (N_5479,In_2070,In_1780);
nor U5480 (N_5480,In_1316,In_659);
or U5481 (N_5481,In_2404,In_1985);
and U5482 (N_5482,In_388,In_2121);
xor U5483 (N_5483,In_1077,In_1348);
nand U5484 (N_5484,In_415,In_2048);
nand U5485 (N_5485,In_917,In_2146);
nand U5486 (N_5486,In_1884,In_929);
nor U5487 (N_5487,In_1054,In_627);
and U5488 (N_5488,In_957,In_417);
nand U5489 (N_5489,In_1652,In_590);
and U5490 (N_5490,In_1041,In_904);
nor U5491 (N_5491,In_1810,In_1750);
or U5492 (N_5492,In_523,In_918);
nor U5493 (N_5493,In_536,In_338);
nand U5494 (N_5494,In_1814,In_551);
or U5495 (N_5495,In_1793,In_804);
nand U5496 (N_5496,In_2272,In_84);
and U5497 (N_5497,In_2335,In_490);
nor U5498 (N_5498,In_1969,In_2405);
nand U5499 (N_5499,In_1849,In_915);
nor U5500 (N_5500,In_1487,In_750);
nand U5501 (N_5501,In_864,In_48);
or U5502 (N_5502,In_1268,In_1142);
or U5503 (N_5503,In_1274,In_557);
nand U5504 (N_5504,In_429,In_2304);
and U5505 (N_5505,In_2148,In_1958);
or U5506 (N_5506,In_862,In_747);
nand U5507 (N_5507,In_544,In_936);
or U5508 (N_5508,In_1070,In_256);
nand U5509 (N_5509,In_2292,In_1929);
nand U5510 (N_5510,In_879,In_282);
or U5511 (N_5511,In_2439,In_1195);
nor U5512 (N_5512,In_2295,In_1409);
or U5513 (N_5513,In_2479,In_1755);
or U5514 (N_5514,In_1382,In_1961);
nor U5515 (N_5515,In_1327,In_1937);
nand U5516 (N_5516,In_1849,In_1801);
nand U5517 (N_5517,In_2337,In_2208);
nand U5518 (N_5518,In_1808,In_2135);
nor U5519 (N_5519,In_2450,In_1030);
xnor U5520 (N_5520,In_1267,In_1811);
nor U5521 (N_5521,In_1230,In_114);
nor U5522 (N_5522,In_290,In_483);
nor U5523 (N_5523,In_133,In_117);
nand U5524 (N_5524,In_422,In_1118);
nor U5525 (N_5525,In_2108,In_1440);
xor U5526 (N_5526,In_492,In_73);
nand U5527 (N_5527,In_324,In_702);
or U5528 (N_5528,In_1391,In_1105);
nor U5529 (N_5529,In_1270,In_1746);
nand U5530 (N_5530,In_2269,In_1897);
and U5531 (N_5531,In_1842,In_1317);
and U5532 (N_5532,In_572,In_12);
and U5533 (N_5533,In_80,In_2196);
or U5534 (N_5534,In_1773,In_1650);
and U5535 (N_5535,In_132,In_353);
and U5536 (N_5536,In_1616,In_1027);
xor U5537 (N_5537,In_528,In_1691);
xnor U5538 (N_5538,In_941,In_2200);
nor U5539 (N_5539,In_1,In_1033);
nand U5540 (N_5540,In_170,In_1876);
or U5541 (N_5541,In_833,In_741);
nand U5542 (N_5542,In_121,In_1106);
nand U5543 (N_5543,In_39,In_1761);
or U5544 (N_5544,In_2107,In_1858);
and U5545 (N_5545,In_2064,In_2424);
and U5546 (N_5546,In_1426,In_916);
and U5547 (N_5547,In_737,In_1095);
or U5548 (N_5548,In_206,In_1855);
and U5549 (N_5549,In_608,In_1304);
nand U5550 (N_5550,In_2333,In_2102);
or U5551 (N_5551,In_1385,In_2027);
nor U5552 (N_5552,In_411,In_1494);
nor U5553 (N_5553,In_2358,In_851);
nor U5554 (N_5554,In_1260,In_2218);
nor U5555 (N_5555,In_149,In_1440);
and U5556 (N_5556,In_2194,In_2263);
nand U5557 (N_5557,In_734,In_1226);
nor U5558 (N_5558,In_2421,In_1398);
and U5559 (N_5559,In_2084,In_1298);
nor U5560 (N_5560,In_1328,In_1810);
nand U5561 (N_5561,In_2243,In_1104);
and U5562 (N_5562,In_2097,In_1884);
nand U5563 (N_5563,In_2279,In_1554);
nand U5564 (N_5564,In_2057,In_1311);
and U5565 (N_5565,In_2263,In_2343);
or U5566 (N_5566,In_2148,In_389);
or U5567 (N_5567,In_143,In_532);
and U5568 (N_5568,In_2211,In_170);
and U5569 (N_5569,In_839,In_1256);
nor U5570 (N_5570,In_2002,In_2188);
and U5571 (N_5571,In_1325,In_2045);
nor U5572 (N_5572,In_1949,In_442);
or U5573 (N_5573,In_256,In_2235);
or U5574 (N_5574,In_252,In_2198);
nand U5575 (N_5575,In_1645,In_1553);
nor U5576 (N_5576,In_202,In_1355);
or U5577 (N_5577,In_118,In_1926);
nand U5578 (N_5578,In_796,In_585);
or U5579 (N_5579,In_942,In_623);
nor U5580 (N_5580,In_632,In_94);
or U5581 (N_5581,In_771,In_1912);
or U5582 (N_5582,In_1765,In_1217);
nand U5583 (N_5583,In_2197,In_1117);
nor U5584 (N_5584,In_2325,In_1090);
or U5585 (N_5585,In_1221,In_1129);
or U5586 (N_5586,In_627,In_2030);
xor U5587 (N_5587,In_2399,In_1738);
nand U5588 (N_5588,In_45,In_852);
and U5589 (N_5589,In_1164,In_460);
nor U5590 (N_5590,In_2304,In_1693);
and U5591 (N_5591,In_1756,In_72);
nand U5592 (N_5592,In_458,In_2108);
or U5593 (N_5593,In_739,In_172);
or U5594 (N_5594,In_850,In_24);
xor U5595 (N_5595,In_2148,In_1169);
nor U5596 (N_5596,In_1213,In_1860);
nand U5597 (N_5597,In_883,In_1155);
and U5598 (N_5598,In_682,In_379);
and U5599 (N_5599,In_97,In_1781);
nor U5600 (N_5600,In_1804,In_528);
nor U5601 (N_5601,In_683,In_1107);
xnor U5602 (N_5602,In_2219,In_2276);
nand U5603 (N_5603,In_1709,In_2183);
or U5604 (N_5604,In_437,In_1197);
or U5605 (N_5605,In_672,In_1528);
xor U5606 (N_5606,In_1613,In_1177);
and U5607 (N_5607,In_476,In_656);
xor U5608 (N_5608,In_543,In_2229);
and U5609 (N_5609,In_1451,In_108);
or U5610 (N_5610,In_1330,In_1696);
and U5611 (N_5611,In_1195,In_575);
and U5612 (N_5612,In_1447,In_1550);
nor U5613 (N_5613,In_357,In_635);
and U5614 (N_5614,In_1701,In_1390);
and U5615 (N_5615,In_2000,In_2113);
and U5616 (N_5616,In_2074,In_61);
nand U5617 (N_5617,In_1202,In_2299);
xor U5618 (N_5618,In_1931,In_1225);
nand U5619 (N_5619,In_1047,In_1686);
nand U5620 (N_5620,In_696,In_2001);
nor U5621 (N_5621,In_501,In_169);
nor U5622 (N_5622,In_1145,In_1904);
nor U5623 (N_5623,In_1542,In_457);
nand U5624 (N_5624,In_695,In_963);
nand U5625 (N_5625,In_2462,In_1882);
xor U5626 (N_5626,In_570,In_2445);
nor U5627 (N_5627,In_454,In_530);
and U5628 (N_5628,In_2324,In_141);
and U5629 (N_5629,In_57,In_2092);
and U5630 (N_5630,In_1295,In_2449);
and U5631 (N_5631,In_1442,In_1411);
nand U5632 (N_5632,In_1365,In_322);
and U5633 (N_5633,In_1101,In_1585);
nand U5634 (N_5634,In_779,In_1476);
nor U5635 (N_5635,In_336,In_1539);
or U5636 (N_5636,In_529,In_1248);
or U5637 (N_5637,In_1706,In_1951);
and U5638 (N_5638,In_2298,In_1911);
and U5639 (N_5639,In_1364,In_1995);
nor U5640 (N_5640,In_1417,In_1513);
and U5641 (N_5641,In_752,In_1345);
and U5642 (N_5642,In_1187,In_1762);
nand U5643 (N_5643,In_655,In_675);
or U5644 (N_5644,In_2158,In_1234);
nand U5645 (N_5645,In_2132,In_1872);
or U5646 (N_5646,In_805,In_1135);
and U5647 (N_5647,In_866,In_832);
nor U5648 (N_5648,In_296,In_804);
and U5649 (N_5649,In_2223,In_908);
or U5650 (N_5650,In_628,In_1940);
nor U5651 (N_5651,In_1853,In_2279);
xor U5652 (N_5652,In_2474,In_234);
nor U5653 (N_5653,In_217,In_2187);
nor U5654 (N_5654,In_946,In_2494);
or U5655 (N_5655,In_874,In_782);
nand U5656 (N_5656,In_1336,In_484);
and U5657 (N_5657,In_528,In_1247);
nand U5658 (N_5658,In_248,In_1846);
nor U5659 (N_5659,In_372,In_2490);
or U5660 (N_5660,In_541,In_1561);
nand U5661 (N_5661,In_361,In_1454);
or U5662 (N_5662,In_2045,In_2448);
and U5663 (N_5663,In_1524,In_30);
xnor U5664 (N_5664,In_821,In_628);
or U5665 (N_5665,In_1984,In_1492);
xor U5666 (N_5666,In_1484,In_2379);
nor U5667 (N_5667,In_1066,In_1312);
nor U5668 (N_5668,In_1815,In_2067);
nor U5669 (N_5669,In_129,In_909);
nor U5670 (N_5670,In_597,In_2464);
nor U5671 (N_5671,In_2109,In_1664);
xor U5672 (N_5672,In_485,In_849);
and U5673 (N_5673,In_1147,In_419);
or U5674 (N_5674,In_418,In_113);
nand U5675 (N_5675,In_1073,In_1749);
and U5676 (N_5676,In_2337,In_427);
or U5677 (N_5677,In_2240,In_1467);
nor U5678 (N_5678,In_2017,In_855);
or U5679 (N_5679,In_671,In_1234);
and U5680 (N_5680,In_422,In_188);
nor U5681 (N_5681,In_1043,In_1654);
and U5682 (N_5682,In_1824,In_583);
or U5683 (N_5683,In_1547,In_1460);
nor U5684 (N_5684,In_1092,In_980);
or U5685 (N_5685,In_2134,In_2179);
or U5686 (N_5686,In_769,In_777);
or U5687 (N_5687,In_1789,In_1060);
and U5688 (N_5688,In_762,In_1436);
or U5689 (N_5689,In_1110,In_1839);
and U5690 (N_5690,In_2159,In_1651);
nor U5691 (N_5691,In_1845,In_2247);
nand U5692 (N_5692,In_2023,In_1717);
xor U5693 (N_5693,In_2072,In_75);
or U5694 (N_5694,In_1467,In_29);
and U5695 (N_5695,In_1719,In_1708);
or U5696 (N_5696,In_315,In_5);
or U5697 (N_5697,In_1898,In_1895);
nand U5698 (N_5698,In_2390,In_1307);
xor U5699 (N_5699,In_1239,In_1581);
or U5700 (N_5700,In_1722,In_95);
xor U5701 (N_5701,In_572,In_1405);
nand U5702 (N_5702,In_2169,In_1174);
nor U5703 (N_5703,In_856,In_1810);
or U5704 (N_5704,In_431,In_531);
and U5705 (N_5705,In_326,In_1169);
and U5706 (N_5706,In_1056,In_1533);
nor U5707 (N_5707,In_2111,In_1899);
and U5708 (N_5708,In_673,In_606);
nor U5709 (N_5709,In_1778,In_1852);
nor U5710 (N_5710,In_684,In_1157);
nor U5711 (N_5711,In_156,In_1532);
nand U5712 (N_5712,In_1981,In_1638);
nor U5713 (N_5713,In_1035,In_2195);
or U5714 (N_5714,In_2301,In_2020);
nor U5715 (N_5715,In_1260,In_2208);
and U5716 (N_5716,In_2047,In_705);
or U5717 (N_5717,In_111,In_1813);
or U5718 (N_5718,In_2268,In_715);
or U5719 (N_5719,In_2010,In_2037);
nor U5720 (N_5720,In_1006,In_1954);
or U5721 (N_5721,In_1697,In_1418);
nand U5722 (N_5722,In_739,In_1807);
and U5723 (N_5723,In_2322,In_2260);
and U5724 (N_5724,In_2093,In_353);
and U5725 (N_5725,In_2023,In_390);
xor U5726 (N_5726,In_1857,In_108);
nand U5727 (N_5727,In_144,In_979);
or U5728 (N_5728,In_1110,In_849);
or U5729 (N_5729,In_2050,In_1752);
nor U5730 (N_5730,In_1822,In_875);
nand U5731 (N_5731,In_1926,In_391);
or U5732 (N_5732,In_631,In_1226);
and U5733 (N_5733,In_1725,In_1350);
nand U5734 (N_5734,In_1859,In_1560);
and U5735 (N_5735,In_2165,In_970);
nor U5736 (N_5736,In_813,In_317);
nand U5737 (N_5737,In_840,In_1666);
or U5738 (N_5738,In_1508,In_271);
and U5739 (N_5739,In_1664,In_2495);
nand U5740 (N_5740,In_1727,In_224);
and U5741 (N_5741,In_1123,In_1098);
nand U5742 (N_5742,In_2373,In_1878);
xnor U5743 (N_5743,In_2107,In_904);
or U5744 (N_5744,In_476,In_1091);
nor U5745 (N_5745,In_1345,In_1171);
and U5746 (N_5746,In_1610,In_287);
xor U5747 (N_5747,In_1375,In_80);
xor U5748 (N_5748,In_47,In_20);
and U5749 (N_5749,In_1818,In_179);
xor U5750 (N_5750,In_225,In_646);
or U5751 (N_5751,In_2355,In_1766);
or U5752 (N_5752,In_1181,In_2336);
xnor U5753 (N_5753,In_346,In_2284);
nor U5754 (N_5754,In_1254,In_270);
xnor U5755 (N_5755,In_1021,In_726);
or U5756 (N_5756,In_1659,In_332);
or U5757 (N_5757,In_625,In_2214);
or U5758 (N_5758,In_1662,In_1958);
or U5759 (N_5759,In_1941,In_1707);
xnor U5760 (N_5760,In_2057,In_20);
or U5761 (N_5761,In_1578,In_2106);
nand U5762 (N_5762,In_1126,In_840);
nand U5763 (N_5763,In_963,In_299);
and U5764 (N_5764,In_1185,In_90);
or U5765 (N_5765,In_27,In_1141);
or U5766 (N_5766,In_1550,In_795);
nand U5767 (N_5767,In_2119,In_1989);
and U5768 (N_5768,In_1720,In_1983);
nand U5769 (N_5769,In_1668,In_1377);
nand U5770 (N_5770,In_2337,In_2136);
nand U5771 (N_5771,In_2404,In_756);
or U5772 (N_5772,In_1207,In_815);
nand U5773 (N_5773,In_842,In_2004);
and U5774 (N_5774,In_225,In_134);
nor U5775 (N_5775,In_1758,In_309);
nand U5776 (N_5776,In_744,In_1364);
nor U5777 (N_5777,In_367,In_2473);
nor U5778 (N_5778,In_759,In_470);
and U5779 (N_5779,In_40,In_1056);
xnor U5780 (N_5780,In_91,In_619);
nor U5781 (N_5781,In_1314,In_689);
nand U5782 (N_5782,In_607,In_573);
xor U5783 (N_5783,In_217,In_621);
nand U5784 (N_5784,In_944,In_1200);
and U5785 (N_5785,In_1726,In_208);
xor U5786 (N_5786,In_224,In_1389);
and U5787 (N_5787,In_592,In_1819);
nand U5788 (N_5788,In_2119,In_454);
and U5789 (N_5789,In_2159,In_1012);
nand U5790 (N_5790,In_355,In_1184);
nand U5791 (N_5791,In_886,In_188);
or U5792 (N_5792,In_2192,In_2071);
or U5793 (N_5793,In_2275,In_1976);
or U5794 (N_5794,In_1771,In_1685);
or U5795 (N_5795,In_1176,In_423);
nand U5796 (N_5796,In_471,In_1229);
or U5797 (N_5797,In_421,In_1180);
or U5798 (N_5798,In_1164,In_1511);
and U5799 (N_5799,In_2130,In_82);
nor U5800 (N_5800,In_1091,In_261);
xnor U5801 (N_5801,In_1353,In_2089);
nand U5802 (N_5802,In_576,In_795);
nand U5803 (N_5803,In_2476,In_1508);
or U5804 (N_5804,In_1071,In_2031);
nand U5805 (N_5805,In_2020,In_1387);
nand U5806 (N_5806,In_1913,In_1922);
nand U5807 (N_5807,In_1366,In_45);
nand U5808 (N_5808,In_263,In_32);
or U5809 (N_5809,In_2297,In_1657);
nand U5810 (N_5810,In_1986,In_29);
nor U5811 (N_5811,In_585,In_488);
and U5812 (N_5812,In_1146,In_2104);
nand U5813 (N_5813,In_653,In_583);
nor U5814 (N_5814,In_1427,In_1871);
xor U5815 (N_5815,In_1615,In_1940);
or U5816 (N_5816,In_1694,In_879);
nor U5817 (N_5817,In_1667,In_2211);
and U5818 (N_5818,In_405,In_84);
nor U5819 (N_5819,In_565,In_846);
nand U5820 (N_5820,In_2287,In_1123);
nor U5821 (N_5821,In_2167,In_1532);
and U5822 (N_5822,In_1934,In_1580);
nor U5823 (N_5823,In_1349,In_2388);
xor U5824 (N_5824,In_488,In_391);
or U5825 (N_5825,In_1369,In_173);
and U5826 (N_5826,In_677,In_328);
or U5827 (N_5827,In_2096,In_436);
nor U5828 (N_5828,In_715,In_1776);
or U5829 (N_5829,In_1199,In_1363);
and U5830 (N_5830,In_1501,In_2);
nor U5831 (N_5831,In_387,In_1259);
nor U5832 (N_5832,In_466,In_1356);
xnor U5833 (N_5833,In_1044,In_913);
and U5834 (N_5834,In_2173,In_1319);
nor U5835 (N_5835,In_1255,In_1181);
or U5836 (N_5836,In_2313,In_87);
or U5837 (N_5837,In_760,In_1529);
or U5838 (N_5838,In_361,In_2384);
nand U5839 (N_5839,In_1866,In_1631);
or U5840 (N_5840,In_760,In_1684);
xnor U5841 (N_5841,In_1111,In_490);
or U5842 (N_5842,In_2314,In_1162);
nor U5843 (N_5843,In_908,In_1959);
xor U5844 (N_5844,In_742,In_1278);
xor U5845 (N_5845,In_836,In_2028);
nand U5846 (N_5846,In_423,In_1462);
and U5847 (N_5847,In_1977,In_574);
and U5848 (N_5848,In_2311,In_1604);
nor U5849 (N_5849,In_1093,In_800);
and U5850 (N_5850,In_1516,In_1900);
and U5851 (N_5851,In_341,In_491);
nand U5852 (N_5852,In_165,In_1603);
nand U5853 (N_5853,In_2316,In_2260);
nor U5854 (N_5854,In_1117,In_1317);
nor U5855 (N_5855,In_262,In_2438);
nor U5856 (N_5856,In_2364,In_1807);
xor U5857 (N_5857,In_2038,In_1008);
xor U5858 (N_5858,In_2236,In_1119);
nand U5859 (N_5859,In_1749,In_1242);
and U5860 (N_5860,In_2182,In_490);
and U5861 (N_5861,In_839,In_428);
and U5862 (N_5862,In_359,In_1535);
nand U5863 (N_5863,In_383,In_2170);
or U5864 (N_5864,In_948,In_393);
nand U5865 (N_5865,In_3,In_2496);
or U5866 (N_5866,In_1907,In_661);
or U5867 (N_5867,In_344,In_48);
nor U5868 (N_5868,In_1064,In_2457);
or U5869 (N_5869,In_506,In_2033);
nand U5870 (N_5870,In_1218,In_1913);
nand U5871 (N_5871,In_1254,In_541);
xnor U5872 (N_5872,In_1767,In_1195);
and U5873 (N_5873,In_1277,In_2214);
nand U5874 (N_5874,In_1462,In_260);
xor U5875 (N_5875,In_1102,In_2069);
nor U5876 (N_5876,In_109,In_998);
nand U5877 (N_5877,In_960,In_2372);
nor U5878 (N_5878,In_1754,In_766);
xor U5879 (N_5879,In_1227,In_1095);
nor U5880 (N_5880,In_1150,In_2485);
xnor U5881 (N_5881,In_961,In_1161);
nor U5882 (N_5882,In_584,In_680);
nand U5883 (N_5883,In_543,In_1725);
nand U5884 (N_5884,In_1430,In_1565);
xor U5885 (N_5885,In_711,In_425);
nand U5886 (N_5886,In_2194,In_987);
and U5887 (N_5887,In_1058,In_942);
nor U5888 (N_5888,In_1781,In_1944);
or U5889 (N_5889,In_1398,In_2492);
nand U5890 (N_5890,In_940,In_868);
nor U5891 (N_5891,In_67,In_2386);
nand U5892 (N_5892,In_1030,In_1567);
or U5893 (N_5893,In_1742,In_994);
and U5894 (N_5894,In_1488,In_2499);
and U5895 (N_5895,In_661,In_2384);
xor U5896 (N_5896,In_1784,In_2497);
or U5897 (N_5897,In_1303,In_556);
nand U5898 (N_5898,In_57,In_666);
nor U5899 (N_5899,In_2348,In_1731);
nand U5900 (N_5900,In_380,In_1917);
xor U5901 (N_5901,In_901,In_124);
nor U5902 (N_5902,In_2240,In_1280);
or U5903 (N_5903,In_77,In_619);
or U5904 (N_5904,In_701,In_554);
nand U5905 (N_5905,In_1037,In_1364);
and U5906 (N_5906,In_1685,In_2258);
nand U5907 (N_5907,In_285,In_1430);
or U5908 (N_5908,In_822,In_1278);
nand U5909 (N_5909,In_904,In_712);
and U5910 (N_5910,In_1067,In_1857);
nand U5911 (N_5911,In_1880,In_362);
nand U5912 (N_5912,In_1341,In_1825);
and U5913 (N_5913,In_651,In_1151);
or U5914 (N_5914,In_2330,In_1665);
or U5915 (N_5915,In_1956,In_561);
or U5916 (N_5916,In_281,In_252);
xnor U5917 (N_5917,In_1739,In_663);
nor U5918 (N_5918,In_491,In_704);
or U5919 (N_5919,In_235,In_1427);
and U5920 (N_5920,In_1944,In_2395);
or U5921 (N_5921,In_494,In_1840);
or U5922 (N_5922,In_785,In_543);
and U5923 (N_5923,In_983,In_2135);
nand U5924 (N_5924,In_2366,In_2174);
and U5925 (N_5925,In_597,In_826);
nand U5926 (N_5926,In_1068,In_1428);
or U5927 (N_5927,In_2071,In_588);
and U5928 (N_5928,In_58,In_1751);
or U5929 (N_5929,In_2041,In_2319);
or U5930 (N_5930,In_623,In_191);
xor U5931 (N_5931,In_2252,In_63);
nor U5932 (N_5932,In_233,In_2240);
or U5933 (N_5933,In_1923,In_1381);
or U5934 (N_5934,In_97,In_2282);
nand U5935 (N_5935,In_1226,In_558);
nand U5936 (N_5936,In_1072,In_1126);
and U5937 (N_5937,In_262,In_1400);
nand U5938 (N_5938,In_734,In_1275);
nor U5939 (N_5939,In_1611,In_1271);
or U5940 (N_5940,In_109,In_53);
nand U5941 (N_5941,In_338,In_606);
or U5942 (N_5942,In_737,In_467);
nand U5943 (N_5943,In_439,In_1302);
nor U5944 (N_5944,In_500,In_731);
or U5945 (N_5945,In_319,In_366);
nor U5946 (N_5946,In_1189,In_1798);
xnor U5947 (N_5947,In_1801,In_1911);
nor U5948 (N_5948,In_43,In_794);
nand U5949 (N_5949,In_480,In_519);
xnor U5950 (N_5950,In_383,In_1846);
or U5951 (N_5951,In_1013,In_1759);
or U5952 (N_5952,In_275,In_2124);
nor U5953 (N_5953,In_515,In_762);
nand U5954 (N_5954,In_1006,In_1791);
and U5955 (N_5955,In_880,In_2142);
nor U5956 (N_5956,In_2159,In_2162);
nand U5957 (N_5957,In_1959,In_959);
xnor U5958 (N_5958,In_1219,In_205);
and U5959 (N_5959,In_2251,In_1823);
nor U5960 (N_5960,In_2019,In_1547);
or U5961 (N_5961,In_157,In_2456);
xnor U5962 (N_5962,In_1035,In_1613);
nand U5963 (N_5963,In_1197,In_1919);
and U5964 (N_5964,In_1587,In_350);
nand U5965 (N_5965,In_2205,In_1535);
and U5966 (N_5966,In_2098,In_454);
nand U5967 (N_5967,In_2149,In_990);
and U5968 (N_5968,In_569,In_1417);
and U5969 (N_5969,In_1469,In_2231);
or U5970 (N_5970,In_2398,In_372);
nand U5971 (N_5971,In_2250,In_1559);
and U5972 (N_5972,In_372,In_53);
and U5973 (N_5973,In_2114,In_403);
nand U5974 (N_5974,In_1357,In_1182);
and U5975 (N_5975,In_1964,In_2365);
nor U5976 (N_5976,In_344,In_982);
nand U5977 (N_5977,In_1492,In_821);
and U5978 (N_5978,In_1592,In_1796);
nor U5979 (N_5979,In_1170,In_1076);
or U5980 (N_5980,In_2376,In_2283);
nand U5981 (N_5981,In_2002,In_1328);
nor U5982 (N_5982,In_1665,In_2495);
nor U5983 (N_5983,In_1028,In_477);
or U5984 (N_5984,In_1697,In_913);
or U5985 (N_5985,In_2018,In_2154);
or U5986 (N_5986,In_2480,In_2196);
or U5987 (N_5987,In_2107,In_94);
and U5988 (N_5988,In_1478,In_962);
nand U5989 (N_5989,In_784,In_271);
nor U5990 (N_5990,In_848,In_2457);
and U5991 (N_5991,In_1274,In_917);
nor U5992 (N_5992,In_867,In_1018);
nand U5993 (N_5993,In_1419,In_1594);
or U5994 (N_5994,In_637,In_593);
nand U5995 (N_5995,In_935,In_990);
nand U5996 (N_5996,In_1185,In_551);
and U5997 (N_5997,In_1090,In_769);
nand U5998 (N_5998,In_1993,In_1198);
and U5999 (N_5999,In_2189,In_1856);
nand U6000 (N_6000,In_2166,In_684);
xor U6001 (N_6001,In_2066,In_1427);
nand U6002 (N_6002,In_1433,In_1805);
and U6003 (N_6003,In_1412,In_1430);
xnor U6004 (N_6004,In_793,In_135);
or U6005 (N_6005,In_1121,In_1089);
xnor U6006 (N_6006,In_1576,In_1196);
or U6007 (N_6007,In_443,In_278);
nand U6008 (N_6008,In_477,In_1511);
and U6009 (N_6009,In_2251,In_339);
and U6010 (N_6010,In_1447,In_1279);
nand U6011 (N_6011,In_1434,In_1445);
or U6012 (N_6012,In_2421,In_497);
and U6013 (N_6013,In_1877,In_428);
xnor U6014 (N_6014,In_43,In_2494);
nor U6015 (N_6015,In_1464,In_734);
nor U6016 (N_6016,In_509,In_1748);
nand U6017 (N_6017,In_1455,In_607);
or U6018 (N_6018,In_2355,In_153);
nand U6019 (N_6019,In_2395,In_797);
and U6020 (N_6020,In_1062,In_1242);
nor U6021 (N_6021,In_981,In_1737);
or U6022 (N_6022,In_2003,In_2427);
xor U6023 (N_6023,In_1036,In_717);
and U6024 (N_6024,In_777,In_232);
nor U6025 (N_6025,In_968,In_729);
nor U6026 (N_6026,In_1223,In_1911);
nor U6027 (N_6027,In_2404,In_659);
nand U6028 (N_6028,In_513,In_2372);
nand U6029 (N_6029,In_1267,In_771);
and U6030 (N_6030,In_1450,In_934);
or U6031 (N_6031,In_702,In_360);
nand U6032 (N_6032,In_1037,In_2158);
nor U6033 (N_6033,In_2182,In_285);
or U6034 (N_6034,In_846,In_1963);
nor U6035 (N_6035,In_1369,In_2257);
nand U6036 (N_6036,In_1633,In_671);
nand U6037 (N_6037,In_874,In_1770);
nand U6038 (N_6038,In_2466,In_1709);
nor U6039 (N_6039,In_119,In_623);
nand U6040 (N_6040,In_2012,In_1180);
or U6041 (N_6041,In_1479,In_303);
and U6042 (N_6042,In_385,In_655);
or U6043 (N_6043,In_1534,In_45);
and U6044 (N_6044,In_1115,In_1122);
and U6045 (N_6045,In_902,In_1147);
and U6046 (N_6046,In_585,In_1739);
and U6047 (N_6047,In_451,In_32);
xnor U6048 (N_6048,In_2026,In_2063);
xnor U6049 (N_6049,In_879,In_1324);
and U6050 (N_6050,In_2215,In_702);
and U6051 (N_6051,In_1506,In_450);
nor U6052 (N_6052,In_155,In_2241);
or U6053 (N_6053,In_1534,In_2168);
and U6054 (N_6054,In_1035,In_1786);
nand U6055 (N_6055,In_1658,In_1858);
nor U6056 (N_6056,In_517,In_2088);
nand U6057 (N_6057,In_186,In_584);
or U6058 (N_6058,In_1027,In_1990);
and U6059 (N_6059,In_400,In_2344);
nand U6060 (N_6060,In_2235,In_1573);
xor U6061 (N_6061,In_1775,In_2447);
or U6062 (N_6062,In_1222,In_1223);
or U6063 (N_6063,In_1219,In_2321);
nor U6064 (N_6064,In_1400,In_1325);
or U6065 (N_6065,In_1934,In_1181);
or U6066 (N_6066,In_1105,In_131);
nor U6067 (N_6067,In_45,In_343);
nor U6068 (N_6068,In_1704,In_2435);
nand U6069 (N_6069,In_1256,In_452);
or U6070 (N_6070,In_1581,In_1727);
nand U6071 (N_6071,In_1122,In_1760);
nand U6072 (N_6072,In_128,In_456);
nor U6073 (N_6073,In_541,In_1086);
nor U6074 (N_6074,In_1620,In_2217);
or U6075 (N_6075,In_192,In_472);
nor U6076 (N_6076,In_2086,In_266);
and U6077 (N_6077,In_681,In_232);
or U6078 (N_6078,In_654,In_1134);
and U6079 (N_6079,In_322,In_539);
nand U6080 (N_6080,In_2395,In_2438);
or U6081 (N_6081,In_1456,In_526);
or U6082 (N_6082,In_603,In_699);
xor U6083 (N_6083,In_377,In_508);
and U6084 (N_6084,In_1176,In_824);
nor U6085 (N_6085,In_2330,In_2497);
nand U6086 (N_6086,In_359,In_2063);
nand U6087 (N_6087,In_2217,In_2088);
and U6088 (N_6088,In_2095,In_2016);
and U6089 (N_6089,In_1024,In_1058);
nor U6090 (N_6090,In_1960,In_1377);
nor U6091 (N_6091,In_538,In_674);
nor U6092 (N_6092,In_950,In_1954);
and U6093 (N_6093,In_1966,In_1562);
nor U6094 (N_6094,In_2157,In_1812);
or U6095 (N_6095,In_270,In_1225);
nor U6096 (N_6096,In_2160,In_110);
or U6097 (N_6097,In_569,In_821);
nand U6098 (N_6098,In_1548,In_2221);
nor U6099 (N_6099,In_2148,In_644);
and U6100 (N_6100,In_667,In_1326);
and U6101 (N_6101,In_1065,In_2480);
or U6102 (N_6102,In_148,In_2308);
and U6103 (N_6103,In_1591,In_1336);
or U6104 (N_6104,In_1395,In_227);
nand U6105 (N_6105,In_1647,In_2117);
nand U6106 (N_6106,In_2199,In_1278);
xor U6107 (N_6107,In_1208,In_2066);
and U6108 (N_6108,In_1440,In_460);
or U6109 (N_6109,In_1241,In_635);
xor U6110 (N_6110,In_568,In_1438);
and U6111 (N_6111,In_586,In_1012);
nor U6112 (N_6112,In_129,In_2256);
and U6113 (N_6113,In_1508,In_13);
or U6114 (N_6114,In_1320,In_818);
nand U6115 (N_6115,In_2425,In_2074);
xnor U6116 (N_6116,In_2377,In_1568);
nand U6117 (N_6117,In_1590,In_1565);
nand U6118 (N_6118,In_448,In_523);
or U6119 (N_6119,In_86,In_863);
nand U6120 (N_6120,In_1820,In_2352);
or U6121 (N_6121,In_426,In_1290);
or U6122 (N_6122,In_1487,In_1385);
nor U6123 (N_6123,In_1463,In_550);
nand U6124 (N_6124,In_786,In_369);
or U6125 (N_6125,In_1094,In_384);
or U6126 (N_6126,In_2122,In_1136);
or U6127 (N_6127,In_924,In_98);
or U6128 (N_6128,In_444,In_935);
and U6129 (N_6129,In_762,In_1091);
or U6130 (N_6130,In_1752,In_1987);
xor U6131 (N_6131,In_787,In_688);
nand U6132 (N_6132,In_374,In_273);
nor U6133 (N_6133,In_2487,In_2289);
and U6134 (N_6134,In_1308,In_455);
nand U6135 (N_6135,In_993,In_602);
and U6136 (N_6136,In_1643,In_1382);
xnor U6137 (N_6137,In_1635,In_605);
nand U6138 (N_6138,In_1916,In_393);
xnor U6139 (N_6139,In_2234,In_2490);
nand U6140 (N_6140,In_1473,In_1743);
or U6141 (N_6141,In_763,In_618);
and U6142 (N_6142,In_583,In_1146);
or U6143 (N_6143,In_818,In_2068);
and U6144 (N_6144,In_1947,In_756);
nor U6145 (N_6145,In_2150,In_2174);
and U6146 (N_6146,In_775,In_2199);
nor U6147 (N_6147,In_2121,In_1284);
nor U6148 (N_6148,In_36,In_527);
nor U6149 (N_6149,In_946,In_2206);
nor U6150 (N_6150,In_513,In_999);
and U6151 (N_6151,In_2438,In_1249);
and U6152 (N_6152,In_2257,In_2044);
or U6153 (N_6153,In_1410,In_1760);
xor U6154 (N_6154,In_2489,In_144);
nor U6155 (N_6155,In_1900,In_530);
and U6156 (N_6156,In_601,In_1199);
nand U6157 (N_6157,In_563,In_414);
or U6158 (N_6158,In_683,In_1031);
and U6159 (N_6159,In_1338,In_153);
nor U6160 (N_6160,In_1823,In_0);
nand U6161 (N_6161,In_821,In_1383);
nor U6162 (N_6162,In_1755,In_966);
xor U6163 (N_6163,In_430,In_2298);
xor U6164 (N_6164,In_1121,In_2175);
or U6165 (N_6165,In_1113,In_39);
nor U6166 (N_6166,In_885,In_296);
nand U6167 (N_6167,In_848,In_1105);
nor U6168 (N_6168,In_1248,In_717);
nor U6169 (N_6169,In_2055,In_1419);
xnor U6170 (N_6170,In_1548,In_2025);
or U6171 (N_6171,In_1954,In_1012);
and U6172 (N_6172,In_162,In_407);
and U6173 (N_6173,In_1850,In_2266);
or U6174 (N_6174,In_1492,In_966);
and U6175 (N_6175,In_1004,In_1677);
nand U6176 (N_6176,In_1449,In_9);
nand U6177 (N_6177,In_1819,In_387);
nand U6178 (N_6178,In_1723,In_1991);
nand U6179 (N_6179,In_1780,In_525);
nor U6180 (N_6180,In_426,In_1591);
or U6181 (N_6181,In_1519,In_27);
nor U6182 (N_6182,In_815,In_1198);
nor U6183 (N_6183,In_1435,In_141);
nor U6184 (N_6184,In_987,In_2246);
nor U6185 (N_6185,In_2159,In_1142);
or U6186 (N_6186,In_2243,In_442);
nand U6187 (N_6187,In_438,In_513);
nor U6188 (N_6188,In_1578,In_1304);
and U6189 (N_6189,In_766,In_271);
nand U6190 (N_6190,In_2305,In_2006);
nor U6191 (N_6191,In_1827,In_1392);
and U6192 (N_6192,In_917,In_2377);
or U6193 (N_6193,In_954,In_874);
or U6194 (N_6194,In_823,In_1130);
nor U6195 (N_6195,In_1848,In_2490);
xor U6196 (N_6196,In_967,In_861);
or U6197 (N_6197,In_527,In_331);
or U6198 (N_6198,In_1741,In_1159);
or U6199 (N_6199,In_1992,In_1916);
and U6200 (N_6200,In_1282,In_1288);
nor U6201 (N_6201,In_2027,In_2084);
or U6202 (N_6202,In_1434,In_2474);
nand U6203 (N_6203,In_286,In_1780);
nor U6204 (N_6204,In_1359,In_912);
nand U6205 (N_6205,In_2422,In_225);
and U6206 (N_6206,In_404,In_951);
nand U6207 (N_6207,In_436,In_706);
or U6208 (N_6208,In_1880,In_1905);
nand U6209 (N_6209,In_2024,In_459);
nor U6210 (N_6210,In_1092,In_416);
xnor U6211 (N_6211,In_795,In_200);
nand U6212 (N_6212,In_247,In_178);
xnor U6213 (N_6213,In_1317,In_1531);
or U6214 (N_6214,In_1826,In_1719);
nand U6215 (N_6215,In_1052,In_657);
or U6216 (N_6216,In_356,In_1532);
nand U6217 (N_6217,In_855,In_1504);
nor U6218 (N_6218,In_1434,In_641);
or U6219 (N_6219,In_2242,In_900);
or U6220 (N_6220,In_779,In_2244);
nand U6221 (N_6221,In_66,In_1792);
or U6222 (N_6222,In_1179,In_366);
or U6223 (N_6223,In_1046,In_1597);
and U6224 (N_6224,In_875,In_510);
nand U6225 (N_6225,In_2146,In_2194);
nand U6226 (N_6226,In_1798,In_317);
nand U6227 (N_6227,In_1292,In_2308);
and U6228 (N_6228,In_741,In_1619);
and U6229 (N_6229,In_2146,In_1086);
and U6230 (N_6230,In_2379,In_147);
or U6231 (N_6231,In_1006,In_1547);
nor U6232 (N_6232,In_691,In_1366);
or U6233 (N_6233,In_2300,In_225);
or U6234 (N_6234,In_586,In_1070);
nor U6235 (N_6235,In_2312,In_242);
nand U6236 (N_6236,In_1090,In_869);
or U6237 (N_6237,In_2027,In_2220);
and U6238 (N_6238,In_1568,In_97);
nor U6239 (N_6239,In_1320,In_893);
nand U6240 (N_6240,In_416,In_2190);
and U6241 (N_6241,In_100,In_1047);
or U6242 (N_6242,In_2390,In_2281);
nor U6243 (N_6243,In_38,In_1441);
or U6244 (N_6244,In_1587,In_237);
nor U6245 (N_6245,In_1810,In_1259);
xnor U6246 (N_6246,In_1389,In_2483);
and U6247 (N_6247,In_314,In_1382);
nand U6248 (N_6248,In_803,In_109);
nand U6249 (N_6249,In_765,In_1700);
nor U6250 (N_6250,N_1551,N_349);
nor U6251 (N_6251,N_1991,N_6078);
or U6252 (N_6252,N_3602,N_5576);
and U6253 (N_6253,N_3004,N_3507);
or U6254 (N_6254,N_4767,N_5348);
or U6255 (N_6255,N_5251,N_1772);
or U6256 (N_6256,N_21,N_2750);
nand U6257 (N_6257,N_633,N_918);
or U6258 (N_6258,N_4776,N_1065);
nand U6259 (N_6259,N_1862,N_4489);
nor U6260 (N_6260,N_4898,N_3784);
nand U6261 (N_6261,N_269,N_2556);
nand U6262 (N_6262,N_2678,N_835);
or U6263 (N_6263,N_5708,N_4473);
nand U6264 (N_6264,N_3181,N_4354);
nand U6265 (N_6265,N_1774,N_3814);
nor U6266 (N_6266,N_2316,N_4239);
or U6267 (N_6267,N_1653,N_782);
nand U6268 (N_6268,N_2421,N_3709);
nor U6269 (N_6269,N_5009,N_1880);
xor U6270 (N_6270,N_4412,N_4843);
or U6271 (N_6271,N_91,N_1342);
and U6272 (N_6272,N_4927,N_39);
and U6273 (N_6273,N_1596,N_26);
nor U6274 (N_6274,N_2109,N_1975);
nor U6275 (N_6275,N_6167,N_5916);
and U6276 (N_6276,N_4557,N_3262);
nand U6277 (N_6277,N_2136,N_2143);
nor U6278 (N_6278,N_4752,N_6107);
and U6279 (N_6279,N_1703,N_4755);
xnor U6280 (N_6280,N_728,N_3137);
or U6281 (N_6281,N_5652,N_3831);
and U6282 (N_6282,N_2955,N_2732);
nor U6283 (N_6283,N_4186,N_5815);
or U6284 (N_6284,N_3572,N_4913);
nor U6285 (N_6285,N_2008,N_5804);
or U6286 (N_6286,N_1013,N_1256);
nand U6287 (N_6287,N_669,N_5854);
nor U6288 (N_6288,N_2058,N_4789);
and U6289 (N_6289,N_5012,N_5803);
nand U6290 (N_6290,N_3926,N_5199);
nand U6291 (N_6291,N_5465,N_2402);
nor U6292 (N_6292,N_2961,N_994);
xnor U6293 (N_6293,N_376,N_4464);
or U6294 (N_6294,N_857,N_997);
or U6295 (N_6295,N_1001,N_4121);
xnor U6296 (N_6296,N_5182,N_1313);
or U6297 (N_6297,N_5520,N_1961);
nand U6298 (N_6298,N_625,N_3558);
nor U6299 (N_6299,N_1810,N_822);
nand U6300 (N_6300,N_69,N_4096);
and U6301 (N_6301,N_2128,N_1701);
nor U6302 (N_6302,N_3578,N_5136);
or U6303 (N_6303,N_5851,N_3542);
and U6304 (N_6304,N_4891,N_495);
and U6305 (N_6305,N_843,N_893);
nor U6306 (N_6306,N_605,N_1489);
xnor U6307 (N_6307,N_972,N_525);
nand U6308 (N_6308,N_6025,N_304);
nor U6309 (N_6309,N_4504,N_1400);
nor U6310 (N_6310,N_823,N_4350);
nand U6311 (N_6311,N_1927,N_2204);
nor U6312 (N_6312,N_5402,N_4108);
xnor U6313 (N_6313,N_1276,N_4911);
nand U6314 (N_6314,N_510,N_5558);
and U6315 (N_6315,N_3892,N_3626);
nor U6316 (N_6316,N_384,N_4631);
nor U6317 (N_6317,N_865,N_6171);
nand U6318 (N_6318,N_4285,N_1467);
or U6319 (N_6319,N_4523,N_938);
nand U6320 (N_6320,N_3163,N_852);
nor U6321 (N_6321,N_1988,N_4830);
nand U6322 (N_6322,N_2981,N_1082);
or U6323 (N_6323,N_4932,N_5322);
nand U6324 (N_6324,N_4785,N_4779);
nor U6325 (N_6325,N_223,N_3806);
nand U6326 (N_6326,N_2183,N_4971);
and U6327 (N_6327,N_3436,N_3951);
nor U6328 (N_6328,N_2394,N_2775);
nand U6329 (N_6329,N_330,N_3655);
nor U6330 (N_6330,N_2671,N_3724);
nor U6331 (N_6331,N_3884,N_5670);
and U6332 (N_6332,N_5481,N_806);
xor U6333 (N_6333,N_1511,N_1817);
nand U6334 (N_6334,N_1732,N_3071);
nor U6335 (N_6335,N_1149,N_1014);
nor U6336 (N_6336,N_2879,N_887);
and U6337 (N_6337,N_1830,N_2539);
nand U6338 (N_6338,N_4696,N_2674);
and U6339 (N_6339,N_3915,N_2299);
or U6340 (N_6340,N_1788,N_780);
nand U6341 (N_6341,N_1214,N_1197);
nor U6342 (N_6342,N_2505,N_5113);
nand U6343 (N_6343,N_5840,N_1818);
nand U6344 (N_6344,N_3595,N_5478);
nor U6345 (N_6345,N_472,N_4520);
xor U6346 (N_6346,N_2697,N_4878);
or U6347 (N_6347,N_5073,N_1283);
or U6348 (N_6348,N_2059,N_597);
nor U6349 (N_6349,N_18,N_3868);
nor U6350 (N_6350,N_1016,N_5215);
or U6351 (N_6351,N_5446,N_5862);
nand U6352 (N_6352,N_3383,N_1393);
nand U6353 (N_6353,N_2564,N_3410);
and U6354 (N_6354,N_3415,N_2384);
nand U6355 (N_6355,N_42,N_4259);
or U6356 (N_6356,N_3032,N_2174);
and U6357 (N_6357,N_3451,N_1883);
or U6358 (N_6358,N_5109,N_4431);
nor U6359 (N_6359,N_3699,N_3962);
nor U6360 (N_6360,N_1017,N_3250);
and U6361 (N_6361,N_2822,N_621);
nand U6362 (N_6362,N_2129,N_619);
nor U6363 (N_6363,N_3473,N_5989);
nor U6364 (N_6364,N_4801,N_3466);
nor U6365 (N_6365,N_4562,N_1757);
or U6366 (N_6366,N_1325,N_4495);
and U6367 (N_6367,N_3036,N_3793);
nand U6368 (N_6368,N_638,N_6066);
and U6369 (N_6369,N_5150,N_6026);
nand U6370 (N_6370,N_5984,N_5356);
and U6371 (N_6371,N_5819,N_3117);
and U6372 (N_6372,N_4022,N_4331);
xnor U6373 (N_6373,N_3885,N_3371);
nand U6374 (N_6374,N_5195,N_3061);
nor U6375 (N_6375,N_6208,N_575);
xnor U6376 (N_6376,N_1643,N_413);
and U6377 (N_6377,N_3051,N_880);
nand U6378 (N_6378,N_3388,N_2507);
xor U6379 (N_6379,N_4769,N_2097);
and U6380 (N_6380,N_3337,N_2841);
nand U6381 (N_6381,N_1078,N_5865);
nand U6382 (N_6382,N_2454,N_2483);
and U6383 (N_6383,N_1417,N_2293);
or U6384 (N_6384,N_3168,N_5323);
xnor U6385 (N_6385,N_5740,N_5618);
and U6386 (N_6386,N_2550,N_5406);
nor U6387 (N_6387,N_4221,N_3936);
or U6388 (N_6388,N_2498,N_3299);
and U6389 (N_6389,N_4372,N_2622);
nand U6390 (N_6390,N_5718,N_5650);
or U6391 (N_6391,N_58,N_1168);
nor U6392 (N_6392,N_352,N_2116);
or U6393 (N_6393,N_3971,N_4536);
nor U6394 (N_6394,N_5660,N_2340);
nand U6395 (N_6395,N_1076,N_2496);
nand U6396 (N_6396,N_5237,N_1952);
nor U6397 (N_6397,N_1327,N_2971);
nand U6398 (N_6398,N_1754,N_5257);
nor U6399 (N_6399,N_2709,N_3556);
and U6400 (N_6400,N_4440,N_4027);
and U6401 (N_6401,N_3281,N_1372);
and U6402 (N_6402,N_6005,N_524);
and U6403 (N_6403,N_1437,N_4867);
nor U6404 (N_6404,N_2921,N_2253);
and U6405 (N_6405,N_3209,N_238);
nand U6406 (N_6406,N_423,N_3767);
and U6407 (N_6407,N_3654,N_2032);
and U6408 (N_6408,N_1411,N_533);
xor U6409 (N_6409,N_315,N_5357);
or U6410 (N_6410,N_916,N_5358);
xnor U6411 (N_6411,N_2292,N_4255);
nand U6412 (N_6412,N_2309,N_5492);
xnor U6413 (N_6413,N_3552,N_3332);
or U6414 (N_6414,N_5959,N_1849);
nand U6415 (N_6415,N_5169,N_3992);
nor U6416 (N_6416,N_1318,N_3873);
xnor U6417 (N_6417,N_2267,N_4863);
or U6418 (N_6418,N_1440,N_4584);
or U6419 (N_6419,N_4685,N_729);
nor U6420 (N_6420,N_2144,N_3840);
nand U6421 (N_6421,N_3576,N_4647);
and U6422 (N_6422,N_4589,N_4370);
and U6423 (N_6423,N_145,N_785);
xnor U6424 (N_6424,N_3227,N_5080);
xor U6425 (N_6425,N_3681,N_1780);
nor U6426 (N_6426,N_1403,N_5196);
or U6427 (N_6427,N_4569,N_382);
or U6428 (N_6428,N_2517,N_1783);
xor U6429 (N_6429,N_4157,N_32);
and U6430 (N_6430,N_3630,N_2432);
and U6431 (N_6431,N_4147,N_5645);
and U6432 (N_6432,N_694,N_2853);
nor U6433 (N_6433,N_159,N_2937);
or U6434 (N_6434,N_1941,N_2462);
xor U6435 (N_6435,N_1904,N_607);
or U6436 (N_6436,N_1264,N_153);
nor U6437 (N_6437,N_5760,N_4364);
or U6438 (N_6438,N_1282,N_5394);
or U6439 (N_6439,N_6145,N_6214);
and U6440 (N_6440,N_6010,N_5936);
and U6441 (N_6441,N_2552,N_2005);
or U6442 (N_6442,N_1965,N_3592);
nor U6443 (N_6443,N_415,N_5850);
or U6444 (N_6444,N_883,N_5780);
nand U6445 (N_6445,N_82,N_190);
and U6446 (N_6446,N_836,N_5370);
or U6447 (N_6447,N_1535,N_3217);
nand U6448 (N_6448,N_5793,N_1233);
and U6449 (N_6449,N_6109,N_3346);
and U6450 (N_6450,N_5194,N_6084);
nor U6451 (N_6451,N_5747,N_2371);
or U6452 (N_6452,N_2904,N_5299);
xnor U6453 (N_6453,N_2436,N_5482);
and U6454 (N_6454,N_4109,N_2348);
or U6455 (N_6455,N_2696,N_2272);
or U6456 (N_6456,N_3961,N_5430);
nand U6457 (N_6457,N_3698,N_4635);
nor U6458 (N_6458,N_5509,N_4312);
xor U6459 (N_6459,N_1486,N_83);
and U6460 (N_6460,N_1390,N_6162);
nand U6461 (N_6461,N_4173,N_3820);
and U6462 (N_6462,N_1695,N_2854);
nor U6463 (N_6463,N_1879,N_684);
and U6464 (N_6464,N_4057,N_344);
and U6465 (N_6465,N_6118,N_5824);
or U6466 (N_6466,N_3588,N_1636);
nand U6467 (N_6467,N_2731,N_1442);
nor U6468 (N_6468,N_1228,N_3018);
nand U6469 (N_6469,N_2185,N_1742);
xor U6470 (N_6470,N_4053,N_3746);
and U6471 (N_6471,N_2708,N_3092);
or U6472 (N_6472,N_5990,N_1932);
and U6473 (N_6473,N_6058,N_3494);
nand U6474 (N_6474,N_278,N_6095);
and U6475 (N_6475,N_2780,N_3252);
nand U6476 (N_6476,N_0,N_1550);
and U6477 (N_6477,N_648,N_3932);
or U6478 (N_6478,N_1131,N_3967);
nand U6479 (N_6479,N_3710,N_5894);
and U6480 (N_6480,N_568,N_3505);
nand U6481 (N_6481,N_2273,N_3854);
nand U6482 (N_6482,N_4050,N_794);
nand U6483 (N_6483,N_580,N_1051);
nor U6484 (N_6484,N_2627,N_2077);
nand U6485 (N_6485,N_2905,N_3104);
nand U6486 (N_6486,N_3502,N_1169);
nor U6487 (N_6487,N_2343,N_4196);
and U6488 (N_6488,N_201,N_1007);
xnor U6489 (N_6489,N_1552,N_4585);
nand U6490 (N_6490,N_4895,N_4518);
nor U6491 (N_6491,N_5971,N_1431);
and U6492 (N_6492,N_1706,N_2249);
or U6493 (N_6493,N_559,N_4949);
xor U6494 (N_6494,N_1516,N_2798);
or U6495 (N_6495,N_1566,N_2886);
or U6496 (N_6496,N_6038,N_4226);
or U6497 (N_6497,N_287,N_3070);
or U6498 (N_6498,N_1728,N_1262);
nor U6499 (N_6499,N_5565,N_3562);
xor U6500 (N_6500,N_1979,N_5425);
xnor U6501 (N_6501,N_2598,N_2495);
nor U6502 (N_6502,N_3839,N_5519);
and U6503 (N_6503,N_2719,N_1167);
xor U6504 (N_6504,N_252,N_2061);
nand U6505 (N_6505,N_36,N_1165);
nand U6506 (N_6506,N_6238,N_4244);
nor U6507 (N_6507,N_4385,N_1092);
xor U6508 (N_6508,N_10,N_2982);
nand U6509 (N_6509,N_1998,N_3886);
and U6510 (N_6510,N_4883,N_3215);
and U6511 (N_6511,N_4737,N_4343);
nor U6512 (N_6512,N_5786,N_692);
nand U6513 (N_6513,N_4527,N_3644);
or U6514 (N_6514,N_5381,N_140);
nand U6515 (N_6515,N_3666,N_2653);
nor U6516 (N_6516,N_810,N_4903);
nand U6517 (N_6517,N_2198,N_4279);
nor U6518 (N_6518,N_355,N_3234);
xnor U6519 (N_6519,N_4939,N_4339);
and U6520 (N_6520,N_2132,N_564);
and U6521 (N_6521,N_2624,N_889);
nor U6522 (N_6522,N_3786,N_1586);
nand U6523 (N_6523,N_3596,N_5434);
nor U6524 (N_6524,N_5426,N_4115);
nand U6525 (N_6525,N_5068,N_954);
or U6526 (N_6526,N_1814,N_5676);
and U6527 (N_6527,N_2339,N_2861);
xor U6528 (N_6528,N_5077,N_645);
or U6529 (N_6529,N_3665,N_2929);
and U6530 (N_6530,N_4969,N_3445);
nor U6531 (N_6531,N_763,N_672);
xor U6532 (N_6532,N_2560,N_1617);
or U6533 (N_6533,N_264,N_1791);
nor U6534 (N_6534,N_4695,N_5452);
nor U6535 (N_6535,N_1377,N_901);
nor U6536 (N_6536,N_5996,N_1920);
and U6537 (N_6537,N_5141,N_3583);
or U6538 (N_6538,N_5023,N_5928);
nand U6539 (N_6539,N_2933,N_5052);
nor U6540 (N_6540,N_1631,N_3910);
nand U6541 (N_6541,N_233,N_3310);
and U6542 (N_6542,N_4291,N_5217);
or U6543 (N_6543,N_1000,N_1958);
nand U6544 (N_6544,N_2226,N_1216);
or U6545 (N_6545,N_1490,N_113);
nand U6546 (N_6546,N_129,N_4297);
nand U6547 (N_6547,N_5705,N_793);
and U6548 (N_6548,N_3449,N_5884);
or U6549 (N_6549,N_4497,N_2930);
or U6550 (N_6550,N_1996,N_4533);
and U6551 (N_6551,N_1127,N_5255);
xnor U6552 (N_6552,N_4321,N_3409);
nor U6553 (N_6553,N_5311,N_760);
nand U6554 (N_6554,N_986,N_929);
nand U6555 (N_6555,N_3862,N_6157);
and U6556 (N_6556,N_3469,N_2197);
nand U6557 (N_6557,N_1488,N_5308);
nor U6558 (N_6558,N_6142,N_2802);
or U6559 (N_6559,N_3619,N_1844);
nand U6560 (N_6560,N_3925,N_1937);
nand U6561 (N_6561,N_3351,N_281);
and U6562 (N_6562,N_3264,N_4966);
and U6563 (N_6563,N_1948,N_3513);
and U6564 (N_6564,N_2170,N_3703);
and U6565 (N_6565,N_5893,N_3541);
nor U6566 (N_6566,N_1751,N_2338);
or U6567 (N_6567,N_501,N_5516);
nor U6568 (N_6568,N_774,N_2881);
and U6569 (N_6569,N_4019,N_570);
xnor U6570 (N_6570,N_4942,N_4828);
nor U6571 (N_6571,N_802,N_683);
nor U6572 (N_6572,N_5028,N_1546);
nor U6573 (N_6573,N_1093,N_1603);
or U6574 (N_6574,N_3269,N_1825);
or U6575 (N_6575,N_995,N_5991);
xnor U6576 (N_6576,N_4806,N_1089);
nand U6577 (N_6577,N_5778,N_4723);
nand U6578 (N_6578,N_4783,N_4796);
and U6579 (N_6579,N_491,N_1856);
or U6580 (N_6580,N_4835,N_1660);
and U6581 (N_6581,N_1005,N_6144);
or U6582 (N_6582,N_2034,N_2230);
and U6583 (N_6583,N_4131,N_1936);
and U6584 (N_6584,N_1408,N_1401);
and U6585 (N_6585,N_879,N_1881);
xor U6586 (N_6586,N_1555,N_4603);
nand U6587 (N_6587,N_5571,N_3);
and U6588 (N_6588,N_3816,N_2374);
and U6589 (N_6589,N_6130,N_5048);
nand U6590 (N_6590,N_1659,N_1497);
xnor U6591 (N_6591,N_4149,N_237);
and U6592 (N_6592,N_5721,N_17);
xnor U6593 (N_6593,N_5629,N_2289);
nand U6594 (N_6594,N_1134,N_5297);
nor U6595 (N_6595,N_4705,N_195);
nor U6596 (N_6596,N_6081,N_3567);
xor U6597 (N_6597,N_327,N_1741);
xor U6598 (N_6598,N_4420,N_4066);
or U6599 (N_6599,N_674,N_3606);
and U6600 (N_6600,N_1985,N_3470);
or U6601 (N_6601,N_5334,N_5798);
and U6602 (N_6602,N_766,N_5677);
or U6603 (N_6603,N_6076,N_5902);
nor U6604 (N_6604,N_2831,N_1986);
nor U6605 (N_6605,N_5970,N_3246);
and U6606 (N_6606,N_3255,N_5530);
or U6607 (N_6607,N_3969,N_5045);
xnor U6608 (N_6608,N_3518,N_6114);
nand U6609 (N_6609,N_4181,N_40);
nand U6610 (N_6610,N_795,N_1439);
nand U6611 (N_6611,N_4896,N_1355);
and U6612 (N_6612,N_2363,N_4020);
nand U6613 (N_6613,N_1840,N_3173);
nor U6614 (N_6614,N_5941,N_5062);
nand U6615 (N_6615,N_3008,N_1358);
and U6616 (N_6616,N_3352,N_2050);
nor U6617 (N_6617,N_3189,N_2745);
and U6618 (N_6618,N_4645,N_3210);
nor U6619 (N_6619,N_4390,N_624);
or U6620 (N_6620,N_4706,N_4588);
nor U6621 (N_6621,N_2012,N_411);
nand U6622 (N_6622,N_5281,N_1529);
and U6623 (N_6623,N_4854,N_3199);
or U6624 (N_6624,N_900,N_2416);
or U6625 (N_6625,N_3922,N_710);
and U6626 (N_6626,N_2200,N_3062);
xor U6627 (N_6627,N_357,N_4310);
xor U6628 (N_6628,N_1652,N_4151);
and U6629 (N_6629,N_2238,N_5019);
nor U6630 (N_6630,N_5918,N_1733);
xor U6631 (N_6631,N_3731,N_1745);
and U6632 (N_6632,N_4357,N_557);
nand U6633 (N_6633,N_2789,N_3373);
xor U6634 (N_6634,N_1392,N_1462);
nand U6635 (N_6635,N_5646,N_3824);
nand U6636 (N_6636,N_1435,N_1521);
xnor U6637 (N_6637,N_417,N_5716);
and U6638 (N_6638,N_2234,N_2779);
xnor U6639 (N_6639,N_530,N_5992);
nand U6640 (N_6640,N_3005,N_1931);
and U6641 (N_6641,N_5157,N_5692);
and U6642 (N_6642,N_461,N_276);
nand U6643 (N_6643,N_5352,N_2614);
nor U6644 (N_6644,N_1646,N_1252);
nor U6645 (N_6645,N_2544,N_2536);
xnor U6646 (N_6646,N_4424,N_4494);
and U6647 (N_6647,N_2332,N_5829);
nand U6648 (N_6648,N_3280,N_4940);
nor U6649 (N_6649,N_926,N_574);
and U6650 (N_6650,N_362,N_2127);
xnor U6651 (N_6651,N_6064,N_6224);
nor U6652 (N_6652,N_2395,N_4491);
and U6653 (N_6653,N_5764,N_2855);
or U6654 (N_6654,N_3114,N_2212);
or U6655 (N_6655,N_2563,N_5181);
nor U6656 (N_6656,N_3879,N_5120);
and U6657 (N_6657,N_4185,N_5514);
or U6658 (N_6658,N_778,N_4237);
nor U6659 (N_6659,N_2767,N_2549);
or U6660 (N_6660,N_5277,N_3870);
nand U6661 (N_6661,N_1678,N_5060);
nor U6662 (N_6662,N_5282,N_2533);
or U6663 (N_6663,N_3601,N_1487);
and U6664 (N_6664,N_671,N_1257);
or U6665 (N_6665,N_1020,N_3535);
nor U6666 (N_6666,N_4791,N_4383);
and U6667 (N_6667,N_2915,N_92);
or U6668 (N_6668,N_1345,N_1281);
nor U6669 (N_6669,N_732,N_2187);
nand U6670 (N_6670,N_892,N_6027);
nand U6671 (N_6671,N_3621,N_4272);
and U6672 (N_6672,N_3286,N_2070);
and U6673 (N_6673,N_482,N_2874);
or U6674 (N_6674,N_5147,N_3830);
or U6675 (N_6675,N_5805,N_905);
nor U6676 (N_6676,N_3256,N_4967);
nand U6677 (N_6677,N_2687,N_2192);
and U6678 (N_6678,N_3590,N_3347);
nand U6679 (N_6679,N_5171,N_2442);
or U6680 (N_6680,N_1402,N_4248);
xor U6681 (N_6681,N_3164,N_6001);
nand U6682 (N_6682,N_5673,N_4251);
nor U6683 (N_6683,N_5545,N_2172);
nor U6684 (N_6684,N_1104,N_3198);
and U6685 (N_6685,N_2972,N_2345);
nor U6686 (N_6686,N_401,N_1476);
or U6687 (N_6687,N_2047,N_2443);
nand U6688 (N_6688,N_3491,N_4238);
or U6689 (N_6689,N_1297,N_3381);
xor U6690 (N_6690,N_2582,N_2110);
and U6691 (N_6691,N_1997,N_392);
xor U6692 (N_6692,N_4751,N_2571);
nor U6693 (N_6693,N_5144,N_661);
and U6694 (N_6694,N_3127,N_4764);
or U6695 (N_6695,N_2445,N_4514);
or U6696 (N_6696,N_5763,N_649);
nor U6697 (N_6697,N_4199,N_5130);
or U6698 (N_6698,N_4119,N_6055);
nand U6699 (N_6699,N_639,N_2898);
nand U6700 (N_6700,N_3006,N_4069);
nand U6701 (N_6701,N_6217,N_1177);
xor U6702 (N_6702,N_1781,N_4701);
or U6703 (N_6703,N_5695,N_725);
and U6704 (N_6704,N_1222,N_2561);
nor U6705 (N_6705,N_945,N_2328);
nor U6706 (N_6706,N_3894,N_1038);
nand U6707 (N_6707,N_1136,N_1563);
and U6708 (N_6708,N_3203,N_318);
nand U6709 (N_6709,N_1887,N_4104);
nor U6710 (N_6710,N_4299,N_2297);
nand U6711 (N_6711,N_6175,N_3627);
nor U6712 (N_6712,N_731,N_5159);
and U6713 (N_6713,N_2527,N_3150);
nor U6714 (N_6714,N_4732,N_95);
nand U6715 (N_6715,N_1949,N_741);
nand U6716 (N_6716,N_6222,N_5539);
or U6717 (N_6717,N_4450,N_1559);
and U6718 (N_6718,N_4811,N_2907);
xor U6719 (N_6719,N_1908,N_5375);
nand U6720 (N_6720,N_828,N_745);
xor U6721 (N_6721,N_1650,N_5952);
or U6722 (N_6722,N_2852,N_4389);
nand U6723 (N_6723,N_4521,N_1715);
or U6724 (N_6724,N_5898,N_1620);
nor U6725 (N_6725,N_1983,N_4375);
or U6726 (N_6726,N_2283,N_4807);
xor U6727 (N_6727,N_3774,N_5455);
nand U6728 (N_6728,N_679,N_1923);
or U6729 (N_6729,N_5106,N_3033);
xor U6730 (N_6730,N_182,N_2487);
nor U6731 (N_6731,N_4072,N_5822);
and U6732 (N_6732,N_3722,N_4264);
nand U6733 (N_6733,N_636,N_2811);
nor U6734 (N_6734,N_3160,N_4613);
nor U6735 (N_6735,N_5653,N_4713);
and U6736 (N_6736,N_2209,N_6151);
nand U6737 (N_6737,N_1698,N_3003);
xnor U6738 (N_6738,N_5387,N_4148);
and U6739 (N_6739,N_5785,N_691);
nand U6740 (N_6740,N_6148,N_312);
and U6741 (N_6741,N_777,N_2526);
and U6742 (N_6742,N_5428,N_4710);
and U6743 (N_6743,N_3539,N_5599);
nand U6744 (N_6744,N_5267,N_1303);
and U6745 (N_6745,N_488,N_5588);
nand U6746 (N_6746,N_5209,N_4163);
nor U6747 (N_6747,N_248,N_2287);
nor U6748 (N_6748,N_5066,N_961);
nor U6749 (N_6749,N_4682,N_5184);
nand U6750 (N_6750,N_4156,N_5668);
nor U6751 (N_6751,N_743,N_2011);
and U6752 (N_6752,N_2511,N_1096);
nor U6753 (N_6753,N_4326,N_4033);
or U6754 (N_6754,N_4268,N_759);
nor U6755 (N_6755,N_4062,N_2094);
or U6756 (N_6756,N_3480,N_4866);
nand U6757 (N_6757,N_2838,N_3843);
nand U6758 (N_6758,N_2346,N_3524);
nand U6759 (N_6759,N_2638,N_6242);
nor U6760 (N_6760,N_4483,N_2959);
nor U6761 (N_6761,N_5046,N_2589);
or U6762 (N_6762,N_3653,N_3861);
or U6763 (N_6763,N_1637,N_1049);
xnor U6764 (N_6764,N_1441,N_2817);
nor U6765 (N_6765,N_924,N_4654);
and U6766 (N_6766,N_5466,N_361);
xor U6767 (N_6767,N_1919,N_6097);
nand U6768 (N_6768,N_4439,N_2479);
nand U6769 (N_6769,N_440,N_164);
or U6770 (N_6770,N_3849,N_4073);
and U6771 (N_6771,N_3434,N_4747);
xor U6772 (N_6772,N_4182,N_4614);
xnor U6773 (N_6773,N_2155,N_5056);
and U6774 (N_6774,N_6124,N_2474);
xor U6775 (N_6775,N_3421,N_4488);
xor U6776 (N_6776,N_3794,N_2036);
and U6777 (N_6777,N_6169,N_2823);
nand U6778 (N_6778,N_1538,N_5974);
nand U6779 (N_6779,N_2579,N_3852);
and U6780 (N_6780,N_1023,N_2023);
or U6781 (N_6781,N_753,N_1835);
xor U6782 (N_6782,N_465,N_730);
and U6783 (N_6783,N_1394,N_5934);
nand U6784 (N_6784,N_6057,N_270);
nor U6785 (N_6785,N_460,N_1851);
or U6786 (N_6786,N_4017,N_3579);
nor U6787 (N_6787,N_138,N_4006);
nand U6788 (N_6788,N_663,N_1615);
nor U6789 (N_6789,N_99,N_259);
nor U6790 (N_6790,N_5950,N_4427);
nand U6791 (N_6791,N_4954,N_5140);
nand U6792 (N_6792,N_1523,N_1011);
nand U6793 (N_6793,N_418,N_3860);
nor U6794 (N_6794,N_4270,N_4646);
and U6795 (N_6795,N_3404,N_554);
nand U6796 (N_6796,N_4659,N_5315);
xnor U6797 (N_6797,N_5269,N_2606);
and U6798 (N_6798,N_5367,N_2509);
nor U6799 (N_6799,N_1806,N_3461);
or U6800 (N_6800,N_660,N_4496);
and U6801 (N_6801,N_3772,N_78);
nand U6802 (N_6802,N_320,N_1054);
or U6803 (N_6803,N_2265,N_2104);
nand U6804 (N_6804,N_2264,N_5727);
nand U6805 (N_6805,N_943,N_2501);
and U6806 (N_6806,N_737,N_210);
or U6807 (N_6807,N_5689,N_1707);
nor U6808 (N_6808,N_5467,N_6204);
nand U6809 (N_6809,N_86,N_5138);
and U6810 (N_6810,N_1376,N_1500);
and U6811 (N_6811,N_3367,N_3113);
or U6812 (N_6812,N_5532,N_5883);
nand U6813 (N_6813,N_1700,N_3933);
or U6814 (N_6814,N_3705,N_1590);
and U6815 (N_6815,N_6015,N_5293);
and U6816 (N_6816,N_5647,N_1713);
and U6817 (N_6817,N_5948,N_2894);
nand U6818 (N_6818,N_2938,N_4016);
nor U6819 (N_6819,N_4855,N_4735);
xor U6820 (N_6820,N_2518,N_1704);
xor U6821 (N_6821,N_4555,N_3713);
or U6822 (N_6822,N_4824,N_3349);
nor U6823 (N_6823,N_5988,N_3475);
and U6824 (N_6824,N_1589,N_2530);
and U6825 (N_6825,N_3391,N_3847);
nand U6826 (N_6826,N_1503,N_714);
or U6827 (N_6827,N_2041,N_5095);
nor U6828 (N_6828,N_2591,N_2269);
xnor U6829 (N_6829,N_6031,N_5276);
nor U6830 (N_6830,N_126,N_3612);
nor U6831 (N_6831,N_2396,N_2827);
nor U6832 (N_6832,N_4143,N_3154);
nand U6833 (N_6833,N_3110,N_2661);
or U6834 (N_6834,N_6131,N_93);
or U6835 (N_6835,N_2239,N_4928);
and U6836 (N_6836,N_3275,N_1352);
nand U6837 (N_6837,N_1326,N_6065);
nand U6838 (N_6838,N_5180,N_3344);
nand U6839 (N_6839,N_2149,N_4348);
and U6840 (N_6840,N_4917,N_5291);
xor U6841 (N_6841,N_1581,N_2409);
or U6842 (N_6842,N_5038,N_4401);
and U6843 (N_6843,N_4524,N_428);
xnor U6844 (N_6844,N_2373,N_5960);
and U6845 (N_6845,N_2635,N_3838);
and U6846 (N_6846,N_354,N_2068);
nand U6847 (N_6847,N_5875,N_4686);
or U6848 (N_6848,N_2969,N_1061);
or U6849 (N_6849,N_1577,N_5307);
or U6850 (N_6850,N_6189,N_5207);
nor U6851 (N_6851,N_5575,N_3093);
nor U6852 (N_6852,N_3440,N_1247);
or U6853 (N_6853,N_288,N_4859);
or U6854 (N_6854,N_3272,N_2873);
and U6855 (N_6855,N_5316,N_6194);
nor U6856 (N_6856,N_3533,N_5253);
and U6857 (N_6857,N_592,N_5642);
and U6858 (N_6858,N_4295,N_2319);
xnor U6859 (N_6859,N_5577,N_3244);
nor U6860 (N_6860,N_4026,N_3799);
nor U6861 (N_6861,N_2913,N_3687);
xnor U6862 (N_6862,N_1719,N_863);
nand U6863 (N_6863,N_5266,N_1219);
and U6864 (N_6864,N_1644,N_5256);
or U6865 (N_6865,N_869,N_2926);
nor U6866 (N_6866,N_5407,N_5298);
nand U6867 (N_6867,N_257,N_3991);
nor U6868 (N_6868,N_5067,N_68);
nor U6869 (N_6869,N_317,N_6244);
or U6870 (N_6870,N_5491,N_516);
nand U6871 (N_6871,N_5445,N_3225);
and U6872 (N_6872,N_682,N_3363);
and U6873 (N_6873,N_4535,N_1542);
nor U6874 (N_6874,N_73,N_5582);
or U6875 (N_6875,N_1506,N_131);
and U6876 (N_6876,N_5039,N_1890);
and U6877 (N_6877,N_3105,N_2461);
nor U6878 (N_6878,N_5354,N_4211);
nand U6879 (N_6879,N_830,N_2457);
and U6880 (N_6880,N_6176,N_5675);
nor U6881 (N_6881,N_4402,N_4229);
nor U6882 (N_6882,N_2203,N_435);
or U6883 (N_6883,N_3046,N_4529);
nand U6884 (N_6884,N_4388,N_249);
nand U6885 (N_6885,N_4697,N_2689);
nor U6886 (N_6886,N_1456,N_4651);
and U6887 (N_6887,N_5871,N_3909);
and U6888 (N_6888,N_55,N_4296);
or U6889 (N_6889,N_3075,N_247);
nand U6890 (N_6890,N_4384,N_3455);
or U6891 (N_6891,N_2691,N_1351);
nor U6892 (N_6892,N_553,N_3216);
nor U6893 (N_6893,N_5137,N_2562);
xnor U6894 (N_6894,N_115,N_5353);
nand U6895 (N_6895,N_1540,N_3733);
and U6896 (N_6896,N_5286,N_1080);
nand U6897 (N_6897,N_3519,N_2753);
and U6898 (N_6898,N_2872,N_4231);
nor U6899 (N_6899,N_2379,N_1962);
and U6900 (N_6900,N_1347,N_2295);
and U6901 (N_6901,N_3285,N_1073);
and U6902 (N_6902,N_2458,N_5878);
or U6903 (N_6903,N_333,N_2931);
or U6904 (N_6904,N_202,N_5769);
or U6905 (N_6905,N_4922,N_1598);
nand U6906 (N_6906,N_623,N_127);
nand U6907 (N_6907,N_4582,N_1519);
xor U6908 (N_6908,N_4198,N_2399);
nand U6909 (N_6909,N_1120,N_1004);
nand U6910 (N_6910,N_2086,N_1805);
xnor U6911 (N_6911,N_6161,N_1277);
or U6912 (N_6912,N_420,N_4052);
xor U6913 (N_6913,N_2331,N_2728);
or U6914 (N_6914,N_4698,N_4203);
nand U6915 (N_6915,N_3378,N_2232);
nand U6916 (N_6916,N_1196,N_2868);
nand U6917 (N_6917,N_2105,N_5337);
or U6918 (N_6918,N_4294,N_5024);
nor U6919 (N_6919,N_4957,N_2590);
or U6920 (N_6920,N_6234,N_859);
and U6921 (N_6921,N_3921,N_4308);
nor U6922 (N_6922,N_2803,N_3248);
and U6923 (N_6923,N_1808,N_1340);
nor U6924 (N_6924,N_4616,N_3901);
nor U6925 (N_6925,N_3624,N_3593);
and U6926 (N_6926,N_175,N_4177);
nor U6927 (N_6927,N_5944,N_1397);
nand U6928 (N_6928,N_5810,N_4498);
and U6929 (N_6929,N_2049,N_3708);
or U6930 (N_6930,N_4038,N_4775);
nand U6931 (N_6931,N_3952,N_2729);
or U6932 (N_6932,N_5399,N_3509);
or U6933 (N_6933,N_1882,N_1547);
and U6934 (N_6934,N_1656,N_323);
nand U6935 (N_6935,N_3400,N_5006);
and U6936 (N_6936,N_3982,N_4950);
or U6937 (N_6937,N_5235,N_87);
or U6938 (N_6938,N_4162,N_1614);
xor U6939 (N_6939,N_5003,N_4897);
nand U6940 (N_6940,N_837,N_3484);
or U6941 (N_6941,N_2506,N_5754);
or U6942 (N_6942,N_2075,N_1162);
nand U6943 (N_6943,N_647,N_548);
xnor U6944 (N_6944,N_1539,N_5688);
nand U6945 (N_6945,N_950,N_5386);
nor U6946 (N_6946,N_3336,N_5818);
or U6947 (N_6947,N_1716,N_457);
or U6948 (N_6948,N_3429,N_5349);
nor U6949 (N_6949,N_3717,N_4002);
nor U6950 (N_6950,N_3645,N_3757);
nand U6951 (N_6951,N_1874,N_345);
nand U6952 (N_6952,N_6000,N_983);
xor U6953 (N_6953,N_2057,N_4323);
nand U6954 (N_6954,N_2390,N_303);
and U6955 (N_6955,N_3029,N_4741);
nand U6956 (N_6956,N_626,N_2456);
nor U6957 (N_6957,N_4825,N_1175);
nor U6958 (N_6958,N_1062,N_4861);
or U6959 (N_6959,N_6212,N_1570);
xnor U6960 (N_6960,N_3883,N_1939);
or U6961 (N_6961,N_6125,N_1155);
and U6962 (N_6962,N_5190,N_2377);
xnor U6963 (N_6963,N_5143,N_4102);
and U6964 (N_6964,N_2106,N_168);
and U6965 (N_6965,N_1957,N_5566);
nor U6966 (N_6966,N_4085,N_4505);
or U6967 (N_6967,N_1787,N_3819);
nand U6968 (N_6968,N_1258,N_2983);
or U6969 (N_6969,N_262,N_3017);
xor U6970 (N_6970,N_4900,N_3265);
and U6971 (N_6971,N_235,N_2889);
xor U6972 (N_6972,N_4722,N_596);
or U6973 (N_6973,N_1170,N_4228);
or U6974 (N_6974,N_12,N_4795);
nor U6975 (N_6975,N_3453,N_5125);
nor U6976 (N_6976,N_6052,N_2246);
and U6977 (N_6977,N_5411,N_4470);
nor U6978 (N_6978,N_1959,N_680);
nor U6979 (N_6979,N_6190,N_4309);
or U6980 (N_6980,N_97,N_915);
nand U6981 (N_6981,N_4515,N_4709);
xor U6982 (N_6982,N_1621,N_752);
xor U6983 (N_6983,N_5540,N_2541);
or U6984 (N_6984,N_3002,N_5817);
or U6985 (N_6985,N_541,N_1221);
or U6986 (N_6986,N_4623,N_1595);
or U6987 (N_6987,N_100,N_2037);
or U6988 (N_6988,N_4544,N_2422);
nand U6989 (N_6989,N_1148,N_5597);
or U6990 (N_6990,N_54,N_2568);
or U6991 (N_6991,N_5206,N_5391);
xnor U6992 (N_6992,N_5926,N_1749);
or U6993 (N_6993,N_2387,N_1622);
and U6994 (N_6994,N_6226,N_4443);
xnor U6995 (N_6995,N_5270,N_1925);
nor U6996 (N_6996,N_5518,N_2213);
or U6997 (N_6997,N_5112,N_1205);
xor U6998 (N_6998,N_5163,N_2644);
nand U6999 (N_6999,N_5226,N_125);
or U7000 (N_7000,N_3740,N_3917);
or U7001 (N_7001,N_1336,N_3928);
nand U7002 (N_7002,N_5681,N_5026);
and U7003 (N_7003,N_3000,N_2698);
nand U7004 (N_7004,N_5230,N_203);
nor U7005 (N_7005,N_1574,N_5999);
or U7006 (N_7006,N_3721,N_6112);
or U7007 (N_7007,N_1048,N_157);
or U7008 (N_7008,N_3537,N_3431);
and U7009 (N_7009,N_4414,N_4008);
and U7010 (N_7010,N_946,N_2813);
xor U7011 (N_7011,N_3563,N_2375);
xnor U7012 (N_7012,N_4453,N_5320);
and U7013 (N_7013,N_5957,N_3028);
or U7014 (N_7014,N_641,N_5938);
nor U7015 (N_7015,N_3437,N_3550);
and U7016 (N_7016,N_5110,N_1203);
and U7017 (N_7017,N_6074,N_4522);
or U7018 (N_7018,N_5027,N_4035);
and U7019 (N_7019,N_412,N_690);
xnor U7020 (N_7020,N_3907,N_1672);
nand U7021 (N_7021,N_2654,N_1980);
nor U7022 (N_7022,N_2277,N_6173);
or U7023 (N_7023,N_4049,N_4127);
nor U7024 (N_7024,N_3144,N_4381);
nor U7025 (N_7025,N_2686,N_337);
nand U7026 (N_7026,N_424,N_5528);
and U7027 (N_7027,N_1746,N_2233);
nor U7028 (N_7028,N_3320,N_5703);
and U7029 (N_7029,N_984,N_6117);
nor U7030 (N_7030,N_6013,N_1915);
xnor U7031 (N_7031,N_4658,N_2943);
or U7032 (N_7032,N_1099,N_5409);
nor U7033 (N_7033,N_2778,N_1311);
nand U7034 (N_7034,N_4142,N_6136);
nor U7035 (N_7035,N_3439,N_2166);
or U7036 (N_7036,N_2617,N_2000);
and U7037 (N_7037,N_2329,N_980);
or U7038 (N_7038,N_2173,N_4858);
or U7039 (N_7039,N_2188,N_2123);
and U7040 (N_7040,N_4080,N_1188);
nor U7041 (N_7041,N_5336,N_2065);
or U7042 (N_7042,N_4225,N_3338);
xnor U7043 (N_7043,N_6049,N_4091);
nor U7044 (N_7044,N_3095,N_3447);
or U7045 (N_7045,N_4851,N_3357);
nand U7046 (N_7046,N_2863,N_1926);
nor U7047 (N_7047,N_1235,N_4892);
nand U7048 (N_7048,N_4074,N_5254);
nor U7049 (N_7049,N_60,N_5870);
or U7050 (N_7050,N_1195,N_769);
nor U7051 (N_7051,N_1532,N_3063);
or U7052 (N_7052,N_5392,N_3997);
or U7053 (N_7053,N_3300,N_4597);
nor U7054 (N_7054,N_2593,N_1767);
nor U7055 (N_7055,N_1184,N_2521);
or U7056 (N_7056,N_151,N_5521);
or U7057 (N_7057,N_1869,N_3171);
nand U7058 (N_7058,N_3727,N_5920);
nor U7059 (N_7059,N_3782,N_919);
and U7060 (N_7060,N_913,N_4935);
nand U7061 (N_7061,N_1338,N_3779);
and U7062 (N_7062,N_1995,N_5847);
nand U7063 (N_7063,N_458,N_2);
or U7064 (N_7064,N_3249,N_104);
nor U7065 (N_7065,N_1480,N_2946);
nor U7066 (N_7066,N_2901,N_5013);
xor U7067 (N_7067,N_1457,N_1674);
nand U7068 (N_7068,N_4134,N_5698);
and U7069 (N_7069,N_2219,N_5639);
nor U7070 (N_7070,N_2532,N_979);
or U7071 (N_7071,N_2290,N_2397);
and U7072 (N_7072,N_566,N_3841);
nor U7073 (N_7073,N_1265,N_4210);
nor U7074 (N_7074,N_5700,N_5636);
nor U7075 (N_7075,N_3825,N_2870);
or U7076 (N_7076,N_2196,N_3972);
nor U7077 (N_7077,N_2081,N_1418);
nand U7078 (N_7078,N_2288,N_1034);
nor U7079 (N_7079,N_4926,N_5369);
and U7080 (N_7080,N_414,N_119);
or U7081 (N_7081,N_5473,N_5343);
or U7082 (N_7082,N_4220,N_5324);
and U7083 (N_7083,N_4876,N_4610);
nor U7084 (N_7084,N_4673,N_2824);
or U7085 (N_7085,N_3023,N_2680);
and U7086 (N_7086,N_431,N_4592);
nor U7087 (N_7087,N_5170,N_5423);
xor U7088 (N_7088,N_5090,N_477);
or U7089 (N_7089,N_4469,N_4123);
or U7090 (N_7090,N_5418,N_1892);
nor U7091 (N_7091,N_2694,N_5283);
nor U7092 (N_7092,N_4906,N_1116);
nand U7093 (N_7093,N_571,N_1290);
or U7094 (N_7094,N_5994,N_3193);
and U7095 (N_7095,N_4733,N_1396);
nand U7096 (N_7096,N_5302,N_229);
xnor U7097 (N_7097,N_4993,N_637);
or U7098 (N_7098,N_6152,N_230);
nor U7099 (N_7099,N_432,N_1968);
nor U7100 (N_7100,N_266,N_2554);
nor U7101 (N_7101,N_2141,N_722);
and U7102 (N_7102,N_2919,N_5551);
nor U7103 (N_7103,N_3530,N_5672);
nand U7104 (N_7104,N_816,N_775);
xor U7105 (N_7105,N_498,N_2191);
and U7106 (N_7106,N_6028,N_137);
or U7107 (N_7107,N_3121,N_989);
nand U7108 (N_7108,N_4833,N_4813);
nor U7109 (N_7109,N_3790,N_707);
nand U7110 (N_7110,N_2333,N_1661);
or U7111 (N_7111,N_5963,N_2455);
and U7112 (N_7112,N_4781,N_4168);
or U7113 (N_7113,N_6102,N_282);
nand U7114 (N_7114,N_3517,N_572);
nand U7115 (N_7115,N_192,N_4905);
and U7116 (N_7116,N_5342,N_5836);
nor U7117 (N_7117,N_4333,N_3610);
nand U7118 (N_7118,N_456,N_3343);
xnor U7119 (N_7119,N_4273,N_220);
xnor U7120 (N_7120,N_5917,N_4650);
nor U7121 (N_7121,N_736,N_5549);
xnor U7122 (N_7122,N_5156,N_3066);
or U7123 (N_7123,N_2307,N_6037);
and U7124 (N_7124,N_110,N_1907);
or U7125 (N_7125,N_2986,N_4169);
nor U7126 (N_7126,N_4772,N_656);
or U7127 (N_7127,N_5659,N_1686);
or U7128 (N_7128,N_3034,N_346);
or U7129 (N_7129,N_2475,N_3506);
nand U7130 (N_7130,N_1019,N_4758);
or U7131 (N_7131,N_5462,N_1642);
or U7132 (N_7132,N_4322,N_4023);
nand U7133 (N_7133,N_4111,N_5861);
nand U7134 (N_7134,N_851,N_3257);
nand U7135 (N_7135,N_213,N_2256);
and U7136 (N_7136,N_3496,N_4672);
or U7137 (N_7137,N_5289,N_5054);
or U7138 (N_7138,N_2014,N_6087);
or U7139 (N_7139,N_2089,N_437);
or U7140 (N_7140,N_2365,N_2692);
and U7141 (N_7141,N_4532,N_3015);
and U7142 (N_7142,N_5723,N_5542);
nand U7143 (N_7143,N_5503,N_5555);
and U7144 (N_7144,N_6165,N_4171);
and U7145 (N_7145,N_2079,N_5525);
or U7146 (N_7146,N_4531,N_3204);
and U7147 (N_7147,N_3515,N_342);
nand U7148 (N_7148,N_2965,N_962);
nand U7149 (N_7149,N_4593,N_4959);
or U7150 (N_7150,N_3560,N_2088);
nand U7151 (N_7151,N_388,N_5347);
nand U7152 (N_7152,N_2076,N_4078);
xnor U7153 (N_7153,N_3649,N_4044);
or U7154 (N_7154,N_2490,N_6237);
nand U7155 (N_7155,N_3048,N_2320);
nor U7156 (N_7156,N_3525,N_1232);
or U7157 (N_7157,N_3098,N_6108);
and U7158 (N_7158,N_963,N_1353);
nand U7159 (N_7159,N_6195,N_6128);
nand U7160 (N_7160,N_923,N_4301);
nand U7161 (N_7161,N_1484,N_5091);
and U7162 (N_7162,N_4548,N_4990);
or U7163 (N_7163,N_1368,N_2266);
or U7164 (N_7164,N_3042,N_4360);
nor U7165 (N_7165,N_6202,N_4214);
or U7166 (N_7166,N_2783,N_1124);
nor U7167 (N_7167,N_4844,N_4135);
nor U7168 (N_7168,N_1709,N_4680);
nand U7169 (N_7169,N_3212,N_850);
nor U7170 (N_7170,N_1399,N_2038);
nor U7171 (N_7171,N_3990,N_1930);
xor U7172 (N_7172,N_3865,N_4573);
or U7173 (N_7173,N_5203,N_4355);
or U7174 (N_7174,N_5097,N_4164);
and U7175 (N_7175,N_466,N_5906);
xnor U7176 (N_7176,N_3620,N_2378);
nor U7177 (N_7177,N_4952,N_2962);
xnor U7178 (N_7178,N_1850,N_2703);
or U7179 (N_7179,N_4693,N_1610);
and U7180 (N_7180,N_610,N_232);
nor U7181 (N_7181,N_2715,N_5732);
and U7182 (N_7182,N_1956,N_1180);
or U7183 (N_7183,N_2566,N_1922);
nand U7184 (N_7184,N_2497,N_2484);
or U7185 (N_7185,N_1496,N_1421);
and U7186 (N_7186,N_5876,N_3223);
or U7187 (N_7187,N_1198,N_5373);
and U7188 (N_7188,N_1126,N_5745);
nor U7189 (N_7189,N_1872,N_1670);
nand U7190 (N_7190,N_5098,N_3100);
xnor U7191 (N_7191,N_2326,N_4934);
nand U7192 (N_7192,N_4748,N_4176);
nor U7193 (N_7193,N_5863,N_5295);
and U7194 (N_7194,N_193,N_1429);
nor U7195 (N_7195,N_4873,N_3608);
nand U7196 (N_7196,N_2013,N_3011);
nor U7197 (N_7197,N_2812,N_4794);
nor U7198 (N_7198,N_1135,N_3402);
nand U7199 (N_7199,N_1365,N_302);
and U7200 (N_7200,N_80,N_6082);
nor U7201 (N_7201,N_3911,N_1052);
nand U7202 (N_7202,N_5317,N_5366);
and U7203 (N_7203,N_2762,N_2084);
xnor U7204 (N_7204,N_178,N_3211);
xor U7205 (N_7205,N_4512,N_3850);
nand U7206 (N_7206,N_4258,N_170);
nand U7207 (N_7207,N_681,N_5301);
nand U7208 (N_7208,N_3801,N_176);
or U7209 (N_7209,N_3107,N_627);
and U7210 (N_7210,N_1863,N_6196);
or U7211 (N_7211,N_4609,N_1482);
and U7212 (N_7212,N_5410,N_1183);
or U7213 (N_7213,N_761,N_5845);
or U7214 (N_7214,N_5278,N_3827);
nor U7215 (N_7215,N_2382,N_2987);
nand U7216 (N_7216,N_2547,N_4992);
nor U7217 (N_7217,N_4644,N_1208);
or U7218 (N_7218,N_2922,N_4549);
nor U7219 (N_7219,N_5447,N_3859);
nand U7220 (N_7220,N_4487,N_1604);
and U7221 (N_7221,N_2437,N_3983);
or U7222 (N_7222,N_3206,N_4058);
or U7223 (N_7223,N_4043,N_244);
or U7224 (N_7224,N_4731,N_5690);
nand U7225 (N_7225,N_6178,N_1223);
nor U7226 (N_7226,N_1527,N_5498);
nand U7227 (N_7227,N_3872,N_1725);
nor U7228 (N_7228,N_4460,N_6135);
and U7229 (N_7229,N_2313,N_528);
and U7230 (N_7230,N_4530,N_3463);
and U7231 (N_7231,N_4466,N_4133);
xnor U7232 (N_7232,N_1602,N_4690);
xor U7233 (N_7233,N_4916,N_3313);
xnor U7234 (N_7234,N_2755,N_3876);
xor U7235 (N_7235,N_3845,N_4325);
and U7236 (N_7236,N_2883,N_96);
nand U7237 (N_7237,N_377,N_5531);
nor U7238 (N_7238,N_2467,N_4558);
nor U7239 (N_7239,N_243,N_3780);
or U7240 (N_7240,N_5726,N_2893);
or U7241 (N_7241,N_2156,N_2949);
and U7242 (N_7242,N_265,N_4541);
and U7243 (N_7243,N_3573,N_2353);
or U7244 (N_7244,N_57,N_1302);
nor U7245 (N_7245,N_4869,N_311);
or U7246 (N_7246,N_5420,N_4831);
and U7247 (N_7247,N_3053,N_3021);
or U7248 (N_7248,N_5376,N_1894);
nor U7249 (N_7249,N_3435,N_6174);
and U7250 (N_7250,N_289,N_2605);
or U7251 (N_7251,N_4191,N_4284);
nand U7252 (N_7252,N_4422,N_3500);
nor U7253 (N_7253,N_2660,N_3968);
or U7254 (N_7254,N_942,N_5587);
nor U7255 (N_7255,N_698,N_4987);
nor U7256 (N_7256,N_4893,N_5100);
nand U7257 (N_7257,N_1009,N_1823);
nand U7258 (N_7258,N_2389,N_517);
nor U7259 (N_7259,N_5072,N_4629);
or U7260 (N_7260,N_5176,N_3664);
or U7261 (N_7261,N_1337,N_3220);
xor U7262 (N_7262,N_5064,N_3340);
xor U7263 (N_7263,N_1225,N_1119);
xor U7264 (N_7264,N_4947,N_5133);
xor U7265 (N_7265,N_1274,N_4738);
nor U7266 (N_7266,N_1978,N_3935);
and U7267 (N_7267,N_2357,N_2391);
nand U7268 (N_7268,N_3303,N_2601);
nand U7269 (N_7269,N_3635,N_5431);
nor U7270 (N_7270,N_3896,N_5413);
xor U7271 (N_7271,N_2882,N_2616);
nand U7272 (N_7272,N_4790,N_4387);
nor U7273 (N_7273,N_3676,N_579);
or U7274 (N_7274,N_3716,N_4970);
nand U7275 (N_7275,N_1152,N_167);
nand U7276 (N_7276,N_2695,N_2748);
or U7277 (N_7277,N_6139,N_5332);
nand U7278 (N_7278,N_3682,N_263);
nand U7279 (N_7279,N_105,N_5359);
nand U7280 (N_7280,N_5485,N_1974);
nor U7281 (N_7281,N_5812,N_1572);
and U7282 (N_7282,N_1455,N_3981);
nand U7283 (N_7283,N_1504,N_419);
and U7284 (N_7284,N_292,N_2832);
nand U7285 (N_7285,N_2386,N_497);
nand U7286 (N_7286,N_4884,N_1813);
nor U7287 (N_7287,N_5686,N_427);
nand U7288 (N_7288,N_3770,N_2347);
nor U7289 (N_7289,N_4009,N_1891);
xor U7290 (N_7290,N_1640,N_1021);
nor U7291 (N_7291,N_5192,N_2216);
and U7292 (N_7292,N_2608,N_4218);
or U7293 (N_7293,N_4944,N_5568);
or U7294 (N_7294,N_5678,N_250);
and U7295 (N_7295,N_3116,N_338);
nor U7296 (N_7296,N_3293,N_827);
nor U7297 (N_7297,N_283,N_968);
or U7298 (N_7298,N_5535,N_4688);
nor U7299 (N_7299,N_5435,N_2424);
nor U7300 (N_7300,N_3035,N_3696);
nand U7301 (N_7301,N_4490,N_481);
nor U7302 (N_7302,N_3902,N_2718);
nand U7303 (N_7303,N_3955,N_800);
nand U7304 (N_7304,N_336,N_5742);
nor U7305 (N_7305,N_4652,N_2491);
nor U7306 (N_7306,N_3775,N_3025);
nor U7307 (N_7307,N_5579,N_6103);
and U7308 (N_7308,N_4253,N_439);
and U7309 (N_7309,N_2741,N_5259);
or U7310 (N_7310,N_150,N_4792);
nor U7311 (N_7311,N_949,N_2951);
nor U7312 (N_7312,N_332,N_4337);
nor U7313 (N_7313,N_3147,N_272);
and U7314 (N_7314,N_4580,N_3218);
xor U7315 (N_7315,N_152,N_5318);
or U7316 (N_7316,N_408,N_5512);
or U7317 (N_7317,N_5129,N_1057);
nor U7318 (N_7318,N_4263,N_499);
nor U7319 (N_7319,N_4061,N_4809);
and U7320 (N_7320,N_976,N_331);
nand U7321 (N_7321,N_5787,N_454);
or U7322 (N_7322,N_1031,N_1301);
nand U7323 (N_7323,N_6111,N_2469);
nor U7324 (N_7324,N_5612,N_5004);
nand U7325 (N_7325,N_4419,N_5616);
or U7326 (N_7326,N_165,N_3259);
nand U7327 (N_7327,N_3412,N_2364);
nand U7328 (N_7328,N_360,N_2800);
nand U7329 (N_7329,N_3106,N_5372);
or U7330 (N_7330,N_2208,N_545);
and U7331 (N_7331,N_1270,N_4586);
nand U7332 (N_7332,N_6068,N_5351);
or U7333 (N_7333,N_744,N_1328);
nor U7334 (N_7334,N_4564,N_5111);
and U7335 (N_7335,N_1371,N_4662);
nand U7336 (N_7336,N_5264,N_63);
or U7337 (N_7337,N_3514,N_951);
and U7338 (N_7338,N_1449,N_3980);
nor U7339 (N_7339,N_2025,N_2594);
nand U7340 (N_7340,N_3504,N_2083);
and U7341 (N_7341,N_3638,N_1471);
or U7342 (N_7342,N_5595,N_4671);
and U7343 (N_7343,N_5560,N_5477);
and U7344 (N_7344,N_2744,N_2186);
nand U7345 (N_7345,N_3625,N_6070);
nand U7346 (N_7346,N_3656,N_6093);
nand U7347 (N_7347,N_6180,N_1284);
xnor U7348 (N_7348,N_4444,N_5522);
nor U7349 (N_7349,N_4034,N_3763);
and U7350 (N_7350,N_5033,N_3836);
nor U7351 (N_7351,N_3050,N_2906);
nor U7352 (N_7352,N_2917,N_1778);
or U7353 (N_7353,N_1554,N_5327);
nor U7354 (N_7354,N_772,N_5075);
nor U7355 (N_7355,N_494,N_5596);
nor U7356 (N_7356,N_5648,N_4172);
nor U7357 (N_7357,N_3416,N_4342);
nand U7358 (N_7358,N_4894,N_4649);
nor U7359 (N_7359,N_1638,N_3386);
and U7360 (N_7360,N_1464,N_3325);
nor U7361 (N_7361,N_1608,N_2860);
and U7362 (N_7362,N_395,N_5005);
or U7363 (N_7363,N_783,N_5749);
nor U7364 (N_7364,N_3543,N_5788);
and U7365 (N_7365,N_5201,N_5213);
and U7366 (N_7366,N_3027,N_3342);
or U7367 (N_7367,N_5869,N_3283);
nand U7368 (N_7368,N_3773,N_5644);
or U7369 (N_7369,N_4194,N_4438);
and U7370 (N_7370,N_5161,N_2837);
and U7371 (N_7371,N_3575,N_831);
nor U7372 (N_7372,N_4392,N_4624);
nor U7373 (N_7373,N_5222,N_3988);
or U7374 (N_7374,N_1111,N_5151);
nor U7375 (N_7375,N_2615,N_2147);
or U7376 (N_7376,N_4261,N_5490);
nor U7377 (N_7377,N_2607,N_1724);
and U7378 (N_7378,N_4417,N_3887);
nor U7379 (N_7379,N_3778,N_3375);
nor U7380 (N_7380,N_5931,N_2829);
or U7381 (N_7381,N_4025,N_650);
or U7382 (N_7382,N_6248,N_1687);
or U7383 (N_7383,N_5903,N_2761);
nor U7384 (N_7384,N_6241,N_2636);
nand U7385 (N_7385,N_3690,N_1889);
or U7386 (N_7386,N_2022,N_4070);
nor U7387 (N_7387,N_3175,N_3930);
or U7388 (N_7388,N_207,N_4568);
nand U7389 (N_7389,N_3766,N_3319);
and U7390 (N_7390,N_5043,N_98);
nor U7391 (N_7391,N_6182,N_5309);
nand U7392 (N_7392,N_3807,N_4200);
nor U7393 (N_7393,N_4865,N_3747);
nor U7394 (N_7394,N_4425,N_4418);
and U7395 (N_7395,N_5244,N_5249);
or U7396 (N_7396,N_4675,N_1509);
xnor U7397 (N_7397,N_3752,N_1220);
xnor U7398 (N_7398,N_529,N_1557);
and U7399 (N_7399,N_5114,N_5280);
and U7400 (N_7400,N_3672,N_4094);
nor U7401 (N_7401,N_5746,N_2225);
nand U7402 (N_7402,N_4224,N_143);
nand U7403 (N_7403,N_2522,N_6170);
or U7404 (N_7404,N_550,N_5495);
or U7405 (N_7405,N_4076,N_2111);
nor U7406 (N_7406,N_3693,N_4985);
and U7407 (N_7407,N_5055,N_1865);
or U7408 (N_7408,N_1896,N_3049);
and U7409 (N_7409,N_2626,N_3056);
nand U7410 (N_7410,N_2899,N_6150);
or U7411 (N_7411,N_2046,N_4754);
nor U7412 (N_7412,N_4933,N_2760);
and U7413 (N_7413,N_3660,N_2415);
nand U7414 (N_7414,N_3570,N_4930);
nand U7415 (N_7415,N_5940,N_6030);
xnor U7416 (N_7416,N_2030,N_1341);
nor U7417 (N_7417,N_1321,N_4441);
nand U7418 (N_7418,N_8,N_3667);
xor U7419 (N_7419,N_808,N_1726);
nand U7420 (N_7420,N_4914,N_3657);
or U7421 (N_7421,N_2095,N_3454);
nand U7422 (N_7422,N_70,N_3874);
nand U7423 (N_7423,N_6223,N_3791);
and U7424 (N_7424,N_4909,N_3202);
and U7425 (N_7425,N_1575,N_4122);
and U7426 (N_7426,N_4327,N_4467);
or U7427 (N_7427,N_4391,N_6069);
or U7428 (N_7428,N_4872,N_5606);
and U7429 (N_7429,N_2612,N_4305);
nor U7430 (N_7430,N_1766,N_297);
and U7431 (N_7431,N_4823,N_35);
nor U7432 (N_7432,N_2069,N_1954);
nand U7433 (N_7433,N_4124,N_1782);
nor U7434 (N_7434,N_1307,N_2451);
nor U7435 (N_7435,N_2600,N_3615);
nand U7436 (N_7436,N_4510,N_2066);
and U7437 (N_7437,N_4189,N_85);
or U7438 (N_7438,N_425,N_6036);
nor U7439 (N_7439,N_4445,N_2181);
and U7440 (N_7440,N_4179,N_3704);
nor U7441 (N_7441,N_5442,N_1838);
or U7442 (N_7442,N_2236,N_2902);
nand U7443 (N_7443,N_936,N_3689);
or U7444 (N_7444,N_1826,N_4627);
nor U7445 (N_7445,N_1876,N_319);
or U7446 (N_7446,N_2119,N_2138);
nor U7447 (N_7447,N_4463,N_3039);
or U7448 (N_7448,N_4840,N_4081);
xnor U7449 (N_7449,N_1045,N_1619);
or U7450 (N_7450,N_5977,N_4410);
nor U7451 (N_7451,N_1250,N_988);
nor U7452 (N_7452,N_1130,N_652);
xor U7453 (N_7453,N_3762,N_6240);
or U7454 (N_7454,N_4641,N_1382);
or U7455 (N_7455,N_387,N_897);
or U7456 (N_7456,N_520,N_5500);
or U7457 (N_7457,N_5814,N_3149);
xnor U7458 (N_7458,N_1161,N_1349);
and U7459 (N_7459,N_4679,N_2646);
xnor U7460 (N_7460,N_5015,N_838);
or U7461 (N_7461,N_2362,N_447);
and U7462 (N_7462,N_3899,N_5059);
nor U7463 (N_7463,N_2411,N_4178);
or U7464 (N_7464,N_490,N_3986);
nor U7465 (N_7465,N_4800,N_3783);
and U7466 (N_7466,N_3711,N_1384);
nand U7467 (N_7467,N_2131,N_1971);
nand U7468 (N_7468,N_4014,N_3187);
nor U7469 (N_7469,N_1299,N_5801);
nor U7470 (N_7470,N_6053,N_911);
nand U7471 (N_7471,N_544,N_2538);
nand U7472 (N_7472,N_5084,N_3321);
or U7473 (N_7473,N_3714,N_1422);
nor U7474 (N_7474,N_101,N_1583);
nand U7475 (N_7475,N_6179,N_5210);
or U7476 (N_7476,N_906,N_4740);
xor U7477 (N_7477,N_1025,N_588);
or U7478 (N_7478,N_6188,N_2604);
and U7479 (N_7479,N_109,N_5937);
nand U7480 (N_7480,N_3586,N_2318);
and U7481 (N_7481,N_254,N_5915);
and U7482 (N_7482,N_1839,N_3547);
or U7483 (N_7483,N_5135,N_2018);
nand U7484 (N_7484,N_4605,N_3851);
nor U7485 (N_7485,N_5378,N_5837);
nor U7486 (N_7486,N_6012,N_2055);
or U7487 (N_7487,N_749,N_47);
nand U7488 (N_7488,N_2722,N_5242);
and U7489 (N_7489,N_1953,N_4963);
nand U7490 (N_7490,N_3331,N_4665);
nor U7491 (N_7491,N_1389,N_3728);
xor U7492 (N_7492,N_6003,N_2021);
xnor U7493 (N_7493,N_2426,N_1736);
or U7494 (N_7494,N_4306,N_2945);
or U7495 (N_7495,N_2214,N_2115);
xnor U7496 (N_7496,N_5325,N_532);
or U7497 (N_7497,N_4361,N_2581);
xor U7498 (N_7498,N_719,N_6183);
and U7499 (N_7499,N_1354,N_2251);
nor U7500 (N_7500,N_5607,N_534);
and U7501 (N_7501,N_5563,N_4461);
or U7502 (N_7502,N_4539,N_2966);
and U7503 (N_7503,N_5594,N_5720);
and U7504 (N_7504,N_2820,N_3397);
or U7505 (N_7505,N_4346,N_2355);
nand U7506 (N_7506,N_4042,N_3043);
or U7507 (N_7507,N_2263,N_4882);
nand U7508 (N_7508,N_3634,N_5864);
nor U7509 (N_7509,N_4994,N_4366);
xnor U7510 (N_7510,N_3818,N_5330);
or U7511 (N_7511,N_872,N_2989);
nand U7512 (N_7512,N_2334,N_6228);
and U7513 (N_7513,N_1914,N_3291);
nor U7514 (N_7514,N_3939,N_1520);
xor U7515 (N_7515,N_3764,N_2254);
and U7516 (N_7516,N_2400,N_521);
and U7517 (N_7517,N_2845,N_4480);
and U7518 (N_7518,N_3369,N_5655);
xnor U7519 (N_7519,N_668,N_155);
or U7520 (N_7520,N_5559,N_6083);
nor U7521 (N_7521,N_3497,N_4482);
nor U7522 (N_7522,N_1731,N_2932);
nor U7523 (N_7523,N_4379,N_3529);
nand U7524 (N_7524,N_4547,N_3566);
and U7525 (N_7525,N_4766,N_4829);
xor U7526 (N_7526,N_5188,N_6156);
xor U7527 (N_7527,N_2991,N_14);
or U7528 (N_7528,N_2525,N_5160);
nor U7529 (N_7529,N_4174,N_348);
or U7530 (N_7530,N_5995,N_3452);
nor U7531 (N_7531,N_1285,N_2040);
nand U7532 (N_7532,N_2224,N_1729);
xnor U7533 (N_7533,N_1317,N_3236);
nor U7534 (N_7534,N_3462,N_3605);
or U7535 (N_7535,N_6021,N_1344);
and U7536 (N_7536,N_3686,N_1386);
xnor U7537 (N_7537,N_2351,N_4462);
xor U7538 (N_7538,N_1679,N_5149);
nand U7539 (N_7539,N_1312,N_2618);
or U7540 (N_7540,N_2417,N_3755);
nand U7541 (N_7541,N_5076,N_3282);
nor U7542 (N_7542,N_5843,N_426);
and U7543 (N_7543,N_2118,N_1655);
and U7544 (N_7544,N_1730,N_2158);
nand U7545 (N_7545,N_1768,N_2184);
nor U7546 (N_7546,N_2393,N_3754);
xor U7547 (N_7547,N_5913,N_4637);
nor U7548 (N_7548,N_2996,N_4018);
nand U7549 (N_7549,N_3109,N_5168);
or U7550 (N_7550,N_1153,N_1436);
nor U7551 (N_7551,N_2404,N_1360);
xnor U7552 (N_7552,N_3551,N_5627);
nor U7553 (N_7553,N_2321,N_1015);
xor U7554 (N_7554,N_3308,N_5604);
nand U7555 (N_7555,N_2749,N_1357);
or U7556 (N_7556,N_5797,N_2805);
or U7557 (N_7557,N_3268,N_4150);
nand U7558 (N_7558,N_3243,N_2447);
and U7559 (N_7559,N_593,N_3184);
nand U7560 (N_7560,N_5643,N_1605);
nor U7561 (N_7561,N_2250,N_4919);
and U7562 (N_7562,N_5912,N_1804);
and U7563 (N_7563,N_1112,N_1626);
nor U7564 (N_7564,N_479,N_2435);
nor U7565 (N_7565,N_1584,N_878);
or U7566 (N_7566,N_2410,N_2053);
and U7567 (N_7567,N_2367,N_1860);
and U7568 (N_7568,N_313,N_1409);
and U7569 (N_7569,N_1982,N_5384);
nor U7570 (N_7570,N_3701,N_3010);
or U7571 (N_7571,N_4661,N_2508);
and U7572 (N_7572,N_3129,N_5074);
and U7573 (N_7573,N_4976,N_2880);
nand U7574 (N_7574,N_2135,N_884);
xnor U7575 (N_7575,N_4028,N_5557);
or U7576 (N_7576,N_540,N_925);
xor U7577 (N_7577,N_3001,N_4979);
or U7578 (N_7578,N_5935,N_1479);
and U7579 (N_7579,N_912,N_3213);
nand U7580 (N_7580,N_4978,N_4269);
nor U7581 (N_7581,N_434,N_81);
and U7582 (N_7582,N_350,N_4479);
or U7583 (N_7583,N_2052,N_396);
nor U7584 (N_7584,N_1964,N_4352);
nor U7585 (N_7585,N_712,N_5866);
or U7586 (N_7586,N_5008,N_4736);
nor U7587 (N_7587,N_5609,N_5685);
or U7588 (N_7588,N_3094,N_5953);
nor U7589 (N_7589,N_1366,N_4694);
or U7590 (N_7590,N_1334,N_2542);
nand U7591 (N_7591,N_3743,N_3133);
nor U7592 (N_7592,N_4743,N_5250);
nor U7593 (N_7593,N_5214,N_2342);
nor U7594 (N_7594,N_3897,N_4975);
xnor U7595 (N_7595,N_3208,N_3700);
or U7596 (N_7596,N_4745,N_5032);
or U7597 (N_7597,N_4526,N_4707);
nand U7598 (N_7598,N_1824,N_576);
and U7599 (N_7599,N_5833,N_3196);
or U7600 (N_7600,N_1702,N_3185);
nor U7601 (N_7601,N_4165,N_3594);
or U7602 (N_7602,N_5637,N_5547);
or U7603 (N_7603,N_5641,N_3393);
nor U7604 (N_7604,N_537,N_1800);
nand U7605 (N_7605,N_1305,N_1545);
nand U7606 (N_7606,N_4880,N_2452);
xnor U7607 (N_7607,N_3372,N_2954);
and U7608 (N_7608,N_5578,N_5887);
or U7609 (N_7609,N_4625,N_5621);
xor U7610 (N_7610,N_2903,N_5424);
xor U7611 (N_7611,N_3718,N_4572);
xor U7612 (N_7612,N_5813,N_5826);
or U7613 (N_7613,N_1864,N_4670);
or U7614 (N_7614,N_1717,N_4099);
nor U7615 (N_7615,N_4761,N_3516);
or U7616 (N_7616,N_947,N_5220);
and U7617 (N_7617,N_2578,N_4506);
nor U7618 (N_7618,N_894,N_4429);
nor U7619 (N_7619,N_5807,N_2151);
or U7620 (N_7620,N_4029,N_4386);
or U7621 (N_7621,N_2350,N_2944);
nor U7622 (N_7622,N_6147,N_4634);
nand U7623 (N_7623,N_825,N_5233);
nand U7624 (N_7624,N_1102,N_4007);
or U7625 (N_7625,N_711,N_1573);
and U7626 (N_7626,N_6033,N_325);
xor U7627 (N_7627,N_4814,N_2707);
or U7628 (N_7628,N_5564,N_5633);
or U7629 (N_7629,N_2392,N_5748);
nand U7630 (N_7630,N_4106,N_5954);
nand U7631 (N_7631,N_5132,N_2828);
nor U7632 (N_7632,N_4565,N_128);
xor U7633 (N_7633,N_535,N_5622);
xnor U7634 (N_7634,N_4227,N_560);
nor U7635 (N_7635,N_3628,N_5770);
nor U7636 (N_7636,N_5212,N_149);
nor U7637 (N_7637,N_4786,N_2091);
and U7638 (N_7638,N_3833,N_1253);
or U7639 (N_7639,N_2891,N_4750);
nand U7640 (N_7640,N_3115,N_5187);
or U7641 (N_7641,N_274,N_4329);
nand U7642 (N_7642,N_1651,N_708);
nor U7643 (N_7643,N_3977,N_5759);
or U7644 (N_7644,N_3103,N_492);
and U7645 (N_7645,N_1292,N_2039);
or U7646 (N_7646,N_1524,N_3792);
nor U7647 (N_7647,N_1333,N_3574);
and U7648 (N_7648,N_364,N_6085);
or U7649 (N_7649,N_506,N_896);
and U7650 (N_7650,N_2975,N_2247);
and U7651 (N_7651,N_1171,N_3811);
nor U7652 (N_7652,N_5538,N_2711);
nor U7653 (N_7653,N_1259,N_6168);
or U7654 (N_7654,N_3954,N_5733);
nor U7655 (N_7655,N_5263,N_5225);
or U7656 (N_7656,N_4160,N_6210);
and U7657 (N_7657,N_1966,N_978);
and U7658 (N_7658,N_3538,N_2510);
xnor U7659 (N_7659,N_1871,N_1159);
xor U7660 (N_7660,N_2701,N_3065);
nor U7661 (N_7661,N_4241,N_1193);
xor U7662 (N_7662,N_3598,N_2520);
nor U7663 (N_7663,N_4797,N_2090);
and U7664 (N_7664,N_6126,N_515);
nor U7665 (N_7665,N_487,N_634);
or U7666 (N_7666,N_3633,N_3464);
nor U7667 (N_7667,N_3406,N_6132);
and U7668 (N_7668,N_6200,N_5923);
nand U7669 (N_7669,N_3798,N_3156);
or U7670 (N_7670,N_3408,N_6104);
nand U7671 (N_7671,N_79,N_1592);
or U7672 (N_7672,N_5762,N_6123);
nand U7673 (N_7673,N_4770,N_3471);
or U7674 (N_7674,N_2177,N_6035);
or U7675 (N_7675,N_2130,N_1665);
and U7676 (N_7676,N_227,N_4234);
nand U7677 (N_7677,N_4213,N_549);
xor U7678 (N_7678,N_2912,N_2317);
and U7679 (N_7679,N_3301,N_755);
nand U7680 (N_7680,N_5173,N_618);
xnor U7681 (N_7681,N_2667,N_5725);
nor U7682 (N_7682,N_234,N_180);
or U7683 (N_7683,N_3045,N_3546);
or U7684 (N_7684,N_1107,N_5486);
nor U7685 (N_7685,N_3324,N_5536);
or U7686 (N_7686,N_2489,N_5842);
or U7687 (N_7687,N_5603,N_1032);
nor U7688 (N_7688,N_1799,N_6245);
nor U7689 (N_7689,N_429,N_294);
and U7690 (N_7690,N_206,N_6177);
nor U7691 (N_7691,N_310,N_5153);
nand U7692 (N_7692,N_1943,N_365);
or U7693 (N_7693,N_3058,N_6143);
or U7694 (N_7694,N_1578,N_1556);
xnor U7695 (N_7695,N_5921,N_3245);
nor U7696 (N_7696,N_2559,N_1453);
xnor U7697 (N_7697,N_4345,N_5908);
nor U7698 (N_7698,N_3520,N_5234);
or U7699 (N_7699,N_4575,N_4827);
or U7700 (N_7700,N_2368,N_5667);
and U7701 (N_7701,N_5344,N_1348);
nand U7702 (N_7702,N_2551,N_3472);
nor U7703 (N_7703,N_5001,N_4656);
nand U7704 (N_7704,N_5782,N_1822);
and U7705 (N_7705,N_2020,N_2871);
nor U7706 (N_7706,N_197,N_3882);
nand U7707 (N_7707,N_1945,N_2716);
nand U7708 (N_7708,N_1845,N_3424);
and U7709 (N_7709,N_2009,N_2073);
or U7710 (N_7710,N_5827,N_5287);
nand U7711 (N_7711,N_727,N_4368);
nor U7712 (N_7712,N_4718,N_1514);
xnor U7713 (N_7713,N_3041,N_4404);
and U7714 (N_7714,N_343,N_4260);
nand U7715 (N_7715,N_1708,N_1694);
nand U7716 (N_7716,N_1027,N_1172);
nand U7717 (N_7717,N_1967,N_4508);
nor U7718 (N_7718,N_219,N_3456);
and U7719 (N_7719,N_88,N_2478);
nor U7720 (N_7720,N_1597,N_5041);
nand U7721 (N_7721,N_1363,N_839);
and U7722 (N_7722,N_2814,N_194);
nand U7723 (N_7723,N_2864,N_2739);
nor U7724 (N_7724,N_5846,N_4307);
or U7725 (N_7725,N_146,N_3976);
nor U7726 (N_7726,N_5791,N_1940);
or U7727 (N_7727,N_1633,N_2159);
and U7728 (N_7728,N_3354,N_3937);
nand U7729 (N_7729,N_3521,N_2503);
and U7730 (N_7730,N_4907,N_1491);
nand U7731 (N_7731,N_5661,N_6233);
nand U7732 (N_7732,N_5752,N_2586);
xor U7733 (N_7733,N_4778,N_695);
and U7734 (N_7734,N_2336,N_5590);
and U7735 (N_7735,N_1204,N_4287);
nor U7736 (N_7736,N_422,N_4400);
nor U7737 (N_7737,N_3364,N_622);
and U7738 (N_7738,N_2947,N_2107);
nand U7739 (N_7739,N_24,N_4476);
or U7740 (N_7740,N_3522,N_5197);
nand U7741 (N_7741,N_3642,N_3221);
nor U7742 (N_7742,N_4845,N_2344);
or U7743 (N_7743,N_33,N_1028);
nand U7744 (N_7744,N_363,N_5600);
nand U7745 (N_7745,N_3157,N_6225);
nor U7746 (N_7746,N_5385,N_4996);
or U7747 (N_7747,N_5709,N_3912);
nand U7748 (N_7748,N_2493,N_4982);
and U7749 (N_7749,N_2211,N_6024);
and U7750 (N_7750,N_3355,N_5104);
and U7751 (N_7751,N_1905,N_797);
or U7752 (N_7752,N_3253,N_4689);
or U7753 (N_7753,N_5929,N_2210);
and U7754 (N_7754,N_2352,N_4724);
nor U7755 (N_7755,N_2546,N_4358);
or U7756 (N_7756,N_5605,N_493);
and U7757 (N_7757,N_2015,N_251);
or U7758 (N_7758,N_2529,N_2408);
and U7759 (N_7759,N_1463,N_3999);
nand U7760 (N_7760,N_5683,N_4691);
or U7761 (N_7761,N_2856,N_407);
and U7762 (N_7762,N_2858,N_5980);
or U7763 (N_7763,N_558,N_3088);
nand U7764 (N_7764,N_5162,N_2772);
nand U7765 (N_7765,N_4170,N_3663);
or U7766 (N_7766,N_4720,N_5638);
nand U7767 (N_7767,N_3785,N_5973);
and U7768 (N_7768,N_931,N_3749);
or U7769 (N_7769,N_3691,N_3760);
xnor U7770 (N_7770,N_1607,N_1350);
nor U7771 (N_7771,N_5260,N_4669);
xnor U7772 (N_7772,N_2162,N_3030);
and U7773 (N_7773,N_2366,N_1886);
nor U7774 (N_7774,N_5139,N_2453);
nand U7775 (N_7775,N_615,N_2082);
nand U7776 (N_7776,N_798,N_5469);
nand U7777 (N_7777,N_756,N_1558);
nor U7778 (N_7778,N_1544,N_1095);
nor U7779 (N_7779,N_4777,N_1339);
nor U7780 (N_7780,N_5877,N_2245);
and U7781 (N_7781,N_1623,N_6050);
nor U7782 (N_7782,N_4451,N_1903);
nand U7783 (N_7783,N_353,N_1288);
and U7784 (N_7784,N_4753,N_716);
and U7785 (N_7785,N_4826,N_5925);
and U7786 (N_7786,N_2205,N_6141);
xor U7787 (N_7787,N_1242,N_3418);
xnor U7788 (N_7788,N_4663,N_5674);
nand U7789 (N_7789,N_5124,N_4887);
nor U7790 (N_7790,N_2108,N_2182);
and U7791 (N_7791,N_796,N_595);
or U7792 (N_7792,N_6018,N_3817);
or U7793 (N_7793,N_1831,N_3328);
nand U7794 (N_7794,N_646,N_3809);
nand U7795 (N_7795,N_28,N_1664);
and U7796 (N_7796,N_5546,N_2101);
nand U7797 (N_7797,N_4571,N_5623);
nor U7798 (N_7798,N_4538,N_228);
nor U7799 (N_7799,N_261,N_4999);
or U7800 (N_7800,N_1775,N_6014);
nand U7801 (N_7801,N_4266,N_4567);
nand U7802 (N_7802,N_1133,N_3835);
nand U7803 (N_7803,N_5457,N_1237);
or U7804 (N_7804,N_5890,N_199);
or U7805 (N_7805,N_5453,N_5088);
nor U7806 (N_7806,N_273,N_536);
or U7807 (N_7807,N_4046,N_4664);
or U7808 (N_7808,N_4084,N_5955);
xor U7809 (N_7809,N_1215,N_1185);
nand U7810 (N_7810,N_1037,N_4881);
nor U7811 (N_7811,N_2099,N_1053);
and U7812 (N_7812,N_3134,N_6020);
or U7813 (N_7813,N_5081,N_2385);
nand U7814 (N_7814,N_5949,N_3086);
and U7815 (N_7815,N_4639,N_3557);
nand U7816 (N_7816,N_3073,N_1100);
and U7817 (N_7817,N_4591,N_762);
and U7818 (N_7818,N_2574,N_3739);
nand U7819 (N_7819,N_614,N_2112);
or U7820 (N_7820,N_3079,N_3877);
and U7821 (N_7821,N_3581,N_6004);
and U7822 (N_7822,N_1809,N_2064);
and U7823 (N_7823,N_665,N_4059);
or U7824 (N_7824,N_2651,N_1209);
nand U7825 (N_7825,N_5755,N_4648);
or U7826 (N_7826,N_367,N_4793);
or U7827 (N_7827,N_4965,N_5480);
nor U7828 (N_7828,N_3559,N_5288);
nor U7829 (N_7829,N_5472,N_4413);
or U7830 (N_7830,N_3931,N_5049);
and U7831 (N_7831,N_4152,N_3474);
or U7832 (N_7832,N_849,N_1666);
nor U7833 (N_7833,N_1018,N_975);
or U7834 (N_7834,N_582,N_231);
and U7835 (N_7835,N_2784,N_4136);
nor U7836 (N_7836,N_5208,N_1924);
or U7837 (N_7837,N_5593,N_4643);
or U7838 (N_7838,N_291,N_453);
and U7839 (N_7839,N_4222,N_2093);
xor U7840 (N_7840,N_6071,N_200);
and U7841 (N_7841,N_2201,N_1395);
nand U7842 (N_7842,N_4338,N_2782);
nor U7843 (N_7843,N_2724,N_5580);
and U7844 (N_7844,N_653,N_3726);
or U7845 (N_7845,N_3753,N_693);
xor U7846 (N_7846,N_4583,N_1893);
xnor U7847 (N_7847,N_2324,N_5294);
nor U7848 (N_7848,N_3235,N_2583);
and U7849 (N_7849,N_3890,N_3744);
nor U7850 (N_7850,N_391,N_3741);
and U7851 (N_7851,N_702,N_1072);
xnor U7852 (N_7852,N_5029,N_3668);
or U7853 (N_7853,N_658,N_4868);
nor U7854 (N_7854,N_2746,N_3292);
nand U7855 (N_7855,N_5506,N_2768);
nor U7856 (N_7856,N_1663,N_3771);
nand U7857 (N_7857,N_3468,N_1160);
and U7858 (N_7858,N_518,N_5078);
and U7859 (N_7859,N_459,N_3678);
or U7860 (N_7860,N_1458,N_5924);
or U7861 (N_7861,N_121,N_4010);
nand U7862 (N_7862,N_5329,N_3707);
nand U7863 (N_7863,N_433,N_3111);
nor U7864 (N_7864,N_4864,N_3183);
xnor U7865 (N_7865,N_5537,N_854);
nor U7866 (N_7866,N_1255,N_1669);
xnor U7867 (N_7867,N_4436,N_4435);
and U7868 (N_7868,N_1415,N_584);
nor U7869 (N_7869,N_2285,N_3287);
nor U7870 (N_7870,N_160,N_3914);
or U7871 (N_7871,N_3166,N_6088);
and U7872 (N_7872,N_4110,N_5965);
or U7873 (N_7873,N_30,N_4499);
nand U7874 (N_7874,N_5449,N_5284);
and U7875 (N_7875,N_2648,N_2613);
nand U7876 (N_7876,N_5756,N_6092);
and U7877 (N_7877,N_2146,N_4045);
or U7878 (N_7878,N_2896,N_3975);
nor U7879 (N_7879,N_3360,N_5191);
nand U7880 (N_7880,N_2979,N_3317);
nand U7881 (N_7881,N_2121,N_2315);
and U7882 (N_7882,N_5117,N_2909);
and U7883 (N_7883,N_147,N_4202);
and U7884 (N_7884,N_1472,N_4819);
nand U7885 (N_7885,N_1828,N_20);
and U7886 (N_7886,N_616,N_3611);
or U7887 (N_7887,N_4158,N_970);
nor U7888 (N_7888,N_5400,N_5154);
or U7889 (N_7889,N_3669,N_5658);
nand U7890 (N_7890,N_1022,N_5591);
xnor U7891 (N_7891,N_2998,N_4581);
nand U7892 (N_7892,N_2176,N_3706);
nand U7893 (N_7893,N_5093,N_1030);
or U7894 (N_7894,N_5529,N_5248);
xnor U7895 (N_7895,N_2797,N_1811);
or U7896 (N_7896,N_944,N_4808);
nor U7897 (N_7897,N_3161,N_613);
nand U7898 (N_7898,N_2001,N_245);
and U7899 (N_7899,N_4437,N_5107);
nor U7900 (N_7900,N_4281,N_3356);
nor U7901 (N_7901,N_2153,N_4428);
and U7902 (N_7902,N_2942,N_4324);
nand U7903 (N_7903,N_842,N_2994);
and U7904 (N_7904,N_2999,N_3758);
and U7905 (N_7905,N_5479,N_4481);
nand U7906 (N_7906,N_5061,N_4477);
nor U7907 (N_7907,N_3503,N_3278);
and U7908 (N_7908,N_3495,N_2920);
nand U7909 (N_7909,N_5395,N_3450);
xnor U7910 (N_7910,N_3715,N_5775);
and U7911 (N_7911,N_5907,N_3864);
nand U7912 (N_7912,N_2774,N_3719);
nor U7913 (N_7913,N_4278,N_5796);
nor U7914 (N_7914,N_2078,N_4576);
xor U7915 (N_7915,N_3787,N_3395);
nand U7916 (N_7916,N_739,N_612);
nor U7917 (N_7917,N_2125,N_5662);
and U7918 (N_7918,N_4271,N_881);
xor U7919 (N_7919,N_2577,N_2747);
nand U7920 (N_7920,N_5816,N_742);
or U7921 (N_7921,N_2652,N_3261);
nand U7922 (N_7922,N_6138,N_1739);
and U7923 (N_7923,N_2190,N_5243);
xor U7924 (N_7924,N_4056,N_2890);
xnor U7925 (N_7925,N_2693,N_1438);
and U7926 (N_7926,N_4525,N_1508);
and U7927 (N_7927,N_2665,N_509);
nand U7928 (N_7928,N_5065,N_1796);
and U7929 (N_7929,N_1842,N_5241);
nand U7930 (N_7930,N_1734,N_4267);
nand U7931 (N_7931,N_356,N_2412);
or U7932 (N_7932,N_1003,N_4356);
and U7933 (N_7933,N_5635,N_3125);
xor U7934 (N_7934,N_1029,N_2717);
or U7935 (N_7935,N_651,N_3228);
nand U7936 (N_7936,N_5273,N_1145);
and U7937 (N_7937,N_4687,N_5712);
and U7938 (N_7938,N_1060,N_4);
and U7939 (N_7939,N_1507,N_393);
or U7940 (N_7940,N_4293,N_5820);
xor U7941 (N_7941,N_2850,N_4636);
nor U7942 (N_7942,N_6185,N_378);
and U7943 (N_7943,N_2380,N_368);
nand U7944 (N_7944,N_4953,N_2480);
or U7945 (N_7945,N_51,N_902);
xor U7946 (N_7946,N_3428,N_3179);
nor U7947 (N_7947,N_4132,N_4997);
and U7948 (N_7948,N_1444,N_1531);
nor U7949 (N_7949,N_981,N_2401);
nand U7950 (N_7950,N_5958,N_1973);
or U7951 (N_7951,N_1690,N_1304);
or U7952 (N_7952,N_4474,N_5682);
or U7953 (N_7953,N_3856,N_2963);
nand U7954 (N_7954,N_3080,N_1385);
and U7955 (N_7955,N_1885,N_2799);
nand U7956 (N_7956,N_4175,N_1727);
and U7957 (N_7957,N_1536,N_2466);
and U7958 (N_7958,N_5541,N_4065);
nor U7959 (N_7959,N_2662,N_4154);
nor U7960 (N_7960,N_890,N_3112);
nor U7961 (N_7961,N_75,N_1612);
nor U7962 (N_7962,N_1858,N_2026);
nand U7963 (N_7963,N_3591,N_3458);
or U7964 (N_7964,N_600,N_2486);
nor U7965 (N_7965,N_218,N_4802);
nand U7966 (N_7966,N_403,N_1067);
and U7967 (N_7967,N_1929,N_5548);
or U7968 (N_7968,N_5051,N_3353);
and U7969 (N_7969,N_2597,N_2500);
or U7970 (N_7970,N_3153,N_832);
or U7971 (N_7971,N_485,N_3226);
nand U7972 (N_7972,N_2585,N_4937);
and U7973 (N_7973,N_631,N_3479);
nor U7974 (N_7974,N_130,N_3927);
or U7975 (N_7975,N_1977,N_1190);
and U7976 (N_7976,N_45,N_2545);
nor U7977 (N_7977,N_6209,N_4910);
nand U7978 (N_7978,N_5476,N_5811);
or U7979 (N_7979,N_2113,N_5779);
nor U7980 (N_7980,N_5964,N_5691);
xnor U7981 (N_7981,N_2910,N_4889);
xor U7982 (N_7982,N_1855,N_4393);
nor U7983 (N_7983,N_5300,N_1802);
nand U7984 (N_7984,N_2958,N_5236);
and U7985 (N_7985,N_2670,N_3880);
or U7986 (N_7986,N_3457,N_1106);
and U7987 (N_7987,N_225,N_3090);
nand U7988 (N_7988,N_1450,N_471);
or U7989 (N_7989,N_3019,N_1769);
and U7990 (N_7990,N_678,N_5777);
or U7991 (N_7991,N_2114,N_1684);
and U7992 (N_7992,N_3345,N_1759);
nand U7993 (N_7993,N_2948,N_3362);
or U7994 (N_7994,N_4561,N_1332);
or U7995 (N_7995,N_1576,N_4032);
or U7996 (N_7996,N_4961,N_4403);
or U7997 (N_7997,N_3350,N_5474);
or U7998 (N_7998,N_1154,N_5665);
nor U7999 (N_7999,N_3998,N_2592);
or U8000 (N_8000,N_181,N_154);
or U8001 (N_8001,N_5885,N_2911);
nand U8002 (N_8002,N_5880,N_1902);
or U8003 (N_8003,N_2916,N_1194);
or U8004 (N_8004,N_5363,N_3052);
nand U8005 (N_8005,N_4155,N_4628);
nand U8006 (N_8006,N_3145,N_4120);
and U8007 (N_8007,N_5459,N_2960);
nor U8008 (N_8008,N_117,N_2645);
or U8009 (N_8009,N_2842,N_1722);
xor U8010 (N_8010,N_4093,N_5178);
nand U8011 (N_8011,N_3738,N_2650);
and U8012 (N_8012,N_2029,N_3554);
and U8013 (N_8013,N_6199,N_1113);
or U8014 (N_8014,N_1314,N_2990);
and U8015 (N_8015,N_4560,N_5377);
nand U8016 (N_8016,N_1981,N_620);
nand U8017 (N_8017,N_475,N_3012);
nand U8018 (N_8018,N_1217,N_4274);
nor U8019 (N_8019,N_2569,N_3597);
and U8020 (N_8020,N_2869,N_2596);
or U8021 (N_8021,N_5757,N_2303);
or U8022 (N_8022,N_6054,N_3405);
nand U8023 (N_8023,N_1324,N_5146);
xor U8024 (N_8024,N_3751,N_4608);
and U8025 (N_8025,N_1378,N_5855);
nand U8026 (N_8026,N_2643,N_2178);
xnor U8027 (N_8027,N_2964,N_1238);
nor U8028 (N_8028,N_3314,N_3674);
or U8029 (N_8029,N_1776,N_3979);
xor U8030 (N_8030,N_6235,N_2773);
nand U8031 (N_8031,N_3737,N_1123);
nor U8032 (N_8032,N_1568,N_132);
and U8033 (N_8033,N_5615,N_5471);
and U8034 (N_8034,N_3059,N_5360);
nand U8035 (N_8035,N_5069,N_4468);
nor U8036 (N_8036,N_2414,N_1740);
nor U8037 (N_8037,N_3366,N_998);
nor U8038 (N_8038,N_5669,N_421);
or U8039 (N_8039,N_974,N_222);
nor U8040 (N_8040,N_4517,N_1938);
or U8041 (N_8041,N_4711,N_814);
or U8042 (N_8042,N_4962,N_2846);
nand U8043 (N_8043,N_3906,N_5198);
or U8044 (N_8044,N_3823,N_4250);
nand U8045 (N_8045,N_4972,N_2002);
nor U8046 (N_8046,N_5252,N_2807);
nor U8047 (N_8047,N_3855,N_449);
xnor U8048 (N_8048,N_5057,N_4726);
nand U8049 (N_8049,N_4075,N_3750);
and U8050 (N_8050,N_993,N_1423);
and U8051 (N_8051,N_5142,N_306);
nor U8052 (N_8052,N_5018,N_3013);
and U8053 (N_8053,N_2275,N_1448);
nand U8054 (N_8054,N_1900,N_390);
and U8055 (N_8055,N_2471,N_5497);
or U8056 (N_8056,N_5494,N_3186);
xnor U8057 (N_8057,N_1525,N_5730);
xor U8058 (N_8058,N_6236,N_5417);
nand U8059 (N_8059,N_5706,N_1117);
or U8060 (N_8060,N_2570,N_4246);
nor U8061 (N_8061,N_4311,N_299);
nand U8062 (N_8062,N_1899,N_4715);
nand U8063 (N_8063,N_2934,N_3312);
nor U8064 (N_8064,N_504,N_2464);
or U8065 (N_8065,N_5823,N_284);
and U8066 (N_8066,N_3044,N_4964);
and U8067 (N_8067,N_5456,N_3617);
and U8068 (N_8068,N_5101,N_3330);
and U8069 (N_8069,N_5914,N_3680);
or U8070 (N_8070,N_4653,N_1271);
nor U8071 (N_8071,N_4626,N_4423);
nor U8072 (N_8072,N_3143,N_5619);
or U8073 (N_8073,N_821,N_5598);
nor U8074 (N_8074,N_5767,N_5083);
and U8075 (N_8075,N_4599,N_1157);
nor U8076 (N_8076,N_4197,N_2637);
or U8077 (N_8077,N_3294,N_5379);
nor U8078 (N_8078,N_286,N_6110);
nand U8079 (N_8079,N_1517,N_733);
nand U8080 (N_8080,N_4051,N_6115);
and U8081 (N_8081,N_94,N_3510);
nor U8082 (N_8082,N_1087,N_2035);
xnor U8083 (N_8083,N_2306,N_2956);
nand U8084 (N_8084,N_2733,N_5981);
nand U8085 (N_8085,N_3584,N_6072);
and U8086 (N_8086,N_5326,N_5333);
and U8087 (N_8087,N_2376,N_1426);
and U8088 (N_8088,N_5145,N_2459);
nor U8089 (N_8089,N_4371,N_2335);
xnor U8090 (N_8090,N_3871,N_4243);
nor U8091 (N_8091,N_56,N_4667);
nand U8092 (N_8092,N_5656,N_586);
or U8093 (N_8093,N_1244,N_5632);
and U8094 (N_8094,N_2587,N_2897);
and U8095 (N_8095,N_1144,N_3643);
and U8096 (N_8096,N_3788,N_1261);
nand U8097 (N_8097,N_5736,N_2042);
nor U8098 (N_8098,N_3905,N_3026);
or U8099 (N_8099,N_2658,N_5858);
xor U8100 (N_8100,N_3482,N_5089);
xnor U8101 (N_8101,N_768,N_2425);
nand U8102 (N_8102,N_6101,N_5774);
nand U8103 (N_8103,N_608,N_886);
nor U8104 (N_8104,N_4041,N_2647);
and U8105 (N_8105,N_1466,N_6105);
and U8106 (N_8106,N_654,N_2668);
and U8107 (N_8107,N_891,N_1147);
and U8108 (N_8108,N_718,N_4021);
and U8109 (N_8109,N_2630,N_750);
xnor U8110 (N_8110,N_4712,N_1750);
nor U8111 (N_8111,N_4452,N_2787);
or U8112 (N_8112,N_3604,N_1278);
nand U8113 (N_8113,N_4166,N_6099);
and U8114 (N_8114,N_3417,N_4167);
nand U8115 (N_8115,N_1077,N_4201);
or U8116 (N_8116,N_4399,N_462);
nor U8117 (N_8117,N_3924,N_1743);
nor U8118 (N_8118,N_1680,N_4456);
nor U8119 (N_8119,N_3083,N_6121);
or U8120 (N_8120,N_107,N_4092);
and U8121 (N_8121,N_740,N_3919);
and U8122 (N_8122,N_2792,N_5345);
or U8123 (N_8123,N_5904,N_1793);
and U8124 (N_8124,N_542,N_4472);
or U8125 (N_8125,N_4622,N_4485);
xnor U8126 (N_8126,N_3609,N_688);
and U8127 (N_8127,N_3940,N_5910);
nor U8128 (N_8128,N_4550,N_3316);
or U8129 (N_8129,N_4406,N_1807);
and U8130 (N_8130,N_4001,N_790);
or U8131 (N_8131,N_2531,N_2223);
and U8132 (N_8132,N_3060,N_6042);
or U8133 (N_8133,N_3891,N_917);
or U8134 (N_8134,N_1,N_5744);
or U8135 (N_8135,N_556,N_2572);
and U8136 (N_8136,N_2794,N_3742);
nor U8137 (N_8137,N_5947,N_1564);
and U8138 (N_8138,N_1541,N_1815);
nand U8139 (N_8139,N_2354,N_5831);
and U8140 (N_8140,N_1861,N_6100);
and U8141 (N_8141,N_956,N_3368);
xnor U8142 (N_8142,N_3613,N_438);
and U8143 (N_8143,N_2519,N_4816);
nor U8144 (N_8144,N_3214,N_3636);
nand U8145 (N_8145,N_4676,N_635);
nor U8146 (N_8146,N_5362,N_5505);
xor U8147 (N_8147,N_1320,N_1820);
nor U8148 (N_8148,N_184,N_5388);
nor U8149 (N_8149,N_5942,N_5543);
nand U8150 (N_8150,N_4095,N_2786);
nor U8151 (N_8151,N_5601,N_2537);
and U8152 (N_8152,N_5164,N_4509);
nand U8153 (N_8153,N_3142,N_4315);
xor U8154 (N_8154,N_3761,N_2621);
nand U8155 (N_8155,N_214,N_3119);
and U8156 (N_8156,N_6247,N_1895);
and U8157 (N_8157,N_2781,N_2440);
nor U8158 (N_8158,N_3274,N_4037);
and U8159 (N_8159,N_1380,N_2649);
and U8160 (N_8160,N_2092,N_2603);
or U8161 (N_8161,N_3102,N_4082);
nand U8162 (N_8162,N_1356,N_848);
xor U8163 (N_8163,N_2120,N_6197);
nand U8164 (N_8164,N_2071,N_1296);
xnor U8165 (N_8165,N_4699,N_2171);
or U8166 (N_8166,N_3549,N_2279);
and U8167 (N_8167,N_2968,N_1151);
xnor U8168 (N_8168,N_5968,N_1189);
nand U8169 (N_8169,N_3064,N_6080);
and U8170 (N_8170,N_2887,N_985);
xor U8171 (N_8171,N_3124,N_4067);
nand U8172 (N_8172,N_2884,N_4187);
xnor U8173 (N_8173,N_2512,N_2051);
nor U8174 (N_8174,N_4454,N_5331);
or U8175 (N_8175,N_1588,N_5070);
and U8176 (N_8176,N_6239,N_1512);
and U8177 (N_8177,N_4484,N_236);
or U8178 (N_8178,N_3697,N_5868);
xnor U8179 (N_8179,N_4502,N_5527);
xnor U8180 (N_8180,N_4180,N_3141);
and U8181 (N_8181,N_1629,N_5427);
nor U8182 (N_8182,N_5835,N_5722);
or U8183 (N_8183,N_385,N_5945);
nor U8184 (N_8184,N_866,N_2875);
nor U8185 (N_8185,N_1969,N_1407);
xnor U8186 (N_8186,N_6127,N_5701);
nor U8187 (N_8187,N_1181,N_1946);
or U8188 (N_8188,N_590,N_4546);
nor U8189 (N_8189,N_496,N_3759);
xnor U8190 (N_8190,N_4048,N_3631);
and U8191 (N_8191,N_803,N_1601);
and U8192 (N_8192,N_2161,N_1121);
nor U8193 (N_8193,N_643,N_644);
or U8194 (N_8194,N_3531,N_1786);
or U8195 (N_8195,N_6017,N_5729);
xnor U8196 (N_8196,N_1901,N_2372);
nand U8197 (N_8197,N_2673,N_907);
nor U8198 (N_8198,N_5204,N_4183);
nand U8199 (N_8199,N_6009,N_4328);
nor U8200 (N_8200,N_1460,N_5610);
and U8201 (N_8201,N_1298,N_3152);
nand U8202 (N_8202,N_5790,N_4405);
or U8203 (N_8203,N_4566,N_3178);
and U8204 (N_8204,N_776,N_3414);
and U8205 (N_8205,N_4841,N_5693);
xor U8206 (N_8206,N_724,N_1565);
nand U8207 (N_8207,N_5533,N_6060);
xnor U8208 (N_8208,N_2472,N_6106);
and U8209 (N_8209,N_1582,N_2939);
and U8210 (N_8210,N_1867,N_5116);
nor U8211 (N_8211,N_2221,N_655);
nor U8212 (N_8212,N_2157,N_5025);
and U8213 (N_8213,N_6067,N_3151);
nor U8214 (N_8214,N_5034,N_5556);
or U8215 (N_8215,N_2403,N_4139);
nand U8216 (N_8216,N_1955,N_4551);
nand U8217 (N_8217,N_3401,N_2361);
or U8218 (N_8218,N_321,N_2281);
nand U8219 (N_8219,N_1071,N_3869);
or U8220 (N_8220,N_3081,N_3411);
or U8221 (N_8221,N_606,N_5799);
nor U8222 (N_8222,N_3938,N_969);
xnor U8223 (N_8223,N_5800,N_5657);
nor U8224 (N_8224,N_2609,N_3994);
or U8225 (N_8225,N_2742,N_2465);
nand U8226 (N_8226,N_4765,N_1245);
nor U8227 (N_8227,N_4086,N_239);
nand U8228 (N_8228,N_4956,N_5063);
nor U8229 (N_8229,N_1632,N_1026);
and U8230 (N_8230,N_3875,N_6220);
and U8231 (N_8231,N_4782,N_5275);
nand U8232 (N_8232,N_4943,N_4344);
nor U8233 (N_8233,N_3172,N_3326);
xnor U8234 (N_8234,N_3958,N_5339);
and U8235 (N_8235,N_1430,N_4604);
xor U8236 (N_8236,N_3837,N_5664);
and U8237 (N_8237,N_3380,N_3808);
nand U8238 (N_8238,N_1963,N_5951);
and U8239 (N_8239,N_3128,N_3394);
nand U8240 (N_8240,N_3889,N_2679);
and U8241 (N_8241,N_767,N_2481);
and U8242 (N_8242,N_3916,N_2103);
and U8243 (N_8243,N_664,N_5011);
and U8244 (N_8244,N_50,N_856);
nor U8245 (N_8245,N_5986,N_1873);
nor U8246 (N_8246,N_3725,N_4611);
or U8247 (N_8247,N_4590,N_77);
and U8248 (N_8248,N_701,N_49);
or U8249 (N_8249,N_4812,N_1918);
nand U8250 (N_8250,N_4606,N_5007);
or U8251 (N_8251,N_844,N_5312);
or U8252 (N_8252,N_2669,N_174);
or U8253 (N_8253,N_801,N_5438);
nand U8254 (N_8254,N_1445,N_1634);
and U8255 (N_8255,N_657,N_5262);
nand U8256 (N_8256,N_1310,N_6063);
or U8257 (N_8257,N_224,N_4717);
nor U8258 (N_8258,N_4493,N_410);
nor U8259 (N_8259,N_3097,N_2427);
xor U8260 (N_8260,N_5511,N_2776);
or U8261 (N_8261,N_4681,N_3639);
or U8262 (N_8262,N_1697,N_4190);
and U8263 (N_8263,N_3853,N_1756);
nor U8264 (N_8264,N_3422,N_4107);
xor U8265 (N_8265,N_5496,N_5123);
or U8266 (N_8266,N_6160,N_1398);
xor U8267 (N_8267,N_1543,N_2524);
xnor U8268 (N_8268,N_4925,N_5687);
or U8269 (N_8269,N_721,N_5524);
xor U8270 (N_8270,N_59,N_3729);
or U8271 (N_8271,N_6056,N_1315);
or U8272 (N_8272,N_3821,N_5919);
and U8273 (N_8273,N_3311,N_3756);
nand U8274 (N_8274,N_267,N_3881);
xor U8275 (N_8275,N_2231,N_1616);
nand U8276 (N_8276,N_2925,N_452);
and U8277 (N_8277,N_5874,N_717);
nor U8278 (N_8278,N_5961,N_5654);
nor U8279 (N_8279,N_1677,N_2878);
nor U8280 (N_8280,N_2515,N_2978);
and U8281 (N_8281,N_4668,N_738);
xnor U8282 (N_8282,N_3536,N_5436);
nand U8283 (N_8283,N_2276,N_1832);
or U8284 (N_8284,N_5738,N_241);
and U8285 (N_8285,N_5499,N_2140);
nand U8286 (N_8286,N_442,N_3122);
nand U8287 (N_8287,N_3155,N_3399);
or U8288 (N_8288,N_591,N_446);
nand U8289 (N_8289,N_5058,N_2795);
nor U8290 (N_8290,N_1086,N_4055);
xnor U8291 (N_8291,N_4332,N_920);
and U8292 (N_8292,N_5152,N_2261);
or U8293 (N_8293,N_3446,N_2714);
xnor U8294 (N_8294,N_1316,N_212);
nor U8295 (N_8295,N_4013,N_1364);
or U8296 (N_8296,N_5768,N_5305);
and U8297 (N_8297,N_841,N_5040);
or U8298 (N_8298,N_5285,N_2413);
nand U8299 (N_8299,N_4708,N_341);
and U8300 (N_8300,N_4983,N_5451);
nor U8301 (N_8301,N_4852,N_2754);
or U8302 (N_8302,N_1128,N_5997);
or U8303 (N_8303,N_4780,N_67);
nor U8304 (N_8304,N_2757,N_6061);
nor U8305 (N_8305,N_1763,N_1683);
nor U8306 (N_8306,N_1369,N_1657);
and U8307 (N_8307,N_587,N_2764);
nor U8308 (N_8308,N_5631,N_1827);
nand U8309 (N_8309,N_5634,N_372);
nand U8310 (N_8310,N_1515,N_1391);
xor U8311 (N_8311,N_2834,N_279);
and U8312 (N_8312,N_4756,N_5611);
nand U8313 (N_8313,N_2244,N_3648);
and U8314 (N_8314,N_5002,N_5071);
nor U8315 (N_8315,N_3384,N_3276);
nor U8316 (N_8316,N_4421,N_2180);
xnor U8317 (N_8317,N_3277,N_3307);
or U8318 (N_8318,N_2908,N_6218);
nand U8319 (N_8319,N_5585,N_2096);
and U8320 (N_8320,N_2721,N_860);
nor U8321 (N_8321,N_4888,N_1091);
or U8322 (N_8322,N_853,N_4087);
or U8323 (N_8323,N_6045,N_4885);
nor U8324 (N_8324,N_2677,N_2756);
or U8325 (N_8325,N_1269,N_3359);
and U8326 (N_8326,N_400,N_1505);
and U8327 (N_8327,N_148,N_2294);
nor U8328 (N_8328,N_5134,N_5044);
and U8329 (N_8329,N_4430,N_4607);
xor U8330 (N_8330,N_5401,N_930);
nand U8331 (N_8331,N_52,N_1492);
or U8332 (N_8332,N_4846,N_3553);
and U8333 (N_8333,N_3950,N_3038);
nor U8334 (N_8334,N_5766,N_4319);
nor U8335 (N_8335,N_3908,N_3685);
nor U8336 (N_8336,N_1649,N_191);
nand U8337 (N_8337,N_1101,N_2847);
and U8338 (N_8338,N_1984,N_5368);
nand U8339 (N_8339,N_3426,N_2599);
nand U8340 (N_8340,N_2133,N_240);
and U8341 (N_8341,N_324,N_2826);
nor U8342 (N_8342,N_2840,N_4184);
and U8343 (N_8343,N_3444,N_6198);
xnor U8344 (N_8344,N_2006,N_4077);
nor U8345 (N_8345,N_4749,N_6075);
xor U8346 (N_8346,N_2449,N_2045);
nand U8347 (N_8347,N_2640,N_3318);
nand U8348 (N_8348,N_4205,N_1293);
nand U8349 (N_8349,N_2222,N_1857);
xnor U8350 (N_8350,N_2702,N_4353);
or U8351 (N_8351,N_158,N_1747);
nand U8352 (N_8352,N_3963,N_4376);
nor U8353 (N_8353,N_2628,N_4633);
or U8354 (N_8354,N_3365,N_2152);
nor U8355 (N_8355,N_1481,N_903);
or U8356 (N_8356,N_826,N_1459);
nand U8357 (N_8357,N_2867,N_5879);
and U8358 (N_8358,N_874,N_2543);
and U8359 (N_8359,N_4369,N_2337);
or U8360 (N_8360,N_6243,N_2720);
nand U8361 (N_8361,N_2862,N_3055);
and U8362 (N_8362,N_4666,N_2675);
nand U8363 (N_8363,N_196,N_3031);
nand U8364 (N_8364,N_3913,N_5487);
nand U8365 (N_8365,N_144,N_5484);
nor U8366 (N_8366,N_895,N_2237);
or U8367 (N_8367,N_5396,N_2766);
or U8368 (N_8368,N_1012,N_6163);
and U8369 (N_8369,N_404,N_805);
or U8370 (N_8370,N_858,N_604);
and U8371 (N_8371,N_5475,N_3167);
nor U8372 (N_8372,N_3390,N_379);
and U8373 (N_8373,N_2314,N_1179);
and U8374 (N_8374,N_1976,N_3407);
or U8375 (N_8375,N_4382,N_6116);
nor U8376 (N_8376,N_2010,N_507);
xor U8377 (N_8377,N_921,N_6002);
nand U8378 (N_8378,N_4904,N_2485);
or U8379 (N_8379,N_271,N_2830);
and U8380 (N_8380,N_4195,N_685);
nand U8381 (N_8381,N_6016,N_5393);
xor U8382 (N_8382,N_2429,N_2713);
and U8383 (N_8383,N_585,N_5802);
nand U8384 (N_8384,N_5042,N_2043);
or U8385 (N_8385,N_1567,N_4117);
and U8386 (N_8386,N_4153,N_1370);
nand U8387 (N_8387,N_43,N_6006);
nand U8388 (N_8388,N_2936,N_5828);
xor U8389 (N_8389,N_3702,N_1667);
nor U8390 (N_8390,N_4936,N_3650);
and U8391 (N_8391,N_833,N_4097);
nor U8392 (N_8392,N_6203,N_1510);
and U8393 (N_8393,N_1912,N_3637);
nor U8394 (N_8394,N_3232,N_3101);
nor U8395 (N_8395,N_3339,N_1681);
and U8396 (N_8396,N_2260,N_4760);
xor U8397 (N_8397,N_347,N_5082);
and U8398 (N_8398,N_5186,N_5972);
nor U8399 (N_8399,N_5341,N_4302);
or U8400 (N_8400,N_468,N_3205);
nand U8401 (N_8401,N_409,N_771);
or U8402 (N_8402,N_1685,N_1362);
or U8403 (N_8403,N_84,N_2033);
and U8404 (N_8404,N_4411,N_2248);
and U8405 (N_8405,N_990,N_293);
or U8406 (N_8406,N_1143,N_1251);
and U8407 (N_8407,N_4901,N_3188);
nor U8408 (N_8408,N_5306,N_4519);
nand U8409 (N_8409,N_1699,N_3296);
and U8410 (N_8410,N_1841,N_316);
xor U8411 (N_8411,N_2633,N_5510);
nor U8412 (N_8412,N_2843,N_1330);
nand U8413 (N_8413,N_4247,N_4980);
nand U8414 (N_8414,N_6146,N_4105);
or U8415 (N_8415,N_1447,N_2976);
or U8416 (N_8416,N_373,N_973);
and U8417 (N_8417,N_6219,N_1199);
or U8418 (N_8418,N_1108,N_1042);
nor U8419 (N_8419,N_6201,N_489);
or U8420 (N_8420,N_5508,N_3748);
or U8421 (N_8421,N_1241,N_2876);
nor U8422 (N_8422,N_3866,N_3195);
and U8423 (N_8423,N_1606,N_4853);
nand U8424 (N_8424,N_531,N_189);
and U8425 (N_8425,N_2262,N_2967);
nand U8426 (N_8426,N_5183,N_5684);
nor U8427 (N_8427,N_959,N_5714);
nand U8428 (N_8428,N_583,N_2060);
nor U8429 (N_8429,N_1682,N_4313);
nand U8430 (N_8430,N_1762,N_3443);
or U8431 (N_8431,N_3361,N_6096);
nand U8432 (N_8432,N_1103,N_6034);
nor U8433 (N_8433,N_4359,N_4598);
and U8434 (N_8434,N_999,N_4236);
nor U8435 (N_8435,N_436,N_3492);
nand U8436 (N_8436,N_4367,N_1821);
or U8437 (N_8437,N_1367,N_4363);
or U8438 (N_8438,N_1084,N_4298);
xnor U8439 (N_8439,N_4064,N_3810);
nor U8440 (N_8440,N_1999,N_3398);
nand U8441 (N_8441,N_242,N_2516);
nor U8442 (N_8442,N_3481,N_1224);
nor U8443 (N_8443,N_5017,N_1176);
and U8444 (N_8444,N_3306,N_4923);
or U8445 (N_8445,N_2595,N_2957);
xnor U8446 (N_8446,N_5939,N_5231);
nand U8447 (N_8447,N_4632,N_2632);
or U8448 (N_8448,N_3671,N_4602);
or U8449 (N_8449,N_386,N_443);
xnor U8450 (N_8450,N_5789,N_4137);
and U8451 (N_8451,N_3652,N_5437);
xnor U8452 (N_8452,N_4507,N_4047);
and U8453 (N_8453,N_3047,N_1950);
nand U8454 (N_8454,N_38,N_2308);
nand U8455 (N_8455,N_1374,N_1055);
or U8456 (N_8456,N_5421,N_4004);
and U8457 (N_8457,N_4773,N_4703);
or U8458 (N_8458,N_3158,N_1771);
nand U8459 (N_8459,N_2359,N_2381);
nor U8460 (N_8460,N_3898,N_2284);
or U8461 (N_8461,N_5296,N_44);
or U8462 (N_8462,N_845,N_3433);
or U8463 (N_8463,N_1897,N_455);
xnor U8464 (N_8464,N_4040,N_4798);
nor U8465 (N_8465,N_2683,N_885);
nor U8466 (N_8466,N_1319,N_705);
nand U8467 (N_8467,N_1373,N_4416);
nor U8468 (N_8468,N_3512,N_603);
or U8469 (N_8469,N_4031,N_6164);
and U8470 (N_8470,N_3219,N_1230);
nand U8471 (N_8471,N_3222,N_757);
and U8472 (N_8472,N_5979,N_5432);
or U8473 (N_8473,N_939,N_5696);
and U8474 (N_8474,N_2555,N_5881);
xnor U8475 (N_8475,N_162,N_1795);
and U8476 (N_8476,N_2311,N_4455);
nand U8477 (N_8477,N_3614,N_16);
nand U8478 (N_8478,N_2003,N_2199);
nor U8479 (N_8479,N_5321,N_547);
and U8480 (N_8480,N_720,N_1246);
nor U8481 (N_8481,N_3632,N_2849);
or U8482 (N_8482,N_2280,N_675);
nor U8483 (N_8483,N_6134,N_3136);
nand U8484 (N_8484,N_992,N_3577);
nand U8485 (N_8485,N_1951,N_1094);
nand U8486 (N_8486,N_5193,N_3555);
or U8487 (N_8487,N_1446,N_3238);
or U8488 (N_8488,N_4619,N_1593);
nor U8489 (N_8489,N_4692,N_1501);
and U8490 (N_8490,N_941,N_1526);
or U8491 (N_8491,N_1493,N_1721);
nor U8492 (N_8492,N_5713,N_5458);
xnor U8493 (N_8493,N_3565,N_908);
or U8494 (N_8494,N_640,N_2735);
or U8495 (N_8495,N_1115,N_3629);
nor U8496 (N_8496,N_2700,N_4204);
nand U8497 (N_8497,N_4314,N_1714);
nor U8498 (N_8498,N_1187,N_6155);
nand U8499 (N_8499,N_6048,N_4501);
nand U8500 (N_8500,N_4834,N_5860);
or U8501 (N_8501,N_2398,N_2419);
nor U8502 (N_8502,N_3745,N_3945);
or U8503 (N_8503,N_5735,N_450);
xor U8504 (N_8504,N_5932,N_5626);
or U8505 (N_8505,N_5753,N_770);
nor U8506 (N_8506,N_123,N_933);
nand U8507 (N_8507,N_1468,N_1618);
nand U8508 (N_8508,N_3949,N_380);
xor U8509 (N_8509,N_787,N_5930);
xnor U8510 (N_8510,N_4207,N_5223);
and U8511 (N_8511,N_4068,N_3995);
or U8512 (N_8512,N_3387,N_451);
nand U8513 (N_8513,N_6062,N_4245);
nand U8514 (N_8514,N_5177,N_4960);
nor U8515 (N_8515,N_1522,N_713);
and U8516 (N_8516,N_1944,N_3241);
or U8517 (N_8517,N_5711,N_1413);
nand U8518 (N_8518,N_1801,N_4951);
and U8519 (N_8519,N_29,N_6094);
nand U8520 (N_8520,N_809,N_4991);
or U8521 (N_8521,N_4193,N_1562);
nor U8522 (N_8522,N_2405,N_1227);
nand U8523 (N_8523,N_3315,N_4223);
or U8524 (N_8524,N_2418,N_1712);
and U8525 (N_8525,N_3138,N_2941);
or U8526 (N_8526,N_1692,N_3934);
and U8527 (N_8527,N_3239,N_5526);
and U8528 (N_8528,N_2124,N_371);
and U8529 (N_8529,N_4559,N_5128);
nor U8530 (N_8530,N_551,N_1452);
nor U8531 (N_8531,N_478,N_5020);
nand U8532 (N_8532,N_589,N_3545);
xnor U8533 (N_8533,N_5783,N_789);
xnor U8534 (N_8534,N_3720,N_1206);
and U8535 (N_8535,N_4230,N_3174);
and U8536 (N_8536,N_3123,N_1947);
nor U8537 (N_8537,N_598,N_2206);
and U8538 (N_8538,N_599,N_882);
xnor U8539 (N_8539,N_4341,N_4303);
or U8540 (N_8540,N_369,N_4434);
or U8541 (N_8541,N_2240,N_1691);
nor U8542 (N_8542,N_5882,N_6140);
or U8543 (N_8543,N_5174,N_3040);
nor U8544 (N_8544,N_3688,N_971);
and U8545 (N_8545,N_563,N_4398);
nand U8546 (N_8546,N_2682,N_2833);
nand U8547 (N_8547,N_3460,N_6193);
nor U8548 (N_8548,N_277,N_2327);
nand U8549 (N_8549,N_2914,N_169);
nand U8550 (N_8550,N_2528,N_4908);
and U8551 (N_8551,N_1267,N_1513);
nor U8552 (N_8552,N_3692,N_5561);
nand U8553 (N_8553,N_2476,N_5340);
and U8554 (N_8554,N_2168,N_4409);
nor U8555 (N_8555,N_1635,N_2666);
nor U8556 (N_8556,N_3057,N_1150);
nor U8557 (N_8557,N_4071,N_734);
and U8558 (N_8558,N_677,N_5849);
and U8559 (N_8559,N_4288,N_2098);
and U8560 (N_8560,N_3765,N_3082);
nor U8561 (N_8561,N_4563,N_3920);
nor U8562 (N_8562,N_1139,N_5671);
nor U8563 (N_8563,N_4820,N_676);
nand U8564 (N_8564,N_2207,N_5734);
xor U8565 (N_8565,N_3812,N_3493);
nor U8566 (N_8566,N_474,N_3723);
nor U8567 (N_8567,N_2330,N_1758);
xor U8568 (N_8568,N_1294,N_1322);
nor U8569 (N_8569,N_4395,N_3948);
nand U8570 (N_8570,N_3815,N_295);
nand U8571 (N_8571,N_2736,N_1928);
and U8572 (N_8572,N_1868,N_2431);
and U8573 (N_8573,N_5573,N_2296);
nand U8574 (N_8574,N_5809,N_1784);
nor U8575 (N_8575,N_3587,N_958);
nand U8576 (N_8576,N_5772,N_512);
and U8577 (N_8577,N_3640,N_2576);
nand U8578 (N_8578,N_3298,N_5901);
nor U8579 (N_8579,N_1410,N_594);
nand U8580 (N_8580,N_3960,N_3230);
or U8581 (N_8581,N_3478,N_2641);
or U8582 (N_8582,N_2940,N_781);
nand U8583 (N_8583,N_3511,N_1779);
nand U8584 (N_8584,N_4318,N_3797);
nor U8585 (N_8585,N_5461,N_3974);
nand U8586 (N_8586,N_2117,N_4543);
xnor U8587 (N_8587,N_4862,N_1451);
nor U8588 (N_8588,N_5200,N_991);
nand U8589 (N_8589,N_246,N_2952);
nor U8590 (N_8590,N_1063,N_2189);
nor U8591 (N_8591,N_6137,N_1434);
and U8592 (N_8592,N_4486,N_5493);
nor U8593 (N_8593,N_1388,N_1129);
and U8594 (N_8594,N_937,N_166);
nand U8595 (N_8595,N_4700,N_5247);
xnor U8596 (N_8596,N_642,N_2758);
xnor U8597 (N_8597,N_124,N_1375);
and U8598 (N_8598,N_1300,N_1414);
nand U8599 (N_8599,N_3662,N_3540);
xnor U8600 (N_8600,N_4000,N_1243);
nor U8601 (N_8601,N_473,N_4721);
and U8602 (N_8602,N_5127,N_1109);
nand U8603 (N_8603,N_3508,N_3580);
and U8604 (N_8604,N_5335,N_6090);
nand U8605 (N_8605,N_3139,N_5589);
and U8606 (N_8606,N_2681,N_4850);
nor U8607 (N_8607,N_1798,N_1829);
xnor U8608 (N_8608,N_4534,N_4373);
nand U8609 (N_8609,N_2575,N_1461);
nor U8610 (N_8610,N_4030,N_6011);
and U8611 (N_8611,N_5584,N_4618);
or U8612 (N_8612,N_2816,N_2349);
nor U8613 (N_8613,N_177,N_3084);
or U8614 (N_8614,N_2063,N_4621);
or U8615 (N_8615,N_3618,N_3829);
xor U8616 (N_8616,N_1191,N_328);
nor U8617 (N_8617,N_314,N_1765);
nand U8618 (N_8618,N_6051,N_2710);
nor U8619 (N_8619,N_122,N_6211);
or U8620 (N_8620,N_6187,N_5933);
or U8621 (N_8621,N_1033,N_1329);
nor U8622 (N_8622,N_2540,N_5613);
and U8623 (N_8623,N_1989,N_4192);
nor U8624 (N_8624,N_4252,N_3477);
nor U8625 (N_8625,N_5710,N_1518);
nor U8626 (N_8626,N_819,N_1960);
and U8627 (N_8627,N_6230,N_6008);
nand U8628 (N_8628,N_2796,N_4300);
or U8629 (N_8629,N_817,N_111);
nor U8630 (N_8630,N_3054,N_2502);
nand U8631 (N_8631,N_5086,N_723);
and U8632 (N_8632,N_444,N_5108);
and U8633 (N_8633,N_3603,N_260);
and U8634 (N_8634,N_326,N_3074);
and U8635 (N_8635,N_2163,N_3878);
xnor U8636 (N_8636,N_2406,N_1207);
or U8637 (N_8637,N_1854,N_1478);
xnor U8638 (N_8638,N_3229,N_4159);
or U8639 (N_8639,N_1470,N_3068);
xor U8640 (N_8640,N_2024,N_5998);
nand U8641 (N_8641,N_1454,N_2122);
or U8642 (N_8642,N_4377,N_4397);
nand U8643 (N_8643,N_4277,N_818);
nand U8644 (N_8644,N_4003,N_4280);
and U8645 (N_8645,N_65,N_116);
nor U8646 (N_8646,N_1797,N_2142);
or U8647 (N_8647,N_484,N_4968);
or U8648 (N_8648,N_5704,N_1689);
and U8649 (N_8649,N_2126,N_1812);
nand U8650 (N_8650,N_3944,N_3946);
nor U8651 (N_8651,N_76,N_5408);
and U8652 (N_8652,N_2369,N_4918);
and U8653 (N_8653,N_5544,N_2895);
and U8654 (N_8654,N_1137,N_3329);
nor U8655 (N_8655,N_3085,N_4545);
nand U8656 (N_8656,N_909,N_523);
or U8657 (N_8657,N_469,N_1611);
nand U8658 (N_8658,N_5268,N_4912);
or U8659 (N_8659,N_430,N_4984);
or U8660 (N_8660,N_4256,N_1213);
nand U8661 (N_8661,N_5867,N_5975);
or U8662 (N_8662,N_4442,N_1420);
and U8663 (N_8663,N_709,N_280);
nand U8664 (N_8664,N_5739,N_2857);
xor U8665 (N_8665,N_1263,N_1085);
nand U8666 (N_8666,N_3334,N_1006);
nor U8667 (N_8667,N_5118,N_5092);
or U8668 (N_8668,N_1044,N_4088);
nand U8669 (N_8669,N_208,N_3374);
nor U8670 (N_8670,N_2145,N_3176);
or U8671 (N_8671,N_4946,N_5440);
or U8672 (N_8672,N_4684,N_3258);
and U8673 (N_8673,N_1630,N_359);
or U8674 (N_8674,N_4973,N_3266);
or U8675 (N_8675,N_253,N_4282);
nor U8676 (N_8676,N_1074,N_957);
or U8677 (N_8677,N_5050,N_2953);
nor U8678 (N_8678,N_2752,N_1847);
nand U8679 (N_8679,N_1186,N_1040);
nand U8680 (N_8680,N_2301,N_2602);
nor U8681 (N_8681,N_3965,N_6091);
xor U8682 (N_8682,N_3420,N_5625);
nand U8683 (N_8683,N_6184,N_1645);
xor U8684 (N_8684,N_3016,N_4283);
and U8685 (N_8685,N_3735,N_1068);
xor U8686 (N_8686,N_2325,N_480);
and U8687 (N_8687,N_630,N_2611);
or U8688 (N_8688,N_268,N_6079);
nor U8689 (N_8689,N_960,N_3523);
nand U8690 (N_8690,N_275,N_3413);
nand U8691 (N_8691,N_2259,N_3966);
or U8692 (N_8692,N_666,N_2439);
nor U8693 (N_8693,N_4125,N_1138);
nor U8694 (N_8694,N_5702,N_3734);
and U8695 (N_8695,N_704,N_5794);
nand U8696 (N_8696,N_820,N_3089);
xnor U8697 (N_8697,N_1090,N_2993);
xnor U8698 (N_8698,N_296,N_2463);
or U8699 (N_8699,N_4101,N_5927);
and U8700 (N_8700,N_3600,N_1202);
nand U8701 (N_8701,N_1859,N_5460);
or U8702 (N_8702,N_5886,N_64);
nor U8703 (N_8703,N_3146,N_216);
and U8704 (N_8704,N_6040,N_4941);
nor U8705 (N_8705,N_3448,N_1140);
and U8706 (N_8706,N_2194,N_5290);
or U8707 (N_8707,N_4899,N_5663);
nor U8708 (N_8708,N_3803,N_5232);
nor U8709 (N_8709,N_1671,N_3532);
and U8710 (N_8710,N_4842,N_2477);
or U8711 (N_8711,N_3802,N_4989);
and U8712 (N_8712,N_3675,N_876);
or U8713 (N_8713,N_204,N_2446);
or U8714 (N_8714,N_3263,N_186);
nor U8715 (N_8715,N_5956,N_5895);
nand U8716 (N_8716,N_5390,N_2072);
and U8717 (N_8717,N_5463,N_982);
nand U8718 (N_8718,N_4739,N_5795);
nor U8719 (N_8719,N_2488,N_2984);
nand U8720 (N_8720,N_6229,N_934);
nor U8721 (N_8721,N_3970,N_2791);
and U8722 (N_8722,N_5583,N_955);
or U8723 (N_8723,N_2179,N_1752);
nor U8724 (N_8724,N_4316,N_2062);
nor U8725 (N_8725,N_2553,N_5899);
or U8726 (N_8726,N_2160,N_4734);
nor U8727 (N_8727,N_290,N_5569);
nand U8728 (N_8728,N_870,N_792);
and U8729 (N_8729,N_5037,N_6086);
nand U8730 (N_8730,N_4902,N_1587);
or U8731 (N_8731,N_2821,N_2494);
and U8732 (N_8732,N_1098,N_5909);
and U8733 (N_8733,N_662,N_5016);
nor U8734 (N_8734,N_1833,N_1425);
and U8735 (N_8735,N_4100,N_632);
nor U8736 (N_8736,N_543,N_2580);
or U8737 (N_8737,N_5504,N_171);
or U8738 (N_8738,N_1916,N_602);
nor U8739 (N_8739,N_5586,N_952);
xor U8740 (N_8740,N_927,N_3169);
or U8741 (N_8741,N_829,N_5758);
nor U8742 (N_8742,N_2499,N_5502);
or U8743 (N_8743,N_3641,N_629);
or U8744 (N_8744,N_3191,N_3904);
nand U8745 (N_8745,N_3327,N_1432);
and U8746 (N_8746,N_914,N_1218);
and U8747 (N_8747,N_3240,N_66);
or U8748 (N_8748,N_5856,N_964);
or U8749 (N_8749,N_786,N_4465);
nand U8750 (N_8750,N_4347,N_2712);
nand U8751 (N_8751,N_861,N_5922);
and U8752 (N_8752,N_4920,N_1231);
nand U8753 (N_8753,N_3441,N_188);
and U8754 (N_8754,N_3789,N_5175);
nor U8755 (N_8755,N_1309,N_3651);
and U8756 (N_8756,N_3126,N_3382);
or U8757 (N_8757,N_5454,N_4683);
nor U8758 (N_8758,N_1088,N_3467);
nand U8759 (N_8759,N_3486,N_2441);
nor U8760 (N_8760,N_779,N_374);
xnor U8761 (N_8761,N_2220,N_4219);
and U8762 (N_8762,N_706,N_5976);
and U8763 (N_8763,N_3190,N_2450);
and U8764 (N_8764,N_5122,N_2980);
or U8765 (N_8765,N_569,N_4036);
and U8766 (N_8766,N_4856,N_1254);
or U8767 (N_8767,N_5422,N_1933);
nor U8768 (N_8768,N_1381,N_3389);
or U8769 (N_8769,N_3973,N_3284);
or U8770 (N_8770,N_2839,N_3993);
or U8771 (N_8771,N_1848,N_4478);
nor U8772 (N_8772,N_2074,N_5751);
nor U8773 (N_8773,N_1226,N_112);
and U8774 (N_8774,N_1114,N_2997);
and U8775 (N_8775,N_3848,N_815);
nand U8776 (N_8776,N_2663,N_5338);
nand U8777 (N_8777,N_3305,N_4860);
or U8778 (N_8778,N_5346,N_4763);
or U8779 (N_8779,N_2885,N_686);
xnor U8780 (N_8780,N_3528,N_804);
nand U8781 (N_8781,N_3078,N_5897);
xnor U8782 (N_8782,N_2790,N_2848);
or U8783 (N_8783,N_670,N_2388);
xnor U8784 (N_8784,N_1331,N_4746);
xnor U8785 (N_8785,N_2588,N_441);
nand U8786 (N_8786,N_2923,N_4039);
xnor U8787 (N_8787,N_1008,N_3695);
and U8788 (N_8788,N_3270,N_4129);
and U8789 (N_8789,N_1785,N_2229);
nand U8790 (N_8790,N_2642,N_4537);
and U8791 (N_8791,N_1200,N_3067);
nor U8792 (N_8792,N_4574,N_2771);
xor U8793 (N_8793,N_5103,N_4500);
and U8794 (N_8794,N_1534,N_5119);
and U8795 (N_8795,N_6206,N_3947);
and U8796 (N_8796,N_748,N_1789);
xnor U8797 (N_8797,N_5630,N_562);
nand U8798 (N_8798,N_2028,N_1921);
xnor U8799 (N_8799,N_351,N_4336);
and U8800 (N_8800,N_508,N_6215);
xnor U8801 (N_8801,N_5771,N_4128);
and U8802 (N_8802,N_1693,N_6246);
nand U8803 (N_8803,N_6077,N_2664);
or U8804 (N_8804,N_1910,N_689);
or U8805 (N_8805,N_1236,N_1569);
nor U8806 (N_8806,N_5303,N_2918);
or U8807 (N_8807,N_3730,N_2740);
nand U8808 (N_8808,N_5978,N_888);
or U8809 (N_8809,N_1790,N_1911);
nand U8810 (N_8810,N_5857,N_4216);
nand U8811 (N_8811,N_2148,N_3377);
and U8812 (N_8812,N_2298,N_5806);
and U8813 (N_8813,N_1079,N_5148);
xor U8814 (N_8814,N_5628,N_764);
or U8815 (N_8815,N_226,N_5839);
or U8816 (N_8816,N_1498,N_2434);
and U8817 (N_8817,N_1475,N_977);
nor U8818 (N_8818,N_133,N_3623);
nand U8819 (N_8819,N_5272,N_546);
or U8820 (N_8820,N_1125,N_3616);
and U8821 (N_8821,N_5507,N_4114);
and U8822 (N_8822,N_4249,N_5240);
nor U8823 (N_8823,N_3684,N_3297);
xnor U8824 (N_8824,N_5179,N_3131);
nor U8825 (N_8825,N_565,N_6073);
nand U8826 (N_8826,N_5900,N_5966);
or U8827 (N_8827,N_2866,N_765);
nor U8828 (N_8828,N_3432,N_824);
nor U8829 (N_8829,N_555,N_31);
nand U8830 (N_8830,N_4340,N_5261);
nor U8831 (N_8831,N_3857,N_2977);
and U8832 (N_8832,N_1760,N_5310);
and U8833 (N_8833,N_2473,N_5834);
nand U8834 (N_8834,N_2031,N_953);
nor U8835 (N_8835,N_2407,N_2150);
nor U8836 (N_8836,N_503,N_699);
xor U8837 (N_8837,N_339,N_4886);
nand U8838 (N_8838,N_5443,N_1718);
or U8839 (N_8839,N_2808,N_2370);
nand U8840 (N_8840,N_3964,N_2785);
and U8841 (N_8841,N_1469,N_4116);
or U8842 (N_8842,N_5892,N_1990);
xnor U8843 (N_8843,N_5873,N_3358);
and U8844 (N_8844,N_1942,N_3170);
and U8845 (N_8845,N_871,N_3267);
or U8846 (N_8846,N_5985,N_3118);
nand U8847 (N_8847,N_3037,N_2227);
and U8848 (N_8848,N_142,N_3099);
or U8849 (N_8849,N_5350,N_3024);
or U8850 (N_8850,N_527,N_2806);
nand U8851 (N_8851,N_5105,N_987);
nor U8852 (N_8852,N_4832,N_6154);
nor U8853 (N_8853,N_1502,N_4118);
xor U8854 (N_8854,N_205,N_2584);
nor U8855 (N_8855,N_4725,N_4595);
nor U8856 (N_8856,N_4958,N_4974);
or U8857 (N_8857,N_4579,N_5784);
or U8858 (N_8858,N_2818,N_4787);
and U8859 (N_8859,N_1600,N_2558);
and U8860 (N_8860,N_2690,N_3942);
and U8861 (N_8861,N_5221,N_1279);
nor U8862 (N_8862,N_3076,N_370);
or U8863 (N_8863,N_2844,N_3781);
nor U8864 (N_8864,N_1273,N_5429);
and U8865 (N_8865,N_2433,N_1906);
nand U8866 (N_8866,N_5404,N_5581);
nor U8867 (N_8867,N_90,N_5574);
xnor U8868 (N_8868,N_6039,N_4924);
nor U8869 (N_8869,N_4232,N_5211);
and U8870 (N_8870,N_4516,N_2514);
xor U8871 (N_8871,N_2257,N_1192);
nand U8872 (N_8872,N_5218,N_519);
and U8873 (N_8873,N_3813,N_5761);
and U8874 (N_8874,N_3177,N_5962);
or U8875 (N_8875,N_1748,N_3096);
and U8876 (N_8876,N_2704,N_4702);
and U8877 (N_8877,N_3459,N_4836);
or U8878 (N_8878,N_305,N_5731);
or U8879 (N_8879,N_4931,N_3425);
and U8880 (N_8880,N_1553,N_5224);
nand U8881 (N_8881,N_2892,N_1046);
nand U8882 (N_8882,N_1156,N_4784);
or U8883 (N_8883,N_5905,N_5572);
nand U8884 (N_8884,N_3485,N_381);
and U8885 (N_8885,N_3140,N_502);
and U8886 (N_8886,N_5614,N_4257);
nand U8887 (N_8887,N_5697,N_4079);
xor U8888 (N_8888,N_910,N_966);
or U8889 (N_8889,N_754,N_4839);
or U8890 (N_8890,N_5021,N_6032);
or U8891 (N_8891,N_53,N_5666);
and U8892 (N_8892,N_5911,N_3923);
or U8893 (N_8893,N_1675,N_2167);
and U8894 (N_8894,N_1794,N_5737);
or U8895 (N_8895,N_4768,N_15);
nor U8896 (N_8896,N_2835,N_4871);
nand U8897 (N_8897,N_4415,N_5439);
nor U8898 (N_8898,N_334,N_2056);
and U8899 (N_8899,N_5552,N_5765);
and U8900 (N_8900,N_2672,N_867);
or U8901 (N_8901,N_1248,N_1755);
nand U8902 (N_8902,N_5832,N_2054);
and U8903 (N_8903,N_3260,N_1792);
nor U8904 (N_8904,N_3796,N_2300);
and U8905 (N_8905,N_255,N_875);
nand U8906 (N_8906,N_4060,N_106);
nand U8907 (N_8907,N_135,N_1580);
xnor U8908 (N_8908,N_1412,N_1676);
and U8909 (N_8909,N_2770,N_3200);
or U8910 (N_8910,N_5888,N_3957);
nor U8911 (N_8911,N_1105,N_5239);
nand U8912 (N_8912,N_3795,N_2928);
and U8913 (N_8913,N_1404,N_4362);
xnor U8914 (N_8914,N_2765,N_5501);
xnor U8915 (N_8915,N_538,N_552);
nor U8916 (N_8916,N_3148,N_445);
nand U8917 (N_8917,N_1141,N_399);
nand U8918 (N_8918,N_2243,N_5094);
or U8919 (N_8919,N_3396,N_3893);
nor U8920 (N_8920,N_1036,N_5679);
nor U8921 (N_8921,N_2557,N_3069);
nor U8922 (N_8922,N_5365,N_5419);
and U8923 (N_8923,N_4995,N_784);
and U8924 (N_8924,N_3322,N_405);
or U8925 (N_8925,N_2291,N_5216);
nand U8926 (N_8926,N_389,N_2383);
nor U8927 (N_8927,N_5274,N_1816);
xnor U8928 (N_8928,N_4660,N_3483);
nand U8929 (N_8929,N_2195,N_1024);
nand U8930 (N_8930,N_2809,N_416);
and U8931 (N_8931,N_4292,N_5189);
or U8932 (N_8932,N_3135,N_375);
and U8933 (N_8933,N_4849,N_840);
or U8934 (N_8934,N_3984,N_4432);
or U8935 (N_8935,N_1158,N_5010);
nor U8936 (N_8936,N_136,N_1383);
or U8937 (N_8937,N_2793,N_3903);
nor U8938 (N_8938,N_2825,N_715);
nor U8939 (N_8939,N_256,N_2685);
or U8940 (N_8940,N_2215,N_1560);
nor U8941 (N_8941,N_5035,N_2286);
nor U8942 (N_8942,N_2218,N_4447);
nand U8943 (N_8943,N_2730,N_300);
nor U8944 (N_8944,N_5219,N_2865);
or U8945 (N_8945,N_1485,N_5570);
and U8946 (N_8946,N_2268,N_5246);
nor U8947 (N_8947,N_4161,N_4838);
and U8948 (N_8948,N_3182,N_486);
or U8949 (N_8949,N_1853,N_898);
nor U8950 (N_8950,N_4209,N_1870);
and U8951 (N_8951,N_1579,N_1571);
or U8952 (N_8952,N_5416,N_1898);
nand U8953 (N_8953,N_1773,N_1688);
nor U8954 (N_8954,N_4678,N_2706);
or U8955 (N_8955,N_3162,N_847);
xor U8956 (N_8956,N_4945,N_928);
and U8957 (N_8957,N_4235,N_747);
and U8958 (N_8958,N_2950,N_807);
and U8959 (N_8959,N_1201,N_3858);
or U8960 (N_8960,N_2270,N_4744);
nor U8961 (N_8961,N_4657,N_2995);
nor U8962 (N_8962,N_103,N_1494);
and U8963 (N_8963,N_4024,N_3132);
or U8964 (N_8964,N_4540,N_1594);
nand U8965 (N_8965,N_5412,N_561);
nand U8966 (N_8966,N_2271,N_2737);
nor U8967 (N_8967,N_1291,N_1056);
nand U8968 (N_8968,N_2973,N_1178);
nand U8969 (N_8969,N_5102,N_3302);
and U8970 (N_8970,N_5304,N_5468);
nand U8971 (N_8971,N_617,N_5872);
and U8972 (N_8972,N_6159,N_215);
nor U8973 (N_8973,N_6043,N_2235);
nor U8974 (N_8974,N_2659,N_5079);
nand U8975 (N_8975,N_1260,N_4054);
nand U8976 (N_8976,N_1346,N_3548);
or U8977 (N_8977,N_27,N_2217);
xnor U8978 (N_8978,N_5053,N_1777);
or U8979 (N_8979,N_5229,N_2513);
and U8980 (N_8980,N_394,N_2019);
and U8981 (N_8981,N_5523,N_5946);
nor U8982 (N_8982,N_4553,N_3087);
or U8983 (N_8983,N_4335,N_726);
or U8984 (N_8984,N_2430,N_864);
or U8985 (N_8985,N_5319,N_2992);
nand U8986 (N_8986,N_868,N_4542);
xor U8987 (N_8987,N_609,N_1306);
nor U8988 (N_8988,N_5781,N_6181);
or U8989 (N_8989,N_735,N_2228);
nand U8990 (N_8990,N_5649,N_5617);
and U8991 (N_8991,N_5085,N_1548);
nand U8992 (N_8992,N_41,N_846);
xor U8993 (N_8993,N_1624,N_3192);
or U8994 (N_8994,N_1166,N_4317);
nor U8995 (N_8995,N_5155,N_402);
and U8996 (N_8996,N_3072,N_1142);
or U8997 (N_8997,N_3273,N_3800);
xnor U8998 (N_8998,N_4874,N_4630);
or U8999 (N_8999,N_1803,N_4144);
nand U9000 (N_9000,N_329,N_6);
nor U9001 (N_9001,N_4492,N_217);
nor U9002 (N_9002,N_4276,N_4870);
or U9003 (N_9003,N_2302,N_2044);
and U9004 (N_9004,N_1240,N_464);
and U9005 (N_9005,N_2358,N_2634);
nor U9006 (N_9006,N_3834,N_1994);
nor U9007 (N_9007,N_3120,N_3568);
nor U9008 (N_9008,N_1174,N_4596);
and U9009 (N_9009,N_161,N_1416);
nand U9010 (N_9010,N_4759,N_308);
or U9011 (N_9011,N_1720,N_1405);
nor U9012 (N_9012,N_3677,N_102);
nand U9013 (N_9013,N_1069,N_3251);
or U9014 (N_9014,N_285,N_1852);
nand U9015 (N_9015,N_1272,N_4817);
nand U9016 (N_9016,N_5364,N_697);
or U9017 (N_9017,N_3430,N_3488);
and U9018 (N_9018,N_1473,N_3304);
and U9019 (N_9019,N_61,N_1075);
and U9020 (N_9020,N_2888,N_335);
nor U9021 (N_9021,N_2139,N_1010);
nand U9022 (N_9022,N_2734,N_6098);
nor U9023 (N_9023,N_3465,N_2193);
nor U9024 (N_9024,N_811,N_3333);
or U9025 (N_9025,N_2154,N_6129);
or U9026 (N_9026,N_5087,N_6205);
and U9027 (N_9027,N_1308,N_5694);
and U9028 (N_9028,N_628,N_2323);
or U9029 (N_9029,N_4242,N_5982);
nand U9030 (N_9030,N_5567,N_467);
or U9031 (N_9031,N_5515,N_6216);
or U9032 (N_9032,N_4998,N_4612);
nand U9033 (N_9033,N_4145,N_5562);
nand U9034 (N_9034,N_3180,N_6059);
nor U9035 (N_9035,N_5258,N_4857);
nand U9036 (N_9036,N_4374,N_3348);
nand U9037 (N_9037,N_687,N_4815);
and U9038 (N_9038,N_3020,N_567);
xnor U9039 (N_9039,N_5121,N_4098);
nor U9040 (N_9040,N_2763,N_3022);
nand U9041 (N_9041,N_577,N_2482);
or U9042 (N_9042,N_4638,N_2726);
nor U9043 (N_9043,N_11,N_4275);
nor U9044 (N_9044,N_5030,N_2007);
and U9045 (N_9045,N_72,N_1764);
and U9046 (N_9046,N_4821,N_2927);
and U9047 (N_9047,N_3571,N_6213);
nand U9048 (N_9048,N_5371,N_2535);
or U9049 (N_9049,N_1761,N_3659);
nor U9050 (N_9050,N_5983,N_4788);
nand U9051 (N_9051,N_2067,N_5415);
or U9052 (N_9052,N_4570,N_4938);
nor U9053 (N_9053,N_2420,N_5889);
nor U9054 (N_9054,N_1229,N_2137);
and U9055 (N_9055,N_4188,N_3941);
nor U9056 (N_9056,N_1711,N_4805);
xnor U9057 (N_9057,N_4265,N_4141);
or U9058 (N_9058,N_3442,N_5602);
nand U9059 (N_9059,N_5355,N_114);
xnor U9060 (N_9060,N_309,N_1335);
or U9061 (N_9061,N_1819,N_1132);
nand U9062 (N_9062,N_3589,N_5172);
or U9063 (N_9063,N_3309,N_922);
or U9064 (N_9064,N_1081,N_4130);
nor U9065 (N_9065,N_2252,N_5398);
or U9066 (N_9066,N_3888,N_2751);
or U9067 (N_9067,N_2444,N_2523);
nor U9068 (N_9068,N_4212,N_1173);
or U9069 (N_9069,N_2631,N_9);
nand U9070 (N_9070,N_6120,N_4655);
or U9071 (N_9071,N_2304,N_4407);
nor U9072 (N_9072,N_5489,N_3822);
and U9073 (N_9073,N_2448,N_3978);
or U9074 (N_9074,N_3130,N_1917);
nand U9075 (N_9075,N_5776,N_1343);
nor U9076 (N_9076,N_5841,N_5441);
and U9077 (N_9077,N_3585,N_2924);
xor U9078 (N_9078,N_6044,N_4577);
and U9079 (N_9079,N_1875,N_5728);
and U9080 (N_9080,N_4206,N_3607);
or U9081 (N_9081,N_4674,N_788);
and U9082 (N_9082,N_2810,N_4774);
nor U9083 (N_9083,N_4262,N_5680);
nor U9084 (N_9084,N_1118,N_4528);
nor U9085 (N_9085,N_2048,N_5414);
or U9086 (N_9086,N_3658,N_2985);
nor U9087 (N_9087,N_3341,N_7);
nor U9088 (N_9088,N_6221,N_1164);
nor U9089 (N_9089,N_120,N_746);
xnor U9090 (N_9090,N_187,N_3842);
and U9091 (N_9091,N_4890,N_2610);
xnor U9092 (N_9092,N_5859,N_4011);
nor U9093 (N_9093,N_3427,N_4600);
or U9094 (N_9094,N_4113,N_5891);
or U9095 (N_9095,N_2769,N_2460);
and U9096 (N_9096,N_4365,N_3832);
nor U9097 (N_9097,N_74,N_358);
and U9098 (N_9098,N_996,N_4458);
nor U9099 (N_9099,N_3670,N_834);
or U9100 (N_9100,N_2282,N_23);
nand U9101 (N_9101,N_4513,N_5245);
nand U9102 (N_9102,N_6019,N_4742);
and U9103 (N_9103,N_1406,N_3009);
nor U9104 (N_9104,N_2169,N_5115);
nand U9105 (N_9105,N_163,N_1359);
nand U9106 (N_9106,N_2804,N_1609);
and U9107 (N_9107,N_4762,N_799);
nand U9108 (N_9108,N_2085,N_4090);
and U9109 (N_9109,N_5383,N_3900);
and U9110 (N_9110,N_1834,N_1647);
xor U9111 (N_9111,N_4254,N_3646);
and U9112 (N_9112,N_2164,N_5444);
or U9113 (N_9113,N_4810,N_3828);
nand U9114 (N_9114,N_1122,N_4233);
nor U9115 (N_9115,N_3569,N_4552);
or U9116 (N_9116,N_1935,N_1465);
nor U9117 (N_9117,N_3768,N_3419);
and U9118 (N_9118,N_3489,N_6186);
nor U9119 (N_9119,N_366,N_4986);
nor U9120 (N_9120,N_4578,N_1286);
nor U9121 (N_9121,N_1419,N_2004);
or U9122 (N_9122,N_3564,N_4879);
nand U9123 (N_9123,N_1753,N_573);
nor U9124 (N_9124,N_5047,N_2258);
xor U9125 (N_9125,N_2470,N_5448);
and U9126 (N_9126,N_2657,N_4459);
and U9127 (N_9127,N_6047,N_340);
nor U9128 (N_9128,N_1070,N_539);
nor U9129 (N_9129,N_673,N_4601);
nor U9130 (N_9130,N_1058,N_1323);
xnor U9131 (N_9131,N_3987,N_1591);
or U9132 (N_9132,N_5821,N_2974);
nand U9133 (N_9133,N_4640,N_46);
nand U9134 (N_9134,N_5228,N_3159);
nand U9135 (N_9135,N_935,N_4617);
xor U9136 (N_9136,N_5403,N_5993);
nand U9137 (N_9137,N_1110,N_3989);
nor U9138 (N_9138,N_4988,N_2623);
and U9139 (N_9139,N_6007,N_2438);
nor U9140 (N_9140,N_1533,N_463);
nand U9141 (N_9141,N_2859,N_1639);
or U9142 (N_9142,N_1234,N_2656);
or U9143 (N_9143,N_4408,N_1039);
or U9144 (N_9144,N_2851,N_3242);
nor U9145 (N_9145,N_6133,N_5943);
and U9146 (N_9146,N_3237,N_1992);
and U9147 (N_9147,N_5202,N_2255);
or U9148 (N_9148,N_1387,N_1041);
or U9149 (N_9149,N_5450,N_526);
and U9150 (N_9150,N_211,N_5554);
or U9151 (N_9151,N_4089,N_4615);
and U9152 (N_9152,N_6166,N_1287);
nand U9153 (N_9153,N_3197,N_5741);
nand U9154 (N_9154,N_4929,N_5227);
nor U9155 (N_9155,N_511,N_4921);
or U9156 (N_9156,N_108,N_3423);
nor U9157 (N_9157,N_4848,N_25);
xnor U9158 (N_9158,N_4380,N_5205);
xnor U9159 (N_9159,N_22,N_3194);
nand U9160 (N_9160,N_813,N_2492);
nor U9161 (N_9161,N_1530,N_5844);
nand U9162 (N_9162,N_3165,N_6029);
nand U9163 (N_9163,N_5131,N_4448);
nor U9164 (N_9164,N_4012,N_71);
nand U9165 (N_9165,N_2777,N_2629);
nor U9166 (N_9166,N_4757,N_1705);
or U9167 (N_9167,N_2759,N_3290);
nor U9168 (N_9168,N_6046,N_3233);
or U9169 (N_9169,N_48,N_1641);
or U9170 (N_9170,N_2988,N_5553);
and U9171 (N_9171,N_6232,N_4330);
nand U9172 (N_9172,N_5382,N_1993);
and U9173 (N_9173,N_5640,N_1249);
or U9174 (N_9174,N_855,N_2305);
or U9175 (N_9175,N_62,N_3014);
nand U9176 (N_9176,N_5096,N_5969);
or U9177 (N_9177,N_4426,N_4015);
or U9178 (N_9178,N_6022,N_448);
nor U9179 (N_9179,N_2274,N_19);
or U9180 (N_9180,N_3392,N_3943);
nand U9181 (N_9181,N_5825,N_5374);
or U9182 (N_9182,N_483,N_5328);
nand U9183 (N_9183,N_6153,N_1770);
nor U9184 (N_9184,N_1163,N_659);
nand U9185 (N_9185,N_578,N_5750);
nand U9186 (N_9186,N_5185,N_3732);
nand U9187 (N_9187,N_1499,N_965);
nand U9188 (N_9188,N_3254,N_3544);
or U9189 (N_9189,N_5470,N_476);
and U9190 (N_9190,N_5743,N_5014);
nor U9191 (N_9191,N_179,N_932);
or U9192 (N_9192,N_1884,N_2241);
or U9193 (N_9193,N_2655,N_513);
nor U9194 (N_9194,N_4837,N_5651);
or U9195 (N_9195,N_2534,N_5167);
and U9196 (N_9196,N_2743,N_5808);
nor U9197 (N_9197,N_4729,N_5313);
and U9198 (N_9198,N_773,N_2900);
or U9199 (N_9199,N_2102,N_3379);
or U9200 (N_9200,N_1628,N_2819);
nor U9201 (N_9201,N_258,N_4396);
xor U9202 (N_9202,N_696,N_3279);
nor U9203 (N_9203,N_3918,N_1585);
nand U9204 (N_9204,N_2723,N_5031);
nor U9205 (N_9205,N_1047,N_5852);
or U9206 (N_9206,N_4822,N_4378);
or U9207 (N_9207,N_4875,N_2620);
and U9208 (N_9208,N_3826,N_5624);
nor U9209 (N_9209,N_172,N_5036);
nand U9210 (N_9210,N_4716,N_5517);
nand U9211 (N_9211,N_2788,N_2801);
and U9212 (N_9212,N_4138,N_1654);
xnor U9213 (N_9213,N_209,N_1361);
nand U9214 (N_9214,N_3867,N_4140);
and U9215 (N_9215,N_1427,N_2727);
nand U9216 (N_9216,N_4955,N_1043);
nor U9217 (N_9217,N_3335,N_1474);
nand U9218 (N_9218,N_3953,N_4728);
nor U9219 (N_9219,N_2548,N_2087);
and U9220 (N_9220,N_3385,N_3929);
and U9221 (N_9221,N_1210,N_1627);
nand U9222 (N_9222,N_3108,N_4289);
xor U9223 (N_9223,N_3694,N_2935);
or U9224 (N_9224,N_6227,N_1275);
nand U9225 (N_9225,N_1846,N_3777);
or U9226 (N_9226,N_5361,N_3501);
nand U9227 (N_9227,N_6149,N_4063);
and U9228 (N_9228,N_5,N_601);
xor U9229 (N_9229,N_2356,N_940);
nor U9230 (N_9230,N_1483,N_3661);
nand U9231 (N_9231,N_2242,N_3895);
xnor U9232 (N_9232,N_2970,N_5433);
nor U9233 (N_9233,N_1744,N_4240);
nand U9234 (N_9234,N_2341,N_1295);
and U9235 (N_9235,N_3288,N_5166);
and U9236 (N_9236,N_904,N_581);
or U9237 (N_9237,N_1002,N_5405);
nand U9238 (N_9238,N_1280,N_3582);
and U9239 (N_9239,N_700,N_1866);
nor U9240 (N_9240,N_1268,N_3490);
nand U9241 (N_9241,N_173,N_4554);
nand U9242 (N_9242,N_967,N_4304);
nand U9243 (N_9243,N_5158,N_2619);
or U9244 (N_9244,N_1877,N_301);
nand U9245 (N_9245,N_1528,N_3776);
nor U9246 (N_9246,N_1673,N_3526);
and U9247 (N_9247,N_5715,N_3956);
nand U9248 (N_9248,N_4112,N_1836);
nand U9249 (N_9249,N_1658,N_1837);
nand U9250 (N_9250,N_505,N_5707);
and U9251 (N_9251,N_2567,N_3863);
xnor U9252 (N_9252,N_1735,N_2423);
nand U9253 (N_9253,N_1428,N_2815);
nand U9254 (N_9254,N_3498,N_4334);
or U9255 (N_9255,N_4475,N_5380);
nand U9256 (N_9256,N_611,N_2504);
or U9257 (N_9257,N_3683,N_3844);
and U9258 (N_9258,N_5724,N_5238);
nand U9259 (N_9259,N_3499,N_3438);
and U9260 (N_9260,N_2310,N_4771);
nor U9261 (N_9261,N_307,N_2705);
or U9262 (N_9262,N_4719,N_703);
nand U9263 (N_9263,N_6207,N_4818);
or U9264 (N_9264,N_4290,N_812);
nand U9265 (N_9265,N_1059,N_3679);
nor U9266 (N_9266,N_4103,N_134);
or U9267 (N_9267,N_948,N_5292);
and U9268 (N_9268,N_5792,N_1934);
nor U9269 (N_9269,N_2625,N_3959);
nand U9270 (N_9270,N_3247,N_2312);
nor U9271 (N_9271,N_4847,N_5513);
nor U9272 (N_9272,N_4727,N_3527);
xor U9273 (N_9273,N_183,N_4977);
and U9274 (N_9274,N_4877,N_2017);
nand U9275 (N_9275,N_3207,N_6249);
xnor U9276 (N_9276,N_5550,N_1266);
or U9277 (N_9277,N_1668,N_3846);
nor U9278 (N_9278,N_2699,N_6023);
nand U9279 (N_9279,N_34,N_6119);
or U9280 (N_9280,N_198,N_3561);
nand U9281 (N_9281,N_4286,N_3370);
or U9282 (N_9282,N_2877,N_1987);
or U9283 (N_9283,N_2573,N_5719);
and U9284 (N_9284,N_3534,N_3271);
nand U9285 (N_9285,N_2468,N_5830);
xnor U9286 (N_9286,N_3231,N_1424);
xnor U9287 (N_9287,N_3712,N_4803);
or U9288 (N_9288,N_3403,N_3673);
nand U9289 (N_9289,N_383,N_899);
and U9290 (N_9290,N_1843,N_5488);
nand U9291 (N_9291,N_2639,N_4677);
nor U9292 (N_9292,N_1613,N_6089);
or U9293 (N_9293,N_4471,N_470);
nor U9294 (N_9294,N_298,N_5987);
nand U9295 (N_9295,N_3996,N_1648);
or U9296 (N_9296,N_3376,N_2100);
nand U9297 (N_9297,N_1972,N_4804);
nand U9298 (N_9298,N_5271,N_5265);
nand U9299 (N_9299,N_4511,N_1289);
nand U9300 (N_9300,N_1878,N_4587);
nor U9301 (N_9301,N_1599,N_5022);
and U9302 (N_9302,N_3622,N_5483);
or U9303 (N_9303,N_2836,N_1662);
or U9304 (N_9304,N_4351,N_5099);
and U9305 (N_9305,N_89,N_322);
xnor U9306 (N_9306,N_2738,N_1477);
nand U9307 (N_9307,N_514,N_667);
nor U9308 (N_9308,N_185,N_3647);
or U9309 (N_9309,N_4005,N_5773);
nand U9310 (N_9310,N_4349,N_6172);
nand U9311 (N_9311,N_1696,N_522);
or U9312 (N_9312,N_6192,N_3769);
and U9313 (N_9313,N_2165,N_1443);
or U9314 (N_9314,N_118,N_3804);
nand U9315 (N_9315,N_4620,N_5838);
nor U9316 (N_9316,N_3289,N_3805);
and U9317 (N_9317,N_1888,N_13);
nor U9318 (N_9318,N_3224,N_397);
nor U9319 (N_9319,N_2134,N_4449);
or U9320 (N_9320,N_3077,N_6231);
or U9321 (N_9321,N_5165,N_5000);
xnor U9322 (N_9322,N_5534,N_5592);
nand U9323 (N_9323,N_5397,N_1239);
or U9324 (N_9324,N_500,N_1097);
nor U9325 (N_9325,N_4503,N_1066);
nor U9326 (N_9326,N_4083,N_5853);
nand U9327 (N_9327,N_3487,N_3476);
or U9328 (N_9328,N_758,N_5848);
and U9329 (N_9329,N_4126,N_1146);
nor U9330 (N_9330,N_1064,N_4642);
xor U9331 (N_9331,N_3007,N_2016);
xnor U9332 (N_9332,N_2322,N_2676);
nor U9333 (N_9333,N_1211,N_2688);
and U9334 (N_9334,N_4594,N_6113);
nand U9335 (N_9335,N_4556,N_4457);
or U9336 (N_9336,N_1549,N_4217);
or U9337 (N_9337,N_5620,N_1913);
or U9338 (N_9338,N_4714,N_1212);
nand U9339 (N_9339,N_1050,N_3295);
or U9340 (N_9340,N_5314,N_4948);
nand U9341 (N_9341,N_2175,N_2428);
and U9342 (N_9342,N_6041,N_791);
and U9343 (N_9343,N_1738,N_4146);
nand U9344 (N_9344,N_4704,N_2027);
nor U9345 (N_9345,N_1970,N_3091);
nor U9346 (N_9346,N_5608,N_877);
and U9347 (N_9347,N_862,N_5699);
or U9348 (N_9348,N_1379,N_4915);
or U9349 (N_9349,N_406,N_5389);
xnor U9350 (N_9350,N_2360,N_4446);
or U9351 (N_9351,N_37,N_1909);
nor U9352 (N_9352,N_2278,N_2080);
xor U9353 (N_9353,N_1723,N_1625);
nand U9354 (N_9354,N_6158,N_3736);
and U9355 (N_9355,N_1083,N_6191);
and U9356 (N_9356,N_5126,N_2202);
xnor U9357 (N_9357,N_3323,N_873);
nand U9358 (N_9358,N_4433,N_5896);
nor U9359 (N_9359,N_5967,N_4320);
and U9360 (N_9360,N_139,N_3599);
nand U9361 (N_9361,N_4799,N_1561);
nor U9362 (N_9362,N_398,N_1035);
xor U9363 (N_9363,N_2565,N_1537);
or U9364 (N_9364,N_6122,N_4981);
or U9365 (N_9365,N_4208,N_1737);
nor U9366 (N_9366,N_3201,N_5717);
or U9367 (N_9367,N_1433,N_2684);
or U9368 (N_9368,N_221,N_4730);
and U9369 (N_9369,N_156,N_4394);
xnor U9370 (N_9370,N_1495,N_5464);
and U9371 (N_9371,N_751,N_2725);
and U9372 (N_9372,N_1710,N_141);
xnor U9373 (N_9373,N_3985,N_4215);
and U9374 (N_9374,N_1182,N_5279);
or U9375 (N_9375,N_4382,N_5665);
or U9376 (N_9376,N_2299,N_1292);
nand U9377 (N_9377,N_6071,N_1720);
nand U9378 (N_9378,N_1897,N_1510);
and U9379 (N_9379,N_4585,N_4165);
and U9380 (N_9380,N_1286,N_836);
and U9381 (N_9381,N_6225,N_704);
xor U9382 (N_9382,N_4895,N_3320);
and U9383 (N_9383,N_5553,N_339);
or U9384 (N_9384,N_337,N_5303);
nand U9385 (N_9385,N_4969,N_3999);
xor U9386 (N_9386,N_5335,N_3187);
nor U9387 (N_9387,N_5244,N_2076);
or U9388 (N_9388,N_1698,N_384);
or U9389 (N_9389,N_4185,N_1077);
or U9390 (N_9390,N_6122,N_3826);
nand U9391 (N_9391,N_1228,N_2955);
or U9392 (N_9392,N_4809,N_3217);
nor U9393 (N_9393,N_3138,N_2665);
or U9394 (N_9394,N_3286,N_3435);
nor U9395 (N_9395,N_6068,N_5621);
nor U9396 (N_9396,N_1328,N_6224);
nand U9397 (N_9397,N_5448,N_1805);
nand U9398 (N_9398,N_3460,N_3803);
and U9399 (N_9399,N_4410,N_4976);
nor U9400 (N_9400,N_4724,N_752);
and U9401 (N_9401,N_3800,N_4783);
nor U9402 (N_9402,N_1920,N_2289);
nand U9403 (N_9403,N_4212,N_5455);
or U9404 (N_9404,N_1793,N_5779);
or U9405 (N_9405,N_4634,N_647);
nand U9406 (N_9406,N_408,N_3917);
or U9407 (N_9407,N_1863,N_3113);
nand U9408 (N_9408,N_6065,N_4106);
nor U9409 (N_9409,N_776,N_3859);
and U9410 (N_9410,N_2250,N_3634);
nor U9411 (N_9411,N_3395,N_2937);
nor U9412 (N_9412,N_2087,N_973);
nand U9413 (N_9413,N_4330,N_3741);
and U9414 (N_9414,N_954,N_3238);
or U9415 (N_9415,N_5069,N_3066);
and U9416 (N_9416,N_3103,N_2072);
nand U9417 (N_9417,N_555,N_367);
nor U9418 (N_9418,N_31,N_3966);
xor U9419 (N_9419,N_5611,N_1856);
or U9420 (N_9420,N_394,N_1932);
nand U9421 (N_9421,N_1901,N_2457);
nand U9422 (N_9422,N_4697,N_2967);
nor U9423 (N_9423,N_1980,N_441);
nand U9424 (N_9424,N_4374,N_3899);
nand U9425 (N_9425,N_1055,N_3619);
and U9426 (N_9426,N_3871,N_4921);
nor U9427 (N_9427,N_5670,N_2339);
and U9428 (N_9428,N_2336,N_5594);
nand U9429 (N_9429,N_2229,N_4143);
xor U9430 (N_9430,N_249,N_2187);
or U9431 (N_9431,N_4702,N_2587);
or U9432 (N_9432,N_1558,N_4926);
and U9433 (N_9433,N_3805,N_2898);
nand U9434 (N_9434,N_6185,N_971);
nor U9435 (N_9435,N_4925,N_277);
or U9436 (N_9436,N_4262,N_2575);
nand U9437 (N_9437,N_460,N_2535);
nor U9438 (N_9438,N_1266,N_30);
nand U9439 (N_9439,N_5228,N_985);
and U9440 (N_9440,N_1126,N_3051);
and U9441 (N_9441,N_1390,N_353);
nand U9442 (N_9442,N_520,N_4167);
nand U9443 (N_9443,N_2049,N_1865);
or U9444 (N_9444,N_695,N_2782);
and U9445 (N_9445,N_3063,N_354);
nor U9446 (N_9446,N_1179,N_2912);
and U9447 (N_9447,N_5651,N_2132);
nand U9448 (N_9448,N_3512,N_2909);
nand U9449 (N_9449,N_3879,N_2999);
or U9450 (N_9450,N_4146,N_1857);
or U9451 (N_9451,N_2099,N_850);
xor U9452 (N_9452,N_2645,N_1244);
or U9453 (N_9453,N_3423,N_3470);
or U9454 (N_9454,N_3034,N_5184);
nor U9455 (N_9455,N_3286,N_807);
and U9456 (N_9456,N_3187,N_2663);
nand U9457 (N_9457,N_3595,N_5207);
or U9458 (N_9458,N_1658,N_4342);
and U9459 (N_9459,N_5415,N_2805);
nand U9460 (N_9460,N_5564,N_3886);
or U9461 (N_9461,N_2467,N_2840);
and U9462 (N_9462,N_54,N_1933);
or U9463 (N_9463,N_2679,N_5709);
nand U9464 (N_9464,N_5219,N_135);
xor U9465 (N_9465,N_3142,N_754);
or U9466 (N_9466,N_3490,N_6021);
nand U9467 (N_9467,N_3807,N_482);
nor U9468 (N_9468,N_4494,N_3247);
nand U9469 (N_9469,N_5297,N_3508);
xor U9470 (N_9470,N_2262,N_3245);
xnor U9471 (N_9471,N_1409,N_5571);
nor U9472 (N_9472,N_5361,N_1190);
or U9473 (N_9473,N_4500,N_1293);
or U9474 (N_9474,N_1713,N_5592);
nor U9475 (N_9475,N_3957,N_284);
or U9476 (N_9476,N_5402,N_4805);
nand U9477 (N_9477,N_1626,N_435);
nand U9478 (N_9478,N_4604,N_2909);
xnor U9479 (N_9479,N_3183,N_4874);
nor U9480 (N_9480,N_3350,N_121);
and U9481 (N_9481,N_4391,N_4951);
or U9482 (N_9482,N_3636,N_5712);
or U9483 (N_9483,N_5954,N_2079);
or U9484 (N_9484,N_3049,N_4420);
and U9485 (N_9485,N_2311,N_4325);
xor U9486 (N_9486,N_522,N_2663);
nand U9487 (N_9487,N_3397,N_4199);
nand U9488 (N_9488,N_62,N_1586);
or U9489 (N_9489,N_1164,N_2799);
or U9490 (N_9490,N_2979,N_709);
nor U9491 (N_9491,N_2288,N_1164);
xnor U9492 (N_9492,N_2985,N_3984);
or U9493 (N_9493,N_2997,N_3947);
and U9494 (N_9494,N_2648,N_695);
or U9495 (N_9495,N_5201,N_460);
nor U9496 (N_9496,N_2724,N_772);
and U9497 (N_9497,N_635,N_491);
or U9498 (N_9498,N_5375,N_2880);
nor U9499 (N_9499,N_5532,N_835);
nand U9500 (N_9500,N_888,N_1247);
nand U9501 (N_9501,N_2118,N_2769);
nor U9502 (N_9502,N_1797,N_5236);
nand U9503 (N_9503,N_3258,N_1483);
or U9504 (N_9504,N_2421,N_2649);
xnor U9505 (N_9505,N_4826,N_4191);
or U9506 (N_9506,N_5310,N_2188);
or U9507 (N_9507,N_1530,N_1236);
and U9508 (N_9508,N_5619,N_478);
xor U9509 (N_9509,N_1939,N_3543);
or U9510 (N_9510,N_4657,N_2407);
nor U9511 (N_9511,N_5900,N_5771);
and U9512 (N_9512,N_3043,N_3122);
and U9513 (N_9513,N_1325,N_593);
nor U9514 (N_9514,N_3268,N_2482);
nor U9515 (N_9515,N_3787,N_1251);
nand U9516 (N_9516,N_550,N_2510);
xnor U9517 (N_9517,N_3887,N_4839);
or U9518 (N_9518,N_1606,N_1660);
nor U9519 (N_9519,N_5918,N_1796);
or U9520 (N_9520,N_5721,N_4676);
nor U9521 (N_9521,N_4981,N_4257);
or U9522 (N_9522,N_4584,N_2108);
or U9523 (N_9523,N_1957,N_4199);
and U9524 (N_9524,N_4480,N_4350);
or U9525 (N_9525,N_285,N_5408);
or U9526 (N_9526,N_4935,N_201);
and U9527 (N_9527,N_5979,N_3588);
and U9528 (N_9528,N_2489,N_4680);
nor U9529 (N_9529,N_4485,N_3194);
nand U9530 (N_9530,N_1014,N_763);
or U9531 (N_9531,N_5214,N_1048);
and U9532 (N_9532,N_2742,N_333);
and U9533 (N_9533,N_3032,N_1527);
and U9534 (N_9534,N_1893,N_2603);
and U9535 (N_9535,N_1312,N_476);
nor U9536 (N_9536,N_2305,N_3238);
xnor U9537 (N_9537,N_3733,N_3185);
nand U9538 (N_9538,N_850,N_3183);
or U9539 (N_9539,N_2424,N_1835);
or U9540 (N_9540,N_293,N_3327);
and U9541 (N_9541,N_2065,N_3775);
and U9542 (N_9542,N_3042,N_4576);
xor U9543 (N_9543,N_2278,N_2745);
nor U9544 (N_9544,N_3726,N_5108);
nand U9545 (N_9545,N_4727,N_1601);
nand U9546 (N_9546,N_1936,N_2709);
nand U9547 (N_9547,N_3486,N_3197);
or U9548 (N_9548,N_652,N_3253);
and U9549 (N_9549,N_5382,N_3561);
nor U9550 (N_9550,N_2324,N_1506);
xor U9551 (N_9551,N_641,N_5100);
or U9552 (N_9552,N_2294,N_3737);
nand U9553 (N_9553,N_1205,N_2862);
nor U9554 (N_9554,N_3807,N_3924);
nand U9555 (N_9555,N_6223,N_5923);
nor U9556 (N_9556,N_5511,N_4658);
xnor U9557 (N_9557,N_3678,N_1441);
or U9558 (N_9558,N_1911,N_6115);
and U9559 (N_9559,N_4526,N_5132);
or U9560 (N_9560,N_262,N_1345);
or U9561 (N_9561,N_115,N_2004);
or U9562 (N_9562,N_1833,N_3826);
nor U9563 (N_9563,N_3053,N_5909);
or U9564 (N_9564,N_3696,N_877);
or U9565 (N_9565,N_2553,N_5039);
nand U9566 (N_9566,N_5643,N_5306);
nor U9567 (N_9567,N_1320,N_1335);
nor U9568 (N_9568,N_2936,N_2172);
and U9569 (N_9569,N_875,N_3988);
or U9570 (N_9570,N_144,N_5735);
nor U9571 (N_9571,N_3836,N_533);
nor U9572 (N_9572,N_1958,N_2224);
nor U9573 (N_9573,N_452,N_1549);
nand U9574 (N_9574,N_2541,N_3705);
xor U9575 (N_9575,N_2821,N_5762);
or U9576 (N_9576,N_5027,N_104);
and U9577 (N_9577,N_3926,N_4971);
and U9578 (N_9578,N_3772,N_5520);
xnor U9579 (N_9579,N_2311,N_445);
xor U9580 (N_9580,N_1640,N_1103);
nor U9581 (N_9581,N_5380,N_5624);
nor U9582 (N_9582,N_170,N_1393);
nand U9583 (N_9583,N_3503,N_4043);
or U9584 (N_9584,N_5917,N_3604);
or U9585 (N_9585,N_1247,N_6009);
or U9586 (N_9586,N_5773,N_4440);
xor U9587 (N_9587,N_3644,N_1765);
nor U9588 (N_9588,N_3621,N_5640);
or U9589 (N_9589,N_5595,N_4275);
nand U9590 (N_9590,N_2840,N_5256);
xnor U9591 (N_9591,N_598,N_5130);
or U9592 (N_9592,N_4815,N_5063);
nand U9593 (N_9593,N_288,N_735);
or U9594 (N_9594,N_2114,N_5809);
nand U9595 (N_9595,N_3188,N_2243);
nor U9596 (N_9596,N_5031,N_5037);
xor U9597 (N_9597,N_4698,N_5603);
or U9598 (N_9598,N_2993,N_6104);
nand U9599 (N_9599,N_4727,N_134);
or U9600 (N_9600,N_125,N_575);
nand U9601 (N_9601,N_899,N_1951);
nor U9602 (N_9602,N_3812,N_4134);
or U9603 (N_9603,N_4499,N_3874);
or U9604 (N_9604,N_1075,N_1733);
or U9605 (N_9605,N_4748,N_633);
or U9606 (N_9606,N_5013,N_1581);
and U9607 (N_9607,N_3754,N_4405);
and U9608 (N_9608,N_2058,N_849);
nor U9609 (N_9609,N_3159,N_5754);
xnor U9610 (N_9610,N_3773,N_3373);
nand U9611 (N_9611,N_4184,N_1281);
nand U9612 (N_9612,N_1026,N_371);
and U9613 (N_9613,N_5119,N_84);
or U9614 (N_9614,N_1402,N_2453);
or U9615 (N_9615,N_6058,N_5155);
nor U9616 (N_9616,N_540,N_2527);
nand U9617 (N_9617,N_542,N_6180);
nand U9618 (N_9618,N_1240,N_3101);
xor U9619 (N_9619,N_4038,N_2723);
nand U9620 (N_9620,N_3826,N_3947);
or U9621 (N_9621,N_278,N_1172);
nor U9622 (N_9622,N_3912,N_1398);
nor U9623 (N_9623,N_2879,N_3806);
nor U9624 (N_9624,N_2355,N_1606);
and U9625 (N_9625,N_1902,N_6170);
or U9626 (N_9626,N_3759,N_1993);
and U9627 (N_9627,N_2785,N_2337);
or U9628 (N_9628,N_2363,N_2132);
or U9629 (N_9629,N_3216,N_4878);
nor U9630 (N_9630,N_632,N_2305);
nor U9631 (N_9631,N_2219,N_3028);
xor U9632 (N_9632,N_584,N_162);
and U9633 (N_9633,N_1928,N_1251);
nor U9634 (N_9634,N_1223,N_758);
or U9635 (N_9635,N_5054,N_4997);
nor U9636 (N_9636,N_5658,N_3228);
or U9637 (N_9637,N_5846,N_6246);
or U9638 (N_9638,N_421,N_4715);
xnor U9639 (N_9639,N_5762,N_5576);
or U9640 (N_9640,N_2503,N_3982);
nand U9641 (N_9641,N_285,N_3396);
nand U9642 (N_9642,N_2816,N_588);
nand U9643 (N_9643,N_4346,N_4363);
or U9644 (N_9644,N_818,N_2111);
and U9645 (N_9645,N_3902,N_5047);
nor U9646 (N_9646,N_5205,N_5870);
or U9647 (N_9647,N_6025,N_1249);
or U9648 (N_9648,N_5151,N_4652);
nor U9649 (N_9649,N_5296,N_4770);
nor U9650 (N_9650,N_2139,N_5375);
nor U9651 (N_9651,N_2897,N_3393);
nand U9652 (N_9652,N_5144,N_1947);
xnor U9653 (N_9653,N_4820,N_3301);
or U9654 (N_9654,N_1901,N_891);
nand U9655 (N_9655,N_2844,N_527);
nor U9656 (N_9656,N_2076,N_107);
nand U9657 (N_9657,N_4552,N_458);
nand U9658 (N_9658,N_1473,N_3877);
xnor U9659 (N_9659,N_4112,N_6076);
xor U9660 (N_9660,N_5580,N_3994);
and U9661 (N_9661,N_880,N_2184);
or U9662 (N_9662,N_2279,N_5051);
nor U9663 (N_9663,N_2634,N_5453);
and U9664 (N_9664,N_3537,N_2161);
or U9665 (N_9665,N_3771,N_3614);
and U9666 (N_9666,N_3294,N_3344);
and U9667 (N_9667,N_3235,N_5521);
xnor U9668 (N_9668,N_2667,N_3071);
or U9669 (N_9669,N_5418,N_503);
and U9670 (N_9670,N_5398,N_4300);
or U9671 (N_9671,N_3635,N_4556);
and U9672 (N_9672,N_1721,N_3388);
nor U9673 (N_9673,N_149,N_5190);
and U9674 (N_9674,N_4134,N_4225);
nand U9675 (N_9675,N_741,N_5026);
or U9676 (N_9676,N_1816,N_1624);
nand U9677 (N_9677,N_4754,N_3233);
or U9678 (N_9678,N_4125,N_3185);
and U9679 (N_9679,N_748,N_3425);
xor U9680 (N_9680,N_935,N_848);
nor U9681 (N_9681,N_6132,N_2781);
nand U9682 (N_9682,N_1996,N_3295);
or U9683 (N_9683,N_3542,N_2203);
xnor U9684 (N_9684,N_2622,N_1712);
nand U9685 (N_9685,N_4093,N_4543);
or U9686 (N_9686,N_1077,N_3276);
or U9687 (N_9687,N_4067,N_3431);
nand U9688 (N_9688,N_3034,N_4668);
or U9689 (N_9689,N_3003,N_309);
or U9690 (N_9690,N_217,N_495);
nor U9691 (N_9691,N_456,N_5050);
nand U9692 (N_9692,N_5763,N_580);
xor U9693 (N_9693,N_2154,N_4852);
and U9694 (N_9694,N_2917,N_3574);
nand U9695 (N_9695,N_5070,N_5310);
and U9696 (N_9696,N_2565,N_2060);
and U9697 (N_9697,N_5250,N_712);
nand U9698 (N_9698,N_3974,N_2174);
xnor U9699 (N_9699,N_1331,N_5770);
and U9700 (N_9700,N_4690,N_5566);
nand U9701 (N_9701,N_6226,N_590);
nor U9702 (N_9702,N_2586,N_5507);
and U9703 (N_9703,N_4729,N_2731);
and U9704 (N_9704,N_4908,N_185);
nand U9705 (N_9705,N_1398,N_214);
nand U9706 (N_9706,N_1505,N_5461);
nand U9707 (N_9707,N_2869,N_2412);
or U9708 (N_9708,N_4454,N_4883);
nand U9709 (N_9709,N_5307,N_2927);
nor U9710 (N_9710,N_723,N_2876);
and U9711 (N_9711,N_2253,N_2420);
and U9712 (N_9712,N_5157,N_6142);
and U9713 (N_9713,N_3489,N_5205);
and U9714 (N_9714,N_3846,N_5094);
and U9715 (N_9715,N_1973,N_2776);
nor U9716 (N_9716,N_6100,N_4934);
xor U9717 (N_9717,N_5945,N_145);
and U9718 (N_9718,N_5483,N_1431);
and U9719 (N_9719,N_4379,N_2188);
nand U9720 (N_9720,N_2114,N_5102);
nand U9721 (N_9721,N_4273,N_6227);
xor U9722 (N_9722,N_3755,N_3044);
nor U9723 (N_9723,N_6186,N_4639);
nand U9724 (N_9724,N_192,N_2621);
nor U9725 (N_9725,N_5780,N_1808);
and U9726 (N_9726,N_4521,N_753);
or U9727 (N_9727,N_1175,N_1492);
or U9728 (N_9728,N_5889,N_363);
and U9729 (N_9729,N_4837,N_2450);
and U9730 (N_9730,N_4769,N_61);
xor U9731 (N_9731,N_4811,N_4201);
and U9732 (N_9732,N_315,N_3291);
xnor U9733 (N_9733,N_212,N_803);
or U9734 (N_9734,N_5611,N_3622);
nand U9735 (N_9735,N_1691,N_3171);
and U9736 (N_9736,N_2345,N_2294);
nor U9737 (N_9737,N_536,N_3542);
nand U9738 (N_9738,N_6062,N_3894);
xnor U9739 (N_9739,N_1693,N_338);
nand U9740 (N_9740,N_1816,N_3003);
nor U9741 (N_9741,N_5285,N_6070);
nand U9742 (N_9742,N_712,N_659);
nand U9743 (N_9743,N_5867,N_2992);
and U9744 (N_9744,N_5563,N_2020);
nor U9745 (N_9745,N_3183,N_3823);
nand U9746 (N_9746,N_4614,N_5764);
and U9747 (N_9747,N_479,N_5612);
or U9748 (N_9748,N_2542,N_2437);
or U9749 (N_9749,N_1738,N_4620);
nor U9750 (N_9750,N_5015,N_6088);
nor U9751 (N_9751,N_1,N_4887);
nor U9752 (N_9752,N_3994,N_600);
nand U9753 (N_9753,N_4871,N_2873);
or U9754 (N_9754,N_85,N_534);
xor U9755 (N_9755,N_5297,N_6226);
and U9756 (N_9756,N_124,N_2698);
nand U9757 (N_9757,N_4223,N_3316);
xor U9758 (N_9758,N_1822,N_1376);
or U9759 (N_9759,N_2335,N_3101);
or U9760 (N_9760,N_5540,N_278);
and U9761 (N_9761,N_2309,N_3148);
and U9762 (N_9762,N_6118,N_3905);
and U9763 (N_9763,N_1234,N_4512);
xnor U9764 (N_9764,N_1716,N_5509);
nand U9765 (N_9765,N_3526,N_3060);
nand U9766 (N_9766,N_4172,N_1583);
or U9767 (N_9767,N_2617,N_3800);
or U9768 (N_9768,N_2698,N_1546);
and U9769 (N_9769,N_6181,N_435);
or U9770 (N_9770,N_5002,N_5727);
and U9771 (N_9771,N_2071,N_4827);
xnor U9772 (N_9772,N_5878,N_2550);
nand U9773 (N_9773,N_346,N_2359);
xnor U9774 (N_9774,N_5049,N_4603);
nand U9775 (N_9775,N_1059,N_2052);
xor U9776 (N_9776,N_2810,N_4627);
or U9777 (N_9777,N_3698,N_846);
xnor U9778 (N_9778,N_5327,N_4367);
and U9779 (N_9779,N_2836,N_5436);
and U9780 (N_9780,N_6159,N_1840);
and U9781 (N_9781,N_4716,N_3573);
nor U9782 (N_9782,N_2155,N_5093);
nand U9783 (N_9783,N_2801,N_5531);
or U9784 (N_9784,N_2155,N_1568);
or U9785 (N_9785,N_3153,N_6170);
xor U9786 (N_9786,N_4303,N_1417);
or U9787 (N_9787,N_1828,N_1543);
nand U9788 (N_9788,N_5407,N_3494);
or U9789 (N_9789,N_2508,N_3637);
nor U9790 (N_9790,N_599,N_3195);
and U9791 (N_9791,N_4350,N_2308);
or U9792 (N_9792,N_2852,N_1036);
and U9793 (N_9793,N_1345,N_4051);
and U9794 (N_9794,N_4996,N_43);
nand U9795 (N_9795,N_188,N_755);
nand U9796 (N_9796,N_4170,N_77);
and U9797 (N_9797,N_499,N_2710);
nor U9798 (N_9798,N_6104,N_4062);
or U9799 (N_9799,N_5085,N_3885);
and U9800 (N_9800,N_2258,N_455);
nand U9801 (N_9801,N_1711,N_1258);
nor U9802 (N_9802,N_3196,N_3367);
and U9803 (N_9803,N_2905,N_1467);
xor U9804 (N_9804,N_1019,N_1199);
nor U9805 (N_9805,N_4889,N_3697);
nand U9806 (N_9806,N_1006,N_376);
or U9807 (N_9807,N_1174,N_994);
or U9808 (N_9808,N_1254,N_2681);
and U9809 (N_9809,N_5220,N_1949);
xnor U9810 (N_9810,N_4415,N_4817);
nand U9811 (N_9811,N_2161,N_1220);
and U9812 (N_9812,N_3447,N_2424);
and U9813 (N_9813,N_1585,N_4291);
and U9814 (N_9814,N_4600,N_4328);
nor U9815 (N_9815,N_408,N_2157);
nand U9816 (N_9816,N_4818,N_642);
and U9817 (N_9817,N_5681,N_478);
nor U9818 (N_9818,N_60,N_3447);
and U9819 (N_9819,N_2700,N_5631);
and U9820 (N_9820,N_3907,N_2392);
nor U9821 (N_9821,N_6132,N_4919);
nor U9822 (N_9822,N_2369,N_5256);
nor U9823 (N_9823,N_260,N_1450);
or U9824 (N_9824,N_1096,N_234);
nand U9825 (N_9825,N_4690,N_1974);
nor U9826 (N_9826,N_6247,N_3818);
nand U9827 (N_9827,N_5028,N_3851);
nand U9828 (N_9828,N_2725,N_3858);
nor U9829 (N_9829,N_5925,N_6167);
and U9830 (N_9830,N_549,N_1625);
xor U9831 (N_9831,N_2237,N_981);
nand U9832 (N_9832,N_2094,N_3508);
and U9833 (N_9833,N_3544,N_5800);
and U9834 (N_9834,N_1164,N_2736);
and U9835 (N_9835,N_2369,N_5538);
or U9836 (N_9836,N_172,N_1060);
nor U9837 (N_9837,N_3518,N_6179);
nor U9838 (N_9838,N_4586,N_2293);
and U9839 (N_9839,N_6141,N_348);
nand U9840 (N_9840,N_2152,N_2337);
and U9841 (N_9841,N_2431,N_738);
nor U9842 (N_9842,N_529,N_2391);
nor U9843 (N_9843,N_1253,N_818);
or U9844 (N_9844,N_3380,N_780);
and U9845 (N_9845,N_5264,N_4863);
xnor U9846 (N_9846,N_763,N_2987);
nand U9847 (N_9847,N_3995,N_2086);
and U9848 (N_9848,N_735,N_4122);
xor U9849 (N_9849,N_4455,N_2411);
nand U9850 (N_9850,N_4298,N_1113);
nand U9851 (N_9851,N_72,N_3274);
nor U9852 (N_9852,N_4073,N_2809);
nor U9853 (N_9853,N_697,N_5548);
or U9854 (N_9854,N_1790,N_248);
nor U9855 (N_9855,N_3999,N_2520);
nor U9856 (N_9856,N_773,N_3745);
nand U9857 (N_9857,N_6136,N_4331);
nand U9858 (N_9858,N_4389,N_4398);
and U9859 (N_9859,N_2264,N_1395);
nor U9860 (N_9860,N_3586,N_6072);
or U9861 (N_9861,N_1618,N_212);
nor U9862 (N_9862,N_3141,N_1695);
or U9863 (N_9863,N_4403,N_4780);
nor U9864 (N_9864,N_2959,N_2684);
and U9865 (N_9865,N_1750,N_4842);
xor U9866 (N_9866,N_5700,N_3854);
nand U9867 (N_9867,N_4302,N_5048);
nor U9868 (N_9868,N_4841,N_991);
or U9869 (N_9869,N_2730,N_1686);
nor U9870 (N_9870,N_3855,N_178);
xor U9871 (N_9871,N_5700,N_2037);
or U9872 (N_9872,N_4075,N_2068);
nor U9873 (N_9873,N_4609,N_2665);
nand U9874 (N_9874,N_5682,N_5245);
nand U9875 (N_9875,N_4059,N_2402);
nand U9876 (N_9876,N_2080,N_1722);
and U9877 (N_9877,N_5591,N_239);
nand U9878 (N_9878,N_3608,N_25);
nor U9879 (N_9879,N_1232,N_5769);
or U9880 (N_9880,N_2428,N_520);
nor U9881 (N_9881,N_5580,N_3101);
and U9882 (N_9882,N_5311,N_2686);
and U9883 (N_9883,N_4556,N_637);
nand U9884 (N_9884,N_2730,N_5774);
and U9885 (N_9885,N_3747,N_823);
or U9886 (N_9886,N_1420,N_2884);
and U9887 (N_9887,N_268,N_2530);
nand U9888 (N_9888,N_1669,N_4238);
nor U9889 (N_9889,N_3806,N_135);
nor U9890 (N_9890,N_583,N_4036);
or U9891 (N_9891,N_5809,N_4900);
nand U9892 (N_9892,N_2276,N_4283);
nand U9893 (N_9893,N_1137,N_1974);
xnor U9894 (N_9894,N_3050,N_6218);
nor U9895 (N_9895,N_4984,N_5655);
and U9896 (N_9896,N_2159,N_3897);
nand U9897 (N_9897,N_5307,N_3472);
xor U9898 (N_9898,N_129,N_2417);
nand U9899 (N_9899,N_128,N_2645);
and U9900 (N_9900,N_1665,N_4337);
or U9901 (N_9901,N_2883,N_3437);
nor U9902 (N_9902,N_697,N_2333);
and U9903 (N_9903,N_5672,N_4266);
nand U9904 (N_9904,N_5459,N_417);
and U9905 (N_9905,N_3199,N_5417);
nand U9906 (N_9906,N_3228,N_5650);
nand U9907 (N_9907,N_5602,N_1071);
nand U9908 (N_9908,N_1282,N_1929);
nor U9909 (N_9909,N_3752,N_5835);
xnor U9910 (N_9910,N_5982,N_354);
nor U9911 (N_9911,N_4713,N_4726);
nor U9912 (N_9912,N_153,N_4327);
and U9913 (N_9913,N_1554,N_654);
nand U9914 (N_9914,N_741,N_1289);
xor U9915 (N_9915,N_2914,N_5341);
or U9916 (N_9916,N_4608,N_1805);
nand U9917 (N_9917,N_1827,N_4067);
nor U9918 (N_9918,N_2265,N_481);
nor U9919 (N_9919,N_3825,N_5866);
and U9920 (N_9920,N_559,N_1029);
nand U9921 (N_9921,N_94,N_3051);
and U9922 (N_9922,N_4196,N_5972);
and U9923 (N_9923,N_5919,N_1766);
nor U9924 (N_9924,N_102,N_3212);
and U9925 (N_9925,N_859,N_4911);
nand U9926 (N_9926,N_5295,N_3522);
xor U9927 (N_9927,N_5635,N_1922);
nor U9928 (N_9928,N_1718,N_4381);
nor U9929 (N_9929,N_2190,N_3291);
or U9930 (N_9930,N_777,N_3636);
nand U9931 (N_9931,N_3650,N_5804);
nor U9932 (N_9932,N_5281,N_1049);
or U9933 (N_9933,N_4842,N_4424);
or U9934 (N_9934,N_4100,N_4415);
nand U9935 (N_9935,N_3786,N_1704);
nor U9936 (N_9936,N_2196,N_1729);
or U9937 (N_9937,N_4038,N_4803);
nor U9938 (N_9938,N_3658,N_1410);
and U9939 (N_9939,N_5390,N_4489);
xor U9940 (N_9940,N_1441,N_1385);
nand U9941 (N_9941,N_1484,N_3071);
and U9942 (N_9942,N_6070,N_2015);
nand U9943 (N_9943,N_5942,N_2150);
nand U9944 (N_9944,N_2825,N_5365);
xnor U9945 (N_9945,N_2537,N_4956);
nand U9946 (N_9946,N_3596,N_25);
or U9947 (N_9947,N_4771,N_1248);
and U9948 (N_9948,N_3806,N_2354);
nor U9949 (N_9949,N_4951,N_5122);
nor U9950 (N_9950,N_3479,N_1621);
nand U9951 (N_9951,N_4744,N_751);
nor U9952 (N_9952,N_4072,N_5324);
and U9953 (N_9953,N_5287,N_5566);
and U9954 (N_9954,N_5700,N_1551);
and U9955 (N_9955,N_1822,N_4174);
nand U9956 (N_9956,N_6003,N_1425);
and U9957 (N_9957,N_5268,N_3456);
or U9958 (N_9958,N_5744,N_688);
xnor U9959 (N_9959,N_821,N_2264);
or U9960 (N_9960,N_5576,N_6145);
or U9961 (N_9961,N_6208,N_2913);
and U9962 (N_9962,N_4277,N_1950);
and U9963 (N_9963,N_1196,N_2215);
nor U9964 (N_9964,N_5967,N_2182);
or U9965 (N_9965,N_1424,N_5230);
or U9966 (N_9966,N_590,N_4923);
xor U9967 (N_9967,N_1888,N_1445);
and U9968 (N_9968,N_2493,N_960);
and U9969 (N_9969,N_6214,N_4383);
and U9970 (N_9970,N_496,N_2757);
xor U9971 (N_9971,N_4196,N_3793);
and U9972 (N_9972,N_385,N_3023);
nor U9973 (N_9973,N_3113,N_5043);
nand U9974 (N_9974,N_5390,N_3936);
nor U9975 (N_9975,N_1149,N_5858);
nand U9976 (N_9976,N_4311,N_5012);
and U9977 (N_9977,N_4877,N_925);
nand U9978 (N_9978,N_1690,N_2837);
or U9979 (N_9979,N_1904,N_2205);
nor U9980 (N_9980,N_1190,N_3870);
nor U9981 (N_9981,N_4153,N_6198);
and U9982 (N_9982,N_4291,N_4626);
and U9983 (N_9983,N_580,N_276);
and U9984 (N_9984,N_3928,N_5432);
and U9985 (N_9985,N_5089,N_1422);
nor U9986 (N_9986,N_3892,N_5796);
nor U9987 (N_9987,N_6218,N_5384);
and U9988 (N_9988,N_699,N_4361);
xor U9989 (N_9989,N_5299,N_520);
or U9990 (N_9990,N_4271,N_2896);
xnor U9991 (N_9991,N_2431,N_227);
and U9992 (N_9992,N_5039,N_4585);
and U9993 (N_9993,N_1316,N_4353);
nor U9994 (N_9994,N_1548,N_1897);
or U9995 (N_9995,N_3056,N_900);
nor U9996 (N_9996,N_5304,N_1730);
nor U9997 (N_9997,N_3272,N_124);
xnor U9998 (N_9998,N_1607,N_4501);
nand U9999 (N_9999,N_3533,N_293);
xor U10000 (N_10000,N_2388,N_2457);
and U10001 (N_10001,N_1909,N_5932);
nand U10002 (N_10002,N_1227,N_2880);
and U10003 (N_10003,N_3264,N_5210);
nand U10004 (N_10004,N_3793,N_1572);
xor U10005 (N_10005,N_703,N_6118);
xor U10006 (N_10006,N_1851,N_6094);
or U10007 (N_10007,N_5298,N_3825);
and U10008 (N_10008,N_3005,N_413);
nand U10009 (N_10009,N_931,N_2032);
nor U10010 (N_10010,N_213,N_4297);
nor U10011 (N_10011,N_1580,N_5833);
or U10012 (N_10012,N_5805,N_3944);
nor U10013 (N_10013,N_2697,N_863);
or U10014 (N_10014,N_216,N_3944);
nor U10015 (N_10015,N_3556,N_3809);
and U10016 (N_10016,N_1755,N_995);
or U10017 (N_10017,N_4624,N_6131);
nor U10018 (N_10018,N_5320,N_2690);
nand U10019 (N_10019,N_1369,N_4289);
nand U10020 (N_10020,N_5277,N_705);
and U10021 (N_10021,N_3060,N_2857);
and U10022 (N_10022,N_1275,N_6074);
nand U10023 (N_10023,N_5355,N_2312);
nand U10024 (N_10024,N_2458,N_3860);
xor U10025 (N_10025,N_2212,N_193);
xnor U10026 (N_10026,N_271,N_3904);
and U10027 (N_10027,N_6136,N_2327);
nand U10028 (N_10028,N_528,N_3301);
or U10029 (N_10029,N_616,N_2226);
or U10030 (N_10030,N_68,N_3651);
nor U10031 (N_10031,N_736,N_3816);
xor U10032 (N_10032,N_320,N_4774);
nor U10033 (N_10033,N_5500,N_624);
and U10034 (N_10034,N_3032,N_2377);
and U10035 (N_10035,N_4572,N_3263);
or U10036 (N_10036,N_4451,N_2220);
or U10037 (N_10037,N_773,N_27);
or U10038 (N_10038,N_5359,N_685);
or U10039 (N_10039,N_5449,N_1550);
nor U10040 (N_10040,N_5958,N_5702);
and U10041 (N_10041,N_3389,N_4831);
or U10042 (N_10042,N_2270,N_1740);
and U10043 (N_10043,N_279,N_3184);
nand U10044 (N_10044,N_5338,N_5016);
nand U10045 (N_10045,N_2805,N_6151);
or U10046 (N_10046,N_1391,N_4817);
or U10047 (N_10047,N_4437,N_4342);
nand U10048 (N_10048,N_4836,N_2460);
and U10049 (N_10049,N_2394,N_1758);
or U10050 (N_10050,N_1105,N_3309);
or U10051 (N_10051,N_4860,N_4141);
and U10052 (N_10052,N_5194,N_6100);
nand U10053 (N_10053,N_5474,N_5734);
or U10054 (N_10054,N_4462,N_1215);
and U10055 (N_10055,N_3601,N_1594);
or U10056 (N_10056,N_81,N_2366);
and U10057 (N_10057,N_6215,N_2912);
nand U10058 (N_10058,N_4954,N_172);
nor U10059 (N_10059,N_2571,N_4457);
or U10060 (N_10060,N_3885,N_1907);
and U10061 (N_10061,N_628,N_1057);
nor U10062 (N_10062,N_1813,N_4991);
nor U10063 (N_10063,N_4726,N_1385);
or U10064 (N_10064,N_3705,N_3977);
nand U10065 (N_10065,N_1343,N_1739);
nand U10066 (N_10066,N_1003,N_2549);
nor U10067 (N_10067,N_4185,N_1498);
and U10068 (N_10068,N_5279,N_1451);
xnor U10069 (N_10069,N_4392,N_2673);
nand U10070 (N_10070,N_4177,N_2911);
and U10071 (N_10071,N_4836,N_2185);
and U10072 (N_10072,N_6068,N_2390);
or U10073 (N_10073,N_357,N_5450);
nor U10074 (N_10074,N_1811,N_323);
nand U10075 (N_10075,N_3118,N_1421);
and U10076 (N_10076,N_2342,N_1954);
nand U10077 (N_10077,N_3142,N_5042);
nor U10078 (N_10078,N_4120,N_3033);
and U10079 (N_10079,N_2963,N_789);
xnor U10080 (N_10080,N_3596,N_1757);
nand U10081 (N_10081,N_297,N_314);
or U10082 (N_10082,N_2276,N_5589);
or U10083 (N_10083,N_4637,N_305);
or U10084 (N_10084,N_2130,N_2933);
nand U10085 (N_10085,N_5606,N_1828);
and U10086 (N_10086,N_4673,N_1978);
or U10087 (N_10087,N_4979,N_1859);
nand U10088 (N_10088,N_4252,N_1500);
nand U10089 (N_10089,N_590,N_3642);
and U10090 (N_10090,N_3477,N_5981);
and U10091 (N_10091,N_1597,N_1007);
nand U10092 (N_10092,N_1344,N_5825);
and U10093 (N_10093,N_3863,N_2647);
xor U10094 (N_10094,N_1622,N_1784);
nand U10095 (N_10095,N_5591,N_4014);
or U10096 (N_10096,N_5737,N_2055);
and U10097 (N_10097,N_887,N_1776);
or U10098 (N_10098,N_2505,N_3846);
nand U10099 (N_10099,N_567,N_1646);
nand U10100 (N_10100,N_4914,N_950);
xor U10101 (N_10101,N_6032,N_10);
and U10102 (N_10102,N_2392,N_251);
and U10103 (N_10103,N_5975,N_118);
or U10104 (N_10104,N_1872,N_5352);
nor U10105 (N_10105,N_5300,N_4095);
and U10106 (N_10106,N_3044,N_1391);
nor U10107 (N_10107,N_4033,N_5164);
nor U10108 (N_10108,N_282,N_1779);
nand U10109 (N_10109,N_6058,N_1286);
xor U10110 (N_10110,N_2901,N_5684);
nor U10111 (N_10111,N_4236,N_3343);
xnor U10112 (N_10112,N_1717,N_3440);
or U10113 (N_10113,N_4612,N_4799);
nor U10114 (N_10114,N_3722,N_1834);
nor U10115 (N_10115,N_1544,N_4599);
or U10116 (N_10116,N_3318,N_6055);
nand U10117 (N_10117,N_2801,N_1091);
and U10118 (N_10118,N_1463,N_748);
and U10119 (N_10119,N_5550,N_4736);
and U10120 (N_10120,N_2561,N_5568);
nand U10121 (N_10121,N_667,N_598);
nor U10122 (N_10122,N_3413,N_2847);
nand U10123 (N_10123,N_1716,N_3434);
nand U10124 (N_10124,N_2367,N_2189);
xnor U10125 (N_10125,N_3504,N_971);
nor U10126 (N_10126,N_1242,N_5376);
or U10127 (N_10127,N_3162,N_2728);
nand U10128 (N_10128,N_1705,N_1008);
or U10129 (N_10129,N_4972,N_4019);
nor U10130 (N_10130,N_4708,N_2475);
nor U10131 (N_10131,N_5825,N_3601);
nand U10132 (N_10132,N_3438,N_6199);
and U10133 (N_10133,N_1718,N_3878);
and U10134 (N_10134,N_5799,N_4948);
or U10135 (N_10135,N_2012,N_6217);
and U10136 (N_10136,N_3927,N_2297);
nor U10137 (N_10137,N_1316,N_2007);
nand U10138 (N_10138,N_3304,N_5057);
nand U10139 (N_10139,N_3120,N_2403);
nand U10140 (N_10140,N_3917,N_3651);
or U10141 (N_10141,N_1496,N_1052);
and U10142 (N_10142,N_1155,N_5160);
nor U10143 (N_10143,N_2622,N_3911);
and U10144 (N_10144,N_6223,N_1930);
or U10145 (N_10145,N_3253,N_3940);
and U10146 (N_10146,N_3343,N_4256);
or U10147 (N_10147,N_5829,N_937);
or U10148 (N_10148,N_4615,N_1599);
nand U10149 (N_10149,N_3879,N_749);
and U10150 (N_10150,N_2691,N_5329);
nand U10151 (N_10151,N_5786,N_6042);
or U10152 (N_10152,N_4137,N_4651);
nand U10153 (N_10153,N_1694,N_3924);
nor U10154 (N_10154,N_4900,N_1132);
and U10155 (N_10155,N_199,N_548);
or U10156 (N_10156,N_5241,N_3389);
and U10157 (N_10157,N_3337,N_1556);
nor U10158 (N_10158,N_4091,N_1920);
and U10159 (N_10159,N_3426,N_1388);
nor U10160 (N_10160,N_3060,N_3183);
nand U10161 (N_10161,N_826,N_5354);
nand U10162 (N_10162,N_5205,N_2594);
nor U10163 (N_10163,N_4138,N_6072);
nor U10164 (N_10164,N_4719,N_6109);
and U10165 (N_10165,N_1559,N_4213);
or U10166 (N_10166,N_6023,N_1584);
nor U10167 (N_10167,N_4825,N_3535);
and U10168 (N_10168,N_652,N_1326);
and U10169 (N_10169,N_4821,N_5954);
nand U10170 (N_10170,N_5977,N_3422);
and U10171 (N_10171,N_5244,N_1815);
or U10172 (N_10172,N_1987,N_614);
and U10173 (N_10173,N_2035,N_2970);
or U10174 (N_10174,N_4201,N_5012);
and U10175 (N_10175,N_3323,N_1206);
nand U10176 (N_10176,N_3421,N_5063);
xor U10177 (N_10177,N_5961,N_3188);
nand U10178 (N_10178,N_2522,N_1607);
nor U10179 (N_10179,N_705,N_967);
xnor U10180 (N_10180,N_2423,N_6117);
nand U10181 (N_10181,N_3215,N_1570);
and U10182 (N_10182,N_4325,N_2243);
or U10183 (N_10183,N_2475,N_813);
or U10184 (N_10184,N_5951,N_1043);
nor U10185 (N_10185,N_2067,N_2677);
and U10186 (N_10186,N_1015,N_6025);
xor U10187 (N_10187,N_216,N_2927);
xor U10188 (N_10188,N_307,N_5787);
and U10189 (N_10189,N_4066,N_4234);
or U10190 (N_10190,N_876,N_5154);
nand U10191 (N_10191,N_2669,N_1309);
and U10192 (N_10192,N_379,N_2599);
nor U10193 (N_10193,N_618,N_6012);
and U10194 (N_10194,N_4622,N_1589);
xnor U10195 (N_10195,N_3645,N_1849);
or U10196 (N_10196,N_2733,N_4005);
or U10197 (N_10197,N_4645,N_4832);
or U10198 (N_10198,N_5155,N_1420);
or U10199 (N_10199,N_2859,N_4294);
nor U10200 (N_10200,N_4481,N_2802);
nand U10201 (N_10201,N_5144,N_516);
nand U10202 (N_10202,N_4445,N_3118);
and U10203 (N_10203,N_4695,N_286);
or U10204 (N_10204,N_2121,N_5300);
and U10205 (N_10205,N_3056,N_3641);
or U10206 (N_10206,N_3797,N_3505);
or U10207 (N_10207,N_5538,N_3797);
xnor U10208 (N_10208,N_5062,N_3937);
and U10209 (N_10209,N_4294,N_3665);
nand U10210 (N_10210,N_4886,N_5614);
nand U10211 (N_10211,N_1279,N_4303);
and U10212 (N_10212,N_4346,N_2380);
nand U10213 (N_10213,N_3577,N_2955);
nand U10214 (N_10214,N_2240,N_4690);
and U10215 (N_10215,N_6129,N_3189);
xnor U10216 (N_10216,N_4439,N_4080);
or U10217 (N_10217,N_5851,N_902);
nor U10218 (N_10218,N_3630,N_5159);
and U10219 (N_10219,N_3210,N_2235);
nor U10220 (N_10220,N_2831,N_2501);
and U10221 (N_10221,N_90,N_2769);
nand U10222 (N_10222,N_990,N_3085);
xnor U10223 (N_10223,N_2368,N_436);
or U10224 (N_10224,N_90,N_5712);
nand U10225 (N_10225,N_3194,N_6201);
xor U10226 (N_10226,N_2804,N_1837);
nor U10227 (N_10227,N_579,N_2951);
xor U10228 (N_10228,N_1930,N_4987);
and U10229 (N_10229,N_3383,N_12);
xor U10230 (N_10230,N_2757,N_3951);
nor U10231 (N_10231,N_4587,N_6093);
nand U10232 (N_10232,N_4506,N_2364);
or U10233 (N_10233,N_3880,N_3477);
or U10234 (N_10234,N_2969,N_5399);
nor U10235 (N_10235,N_3046,N_4102);
or U10236 (N_10236,N_3318,N_408);
nand U10237 (N_10237,N_4951,N_2037);
nand U10238 (N_10238,N_2603,N_137);
or U10239 (N_10239,N_599,N_3725);
or U10240 (N_10240,N_1105,N_4646);
or U10241 (N_10241,N_826,N_4737);
or U10242 (N_10242,N_269,N_3842);
or U10243 (N_10243,N_134,N_3009);
nor U10244 (N_10244,N_1265,N_5361);
nor U10245 (N_10245,N_253,N_5629);
or U10246 (N_10246,N_3941,N_1945);
and U10247 (N_10247,N_1999,N_3718);
or U10248 (N_10248,N_3017,N_4887);
and U10249 (N_10249,N_602,N_3617);
xnor U10250 (N_10250,N_3700,N_5078);
or U10251 (N_10251,N_390,N_2454);
nor U10252 (N_10252,N_3928,N_2433);
nor U10253 (N_10253,N_4515,N_2375);
or U10254 (N_10254,N_1910,N_5064);
xnor U10255 (N_10255,N_5717,N_61);
and U10256 (N_10256,N_1803,N_1815);
nor U10257 (N_10257,N_3151,N_5272);
nand U10258 (N_10258,N_1156,N_725);
xor U10259 (N_10259,N_1170,N_5530);
and U10260 (N_10260,N_238,N_2711);
and U10261 (N_10261,N_3450,N_2489);
or U10262 (N_10262,N_1458,N_1933);
nand U10263 (N_10263,N_4559,N_5402);
or U10264 (N_10264,N_1434,N_3737);
or U10265 (N_10265,N_3050,N_1111);
xor U10266 (N_10266,N_3884,N_2374);
nand U10267 (N_10267,N_1157,N_2276);
nand U10268 (N_10268,N_1412,N_1118);
nor U10269 (N_10269,N_3037,N_1373);
and U10270 (N_10270,N_5833,N_3291);
nand U10271 (N_10271,N_4451,N_4789);
and U10272 (N_10272,N_2339,N_4869);
and U10273 (N_10273,N_3103,N_1461);
nand U10274 (N_10274,N_3384,N_6016);
or U10275 (N_10275,N_4429,N_5442);
and U10276 (N_10276,N_4448,N_5084);
and U10277 (N_10277,N_1968,N_4754);
and U10278 (N_10278,N_1702,N_1316);
nor U10279 (N_10279,N_989,N_2220);
and U10280 (N_10280,N_11,N_3064);
or U10281 (N_10281,N_3742,N_5225);
nor U10282 (N_10282,N_3660,N_3427);
xnor U10283 (N_10283,N_5425,N_2707);
nor U10284 (N_10284,N_956,N_2887);
nor U10285 (N_10285,N_4681,N_622);
or U10286 (N_10286,N_3094,N_5988);
nand U10287 (N_10287,N_3526,N_4132);
nand U10288 (N_10288,N_1698,N_5844);
or U10289 (N_10289,N_2737,N_478);
xnor U10290 (N_10290,N_1203,N_5671);
or U10291 (N_10291,N_1717,N_2801);
or U10292 (N_10292,N_454,N_2983);
nor U10293 (N_10293,N_1976,N_4079);
nor U10294 (N_10294,N_2069,N_545);
or U10295 (N_10295,N_5111,N_4323);
and U10296 (N_10296,N_4148,N_6127);
nor U10297 (N_10297,N_1125,N_6133);
nor U10298 (N_10298,N_6086,N_685);
nand U10299 (N_10299,N_5156,N_5433);
nor U10300 (N_10300,N_4069,N_3315);
or U10301 (N_10301,N_4746,N_5516);
xnor U10302 (N_10302,N_5697,N_4042);
nand U10303 (N_10303,N_3125,N_5813);
xor U10304 (N_10304,N_3950,N_1995);
or U10305 (N_10305,N_3791,N_2717);
nor U10306 (N_10306,N_5433,N_6143);
or U10307 (N_10307,N_2736,N_3587);
nand U10308 (N_10308,N_2997,N_2075);
nor U10309 (N_10309,N_3796,N_3368);
and U10310 (N_10310,N_3984,N_1123);
nor U10311 (N_10311,N_1453,N_614);
and U10312 (N_10312,N_3400,N_5191);
nand U10313 (N_10313,N_4478,N_5845);
nor U10314 (N_10314,N_5405,N_3794);
nand U10315 (N_10315,N_4761,N_3860);
and U10316 (N_10316,N_5197,N_5618);
or U10317 (N_10317,N_315,N_3321);
and U10318 (N_10318,N_1588,N_2113);
and U10319 (N_10319,N_5975,N_5407);
nand U10320 (N_10320,N_4500,N_845);
or U10321 (N_10321,N_148,N_4521);
and U10322 (N_10322,N_3261,N_4288);
nor U10323 (N_10323,N_5854,N_5979);
nor U10324 (N_10324,N_3432,N_3054);
nand U10325 (N_10325,N_262,N_797);
and U10326 (N_10326,N_1227,N_5388);
nor U10327 (N_10327,N_5898,N_4756);
nor U10328 (N_10328,N_3951,N_3113);
and U10329 (N_10329,N_2314,N_5411);
nor U10330 (N_10330,N_5017,N_2014);
nor U10331 (N_10331,N_2214,N_5589);
nor U10332 (N_10332,N_4403,N_977);
nor U10333 (N_10333,N_4290,N_898);
and U10334 (N_10334,N_5911,N_4600);
or U10335 (N_10335,N_4852,N_5490);
and U10336 (N_10336,N_5429,N_1049);
nor U10337 (N_10337,N_745,N_4820);
nor U10338 (N_10338,N_3396,N_3635);
nor U10339 (N_10339,N_4742,N_5118);
nand U10340 (N_10340,N_3820,N_3261);
and U10341 (N_10341,N_4117,N_6220);
or U10342 (N_10342,N_4254,N_667);
and U10343 (N_10343,N_3325,N_3645);
or U10344 (N_10344,N_1547,N_3278);
or U10345 (N_10345,N_2192,N_1603);
nand U10346 (N_10346,N_1870,N_4141);
nor U10347 (N_10347,N_2826,N_4881);
nor U10348 (N_10348,N_678,N_3492);
and U10349 (N_10349,N_5876,N_867);
or U10350 (N_10350,N_3867,N_2352);
and U10351 (N_10351,N_5124,N_2072);
nor U10352 (N_10352,N_4133,N_445);
and U10353 (N_10353,N_5009,N_3569);
nor U10354 (N_10354,N_1672,N_3549);
nand U10355 (N_10355,N_5208,N_1265);
or U10356 (N_10356,N_3461,N_2066);
xnor U10357 (N_10357,N_3312,N_6169);
and U10358 (N_10358,N_5312,N_253);
nor U10359 (N_10359,N_867,N_6068);
or U10360 (N_10360,N_4305,N_1290);
nor U10361 (N_10361,N_3104,N_4193);
and U10362 (N_10362,N_3422,N_6155);
and U10363 (N_10363,N_4199,N_1874);
or U10364 (N_10364,N_4406,N_1222);
or U10365 (N_10365,N_163,N_1192);
xnor U10366 (N_10366,N_4141,N_2257);
nand U10367 (N_10367,N_1285,N_3276);
nand U10368 (N_10368,N_5513,N_3327);
and U10369 (N_10369,N_2198,N_6079);
nand U10370 (N_10370,N_704,N_3067);
and U10371 (N_10371,N_165,N_6036);
or U10372 (N_10372,N_1297,N_5433);
nand U10373 (N_10373,N_5531,N_5964);
or U10374 (N_10374,N_2332,N_3218);
or U10375 (N_10375,N_4286,N_3412);
nor U10376 (N_10376,N_421,N_5162);
and U10377 (N_10377,N_3948,N_3851);
nor U10378 (N_10378,N_3139,N_3175);
and U10379 (N_10379,N_3743,N_5757);
nand U10380 (N_10380,N_1105,N_5010);
or U10381 (N_10381,N_2088,N_2668);
nand U10382 (N_10382,N_5924,N_3697);
and U10383 (N_10383,N_2195,N_801);
nand U10384 (N_10384,N_5703,N_1921);
nand U10385 (N_10385,N_3961,N_2903);
nand U10386 (N_10386,N_5177,N_1309);
or U10387 (N_10387,N_4017,N_5902);
xnor U10388 (N_10388,N_5077,N_5389);
nand U10389 (N_10389,N_6215,N_1611);
and U10390 (N_10390,N_2087,N_3112);
nand U10391 (N_10391,N_3817,N_2482);
nand U10392 (N_10392,N_505,N_5051);
xor U10393 (N_10393,N_4465,N_3703);
nor U10394 (N_10394,N_5006,N_673);
nor U10395 (N_10395,N_1694,N_1312);
or U10396 (N_10396,N_5183,N_20);
nor U10397 (N_10397,N_3110,N_189);
xor U10398 (N_10398,N_5149,N_4331);
and U10399 (N_10399,N_5127,N_5607);
or U10400 (N_10400,N_4018,N_5724);
and U10401 (N_10401,N_975,N_5330);
nor U10402 (N_10402,N_5299,N_63);
and U10403 (N_10403,N_3362,N_4187);
nor U10404 (N_10404,N_2404,N_1837);
nor U10405 (N_10405,N_5390,N_5401);
and U10406 (N_10406,N_4455,N_5136);
and U10407 (N_10407,N_5800,N_76);
nor U10408 (N_10408,N_1317,N_4580);
and U10409 (N_10409,N_3624,N_5996);
nand U10410 (N_10410,N_2111,N_777);
or U10411 (N_10411,N_830,N_451);
and U10412 (N_10412,N_4369,N_1051);
nor U10413 (N_10413,N_319,N_46);
nor U10414 (N_10414,N_4122,N_4428);
nand U10415 (N_10415,N_5995,N_2169);
nor U10416 (N_10416,N_2371,N_3620);
and U10417 (N_10417,N_3301,N_3007);
and U10418 (N_10418,N_894,N_3804);
and U10419 (N_10419,N_3109,N_2322);
or U10420 (N_10420,N_387,N_2427);
or U10421 (N_10421,N_1475,N_3770);
or U10422 (N_10422,N_4289,N_794);
and U10423 (N_10423,N_2899,N_3536);
and U10424 (N_10424,N_5323,N_2072);
nand U10425 (N_10425,N_601,N_2412);
nor U10426 (N_10426,N_2774,N_1701);
and U10427 (N_10427,N_1926,N_105);
and U10428 (N_10428,N_156,N_6064);
and U10429 (N_10429,N_2201,N_1454);
xor U10430 (N_10430,N_6134,N_390);
and U10431 (N_10431,N_6118,N_68);
nor U10432 (N_10432,N_5455,N_4001);
nand U10433 (N_10433,N_5717,N_37);
nand U10434 (N_10434,N_4557,N_5132);
or U10435 (N_10435,N_922,N_1177);
nand U10436 (N_10436,N_4538,N_2413);
and U10437 (N_10437,N_2919,N_2757);
nand U10438 (N_10438,N_454,N_4568);
or U10439 (N_10439,N_4438,N_5290);
nand U10440 (N_10440,N_4821,N_4380);
and U10441 (N_10441,N_4631,N_167);
nor U10442 (N_10442,N_5531,N_1221);
nor U10443 (N_10443,N_373,N_6242);
and U10444 (N_10444,N_4574,N_3063);
nand U10445 (N_10445,N_2182,N_2303);
nor U10446 (N_10446,N_405,N_1478);
and U10447 (N_10447,N_2572,N_4529);
nand U10448 (N_10448,N_3378,N_5979);
and U10449 (N_10449,N_5413,N_5734);
nor U10450 (N_10450,N_4056,N_691);
nand U10451 (N_10451,N_3663,N_6135);
and U10452 (N_10452,N_219,N_2409);
or U10453 (N_10453,N_641,N_5852);
nor U10454 (N_10454,N_5529,N_771);
or U10455 (N_10455,N_1516,N_3499);
nand U10456 (N_10456,N_5584,N_3804);
nor U10457 (N_10457,N_689,N_1614);
xnor U10458 (N_10458,N_4923,N_616);
nor U10459 (N_10459,N_3712,N_1280);
nor U10460 (N_10460,N_685,N_4150);
nor U10461 (N_10461,N_3276,N_3023);
xnor U10462 (N_10462,N_868,N_5264);
and U10463 (N_10463,N_3461,N_1402);
xnor U10464 (N_10464,N_230,N_2142);
nor U10465 (N_10465,N_5919,N_5547);
and U10466 (N_10466,N_4012,N_28);
and U10467 (N_10467,N_4426,N_184);
nor U10468 (N_10468,N_2098,N_5064);
nor U10469 (N_10469,N_1882,N_2522);
nand U10470 (N_10470,N_5361,N_1840);
and U10471 (N_10471,N_357,N_3145);
or U10472 (N_10472,N_4500,N_5857);
and U10473 (N_10473,N_3525,N_5995);
nand U10474 (N_10474,N_2608,N_1809);
or U10475 (N_10475,N_3383,N_3004);
xnor U10476 (N_10476,N_1481,N_489);
nand U10477 (N_10477,N_424,N_2432);
or U10478 (N_10478,N_133,N_3474);
and U10479 (N_10479,N_441,N_891);
or U10480 (N_10480,N_6202,N_4128);
nand U10481 (N_10481,N_1136,N_1742);
or U10482 (N_10482,N_1810,N_5707);
or U10483 (N_10483,N_899,N_3623);
nand U10484 (N_10484,N_4303,N_6249);
nor U10485 (N_10485,N_1571,N_235);
nor U10486 (N_10486,N_1779,N_3733);
or U10487 (N_10487,N_2687,N_5508);
and U10488 (N_10488,N_2545,N_1570);
and U10489 (N_10489,N_4154,N_3482);
nand U10490 (N_10490,N_511,N_4878);
nor U10491 (N_10491,N_1096,N_1030);
xnor U10492 (N_10492,N_2441,N_3543);
or U10493 (N_10493,N_6210,N_6187);
nand U10494 (N_10494,N_3386,N_760);
nor U10495 (N_10495,N_2926,N_4215);
xor U10496 (N_10496,N_2854,N_5042);
or U10497 (N_10497,N_129,N_1099);
or U10498 (N_10498,N_3457,N_1818);
or U10499 (N_10499,N_4234,N_247);
nor U10500 (N_10500,N_4547,N_2964);
nand U10501 (N_10501,N_3357,N_3163);
and U10502 (N_10502,N_1479,N_2695);
nand U10503 (N_10503,N_3886,N_4251);
and U10504 (N_10504,N_443,N_368);
nand U10505 (N_10505,N_6233,N_176);
nor U10506 (N_10506,N_342,N_5785);
nor U10507 (N_10507,N_2158,N_616);
nor U10508 (N_10508,N_154,N_3319);
and U10509 (N_10509,N_965,N_2164);
xor U10510 (N_10510,N_3681,N_4150);
xor U10511 (N_10511,N_2895,N_5804);
and U10512 (N_10512,N_176,N_3302);
nor U10513 (N_10513,N_5482,N_1458);
and U10514 (N_10514,N_2582,N_4190);
or U10515 (N_10515,N_5450,N_5884);
nand U10516 (N_10516,N_5063,N_930);
nand U10517 (N_10517,N_1601,N_5854);
nor U10518 (N_10518,N_1806,N_4032);
nor U10519 (N_10519,N_3815,N_4130);
nor U10520 (N_10520,N_1121,N_1517);
nand U10521 (N_10521,N_1033,N_5383);
nand U10522 (N_10522,N_2748,N_1621);
and U10523 (N_10523,N_5910,N_899);
or U10524 (N_10524,N_3504,N_1011);
nand U10525 (N_10525,N_1679,N_2265);
nor U10526 (N_10526,N_3004,N_1304);
nand U10527 (N_10527,N_3973,N_2488);
nor U10528 (N_10528,N_5016,N_848);
nand U10529 (N_10529,N_1520,N_5290);
nand U10530 (N_10530,N_1194,N_3133);
nand U10531 (N_10531,N_1498,N_914);
nor U10532 (N_10532,N_2111,N_2734);
and U10533 (N_10533,N_4539,N_2189);
and U10534 (N_10534,N_5110,N_5037);
or U10535 (N_10535,N_1018,N_6006);
nand U10536 (N_10536,N_2676,N_1937);
nand U10537 (N_10537,N_583,N_5597);
and U10538 (N_10538,N_271,N_4754);
and U10539 (N_10539,N_5945,N_5484);
xor U10540 (N_10540,N_3357,N_4433);
or U10541 (N_10541,N_4438,N_5744);
nor U10542 (N_10542,N_2230,N_3581);
and U10543 (N_10543,N_874,N_2263);
nand U10544 (N_10544,N_5239,N_5224);
nor U10545 (N_10545,N_2810,N_2606);
nor U10546 (N_10546,N_5497,N_3067);
nand U10547 (N_10547,N_1204,N_1241);
or U10548 (N_10548,N_4484,N_5642);
xnor U10549 (N_10549,N_4023,N_412);
nor U10550 (N_10550,N_1660,N_411);
or U10551 (N_10551,N_3579,N_4128);
nand U10552 (N_10552,N_335,N_1734);
nand U10553 (N_10553,N_4352,N_3830);
nand U10554 (N_10554,N_986,N_5215);
and U10555 (N_10555,N_4313,N_4484);
or U10556 (N_10556,N_1171,N_539);
nor U10557 (N_10557,N_2893,N_116);
nor U10558 (N_10558,N_1261,N_2729);
or U10559 (N_10559,N_5636,N_2702);
and U10560 (N_10560,N_907,N_66);
nand U10561 (N_10561,N_5593,N_4986);
or U10562 (N_10562,N_4822,N_1855);
or U10563 (N_10563,N_5909,N_2567);
and U10564 (N_10564,N_3036,N_5565);
nand U10565 (N_10565,N_946,N_564);
nand U10566 (N_10566,N_1220,N_1340);
nor U10567 (N_10567,N_5561,N_105);
or U10568 (N_10568,N_2411,N_2918);
nor U10569 (N_10569,N_4087,N_820);
nand U10570 (N_10570,N_2830,N_2116);
or U10571 (N_10571,N_5246,N_4863);
nand U10572 (N_10572,N_5491,N_4226);
or U10573 (N_10573,N_3244,N_5828);
or U10574 (N_10574,N_492,N_3180);
nand U10575 (N_10575,N_4077,N_2386);
nor U10576 (N_10576,N_3356,N_1140);
nand U10577 (N_10577,N_3703,N_3638);
nand U10578 (N_10578,N_593,N_3111);
or U10579 (N_10579,N_558,N_3529);
xor U10580 (N_10580,N_2813,N_4688);
nand U10581 (N_10581,N_5461,N_4755);
or U10582 (N_10582,N_5457,N_616);
and U10583 (N_10583,N_1427,N_168);
nand U10584 (N_10584,N_673,N_615);
nand U10585 (N_10585,N_31,N_3374);
nand U10586 (N_10586,N_5942,N_6055);
nor U10587 (N_10587,N_1914,N_2296);
xnor U10588 (N_10588,N_2856,N_4896);
or U10589 (N_10589,N_1191,N_646);
or U10590 (N_10590,N_4228,N_2781);
nand U10591 (N_10591,N_5219,N_2068);
nor U10592 (N_10592,N_3689,N_6199);
and U10593 (N_10593,N_610,N_5931);
xor U10594 (N_10594,N_2420,N_334);
nor U10595 (N_10595,N_1926,N_3759);
and U10596 (N_10596,N_209,N_652);
or U10597 (N_10597,N_1624,N_2925);
or U10598 (N_10598,N_2597,N_2968);
or U10599 (N_10599,N_574,N_1681);
nor U10600 (N_10600,N_5715,N_5137);
and U10601 (N_10601,N_5442,N_3486);
and U10602 (N_10602,N_77,N_4433);
and U10603 (N_10603,N_3460,N_4860);
nor U10604 (N_10604,N_2260,N_1989);
and U10605 (N_10605,N_4969,N_1054);
nand U10606 (N_10606,N_3306,N_1055);
xor U10607 (N_10607,N_987,N_1542);
nand U10608 (N_10608,N_13,N_1435);
nand U10609 (N_10609,N_3156,N_527);
nor U10610 (N_10610,N_520,N_3755);
nand U10611 (N_10611,N_1805,N_4302);
xor U10612 (N_10612,N_2165,N_2185);
or U10613 (N_10613,N_2544,N_4740);
xor U10614 (N_10614,N_2750,N_727);
or U10615 (N_10615,N_4528,N_798);
nand U10616 (N_10616,N_2050,N_5101);
and U10617 (N_10617,N_4164,N_1063);
or U10618 (N_10618,N_1501,N_3858);
or U10619 (N_10619,N_4384,N_5064);
and U10620 (N_10620,N_5188,N_5338);
nand U10621 (N_10621,N_5608,N_836);
nor U10622 (N_10622,N_1319,N_2776);
and U10623 (N_10623,N_3901,N_4313);
and U10624 (N_10624,N_4032,N_5512);
xor U10625 (N_10625,N_307,N_5465);
xnor U10626 (N_10626,N_5285,N_979);
nand U10627 (N_10627,N_2915,N_2711);
nand U10628 (N_10628,N_762,N_5906);
nand U10629 (N_10629,N_743,N_2010);
nand U10630 (N_10630,N_283,N_2146);
nor U10631 (N_10631,N_266,N_1593);
or U10632 (N_10632,N_5132,N_3482);
and U10633 (N_10633,N_5274,N_6162);
nand U10634 (N_10634,N_2423,N_4492);
or U10635 (N_10635,N_2726,N_2895);
nand U10636 (N_10636,N_2739,N_4987);
nand U10637 (N_10637,N_343,N_5767);
nor U10638 (N_10638,N_1678,N_97);
nor U10639 (N_10639,N_5595,N_5198);
and U10640 (N_10640,N_6084,N_210);
and U10641 (N_10641,N_1155,N_2990);
nand U10642 (N_10642,N_2081,N_933);
or U10643 (N_10643,N_4903,N_5620);
or U10644 (N_10644,N_5268,N_4869);
nor U10645 (N_10645,N_1024,N_756);
nor U10646 (N_10646,N_2988,N_2840);
or U10647 (N_10647,N_1726,N_748);
or U10648 (N_10648,N_819,N_1649);
nor U10649 (N_10649,N_5131,N_2834);
or U10650 (N_10650,N_5491,N_3496);
or U10651 (N_10651,N_1340,N_5773);
or U10652 (N_10652,N_6187,N_3920);
nand U10653 (N_10653,N_3200,N_265);
or U10654 (N_10654,N_3323,N_1831);
nand U10655 (N_10655,N_2286,N_5888);
or U10656 (N_10656,N_3951,N_2459);
and U10657 (N_10657,N_5588,N_1025);
or U10658 (N_10658,N_2889,N_4980);
or U10659 (N_10659,N_2942,N_4998);
nor U10660 (N_10660,N_1065,N_126);
nor U10661 (N_10661,N_3537,N_3615);
nand U10662 (N_10662,N_721,N_3284);
or U10663 (N_10663,N_5687,N_1194);
nor U10664 (N_10664,N_3385,N_4257);
nand U10665 (N_10665,N_104,N_5062);
nand U10666 (N_10666,N_2524,N_4201);
or U10667 (N_10667,N_1168,N_3130);
nand U10668 (N_10668,N_3835,N_5988);
and U10669 (N_10669,N_3905,N_565);
and U10670 (N_10670,N_5070,N_1782);
nor U10671 (N_10671,N_2936,N_4895);
nor U10672 (N_10672,N_5652,N_2581);
or U10673 (N_10673,N_3711,N_4300);
or U10674 (N_10674,N_2527,N_4229);
or U10675 (N_10675,N_35,N_3523);
or U10676 (N_10676,N_2856,N_2414);
or U10677 (N_10677,N_3389,N_2868);
xnor U10678 (N_10678,N_1265,N_1056);
nor U10679 (N_10679,N_3515,N_635);
and U10680 (N_10680,N_4912,N_6114);
nor U10681 (N_10681,N_5546,N_1387);
and U10682 (N_10682,N_669,N_3644);
or U10683 (N_10683,N_5385,N_3926);
nor U10684 (N_10684,N_1022,N_1031);
xor U10685 (N_10685,N_4650,N_3746);
and U10686 (N_10686,N_316,N_536);
and U10687 (N_10687,N_4241,N_4324);
nor U10688 (N_10688,N_755,N_5014);
nor U10689 (N_10689,N_1443,N_4776);
nand U10690 (N_10690,N_2645,N_915);
nand U10691 (N_10691,N_128,N_1611);
nor U10692 (N_10692,N_1077,N_3627);
and U10693 (N_10693,N_2585,N_1039);
and U10694 (N_10694,N_4503,N_5862);
and U10695 (N_10695,N_5762,N_2445);
or U10696 (N_10696,N_3082,N_4118);
nand U10697 (N_10697,N_2785,N_3469);
and U10698 (N_10698,N_5508,N_2043);
nand U10699 (N_10699,N_241,N_2423);
or U10700 (N_10700,N_4711,N_3254);
and U10701 (N_10701,N_4910,N_1745);
nor U10702 (N_10702,N_4212,N_2278);
or U10703 (N_10703,N_4193,N_5808);
nand U10704 (N_10704,N_850,N_3161);
nand U10705 (N_10705,N_1120,N_2211);
or U10706 (N_10706,N_4005,N_2218);
nand U10707 (N_10707,N_2681,N_3063);
or U10708 (N_10708,N_774,N_2684);
nand U10709 (N_10709,N_156,N_1173);
nand U10710 (N_10710,N_5184,N_3628);
nor U10711 (N_10711,N_3411,N_4173);
xnor U10712 (N_10712,N_2452,N_3978);
nand U10713 (N_10713,N_4429,N_1196);
nor U10714 (N_10714,N_2047,N_2838);
and U10715 (N_10715,N_1497,N_81);
nor U10716 (N_10716,N_671,N_2159);
nand U10717 (N_10717,N_2595,N_4978);
nor U10718 (N_10718,N_5879,N_1891);
nand U10719 (N_10719,N_3102,N_3445);
xnor U10720 (N_10720,N_3739,N_4252);
and U10721 (N_10721,N_4844,N_1046);
nor U10722 (N_10722,N_555,N_2837);
nor U10723 (N_10723,N_3194,N_1953);
and U10724 (N_10724,N_3726,N_6217);
nand U10725 (N_10725,N_3034,N_2289);
and U10726 (N_10726,N_3044,N_3975);
or U10727 (N_10727,N_2620,N_3494);
or U10728 (N_10728,N_4446,N_5982);
nor U10729 (N_10729,N_3921,N_4133);
nand U10730 (N_10730,N_6144,N_3345);
xor U10731 (N_10731,N_4307,N_4329);
and U10732 (N_10732,N_2290,N_2799);
nor U10733 (N_10733,N_344,N_607);
or U10734 (N_10734,N_4900,N_6216);
and U10735 (N_10735,N_2330,N_4010);
nand U10736 (N_10736,N_3714,N_1855);
nand U10737 (N_10737,N_1757,N_4682);
nand U10738 (N_10738,N_216,N_6246);
xor U10739 (N_10739,N_317,N_1728);
or U10740 (N_10740,N_4864,N_1542);
nor U10741 (N_10741,N_609,N_166);
nor U10742 (N_10742,N_1555,N_4443);
or U10743 (N_10743,N_3822,N_3107);
and U10744 (N_10744,N_3369,N_76);
nor U10745 (N_10745,N_2678,N_3798);
or U10746 (N_10746,N_1301,N_4164);
or U10747 (N_10747,N_264,N_2346);
nand U10748 (N_10748,N_4643,N_5685);
or U10749 (N_10749,N_2774,N_1117);
and U10750 (N_10750,N_4416,N_1222);
and U10751 (N_10751,N_6224,N_3859);
or U10752 (N_10752,N_3578,N_2657);
nand U10753 (N_10753,N_85,N_1905);
and U10754 (N_10754,N_2017,N_1357);
nand U10755 (N_10755,N_3852,N_2253);
xor U10756 (N_10756,N_3925,N_2826);
nand U10757 (N_10757,N_2129,N_5330);
and U10758 (N_10758,N_2866,N_1281);
or U10759 (N_10759,N_3498,N_2167);
and U10760 (N_10760,N_390,N_4975);
and U10761 (N_10761,N_1701,N_5597);
or U10762 (N_10762,N_1892,N_5821);
and U10763 (N_10763,N_5797,N_321);
nor U10764 (N_10764,N_3058,N_713);
or U10765 (N_10765,N_3775,N_5705);
nand U10766 (N_10766,N_1360,N_5163);
nor U10767 (N_10767,N_2318,N_5079);
nor U10768 (N_10768,N_856,N_11);
and U10769 (N_10769,N_1628,N_2283);
or U10770 (N_10770,N_5473,N_4388);
and U10771 (N_10771,N_3750,N_3761);
nor U10772 (N_10772,N_1583,N_2976);
nand U10773 (N_10773,N_3452,N_4592);
or U10774 (N_10774,N_1418,N_16);
and U10775 (N_10775,N_5912,N_2676);
and U10776 (N_10776,N_6059,N_6147);
nand U10777 (N_10777,N_2403,N_4231);
or U10778 (N_10778,N_4529,N_33);
or U10779 (N_10779,N_2937,N_523);
nor U10780 (N_10780,N_5779,N_2755);
and U10781 (N_10781,N_3786,N_2106);
or U10782 (N_10782,N_4831,N_5703);
nand U10783 (N_10783,N_2614,N_3032);
or U10784 (N_10784,N_3233,N_1104);
nand U10785 (N_10785,N_1833,N_5532);
nand U10786 (N_10786,N_2234,N_5420);
xnor U10787 (N_10787,N_2117,N_5667);
and U10788 (N_10788,N_4373,N_3225);
xor U10789 (N_10789,N_492,N_2576);
or U10790 (N_10790,N_5542,N_2720);
and U10791 (N_10791,N_338,N_2793);
and U10792 (N_10792,N_6243,N_6082);
nand U10793 (N_10793,N_735,N_6242);
xnor U10794 (N_10794,N_4341,N_5907);
nand U10795 (N_10795,N_252,N_4629);
nand U10796 (N_10796,N_1493,N_310);
or U10797 (N_10797,N_223,N_5505);
nor U10798 (N_10798,N_5427,N_939);
and U10799 (N_10799,N_66,N_4245);
nor U10800 (N_10800,N_980,N_341);
and U10801 (N_10801,N_2602,N_5575);
nor U10802 (N_10802,N_4966,N_6039);
nand U10803 (N_10803,N_4460,N_4717);
nor U10804 (N_10804,N_5977,N_4737);
and U10805 (N_10805,N_5314,N_4391);
or U10806 (N_10806,N_142,N_2941);
nor U10807 (N_10807,N_5156,N_460);
and U10808 (N_10808,N_1865,N_3939);
and U10809 (N_10809,N_4532,N_665);
nor U10810 (N_10810,N_3833,N_4011);
xor U10811 (N_10811,N_2478,N_5730);
nor U10812 (N_10812,N_5349,N_2340);
or U10813 (N_10813,N_691,N_3784);
nand U10814 (N_10814,N_3670,N_5663);
or U10815 (N_10815,N_847,N_5886);
nor U10816 (N_10816,N_3761,N_3082);
or U10817 (N_10817,N_5955,N_3219);
nand U10818 (N_10818,N_5505,N_3867);
or U10819 (N_10819,N_1906,N_1608);
nand U10820 (N_10820,N_2590,N_1268);
and U10821 (N_10821,N_3944,N_6148);
or U10822 (N_10822,N_6220,N_1235);
or U10823 (N_10823,N_1662,N_1132);
xnor U10824 (N_10824,N_2826,N_2214);
xor U10825 (N_10825,N_3973,N_3478);
and U10826 (N_10826,N_2864,N_3265);
or U10827 (N_10827,N_2928,N_2134);
nand U10828 (N_10828,N_3153,N_2103);
nor U10829 (N_10829,N_5424,N_5581);
and U10830 (N_10830,N_1084,N_69);
and U10831 (N_10831,N_2592,N_2418);
and U10832 (N_10832,N_2144,N_4285);
or U10833 (N_10833,N_4723,N_1140);
and U10834 (N_10834,N_4853,N_1481);
nand U10835 (N_10835,N_305,N_1856);
nand U10836 (N_10836,N_2475,N_3655);
nor U10837 (N_10837,N_5955,N_5179);
nor U10838 (N_10838,N_2006,N_2580);
nor U10839 (N_10839,N_5658,N_206);
and U10840 (N_10840,N_788,N_1699);
or U10841 (N_10841,N_1332,N_2075);
nor U10842 (N_10842,N_1866,N_5829);
nand U10843 (N_10843,N_1637,N_5583);
or U10844 (N_10844,N_3120,N_1007);
or U10845 (N_10845,N_3412,N_1673);
and U10846 (N_10846,N_218,N_3710);
nand U10847 (N_10847,N_5621,N_3970);
nor U10848 (N_10848,N_2578,N_5481);
and U10849 (N_10849,N_4714,N_3430);
nand U10850 (N_10850,N_816,N_852);
nor U10851 (N_10851,N_6112,N_4228);
or U10852 (N_10852,N_3311,N_2937);
and U10853 (N_10853,N_1243,N_4492);
and U10854 (N_10854,N_4132,N_4055);
and U10855 (N_10855,N_1780,N_1666);
xor U10856 (N_10856,N_1008,N_4368);
and U10857 (N_10857,N_997,N_3896);
nor U10858 (N_10858,N_2695,N_2822);
nor U10859 (N_10859,N_5438,N_4043);
or U10860 (N_10860,N_5880,N_4148);
and U10861 (N_10861,N_378,N_4383);
and U10862 (N_10862,N_1466,N_3505);
xor U10863 (N_10863,N_5299,N_2390);
nor U10864 (N_10864,N_962,N_2059);
nor U10865 (N_10865,N_153,N_4381);
and U10866 (N_10866,N_3381,N_3379);
nand U10867 (N_10867,N_2276,N_2759);
nor U10868 (N_10868,N_5504,N_2187);
nand U10869 (N_10869,N_213,N_5131);
and U10870 (N_10870,N_1877,N_2873);
nand U10871 (N_10871,N_681,N_4202);
nor U10872 (N_10872,N_3742,N_4994);
and U10873 (N_10873,N_512,N_5038);
nand U10874 (N_10874,N_3567,N_2732);
or U10875 (N_10875,N_2628,N_535);
or U10876 (N_10876,N_1228,N_526);
and U10877 (N_10877,N_273,N_2188);
nand U10878 (N_10878,N_3196,N_809);
nand U10879 (N_10879,N_4700,N_6240);
and U10880 (N_10880,N_4944,N_1764);
nand U10881 (N_10881,N_5934,N_501);
or U10882 (N_10882,N_1202,N_4094);
nand U10883 (N_10883,N_5729,N_4314);
or U10884 (N_10884,N_2877,N_6155);
or U10885 (N_10885,N_2106,N_2770);
nor U10886 (N_10886,N_1007,N_5276);
or U10887 (N_10887,N_2615,N_428);
nand U10888 (N_10888,N_2531,N_4933);
nor U10889 (N_10889,N_3203,N_1621);
nor U10890 (N_10890,N_2109,N_5544);
and U10891 (N_10891,N_4667,N_3883);
nand U10892 (N_10892,N_548,N_407);
and U10893 (N_10893,N_2357,N_4840);
xnor U10894 (N_10894,N_6015,N_5480);
nor U10895 (N_10895,N_6084,N_5821);
nor U10896 (N_10896,N_5219,N_5197);
nand U10897 (N_10897,N_5087,N_2104);
or U10898 (N_10898,N_5888,N_1543);
or U10899 (N_10899,N_908,N_2318);
and U10900 (N_10900,N_3409,N_780);
and U10901 (N_10901,N_966,N_5504);
and U10902 (N_10902,N_603,N_1878);
nor U10903 (N_10903,N_6126,N_3547);
xor U10904 (N_10904,N_4523,N_1189);
nor U10905 (N_10905,N_3443,N_463);
nor U10906 (N_10906,N_4117,N_4237);
nand U10907 (N_10907,N_307,N_3787);
and U10908 (N_10908,N_3470,N_987);
xor U10909 (N_10909,N_1017,N_4202);
or U10910 (N_10910,N_5531,N_6095);
and U10911 (N_10911,N_241,N_177);
or U10912 (N_10912,N_4254,N_6061);
and U10913 (N_10913,N_5215,N_5320);
nand U10914 (N_10914,N_1325,N_3332);
and U10915 (N_10915,N_4952,N_4157);
nor U10916 (N_10916,N_3628,N_1541);
nor U10917 (N_10917,N_978,N_4714);
xor U10918 (N_10918,N_4150,N_2893);
and U10919 (N_10919,N_2228,N_3770);
xor U10920 (N_10920,N_4842,N_3372);
or U10921 (N_10921,N_1862,N_2722);
or U10922 (N_10922,N_2732,N_6214);
or U10923 (N_10923,N_1752,N_863);
nor U10924 (N_10924,N_2697,N_1272);
nor U10925 (N_10925,N_400,N_1243);
and U10926 (N_10926,N_5323,N_2004);
xor U10927 (N_10927,N_4011,N_3976);
and U10928 (N_10928,N_6064,N_4376);
xor U10929 (N_10929,N_4425,N_3667);
or U10930 (N_10930,N_2624,N_2662);
nor U10931 (N_10931,N_5285,N_346);
and U10932 (N_10932,N_5205,N_1950);
nor U10933 (N_10933,N_2241,N_2883);
and U10934 (N_10934,N_4724,N_2090);
or U10935 (N_10935,N_582,N_1421);
nand U10936 (N_10936,N_3995,N_1598);
xor U10937 (N_10937,N_3064,N_3863);
or U10938 (N_10938,N_2938,N_1878);
nor U10939 (N_10939,N_970,N_1003);
and U10940 (N_10940,N_2626,N_4360);
and U10941 (N_10941,N_1567,N_349);
or U10942 (N_10942,N_2387,N_1043);
nand U10943 (N_10943,N_3657,N_730);
xnor U10944 (N_10944,N_5574,N_3801);
nor U10945 (N_10945,N_51,N_3898);
xnor U10946 (N_10946,N_5997,N_3546);
or U10947 (N_10947,N_3237,N_3788);
nand U10948 (N_10948,N_6143,N_695);
nand U10949 (N_10949,N_5693,N_2908);
or U10950 (N_10950,N_3606,N_4811);
or U10951 (N_10951,N_576,N_6192);
or U10952 (N_10952,N_2641,N_1241);
xnor U10953 (N_10953,N_2086,N_2463);
nor U10954 (N_10954,N_6084,N_1825);
nand U10955 (N_10955,N_1548,N_4502);
or U10956 (N_10956,N_3108,N_5943);
or U10957 (N_10957,N_6014,N_760);
or U10958 (N_10958,N_6028,N_1466);
nand U10959 (N_10959,N_4616,N_5482);
or U10960 (N_10960,N_3729,N_1797);
nor U10961 (N_10961,N_5649,N_3292);
nor U10962 (N_10962,N_4325,N_4443);
and U10963 (N_10963,N_3974,N_4066);
nor U10964 (N_10964,N_3428,N_2715);
nor U10965 (N_10965,N_1006,N_205);
nand U10966 (N_10966,N_3904,N_3578);
nor U10967 (N_10967,N_3429,N_5695);
and U10968 (N_10968,N_374,N_5351);
nand U10969 (N_10969,N_1102,N_1504);
or U10970 (N_10970,N_651,N_4476);
xnor U10971 (N_10971,N_474,N_3487);
or U10972 (N_10972,N_823,N_370);
or U10973 (N_10973,N_4659,N_914);
nor U10974 (N_10974,N_2545,N_4461);
nor U10975 (N_10975,N_5048,N_6141);
or U10976 (N_10976,N_1871,N_4007);
nand U10977 (N_10977,N_2875,N_5694);
or U10978 (N_10978,N_3208,N_5122);
nand U10979 (N_10979,N_1204,N_6108);
or U10980 (N_10980,N_4775,N_347);
xnor U10981 (N_10981,N_924,N_1044);
nand U10982 (N_10982,N_2097,N_5915);
and U10983 (N_10983,N_4110,N_1788);
nand U10984 (N_10984,N_2717,N_3597);
nand U10985 (N_10985,N_5866,N_3232);
or U10986 (N_10986,N_2501,N_6107);
nor U10987 (N_10987,N_18,N_4945);
or U10988 (N_10988,N_4119,N_5266);
or U10989 (N_10989,N_6097,N_2269);
nor U10990 (N_10990,N_4434,N_4549);
nand U10991 (N_10991,N_2130,N_6226);
or U10992 (N_10992,N_2065,N_2135);
nor U10993 (N_10993,N_1360,N_2948);
or U10994 (N_10994,N_4611,N_3903);
or U10995 (N_10995,N_1382,N_4955);
or U10996 (N_10996,N_1866,N_4831);
or U10997 (N_10997,N_763,N_4762);
and U10998 (N_10998,N_5182,N_2253);
nor U10999 (N_10999,N_2715,N_4886);
nand U11000 (N_11000,N_4703,N_1803);
nor U11001 (N_11001,N_5102,N_4686);
or U11002 (N_11002,N_2646,N_81);
nand U11003 (N_11003,N_2807,N_505);
nand U11004 (N_11004,N_3369,N_1074);
nand U11005 (N_11005,N_5900,N_1943);
nand U11006 (N_11006,N_5369,N_2735);
and U11007 (N_11007,N_90,N_5035);
and U11008 (N_11008,N_5693,N_4242);
nand U11009 (N_11009,N_2796,N_5096);
nor U11010 (N_11010,N_667,N_3617);
or U11011 (N_11011,N_4899,N_4023);
xor U11012 (N_11012,N_5903,N_2437);
or U11013 (N_11013,N_1851,N_292);
nor U11014 (N_11014,N_2644,N_4877);
nor U11015 (N_11015,N_5903,N_405);
xor U11016 (N_11016,N_2457,N_486);
and U11017 (N_11017,N_2574,N_6161);
and U11018 (N_11018,N_1220,N_4090);
and U11019 (N_11019,N_2023,N_5239);
nand U11020 (N_11020,N_446,N_6133);
or U11021 (N_11021,N_1315,N_1907);
xor U11022 (N_11022,N_1098,N_2937);
nand U11023 (N_11023,N_5882,N_2974);
and U11024 (N_11024,N_1031,N_4219);
nand U11025 (N_11025,N_5789,N_5514);
and U11026 (N_11026,N_4745,N_4495);
nand U11027 (N_11027,N_6152,N_2375);
and U11028 (N_11028,N_5412,N_5611);
or U11029 (N_11029,N_4341,N_1544);
nand U11030 (N_11030,N_1711,N_5405);
nor U11031 (N_11031,N_2529,N_2874);
nor U11032 (N_11032,N_3176,N_4368);
nor U11033 (N_11033,N_5518,N_3476);
xor U11034 (N_11034,N_4093,N_4136);
and U11035 (N_11035,N_4208,N_3461);
and U11036 (N_11036,N_1881,N_2304);
nor U11037 (N_11037,N_2203,N_2489);
xor U11038 (N_11038,N_6154,N_5801);
nand U11039 (N_11039,N_3094,N_1115);
nor U11040 (N_11040,N_1596,N_4309);
nor U11041 (N_11041,N_640,N_5085);
and U11042 (N_11042,N_159,N_2095);
nand U11043 (N_11043,N_5455,N_2753);
and U11044 (N_11044,N_3320,N_5126);
xor U11045 (N_11045,N_5700,N_2754);
nor U11046 (N_11046,N_4229,N_282);
xor U11047 (N_11047,N_5669,N_4379);
nor U11048 (N_11048,N_5794,N_1923);
or U11049 (N_11049,N_1398,N_5427);
and U11050 (N_11050,N_4721,N_5502);
and U11051 (N_11051,N_507,N_4044);
nand U11052 (N_11052,N_3819,N_4239);
nor U11053 (N_11053,N_1060,N_3034);
nand U11054 (N_11054,N_3568,N_4436);
and U11055 (N_11055,N_960,N_916);
nand U11056 (N_11056,N_2424,N_1654);
or U11057 (N_11057,N_687,N_5061);
xor U11058 (N_11058,N_1351,N_1905);
xnor U11059 (N_11059,N_4975,N_4981);
and U11060 (N_11060,N_5811,N_4099);
nor U11061 (N_11061,N_408,N_2039);
nand U11062 (N_11062,N_6176,N_5605);
nand U11063 (N_11063,N_4915,N_293);
nor U11064 (N_11064,N_2284,N_4671);
nor U11065 (N_11065,N_5553,N_1818);
nand U11066 (N_11066,N_654,N_1154);
nor U11067 (N_11067,N_6133,N_3163);
and U11068 (N_11068,N_873,N_4485);
nand U11069 (N_11069,N_5073,N_6182);
and U11070 (N_11070,N_6042,N_3630);
nand U11071 (N_11071,N_2695,N_5259);
nand U11072 (N_11072,N_3739,N_2960);
and U11073 (N_11073,N_79,N_1478);
nand U11074 (N_11074,N_6119,N_6008);
or U11075 (N_11075,N_3506,N_2355);
and U11076 (N_11076,N_6169,N_4604);
nand U11077 (N_11077,N_4332,N_1530);
nand U11078 (N_11078,N_568,N_2393);
and U11079 (N_11079,N_5651,N_3342);
and U11080 (N_11080,N_6082,N_3112);
and U11081 (N_11081,N_4187,N_671);
nand U11082 (N_11082,N_5111,N_2591);
nand U11083 (N_11083,N_4168,N_2724);
nor U11084 (N_11084,N_1796,N_2559);
nor U11085 (N_11085,N_3148,N_2315);
or U11086 (N_11086,N_2369,N_3903);
and U11087 (N_11087,N_5834,N_30);
nor U11088 (N_11088,N_5895,N_862);
nor U11089 (N_11089,N_4047,N_2099);
nor U11090 (N_11090,N_5992,N_1687);
nand U11091 (N_11091,N_4670,N_4159);
nor U11092 (N_11092,N_4423,N_2916);
or U11093 (N_11093,N_2687,N_1619);
nor U11094 (N_11094,N_401,N_2766);
nor U11095 (N_11095,N_473,N_3322);
xor U11096 (N_11096,N_1043,N_5362);
xnor U11097 (N_11097,N_5378,N_1217);
or U11098 (N_11098,N_2022,N_5963);
nor U11099 (N_11099,N_2597,N_3048);
and U11100 (N_11100,N_5668,N_1576);
or U11101 (N_11101,N_1332,N_5073);
and U11102 (N_11102,N_4697,N_1457);
nor U11103 (N_11103,N_4314,N_2473);
xor U11104 (N_11104,N_172,N_4380);
nor U11105 (N_11105,N_2709,N_2456);
nor U11106 (N_11106,N_4167,N_354);
and U11107 (N_11107,N_3774,N_4035);
or U11108 (N_11108,N_3652,N_4217);
and U11109 (N_11109,N_2352,N_261);
nand U11110 (N_11110,N_5160,N_3446);
nor U11111 (N_11111,N_1193,N_3526);
nand U11112 (N_11112,N_154,N_5635);
nor U11113 (N_11113,N_1667,N_1254);
and U11114 (N_11114,N_3431,N_2513);
or U11115 (N_11115,N_1618,N_3038);
nor U11116 (N_11116,N_1974,N_4358);
nor U11117 (N_11117,N_2281,N_4433);
xnor U11118 (N_11118,N_122,N_2204);
nor U11119 (N_11119,N_5231,N_970);
xor U11120 (N_11120,N_3005,N_2587);
and U11121 (N_11121,N_263,N_1245);
nor U11122 (N_11122,N_5951,N_2514);
or U11123 (N_11123,N_1334,N_3985);
and U11124 (N_11124,N_1347,N_6081);
or U11125 (N_11125,N_3776,N_2405);
nor U11126 (N_11126,N_2154,N_4488);
or U11127 (N_11127,N_884,N_1043);
nand U11128 (N_11128,N_5269,N_2040);
nand U11129 (N_11129,N_3914,N_5644);
and U11130 (N_11130,N_1119,N_2527);
and U11131 (N_11131,N_1864,N_4103);
or U11132 (N_11132,N_5793,N_1526);
nor U11133 (N_11133,N_5545,N_715);
and U11134 (N_11134,N_2850,N_4813);
nand U11135 (N_11135,N_212,N_2415);
and U11136 (N_11136,N_2668,N_5767);
or U11137 (N_11137,N_842,N_4866);
nor U11138 (N_11138,N_5087,N_1506);
nor U11139 (N_11139,N_2191,N_5275);
and U11140 (N_11140,N_3613,N_3512);
or U11141 (N_11141,N_3612,N_2095);
nor U11142 (N_11142,N_2148,N_2841);
nand U11143 (N_11143,N_4162,N_3212);
nor U11144 (N_11144,N_761,N_1961);
nand U11145 (N_11145,N_3940,N_5054);
nor U11146 (N_11146,N_2642,N_3931);
nor U11147 (N_11147,N_607,N_2010);
nand U11148 (N_11148,N_624,N_2587);
nand U11149 (N_11149,N_103,N_5239);
and U11150 (N_11150,N_428,N_394);
xor U11151 (N_11151,N_3003,N_2736);
or U11152 (N_11152,N_278,N_2362);
xnor U11153 (N_11153,N_2914,N_5006);
nor U11154 (N_11154,N_5362,N_3675);
or U11155 (N_11155,N_115,N_3521);
nor U11156 (N_11156,N_89,N_613);
and U11157 (N_11157,N_3063,N_3269);
nand U11158 (N_11158,N_1976,N_4412);
xnor U11159 (N_11159,N_3761,N_123);
nand U11160 (N_11160,N_887,N_4025);
or U11161 (N_11161,N_446,N_1902);
or U11162 (N_11162,N_2055,N_5401);
nor U11163 (N_11163,N_2746,N_876);
or U11164 (N_11164,N_5416,N_763);
xor U11165 (N_11165,N_1040,N_212);
nor U11166 (N_11166,N_1552,N_5672);
or U11167 (N_11167,N_44,N_2551);
or U11168 (N_11168,N_2233,N_1745);
or U11169 (N_11169,N_1624,N_75);
nor U11170 (N_11170,N_5129,N_5705);
nand U11171 (N_11171,N_6159,N_4571);
xnor U11172 (N_11172,N_437,N_2374);
or U11173 (N_11173,N_3059,N_3262);
nand U11174 (N_11174,N_5973,N_904);
and U11175 (N_11175,N_4251,N_5956);
and U11176 (N_11176,N_5926,N_434);
nor U11177 (N_11177,N_1109,N_6187);
nor U11178 (N_11178,N_1287,N_3205);
and U11179 (N_11179,N_1807,N_5362);
nand U11180 (N_11180,N_4541,N_31);
nor U11181 (N_11181,N_5049,N_3968);
nor U11182 (N_11182,N_4858,N_1165);
and U11183 (N_11183,N_2397,N_5996);
and U11184 (N_11184,N_4774,N_6035);
nor U11185 (N_11185,N_2915,N_1392);
nand U11186 (N_11186,N_6002,N_1643);
and U11187 (N_11187,N_3060,N_507);
nor U11188 (N_11188,N_2337,N_1038);
or U11189 (N_11189,N_4858,N_3063);
or U11190 (N_11190,N_2213,N_3079);
or U11191 (N_11191,N_5874,N_3168);
and U11192 (N_11192,N_2884,N_2493);
and U11193 (N_11193,N_5193,N_309);
and U11194 (N_11194,N_2501,N_2756);
nor U11195 (N_11195,N_4731,N_3386);
and U11196 (N_11196,N_2845,N_553);
xor U11197 (N_11197,N_5950,N_4485);
and U11198 (N_11198,N_4861,N_3616);
nand U11199 (N_11199,N_5642,N_4960);
or U11200 (N_11200,N_2885,N_1457);
and U11201 (N_11201,N_5033,N_223);
and U11202 (N_11202,N_3148,N_4418);
nand U11203 (N_11203,N_1522,N_5136);
nor U11204 (N_11204,N_766,N_5120);
or U11205 (N_11205,N_1007,N_450);
nor U11206 (N_11206,N_537,N_2769);
xor U11207 (N_11207,N_631,N_2785);
or U11208 (N_11208,N_4150,N_1709);
nor U11209 (N_11209,N_415,N_4137);
or U11210 (N_11210,N_6028,N_1343);
or U11211 (N_11211,N_896,N_6116);
xnor U11212 (N_11212,N_1156,N_2556);
nor U11213 (N_11213,N_5589,N_2304);
xor U11214 (N_11214,N_4785,N_5761);
or U11215 (N_11215,N_2551,N_5663);
nor U11216 (N_11216,N_5248,N_4972);
or U11217 (N_11217,N_5408,N_2478);
and U11218 (N_11218,N_2755,N_1309);
nand U11219 (N_11219,N_2768,N_2897);
or U11220 (N_11220,N_1067,N_754);
xnor U11221 (N_11221,N_2043,N_3708);
and U11222 (N_11222,N_393,N_2058);
nor U11223 (N_11223,N_1784,N_5182);
nand U11224 (N_11224,N_1002,N_1433);
or U11225 (N_11225,N_3541,N_5373);
nand U11226 (N_11226,N_3863,N_5854);
or U11227 (N_11227,N_3397,N_3944);
nor U11228 (N_11228,N_4185,N_2573);
or U11229 (N_11229,N_3277,N_813);
nand U11230 (N_11230,N_4645,N_310);
or U11231 (N_11231,N_1526,N_4014);
and U11232 (N_11232,N_3166,N_1915);
and U11233 (N_11233,N_1481,N_1659);
nand U11234 (N_11234,N_1843,N_2323);
nand U11235 (N_11235,N_5212,N_5314);
xor U11236 (N_11236,N_1752,N_485);
nor U11237 (N_11237,N_6014,N_4289);
and U11238 (N_11238,N_1356,N_720);
or U11239 (N_11239,N_1111,N_3130);
nor U11240 (N_11240,N_4539,N_2424);
or U11241 (N_11241,N_482,N_3626);
nand U11242 (N_11242,N_6164,N_675);
or U11243 (N_11243,N_3349,N_1085);
or U11244 (N_11244,N_4093,N_5691);
and U11245 (N_11245,N_1957,N_3932);
or U11246 (N_11246,N_1026,N_1138);
or U11247 (N_11247,N_3758,N_2950);
and U11248 (N_11248,N_4722,N_1124);
nor U11249 (N_11249,N_2653,N_316);
or U11250 (N_11250,N_4306,N_1004);
nand U11251 (N_11251,N_4789,N_5450);
nor U11252 (N_11252,N_5686,N_6143);
nor U11253 (N_11253,N_4843,N_5493);
nand U11254 (N_11254,N_1534,N_4317);
nor U11255 (N_11255,N_1350,N_1467);
or U11256 (N_11256,N_294,N_1554);
and U11257 (N_11257,N_3834,N_1080);
and U11258 (N_11258,N_2131,N_430);
and U11259 (N_11259,N_2558,N_701);
nand U11260 (N_11260,N_1309,N_5314);
or U11261 (N_11261,N_2297,N_5144);
nor U11262 (N_11262,N_1176,N_4523);
nand U11263 (N_11263,N_2296,N_2182);
or U11264 (N_11264,N_1902,N_2671);
or U11265 (N_11265,N_3814,N_2020);
or U11266 (N_11266,N_1772,N_114);
nor U11267 (N_11267,N_2401,N_3308);
and U11268 (N_11268,N_3608,N_1942);
and U11269 (N_11269,N_2437,N_2558);
nor U11270 (N_11270,N_6044,N_2426);
xor U11271 (N_11271,N_503,N_3707);
nor U11272 (N_11272,N_1547,N_283);
or U11273 (N_11273,N_3218,N_3091);
nor U11274 (N_11274,N_4089,N_3894);
nand U11275 (N_11275,N_3395,N_5672);
nor U11276 (N_11276,N_4338,N_5064);
nor U11277 (N_11277,N_1184,N_547);
nand U11278 (N_11278,N_3055,N_5251);
and U11279 (N_11279,N_1699,N_3986);
or U11280 (N_11280,N_236,N_3543);
and U11281 (N_11281,N_4371,N_2387);
nand U11282 (N_11282,N_5444,N_2169);
or U11283 (N_11283,N_975,N_3247);
nand U11284 (N_11284,N_1465,N_4084);
nor U11285 (N_11285,N_241,N_5528);
nor U11286 (N_11286,N_2900,N_513);
nor U11287 (N_11287,N_1677,N_255);
and U11288 (N_11288,N_3816,N_3314);
and U11289 (N_11289,N_5920,N_1330);
and U11290 (N_11290,N_4343,N_5256);
or U11291 (N_11291,N_5098,N_3549);
nand U11292 (N_11292,N_2258,N_526);
nor U11293 (N_11293,N_2057,N_5360);
nand U11294 (N_11294,N_748,N_3466);
or U11295 (N_11295,N_3644,N_5289);
xnor U11296 (N_11296,N_4093,N_3732);
xor U11297 (N_11297,N_1717,N_1636);
nor U11298 (N_11298,N_10,N_934);
and U11299 (N_11299,N_1904,N_6215);
nor U11300 (N_11300,N_2125,N_1064);
or U11301 (N_11301,N_5624,N_2473);
nand U11302 (N_11302,N_1255,N_3849);
nor U11303 (N_11303,N_1274,N_1001);
nand U11304 (N_11304,N_4830,N_5806);
nor U11305 (N_11305,N_5744,N_923);
nor U11306 (N_11306,N_4888,N_3792);
nand U11307 (N_11307,N_4499,N_2628);
and U11308 (N_11308,N_3596,N_5869);
nand U11309 (N_11309,N_3269,N_652);
or U11310 (N_11310,N_2738,N_4867);
and U11311 (N_11311,N_4269,N_6043);
nor U11312 (N_11312,N_3639,N_1009);
and U11313 (N_11313,N_5044,N_3623);
nand U11314 (N_11314,N_3565,N_280);
nand U11315 (N_11315,N_1735,N_5941);
nor U11316 (N_11316,N_68,N_4388);
nand U11317 (N_11317,N_410,N_379);
nor U11318 (N_11318,N_2804,N_2155);
xor U11319 (N_11319,N_1373,N_4790);
and U11320 (N_11320,N_4346,N_814);
nor U11321 (N_11321,N_6061,N_2213);
nor U11322 (N_11322,N_1033,N_3265);
nor U11323 (N_11323,N_2494,N_592);
nand U11324 (N_11324,N_641,N_2567);
nor U11325 (N_11325,N_4790,N_2985);
or U11326 (N_11326,N_1673,N_5882);
xnor U11327 (N_11327,N_1173,N_5060);
or U11328 (N_11328,N_5524,N_1374);
or U11329 (N_11329,N_2853,N_1740);
nand U11330 (N_11330,N_637,N_532);
nand U11331 (N_11331,N_4250,N_4272);
and U11332 (N_11332,N_167,N_848);
xnor U11333 (N_11333,N_615,N_2197);
nand U11334 (N_11334,N_2269,N_3300);
and U11335 (N_11335,N_4267,N_1246);
nor U11336 (N_11336,N_4235,N_2907);
nand U11337 (N_11337,N_2570,N_5800);
or U11338 (N_11338,N_3132,N_840);
xor U11339 (N_11339,N_3551,N_4435);
and U11340 (N_11340,N_22,N_3823);
or U11341 (N_11341,N_3653,N_3060);
nor U11342 (N_11342,N_923,N_2516);
and U11343 (N_11343,N_3710,N_1185);
nand U11344 (N_11344,N_545,N_5440);
and U11345 (N_11345,N_2972,N_6049);
nor U11346 (N_11346,N_4944,N_3088);
nand U11347 (N_11347,N_6165,N_5753);
and U11348 (N_11348,N_955,N_3025);
or U11349 (N_11349,N_1857,N_5463);
and U11350 (N_11350,N_2801,N_2396);
nand U11351 (N_11351,N_388,N_74);
or U11352 (N_11352,N_2362,N_3575);
nor U11353 (N_11353,N_2391,N_2291);
or U11354 (N_11354,N_5278,N_2756);
nand U11355 (N_11355,N_939,N_5232);
or U11356 (N_11356,N_3050,N_1497);
nor U11357 (N_11357,N_2818,N_4120);
nand U11358 (N_11358,N_4951,N_1703);
xor U11359 (N_11359,N_5511,N_2100);
xor U11360 (N_11360,N_4592,N_4783);
and U11361 (N_11361,N_3755,N_325);
nand U11362 (N_11362,N_4948,N_2710);
or U11363 (N_11363,N_6013,N_4343);
and U11364 (N_11364,N_4145,N_286);
nand U11365 (N_11365,N_5221,N_3701);
or U11366 (N_11366,N_1931,N_856);
nor U11367 (N_11367,N_267,N_4693);
nand U11368 (N_11368,N_188,N_6244);
or U11369 (N_11369,N_3195,N_4690);
and U11370 (N_11370,N_3164,N_948);
or U11371 (N_11371,N_2821,N_1199);
nor U11372 (N_11372,N_3382,N_4778);
or U11373 (N_11373,N_2413,N_3895);
and U11374 (N_11374,N_381,N_1540);
and U11375 (N_11375,N_4751,N_2333);
or U11376 (N_11376,N_5363,N_6184);
nand U11377 (N_11377,N_2373,N_5756);
and U11378 (N_11378,N_5267,N_4620);
xnor U11379 (N_11379,N_3010,N_81);
nor U11380 (N_11380,N_6040,N_6192);
nor U11381 (N_11381,N_884,N_5290);
and U11382 (N_11382,N_3057,N_1460);
xnor U11383 (N_11383,N_366,N_2815);
nand U11384 (N_11384,N_1273,N_3072);
xor U11385 (N_11385,N_477,N_5846);
nor U11386 (N_11386,N_4283,N_3545);
nor U11387 (N_11387,N_2639,N_2961);
xnor U11388 (N_11388,N_1267,N_1754);
nor U11389 (N_11389,N_6192,N_3292);
nor U11390 (N_11390,N_3498,N_5947);
and U11391 (N_11391,N_3758,N_3451);
or U11392 (N_11392,N_1236,N_1391);
nand U11393 (N_11393,N_6126,N_3114);
nand U11394 (N_11394,N_5217,N_1840);
or U11395 (N_11395,N_5199,N_4132);
nor U11396 (N_11396,N_3763,N_4998);
nand U11397 (N_11397,N_113,N_636);
xnor U11398 (N_11398,N_1636,N_3550);
or U11399 (N_11399,N_4091,N_1466);
or U11400 (N_11400,N_2516,N_3934);
nand U11401 (N_11401,N_3374,N_5662);
nand U11402 (N_11402,N_2753,N_2215);
nand U11403 (N_11403,N_1257,N_312);
xnor U11404 (N_11404,N_2999,N_660);
nand U11405 (N_11405,N_2442,N_5784);
nor U11406 (N_11406,N_3609,N_425);
nor U11407 (N_11407,N_5054,N_697);
or U11408 (N_11408,N_4640,N_1197);
nand U11409 (N_11409,N_1369,N_5231);
or U11410 (N_11410,N_3313,N_6160);
and U11411 (N_11411,N_1770,N_4990);
or U11412 (N_11412,N_3199,N_4186);
and U11413 (N_11413,N_2127,N_5244);
or U11414 (N_11414,N_3755,N_772);
nand U11415 (N_11415,N_3082,N_2312);
or U11416 (N_11416,N_1402,N_3868);
xnor U11417 (N_11417,N_743,N_5694);
xnor U11418 (N_11418,N_262,N_3448);
and U11419 (N_11419,N_6231,N_5878);
nand U11420 (N_11420,N_1930,N_5021);
nor U11421 (N_11421,N_1668,N_2746);
nand U11422 (N_11422,N_5985,N_3572);
or U11423 (N_11423,N_1270,N_1719);
nand U11424 (N_11424,N_3163,N_3442);
and U11425 (N_11425,N_3698,N_4858);
and U11426 (N_11426,N_3921,N_5632);
nand U11427 (N_11427,N_1133,N_740);
or U11428 (N_11428,N_1159,N_1438);
and U11429 (N_11429,N_2352,N_575);
nand U11430 (N_11430,N_3569,N_6000);
nand U11431 (N_11431,N_3823,N_3470);
xor U11432 (N_11432,N_919,N_3820);
nand U11433 (N_11433,N_1167,N_3267);
xor U11434 (N_11434,N_389,N_2618);
nor U11435 (N_11435,N_4250,N_5744);
and U11436 (N_11436,N_5756,N_4917);
nand U11437 (N_11437,N_4574,N_1229);
nor U11438 (N_11438,N_5609,N_4954);
nand U11439 (N_11439,N_4211,N_3724);
nor U11440 (N_11440,N_3281,N_2844);
nor U11441 (N_11441,N_153,N_2256);
nand U11442 (N_11442,N_5694,N_4208);
or U11443 (N_11443,N_4100,N_2797);
and U11444 (N_11444,N_3017,N_727);
nor U11445 (N_11445,N_3612,N_3722);
or U11446 (N_11446,N_3049,N_4794);
and U11447 (N_11447,N_3035,N_1195);
nand U11448 (N_11448,N_2117,N_5438);
nand U11449 (N_11449,N_4811,N_609);
nand U11450 (N_11450,N_4592,N_669);
and U11451 (N_11451,N_5176,N_485);
xnor U11452 (N_11452,N_3077,N_798);
xor U11453 (N_11453,N_5925,N_1747);
and U11454 (N_11454,N_6158,N_1671);
and U11455 (N_11455,N_313,N_5504);
nand U11456 (N_11456,N_124,N_2196);
nand U11457 (N_11457,N_3015,N_1759);
nand U11458 (N_11458,N_3843,N_3245);
nand U11459 (N_11459,N_1039,N_5117);
nor U11460 (N_11460,N_1491,N_202);
and U11461 (N_11461,N_5710,N_811);
nor U11462 (N_11462,N_4442,N_451);
xnor U11463 (N_11463,N_5490,N_75);
nor U11464 (N_11464,N_5381,N_636);
nand U11465 (N_11465,N_1417,N_3291);
and U11466 (N_11466,N_2089,N_2631);
nor U11467 (N_11467,N_2577,N_1552);
xor U11468 (N_11468,N_1350,N_2559);
nor U11469 (N_11469,N_5152,N_1856);
or U11470 (N_11470,N_5983,N_364);
nand U11471 (N_11471,N_3545,N_3342);
nor U11472 (N_11472,N_6028,N_5261);
xnor U11473 (N_11473,N_3487,N_3687);
or U11474 (N_11474,N_4150,N_404);
xor U11475 (N_11475,N_5072,N_320);
nand U11476 (N_11476,N_1680,N_3217);
nor U11477 (N_11477,N_5007,N_617);
nand U11478 (N_11478,N_3030,N_725);
nor U11479 (N_11479,N_3928,N_2039);
nand U11480 (N_11480,N_462,N_4130);
xor U11481 (N_11481,N_1299,N_1822);
nand U11482 (N_11482,N_5949,N_995);
and U11483 (N_11483,N_4906,N_2794);
or U11484 (N_11484,N_1927,N_431);
nor U11485 (N_11485,N_4404,N_5984);
and U11486 (N_11486,N_3453,N_1412);
nor U11487 (N_11487,N_4752,N_2088);
or U11488 (N_11488,N_1953,N_3808);
nand U11489 (N_11489,N_4108,N_4554);
nor U11490 (N_11490,N_516,N_1465);
xnor U11491 (N_11491,N_5120,N_4858);
xor U11492 (N_11492,N_2929,N_4099);
or U11493 (N_11493,N_679,N_3135);
or U11494 (N_11494,N_5018,N_1518);
nand U11495 (N_11495,N_856,N_2592);
and U11496 (N_11496,N_1080,N_3826);
or U11497 (N_11497,N_803,N_1290);
or U11498 (N_11498,N_5558,N_2192);
xor U11499 (N_11499,N_3396,N_2845);
nand U11500 (N_11500,N_2494,N_4588);
nand U11501 (N_11501,N_862,N_5700);
xor U11502 (N_11502,N_389,N_3675);
and U11503 (N_11503,N_6115,N_55);
and U11504 (N_11504,N_5637,N_3457);
or U11505 (N_11505,N_1730,N_1659);
nand U11506 (N_11506,N_5308,N_2439);
nand U11507 (N_11507,N_3580,N_4290);
nand U11508 (N_11508,N_1846,N_6078);
nor U11509 (N_11509,N_1088,N_5541);
or U11510 (N_11510,N_3254,N_4562);
and U11511 (N_11511,N_4888,N_2129);
nand U11512 (N_11512,N_5023,N_5232);
or U11513 (N_11513,N_1314,N_2155);
nor U11514 (N_11514,N_105,N_5499);
nand U11515 (N_11515,N_5799,N_3728);
nor U11516 (N_11516,N_3442,N_3688);
or U11517 (N_11517,N_387,N_5878);
and U11518 (N_11518,N_5847,N_404);
xor U11519 (N_11519,N_5259,N_4262);
nand U11520 (N_11520,N_2288,N_3188);
nand U11521 (N_11521,N_3136,N_2828);
nor U11522 (N_11522,N_2538,N_1896);
nand U11523 (N_11523,N_3055,N_1869);
nor U11524 (N_11524,N_2317,N_2236);
nand U11525 (N_11525,N_5894,N_3376);
xnor U11526 (N_11526,N_3619,N_3854);
or U11527 (N_11527,N_3678,N_2882);
or U11528 (N_11528,N_1008,N_5406);
nor U11529 (N_11529,N_5569,N_1714);
xor U11530 (N_11530,N_2228,N_1674);
or U11531 (N_11531,N_3966,N_1177);
nand U11532 (N_11532,N_721,N_5134);
nand U11533 (N_11533,N_5718,N_3634);
or U11534 (N_11534,N_5565,N_2);
nand U11535 (N_11535,N_2934,N_2606);
and U11536 (N_11536,N_5727,N_3993);
and U11537 (N_11537,N_3466,N_4108);
nand U11538 (N_11538,N_5357,N_2740);
and U11539 (N_11539,N_3279,N_6231);
and U11540 (N_11540,N_4655,N_2467);
nor U11541 (N_11541,N_4457,N_5701);
and U11542 (N_11542,N_6238,N_3597);
xor U11543 (N_11543,N_2335,N_1570);
nand U11544 (N_11544,N_6216,N_4717);
and U11545 (N_11545,N_3190,N_5555);
or U11546 (N_11546,N_2561,N_5891);
nand U11547 (N_11547,N_3345,N_2962);
and U11548 (N_11548,N_3444,N_4787);
nand U11549 (N_11549,N_1065,N_1968);
and U11550 (N_11550,N_995,N_4074);
nor U11551 (N_11551,N_4187,N_3781);
nor U11552 (N_11552,N_4159,N_3241);
xor U11553 (N_11553,N_2697,N_2125);
and U11554 (N_11554,N_6184,N_5923);
nand U11555 (N_11555,N_843,N_5000);
nor U11556 (N_11556,N_1862,N_1477);
and U11557 (N_11557,N_4543,N_3427);
and U11558 (N_11558,N_3789,N_2163);
or U11559 (N_11559,N_4569,N_1462);
nand U11560 (N_11560,N_2564,N_2162);
and U11561 (N_11561,N_81,N_2924);
nand U11562 (N_11562,N_4800,N_3440);
nor U11563 (N_11563,N_1350,N_2332);
xnor U11564 (N_11564,N_2559,N_3789);
and U11565 (N_11565,N_337,N_1800);
or U11566 (N_11566,N_4290,N_725);
or U11567 (N_11567,N_6115,N_3803);
xor U11568 (N_11568,N_5255,N_1585);
nand U11569 (N_11569,N_464,N_6207);
nor U11570 (N_11570,N_2533,N_4109);
or U11571 (N_11571,N_1593,N_2699);
and U11572 (N_11572,N_5876,N_6027);
or U11573 (N_11573,N_4803,N_881);
nor U11574 (N_11574,N_3293,N_1177);
and U11575 (N_11575,N_2170,N_1729);
xnor U11576 (N_11576,N_1605,N_409);
or U11577 (N_11577,N_5610,N_4513);
or U11578 (N_11578,N_1079,N_5555);
nand U11579 (N_11579,N_3663,N_983);
xor U11580 (N_11580,N_2849,N_2907);
or U11581 (N_11581,N_5255,N_2203);
xnor U11582 (N_11582,N_1154,N_2042);
nand U11583 (N_11583,N_578,N_5001);
nand U11584 (N_11584,N_5732,N_890);
nand U11585 (N_11585,N_4644,N_1239);
or U11586 (N_11586,N_28,N_1097);
or U11587 (N_11587,N_708,N_3737);
or U11588 (N_11588,N_2737,N_5203);
nand U11589 (N_11589,N_2765,N_1231);
or U11590 (N_11590,N_3819,N_5485);
nand U11591 (N_11591,N_5558,N_904);
xor U11592 (N_11592,N_2365,N_6054);
and U11593 (N_11593,N_1774,N_2485);
or U11594 (N_11594,N_6136,N_4337);
xnor U11595 (N_11595,N_1323,N_2901);
nor U11596 (N_11596,N_456,N_2356);
and U11597 (N_11597,N_943,N_733);
and U11598 (N_11598,N_3543,N_5324);
and U11599 (N_11599,N_2318,N_2508);
nand U11600 (N_11600,N_4226,N_5953);
and U11601 (N_11601,N_201,N_2176);
or U11602 (N_11602,N_3743,N_430);
and U11603 (N_11603,N_2271,N_325);
nor U11604 (N_11604,N_1062,N_1377);
nand U11605 (N_11605,N_2540,N_4214);
or U11606 (N_11606,N_322,N_2777);
nor U11607 (N_11607,N_4373,N_3778);
nand U11608 (N_11608,N_4480,N_5298);
nand U11609 (N_11609,N_5878,N_4639);
or U11610 (N_11610,N_3854,N_3959);
nor U11611 (N_11611,N_5346,N_2263);
nand U11612 (N_11612,N_5007,N_2901);
nor U11613 (N_11613,N_5908,N_2467);
and U11614 (N_11614,N_133,N_3837);
or U11615 (N_11615,N_5445,N_5094);
and U11616 (N_11616,N_2176,N_2961);
and U11617 (N_11617,N_924,N_2610);
xor U11618 (N_11618,N_1788,N_4061);
or U11619 (N_11619,N_1549,N_5190);
nand U11620 (N_11620,N_201,N_4876);
and U11621 (N_11621,N_3393,N_4891);
or U11622 (N_11622,N_652,N_2665);
nor U11623 (N_11623,N_4626,N_2013);
nand U11624 (N_11624,N_3186,N_2087);
or U11625 (N_11625,N_5629,N_6051);
nand U11626 (N_11626,N_2173,N_3467);
or U11627 (N_11627,N_3678,N_170);
and U11628 (N_11628,N_1418,N_5083);
xor U11629 (N_11629,N_1152,N_2169);
and U11630 (N_11630,N_2095,N_5361);
and U11631 (N_11631,N_3638,N_219);
nor U11632 (N_11632,N_4070,N_1410);
or U11633 (N_11633,N_3207,N_4193);
nand U11634 (N_11634,N_3234,N_1266);
nor U11635 (N_11635,N_2419,N_530);
nand U11636 (N_11636,N_827,N_1450);
and U11637 (N_11637,N_5008,N_4745);
nor U11638 (N_11638,N_3597,N_5788);
or U11639 (N_11639,N_445,N_5222);
or U11640 (N_11640,N_2172,N_444);
and U11641 (N_11641,N_4397,N_4009);
and U11642 (N_11642,N_4701,N_2124);
nor U11643 (N_11643,N_5134,N_3200);
and U11644 (N_11644,N_106,N_5895);
or U11645 (N_11645,N_743,N_4572);
nand U11646 (N_11646,N_3329,N_1243);
xnor U11647 (N_11647,N_1403,N_519);
and U11648 (N_11648,N_4840,N_2486);
nand U11649 (N_11649,N_430,N_4943);
nor U11650 (N_11650,N_4396,N_4229);
and U11651 (N_11651,N_5717,N_5183);
nor U11652 (N_11652,N_205,N_3536);
or U11653 (N_11653,N_5744,N_1261);
nor U11654 (N_11654,N_409,N_1874);
or U11655 (N_11655,N_5972,N_1689);
nand U11656 (N_11656,N_345,N_1144);
xor U11657 (N_11657,N_4976,N_5305);
xor U11658 (N_11658,N_4868,N_6240);
nor U11659 (N_11659,N_4218,N_777);
nor U11660 (N_11660,N_4314,N_3951);
xor U11661 (N_11661,N_4634,N_4839);
or U11662 (N_11662,N_689,N_2951);
nand U11663 (N_11663,N_3900,N_2657);
or U11664 (N_11664,N_4212,N_4964);
and U11665 (N_11665,N_3424,N_335);
or U11666 (N_11666,N_3449,N_1637);
xnor U11667 (N_11667,N_4285,N_4820);
nor U11668 (N_11668,N_5217,N_5664);
or U11669 (N_11669,N_2398,N_1643);
or U11670 (N_11670,N_3116,N_1780);
nor U11671 (N_11671,N_619,N_474);
nand U11672 (N_11672,N_4310,N_3729);
nor U11673 (N_11673,N_5415,N_1195);
xor U11674 (N_11674,N_2466,N_979);
xnor U11675 (N_11675,N_2019,N_1381);
or U11676 (N_11676,N_5261,N_1912);
or U11677 (N_11677,N_4821,N_1193);
xnor U11678 (N_11678,N_5906,N_22);
nor U11679 (N_11679,N_5778,N_860);
nand U11680 (N_11680,N_5140,N_4637);
and U11681 (N_11681,N_2422,N_258);
nor U11682 (N_11682,N_4101,N_5528);
nor U11683 (N_11683,N_1734,N_1981);
and U11684 (N_11684,N_3813,N_6040);
nand U11685 (N_11685,N_37,N_2245);
nand U11686 (N_11686,N_677,N_2152);
and U11687 (N_11687,N_5143,N_677);
nand U11688 (N_11688,N_4343,N_4884);
nor U11689 (N_11689,N_4503,N_5563);
nor U11690 (N_11690,N_376,N_4690);
or U11691 (N_11691,N_4445,N_990);
xnor U11692 (N_11692,N_6224,N_4913);
or U11693 (N_11693,N_2841,N_3944);
xor U11694 (N_11694,N_4815,N_4935);
or U11695 (N_11695,N_5894,N_978);
nor U11696 (N_11696,N_966,N_6042);
and U11697 (N_11697,N_245,N_467);
nand U11698 (N_11698,N_6097,N_1464);
nor U11699 (N_11699,N_5485,N_1920);
nor U11700 (N_11700,N_4159,N_1585);
and U11701 (N_11701,N_464,N_2981);
or U11702 (N_11702,N_3145,N_397);
nor U11703 (N_11703,N_3365,N_93);
or U11704 (N_11704,N_1650,N_2955);
nand U11705 (N_11705,N_5351,N_3781);
xor U11706 (N_11706,N_1371,N_1963);
nand U11707 (N_11707,N_1885,N_4680);
nand U11708 (N_11708,N_1745,N_569);
nor U11709 (N_11709,N_2710,N_4416);
nand U11710 (N_11710,N_5073,N_3645);
or U11711 (N_11711,N_2460,N_4356);
nand U11712 (N_11712,N_3323,N_4286);
or U11713 (N_11713,N_5586,N_923);
and U11714 (N_11714,N_3932,N_2253);
nor U11715 (N_11715,N_3449,N_413);
and U11716 (N_11716,N_3387,N_5330);
nand U11717 (N_11717,N_5657,N_3253);
nand U11718 (N_11718,N_3903,N_989);
nor U11719 (N_11719,N_5932,N_4156);
nand U11720 (N_11720,N_350,N_2317);
or U11721 (N_11721,N_1201,N_6237);
and U11722 (N_11722,N_724,N_189);
xnor U11723 (N_11723,N_2595,N_142);
or U11724 (N_11724,N_2939,N_4918);
nor U11725 (N_11725,N_3780,N_5831);
or U11726 (N_11726,N_3634,N_3389);
nor U11727 (N_11727,N_5399,N_4428);
or U11728 (N_11728,N_436,N_293);
nor U11729 (N_11729,N_3146,N_5117);
and U11730 (N_11730,N_2245,N_1897);
nor U11731 (N_11731,N_1296,N_3680);
and U11732 (N_11732,N_5574,N_4957);
and U11733 (N_11733,N_6160,N_2568);
xnor U11734 (N_11734,N_1171,N_1887);
or U11735 (N_11735,N_2091,N_2133);
nor U11736 (N_11736,N_3370,N_2018);
nand U11737 (N_11737,N_4327,N_1801);
nor U11738 (N_11738,N_5242,N_5231);
xor U11739 (N_11739,N_1101,N_4706);
nand U11740 (N_11740,N_2386,N_1917);
and U11741 (N_11741,N_1862,N_3771);
xor U11742 (N_11742,N_4068,N_1584);
xor U11743 (N_11743,N_416,N_520);
and U11744 (N_11744,N_295,N_1689);
or U11745 (N_11745,N_295,N_4036);
nor U11746 (N_11746,N_4207,N_6022);
nor U11747 (N_11747,N_2088,N_758);
nand U11748 (N_11748,N_6209,N_3011);
or U11749 (N_11749,N_2348,N_1504);
and U11750 (N_11750,N_2930,N_6043);
nand U11751 (N_11751,N_865,N_4590);
and U11752 (N_11752,N_973,N_5401);
and U11753 (N_11753,N_2306,N_3298);
xor U11754 (N_11754,N_3678,N_5127);
and U11755 (N_11755,N_1125,N_1343);
and U11756 (N_11756,N_611,N_5926);
or U11757 (N_11757,N_2855,N_4920);
nor U11758 (N_11758,N_896,N_1934);
nor U11759 (N_11759,N_1949,N_910);
or U11760 (N_11760,N_4987,N_4447);
nand U11761 (N_11761,N_1158,N_5621);
nor U11762 (N_11762,N_3622,N_4615);
nor U11763 (N_11763,N_4668,N_1695);
nand U11764 (N_11764,N_3585,N_1350);
and U11765 (N_11765,N_1857,N_4119);
nand U11766 (N_11766,N_6014,N_920);
and U11767 (N_11767,N_2151,N_1485);
xnor U11768 (N_11768,N_4076,N_475);
nor U11769 (N_11769,N_2492,N_5965);
nor U11770 (N_11770,N_839,N_103);
nor U11771 (N_11771,N_6203,N_4330);
or U11772 (N_11772,N_3420,N_5025);
and U11773 (N_11773,N_1565,N_5509);
or U11774 (N_11774,N_3234,N_3548);
nor U11775 (N_11775,N_2265,N_4176);
xnor U11776 (N_11776,N_4852,N_4376);
nor U11777 (N_11777,N_4918,N_6038);
nand U11778 (N_11778,N_3661,N_2451);
nor U11779 (N_11779,N_3027,N_568);
or U11780 (N_11780,N_4134,N_595);
or U11781 (N_11781,N_4046,N_5899);
or U11782 (N_11782,N_5072,N_5295);
or U11783 (N_11783,N_4102,N_3173);
nor U11784 (N_11784,N_1110,N_549);
nor U11785 (N_11785,N_4663,N_2981);
xnor U11786 (N_11786,N_4851,N_2585);
nand U11787 (N_11787,N_6011,N_2678);
and U11788 (N_11788,N_2384,N_4027);
or U11789 (N_11789,N_5621,N_2527);
and U11790 (N_11790,N_3528,N_1493);
nor U11791 (N_11791,N_937,N_1944);
and U11792 (N_11792,N_2289,N_5467);
nand U11793 (N_11793,N_752,N_3266);
and U11794 (N_11794,N_4423,N_5299);
nand U11795 (N_11795,N_1948,N_4566);
nand U11796 (N_11796,N_2179,N_1240);
nand U11797 (N_11797,N_1220,N_3767);
or U11798 (N_11798,N_1688,N_5140);
nand U11799 (N_11799,N_4912,N_2244);
and U11800 (N_11800,N_6176,N_5361);
or U11801 (N_11801,N_5900,N_1251);
nor U11802 (N_11802,N_1250,N_4494);
nor U11803 (N_11803,N_4337,N_5885);
nor U11804 (N_11804,N_5453,N_3098);
nand U11805 (N_11805,N_4154,N_3959);
nand U11806 (N_11806,N_3111,N_5052);
or U11807 (N_11807,N_431,N_5950);
and U11808 (N_11808,N_3286,N_317);
and U11809 (N_11809,N_2825,N_6246);
nor U11810 (N_11810,N_2543,N_6210);
nand U11811 (N_11811,N_3806,N_3078);
nand U11812 (N_11812,N_5133,N_6142);
or U11813 (N_11813,N_1263,N_2448);
nand U11814 (N_11814,N_5807,N_4181);
nand U11815 (N_11815,N_6019,N_1897);
and U11816 (N_11816,N_656,N_6212);
nor U11817 (N_11817,N_5547,N_557);
nor U11818 (N_11818,N_871,N_569);
and U11819 (N_11819,N_1895,N_4998);
xnor U11820 (N_11820,N_4507,N_487);
nor U11821 (N_11821,N_5005,N_5321);
nor U11822 (N_11822,N_4635,N_2437);
or U11823 (N_11823,N_2500,N_1695);
nand U11824 (N_11824,N_4850,N_2691);
nand U11825 (N_11825,N_1241,N_5202);
xor U11826 (N_11826,N_6104,N_403);
and U11827 (N_11827,N_1586,N_5886);
or U11828 (N_11828,N_3889,N_3169);
and U11829 (N_11829,N_4361,N_4431);
nor U11830 (N_11830,N_4232,N_3560);
nor U11831 (N_11831,N_591,N_4104);
and U11832 (N_11832,N_1376,N_1955);
and U11833 (N_11833,N_4970,N_3580);
xnor U11834 (N_11834,N_1312,N_3525);
nand U11835 (N_11835,N_2458,N_1239);
and U11836 (N_11836,N_5628,N_6093);
xnor U11837 (N_11837,N_837,N_3947);
and U11838 (N_11838,N_5960,N_5491);
nand U11839 (N_11839,N_1514,N_2798);
nand U11840 (N_11840,N_897,N_2756);
or U11841 (N_11841,N_4746,N_2989);
xnor U11842 (N_11842,N_4535,N_4683);
and U11843 (N_11843,N_1048,N_2807);
xor U11844 (N_11844,N_1624,N_919);
and U11845 (N_11845,N_1842,N_673);
and U11846 (N_11846,N_4129,N_2618);
nor U11847 (N_11847,N_3827,N_2710);
nor U11848 (N_11848,N_4780,N_2134);
nor U11849 (N_11849,N_4105,N_2404);
nand U11850 (N_11850,N_4085,N_4753);
nand U11851 (N_11851,N_4059,N_5303);
or U11852 (N_11852,N_6112,N_1642);
xnor U11853 (N_11853,N_4615,N_4971);
nand U11854 (N_11854,N_2222,N_2201);
nor U11855 (N_11855,N_3617,N_3219);
nand U11856 (N_11856,N_2377,N_4552);
nand U11857 (N_11857,N_5378,N_5598);
xnor U11858 (N_11858,N_5887,N_870);
nor U11859 (N_11859,N_3783,N_1879);
xnor U11860 (N_11860,N_5851,N_112);
nand U11861 (N_11861,N_721,N_4111);
nand U11862 (N_11862,N_3089,N_3747);
or U11863 (N_11863,N_2828,N_3814);
nand U11864 (N_11864,N_6068,N_5427);
nand U11865 (N_11865,N_1680,N_4477);
nand U11866 (N_11866,N_4094,N_3744);
or U11867 (N_11867,N_2246,N_5406);
or U11868 (N_11868,N_4907,N_2554);
or U11869 (N_11869,N_1249,N_587);
nor U11870 (N_11870,N_5709,N_2339);
nor U11871 (N_11871,N_3921,N_3429);
and U11872 (N_11872,N_2124,N_4945);
nor U11873 (N_11873,N_2147,N_5205);
nand U11874 (N_11874,N_3768,N_2032);
xnor U11875 (N_11875,N_619,N_1340);
nor U11876 (N_11876,N_4873,N_5302);
or U11877 (N_11877,N_4249,N_1654);
nor U11878 (N_11878,N_5771,N_1783);
nor U11879 (N_11879,N_2580,N_6171);
nand U11880 (N_11880,N_1312,N_1522);
nor U11881 (N_11881,N_3252,N_2258);
and U11882 (N_11882,N_3335,N_2149);
xor U11883 (N_11883,N_3344,N_2243);
or U11884 (N_11884,N_1921,N_125);
or U11885 (N_11885,N_4937,N_2817);
xnor U11886 (N_11886,N_5365,N_6213);
or U11887 (N_11887,N_5793,N_2355);
and U11888 (N_11888,N_1262,N_880);
nand U11889 (N_11889,N_5030,N_260);
and U11890 (N_11890,N_5955,N_2693);
xnor U11891 (N_11891,N_5394,N_5158);
and U11892 (N_11892,N_5304,N_925);
nor U11893 (N_11893,N_5309,N_857);
or U11894 (N_11894,N_5466,N_5685);
nor U11895 (N_11895,N_3035,N_1543);
and U11896 (N_11896,N_5650,N_1820);
nand U11897 (N_11897,N_647,N_5369);
xnor U11898 (N_11898,N_767,N_1490);
nor U11899 (N_11899,N_6018,N_5044);
and U11900 (N_11900,N_1431,N_4571);
nor U11901 (N_11901,N_4824,N_2700);
or U11902 (N_11902,N_5696,N_5347);
and U11903 (N_11903,N_1268,N_3673);
or U11904 (N_11904,N_4279,N_1427);
nand U11905 (N_11905,N_5606,N_4652);
xnor U11906 (N_11906,N_1545,N_895);
or U11907 (N_11907,N_1490,N_645);
nor U11908 (N_11908,N_5279,N_5785);
and U11909 (N_11909,N_4381,N_4488);
nor U11910 (N_11910,N_4156,N_2913);
and U11911 (N_11911,N_1995,N_2674);
or U11912 (N_11912,N_745,N_2508);
and U11913 (N_11913,N_5317,N_4126);
nand U11914 (N_11914,N_5349,N_896);
nand U11915 (N_11915,N_2130,N_6234);
xnor U11916 (N_11916,N_5990,N_1601);
xnor U11917 (N_11917,N_3176,N_4940);
nor U11918 (N_11918,N_3792,N_3337);
nand U11919 (N_11919,N_5428,N_3191);
nand U11920 (N_11920,N_718,N_2869);
nand U11921 (N_11921,N_6074,N_3547);
nor U11922 (N_11922,N_2793,N_1307);
or U11923 (N_11923,N_1482,N_1147);
nor U11924 (N_11924,N_122,N_6043);
nand U11925 (N_11925,N_2207,N_1987);
nand U11926 (N_11926,N_4891,N_1937);
and U11927 (N_11927,N_5927,N_1575);
and U11928 (N_11928,N_2590,N_5485);
xor U11929 (N_11929,N_3714,N_1660);
and U11930 (N_11930,N_5783,N_909);
nor U11931 (N_11931,N_2270,N_1846);
or U11932 (N_11932,N_213,N_347);
nor U11933 (N_11933,N_4857,N_1706);
nand U11934 (N_11934,N_4474,N_4244);
xnor U11935 (N_11935,N_1962,N_3502);
or U11936 (N_11936,N_5076,N_5063);
or U11937 (N_11937,N_1388,N_2152);
or U11938 (N_11938,N_5113,N_1247);
nor U11939 (N_11939,N_432,N_2017);
nor U11940 (N_11940,N_3906,N_728);
or U11941 (N_11941,N_2391,N_5318);
or U11942 (N_11942,N_718,N_1322);
xnor U11943 (N_11943,N_1737,N_1213);
nor U11944 (N_11944,N_2365,N_824);
nand U11945 (N_11945,N_2146,N_5042);
and U11946 (N_11946,N_3767,N_5783);
nand U11947 (N_11947,N_4616,N_4777);
and U11948 (N_11948,N_4704,N_5581);
or U11949 (N_11949,N_1449,N_698);
or U11950 (N_11950,N_4698,N_3133);
nand U11951 (N_11951,N_5685,N_4653);
nand U11952 (N_11952,N_3656,N_5127);
nor U11953 (N_11953,N_2931,N_1024);
or U11954 (N_11954,N_3100,N_5659);
or U11955 (N_11955,N_2339,N_4013);
and U11956 (N_11956,N_5104,N_329);
and U11957 (N_11957,N_5757,N_5321);
and U11958 (N_11958,N_4181,N_2800);
nor U11959 (N_11959,N_4429,N_1291);
or U11960 (N_11960,N_6197,N_3512);
nand U11961 (N_11961,N_5371,N_1056);
and U11962 (N_11962,N_2077,N_928);
nor U11963 (N_11963,N_1271,N_5823);
or U11964 (N_11964,N_3448,N_2070);
or U11965 (N_11965,N_100,N_4196);
xnor U11966 (N_11966,N_3918,N_5151);
and U11967 (N_11967,N_1114,N_3071);
nor U11968 (N_11968,N_4192,N_4041);
and U11969 (N_11969,N_2862,N_3168);
nand U11970 (N_11970,N_723,N_2639);
and U11971 (N_11971,N_5338,N_5372);
or U11972 (N_11972,N_4672,N_1359);
xor U11973 (N_11973,N_2300,N_5456);
nand U11974 (N_11974,N_2921,N_3635);
and U11975 (N_11975,N_891,N_1346);
nand U11976 (N_11976,N_1629,N_2925);
and U11977 (N_11977,N_4785,N_3684);
and U11978 (N_11978,N_201,N_2949);
xnor U11979 (N_11979,N_3126,N_1850);
nand U11980 (N_11980,N_6124,N_268);
nand U11981 (N_11981,N_1630,N_322);
and U11982 (N_11982,N_4076,N_5469);
and U11983 (N_11983,N_4931,N_2204);
nor U11984 (N_11984,N_5801,N_19);
or U11985 (N_11985,N_2989,N_2813);
nand U11986 (N_11986,N_936,N_5520);
and U11987 (N_11987,N_5682,N_3296);
or U11988 (N_11988,N_948,N_5044);
nor U11989 (N_11989,N_5398,N_3988);
nor U11990 (N_11990,N_3346,N_5844);
nand U11991 (N_11991,N_2710,N_3703);
xnor U11992 (N_11992,N_4674,N_3166);
or U11993 (N_11993,N_5378,N_809);
and U11994 (N_11994,N_1650,N_5784);
nand U11995 (N_11995,N_2769,N_4367);
nand U11996 (N_11996,N_2970,N_2460);
nor U11997 (N_11997,N_1096,N_4801);
and U11998 (N_11998,N_1045,N_3103);
nand U11999 (N_11999,N_1861,N_304);
nor U12000 (N_12000,N_4424,N_2782);
or U12001 (N_12001,N_4373,N_2640);
and U12002 (N_12002,N_3417,N_3516);
and U12003 (N_12003,N_3556,N_4464);
or U12004 (N_12004,N_2811,N_3593);
and U12005 (N_12005,N_5230,N_4476);
and U12006 (N_12006,N_4274,N_4679);
nand U12007 (N_12007,N_4122,N_3725);
and U12008 (N_12008,N_180,N_5991);
xnor U12009 (N_12009,N_538,N_798);
and U12010 (N_12010,N_951,N_3032);
or U12011 (N_12011,N_4052,N_3842);
nand U12012 (N_12012,N_2298,N_1725);
and U12013 (N_12013,N_1911,N_4042);
or U12014 (N_12014,N_2121,N_3904);
nand U12015 (N_12015,N_673,N_1233);
and U12016 (N_12016,N_1039,N_1659);
nand U12017 (N_12017,N_4832,N_4542);
or U12018 (N_12018,N_3589,N_2877);
xnor U12019 (N_12019,N_2195,N_5975);
and U12020 (N_12020,N_2140,N_603);
and U12021 (N_12021,N_961,N_2103);
or U12022 (N_12022,N_3743,N_5797);
or U12023 (N_12023,N_1228,N_5113);
and U12024 (N_12024,N_5379,N_2366);
and U12025 (N_12025,N_2118,N_4727);
nand U12026 (N_12026,N_4909,N_2352);
and U12027 (N_12027,N_5459,N_4253);
nand U12028 (N_12028,N_3867,N_5241);
or U12029 (N_12029,N_313,N_5713);
or U12030 (N_12030,N_3702,N_1364);
xor U12031 (N_12031,N_4988,N_1539);
or U12032 (N_12032,N_422,N_2670);
or U12033 (N_12033,N_2205,N_2660);
nor U12034 (N_12034,N_5724,N_2210);
xor U12035 (N_12035,N_5904,N_2183);
or U12036 (N_12036,N_2960,N_913);
or U12037 (N_12037,N_5736,N_2363);
or U12038 (N_12038,N_3168,N_4264);
or U12039 (N_12039,N_1287,N_4884);
or U12040 (N_12040,N_4971,N_5500);
or U12041 (N_12041,N_1067,N_1106);
and U12042 (N_12042,N_2493,N_5536);
or U12043 (N_12043,N_5606,N_2708);
or U12044 (N_12044,N_6167,N_4755);
and U12045 (N_12045,N_5796,N_701);
nand U12046 (N_12046,N_517,N_6180);
and U12047 (N_12047,N_1215,N_3419);
and U12048 (N_12048,N_3869,N_1541);
nand U12049 (N_12049,N_338,N_1931);
or U12050 (N_12050,N_675,N_2786);
and U12051 (N_12051,N_4550,N_1980);
nand U12052 (N_12052,N_1574,N_6022);
nand U12053 (N_12053,N_3992,N_5686);
xor U12054 (N_12054,N_1749,N_4517);
or U12055 (N_12055,N_5505,N_5538);
and U12056 (N_12056,N_1231,N_5400);
xor U12057 (N_12057,N_532,N_747);
xnor U12058 (N_12058,N_2911,N_6111);
nand U12059 (N_12059,N_3821,N_5334);
nor U12060 (N_12060,N_1361,N_1062);
nand U12061 (N_12061,N_2003,N_1685);
xor U12062 (N_12062,N_6193,N_5857);
and U12063 (N_12063,N_5663,N_2841);
nand U12064 (N_12064,N_4488,N_5971);
nor U12065 (N_12065,N_1506,N_2175);
nand U12066 (N_12066,N_5279,N_4044);
and U12067 (N_12067,N_839,N_1109);
or U12068 (N_12068,N_3433,N_6067);
xor U12069 (N_12069,N_2283,N_3205);
and U12070 (N_12070,N_3546,N_4645);
nor U12071 (N_12071,N_527,N_786);
or U12072 (N_12072,N_1489,N_3018);
xor U12073 (N_12073,N_1650,N_2968);
and U12074 (N_12074,N_2396,N_4865);
nand U12075 (N_12075,N_5047,N_3797);
or U12076 (N_12076,N_1078,N_2061);
or U12077 (N_12077,N_2153,N_5618);
nor U12078 (N_12078,N_4486,N_2096);
or U12079 (N_12079,N_664,N_4863);
or U12080 (N_12080,N_1421,N_1122);
or U12081 (N_12081,N_1376,N_2425);
nor U12082 (N_12082,N_5090,N_3038);
or U12083 (N_12083,N_4478,N_299);
xnor U12084 (N_12084,N_5275,N_4971);
nor U12085 (N_12085,N_4422,N_4707);
and U12086 (N_12086,N_2025,N_2787);
and U12087 (N_12087,N_459,N_5133);
and U12088 (N_12088,N_3969,N_2925);
or U12089 (N_12089,N_3412,N_3468);
or U12090 (N_12090,N_4616,N_4530);
nor U12091 (N_12091,N_4376,N_1786);
and U12092 (N_12092,N_3140,N_214);
nor U12093 (N_12093,N_5334,N_2566);
and U12094 (N_12094,N_2263,N_1895);
nor U12095 (N_12095,N_5485,N_73);
or U12096 (N_12096,N_2197,N_4421);
nand U12097 (N_12097,N_796,N_2918);
or U12098 (N_12098,N_575,N_1297);
or U12099 (N_12099,N_3851,N_879);
and U12100 (N_12100,N_1307,N_5464);
xnor U12101 (N_12101,N_5813,N_644);
or U12102 (N_12102,N_3902,N_5625);
nand U12103 (N_12103,N_2564,N_228);
or U12104 (N_12104,N_1622,N_1656);
and U12105 (N_12105,N_2428,N_2609);
and U12106 (N_12106,N_250,N_3703);
or U12107 (N_12107,N_4863,N_5386);
nand U12108 (N_12108,N_3266,N_2824);
nor U12109 (N_12109,N_5506,N_237);
or U12110 (N_12110,N_1857,N_5196);
nand U12111 (N_12111,N_922,N_5929);
xor U12112 (N_12112,N_5782,N_2616);
and U12113 (N_12113,N_2543,N_2272);
nand U12114 (N_12114,N_952,N_284);
nor U12115 (N_12115,N_2529,N_5530);
and U12116 (N_12116,N_4406,N_4009);
and U12117 (N_12117,N_5070,N_5993);
nand U12118 (N_12118,N_4572,N_5411);
or U12119 (N_12119,N_304,N_2343);
or U12120 (N_12120,N_2138,N_1330);
nor U12121 (N_12121,N_3541,N_896);
or U12122 (N_12122,N_770,N_5275);
and U12123 (N_12123,N_5761,N_532);
or U12124 (N_12124,N_6247,N_556);
or U12125 (N_12125,N_4343,N_2003);
and U12126 (N_12126,N_1698,N_4591);
or U12127 (N_12127,N_292,N_3531);
nor U12128 (N_12128,N_4316,N_3873);
or U12129 (N_12129,N_5130,N_5184);
or U12130 (N_12130,N_1382,N_1954);
nor U12131 (N_12131,N_2562,N_4926);
and U12132 (N_12132,N_5207,N_3976);
and U12133 (N_12133,N_3895,N_1784);
xnor U12134 (N_12134,N_5664,N_4279);
and U12135 (N_12135,N_5972,N_5449);
and U12136 (N_12136,N_4166,N_2800);
and U12137 (N_12137,N_3351,N_4953);
and U12138 (N_12138,N_4896,N_2981);
and U12139 (N_12139,N_32,N_3613);
nor U12140 (N_12140,N_885,N_2008);
nor U12141 (N_12141,N_5796,N_5022);
nand U12142 (N_12142,N_69,N_2417);
nor U12143 (N_12143,N_901,N_4233);
or U12144 (N_12144,N_4835,N_1345);
and U12145 (N_12145,N_3272,N_1249);
and U12146 (N_12146,N_3825,N_1465);
nor U12147 (N_12147,N_4362,N_2213);
or U12148 (N_12148,N_3605,N_4881);
and U12149 (N_12149,N_513,N_2812);
or U12150 (N_12150,N_5553,N_745);
or U12151 (N_12151,N_3863,N_2772);
nand U12152 (N_12152,N_5427,N_1970);
nor U12153 (N_12153,N_384,N_3775);
xnor U12154 (N_12154,N_3025,N_1456);
or U12155 (N_12155,N_1868,N_5742);
nor U12156 (N_12156,N_754,N_4226);
or U12157 (N_12157,N_2515,N_324);
nand U12158 (N_12158,N_3304,N_5972);
or U12159 (N_12159,N_2695,N_241);
nand U12160 (N_12160,N_2174,N_1231);
nand U12161 (N_12161,N_1157,N_5981);
and U12162 (N_12162,N_957,N_2262);
or U12163 (N_12163,N_1099,N_4937);
nor U12164 (N_12164,N_2868,N_4228);
or U12165 (N_12165,N_2609,N_170);
nand U12166 (N_12166,N_4308,N_6086);
xnor U12167 (N_12167,N_1768,N_6098);
and U12168 (N_12168,N_4287,N_2303);
and U12169 (N_12169,N_2590,N_1592);
or U12170 (N_12170,N_6041,N_3155);
and U12171 (N_12171,N_4269,N_1820);
xor U12172 (N_12172,N_1098,N_881);
xnor U12173 (N_12173,N_97,N_302);
or U12174 (N_12174,N_5510,N_4623);
and U12175 (N_12175,N_5100,N_460);
and U12176 (N_12176,N_3113,N_1320);
or U12177 (N_12177,N_2271,N_5246);
and U12178 (N_12178,N_260,N_2799);
and U12179 (N_12179,N_5659,N_2308);
nand U12180 (N_12180,N_3886,N_4068);
nand U12181 (N_12181,N_3706,N_1448);
or U12182 (N_12182,N_1637,N_2266);
or U12183 (N_12183,N_3463,N_1927);
nor U12184 (N_12184,N_2758,N_3036);
xor U12185 (N_12185,N_976,N_6163);
or U12186 (N_12186,N_2117,N_665);
and U12187 (N_12187,N_5273,N_2327);
nor U12188 (N_12188,N_4924,N_9);
or U12189 (N_12189,N_850,N_3614);
or U12190 (N_12190,N_5713,N_2407);
nor U12191 (N_12191,N_5711,N_5254);
nor U12192 (N_12192,N_1912,N_1543);
nand U12193 (N_12193,N_4272,N_4731);
and U12194 (N_12194,N_5745,N_2654);
nor U12195 (N_12195,N_4675,N_3522);
nand U12196 (N_12196,N_4489,N_1816);
nor U12197 (N_12197,N_5300,N_1445);
and U12198 (N_12198,N_5937,N_3016);
nand U12199 (N_12199,N_5111,N_2896);
and U12200 (N_12200,N_2261,N_2596);
and U12201 (N_12201,N_2897,N_2284);
nand U12202 (N_12202,N_4514,N_973);
nand U12203 (N_12203,N_5895,N_1927);
nand U12204 (N_12204,N_1996,N_3332);
nand U12205 (N_12205,N_3804,N_3322);
or U12206 (N_12206,N_397,N_865);
nand U12207 (N_12207,N_2610,N_5405);
and U12208 (N_12208,N_4799,N_1884);
nand U12209 (N_12209,N_2309,N_2105);
or U12210 (N_12210,N_1722,N_2030);
nor U12211 (N_12211,N_1891,N_2212);
nand U12212 (N_12212,N_5258,N_5037);
nor U12213 (N_12213,N_3480,N_1505);
nand U12214 (N_12214,N_1788,N_6093);
nand U12215 (N_12215,N_5667,N_2934);
nor U12216 (N_12216,N_2684,N_4801);
and U12217 (N_12217,N_6220,N_2047);
nand U12218 (N_12218,N_1548,N_4933);
xnor U12219 (N_12219,N_3941,N_5664);
xnor U12220 (N_12220,N_1848,N_49);
xor U12221 (N_12221,N_4891,N_5617);
nand U12222 (N_12222,N_1384,N_375);
nand U12223 (N_12223,N_759,N_2944);
nor U12224 (N_12224,N_6145,N_1667);
nor U12225 (N_12225,N_1949,N_3274);
nand U12226 (N_12226,N_6209,N_2646);
nor U12227 (N_12227,N_487,N_4339);
nor U12228 (N_12228,N_1354,N_5388);
and U12229 (N_12229,N_1159,N_1376);
and U12230 (N_12230,N_4492,N_4618);
and U12231 (N_12231,N_2573,N_6195);
nand U12232 (N_12232,N_3740,N_1341);
xor U12233 (N_12233,N_5247,N_3847);
xor U12234 (N_12234,N_3278,N_3765);
and U12235 (N_12235,N_5969,N_2280);
and U12236 (N_12236,N_1757,N_6009);
nor U12237 (N_12237,N_5350,N_4167);
and U12238 (N_12238,N_4761,N_281);
nand U12239 (N_12239,N_2503,N_1725);
or U12240 (N_12240,N_4505,N_308);
xor U12241 (N_12241,N_218,N_5756);
nand U12242 (N_12242,N_483,N_406);
nor U12243 (N_12243,N_75,N_5793);
nor U12244 (N_12244,N_2401,N_2106);
nor U12245 (N_12245,N_2700,N_4037);
nor U12246 (N_12246,N_622,N_3253);
nand U12247 (N_12247,N_5945,N_3276);
xnor U12248 (N_12248,N_2422,N_2206);
and U12249 (N_12249,N_737,N_5054);
and U12250 (N_12250,N_5382,N_3388);
nor U12251 (N_12251,N_2682,N_4175);
and U12252 (N_12252,N_5973,N_2102);
and U12253 (N_12253,N_2605,N_2653);
or U12254 (N_12254,N_3303,N_1965);
or U12255 (N_12255,N_2930,N_5287);
and U12256 (N_12256,N_5504,N_6151);
xnor U12257 (N_12257,N_5427,N_4487);
xor U12258 (N_12258,N_2558,N_4732);
or U12259 (N_12259,N_1474,N_3501);
and U12260 (N_12260,N_1724,N_2151);
and U12261 (N_12261,N_3409,N_3562);
and U12262 (N_12262,N_2708,N_1449);
or U12263 (N_12263,N_2779,N_4313);
and U12264 (N_12264,N_2489,N_2287);
or U12265 (N_12265,N_2441,N_2271);
xnor U12266 (N_12266,N_2651,N_137);
and U12267 (N_12267,N_156,N_3279);
nor U12268 (N_12268,N_4754,N_0);
and U12269 (N_12269,N_6172,N_4005);
and U12270 (N_12270,N_2423,N_4916);
or U12271 (N_12271,N_6018,N_3290);
and U12272 (N_12272,N_5647,N_5311);
nand U12273 (N_12273,N_3445,N_6053);
or U12274 (N_12274,N_3871,N_3253);
or U12275 (N_12275,N_876,N_3194);
or U12276 (N_12276,N_5786,N_5701);
and U12277 (N_12277,N_2421,N_4357);
and U12278 (N_12278,N_2220,N_3991);
nand U12279 (N_12279,N_2421,N_377);
nand U12280 (N_12280,N_5247,N_5978);
xor U12281 (N_12281,N_2985,N_1185);
and U12282 (N_12282,N_819,N_6175);
nor U12283 (N_12283,N_4757,N_4623);
nor U12284 (N_12284,N_5562,N_5895);
nor U12285 (N_12285,N_4016,N_3609);
xnor U12286 (N_12286,N_5713,N_2274);
or U12287 (N_12287,N_4846,N_3547);
or U12288 (N_12288,N_2000,N_1449);
and U12289 (N_12289,N_246,N_3466);
nand U12290 (N_12290,N_1599,N_3689);
nor U12291 (N_12291,N_1343,N_7);
nand U12292 (N_12292,N_4031,N_3633);
or U12293 (N_12293,N_4658,N_3081);
nor U12294 (N_12294,N_2422,N_3952);
nand U12295 (N_12295,N_1203,N_5616);
and U12296 (N_12296,N_1287,N_1444);
nor U12297 (N_12297,N_3161,N_5176);
or U12298 (N_12298,N_2236,N_2715);
xor U12299 (N_12299,N_183,N_873);
or U12300 (N_12300,N_2560,N_5854);
nand U12301 (N_12301,N_3342,N_1242);
and U12302 (N_12302,N_3873,N_558);
xor U12303 (N_12303,N_3069,N_4649);
nor U12304 (N_12304,N_1890,N_1704);
nand U12305 (N_12305,N_3849,N_1003);
nand U12306 (N_12306,N_1458,N_1300);
or U12307 (N_12307,N_5937,N_4821);
and U12308 (N_12308,N_948,N_1682);
and U12309 (N_12309,N_3335,N_2979);
xnor U12310 (N_12310,N_771,N_3053);
nand U12311 (N_12311,N_2276,N_5110);
nor U12312 (N_12312,N_3140,N_454);
and U12313 (N_12313,N_3637,N_6234);
nand U12314 (N_12314,N_4186,N_4121);
and U12315 (N_12315,N_2779,N_4868);
xnor U12316 (N_12316,N_2182,N_4747);
or U12317 (N_12317,N_4901,N_402);
nand U12318 (N_12318,N_5245,N_3790);
xnor U12319 (N_12319,N_6015,N_3724);
and U12320 (N_12320,N_5761,N_2418);
and U12321 (N_12321,N_4595,N_4494);
nor U12322 (N_12322,N_2569,N_5292);
or U12323 (N_12323,N_2802,N_4007);
nor U12324 (N_12324,N_3661,N_5203);
or U12325 (N_12325,N_5998,N_2945);
and U12326 (N_12326,N_77,N_6202);
and U12327 (N_12327,N_4588,N_2553);
nand U12328 (N_12328,N_1501,N_3990);
and U12329 (N_12329,N_5791,N_822);
xor U12330 (N_12330,N_3076,N_960);
or U12331 (N_12331,N_1535,N_660);
nand U12332 (N_12332,N_1796,N_540);
xor U12333 (N_12333,N_5916,N_2768);
nor U12334 (N_12334,N_5383,N_4283);
xnor U12335 (N_12335,N_4981,N_1648);
or U12336 (N_12336,N_469,N_4548);
nand U12337 (N_12337,N_2291,N_5509);
and U12338 (N_12338,N_5508,N_5603);
nand U12339 (N_12339,N_733,N_3586);
or U12340 (N_12340,N_911,N_1462);
nor U12341 (N_12341,N_5866,N_5734);
nor U12342 (N_12342,N_4646,N_4358);
and U12343 (N_12343,N_720,N_478);
and U12344 (N_12344,N_4974,N_4518);
nand U12345 (N_12345,N_1999,N_3476);
nor U12346 (N_12346,N_275,N_3594);
nand U12347 (N_12347,N_6006,N_1299);
nand U12348 (N_12348,N_244,N_4629);
and U12349 (N_12349,N_6093,N_5564);
and U12350 (N_12350,N_1742,N_3622);
and U12351 (N_12351,N_1853,N_3250);
or U12352 (N_12352,N_4963,N_957);
nand U12353 (N_12353,N_6095,N_528);
nor U12354 (N_12354,N_1736,N_1353);
nand U12355 (N_12355,N_2106,N_2780);
nor U12356 (N_12356,N_1227,N_749);
nor U12357 (N_12357,N_1889,N_4521);
nor U12358 (N_12358,N_4326,N_234);
nor U12359 (N_12359,N_5064,N_2115);
nor U12360 (N_12360,N_5339,N_3011);
nand U12361 (N_12361,N_4685,N_6050);
or U12362 (N_12362,N_4247,N_341);
nand U12363 (N_12363,N_66,N_464);
or U12364 (N_12364,N_5258,N_625);
nand U12365 (N_12365,N_3753,N_294);
nor U12366 (N_12366,N_2310,N_1637);
and U12367 (N_12367,N_5409,N_6245);
or U12368 (N_12368,N_4018,N_1268);
nor U12369 (N_12369,N_1030,N_294);
xor U12370 (N_12370,N_2649,N_4670);
nor U12371 (N_12371,N_2860,N_5381);
nor U12372 (N_12372,N_5258,N_2413);
nor U12373 (N_12373,N_6213,N_3127);
nand U12374 (N_12374,N_5814,N_108);
nor U12375 (N_12375,N_1072,N_3448);
nand U12376 (N_12376,N_3266,N_5894);
or U12377 (N_12377,N_1383,N_3836);
or U12378 (N_12378,N_3648,N_2319);
nor U12379 (N_12379,N_3447,N_1921);
xnor U12380 (N_12380,N_4601,N_147);
and U12381 (N_12381,N_3984,N_300);
or U12382 (N_12382,N_1989,N_4945);
nand U12383 (N_12383,N_1035,N_2829);
or U12384 (N_12384,N_3176,N_2669);
and U12385 (N_12385,N_3809,N_1957);
or U12386 (N_12386,N_533,N_1343);
nand U12387 (N_12387,N_665,N_1911);
nand U12388 (N_12388,N_5755,N_2457);
or U12389 (N_12389,N_4736,N_3178);
or U12390 (N_12390,N_2348,N_3836);
nand U12391 (N_12391,N_2770,N_5314);
xor U12392 (N_12392,N_2958,N_589);
nand U12393 (N_12393,N_293,N_1319);
nand U12394 (N_12394,N_4866,N_4435);
and U12395 (N_12395,N_959,N_936);
nor U12396 (N_12396,N_5479,N_4755);
nor U12397 (N_12397,N_380,N_4308);
or U12398 (N_12398,N_4733,N_4071);
and U12399 (N_12399,N_5451,N_5064);
nand U12400 (N_12400,N_5852,N_4401);
or U12401 (N_12401,N_4959,N_2548);
nor U12402 (N_12402,N_2102,N_6122);
and U12403 (N_12403,N_3567,N_740);
nor U12404 (N_12404,N_87,N_4496);
nand U12405 (N_12405,N_4079,N_2006);
or U12406 (N_12406,N_5825,N_2798);
and U12407 (N_12407,N_4080,N_557);
or U12408 (N_12408,N_2652,N_4347);
and U12409 (N_12409,N_293,N_4712);
nand U12410 (N_12410,N_4450,N_1213);
nor U12411 (N_12411,N_5701,N_2754);
or U12412 (N_12412,N_2998,N_5617);
xor U12413 (N_12413,N_1043,N_1410);
nor U12414 (N_12414,N_5133,N_1144);
and U12415 (N_12415,N_2359,N_3375);
and U12416 (N_12416,N_5603,N_1351);
or U12417 (N_12417,N_462,N_5486);
and U12418 (N_12418,N_233,N_4274);
nand U12419 (N_12419,N_76,N_3157);
nor U12420 (N_12420,N_3476,N_1742);
or U12421 (N_12421,N_1428,N_155);
nor U12422 (N_12422,N_3199,N_1589);
xnor U12423 (N_12423,N_643,N_1919);
nand U12424 (N_12424,N_2459,N_4796);
and U12425 (N_12425,N_5260,N_4236);
nor U12426 (N_12426,N_4142,N_1073);
and U12427 (N_12427,N_837,N_45);
xor U12428 (N_12428,N_1908,N_770);
nor U12429 (N_12429,N_2755,N_1254);
or U12430 (N_12430,N_1268,N_4203);
xnor U12431 (N_12431,N_5477,N_4492);
xor U12432 (N_12432,N_3822,N_3940);
nand U12433 (N_12433,N_1093,N_867);
or U12434 (N_12434,N_2,N_4089);
xor U12435 (N_12435,N_5354,N_5049);
nor U12436 (N_12436,N_3446,N_1195);
or U12437 (N_12437,N_56,N_484);
and U12438 (N_12438,N_4175,N_51);
nand U12439 (N_12439,N_3726,N_2197);
nor U12440 (N_12440,N_220,N_1749);
and U12441 (N_12441,N_3181,N_5039);
xor U12442 (N_12442,N_2034,N_932);
or U12443 (N_12443,N_2485,N_5907);
and U12444 (N_12444,N_3884,N_50);
or U12445 (N_12445,N_2959,N_250);
or U12446 (N_12446,N_4575,N_1787);
nor U12447 (N_12447,N_2738,N_2018);
and U12448 (N_12448,N_4637,N_416);
and U12449 (N_12449,N_4622,N_5775);
and U12450 (N_12450,N_1609,N_3592);
or U12451 (N_12451,N_2005,N_1351);
or U12452 (N_12452,N_3883,N_5376);
and U12453 (N_12453,N_1864,N_4667);
and U12454 (N_12454,N_5718,N_1631);
or U12455 (N_12455,N_2242,N_4006);
and U12456 (N_12456,N_1880,N_3242);
nor U12457 (N_12457,N_368,N_5540);
nand U12458 (N_12458,N_867,N_717);
nor U12459 (N_12459,N_6140,N_4890);
nor U12460 (N_12460,N_41,N_1931);
or U12461 (N_12461,N_375,N_3626);
nor U12462 (N_12462,N_1856,N_5529);
or U12463 (N_12463,N_1563,N_60);
xnor U12464 (N_12464,N_2169,N_2280);
and U12465 (N_12465,N_4662,N_5307);
nor U12466 (N_12466,N_1388,N_1214);
nor U12467 (N_12467,N_5919,N_600);
nand U12468 (N_12468,N_4353,N_414);
nand U12469 (N_12469,N_5670,N_5022);
nor U12470 (N_12470,N_429,N_2735);
nand U12471 (N_12471,N_1185,N_2067);
or U12472 (N_12472,N_699,N_1482);
nand U12473 (N_12473,N_6146,N_5805);
nand U12474 (N_12474,N_1513,N_3937);
and U12475 (N_12475,N_514,N_196);
nor U12476 (N_12476,N_1667,N_4283);
nor U12477 (N_12477,N_3441,N_3092);
and U12478 (N_12478,N_355,N_5566);
or U12479 (N_12479,N_1038,N_888);
and U12480 (N_12480,N_1240,N_3019);
nor U12481 (N_12481,N_4127,N_237);
nand U12482 (N_12482,N_5288,N_1299);
and U12483 (N_12483,N_6206,N_492);
or U12484 (N_12484,N_1655,N_44);
and U12485 (N_12485,N_1842,N_1437);
nand U12486 (N_12486,N_5212,N_3869);
nand U12487 (N_12487,N_5223,N_2165);
or U12488 (N_12488,N_376,N_1466);
or U12489 (N_12489,N_1714,N_4924);
xor U12490 (N_12490,N_4731,N_1446);
nand U12491 (N_12491,N_1459,N_2754);
nand U12492 (N_12492,N_280,N_731);
nor U12493 (N_12493,N_87,N_4564);
nor U12494 (N_12494,N_3187,N_5617);
or U12495 (N_12495,N_2522,N_5967);
and U12496 (N_12496,N_328,N_2541);
nor U12497 (N_12497,N_5162,N_135);
or U12498 (N_12498,N_4649,N_4461);
nor U12499 (N_12499,N_5315,N_914);
or U12500 (N_12500,N_9250,N_7785);
and U12501 (N_12501,N_7275,N_7445);
and U12502 (N_12502,N_11304,N_9429);
or U12503 (N_12503,N_6681,N_9593);
or U12504 (N_12504,N_8500,N_12091);
or U12505 (N_12505,N_8509,N_10682);
and U12506 (N_12506,N_8978,N_6773);
or U12507 (N_12507,N_12167,N_8737);
and U12508 (N_12508,N_9057,N_11889);
nor U12509 (N_12509,N_11034,N_6404);
nand U12510 (N_12510,N_10752,N_7892);
nor U12511 (N_12511,N_9446,N_7357);
nor U12512 (N_12512,N_8859,N_8204);
or U12513 (N_12513,N_8454,N_11052);
nor U12514 (N_12514,N_9142,N_11371);
nand U12515 (N_12515,N_8185,N_7551);
or U12516 (N_12516,N_6759,N_10240);
nor U12517 (N_12517,N_9392,N_10253);
xnor U12518 (N_12518,N_11769,N_8771);
or U12519 (N_12519,N_6441,N_8106);
or U12520 (N_12520,N_9670,N_8161);
nor U12521 (N_12521,N_8570,N_7817);
nand U12522 (N_12522,N_7321,N_6811);
xor U12523 (N_12523,N_7157,N_7594);
or U12524 (N_12524,N_10563,N_6419);
and U12525 (N_12525,N_8826,N_9104);
and U12526 (N_12526,N_7718,N_8680);
xnor U12527 (N_12527,N_6326,N_9710);
nor U12528 (N_12528,N_7988,N_8007);
nand U12529 (N_12529,N_11100,N_6855);
or U12530 (N_12530,N_10156,N_9943);
or U12531 (N_12531,N_8095,N_9186);
and U12532 (N_12532,N_9395,N_7710);
or U12533 (N_12533,N_10641,N_7158);
nand U12534 (N_12534,N_7093,N_7532);
nor U12535 (N_12535,N_7136,N_9424);
and U12536 (N_12536,N_7244,N_6955);
and U12537 (N_12537,N_8023,N_8723);
and U12538 (N_12538,N_9839,N_6286);
or U12539 (N_12539,N_7316,N_6804);
or U12540 (N_12540,N_10834,N_8100);
or U12541 (N_12541,N_8034,N_7847);
and U12542 (N_12542,N_10890,N_7754);
nand U12543 (N_12543,N_11541,N_10374);
nor U12544 (N_12544,N_10502,N_12027);
nor U12545 (N_12545,N_11649,N_12088);
nand U12546 (N_12546,N_10981,N_9569);
xnor U12547 (N_12547,N_11526,N_11033);
xnor U12548 (N_12548,N_9265,N_9366);
or U12549 (N_12549,N_10941,N_9354);
and U12550 (N_12550,N_12460,N_10866);
or U12551 (N_12551,N_10059,N_10996);
nand U12552 (N_12552,N_8693,N_10933);
nor U12553 (N_12553,N_8805,N_9739);
nor U12554 (N_12554,N_11922,N_11881);
xnor U12555 (N_12555,N_11528,N_7002);
and U12556 (N_12556,N_8507,N_12001);
or U12557 (N_12557,N_11116,N_11815);
or U12558 (N_12558,N_9609,N_11720);
nor U12559 (N_12559,N_9263,N_9717);
nor U12560 (N_12560,N_6726,N_10131);
or U12561 (N_12561,N_7620,N_10318);
or U12562 (N_12562,N_10212,N_7286);
nand U12563 (N_12563,N_7600,N_9008);
nand U12564 (N_12564,N_11647,N_10736);
nand U12565 (N_12565,N_11704,N_10602);
nand U12566 (N_12566,N_7082,N_10688);
nand U12567 (N_12567,N_8388,N_9464);
nand U12568 (N_12568,N_12262,N_9039);
or U12569 (N_12569,N_8225,N_9381);
nor U12570 (N_12570,N_11746,N_7723);
or U12571 (N_12571,N_10761,N_7593);
and U12572 (N_12572,N_10976,N_11002);
nor U12573 (N_12573,N_7577,N_11474);
and U12574 (N_12574,N_9854,N_11775);
and U12575 (N_12575,N_11384,N_8849);
nand U12576 (N_12576,N_9514,N_11787);
xnor U12577 (N_12577,N_7276,N_11478);
nor U12578 (N_12578,N_8439,N_11551);
nor U12579 (N_12579,N_8801,N_12463);
nand U12580 (N_12580,N_12319,N_7438);
or U12581 (N_12581,N_7787,N_11493);
and U12582 (N_12582,N_7161,N_12208);
nor U12583 (N_12583,N_12186,N_11359);
or U12584 (N_12584,N_6716,N_11098);
and U12585 (N_12585,N_11657,N_6546);
nor U12586 (N_12586,N_11328,N_8900);
nor U12587 (N_12587,N_11128,N_6826);
nor U12588 (N_12588,N_9603,N_6575);
and U12589 (N_12589,N_7356,N_10673);
nand U12590 (N_12590,N_10725,N_8206);
nor U12591 (N_12591,N_9965,N_10578);
nand U12592 (N_12592,N_7673,N_7665);
nor U12593 (N_12593,N_8514,N_9258);
and U12594 (N_12594,N_10064,N_9630);
and U12595 (N_12595,N_8700,N_9437);
or U12596 (N_12596,N_12295,N_11927);
xor U12597 (N_12597,N_11642,N_7826);
nor U12598 (N_12598,N_8262,N_9393);
and U12599 (N_12599,N_10877,N_7070);
nor U12600 (N_12600,N_6915,N_10629);
nand U12601 (N_12601,N_8729,N_6987);
nor U12602 (N_12602,N_7654,N_7343);
and U12603 (N_12603,N_10407,N_7549);
nor U12604 (N_12604,N_6983,N_6843);
or U12605 (N_12605,N_11874,N_11710);
and U12606 (N_12606,N_9802,N_7587);
and U12607 (N_12607,N_10119,N_12453);
nor U12608 (N_12608,N_9114,N_11693);
or U12609 (N_12609,N_10946,N_6485);
nor U12610 (N_12610,N_6999,N_9984);
and U12611 (N_12611,N_6814,N_9023);
xnor U12612 (N_12612,N_9279,N_7838);
nand U12613 (N_12613,N_11228,N_7698);
nand U12614 (N_12614,N_6293,N_11618);
or U12615 (N_12615,N_12024,N_12259);
nand U12616 (N_12616,N_9301,N_11736);
nand U12617 (N_12617,N_6686,N_12289);
nand U12618 (N_12618,N_6638,N_11149);
or U12619 (N_12619,N_7005,N_8854);
nand U12620 (N_12620,N_6619,N_7870);
xor U12621 (N_12621,N_6437,N_9151);
nand U12622 (N_12622,N_7498,N_10395);
xnor U12623 (N_12623,N_9410,N_10537);
nand U12624 (N_12624,N_8725,N_12403);
and U12625 (N_12625,N_9241,N_9225);
nand U12626 (N_12626,N_7573,N_7131);
nor U12627 (N_12627,N_9870,N_11409);
and U12628 (N_12628,N_9618,N_7644);
and U12629 (N_12629,N_11534,N_10277);
nand U12630 (N_12630,N_11561,N_7607);
nor U12631 (N_12631,N_8170,N_11792);
nor U12632 (N_12632,N_9064,N_8977);
nor U12633 (N_12633,N_11107,N_12444);
nor U12634 (N_12634,N_10010,N_12471);
or U12635 (N_12635,N_9999,N_9626);
xnor U12636 (N_12636,N_11588,N_11878);
nand U12637 (N_12637,N_11961,N_10450);
and U12638 (N_12638,N_10485,N_8236);
nor U12639 (N_12639,N_8132,N_11646);
or U12640 (N_12640,N_11663,N_10307);
and U12641 (N_12641,N_10842,N_7065);
nor U12642 (N_12642,N_10052,N_8409);
nand U12643 (N_12643,N_11249,N_11799);
nor U12644 (N_12644,N_10704,N_9841);
or U12645 (N_12645,N_10935,N_6787);
nor U12646 (N_12646,N_6539,N_9146);
and U12647 (N_12647,N_9314,N_9408);
and U12648 (N_12648,N_12323,N_6721);
or U12649 (N_12649,N_11739,N_11542);
or U12650 (N_12650,N_6518,N_6418);
nor U12651 (N_12651,N_10302,N_8656);
and U12652 (N_12652,N_10191,N_11932);
nor U12653 (N_12653,N_6699,N_6675);
or U12654 (N_12654,N_9772,N_10655);
nand U12655 (N_12655,N_6535,N_7642);
nand U12656 (N_12656,N_11712,N_11059);
and U12657 (N_12657,N_8630,N_7127);
nor U12658 (N_12658,N_10295,N_8765);
xnor U12659 (N_12659,N_9500,N_9116);
nor U12660 (N_12660,N_6550,N_9905);
or U12661 (N_12661,N_12160,N_8406);
nor U12662 (N_12662,N_8542,N_10367);
nand U12663 (N_12663,N_8646,N_12228);
nand U12664 (N_12664,N_7084,N_11141);
nor U12665 (N_12665,N_8193,N_8836);
nor U12666 (N_12666,N_8589,N_8713);
xor U12667 (N_12667,N_9445,N_6301);
nor U12668 (N_12668,N_8548,N_10837);
xnor U12669 (N_12669,N_10544,N_8954);
xnor U12670 (N_12670,N_11515,N_10244);
and U12671 (N_12671,N_9819,N_7201);
and U12672 (N_12672,N_6319,N_11833);
or U12673 (N_12673,N_10534,N_8026);
nand U12674 (N_12674,N_8947,N_7552);
xor U12675 (N_12675,N_7477,N_11826);
or U12676 (N_12676,N_9305,N_9480);
xnor U12677 (N_12677,N_9188,N_12122);
nor U12678 (N_12678,N_11948,N_10097);
and U12679 (N_12679,N_9721,N_9471);
nor U12680 (N_12680,N_6421,N_10880);
nor U12681 (N_12681,N_9953,N_11397);
nand U12682 (N_12682,N_9047,N_10232);
and U12683 (N_12683,N_9954,N_6931);
nand U12684 (N_12684,N_10488,N_11524);
nor U12685 (N_12685,N_6362,N_11613);
or U12686 (N_12686,N_8041,N_9482);
nor U12687 (N_12687,N_9028,N_6701);
nor U12688 (N_12688,N_11929,N_7079);
nand U12689 (N_12689,N_11206,N_7930);
nand U12690 (N_12690,N_6685,N_10854);
xor U12691 (N_12691,N_6742,N_11594);
and U12692 (N_12692,N_7020,N_10158);
and U12693 (N_12693,N_12318,N_7443);
xor U12694 (N_12694,N_12180,N_11740);
nor U12695 (N_12695,N_7175,N_8112);
nor U12696 (N_12696,N_12000,N_10762);
nor U12697 (N_12697,N_8345,N_11216);
or U12698 (N_12698,N_11157,N_10972);
or U12699 (N_12699,N_10749,N_9858);
or U12700 (N_12700,N_6310,N_11827);
and U12701 (N_12701,N_7729,N_8728);
or U12702 (N_12702,N_9950,N_7394);
and U12703 (N_12703,N_11911,N_12350);
nand U12704 (N_12704,N_6981,N_12406);
xnor U12705 (N_12705,N_8203,N_12164);
nor U12706 (N_12706,N_7756,N_10118);
and U12707 (N_12707,N_8412,N_6592);
or U12708 (N_12708,N_9293,N_7764);
xor U12709 (N_12709,N_11880,N_11131);
or U12710 (N_12710,N_6659,N_9848);
xnor U12711 (N_12711,N_7882,N_9503);
or U12712 (N_12712,N_11448,N_8941);
nor U12713 (N_12713,N_6979,N_10329);
xor U12714 (N_12714,N_10216,N_6464);
or U12715 (N_12715,N_11473,N_11234);
xor U12716 (N_12716,N_9896,N_8319);
and U12717 (N_12717,N_6745,N_9853);
or U12718 (N_12718,N_11010,N_10867);
nand U12719 (N_12719,N_10897,N_12333);
nand U12720 (N_12720,N_11521,N_11089);
nor U12721 (N_12721,N_12263,N_7991);
or U12722 (N_12722,N_12481,N_9576);
or U12723 (N_12723,N_6852,N_9352);
nor U12724 (N_12724,N_7719,N_10963);
nand U12725 (N_12725,N_10994,N_8361);
and U12726 (N_12726,N_7339,N_6824);
or U12727 (N_12727,N_7843,N_10843);
xnor U12728 (N_12728,N_9842,N_9031);
nor U12729 (N_12729,N_11194,N_11835);
xor U12730 (N_12730,N_9409,N_10123);
nand U12731 (N_12731,N_6698,N_9651);
nor U12732 (N_12732,N_7996,N_8435);
nand U12733 (N_12733,N_6356,N_8642);
xor U12734 (N_12734,N_10172,N_10681);
nor U12735 (N_12735,N_11491,N_8964);
xor U12736 (N_12736,N_12108,N_8087);
nand U12737 (N_12737,N_10914,N_9380);
and U12738 (N_12738,N_8149,N_11540);
and U12739 (N_12739,N_10968,N_10040);
or U12740 (N_12740,N_8598,N_8855);
nand U12741 (N_12741,N_7060,N_9535);
or U12742 (N_12742,N_11643,N_8910);
nand U12743 (N_12743,N_11173,N_7500);
or U12744 (N_12744,N_8753,N_11539);
xnor U12745 (N_12745,N_12364,N_7176);
nor U12746 (N_12746,N_8417,N_8788);
nor U12747 (N_12747,N_9234,N_11759);
and U12748 (N_12748,N_6848,N_8842);
and U12749 (N_12749,N_12429,N_8220);
xnor U12750 (N_12750,N_11415,N_6480);
or U12751 (N_12751,N_8721,N_8249);
or U12752 (N_12752,N_10106,N_11580);
or U12753 (N_12753,N_6451,N_8110);
nand U12754 (N_12754,N_6815,N_10584);
or U12755 (N_12755,N_8762,N_8137);
or U12756 (N_12756,N_9518,N_11807);
and U12757 (N_12757,N_7808,N_9013);
and U12758 (N_12758,N_11344,N_10051);
nand U12759 (N_12759,N_10417,N_9659);
nand U12760 (N_12760,N_9978,N_7298);
nor U12761 (N_12761,N_9126,N_9290);
or U12762 (N_12762,N_9784,N_9705);
nor U12763 (N_12763,N_9257,N_9966);
and U12764 (N_12764,N_7667,N_8892);
nand U12765 (N_12765,N_9932,N_12196);
or U12766 (N_12766,N_10004,N_7931);
and U12767 (N_12767,N_6283,N_6545);
nor U12768 (N_12768,N_8191,N_7041);
or U12769 (N_12769,N_12483,N_10891);
nor U12770 (N_12770,N_7491,N_10175);
nor U12771 (N_12771,N_8235,N_10046);
or U12772 (N_12772,N_8092,N_9442);
or U12773 (N_12773,N_8292,N_10943);
or U12774 (N_12774,N_10095,N_12231);
xor U12775 (N_12775,N_11144,N_7341);
nor U12776 (N_12776,N_8541,N_6876);
nand U12777 (N_12777,N_11620,N_7077);
and U12778 (N_12778,N_12170,N_8888);
nor U12779 (N_12779,N_10048,N_7852);
xnor U12780 (N_12780,N_7699,N_6400);
xor U12781 (N_12781,N_10017,N_8463);
xor U12782 (N_12782,N_12029,N_11604);
and U12783 (N_12783,N_9812,N_11706);
xnor U12784 (N_12784,N_6810,N_7350);
xor U12785 (N_12785,N_7714,N_12305);
and U12786 (N_12786,N_7758,N_11320);
nand U12787 (N_12787,N_11471,N_9814);
or U12788 (N_12788,N_7865,N_11220);
nand U12789 (N_12789,N_6869,N_7981);
and U12790 (N_12790,N_6253,N_9001);
xnor U12791 (N_12791,N_12156,N_11965);
or U12792 (N_12792,N_12356,N_12440);
and U12793 (N_12793,N_9731,N_7359);
or U12794 (N_12794,N_7524,N_8317);
or U12795 (N_12795,N_9387,N_11009);
or U12796 (N_12796,N_9649,N_7358);
nor U12797 (N_12797,N_8260,N_10267);
nor U12798 (N_12798,N_10722,N_10524);
nor U12799 (N_12799,N_9046,N_8334);
or U12800 (N_12800,N_6318,N_7210);
nand U12801 (N_12801,N_9245,N_9572);
or U12802 (N_12802,N_11047,N_7720);
and U12803 (N_12803,N_7674,N_10928);
xor U12804 (N_12804,N_9714,N_10683);
or U12805 (N_12805,N_6279,N_9214);
nor U12806 (N_12806,N_12378,N_7649);
nand U12807 (N_12807,N_7195,N_9036);
xnor U12808 (N_12808,N_11259,N_12270);
xor U12809 (N_12809,N_11903,N_12063);
nor U12810 (N_12810,N_8391,N_8821);
nand U12811 (N_12811,N_9097,N_8959);
nor U12812 (N_12812,N_11850,N_9824);
nor U12813 (N_12813,N_12321,N_7536);
nand U12814 (N_12814,N_12168,N_12197);
and U12815 (N_12815,N_9745,N_10706);
or U12816 (N_12816,N_10361,N_10068);
nor U12817 (N_12817,N_10830,N_7514);
and U12818 (N_12818,N_8610,N_9573);
nor U12819 (N_12819,N_8974,N_11057);
and U12820 (N_12820,N_9532,N_11812);
nand U12821 (N_12821,N_8754,N_10530);
and U12822 (N_12822,N_11076,N_7633);
nand U12823 (N_12823,N_10930,N_10822);
nor U12824 (N_12824,N_9306,N_8405);
nand U12825 (N_12825,N_8030,N_11062);
or U12826 (N_12826,N_12239,N_8212);
and U12827 (N_12827,N_10319,N_9270);
nand U12828 (N_12828,N_10679,N_8118);
nand U12829 (N_12829,N_8365,N_6957);
xnor U12830 (N_12830,N_11680,N_9895);
xor U12831 (N_12831,N_12358,N_9223);
nor U12832 (N_12832,N_9902,N_8985);
and U12833 (N_12833,N_10551,N_12003);
and U12834 (N_12834,N_7203,N_8759);
nor U12835 (N_12835,N_8672,N_7533);
or U12836 (N_12836,N_9019,N_12447);
nand U12837 (N_12837,N_7345,N_11197);
and U12838 (N_12838,N_12194,N_12274);
nand U12839 (N_12839,N_6271,N_7483);
or U12840 (N_12840,N_8618,N_10391);
nor U12841 (N_12841,N_6417,N_11803);
xor U12842 (N_12842,N_7288,N_6532);
nand U12843 (N_12843,N_11142,N_8601);
nand U12844 (N_12844,N_7253,N_11527);
and U12845 (N_12845,N_7799,N_8755);
nand U12846 (N_12846,N_11975,N_7389);
xnor U12847 (N_12847,N_8505,N_9222);
xor U12848 (N_12848,N_9699,N_6488);
or U12849 (N_12849,N_6692,N_7290);
or U12850 (N_12850,N_11426,N_7061);
nor U12851 (N_12851,N_7715,N_10304);
nor U12852 (N_12852,N_11702,N_7984);
and U12853 (N_12853,N_7267,N_6368);
or U12854 (N_12854,N_8965,N_8577);
nand U12855 (N_12855,N_8897,N_10627);
nor U12856 (N_12856,N_12470,N_11797);
and U12857 (N_12857,N_8215,N_6474);
nor U12858 (N_12858,N_11614,N_7328);
xor U12859 (N_12859,N_10020,N_9737);
and U12860 (N_12860,N_6431,N_12268);
and U12861 (N_12861,N_10215,N_10847);
and U12862 (N_12862,N_10870,N_7429);
nand U12863 (N_12863,N_11592,N_6743);
or U12864 (N_12864,N_8904,N_10667);
and U12865 (N_12865,N_9233,N_8329);
nand U12866 (N_12866,N_11182,N_12493);
and U12867 (N_12867,N_12140,N_6537);
and U12868 (N_12868,N_8530,N_6323);
nor U12869 (N_12869,N_11346,N_8939);
nor U12870 (N_12870,N_10327,N_7259);
and U12871 (N_12871,N_11793,N_8285);
or U12872 (N_12872,N_12314,N_8767);
nor U12873 (N_12873,N_11627,N_7803);
nand U12874 (N_12874,N_11487,N_7324);
nor U12875 (N_12875,N_10542,N_7293);
and U12876 (N_12876,N_10889,N_9549);
or U12877 (N_12877,N_9928,N_6921);
nand U12878 (N_12878,N_11801,N_11199);
and U12879 (N_12879,N_8572,N_12322);
xnor U12880 (N_12880,N_12080,N_10632);
nand U12881 (N_12881,N_8057,N_11246);
or U12882 (N_12882,N_9583,N_11584);
and U12883 (N_12883,N_8163,N_6627);
nor U12884 (N_12884,N_11694,N_7562);
and U12885 (N_12885,N_8146,N_8366);
nand U12886 (N_12886,N_10671,N_6678);
nor U12887 (N_12887,N_8838,N_10316);
or U12888 (N_12888,N_7215,N_7995);
xor U12889 (N_12889,N_12419,N_6765);
nor U12890 (N_12890,N_6553,N_11930);
and U12891 (N_12891,N_12066,N_11837);
nor U12892 (N_12892,N_11495,N_7905);
or U12893 (N_12893,N_6785,N_8493);
or U12894 (N_12894,N_12416,N_10903);
xor U12895 (N_12895,N_10390,N_6322);
or U12896 (N_12896,N_11678,N_8865);
or U12897 (N_12897,N_11247,N_6806);
and U12898 (N_12898,N_7936,N_10644);
and U12899 (N_12899,N_6605,N_7575);
nor U12900 (N_12900,N_7406,N_11215);
and U12901 (N_12901,N_7953,N_11684);
or U12902 (N_12902,N_9751,N_9575);
nor U12903 (N_12903,N_9135,N_11104);
and U12904 (N_12904,N_8177,N_10593);
nor U12905 (N_12905,N_10099,N_10429);
or U12906 (N_12906,N_9718,N_11139);
nand U12907 (N_12907,N_6623,N_9120);
nor U12908 (N_12908,N_11440,N_11847);
or U12909 (N_12909,N_7545,N_9274);
xnor U12910 (N_12910,N_8072,N_9458);
nand U12911 (N_12911,N_6290,N_7148);
xor U12912 (N_12912,N_9663,N_7006);
and U12913 (N_12913,N_9426,N_12382);
nand U12914 (N_12914,N_12249,N_9300);
xnor U12915 (N_12915,N_10455,N_8823);
xor U12916 (N_12916,N_10043,N_7608);
nor U12917 (N_12917,N_6709,N_7924);
nor U12918 (N_12918,N_10800,N_9697);
and U12919 (N_12919,N_10210,N_8582);
nand U12920 (N_12920,N_9256,N_6969);
and U12921 (N_12921,N_6430,N_11662);
xor U12922 (N_12922,N_11337,N_7822);
or U12923 (N_12923,N_7749,N_12181);
or U12924 (N_12924,N_11412,N_6251);
nor U12925 (N_12925,N_9351,N_7089);
and U12926 (N_12926,N_6782,N_10481);
nor U12927 (N_12927,N_7179,N_8781);
or U12928 (N_12928,N_10734,N_10451);
nor U12929 (N_12929,N_6949,N_7963);
and U12930 (N_12930,N_8004,N_9136);
or U12931 (N_12931,N_7507,N_12462);
and U12932 (N_12932,N_11027,N_7236);
nand U12933 (N_12933,N_12432,N_9684);
xnor U12934 (N_12934,N_9208,N_9373);
and U12935 (N_12935,N_11334,N_12171);
nor U12936 (N_12936,N_10492,N_7909);
and U12937 (N_12937,N_11782,N_8165);
nor U12938 (N_12938,N_8117,N_9648);
nand U12939 (N_12939,N_9880,N_7519);
nand U12940 (N_12940,N_8085,N_10311);
or U12941 (N_12941,N_9828,N_7027);
xnor U12942 (N_12942,N_7771,N_7205);
and U12943 (N_12943,N_8683,N_10886);
nor U12944 (N_12944,N_7589,N_12205);
nor U12945 (N_12945,N_9212,N_10606);
nand U12946 (N_12946,N_6714,N_11365);
or U12947 (N_12947,N_11749,N_7653);
xnor U12948 (N_12948,N_11648,N_9890);
nor U12949 (N_12949,N_11665,N_8848);
or U12950 (N_12950,N_8824,N_11176);
or U12951 (N_12951,N_8616,N_11405);
nand U12952 (N_12952,N_8423,N_8928);
and U12953 (N_12953,N_8238,N_7439);
nor U12954 (N_12954,N_11174,N_6670);
or U12955 (N_12955,N_8169,N_12187);
or U12956 (N_12956,N_9740,N_9620);
and U12957 (N_12957,N_11517,N_9147);
nand U12958 (N_12958,N_12390,N_10234);
and U12959 (N_12959,N_8661,N_8649);
nor U12960 (N_12960,N_7265,N_8956);
or U12961 (N_12961,N_7380,N_10344);
nor U12962 (N_12962,N_11818,N_10613);
or U12963 (N_12963,N_7327,N_12461);
nand U12964 (N_12964,N_12216,N_11755);
and U12965 (N_12965,N_9899,N_11898);
xnor U12966 (N_12966,N_12198,N_10619);
nand U12967 (N_12967,N_9448,N_10998);
and U12968 (N_12968,N_8456,N_7025);
or U12969 (N_12969,N_8099,N_8019);
nor U12970 (N_12970,N_10532,N_12455);
nand U12971 (N_12971,N_6472,N_8520);
nand U12972 (N_12972,N_10419,N_11834);
or U12973 (N_12973,N_8352,N_10075);
and U12974 (N_12974,N_7442,N_10786);
and U12975 (N_12975,N_8551,N_6702);
and U12976 (N_12976,N_9782,N_7782);
xnor U12977 (N_12977,N_7485,N_6505);
nor U12978 (N_12978,N_7130,N_11041);
nor U12979 (N_12979,N_10514,N_6340);
nand U12980 (N_12980,N_6524,N_11306);
xnor U12981 (N_12981,N_7187,N_10339);
nor U12982 (N_12982,N_10711,N_6762);
nor U12983 (N_12983,N_8891,N_11240);
and U12984 (N_12984,N_7509,N_8399);
nor U12985 (N_12985,N_6391,N_7263);
or U12986 (N_12986,N_9391,N_8907);
or U12987 (N_12987,N_9598,N_12281);
nand U12988 (N_12988,N_8351,N_9406);
and U12989 (N_12989,N_9347,N_8491);
xor U12990 (N_12990,N_10709,N_6395);
xor U12991 (N_12991,N_6831,N_12166);
nor U12992 (N_12992,N_11123,N_10664);
nor U12993 (N_12993,N_6603,N_9892);
nand U12994 (N_12994,N_7416,N_11751);
nand U12995 (N_12995,N_6479,N_8279);
or U12996 (N_12996,N_8088,N_12165);
and U12997 (N_12997,N_8931,N_11695);
nor U12998 (N_12998,N_8575,N_7582);
or U12999 (N_12999,N_8267,N_10349);
nand U13000 (N_13000,N_6860,N_12119);
nand U13001 (N_13001,N_6940,N_10337);
and U13002 (N_13002,N_10479,N_12214);
nor U13003 (N_13003,N_9282,N_6384);
nand U13004 (N_13004,N_11288,N_10865);
and U13005 (N_13005,N_8538,N_9809);
and U13006 (N_13006,N_6456,N_6261);
nand U13007 (N_13007,N_9613,N_8643);
and U13008 (N_13008,N_9163,N_11053);
nor U13009 (N_13009,N_7855,N_11981);
or U13010 (N_13010,N_6277,N_10500);
xnor U13011 (N_13011,N_9770,N_6475);
and U13012 (N_13012,N_6708,N_8518);
nand U13013 (N_13013,N_11723,N_9181);
or U13014 (N_13014,N_9465,N_7306);
or U13015 (N_13015,N_10045,N_11439);
and U13016 (N_13016,N_7537,N_11105);
nor U13017 (N_13017,N_11629,N_9995);
xor U13018 (N_13018,N_11086,N_10801);
or U13019 (N_13019,N_11050,N_9836);
nand U13020 (N_13020,N_11951,N_7938);
nor U13021 (N_13021,N_11659,N_8994);
and U13022 (N_13022,N_11441,N_8535);
and U13023 (N_13023,N_7090,N_8293);
nand U13024 (N_13024,N_8814,N_10496);
nor U13025 (N_13025,N_9182,N_9026);
nor U13026 (N_13026,N_7779,N_12337);
or U13027 (N_13027,N_9192,N_7851);
or U13028 (N_13028,N_10796,N_11420);
nor U13029 (N_13029,N_8387,N_9103);
nand U13030 (N_13030,N_8671,N_11970);
and U13031 (N_13031,N_12404,N_11705);
or U13032 (N_13032,N_7024,N_10650);
nor U13033 (N_13033,N_7736,N_9364);
nor U13034 (N_13034,N_12121,N_8628);
or U13035 (N_13035,N_9012,N_10427);
nor U13036 (N_13036,N_6359,N_8414);
and U13037 (N_13037,N_6289,N_11986);
and U13038 (N_13038,N_6793,N_7910);
and U13039 (N_13039,N_9886,N_11783);
and U13040 (N_13040,N_11806,N_10757);
and U13041 (N_13041,N_10723,N_8103);
nor U13042 (N_13042,N_9128,N_6578);
nand U13043 (N_13043,N_9275,N_7780);
and U13044 (N_13044,N_9750,N_8340);
xnor U13045 (N_13045,N_9695,N_12031);
nor U13046 (N_13046,N_11263,N_12245);
xnor U13047 (N_13047,N_10204,N_10397);
and U13048 (N_13048,N_12273,N_7252);
or U13049 (N_13049,N_9523,N_9799);
nand U13050 (N_13050,N_8229,N_8660);
nor U13051 (N_13051,N_10333,N_6382);
and U13052 (N_13052,N_8666,N_7918);
or U13053 (N_13053,N_11163,N_12175);
and U13054 (N_13054,N_6416,N_9320);
nand U13055 (N_13055,N_10330,N_10173);
nand U13056 (N_13056,N_6410,N_12292);
nand U13057 (N_13057,N_9597,N_10183);
xor U13058 (N_13058,N_12225,N_12120);
and U13059 (N_13059,N_12400,N_12478);
nand U13060 (N_13060,N_9205,N_7794);
nand U13061 (N_13061,N_8125,N_8039);
or U13062 (N_13062,N_11475,N_10114);
nor U13063 (N_13063,N_10272,N_11393);
nor U13064 (N_13064,N_6351,N_11950);
xor U13065 (N_13065,N_11083,N_7372);
or U13066 (N_13066,N_6903,N_7903);
or U13067 (N_13067,N_8674,N_6588);
nor U13068 (N_13068,N_8063,N_9400);
nand U13069 (N_13069,N_10936,N_7224);
nand U13070 (N_13070,N_11688,N_8336);
nand U13071 (N_13071,N_6493,N_10190);
nand U13072 (N_13072,N_7518,N_8779);
and U13073 (N_13073,N_9066,N_8893);
nor U13074 (N_13074,N_6967,N_7475);
or U13075 (N_13075,N_9846,N_7617);
nand U13076 (N_13076,N_8176,N_10343);
xnor U13077 (N_13077,N_9359,N_12328);
or U13078 (N_13078,N_10876,N_9834);
nor U13079 (N_13079,N_10025,N_6491);
or U13080 (N_13080,N_9478,N_11358);
and U13081 (N_13081,N_10207,N_11260);
nor U13082 (N_13082,N_9586,N_6856);
nor U13083 (N_13083,N_9668,N_11275);
or U13084 (N_13084,N_6476,N_11867);
or U13085 (N_13085,N_8837,N_12282);
or U13086 (N_13086,N_8578,N_8813);
and U13087 (N_13087,N_9599,N_6613);
nand U13088 (N_13088,N_8316,N_10789);
nand U13089 (N_13089,N_6663,N_10198);
or U13090 (N_13090,N_8341,N_6316);
or U13091 (N_13091,N_8806,N_9253);
and U13092 (N_13092,N_10448,N_10956);
nor U13093 (N_13093,N_11872,N_9388);
xor U13094 (N_13094,N_10355,N_10769);
nor U13095 (N_13095,N_12296,N_9302);
nor U13096 (N_13096,N_10484,N_9869);
xor U13097 (N_13097,N_7313,N_8993);
and U13098 (N_13098,N_9589,N_11938);
nand U13099 (N_13099,N_10315,N_8820);
and U13100 (N_13100,N_10562,N_10162);
xnor U13101 (N_13101,N_10495,N_12430);
nor U13102 (N_13102,N_10651,N_9730);
nand U13103 (N_13103,N_7778,N_7659);
or U13104 (N_13104,N_9052,N_7950);
xor U13105 (N_13105,N_8403,N_11979);
and U13106 (N_13106,N_6295,N_11844);
nand U13107 (N_13107,N_10299,N_10817);
and U13108 (N_13108,N_11976,N_8344);
and U13109 (N_13109,N_9796,N_9153);
and U13110 (N_13110,N_11155,N_6794);
nand U13111 (N_13111,N_7019,N_7663);
or U13112 (N_13112,N_10378,N_8462);
nand U13113 (N_13113,N_8226,N_10308);
nor U13114 (N_13114,N_6703,N_10577);
xor U13115 (N_13115,N_6982,N_12101);
or U13116 (N_13116,N_10387,N_10491);
nand U13117 (N_13117,N_7450,N_11229);
nor U13118 (N_13118,N_7044,N_9759);
and U13119 (N_13119,N_7192,N_7486);
nand U13120 (N_13120,N_7700,N_11094);
and U13121 (N_13121,N_10195,N_9108);
nand U13122 (N_13122,N_11532,N_12386);
nor U13123 (N_13123,N_8283,N_9927);
xnor U13124 (N_13124,N_11191,N_7048);
and U13125 (N_13125,N_11125,N_8306);
and U13126 (N_13126,N_6837,N_6552);
nand U13127 (N_13127,N_7684,N_12310);
nand U13128 (N_13128,N_8211,N_10366);
nand U13129 (N_13129,N_8015,N_7883);
and U13130 (N_13130,N_8209,N_9025);
nand U13131 (N_13131,N_11639,N_12078);
nor U13132 (N_13132,N_8420,N_8946);
or U13133 (N_13133,N_8547,N_11323);
xnor U13134 (N_13134,N_9792,N_11421);
nand U13135 (N_13135,N_6363,N_11460);
and U13136 (N_13136,N_10120,N_9255);
nand U13137 (N_13137,N_10896,N_9991);
nor U13138 (N_13138,N_9526,N_11192);
and U13139 (N_13139,N_11701,N_10044);
nand U13140 (N_13140,N_8915,N_11676);
xnor U13141 (N_13141,N_7482,N_12022);
or U13142 (N_13142,N_9606,N_8374);
or U13143 (N_13143,N_7859,N_8699);
or U13144 (N_13144,N_11280,N_7388);
and U13145 (N_13145,N_6531,N_12087);
or U13146 (N_13146,N_9521,N_11770);
nor U13147 (N_13147,N_9700,N_9085);
nand U13148 (N_13148,N_9081,N_8079);
nand U13149 (N_13149,N_7580,N_7945);
nor U13150 (N_13150,N_7257,N_7925);
nor U13151 (N_13151,N_8914,N_11634);
nor U13152 (N_13152,N_10259,N_8684);
xor U13153 (N_13153,N_6357,N_7655);
nand U13154 (N_13154,N_9553,N_7231);
and U13155 (N_13155,N_9958,N_8216);
and U13156 (N_13156,N_11778,N_10270);
or U13157 (N_13157,N_7053,N_9438);
or U13158 (N_13158,N_6763,N_7128);
nor U13159 (N_13159,N_11983,N_9662);
nor U13160 (N_13160,N_8717,N_8935);
nor U13161 (N_13161,N_9433,N_12174);
nand U13162 (N_13162,N_11355,N_6873);
nand U13163 (N_13163,N_9977,N_9632);
and U13164 (N_13164,N_7269,N_9129);
or U13165 (N_13165,N_8825,N_11013);
nor U13166 (N_13166,N_8780,N_6533);
nor U13167 (N_13167,N_7846,N_10081);
and U13168 (N_13168,N_12412,N_9358);
nand U13169 (N_13169,N_10146,N_9539);
nor U13170 (N_13170,N_10379,N_10797);
or U13171 (N_13171,N_10373,N_11503);
and U13172 (N_13172,N_7092,N_11418);
and U13173 (N_13173,N_9332,N_8544);
nand U13174 (N_13174,N_10691,N_7046);
xnor U13175 (N_13175,N_6314,N_9881);
nand U13176 (N_13176,N_9860,N_9507);
nand U13177 (N_13177,N_6941,N_8870);
xor U13178 (N_13178,N_11284,N_7638);
nand U13179 (N_13179,N_8701,N_8354);
nor U13180 (N_13180,N_10680,N_8309);
nand U13181 (N_13181,N_9893,N_9112);
xnor U13182 (N_13182,N_10236,N_7959);
or U13183 (N_13183,N_6308,N_7247);
nand U13184 (N_13184,N_10838,N_8981);
nor U13185 (N_13185,N_6851,N_6563);
nor U13186 (N_13186,N_7781,N_9217);
nor U13187 (N_13187,N_9083,N_11092);
nor U13188 (N_13188,N_7541,N_10165);
or U13189 (N_13189,N_9474,N_8058);
or U13190 (N_13190,N_7137,N_7382);
and U13191 (N_13191,N_9754,N_8665);
or U13192 (N_13192,N_12076,N_11573);
and U13193 (N_13193,N_12496,N_9470);
and U13194 (N_13194,N_10170,N_6640);
xnor U13195 (N_13195,N_10430,N_8339);
and U13196 (N_13196,N_9107,N_6263);
or U13197 (N_13197,N_9774,N_10285);
or U13198 (N_13198,N_11635,N_8400);
or U13199 (N_13199,N_10919,N_6355);
or U13200 (N_13200,N_8619,N_11341);
and U13201 (N_13201,N_8822,N_6753);
or U13202 (N_13202,N_12402,N_7888);
and U13203 (N_13203,N_9189,N_6554);
nand U13204 (N_13204,N_10564,N_6386);
nand U13205 (N_13205,N_7504,N_10345);
and U13206 (N_13206,N_7166,N_11548);
nand U13207 (N_13207,N_6278,N_9962);
nor U13208 (N_13208,N_9501,N_12242);
or U13209 (N_13209,N_8797,N_11070);
nor U13210 (N_13210,N_9567,N_10790);
and U13211 (N_13211,N_7297,N_9335);
nand U13212 (N_13212,N_10753,N_7102);
or U13213 (N_13213,N_11110,N_6812);
nor U13214 (N_13214,N_6706,N_6549);
and U13215 (N_13215,N_7944,N_10713);
xnor U13216 (N_13216,N_8984,N_7493);
and U13217 (N_13217,N_10083,N_7383);
and U13218 (N_13218,N_6343,N_9228);
or U13219 (N_13219,N_10022,N_9431);
nor U13220 (N_13220,N_10692,N_7103);
nand U13221 (N_13221,N_6281,N_12209);
nor U13222 (N_13222,N_10437,N_9733);
and U13223 (N_13223,N_7941,N_7110);
and U13224 (N_13224,N_7322,N_12450);
xnor U13225 (N_13225,N_10546,N_6626);
and U13226 (N_13226,N_10325,N_6459);
or U13227 (N_13227,N_9677,N_9725);
xnor U13228 (N_13228,N_9919,N_10107);
and U13229 (N_13229,N_6997,N_6526);
and U13230 (N_13230,N_8152,N_11232);
and U13231 (N_13231,N_10642,N_6573);
and U13232 (N_13232,N_7804,N_11957);
or U13233 (N_13233,N_11721,N_7329);
nand U13234 (N_13234,N_8834,N_9313);
or U13235 (N_13235,N_11511,N_8310);
nor U13236 (N_13236,N_8596,N_10294);
nand U13237 (N_13237,N_9040,N_12464);
and U13238 (N_13238,N_7237,N_7923);
nand U13239 (N_13239,N_8817,N_6473);
xor U13240 (N_13240,N_8436,N_11928);
or U13241 (N_13241,N_6565,N_9642);
or U13242 (N_13242,N_10412,N_7034);
or U13243 (N_13243,N_12092,N_12113);
nand U13244 (N_13244,N_9086,N_7226);
or U13245 (N_13245,N_9000,N_7399);
nand U13246 (N_13246,N_8151,N_8051);
nor U13247 (N_13247,N_11403,N_9581);
nand U13248 (N_13248,N_8816,N_8075);
or U13249 (N_13249,N_11578,N_7409);
nand U13250 (N_13250,N_7970,N_6947);
or U13251 (N_13251,N_8592,N_12327);
and U13252 (N_13252,N_11982,N_9154);
xnor U13253 (N_13253,N_6555,N_7078);
nor U13254 (N_13254,N_6650,N_11278);
nand U13255 (N_13255,N_12248,N_7457);
or U13256 (N_13256,N_9811,N_7590);
and U13257 (N_13257,N_11379,N_6622);
or U13258 (N_13258,N_10939,N_6341);
and U13259 (N_13259,N_8561,N_7755);
or U13260 (N_13260,N_12118,N_9897);
and U13261 (N_13261,N_10794,N_9826);
nand U13262 (N_13262,N_6906,N_10755);
or U13263 (N_13263,N_9692,N_11018);
and U13264 (N_13264,N_8253,N_9596);
nand U13265 (N_13265,N_9422,N_8943);
nand U13266 (N_13266,N_7704,N_11761);
and U13267 (N_13267,N_10023,N_10129);
nand U13268 (N_13268,N_12050,N_11544);
nand U13269 (N_13269,N_8123,N_12494);
nand U13270 (N_13270,N_7513,N_9278);
and U13271 (N_13271,N_7777,N_8731);
xnor U13272 (N_13272,N_10122,N_7141);
nand U13273 (N_13273,N_7512,N_10237);
nor U13274 (N_13274,N_12428,N_6482);
or U13275 (N_13275,N_12443,N_11077);
xor U13276 (N_13276,N_12366,N_8905);
xor U13277 (N_13277,N_8473,N_9453);
nor U13278 (N_13278,N_12103,N_8346);
and U13279 (N_13279,N_7885,N_8609);
or U13280 (N_13280,N_6683,N_6574);
and U13281 (N_13281,N_9762,N_8282);
nand U13282 (N_13282,N_12045,N_12437);
nor U13283 (N_13283,N_8494,N_11802);
and U13284 (N_13284,N_11810,N_6352);
nor U13285 (N_13285,N_8757,N_6777);
nand U13286 (N_13286,N_6349,N_11272);
nand U13287 (N_13287,N_7411,N_8028);
nor U13288 (N_13288,N_8466,N_6733);
and U13289 (N_13289,N_11279,N_8690);
and U13290 (N_13290,N_9432,N_9619);
xor U13291 (N_13291,N_9830,N_11170);
xor U13292 (N_13292,N_12012,N_8086);
and U13293 (N_13293,N_6465,N_6428);
xor U13294 (N_13294,N_6965,N_6443);
nor U13295 (N_13295,N_9042,N_8416);
or U13296 (N_13296,N_8523,N_7289);
or U13297 (N_13297,N_11464,N_10987);
xor U13298 (N_13298,N_8231,N_7326);
nand U13299 (N_13299,N_7160,N_8957);
nor U13300 (N_13300,N_8430,N_10788);
and U13301 (N_13301,N_7164,N_7299);
nand U13302 (N_13302,N_9690,N_7948);
nand U13303 (N_13303,N_10151,N_10643);
and U13304 (N_13304,N_12375,N_10388);
or U13305 (N_13305,N_7597,N_10535);
xnor U13306 (N_13306,N_7877,N_9484);
nand U13307 (N_13307,N_10661,N_6477);
and U13308 (N_13308,N_9653,N_7732);
or U13309 (N_13309,N_11560,N_7717);
nand U13310 (N_13310,N_11599,N_6490);
nor U13311 (N_13311,N_12227,N_11717);
or U13312 (N_13312,N_11213,N_11363);
nand U13313 (N_13313,N_7499,N_10006);
xnor U13314 (N_13314,N_11254,N_11840);
xor U13315 (N_13315,N_10531,N_7933);
nand U13316 (N_13316,N_8013,N_10592);
nor U13317 (N_13317,N_10701,N_11088);
or U13318 (N_13318,N_8172,N_6617);
nor U13319 (N_13319,N_6586,N_8901);
nor U13320 (N_13320,N_9346,N_7898);
and U13321 (N_13321,N_12010,N_9350);
and U13322 (N_13322,N_10738,N_9942);
nor U13323 (N_13323,N_11114,N_7949);
or U13324 (N_13324,N_7869,N_7557);
and U13325 (N_13325,N_11082,N_11293);
nor U13326 (N_13326,N_11301,N_12312);
and U13327 (N_13327,N_8421,N_7330);
and U13328 (N_13328,N_10983,N_7618);
nand U13329 (N_13329,N_9156,N_7369);
nor U13330 (N_13330,N_8070,N_11283);
nand U13331 (N_13331,N_7459,N_12250);
and U13332 (N_13332,N_7366,N_11164);
nor U13333 (N_13333,N_11202,N_11851);
nor U13334 (N_13334,N_6754,N_8464);
or U13335 (N_13335,N_10763,N_9468);
or U13336 (N_13336,N_11177,N_11376);
and U13337 (N_13337,N_6881,N_11188);
or U13338 (N_13338,N_12372,N_11877);
nor U13339 (N_13339,N_10221,N_10341);
or U13340 (N_13340,N_9403,N_9864);
nor U13341 (N_13341,N_12006,N_8111);
and U13342 (N_13342,N_7942,N_6611);
and U13343 (N_13343,N_11670,N_9187);
and U13344 (N_13344,N_8968,N_8919);
and U13345 (N_13345,N_10885,N_10543);
and U13346 (N_13346,N_12048,N_10910);
and U13347 (N_13347,N_10238,N_11841);
and U13348 (N_13348,N_12405,N_6397);
or U13349 (N_13349,N_10959,N_11096);
nor U13350 (N_13350,N_12393,N_11813);
and U13351 (N_13351,N_12221,N_8508);
nand U13352 (N_13352,N_12424,N_9708);
nand U13353 (N_13353,N_9094,N_11386);
and U13354 (N_13354,N_11754,N_12039);
or U13355 (N_13355,N_9425,N_11547);
nand U13356 (N_13356,N_11871,N_6598);
or U13357 (N_13357,N_8459,N_7163);
or U13358 (N_13358,N_7683,N_8159);
and U13359 (N_13359,N_11973,N_8263);
or U13360 (N_13360,N_11985,N_9667);
and U13361 (N_13361,N_7431,N_6393);
nor U13362 (N_13362,N_8398,N_8445);
xor U13363 (N_13363,N_11352,N_10702);
or U13364 (N_13364,N_7405,N_8659);
or U13365 (N_13365,N_10473,N_10254);
nand U13366 (N_13366,N_8776,N_10279);
nand U13367 (N_13367,N_9389,N_12085);
or U13368 (N_13368,N_11596,N_6580);
xor U13369 (N_13369,N_11015,N_8254);
or U13370 (N_13370,N_7751,N_7422);
or U13371 (N_13371,N_12232,N_12301);
or U13372 (N_13372,N_11112,N_7556);
and U13373 (N_13373,N_10262,N_8880);
or U13374 (N_13374,N_10773,N_10565);
or U13375 (N_13375,N_6689,N_9543);
nor U13376 (N_13376,N_6509,N_12230);
nand U13377 (N_13377,N_10405,N_12410);
nor U13378 (N_13378,N_7660,N_7858);
nor U13379 (N_13379,N_8011,N_7570);
and U13380 (N_13380,N_11406,N_10953);
nand U13381 (N_13381,N_11854,N_10082);
or U13382 (N_13382,N_9910,N_11600);
nor U13383 (N_13383,N_6250,N_7613);
nor U13384 (N_13384,N_7112,N_10804);
nor U13385 (N_13385,N_9588,N_9891);
nor U13386 (N_13386,N_8208,N_8653);
or U13387 (N_13387,N_7971,N_6311);
nand U13388 (N_13388,N_6506,N_9273);
nor U13389 (N_13389,N_12177,N_11964);
and U13390 (N_13390,N_7424,N_11424);
and U13391 (N_13391,N_10961,N_10452);
or U13392 (N_13392,N_11686,N_9384);
nand U13393 (N_13393,N_11217,N_7844);
or U13394 (N_13394,N_11172,N_7478);
nor U13395 (N_13395,N_6817,N_7427);
or U13396 (N_13396,N_9058,N_7229);
or U13397 (N_13397,N_10323,N_8588);
or U13398 (N_13398,N_10579,N_10009);
and U13399 (N_13399,N_10947,N_7338);
and U13400 (N_13400,N_12089,N_7447);
nor U13401 (N_13401,N_10127,N_9195);
nand U13402 (N_13402,N_11207,N_11968);
or U13403 (N_13403,N_9822,N_11920);
nand U13404 (N_13404,N_8255,N_11236);
or U13405 (N_13405,N_9970,N_12487);
and U13406 (N_13406,N_6591,N_10409);
and U13407 (N_13407,N_7413,N_6958);
xnor U13408 (N_13408,N_11598,N_8277);
and U13409 (N_13409,N_8244,N_11571);
nand U13410 (N_13410,N_11307,N_8468);
nand U13411 (N_13411,N_11354,N_8480);
nor U13412 (N_13412,N_12017,N_9419);
or U13413 (N_13413,N_9494,N_10269);
nor U13414 (N_13414,N_7320,N_6951);
nand U13415 (N_13415,N_9666,N_12137);
xnor U13416 (N_13416,N_11026,N_7068);
nor U13417 (N_13417,N_10468,N_10600);
or U13418 (N_13418,N_9955,N_11566);
nand U13419 (N_13419,N_12300,N_6425);
nand U13420 (N_13420,N_6839,N_12269);
nor U13421 (N_13421,N_8049,N_11978);
nor U13422 (N_13422,N_7695,N_10132);
and U13423 (N_13423,N_10440,N_6407);
and U13424 (N_13424,N_11652,N_10948);
and U13425 (N_13425,N_9685,N_9376);
or U13426 (N_13426,N_6899,N_10365);
nand U13427 (N_13427,N_10301,N_8098);
nand U13428 (N_13428,N_10334,N_8687);
or U13429 (N_13429,N_8488,N_9133);
or U13430 (N_13430,N_6932,N_6769);
nand U13431 (N_13431,N_11763,N_10649);
nor U13432 (N_13432,N_12384,N_8425);
or U13433 (N_13433,N_8898,N_11374);
or U13434 (N_13434,N_10153,N_8296);
or U13435 (N_13435,N_7030,N_9211);
or U13436 (N_13436,N_6822,N_6962);
xnor U13437 (N_13437,N_8008,N_6868);
nand U13438 (N_13438,N_7395,N_7836);
nor U13439 (N_13439,N_9982,N_10917);
or U13440 (N_13440,N_11853,N_10252);
or U13441 (N_13441,N_7230,N_8050);
xnor U13442 (N_13442,N_12344,N_8080);
or U13443 (N_13443,N_9240,N_11248);
and U13444 (N_13444,N_7337,N_7967);
nand U13445 (N_13445,N_12026,N_9788);
and U13446 (N_13446,N_8815,N_9035);
nand U13447 (N_13447,N_9825,N_12284);
and U13448 (N_13448,N_9729,N_8467);
nand U13449 (N_13449,N_11923,N_10879);
nand U13450 (N_13450,N_8778,N_10668);
xnor U13451 (N_13451,N_7656,N_11980);
or U13452 (N_13452,N_6321,N_9496);
nand U13453 (N_13453,N_12008,N_9944);
nor U13454 (N_13454,N_7652,N_6902);
and U13455 (N_13455,N_12158,N_11536);
nor U13456 (N_13456,N_9568,N_7547);
xor U13457 (N_13457,N_9295,N_8877);
xor U13458 (N_13458,N_8224,N_12374);
nand U13459 (N_13459,N_7954,N_7489);
xor U13460 (N_13460,N_7690,N_10825);
nor U13461 (N_13461,N_10460,N_12134);
nand U13462 (N_13462,N_10297,N_10604);
nand U13463 (N_13463,N_10506,N_12381);
nand U13464 (N_13464,N_8389,N_9993);
nor U13465 (N_13465,N_11512,N_8986);
nand U13466 (N_13466,N_9361,N_11698);
xor U13467 (N_13467,N_9852,N_7365);
and U13468 (N_13468,N_11593,N_9562);
nor U13469 (N_13469,N_6332,N_8495);
or U13470 (N_13470,N_8746,N_7303);
and U13471 (N_13471,N_7558,N_9925);
nand U13472 (N_13472,N_8109,N_9315);
xor U13473 (N_13473,N_10065,N_12246);
or U13474 (N_13474,N_10139,N_9180);
and U13475 (N_13475,N_6504,N_12217);
xnor U13476 (N_13476,N_11661,N_10482);
and U13477 (N_13477,N_9210,N_6695);
and U13478 (N_13478,N_10085,N_10721);
nor U13479 (N_13479,N_8926,N_9590);
xor U13480 (N_13480,N_8710,N_7440);
nand U13481 (N_13481,N_9723,N_9363);
or U13482 (N_13482,N_8048,N_9712);
or U13483 (N_13483,N_11899,N_10125);
and U13484 (N_13484,N_11780,N_8982);
nand U13485 (N_13485,N_12178,N_9355);
nor U13486 (N_13486,N_9033,N_7831);
nor U13487 (N_13487,N_8594,N_6977);
nor U13488 (N_13488,N_9963,N_11064);
and U13489 (N_13489,N_11242,N_12306);
and U13490 (N_13490,N_7115,N_10575);
nor U13491 (N_13491,N_9360,N_6766);
nor U13492 (N_13492,N_9455,N_10727);
nor U13493 (N_13493,N_9621,N_10305);
or U13494 (N_13494,N_9124,N_10511);
or U13495 (N_13495,N_7812,N_11370);
and U13496 (N_13496,N_6857,N_6589);
nand U13497 (N_13497,N_6616,N_11895);
and U13498 (N_13498,N_6399,N_8846);
and U13499 (N_13499,N_7937,N_8027);
nor U13500 (N_13500,N_7351,N_9307);
or U13501 (N_13501,N_11257,N_8810);
nor U13502 (N_13502,N_8715,N_11449);
nor U13503 (N_13503,N_7927,N_10582);
and U13504 (N_13504,N_9283,N_8383);
or U13505 (N_13505,N_6712,N_7992);
nand U13506 (N_13506,N_8802,N_10783);
and U13507 (N_13507,N_6291,N_7993);
xnor U13508 (N_13508,N_11789,N_8971);
and U13509 (N_13509,N_6993,N_6499);
nor U13510 (N_13510,N_12082,N_7559);
nand U13511 (N_13511,N_11791,N_10962);
xnor U13512 (N_13512,N_9449,N_7999);
or U13513 (N_13513,N_7553,N_11212);
nand U13514 (N_13514,N_9868,N_9587);
nand U13515 (N_13515,N_10434,N_9284);
nand U13516 (N_13516,N_8681,N_11502);
nand U13517 (N_13517,N_10014,N_8951);
and U13518 (N_13518,N_9560,N_12192);
nor U13519 (N_13519,N_10735,N_7461);
and U13520 (N_13520,N_6306,N_7497);
xor U13521 (N_13521,N_8537,N_11890);
and U13522 (N_13522,N_10335,N_11061);
and U13523 (N_13523,N_8219,N_8139);
nor U13524 (N_13524,N_7856,N_9269);
nand U13525 (N_13525,N_12136,N_8605);
nand U13526 (N_13526,N_10621,N_6548);
or U13527 (N_13527,N_8503,N_6454);
or U13528 (N_13528,N_10399,N_8044);
nor U13529 (N_13529,N_9115,N_11940);
or U13530 (N_13530,N_8261,N_7277);
xnor U13531 (N_13531,N_6313,N_9065);
nand U13532 (N_13532,N_9987,N_7813);
and U13533 (N_13533,N_6495,N_10245);
nand U13534 (N_13534,N_10284,N_11429);
or U13535 (N_13535,N_9007,N_6600);
or U13536 (N_13536,N_10364,N_7612);
and U13537 (N_13537,N_9190,N_9056);
and U13538 (N_13538,N_6429,N_8038);
xor U13539 (N_13539,N_6470,N_10662);
or U13540 (N_13540,N_11046,N_7912);
or U13541 (N_13541,N_7521,N_8432);
or U13542 (N_13542,N_12275,N_11119);
nor U13543 (N_13543,N_11360,N_12009);
nand U13544 (N_13544,N_11716,N_7309);
and U13545 (N_13545,N_11332,N_12276);
nand U13546 (N_13546,N_9149,N_7001);
and U13547 (N_13547,N_7401,N_8673);
nor U13548 (N_13548,N_8698,N_11843);
and U13549 (N_13549,N_8515,N_10126);
xnor U13550 (N_13550,N_12391,N_7565);
nor U13551 (N_13551,N_10100,N_7311);
or U13552 (N_13552,N_7691,N_8010);
or U13553 (N_13553,N_8335,N_10992);
nand U13554 (N_13554,N_6427,N_9259);
nand U13555 (N_13555,N_9829,N_6275);
and U13556 (N_13556,N_7178,N_11766);
and U13557 (N_13557,N_8153,N_10224);
nor U13558 (N_13558,N_8396,N_8308);
nand U13559 (N_13559,N_11622,N_8101);
xnor U13560 (N_13560,N_7280,N_9515);
and U13561 (N_13561,N_8434,N_9452);
nand U13562 (N_13562,N_6502,N_11193);
and U13563 (N_13563,N_9793,N_10818);
xor U13564 (N_13564,N_12169,N_10626);
nand U13565 (N_13565,N_6904,N_10187);
or U13566 (N_13566,N_10394,N_12456);
nand U13567 (N_13567,N_11211,N_7125);
and U13568 (N_13568,N_7733,N_7150);
nand U13569 (N_13569,N_6760,N_12226);
nand U13570 (N_13570,N_9934,N_12049);
and U13571 (N_13571,N_6630,N_7261);
or U13572 (N_13572,N_10105,N_8593);
nand U13573 (N_13573,N_6821,N_8126);
nand U13574 (N_13574,N_10076,N_12102);
or U13575 (N_13575,N_11340,N_9540);
xnor U13576 (N_13576,N_11423,N_10833);
and U13577 (N_13577,N_8958,N_10404);
nand U13578 (N_13578,N_10703,N_11933);
or U13579 (N_13579,N_11838,N_10350);
or U13580 (N_13580,N_6885,N_8532);
nand U13581 (N_13581,N_10675,N_6254);
xnor U13582 (N_13582,N_8777,N_11591);
nor U13583 (N_13583,N_9736,N_9546);
nand U13584 (N_13584,N_10389,N_9640);
or U13585 (N_13585,N_11190,N_7402);
and U13586 (N_13586,N_12151,N_6891);
nor U13587 (N_13587,N_10287,N_10967);
or U13588 (N_13588,N_6795,N_11995);
or U13589 (N_13589,N_9117,N_12395);
and U13590 (N_13590,N_7641,N_12377);
xor U13591 (N_13591,N_11610,N_8274);
nor U13592 (N_13592,N_11357,N_11820);
nand U13593 (N_13593,N_7908,N_7542);
nand U13594 (N_13594,N_7543,N_10087);
and U13595 (N_13595,N_6450,N_8835);
or U13596 (N_13596,N_8148,N_10628);
nor U13597 (N_13597,N_10620,N_6920);
nor U13598 (N_13598,N_11078,N_9218);
nor U13599 (N_13599,N_12204,N_8179);
xor U13600 (N_13600,N_12477,N_6808);
or U13601 (N_13601,N_9327,N_8521);
nor U13602 (N_13602,N_6974,N_7036);
or U13603 (N_13603,N_7168,N_8584);
nor U13604 (N_13604,N_10196,N_8945);
nand U13605 (N_13605,N_9498,N_12280);
or U13606 (N_13606,N_11295,N_10587);
or U13607 (N_13607,N_7272,N_6383);
or U13608 (N_13608,N_11956,N_10425);
xor U13609 (N_13609,N_7446,N_11699);
xnor U13610 (N_13610,N_8650,N_10168);
and U13611 (N_13611,N_8952,N_11896);
or U13612 (N_13612,N_8484,N_7878);
or U13613 (N_13613,N_6664,N_11960);
nand U13614 (N_13614,N_10832,N_10669);
xor U13615 (N_13615,N_9398,N_7238);
and U13616 (N_13616,N_6315,N_12236);
and U13617 (N_13617,N_9657,N_11809);
or U13618 (N_13618,N_10874,N_8266);
and U13619 (N_13619,N_11314,N_10406);
xnor U13620 (N_13620,N_9070,N_10222);
nor U13621 (N_13621,N_8903,N_12490);
and U13622 (N_13622,N_9337,N_9252);
and U13623 (N_13623,N_9771,N_9823);
and U13624 (N_13624,N_12184,N_7775);
or U13625 (N_13625,N_6365,N_8155);
nand U13626 (N_13626,N_7241,N_6656);
and U13627 (N_13627,N_11900,N_8077);
and U13628 (N_13628,N_8093,N_8550);
and U13629 (N_13629,N_8686,N_10346);
or U13630 (N_13630,N_11915,N_9833);
nor U13631 (N_13631,N_8246,N_6933);
nand U13632 (N_13632,N_11876,N_6287);
or U13633 (N_13633,N_11349,N_11178);
nor U13634 (N_13634,N_6863,N_10432);
nand U13635 (N_13635,N_12033,N_7050);
and U13636 (N_13636,N_9900,N_8119);
xnor U13637 (N_13637,N_11004,N_7985);
and U13638 (N_13638,N_10231,N_10670);
or U13639 (N_13639,N_10985,N_8043);
nand U13640 (N_13640,N_10135,N_7629);
nor U13641 (N_13641,N_11150,N_10685);
xor U13642 (N_13642,N_10617,N_8902);
nand U13643 (N_13643,N_11292,N_8428);
nor U13644 (N_13644,N_7693,N_11251);
nand U13645 (N_13645,N_8932,N_7837);
or U13646 (N_13646,N_8385,N_9157);
nor U13647 (N_13647,N_12144,N_7097);
or U13648 (N_13648,N_8239,N_9622);
or U13649 (N_13649,N_7741,N_11760);
nor U13650 (N_13650,N_6972,N_8862);
nand U13651 (N_13651,N_11312,N_8966);
nor U13652 (N_13652,N_7376,N_8772);
nor U13653 (N_13653,N_9878,N_11516);
nand U13654 (N_13654,N_10289,N_9765);
nor U13655 (N_13655,N_12329,N_8625);
and U13656 (N_13656,N_12488,N_7140);
nor U13657 (N_13657,N_6990,N_10047);
nand U13658 (N_13658,N_6937,N_6536);
nand U13659 (N_13659,N_11731,N_8894);
nand U13660 (N_13660,N_6723,N_11289);
and U13661 (N_13661,N_7839,N_7566);
and U13662 (N_13662,N_10154,N_7879);
nand U13663 (N_13663,N_8371,N_9308);
or U13664 (N_13664,N_7468,N_11863);
nand U13665 (N_13665,N_6496,N_12172);
nor U13666 (N_13666,N_6587,N_7488);
nand U13667 (N_13667,N_7455,N_9168);
xor U13668 (N_13668,N_12104,N_8950);
xor U13669 (N_13669,N_8774,N_9450);
nand U13670 (N_13670,N_8730,N_6423);
and U13671 (N_13671,N_10018,N_12098);
and U13672 (N_13672,N_9105,N_7592);
nand U13673 (N_13673,N_7776,N_7939);
and U13674 (N_13674,N_10523,N_7165);
nor U13675 (N_13675,N_12182,N_7323);
and U13676 (N_13676,N_10235,N_9827);
nand U13677 (N_13677,N_7860,N_12013);
nand U13678 (N_13678,N_11497,N_12261);
and U13679 (N_13679,N_9851,N_9091);
nand U13680 (N_13680,N_10893,N_9401);
xor U13681 (N_13681,N_10093,N_10181);
nor U13682 (N_13682,N_10112,N_8129);
or U13683 (N_13683,N_9744,N_11285);
nor U13684 (N_13684,N_9951,N_7367);
nor U13685 (N_13685,N_11946,N_6909);
nor U13686 (N_13686,N_8519,N_7087);
xor U13687 (N_13687,N_11690,N_6672);
or U13688 (N_13688,N_8867,N_7807);
nand U13689 (N_13689,N_7218,N_6813);
and U13690 (N_13690,N_7132,N_9767);
nor U13691 (N_13691,N_9885,N_7921);
or U13692 (N_13692,N_8751,N_7694);
xor U13693 (N_13693,N_7135,N_8055);
or U13694 (N_13694,N_6679,N_8676);
and U13695 (N_13695,N_6312,N_8359);
and U13696 (N_13696,N_8380,N_7538);
nor U13697 (N_13697,N_9949,N_11186);
nor U13698 (N_13698,N_11115,N_8562);
nand U13699 (N_13699,N_11219,N_10290);
or U13700 (N_13700,N_9980,N_11025);
nand U13701 (N_13701,N_6893,N_7784);
nand U13702 (N_13702,N_9143,N_10686);
or U13703 (N_13703,N_7414,N_11939);
or U13704 (N_13704,N_11831,N_7251);
and U13705 (N_13705,N_6914,N_10586);
nor U13706 (N_13706,N_10779,N_10694);
or U13707 (N_13707,N_10348,N_8302);
and U13708 (N_13708,N_11230,N_6934);
or U13709 (N_13709,N_6936,N_12373);
nand U13710 (N_13710,N_10743,N_7285);
nand U13711 (N_13711,N_8450,N_7428);
or U13712 (N_13712,N_12482,N_10166);
or U13713 (N_13713,N_8612,N_11868);
nand U13714 (N_13714,N_7208,N_12357);
or U13715 (N_13715,N_12291,N_11916);
xnor U13716 (N_13716,N_8237,N_6538);
or U13717 (N_13717,N_10326,N_11727);
or U13718 (N_13718,N_8402,N_11037);
nor U13719 (N_13719,N_11821,N_6634);
nand U13720 (N_13720,N_10990,N_9443);
nor U13721 (N_13721,N_8553,N_12043);
and U13722 (N_13722,N_11267,N_7511);
and U13723 (N_13723,N_8719,N_11087);
nand U13724 (N_13724,N_9914,N_11208);
nor U13725 (N_13725,N_7154,N_7951);
and U13726 (N_13726,N_8133,N_7120);
nor U13727 (N_13727,N_9968,N_12107);
and U13728 (N_13728,N_6688,N_9106);
nand U13729 (N_13729,N_10828,N_7074);
and U13730 (N_13730,N_9791,N_12418);
nand U13731 (N_13731,N_7616,N_6734);
and U13732 (N_13732,N_9627,N_11924);
nor U13733 (N_13733,N_8560,N_9415);
nor U13734 (N_13734,N_6498,N_10338);
or U13735 (N_13735,N_6896,N_9215);
nor U13736 (N_13736,N_6952,N_11825);
and U13737 (N_13737,N_10246,N_12238);
and U13738 (N_13738,N_8808,N_10809);
and U13739 (N_13739,N_10354,N_6996);
or U13740 (N_13740,N_9357,N_11722);
or U13741 (N_13741,N_11097,N_10420);
nor U13742 (N_13742,N_9542,N_9867);
and U13743 (N_13743,N_8175,N_11321);
xor U13744 (N_13744,N_10716,N_10549);
xor U13745 (N_13745,N_11063,N_8373);
and U13746 (N_13746,N_10672,N_11014);
nor U13747 (N_13747,N_10411,N_8031);
nor U13748 (N_13748,N_7871,N_12351);
or U13749 (N_13749,N_11811,N_12229);
xnor U13750 (N_13750,N_6959,N_10186);
and U13751 (N_13751,N_9511,N_12399);
or U13752 (N_13752,N_11666,N_8766);
or U13753 (N_13753,N_11282,N_12499);
nand U13754 (N_13754,N_10249,N_11012);
or U13755 (N_13755,N_9888,N_9709);
nor U13756 (N_13756,N_8168,N_10239);
and U13757 (N_13757,N_11447,N_9533);
nand U13758 (N_13758,N_9055,N_9816);
and U13759 (N_13759,N_8791,N_7170);
nor U13760 (N_13760,N_9132,N_12486);
or U13761 (N_13761,N_12046,N_6583);
nor U13762 (N_13762,N_11428,N_8705);
nor U13763 (N_13763,N_8933,N_11750);
or U13764 (N_13764,N_8569,N_7636);
and U13765 (N_13765,N_10037,N_9191);
nor U13766 (N_13766,N_9789,N_10138);
nand U13767 (N_13767,N_10507,N_10164);
or U13768 (N_13768,N_8037,N_9988);
or U13769 (N_13769,N_6542,N_12338);
or U13770 (N_13770,N_9732,N_6645);
and U13771 (N_13771,N_9402,N_12110);
and U13772 (N_13772,N_6285,N_7189);
nor U13773 (N_13773,N_6978,N_10954);
or U13774 (N_13774,N_11180,N_6350);
or U13775 (N_13775,N_6758,N_6528);
nor U13776 (N_13776,N_11040,N_10309);
xor U13777 (N_13777,N_7374,N_9946);
and U13778 (N_13778,N_8756,N_9894);
and U13779 (N_13779,N_11095,N_6953);
nor U13780 (N_13780,N_8890,N_10974);
nand U13781 (N_13781,N_11500,N_11400);
or U13782 (N_13782,N_7334,N_6453);
nor U13783 (N_13783,N_8864,N_10728);
nor U13784 (N_13784,N_9328,N_6614);
and U13785 (N_13785,N_8469,N_8587);
or U13786 (N_13786,N_11673,N_11656);
nor U13787 (N_13787,N_6568,N_8269);
and U13788 (N_13788,N_10091,N_10226);
xor U13789 (N_13789,N_7972,N_10480);
nor U13790 (N_13790,N_6422,N_8740);
nor U13791 (N_13791,N_8192,N_7540);
and U13792 (N_13792,N_7672,N_9926);
and U13793 (N_13793,N_7757,N_7744);
or U13794 (N_13794,N_11434,N_8060);
and U13795 (N_13795,N_9167,N_8571);
and U13796 (N_13796,N_6715,N_6457);
or U13797 (N_13797,N_8276,N_8353);
nor U13798 (N_13798,N_11122,N_8627);
nand U13799 (N_13799,N_6438,N_12283);
or U13800 (N_13800,N_9865,N_6461);
or U13801 (N_13801,N_7567,N_6637);
nor U13802 (N_13802,N_9096,N_7564);
or U13803 (N_13803,N_11873,N_6718);
nand U13804 (N_13804,N_7832,N_12143);
nand U13805 (N_13805,N_10261,N_10147);
nand U13806 (N_13806,N_8800,N_6682);
or U13807 (N_13807,N_9072,N_8178);
nand U13808 (N_13808,N_10214,N_11485);
nand U13809 (N_13809,N_11902,N_10697);
xor U13810 (N_13810,N_8448,N_7767);
nand U13811 (N_13811,N_6353,N_10663);
or U13812 (N_13812,N_8872,N_9285);
nor U13813 (N_13813,N_7979,N_10336);
or U13814 (N_13814,N_6818,N_6309);
nand U13815 (N_13815,N_11380,N_8214);
nor U13816 (N_13816,N_12139,N_12233);
and U13817 (N_13817,N_7471,N_7032);
and U13818 (N_13818,N_11255,N_8540);
xor U13819 (N_13819,N_6582,N_10211);
nor U13820 (N_13820,N_9608,N_12130);
nor U13821 (N_13821,N_10457,N_12415);
or U13822 (N_13822,N_12353,N_7111);
and U13823 (N_13823,N_9044,N_6307);
nand U13824 (N_13824,N_8478,N_11468);
nor U13825 (N_13825,N_6330,N_6898);
nand U13826 (N_13826,N_10314,N_9102);
nor U13827 (N_13827,N_10328,N_9785);
and U13828 (N_13828,N_9735,N_8113);
nor U13829 (N_13829,N_9694,N_10678);
nor U13830 (N_13830,N_9074,N_11556);
and U13831 (N_13831,N_9585,N_12398);
and U13832 (N_13832,N_6512,N_10740);
nor U13833 (N_13833,N_7191,N_8144);
and U13834 (N_13834,N_7742,N_9876);
nand U13835 (N_13835,N_7255,N_8738);
nand U13836 (N_13836,N_10142,N_11011);
nor U13837 (N_13837,N_8074,N_6398);
nand U13838 (N_13838,N_12392,N_10517);
nor U13839 (N_13839,N_6687,N_6521);
nand U13840 (N_13840,N_6747,N_8970);
and U13841 (N_13841,N_10263,N_7256);
nor U13842 (N_13842,N_10375,N_8207);
nand U13843 (N_13843,N_8635,N_8911);
and U13844 (N_13844,N_10777,N_11319);
or U13845 (N_13845,N_7821,N_6668);
nor U13846 (N_13846,N_9646,N_11621);
or U13847 (N_13847,N_11315,N_7626);
xor U13848 (N_13848,N_7340,N_9715);
nor U13849 (N_13849,N_7375,N_8655);
nand U13850 (N_13850,N_11262,N_12058);
or U13851 (N_13851,N_6994,N_6834);
nand U13852 (N_13852,N_10223,N_11531);
or U13853 (N_13853,N_10913,N_7569);
nand U13854 (N_13854,N_12468,N_9531);
nand U13855 (N_13855,N_8830,N_8812);
nor U13856 (N_13856,N_9330,N_8853);
nand U13857 (N_13857,N_6746,N_7174);
nand U13858 (N_13858,N_6803,N_7018);
and U13859 (N_13859,N_7031,N_11454);
nor U13860 (N_13860,N_9844,N_12349);
and U13861 (N_13861,N_9530,N_11952);
nand U13862 (N_13862,N_10712,N_7169);
or U13863 (N_13863,N_9297,N_10645);
or U13864 (N_13864,N_6823,N_7104);
nor U13865 (N_13865,N_10038,N_10607);
xnor U13866 (N_13866,N_9080,N_9859);
nor U13867 (N_13867,N_11043,N_10826);
and U13868 (N_13868,N_10116,N_7531);
xnor U13869 (N_13869,N_7893,N_9118);
nor U13870 (N_13870,N_10863,N_11774);
xnor U13871 (N_13871,N_8677,N_11703);
xor U13872 (N_13872,N_12176,N_7815);
nand U13873 (N_13873,N_8298,N_8474);
or U13874 (N_13874,N_6581,N_8286);
and U13875 (N_13875,N_9624,N_6654);
nand U13876 (N_13876,N_10561,N_11728);
and U13877 (N_13877,N_11085,N_7071);
or U13878 (N_13878,N_12149,N_8410);
xnor U13879 (N_13879,N_7248,N_8976);
and U13880 (N_13880,N_8241,N_11055);
xor U13881 (N_13881,N_7709,N_10855);
nor U13882 (N_13882,N_11214,N_10242);
nor U13883 (N_13883,N_10109,N_8845);
or U13884 (N_13884,N_11653,N_7386);
xor U13885 (N_13885,N_10815,N_10383);
nor U13886 (N_13886,N_10802,N_9460);
and U13887 (N_13887,N_6731,N_7296);
nor U13888 (N_13888,N_9882,N_10614);
and U13889 (N_13889,N_9179,N_6460);
or U13890 (N_13890,N_11451,N_9508);
nor U13891 (N_13891,N_10513,N_7180);
nand U13892 (N_13892,N_11941,N_6950);
and U13893 (N_13893,N_7397,N_8697);
nand U13894 (N_13894,N_10525,N_11032);
or U13895 (N_13895,N_9475,N_8918);
nor U13896 (N_13896,N_7235,N_10442);
nand U13897 (N_13897,N_7730,N_9578);
nand U13898 (N_13898,N_10674,N_12190);
nor U13899 (N_13899,N_10288,N_9545);
and U13900 (N_13900,N_11804,N_9941);
nand U13901 (N_13901,N_6501,N_7384);
nor U13902 (N_13902,N_7333,N_10073);
and U13903 (N_13903,N_10015,N_11579);
nand U13904 (N_13904,N_8342,N_9459);
or U13905 (N_13905,N_12138,N_10781);
and U13906 (N_13906,N_6989,N_10521);
xor U13907 (N_13907,N_10466,N_11798);
xor U13908 (N_13908,N_8367,N_8668);
nand U13909 (N_13909,N_6541,N_9873);
nor U13910 (N_13910,N_10538,N_9992);
nand U13911 (N_13911,N_8980,N_9676);
and U13912 (N_13912,N_9138,N_10079);
nand U13913 (N_13913,N_8372,N_7962);
nand U13914 (N_13914,N_10021,N_7786);
nand U13915 (N_13915,N_11658,N_8623);
nor U13916 (N_13916,N_7083,N_9436);
nand U13917 (N_13917,N_11800,N_7697);
nand U13918 (N_13918,N_11817,N_6725);
or U13919 (N_13919,N_11245,N_7867);
nor U13920 (N_13920,N_10403,N_12056);
or U13921 (N_13921,N_10771,N_7012);
and U13922 (N_13922,N_8065,N_7310);
or U13923 (N_13923,N_7681,N_12387);
and U13924 (N_13924,N_11564,N_12335);
and U13925 (N_13925,N_11771,N_7315);
or U13926 (N_13926,N_9069,N_11700);
nor U13927 (N_13927,N_7884,N_11839);
or U13928 (N_13928,N_11583,N_7727);
nand U13929 (N_13929,N_12069,N_8843);
nor U13930 (N_13930,N_10846,N_8722);
and U13931 (N_13931,N_9299,N_11496);
nor U13932 (N_13932,N_10596,N_11121);
nand U13933 (N_13933,N_9251,N_9527);
or U13934 (N_13934,N_7109,N_8190);
nor U13935 (N_13935,N_9411,N_11377);
or U13936 (N_13936,N_6534,N_10566);
nor U13937 (N_13937,N_8622,N_10850);
nand U13938 (N_13938,N_10368,N_7221);
nor U13939 (N_13939,N_11522,N_8331);
and U13940 (N_13940,N_12309,N_8987);
and U13941 (N_13941,N_12340,N_9901);
and U13942 (N_13942,N_12114,N_6358);
or U13943 (N_13943,N_9160,N_8020);
nand U13944 (N_13944,N_10377,N_9749);
or U13945 (N_13945,N_9469,N_10000);
nand U13946 (N_13946,N_7408,N_7198);
and U13947 (N_13947,N_12127,N_10951);
xor U13948 (N_13948,N_11322,N_9435);
nor U13949 (N_13949,N_9063,N_6772);
xnor U13950 (N_13950,N_11168,N_11668);
and U13951 (N_13951,N_11788,N_10431);
and U13952 (N_13952,N_10033,N_10603);
xnor U13953 (N_13953,N_8496,N_8866);
or U13954 (N_13954,N_7639,N_7530);
xor U13955 (N_13955,N_11127,N_7529);
xnor U13956 (N_13956,N_6880,N_11490);
nand U13957 (N_13957,N_12267,N_11223);
nand U13958 (N_13958,N_10467,N_8685);
nor U13959 (N_13959,N_7957,N_9563);
nand U13960 (N_13960,N_6783,N_12288);
and U13961 (N_13961,N_11175,N_6724);
or U13962 (N_13962,N_6691,N_7043);
nand U13963 (N_13963,N_7186,N_12342);
nor U13964 (N_13964,N_10778,N_9416);
and U13965 (N_13965,N_10408,N_6707);
xnor U13966 (N_13966,N_8557,N_7398);
or U13967 (N_13967,N_11786,N_7974);
and U13968 (N_13968,N_8437,N_12253);
xnor U13969 (N_13969,N_11494,N_12252);
and U13970 (N_13970,N_9247,N_7129);
or U13971 (N_13971,N_6494,N_7798);
nand U13972 (N_13972,N_11612,N_9813);
nor U13973 (N_13973,N_7603,N_8046);
nand U13974 (N_13974,N_11146,N_8549);
and U13975 (N_13975,N_9280,N_10851);
and U13976 (N_13976,N_11417,N_11350);
xor U13977 (N_13977,N_8997,N_6780);
nand U13978 (N_13978,N_11233,N_12005);
xor U13979 (N_13979,N_10912,N_10128);
nor U13980 (N_13980,N_6329,N_10217);
or U13981 (N_13981,N_7952,N_8967);
nand U13982 (N_13982,N_11910,N_6633);
nor U13983 (N_13983,N_9843,N_11942);
nand U13984 (N_13984,N_11084,N_9341);
or U13985 (N_13985,N_11137,N_7271);
nor U13986 (N_13986,N_12153,N_10527);
or U13987 (N_13987,N_6519,N_10136);
or U13988 (N_13988,N_7456,N_7605);
or U13989 (N_13989,N_11195,N_11080);
or U13990 (N_13990,N_7258,N_9318);
and U13991 (N_13991,N_11601,N_7314);
nor U13992 (N_13992,N_8583,N_8850);
xnor U13993 (N_13993,N_9728,N_11514);
and U13994 (N_13994,N_9345,N_12339);
and U13995 (N_13995,N_8733,N_7173);
nor U13996 (N_13996,N_8355,N_7342);
and U13997 (N_13997,N_7990,N_9272);
or U13998 (N_13998,N_6331,N_8482);
and U13999 (N_13999,N_10320,N_9045);
or U14000 (N_14000,N_7632,N_7390);
nor U14001 (N_14001,N_11135,N_10392);
or U14002 (N_14002,N_8696,N_10011);
and U14003 (N_14003,N_11865,N_6628);
xnor U14004 (N_14004,N_10078,N_11281);
or U14005 (N_14005,N_9254,N_8793);
or U14006 (N_14006,N_11567,N_8348);
or U14007 (N_14007,N_8245,N_10515);
or U14008 (N_14008,N_9939,N_12466);
nand U14009 (N_14009,N_8712,N_10152);
nand U14010 (N_14010,N_6666,N_7096);
nand U14011 (N_14011,N_12362,N_11132);
nor U14012 (N_14012,N_7368,N_10157);
or U14013 (N_14013,N_10560,N_7033);
nor U14014 (N_14014,N_7410,N_11954);
nor U14015 (N_14015,N_9849,N_6262);
nor U14016 (N_14016,N_9887,N_6320);
or U14017 (N_14017,N_9673,N_6728);
nor U14018 (N_14018,N_9857,N_11243);
xnor U14019 (N_14019,N_8626,N_7022);
or U14020 (N_14020,N_10441,N_9856);
and U14021 (N_14021,N_10548,N_12141);
xnor U14022 (N_14022,N_9808,N_8349);
nand U14023 (N_14023,N_11361,N_6267);
and U14024 (N_14024,N_9509,N_6469);
nand U14025 (N_14025,N_11108,N_10202);
and U14026 (N_14026,N_9976,N_6913);
or U14027 (N_14027,N_10715,N_7381);
xnor U14028 (N_14028,N_10821,N_12359);
nand U14029 (N_14029,N_9604,N_10169);
or U14030 (N_14030,N_11848,N_8858);
nor U14031 (N_14031,N_12097,N_12146);
or U14032 (N_14032,N_10748,N_9637);
nor U14033 (N_14033,N_11218,N_10536);
and U14034 (N_14034,N_12059,N_10322);
or U14035 (N_14035,N_6388,N_11395);
nand U14036 (N_14036,N_7560,N_8749);
nor U14037 (N_14037,N_10436,N_12213);
or U14038 (N_14038,N_6270,N_9454);
xnor U14039 (N_14039,N_6609,N_12038);
and U14040 (N_14040,N_11030,N_8770);
nand U14041 (N_14041,N_9783,N_7254);
xnor U14042 (N_14042,N_8718,N_6657);
nand U14043 (N_14043,N_10376,N_10413);
nor U14044 (N_14044,N_10571,N_11171);
xnor U14045 (N_14045,N_10526,N_10944);
and U14046 (N_14046,N_11103,N_7421);
nor U14047 (N_14047,N_10652,N_11381);
nand U14048 (N_14048,N_9199,N_10490);
nand U14049 (N_14049,N_9140,N_7915);
nand U14050 (N_14050,N_8314,N_10426);
or U14051 (N_14051,N_6674,N_8166);
or U14052 (N_14052,N_7378,N_11253);
nor U14053 (N_14053,N_8502,N_9216);
nand U14054 (N_14054,N_7528,N_11408);
nand U14055 (N_14055,N_9964,N_8390);
nand U14056 (N_14056,N_10369,N_9079);
nor U14057 (N_14057,N_7385,N_9010);
and U14058 (N_14058,N_8498,N_9061);
or U14059 (N_14059,N_9931,N_8552);
and U14060 (N_14060,N_6593,N_11486);
nor U14061 (N_14061,N_6894,N_10499);
nand U14062 (N_14062,N_11944,N_9101);
nor U14063 (N_14063,N_10631,N_11252);
nand U14064 (N_14064,N_9577,N_11022);
or U14065 (N_14065,N_8135,N_12124);
or U14066 (N_14066,N_11327,N_11507);
nor U14067 (N_14067,N_10504,N_11709);
nand U14068 (N_14068,N_8427,N_8769);
or U14069 (N_14069,N_7133,N_11625);
nand U14070 (N_14070,N_8724,N_10291);
and U14071 (N_14071,N_8567,N_7576);
and U14072 (N_14072,N_10618,N_7805);
and U14073 (N_14073,N_11396,N_9522);
and U14074 (N_14074,N_7239,N_10813);
nor U14075 (N_14075,N_9276,N_8330);
nand U14076 (N_14076,N_9100,N_10647);
and U14077 (N_14077,N_11353,N_6366);
or U14078 (N_14078,N_7331,N_6781);
and U14079 (N_14079,N_10062,N_6544);
and U14080 (N_14080,N_7960,N_11106);
nor U14081 (N_14081,N_11550,N_10036);
nor U14082 (N_14082,N_12040,N_7841);
nor U14083 (N_14083,N_12034,N_11619);
and U14084 (N_14084,N_7810,N_9405);
or U14085 (N_14085,N_6392,N_9206);
nor U14086 (N_14086,N_11394,N_8861);
nor U14087 (N_14087,N_12074,N_10646);
and U14088 (N_14088,N_9310,N_10915);
or U14089 (N_14089,N_7611,N_8084);
xnor U14090 (N_14090,N_7347,N_7099);
nor U14091 (N_14091,N_9989,N_7976);
or U14092 (N_14092,N_8009,N_7481);
nor U14093 (N_14093,N_10469,N_12260);
nor U14094 (N_14094,N_7149,N_8787);
nor U14095 (N_14095,N_8443,N_9625);
nand U14096 (N_14096,N_10300,N_7433);
nand U14097 (N_14097,N_8988,N_11885);
nand U14098 (N_14098,N_7907,N_11609);
nand U14099 (N_14099,N_9582,N_12077);
nand U14100 (N_14100,N_11075,N_9029);
nand U14101 (N_14101,N_6525,N_8758);
nor U14102 (N_14102,N_7766,N_6371);
nor U14103 (N_14103,N_6468,N_7361);
nor U14104 (N_14104,N_10104,N_12191);
nand U14105 (N_14105,N_12251,N_8460);
and U14106 (N_14106,N_8318,N_9650);
or U14107 (N_14107,N_6923,N_10965);
and U14108 (N_14108,N_10926,N_8490);
nor U14109 (N_14109,N_10359,N_7873);
and U14110 (N_14110,N_8325,N_7264);
xnor U14111 (N_14111,N_7802,N_12367);
or U14112 (N_14112,N_7308,N_9264);
nor U14113 (N_14113,N_10908,N_10807);
or U14114 (N_14114,N_9177,N_9804);
or U14115 (N_14115,N_12336,N_6354);
or U14116 (N_14116,N_8844,N_8404);
nor U14117 (N_14117,N_10881,N_8455);
or U14118 (N_14118,N_11538,N_6830);
and U14119 (N_14119,N_8716,N_6871);
nand U14120 (N_14120,N_10094,N_11562);
and U14121 (N_14121,N_10860,N_9267);
and U14122 (N_14122,N_10756,N_7014);
or U14123 (N_14123,N_11081,N_11463);
nand U14124 (N_14124,N_8663,N_10313);
or U14125 (N_14125,N_12324,N_7584);
and U14126 (N_14126,N_12457,N_8973);
and U14127 (N_14127,N_12354,N_9660);
or U14128 (N_14128,N_11336,N_9059);
nand U14129 (N_14129,N_8182,N_6481);
or U14130 (N_14130,N_9997,N_8662);
nand U14131 (N_14131,N_6503,N_11790);
nand U14132 (N_14132,N_8035,N_11196);
and U14133 (N_14133,N_7100,N_8558);
nand U14134 (N_14134,N_8528,N_8512);
nor U14135 (N_14135,N_6378,N_8001);
or U14136 (N_14136,N_9490,N_6770);
nand U14137 (N_14137,N_8222,N_6805);
and U14138 (N_14138,N_10258,N_11824);
or U14139 (N_14139,N_9840,N_7643);
nand U14140 (N_14140,N_8424,N_10816);
nand U14141 (N_14141,N_6624,N_11264);
or U14142 (N_14142,N_11138,N_12062);
nor U14143 (N_14143,N_8841,N_8645);
xnor U14144 (N_14144,N_7064,N_10687);
or U14145 (N_14145,N_7480,N_12469);
nand U14146 (N_14146,N_7415,N_7725);
nand U14147 (N_14147,N_11832,N_8268);
nand U14148 (N_14148,N_11489,N_9121);
or U14149 (N_14149,N_6324,N_10423);
and U14150 (N_14150,N_12084,N_10090);
or U14151 (N_14151,N_6694,N_9060);
and U14152 (N_14152,N_6841,N_11530);
and U14153 (N_14153,N_8938,N_8114);
nor U14154 (N_14154,N_9665,N_9835);
or U14155 (N_14155,N_11747,N_7947);
xor U14156 (N_14156,N_6364,N_7494);
and U14157 (N_14157,N_12016,N_12030);
nor U14158 (N_14158,N_8760,N_7213);
nor U14159 (N_14159,N_7705,N_7393);
and U14160 (N_14160,N_10054,N_12407);
nand U14161 (N_14161,N_6631,N_7980);
and U14162 (N_14162,N_9165,N_10991);
and U14163 (N_14163,N_11681,N_7035);
nand U14164 (N_14164,N_11277,N_10591);
xnor U14165 (N_14165,N_8611,N_10493);
nand U14166 (N_14166,N_10558,N_7214);
xnor U14167 (N_14167,N_7834,N_7647);
and U14168 (N_14168,N_12036,N_8637);
nand U14169 (N_14169,N_7407,N_9766);
or U14170 (N_14170,N_8358,N_7156);
xnor U14171 (N_14171,N_6508,N_11869);
nor U14172 (N_14172,N_6800,N_6970);
and U14173 (N_14173,N_10280,N_8313);
and U14174 (N_14174,N_12159,N_9456);
or U14175 (N_14175,N_7055,N_9221);
and U14176 (N_14176,N_7816,N_7245);
and U14177 (N_14177,N_9652,N_11794);
nor U14178 (N_14178,N_9611,N_7307);
or U14179 (N_14179,N_10351,N_6802);
nand U14180 (N_14180,N_9477,N_8990);
and U14181 (N_14181,N_11886,N_10553);
nor U14182 (N_14182,N_7204,N_6385);
nand U14183 (N_14183,N_12343,N_12397);
or U14184 (N_14184,N_10554,N_6369);
nand U14185 (N_14185,N_6272,N_8585);
nand U14186 (N_14186,N_11383,N_10601);
nand U14187 (N_14187,N_8889,N_11148);
or U14188 (N_14188,N_9244,N_8639);
xnor U14189 (N_14189,N_7795,N_9281);
and U14190 (N_14190,N_9821,N_8408);
nor U14191 (N_14191,N_8675,N_6252);
nand U14192 (N_14192,N_7364,N_11179);
and U14193 (N_14193,N_8300,N_10363);
nand U14194 (N_14194,N_8832,N_7281);
nor U14195 (N_14195,N_10035,N_6705);
nor U14196 (N_14196,N_11897,N_11947);
or U14197 (N_14197,N_7712,N_8073);
nand U14198 (N_14198,N_7916,N_6284);
nor U14199 (N_14199,N_6886,N_8227);
or U14200 (N_14200,N_11345,N_8632);
or U14201 (N_14201,N_9680,N_8839);
xnor U14202 (N_14202,N_12067,N_7126);
and U14203 (N_14203,N_6845,N_6890);
nand U14204 (N_14204,N_8127,N_7601);
nor U14205 (N_14205,N_12002,N_10256);
nor U14206 (N_14206,N_6748,N_8929);
xor U14207 (N_14207,N_9756,N_8607);
nor U14208 (N_14208,N_11431,N_7117);
nand U14209 (N_14209,N_9162,N_10016);
and U14210 (N_14210,N_9917,N_9175);
or U14211 (N_14211,N_7040,N_6584);
nand U14212 (N_14212,N_8036,N_6571);
xnor U14213 (N_14213,N_11372,N_10623);
or U14214 (N_14214,N_10317,N_10257);
or U14215 (N_14215,N_10243,N_10510);
xnor U14216 (N_14216,N_9194,N_8599);
nand U14217 (N_14217,N_9316,N_10184);
and U14218 (N_14218,N_9220,N_7548);
nor U14219 (N_14219,N_7920,N_7578);
nor U14220 (N_14220,N_9617,N_11743);
and U14221 (N_14221,N_8250,N_11101);
and U14222 (N_14222,N_10986,N_8604);
and U14223 (N_14223,N_10422,N_7197);
nand U14224 (N_14224,N_8461,N_8360);
nor U14225 (N_14225,N_11271,N_8969);
xnor U14226 (N_14226,N_7294,N_7679);
nand U14227 (N_14227,N_10857,N_10508);
nor U14228 (N_14228,N_10456,N_9909);
nor U14229 (N_14229,N_6585,N_10952);
nor U14230 (N_14230,N_11822,N_7144);
nand U14231 (N_14231,N_8831,N_10447);
nor U14232 (N_14232,N_11265,N_6462);
nor U14233 (N_14233,N_11294,N_10580);
and U14234 (N_14234,N_10635,N_10312);
nor U14235 (N_14235,N_10892,N_10696);
and U14236 (N_14236,N_11568,N_12345);
or U14237 (N_14237,N_9009,N_11210);
xnor U14238 (N_14238,N_9150,N_9805);
and U14239 (N_14239,N_8752,N_8350);
xor U14240 (N_14240,N_8258,N_7038);
nand U14241 (N_14241,N_8566,N_7098);
and U14242 (N_14242,N_7702,N_9592);
nand U14243 (N_14243,N_7994,N_7373);
nand U14244 (N_14244,N_7295,N_10067);
nand U14245 (N_14245,N_6564,N_7801);
nor U14246 (N_14246,N_8991,N_12467);
or U14247 (N_14247,N_11660,N_10121);
and U14248 (N_14248,N_10555,N_9551);
nand U14249 (N_14249,N_7448,N_9016);
and U14250 (N_14250,N_7435,N_9537);
or U14251 (N_14251,N_10624,N_10362);
nor U14252 (N_14252,N_8764,N_6998);
nor U14253 (N_14253,N_10144,N_9386);
or U14254 (N_14254,N_11126,N_8617);
nand U14255 (N_14255,N_10034,N_10160);
xnor U14256 (N_14256,N_10980,N_11476);
nand U14257 (N_14257,N_12286,N_7561);
nand U14258 (N_14258,N_9166,N_11154);
nand U14259 (N_14259,N_9595,N_10920);
nor U14260 (N_14260,N_7973,N_9329);
nor U14261 (N_14261,N_10248,N_11375);
or U14262 (N_14262,N_9748,N_6919);
nor U14263 (N_14263,N_11967,N_8141);
or U14264 (N_14264,N_7228,N_10200);
nor U14265 (N_14265,N_10505,N_9638);
nand U14266 (N_14266,N_9747,N_10435);
or U14267 (N_14267,N_6344,N_9656);
nand U14268 (N_14268,N_6988,N_10729);
nand U14269 (N_14269,N_9184,N_12473);
xnor U14270 (N_14270,N_9996,N_12020);
and U14271 (N_14271,N_8591,N_10732);
and U14272 (N_14272,N_12451,N_6764);
nand U14273 (N_14273,N_10547,N_9174);
or U14274 (N_14274,N_10424,N_7404);
xor U14275 (N_14275,N_9286,N_7958);
xor U14276 (N_14276,N_7291,N_11908);
or U14277 (N_14277,N_8786,N_12431);
nand U14278 (N_14278,N_12111,N_9326);
nor U14279 (N_14279,N_10298,N_7621);
nor U14280 (N_14280,N_8708,N_12199);
nor U14281 (N_14281,N_7595,N_10449);
and U14282 (N_14282,N_6792,N_12254);
and U14283 (N_14283,N_10225,N_6515);
or U14284 (N_14284,N_7454,N_9547);
nor U14285 (N_14285,N_6594,N_9773);
nor U14286 (N_14286,N_8960,N_11552);
or U14287 (N_14287,N_12421,N_11862);
or U14288 (N_14288,N_6690,N_7142);
nand U14289 (N_14289,N_6973,N_9752);
and U14290 (N_14290,N_7122,N_11020);
xor U14291 (N_14291,N_9289,N_8321);
and U14292 (N_14292,N_8489,N_11068);
nand U14293 (N_14293,N_12420,N_7225);
and U14294 (N_14294,N_6412,N_9053);
or U14295 (N_14295,N_11268,N_8413);
nor U14296 (N_14296,N_11977,N_9087);
nor U14297 (N_14297,N_7108,N_6761);
nand U14298 (N_14298,N_8559,N_11003);
or U14299 (N_14299,N_10785,N_9512);
nand U14300 (N_14300,N_7181,N_10654);
or U14301 (N_14301,N_8807,N_11356);
nor U14302 (N_14302,N_9414,N_10840);
xor U14303 (N_14303,N_9492,N_8819);
nand U14304 (N_14304,N_6963,N_10019);
or U14305 (N_14305,N_11725,N_7526);
or U14306 (N_14306,N_6484,N_10900);
nand U14307 (N_14307,N_8392,N_8768);
or U14308 (N_14308,N_11719,N_11074);
nand U14309 (N_14309,N_12316,N_8925);
and U14310 (N_14310,N_6547,N_12256);
nor U14311 (N_14311,N_9798,N_9855);
nand U14312 (N_14312,N_12079,N_11416);
or U14313 (N_14313,N_12277,N_10784);
nor U14314 (N_14314,N_9519,N_10197);
and U14315 (N_14315,N_11935,N_12304);
and U14316 (N_14316,N_10795,N_8223);
nor U14317 (N_14317,N_11362,N_10689);
and U14318 (N_14318,N_7848,N_12055);
and U14319 (N_14319,N_9204,N_10283);
xnor U14320 (N_14320,N_11435,N_8089);
and U14321 (N_14321,N_10347,N_10950);
or U14322 (N_14322,N_11492,N_10247);
and U14323 (N_14323,N_11632,N_7760);
or U14324 (N_14324,N_10717,N_9396);
nand U14325 (N_14325,N_7490,N_6956);
xor U14326 (N_14326,N_7234,N_11311);
nor U14327 (N_14327,N_7051,N_7964);
or U14328 (N_14328,N_7523,N_8556);
xnor U14329 (N_14329,N_12394,N_12247);
xor U14330 (N_14330,N_7370,N_6373);
nand U14331 (N_14331,N_11227,N_12408);
xnor U14332 (N_14332,N_11756,N_8327);
and U14333 (N_14333,N_10776,N_6901);
or U14334 (N_14334,N_9763,N_10494);
and U14335 (N_14335,N_7828,N_11737);
nor U14336 (N_14336,N_6767,N_11399);
and U14337 (N_14337,N_9159,N_8510);
and U14338 (N_14338,N_6570,N_11773);
nor U14339 (N_14339,N_9889,N_7016);
or U14340 (N_14340,N_9374,N_11450);
or U14341 (N_14341,N_7441,N_8499);
and U14342 (N_14342,N_10616,N_9755);
and U14343 (N_14343,N_11870,N_9323);
xnor U14344 (N_14344,N_10028,N_9017);
nor U14345 (N_14345,N_8021,N_9483);
and U14346 (N_14346,N_10894,N_7400);
and U14347 (N_14347,N_11692,N_11664);
and U14348 (N_14348,N_11005,N_10251);
nand U14349 (N_14349,N_10174,N_11459);
nand U14350 (N_14350,N_7262,N_11860);
nand U14351 (N_14351,N_11481,N_12449);
and U14352 (N_14352,N_8337,N_10810);
or U14353 (N_14353,N_8247,N_6917);
and U14354 (N_14354,N_12135,N_8727);
and U14355 (N_14355,N_7522,N_10775);
nor U14356 (N_14356,N_6527,N_11458);
and U14357 (N_14357,N_8136,N_11286);
and U14358 (N_14358,N_11943,N_12299);
or U14359 (N_14359,N_8792,N_8703);
nand U14360 (N_14360,N_10148,N_9506);
nand U14361 (N_14361,N_10077,N_8294);
or U14362 (N_14362,N_10292,N_9209);
nor U14363 (N_14363,N_7880,N_8615);
or U14364 (N_14364,N_12368,N_12018);
and U14365 (N_14365,N_6405,N_8047);
or U14366 (N_14366,N_11671,N_8082);
or U14367 (N_14367,N_10486,N_11546);
and U14368 (N_14368,N_12093,N_9343);
xnor U14369 (N_14369,N_7765,N_11329);
nor U14370 (N_14370,N_11401,N_12479);
xor U14371 (N_14371,N_7708,N_11209);
nor U14372 (N_14372,N_7622,N_11856);
and U14373 (N_14373,N_12155,N_6968);
or U14374 (N_14374,N_9800,N_12290);
nand U14375 (N_14375,N_10013,N_7219);
or U14376 (N_14376,N_8811,N_7049);
xnor U14377 (N_14377,N_11201,N_6264);
and U14378 (N_14378,N_10501,N_9974);
and U14379 (N_14379,N_7563,N_9675);
nand U14380 (N_14380,N_7726,N_11305);
nand U14381 (N_14381,N_10793,N_10733);
or U14382 (N_14382,N_11628,N_6606);
and U14383 (N_14383,N_11506,N_7047);
and U14384 (N_14384,N_6432,N_12265);
xor U14385 (N_14385,N_7403,N_9073);
and U14386 (N_14386,N_10630,N_9421);
nand U14387 (N_14387,N_7232,N_10060);
nor U14388 (N_14388,N_8739,N_9702);
nor U14389 (N_14389,N_8138,N_8909);
nand U14390 (N_14390,N_8240,N_8379);
nor U14391 (N_14391,N_7713,N_7246);
and U14392 (N_14392,N_11021,N_8324);
or U14393 (N_14393,N_10942,N_11453);
xor U14394 (N_14394,N_6905,N_11058);
and U14395 (N_14395,N_11513,N_10923);
and U14396 (N_14396,N_7467,N_6943);
nor U14397 (N_14397,N_8682,N_8747);
xor U14398 (N_14398,N_7796,N_11498);
or U14399 (N_14399,N_12125,N_10206);
nor U14400 (N_14400,N_9761,N_12154);
nor U14401 (N_14401,N_11894,N_10276);
and U14402 (N_14402,N_8940,N_8270);
nand U14403 (N_14403,N_10767,N_8105);
or U14404 (N_14404,N_9786,N_10869);
nor U14405 (N_14405,N_10439,N_12492);
xor U14406 (N_14406,N_11883,N_6796);
xnor U14407 (N_14407,N_12414,N_7864);
xor U14408 (N_14408,N_9466,N_11669);
nor U14409 (N_14409,N_6599,N_11718);
nand U14410 (N_14410,N_7682,N_9353);
xnor U14411 (N_14411,N_8525,N_8107);
nor U14412 (N_14412,N_8633,N_8851);
and U14413 (N_14413,N_8362,N_7680);
nor U14414 (N_14414,N_11462,N_9068);
xor U14415 (N_14415,N_7354,N_9780);
nand U14416 (N_14416,N_6569,N_8451);
nand U14417 (N_14417,N_7625,N_9922);
nor U14418 (N_14418,N_9990,N_9304);
or U14419 (N_14419,N_7458,N_7596);
and U14420 (N_14420,N_10199,N_7426);
xor U14421 (N_14421,N_9473,N_9048);
nand U14422 (N_14422,N_10559,N_7896);
nand U14423 (N_14423,N_11637,N_6424);
nor U14424 (N_14424,N_7853,N_9920);
nand U14425 (N_14425,N_10921,N_8124);
nor U14426 (N_14426,N_6374,N_7968);
and U14427 (N_14427,N_11962,N_6735);
or U14428 (N_14428,N_9602,N_7243);
nand U14429 (N_14429,N_7086,N_9644);
nor U14430 (N_14430,N_9333,N_7983);
nor U14431 (N_14431,N_11309,N_7581);
and U14432 (N_14432,N_11165,N_10609);
and U14433 (N_14433,N_7227,N_11160);
nand U14434 (N_14434,N_7819,N_9144);
nand U14435 (N_14435,N_10031,N_9171);
or U14436 (N_14436,N_9238,N_8381);
xnor U14437 (N_14437,N_11846,N_7535);
nor U14438 (N_14438,N_6379,N_9850);
nor U14439 (N_14439,N_8157,N_10483);
nand U14440 (N_14440,N_7739,N_7106);
xor U14441 (N_14441,N_6662,N_12298);
nor U14442 (N_14442,N_8275,N_6673);
and U14443 (N_14443,N_9967,N_10612);
nor U14444 (N_14444,N_9565,N_11093);
or U14445 (N_14445,N_7095,N_12065);
nor U14446 (N_14446,N_10464,N_10360);
or U14447 (N_14447,N_9738,N_12064);
nor U14448 (N_14448,N_8975,N_6737);
or U14449 (N_14449,N_11959,N_11016);
or U14450 (N_14450,N_7604,N_6282);
or U14451 (N_14451,N_11972,N_8369);
nor U14452 (N_14452,N_12497,N_7371);
and U14453 (N_14453,N_9232,N_11955);
xor U14454 (N_14454,N_6887,N_7630);
xor U14455 (N_14455,N_10402,N_10964);
nor U14456 (N_14456,N_8702,N_11893);
or U14457 (N_14457,N_10665,N_11683);
xor U14458 (N_14458,N_11724,N_8457);
nand U14459 (N_14459,N_11117,N_11099);
and U14460 (N_14460,N_11205,N_11446);
and U14461 (N_14461,N_7462,N_8501);
nor U14462 (N_14462,N_9054,N_10282);
nand U14463 (N_14463,N_12023,N_6497);
nor U14464 (N_14464,N_7759,N_7768);
and U14465 (N_14465,N_8256,N_11073);
and U14466 (N_14466,N_9368,N_6713);
nand U14467 (N_14467,N_8303,N_9696);
or U14468 (N_14468,N_7574,N_7631);
nand U14469 (N_14469,N_8763,N_7155);
nand U14470 (N_14470,N_7003,N_8513);
or U14471 (N_14471,N_11326,N_11444);
nand U14472 (N_14472,N_10918,N_9011);
nor U14473 (N_14473,N_7657,N_11713);
and U14474 (N_14474,N_6732,N_6938);
and U14475 (N_14475,N_8347,N_9463);
xnor U14476 (N_14476,N_10774,N_7525);
or U14477 (N_14477,N_10098,N_8852);
nor U14478 (N_14478,N_7242,N_9434);
and U14479 (N_14479,N_8081,N_9579);
nor U14480 (N_14480,N_7220,N_6954);
nor U14481 (N_14481,N_7586,N_9758);
or U14482 (N_14482,N_9556,N_11338);
nand U14483 (N_14483,N_11997,N_11553);
and U14484 (N_14484,N_6333,N_11330);
xnor U14485 (N_14485,N_11640,N_8032);
and U14486 (N_14486,N_8887,N_9554);
nand U14487 (N_14487,N_11633,N_7146);
nand U14488 (N_14488,N_8679,N_11864);
xor U14489 (N_14489,N_10988,N_8912);
and U14490 (N_14490,N_7872,N_10356);
nand U14491 (N_14491,N_10853,N_6835);
nand U14492 (N_14492,N_12454,N_7349);
xnor U14493 (N_14493,N_10638,N_9544);
or U14494 (N_14494,N_11505,N_6779);
nor U14495 (N_14495,N_6704,N_12096);
nand U14496 (N_14496,N_11156,N_10583);
or U14497 (N_14497,N_12389,N_10306);
or U14498 (N_14498,N_11038,N_10581);
or U14499 (N_14499,N_8395,N_9703);
nand U14500 (N_14500,N_7627,N_7496);
xnor U14501 (N_14501,N_11606,N_10266);
or U14502 (N_14502,N_10969,N_7506);
or U14503 (N_14503,N_10358,N_12498);
nand U14504 (N_14504,N_10007,N_9832);
nand U14505 (N_14505,N_11203,N_11555);
and U14506 (N_14506,N_6850,N_9235);
xor U14507 (N_14507,N_9874,N_10819);
nand U14508 (N_14508,N_9183,N_12474);
or U14509 (N_14509,N_6406,N_6339);
or U14510 (N_14510,N_6260,N_9769);
and U14511 (N_14511,N_7685,N_9654);
nand U14512 (N_14512,N_11501,N_7989);
or U14513 (N_14513,N_10861,N_7436);
nor U14514 (N_14514,N_9600,N_10130);
nor U14515 (N_14515,N_8522,N_7747);
or U14516 (N_14516,N_12223,N_9336);
nor U14517 (N_14517,N_10428,N_7591);
nand U14518 (N_14518,N_7814,N_6775);
xor U14519 (N_14519,N_8868,N_11308);
and U14520 (N_14520,N_6513,N_10264);
nor U14521 (N_14521,N_6632,N_12491);
xnor U14522 (N_14522,N_7692,N_11239);
and U14523 (N_14523,N_7392,N_10640);
and U14524 (N_14524,N_9137,N_9321);
nand U14525 (N_14525,N_11445,N_6756);
or U14526 (N_14526,N_9002,N_9971);
and U14527 (N_14527,N_12202,N_11953);
or U14528 (N_14528,N_7752,N_9904);
nand U14529 (N_14529,N_8930,N_7722);
xnor U14530 (N_14530,N_9219,N_11069);
nand U14531 (N_14531,N_7134,N_8014);
nand U14532 (N_14532,N_9268,N_11347);
and U14533 (N_14533,N_10331,N_12028);
or U14534 (N_14534,N_8407,N_6838);
or U14535 (N_14535,N_11994,N_6642);
nor U14536 (N_14536,N_9536,N_10835);
or U14537 (N_14537,N_7640,N_10570);
nand U14538 (N_14538,N_8297,N_6874);
and U14539 (N_14539,N_11457,N_7352);
nor U14540 (N_14540,N_7081,N_9202);
nor U14541 (N_14541,N_8734,N_9960);
and U14542 (N_14542,N_10414,N_9261);
and U14543 (N_14543,N_12332,N_8278);
or U14544 (N_14544,N_6579,N_11019);
nor U14545 (N_14545,N_8248,N_9706);
nor U14546 (N_14546,N_11060,N_9309);
and U14547 (N_14547,N_11300,N_10907);
and U14548 (N_14548,N_11298,N_7121);
nor U14549 (N_14549,N_8796,N_6335);
nand U14550 (N_14550,N_7550,N_6660);
or U14551 (N_14551,N_12150,N_10241);
nand U14552 (N_14552,N_8856,N_6646);
and U14553 (N_14553,N_6853,N_6832);
xor U14554 (N_14554,N_7863,N_12117);
and U14555 (N_14555,N_8773,N_7418);
nand U14556 (N_14556,N_6625,N_10859);
nor U14557 (N_14557,N_11925,N_11758);
nand U14558 (N_14558,N_10827,N_12484);
nor U14559 (N_14559,N_9088,N_9790);
xor U14560 (N_14560,N_12294,N_10066);
or U14561 (N_14561,N_10141,N_12446);
or U14562 (N_14562,N_12147,N_11302);
nor U14563 (N_14563,N_10746,N_9956);
or U14564 (N_14564,N_12035,N_10605);
nor U14565 (N_14565,N_8871,N_10741);
or U14566 (N_14566,N_10569,N_10925);
or U14567 (N_14567,N_6299,N_8375);
nor U14568 (N_14568,N_10708,N_11147);
and U14569 (N_14569,N_6930,N_8983);
xor U14570 (N_14570,N_6487,N_9196);
nand U14571 (N_14571,N_10737,N_9704);
or U14572 (N_14572,N_9871,N_8714);
nor U14573 (N_14573,N_10916,N_9906);
and U14574 (N_14574,N_7650,N_11919);
and U14575 (N_14575,N_10463,N_8565);
or U14576 (N_14576,N_10973,N_8927);
xor U14577 (N_14577,N_9734,N_8608);
or U14578 (N_14578,N_12126,N_11966);
and U14579 (N_14579,N_10608,N_8271);
or U14580 (N_14580,N_8452,N_7956);
nand U14581 (N_14581,N_12369,N_11079);
or U14582 (N_14582,N_9631,N_8122);
nand U14583 (N_14583,N_10858,N_7806);
or U14584 (N_14584,N_6778,N_10029);
and U14585 (N_14585,N_7190,N_7124);
nand U14586 (N_14586,N_8332,N_11225);
and U14587 (N_14587,N_10462,N_7861);
or U14588 (N_14588,N_6872,N_9682);
nor U14589 (N_14589,N_7209,N_7029);
nor U14590 (N_14590,N_6995,N_11140);
nand U14591 (N_14591,N_8694,N_8860);
and U14592 (N_14592,N_11845,N_6798);
nor U14593 (N_14593,N_8761,N_6710);
nand U14594 (N_14594,N_11630,N_10937);
nand U14595 (N_14595,N_7874,N_10167);
nor U14596 (N_14596,N_9664,N_10477);
nor U14597 (N_14597,N_7823,N_10497);
xor U14598 (N_14598,N_6408,N_9921);
nand U14599 (N_14599,N_10848,N_6960);
nand U14600 (N_14600,N_11162,N_8096);
nor U14601 (N_14601,N_6752,N_10589);
and U14602 (N_14602,N_9394,N_7266);
nor U14603 (N_14603,N_12222,N_6984);
and U14604 (N_14604,N_6847,N_10268);
nand U14605 (N_14605,N_8232,N_10744);
and U14606 (N_14606,N_9671,N_6466);
or U14607 (N_14607,N_12308,N_11623);
nand U14608 (N_14608,N_9742,N_6883);
and U14609 (N_14609,N_8196,N_12106);
xnor U14610 (N_14610,N_10161,N_9486);
and U14611 (N_14611,N_10203,N_11852);
and U14612 (N_14612,N_11672,N_6602);
or U14613 (N_14613,N_6590,N_7774);
and U14614 (N_14614,N_7833,N_10529);
or U14615 (N_14615,N_6334,N_7284);
nor U14616 (N_14616,N_9051,N_10545);
nor U14617 (N_14617,N_6266,N_10931);
nand U14618 (N_14618,N_12363,N_11158);
nor U14619 (N_14619,N_10219,N_8094);
nor U14620 (N_14620,N_6751,N_9022);
and U14621 (N_14621,N_10278,N_9923);
nor U14622 (N_14622,N_6390,N_7614);
xor U14623 (N_14623,N_6677,N_9571);
nand U14624 (N_14624,N_10340,N_9743);
nor U14625 (N_14625,N_6861,N_7965);
nor U14626 (N_14626,N_7325,N_9566);
or U14627 (N_14627,N_8059,N_9616);
or U14628 (N_14628,N_6556,N_12303);
or U14629 (N_14629,N_9371,N_10255);
xnor U14630 (N_14630,N_12320,N_6325);
xnor U14631 (N_14631,N_6980,N_9145);
and U14632 (N_14632,N_6292,N_7199);
nor U14633 (N_14633,N_10750,N_9034);
nor U14634 (N_14634,N_7200,N_10611);
and U14635 (N_14635,N_11535,N_9591);
and U14636 (N_14636,N_10461,N_9559);
nor U14637 (N_14637,N_7147,N_11297);
or U14638 (N_14638,N_6377,N_10102);
or U14639 (N_14639,N_9558,N_6305);
and U14640 (N_14640,N_9701,N_6387);
nand U14641 (N_14641,N_6797,N_7969);
nand U14642 (N_14642,N_6884,N_9957);
or U14643 (N_14643,N_10799,N_8961);
xnor U14644 (N_14644,N_6342,N_6647);
or U14645 (N_14645,N_11624,N_9529);
and U14646 (N_14646,N_9005,N_11805);
or U14647 (N_14647,N_7829,N_10008);
and U14648 (N_14648,N_10568,N_10751);
and U14649 (N_14649,N_10180,N_10806);
nor U14650 (N_14650,N_7476,N_8164);
nor U14651 (N_14651,N_8706,N_10188);
nor U14652 (N_14652,N_9319,N_10567);
xor U14653 (N_14653,N_8568,N_8311);
nor U14654 (N_14654,N_10177,N_8012);
and U14655 (N_14655,N_10971,N_7172);
or U14656 (N_14656,N_8221,N_11313);
nand U14657 (N_14657,N_11136,N_12037);
nor U14658 (N_14658,N_11708,N_8647);
and U14659 (N_14659,N_8896,N_9334);
and U14660 (N_14660,N_7615,N_10929);
nand U14661 (N_14661,N_8217,N_9090);
nand U14662 (N_14662,N_7820,N_6576);
nor U14663 (N_14663,N_10792,N_11987);
xnor U14664 (N_14664,N_7688,N_11390);
and U14665 (N_14665,N_9049,N_7425);
or U14666 (N_14666,N_9178,N_9615);
xnor U14667 (N_14667,N_8040,N_9479);
and U14668 (N_14668,N_11378,N_11413);
nand U14669 (N_14669,N_11707,N_8083);
or U14670 (N_14670,N_10557,N_7886);
nand U14671 (N_14671,N_11616,N_12057);
xnor U14672 (N_14672,N_11753,N_10791);
and U14673 (N_14673,N_11391,N_8291);
nand U14674 (N_14674,N_6653,N_8397);
nand U14675 (N_14675,N_7703,N_12379);
or U14676 (N_14676,N_11569,N_10027);
or U14677 (N_14677,N_10096,N_9538);
or U14678 (N_14678,N_9815,N_12489);
nor U14679 (N_14679,N_11631,N_6530);
or U14680 (N_14680,N_11256,N_6268);
xnor U14681 (N_14681,N_6862,N_12365);
nor U14682 (N_14682,N_10878,N_8384);
nand U14683 (N_14683,N_10724,N_10989);
and U14684 (N_14684,N_12485,N_10945);
or U14685 (N_14685,N_8989,N_12441);
or U14686 (N_14686,N_9339,N_12458);
nor U14687 (N_14687,N_6347,N_9505);
or U14688 (N_14688,N_6257,N_6376);
nor U14689 (N_14689,N_7875,N_10693);
and U14690 (N_14690,N_6665,N_7854);
and U14691 (N_14691,N_10063,N_8472);
or U14692 (N_14692,N_9075,N_12445);
nor U14693 (N_14693,N_11735,N_8923);
or U14694 (N_14694,N_7517,N_8078);
nor U14695 (N_14695,N_9959,N_7906);
and U14696 (N_14696,N_11488,N_6859);
and U14697 (N_14697,N_8963,N_8711);
or U14698 (N_14698,N_8052,N_8704);
nand U14699 (N_14699,N_7437,N_11258);
or U14700 (N_14700,N_7986,N_12163);
and U14701 (N_14701,N_8545,N_7336);
nor U14702 (N_14702,N_11438,N_12218);
or U14703 (N_14703,N_10588,N_12438);
and U14704 (N_14704,N_8652,N_9390);
and U14705 (N_14705,N_7185,N_11677);
and U14706 (N_14706,N_9041,N_7651);
or U14707 (N_14707,N_8874,N_9172);
or U14708 (N_14708,N_11402,N_9779);
or U14709 (N_14709,N_12240,N_9169);
nor U14710 (N_14710,N_11742,N_9907);
and U14711 (N_14711,N_9249,N_6875);
or U14712 (N_14712,N_7790,N_7188);
and U14713 (N_14713,N_9504,N_6944);
nand U14714 (N_14714,N_11597,N_10765);
or U14715 (N_14715,N_11518,N_10955);
or U14716 (N_14716,N_9552,N_7007);
or U14717 (N_14717,N_6833,N_10178);
and U14718 (N_14718,N_6327,N_7645);
or U14719 (N_14719,N_9119,N_11250);
nand U14720 (N_14720,N_10393,N_11342);
nor U14721 (N_14721,N_8790,N_9127);
nor U14722 (N_14722,N_6420,N_6892);
or U14723 (N_14723,N_8775,N_10179);
and U14724 (N_14724,N_8576,N_7546);
and U14725 (N_14725,N_7599,N_12346);
nor U14726 (N_14726,N_12315,N_6649);
or U14727 (N_14727,N_6946,N_12472);
nor U14728 (N_14728,N_6925,N_12210);
and U14729 (N_14729,N_8620,N_12115);
or U14730 (N_14730,N_8736,N_10088);
nor U14731 (N_14731,N_8516,N_11655);
nor U14732 (N_14732,N_7849,N_6629);
nor U14733 (N_14733,N_11000,N_11509);
nand U14734 (N_14734,N_9722,N_10163);
nand U14735 (N_14735,N_6601,N_6298);
nand U14736 (N_14736,N_11071,N_9936);
and U14737 (N_14737,N_10519,N_8154);
or U14738 (N_14738,N_12116,N_10909);
or U14739 (N_14739,N_8533,N_12258);
or U14740 (N_14740,N_6840,N_9071);
nand U14741 (N_14741,N_11748,N_6744);
nor U14742 (N_14742,N_8603,N_8539);
nor U14743 (N_14743,N_8934,N_6529);
nor U14744 (N_14744,N_11907,N_10205);
or U14745 (N_14745,N_6436,N_8187);
nor U14746 (N_14746,N_7017,N_9084);
and U14747 (N_14747,N_11858,N_8782);
or U14748 (N_14748,N_9513,N_9037);
nor U14749 (N_14749,N_12417,N_10873);
and U14750 (N_14750,N_10003,N_11436);
and U14751 (N_14751,N_8104,N_11310);
nand U14752 (N_14752,N_11455,N_10030);
xnor U14753 (N_14753,N_9236,N_9502);
and U14754 (N_14754,N_9430,N_10194);
or U14755 (N_14755,N_8745,N_10092);
nand U14756 (N_14756,N_10798,N_8638);
or U14757 (N_14757,N_6618,N_10758);
xnor U14758 (N_14758,N_9457,N_7184);
nand U14759 (N_14759,N_9340,N_9716);
and U14760 (N_14760,N_8667,N_10782);
nor U14761 (N_14761,N_11120,N_10814);
nand U14762 (N_14762,N_12331,N_8742);
xnor U14763 (N_14763,N_8629,N_11651);
and U14764 (N_14764,N_12376,N_11557);
nand U14765 (N_14765,N_9288,N_6667);
nand U14766 (N_14766,N_7011,N_12071);
or U14767 (N_14767,N_7740,N_12439);
nor U14768 (N_14768,N_6644,N_11607);
or U14769 (N_14769,N_11369,N_11456);
or U14770 (N_14770,N_11235,N_7080);
or U14771 (N_14771,N_7997,N_9924);
or U14772 (N_14772,N_7588,N_8972);
and U14773 (N_14773,N_7432,N_8543);
xnor U14774 (N_14774,N_7724,N_9930);
xor U14775 (N_14775,N_6288,N_9912);
nand U14776 (N_14776,N_9158,N_7935);
and U14777 (N_14777,N_7862,N_8586);
and U14778 (N_14778,N_12433,N_11905);
nor U14779 (N_14779,N_11427,N_8486);
nand U14780 (N_14780,N_8287,N_12334);
nand U14781 (N_14781,N_6561,N_7676);
or U14782 (N_14782,N_8415,N_9875);
or U14783 (N_14783,N_8368,N_11679);
nor U14784 (N_14784,N_10899,N_6858);
or U14785 (N_14785,N_9757,N_9986);
and U14786 (N_14786,N_8025,N_11891);
or U14787 (N_14787,N_6265,N_7139);
xnor U14788 (N_14788,N_8115,N_8280);
nand U14789 (N_14789,N_11118,N_9213);
xor U14790 (N_14790,N_6566,N_11969);
nand U14791 (N_14791,N_11045,N_8440);
and U14792 (N_14792,N_7116,N_9447);
nand U14793 (N_14793,N_9806,N_9125);
nand U14794 (N_14794,N_8602,N_8564);
or U14795 (N_14795,N_11198,N_8886);
or U14796 (N_14796,N_10747,N_9872);
and U14797 (N_14797,N_12425,N_11056);
nor U14798 (N_14798,N_8230,N_10975);
nor U14799 (N_14799,N_9266,N_9837);
nor U14800 (N_14800,N_7469,N_6719);
nor U14801 (N_14801,N_12179,N_6337);
nor U14802 (N_14802,N_11732,N_7419);
nor U14803 (N_14803,N_9379,N_7353);
and U14804 (N_14804,N_11808,N_12423);
nor U14805 (N_14805,N_9698,N_8442);
nor U14806 (N_14806,N_9134,N_8555);
nand U14807 (N_14807,N_11991,N_7423);
and U14808 (N_14808,N_7363,N_11189);
nand U14809 (N_14809,N_7118,N_6577);
or U14810 (N_14810,N_6486,N_9794);
or U14811 (N_14811,N_8511,N_8999);
and U14812 (N_14812,N_11752,N_12044);
nand U14813 (N_14813,N_8803,N_9317);
or U14814 (N_14814,N_11159,N_11855);
and U14815 (N_14815,N_11576,N_10396);
and U14816 (N_14816,N_9342,N_7940);
and U14817 (N_14817,N_12053,N_8944);
nand U14818 (N_14818,N_9412,N_10342);
and U14819 (N_14819,N_9918,N_9311);
nor U14820 (N_14820,N_7067,N_10415);
nor U14821 (N_14821,N_9248,N_9952);
and U14822 (N_14822,N_7487,N_6302);
xor U14823 (N_14823,N_10924,N_10966);
or U14824 (N_14824,N_8199,N_12442);
nand U14825 (N_14825,N_10636,N_6736);
and U14826 (N_14826,N_11499,N_12243);
nor U14827 (N_14827,N_11480,N_12385);
nand U14828 (N_14828,N_8134,N_7783);
xor U14829 (N_14829,N_10633,N_11605);
or U14830 (N_14830,N_7866,N_7731);
nand U14831 (N_14831,N_10220,N_11785);
and U14832 (N_14832,N_6927,N_6900);
nand U14833 (N_14833,N_11145,N_10573);
and U14834 (N_14834,N_8140,N_11200);
nand U14835 (N_14835,N_7811,N_9678);
or U14836 (N_14836,N_12189,N_11432);
and U14837 (N_14837,N_9441,N_12014);
or U14838 (N_14838,N_11244,N_11166);
or U14839 (N_14839,N_12129,N_8197);
xnor U14840 (N_14840,N_8290,N_8062);
nand U14841 (N_14841,N_11066,N_9935);
and U14842 (N_14842,N_11762,N_7177);
or U14843 (N_14843,N_11574,N_10321);
and U14844 (N_14844,N_9550,N_11590);
and U14845 (N_14845,N_7143,N_6596);
nor U14846 (N_14846,N_9356,N_6757);
nor U14847 (N_14847,N_9200,N_9903);
and U14848 (N_14848,N_11351,N_7495);
nand U14849 (N_14849,N_11667,N_6945);
nor U14850 (N_14850,N_6348,N_7572);
and U14851 (N_14851,N_10061,N_7914);
nand U14852 (N_14852,N_9911,N_8613);
or U14853 (N_14853,N_6786,N_8809);
and U14854 (N_14854,N_8784,N_8597);
or U14855 (N_14855,N_7004,N_6966);
or U14856 (N_14856,N_7501,N_6991);
and U14857 (N_14857,N_7919,N_9820);
or U14858 (N_14858,N_9365,N_9778);
or U14859 (N_14859,N_7028,N_10058);
and U14860 (N_14860,N_6935,N_7728);
xor U14861 (N_14861,N_9497,N_11367);
nand U14862 (N_14862,N_6888,N_9489);
or U14863 (N_14863,N_10905,N_11570);
or U14864 (N_14864,N_7539,N_10057);
and U14865 (N_14865,N_11385,N_9113);
and U14866 (N_14866,N_9407,N_8441);
nand U14867 (N_14867,N_9111,N_9724);
or U14868 (N_14868,N_10882,N_11318);
nor U14869 (N_14869,N_7761,N_9525);
and U14870 (N_14870,N_8783,N_11830);
nor U14871 (N_14871,N_9095,N_11993);
nand U14872 (N_14872,N_6911,N_11879);
nand U14873 (N_14873,N_11917,N_11430);
nor U14874 (N_14874,N_10705,N_10453);
or U14875 (N_14875,N_6478,N_6557);
and U14876 (N_14876,N_12341,N_12371);
and U14877 (N_14877,N_9534,N_9207);
nand U14878 (N_14878,N_10055,N_11467);
and U14879 (N_14879,N_7302,N_11422);
and U14880 (N_14880,N_6345,N_11595);
and U14881 (N_14881,N_6274,N_6816);
and U14882 (N_14882,N_11204,N_7282);
and U14883 (N_14883,N_8996,N_10518);
or U14884 (N_14884,N_8913,N_8305);
nor U14885 (N_14885,N_12195,N_6543);
nand U14886 (N_14886,N_9197,N_9176);
and U14887 (N_14887,N_7273,N_8580);
and U14888 (N_14888,N_12019,N_10690);
nor U14889 (N_14889,N_8992,N_7619);
and U14890 (N_14890,N_10700,N_8998);
and U14891 (N_14891,N_6455,N_8875);
nand U14892 (N_14892,N_6361,N_8210);
nor U14893 (N_14893,N_8658,N_8394);
xnor U14894 (N_14894,N_8370,N_8732);
nor U14895 (N_14895,N_7466,N_8878);
nor U14896 (N_14896,N_7460,N_7900);
nand U14897 (N_14897,N_12219,N_8798);
or U14898 (N_14898,N_12302,N_9719);
and U14899 (N_14899,N_6452,N_10657);
nor U14900 (N_14900,N_10556,N_10533);
xor U14901 (N_14901,N_12157,N_12293);
nor U14902 (N_14902,N_8143,N_12133);
nand U14903 (N_14903,N_6648,N_11008);
and U14904 (N_14904,N_6828,N_6889);
and U14905 (N_14905,N_9672,N_7707);
nor U14906 (N_14906,N_11989,N_9847);
or U14907 (N_14907,N_6789,N_6304);
nor U14908 (N_14908,N_7966,N_9377);
or U14909 (N_14909,N_8022,N_10622);
nor U14910 (N_14910,N_12173,N_8600);
or U14911 (N_14911,N_11974,N_9645);
nor U14912 (N_14912,N_9528,N_12073);
and U14913 (N_14913,N_7894,N_7270);
or U14914 (N_14914,N_7473,N_7069);
nand U14915 (N_14915,N_8257,N_11988);
nor U14916 (N_14916,N_6520,N_6680);
and U14917 (N_14917,N_6784,N_11364);
or U14918 (N_14918,N_7387,N_10625);
nand U14919 (N_14919,N_6540,N_11738);
and U14920 (N_14920,N_8847,N_9883);
or U14921 (N_14921,N_10770,N_7598);
nand U14922 (N_14922,N_12206,N_8323);
or U14923 (N_14923,N_12361,N_12185);
and U14924 (N_14924,N_8120,N_11587);
or U14925 (N_14925,N_10229,N_9574);
and U14926 (N_14926,N_8431,N_11031);
xnor U14927 (N_14927,N_9711,N_7792);
or U14928 (N_14928,N_10772,N_9691);
nand U14929 (N_14929,N_8195,N_8299);
and U14930 (N_14930,N_11051,N_10113);
xnor U14931 (N_14931,N_7505,N_10960);
and U14932 (N_14932,N_12255,N_10812);
xor U14933 (N_14933,N_9362,N_8228);
nand U14934 (N_14934,N_12032,N_12257);
or U14935 (N_14935,N_7152,N_8259);
xnor U14936 (N_14936,N_9062,N_8201);
and U14937 (N_14937,N_10653,N_6776);
nand U14938 (N_14938,N_7857,N_9131);
and U14939 (N_14939,N_10585,N_7881);
or U14940 (N_14940,N_9093,N_7430);
nand U14941 (N_14941,N_6916,N_6439);
nor U14942 (N_14942,N_6986,N_9024);
nor U14943 (N_14943,N_11918,N_10984);
nand U14944 (N_14944,N_6717,N_11781);
or U14945 (N_14945,N_9517,N_10072);
or U14946 (N_14946,N_12224,N_7508);
nor U14947 (N_14947,N_8483,N_6849);
or U14948 (N_14948,N_11443,N_11687);
and U14949 (N_14949,N_12052,N_8869);
nand U14950 (N_14950,N_11133,N_12090);
nand U14951 (N_14951,N_6897,N_10572);
or U14952 (N_14952,N_11914,N_12355);
xnor U14953 (N_14953,N_12215,N_10528);
xnor U14954 (N_14954,N_8917,N_7479);
nand U14955 (N_14955,N_6380,N_8695);
and U14956 (N_14956,N_10208,N_8184);
nor U14957 (N_14957,N_10720,N_9372);
nand U14958 (N_14958,N_11331,N_10730);
nand U14959 (N_14959,N_8364,N_9122);
nor U14960 (N_14960,N_10115,N_11039);
or U14961 (N_14961,N_10911,N_9985);
and U14962 (N_14962,N_11479,N_10474);
or U14963 (N_14963,N_6918,N_10754);
nor U14964 (N_14964,N_11006,N_9231);
and U14965 (N_14965,N_11398,N_10357);
and U14966 (N_14966,N_6867,N_8497);
nand U14967 (N_14967,N_6297,N_10550);
xnor U14968 (N_14968,N_7773,N_6799);
nand U14969 (N_14969,N_7648,N_9485);
and U14970 (N_14970,N_7661,N_8449);
and U14971 (N_14971,N_11153,N_11819);
nor U14972 (N_14972,N_12388,N_7818);
nor U14973 (N_14973,N_6740,N_10471);
or U14974 (N_14974,N_11734,N_8333);
xnor U14975 (N_14975,N_9021,N_10823);
nand U14976 (N_14976,N_7891,N_11650);
nand U14977 (N_14977,N_9524,N_12061);
xnor U14978 (N_14978,N_7379,N_8108);
nand U14979 (N_14979,N_7583,N_10760);
and U14980 (N_14980,N_9693,N_12041);
and U14981 (N_14981,N_9237,N_11392);
nand U14982 (N_14982,N_12011,N_6635);
nand U14983 (N_14983,N_9375,N_10071);
nand U14984 (N_14984,N_10275,N_9655);
nor U14985 (N_14985,N_11875,N_10117);
and U14986 (N_14986,N_11465,N_11730);
or U14987 (N_14987,N_10516,N_11523);
nand U14988 (N_14988,N_6444,N_9818);
or U14989 (N_14989,N_12348,N_6511);
and U14990 (N_14990,N_8234,N_9795);
nor U14991 (N_14991,N_11238,N_10932);
or U14992 (N_14992,N_9491,N_10159);
and U14993 (N_14993,N_8476,N_10401);
or U14994 (N_14994,N_7711,N_9612);
nor U14995 (N_14995,N_11111,N_9541);
nand U14996 (N_14996,N_7686,N_7623);
nor U14997 (N_14997,N_8833,N_11510);
nor U14998 (N_14998,N_8186,N_12317);
nor U14999 (N_14999,N_9226,N_10970);
nand U15000 (N_15000,N_8233,N_7868);
nand U15001 (N_15001,N_9242,N_6661);
nand U15002 (N_15002,N_9089,N_11963);
xnor U15003 (N_15003,N_11130,N_10111);
and U15004 (N_15004,N_11484,N_9015);
and U15005 (N_15005,N_10871,N_11565);
or U15006 (N_15006,N_7167,N_8526);
nand U15007 (N_15007,N_6514,N_11887);
or U15008 (N_15008,N_12042,N_8180);
and U15009 (N_15009,N_8657,N_7396);
and U15010 (N_15010,N_11836,N_6413);
and U15011 (N_15011,N_8573,N_9294);
xor U15012 (N_15012,N_8056,N_10293);
or U15013 (N_15013,N_11828,N_12152);
or U15014 (N_15014,N_8053,N_7094);
xnor U15015 (N_15015,N_7516,N_8735);
nor U15016 (N_15016,N_9032,N_6273);
nand U15017 (N_15017,N_12409,N_7355);
or U15018 (N_15018,N_9203,N_9669);
and U15019 (N_15019,N_8743,N_11469);
xnor U15020 (N_15020,N_9078,N_12109);
nor U15021 (N_15021,N_10829,N_8744);
and U15022 (N_15022,N_8156,N_11992);
nor U15023 (N_15023,N_11382,N_7646);
nand U15024 (N_15024,N_8908,N_10839);
nor U15025 (N_15025,N_8071,N_10476);
and U15026 (N_15026,N_9369,N_11859);
nor U15027 (N_15027,N_11585,N_8882);
nor U15028 (N_15028,N_6620,N_9004);
nor U15029 (N_15029,N_9641,N_10841);
nor U15030 (N_15030,N_9043,N_6458);
nor U15031 (N_15031,N_9493,N_11017);
and U15032 (N_15032,N_8242,N_11129);
nand U15033 (N_15033,N_8288,N_11697);
or U15034 (N_15034,N_10227,N_10303);
nand U15035 (N_15035,N_7520,N_10824);
nand U15036 (N_15036,N_7085,N_11823);
and U15037 (N_15037,N_11696,N_11912);
nand U15038 (N_15038,N_10698,N_9861);
and U15039 (N_15039,N_11617,N_7076);
nand U15040 (N_15040,N_7088,N_12427);
nor U15041 (N_15041,N_7279,N_10927);
and U15042 (N_15042,N_7606,N_6693);
nand U15043 (N_15043,N_8458,N_12237);
nor U15044 (N_15044,N_11525,N_12047);
nand U15045 (N_15045,N_6446,N_10648);
nand U15046 (N_15046,N_8922,N_11572);
or U15047 (N_15047,N_9594,N_7194);
and U15048 (N_15048,N_11958,N_11151);
or U15049 (N_15049,N_7840,N_11645);
nor U15050 (N_15050,N_10398,N_7830);
and U15051 (N_15051,N_10883,N_7669);
nand U15052 (N_15052,N_8401,N_11067);
xor U15053 (N_15053,N_10145,N_11325);
and U15054 (N_15054,N_11999,N_6259);
nor U15055 (N_15055,N_10875,N_8054);
nor U15056 (N_15056,N_11044,N_9916);
or U15057 (N_15057,N_8281,N_8205);
and U15058 (N_15058,N_8097,N_11971);
nand U15059 (N_15059,N_7677,N_10509);
nor U15060 (N_15060,N_10598,N_11466);
or U15061 (N_15061,N_8066,N_8634);
or U15062 (N_15062,N_8873,N_6907);
or U15063 (N_15063,N_7743,N_10433);
nand U15064 (N_15064,N_12142,N_7762);
xnor U15065 (N_15065,N_9423,N_6700);
nand U15066 (N_15066,N_10958,N_10444);
xor U15067 (N_15067,N_6771,N_10949);
nor U15068 (N_15068,N_10069,N_7211);
nand U15069 (N_15069,N_10384,N_10458);
and U15070 (N_15070,N_11317,N_10977);
nand U15071 (N_15071,N_8067,N_6296);
nand U15072 (N_15072,N_7283,N_10201);
xnor U15073 (N_15073,N_12411,N_7105);
nor U15074 (N_15074,N_12422,N_9155);
xnor U15075 (N_15075,N_9979,N_12128);
nand U15076 (N_15076,N_6615,N_10400);
nand U15077 (N_15077,N_9817,N_9170);
nand U15078 (N_15078,N_8419,N_12330);
nor U15079 (N_15079,N_7304,N_9689);
nand U15080 (N_15080,N_8198,N_11419);
xor U15081 (N_15081,N_11143,N_11343);
nor U15082 (N_15082,N_7451,N_6697);
and U15083 (N_15083,N_7628,N_8942);
or U15084 (N_15084,N_9014,N_12495);
nand U15085 (N_15085,N_9746,N_8979);
or U15086 (N_15086,N_9908,N_10849);
xnor U15087 (N_15087,N_10707,N_6854);
or U15088 (N_15088,N_11368,N_8251);
or U15089 (N_15089,N_6827,N_10884);
nor U15090 (N_15090,N_10759,N_11936);
or U15091 (N_15091,N_11776,N_12307);
nor U15092 (N_15092,N_10731,N_8045);
or U15093 (N_15093,N_9753,N_11945);
xnor U15094 (N_15094,N_9831,N_7151);
xor U15095 (N_15095,N_9382,N_9862);
and U15096 (N_15096,N_12201,N_6597);
and U15097 (N_15097,N_9277,N_8546);
nor U15098 (N_15098,N_6402,N_7668);
and U15099 (N_15099,N_12271,N_6864);
nand U15100 (N_15100,N_9838,N_7678);
nor U15101 (N_15101,N_8284,N_12162);
and U15102 (N_15102,N_9687,N_6447);
nand U15103 (N_15103,N_11882,N_9224);
or U15104 (N_15104,N_9291,N_9077);
nor U15105 (N_15105,N_12054,N_7453);
or U15106 (N_15106,N_11054,N_11559);
nand U15107 (N_15107,N_12183,N_6820);
xnor U15108 (N_15108,N_10811,N_9681);
nand U15109 (N_15109,N_7274,N_10852);
nor U15110 (N_15110,N_7571,N_10352);
or U15111 (N_15111,N_11183,N_9975);
or U15112 (N_15112,N_6669,N_12203);
xor U15113 (N_15113,N_9303,N_11998);
and U15114 (N_15114,N_9803,N_6992);
nand U15115 (N_15115,N_7687,N_8789);
or U15116 (N_15116,N_8648,N_7753);
nor U15117 (N_15117,N_8937,N_11866);
nor U15118 (N_15118,N_9481,N_11090);
or U15119 (N_15119,N_10868,N_8444);
nand U15120 (N_15120,N_8158,N_8995);
nand U15121 (N_15121,N_8651,N_10371);
or U15122 (N_15122,N_9383,N_9030);
nor U15123 (N_15123,N_10922,N_9130);
and U15124 (N_15124,N_7013,N_11187);
or U15125 (N_15125,N_9707,N_8899);
nand U15126 (N_15126,N_7515,N_7721);
and U15127 (N_15127,N_7207,N_7062);
or U15128 (N_15128,N_6500,N_8102);
nand U15129 (N_15129,N_8160,N_10386);
nand U15130 (N_15130,N_8691,N_10445);
nand U15131 (N_15131,N_7042,N_7305);
and U15132 (N_15132,N_7734,N_9933);
nor U15133 (N_15133,N_9239,N_8002);
or U15134 (N_15134,N_6929,N_7470);
nand U15135 (N_15135,N_12193,N_7260);
nor U15136 (N_15136,N_6971,N_9292);
nand U15137 (N_15137,N_6449,N_7748);
nand U15138 (N_15138,N_10780,N_11042);
nor U15139 (N_15139,N_10230,N_9141);
and U15140 (N_15140,N_9495,N_11816);
nor U15141 (N_15141,N_9775,N_7716);
nor U15142 (N_15142,N_7745,N_6684);
or U15143 (N_15143,N_6280,N_6516);
xor U15144 (N_15144,N_8720,N_6256);
nand U15145 (N_15145,N_6985,N_7735);
and U15146 (N_15146,N_12015,N_7887);
nor U15147 (N_15147,N_7153,N_12347);
nor U15148 (N_15148,N_7904,N_9561);
nor U15149 (N_15149,N_10041,N_9557);
nor U15150 (N_15150,N_9098,N_10089);
or U15151 (N_15151,N_9260,N_11433);
nand U15152 (N_15152,N_10898,N_9472);
and U15153 (N_15153,N_7114,N_11909);
nor U15154 (N_15154,N_6360,N_7658);
or U15155 (N_15155,N_7344,N_10831);
nor U15156 (N_15156,N_10134,N_11757);
and U15157 (N_15157,N_10176,N_9109);
or U15158 (N_15158,N_6394,N_7895);
nand U15159 (N_15159,N_8741,N_11339);
and U15160 (N_15160,N_8863,N_12095);
and U15161 (N_15161,N_6720,N_6336);
or U15162 (N_15162,N_7634,N_9123);
xor U15163 (N_15163,N_10421,N_10522);
or U15164 (N_15164,N_10595,N_7052);
and U15165 (N_15165,N_10887,N_10539);
and U15166 (N_15166,N_7926,N_9713);
nor U15167 (N_15167,N_9312,N_7929);
or U15168 (N_15168,N_9674,N_9173);
nand U15169 (N_15169,N_11675,N_7216);
and U15170 (N_15170,N_11764,N_9658);
or U15171 (N_15171,N_12200,N_8579);
or U15172 (N_15172,N_10274,N_11901);
nor U15173 (N_15173,N_10576,N_6414);
nand U15174 (N_15174,N_10005,N_10999);
nand U15175 (N_15175,N_9947,N_8252);
nor U15176 (N_15176,N_7107,N_7000);
nor U15177 (N_15177,N_8895,N_12241);
and U15178 (N_15178,N_7568,N_10410);
nand U15179 (N_15179,N_8446,N_11777);
nor U15180 (N_15180,N_8017,N_10108);
nor U15181 (N_15181,N_11109,N_10768);
nand U15182 (N_15182,N_8116,N_10281);
and U15183 (N_15183,N_7039,N_8595);
and U15184 (N_15184,N_8818,N_12105);
or U15185 (N_15185,N_11913,N_8003);
xnor U15186 (N_15186,N_11072,N_10512);
nand U15187 (N_15187,N_8726,N_10745);
nor U15188 (N_15188,N_7222,N_9385);
xnor U15189 (N_15189,N_6829,N_10856);
nor U15190 (N_15190,N_6926,N_10150);
and U15191 (N_15191,N_8678,N_10766);
or U15192 (N_15192,N_12396,N_9440);
nor U15193 (N_15193,N_6922,N_9378);
nand U15194 (N_15194,N_12207,N_11266);
and U15195 (N_15195,N_6463,N_11028);
nor U15196 (N_15196,N_8301,N_8688);
or U15197 (N_15197,N_10143,N_8879);
xnor U15198 (N_15198,N_11892,N_11779);
xnor U15199 (N_15199,N_6303,N_9807);
or U15200 (N_15200,N_10149,N_6844);
or U15201 (N_15201,N_8590,N_10599);
or U15202 (N_15202,N_12112,N_11388);
nor U15203 (N_15203,N_8200,N_11741);
nor U15204 (N_15204,N_10271,N_11711);
or U15205 (N_15205,N_11299,N_8485);
and U15206 (N_15206,N_10594,N_10286);
nor U15207 (N_15207,N_11269,N_11949);
nand U15208 (N_15208,N_8924,N_6559);
nor U15209 (N_15209,N_12435,N_8574);
or U15210 (N_15210,N_9322,N_7319);
or U15211 (N_15211,N_9201,N_10503);
nor U15212 (N_15212,N_10997,N_6878);
nand U15213 (N_15213,N_9185,N_8906);
nor U15214 (N_15214,N_9683,N_8090);
xor U15215 (N_15215,N_9076,N_9404);
and U15216 (N_15216,N_10265,N_11685);
and U15217 (N_15217,N_6671,N_10070);
or U15218 (N_15218,N_11134,N_11442);
nor U15219 (N_15219,N_11765,N_7223);
or U15220 (N_15220,N_6621,N_11784);
or U15221 (N_15221,N_8631,N_6942);
nor U15222 (N_15222,N_8422,N_6567);
or U15223 (N_15223,N_7492,N_6367);
nor U15224 (N_15224,N_6612,N_9636);
or U15225 (N_15225,N_10540,N_7123);
or U15226 (N_15226,N_7465,N_9661);
nand U15227 (N_15227,N_10050,N_11366);
or U15228 (N_15228,N_10233,N_10049);
nand U15229 (N_15229,N_12132,N_11996);
xor U15230 (N_15230,N_7955,N_7318);
xnor U15231 (N_15231,N_6442,N_8202);
and U15232 (N_15232,N_10872,N_12476);
nor U15233 (N_15233,N_8453,N_9741);
or U15234 (N_15234,N_7842,N_7696);
or U15235 (N_15235,N_10656,N_10002);
nor U15236 (N_15236,N_11589,N_6558);
xnor U15237 (N_15237,N_10171,N_9720);
or U15238 (N_15238,N_6652,N_7037);
or U15239 (N_15239,N_6507,N_10610);
nor U15240 (N_15240,N_7901,N_9994);
or U15241 (N_15241,N_11554,N_10103);
and U15242 (N_15242,N_9110,N_7182);
nand U15243 (N_15243,N_7026,N_12475);
nor U15244 (N_15244,N_10026,N_11904);
nand U15245 (N_15245,N_7171,N_9428);
or U15246 (N_15246,N_12313,N_11744);
nand U15247 (N_15247,N_10182,N_8804);
nand U15248 (N_15248,N_8624,N_8315);
or U15249 (N_15249,N_6551,N_7503);
nor U15250 (N_15250,N_11537,N_12070);
nand U15251 (N_15251,N_10189,N_9623);
nor U15252 (N_15252,N_10324,N_9726);
and U15253 (N_15253,N_6788,N_8885);
nor U15254 (N_15254,N_11581,N_11582);
or U15255 (N_15255,N_11113,N_7312);
and U15256 (N_15256,N_10695,N_8640);
and U15257 (N_15257,N_11796,N_9349);
nor U15258 (N_15258,N_6448,N_7666);
and U15259 (N_15259,N_12161,N_7793);
and U15260 (N_15260,N_9287,N_9948);
xnor U15261 (N_15261,N_6608,N_8162);
nand U15262 (N_15262,N_8418,N_12380);
xor U15263 (N_15263,N_7072,N_7348);
nor U15264 (N_15264,N_12401,N_10888);
or U15265 (N_15265,N_6636,N_8377);
nand U15266 (N_15266,N_7193,N_8016);
nand U15267 (N_15267,N_8411,N_8076);
or U15268 (N_15268,N_10416,N_7987);
nor U15269 (N_15269,N_8006,N_6948);
nor U15270 (N_15270,N_6396,N_12370);
nand U15271 (N_15271,N_8465,N_10719);
and U15272 (N_15272,N_7240,N_8953);
nand U15273 (N_15273,N_6976,N_6560);
nand U15274 (N_15274,N_10934,N_11291);
nand U15275 (N_15275,N_11270,N_12272);
or U15276 (N_15276,N_6741,N_7738);
nand U15277 (N_15277,N_9152,N_7555);
and U15278 (N_15278,N_9050,N_9520);
nand U15279 (N_15279,N_10906,N_8121);
nor U15280 (N_15280,N_7196,N_6317);
or U15281 (N_15281,N_12434,N_6964);
or U15282 (N_15282,N_10372,N_7212);
or U15283 (N_15283,N_12459,N_8312);
or U15284 (N_15284,N_10590,N_10273);
nand U15285 (N_15285,N_9488,N_11921);
xor U15286 (N_15286,N_12264,N_6403);
xnor U15287 (N_15287,N_9972,N_7510);
and U15288 (N_15288,N_9686,N_12234);
or U15289 (N_15289,N_7063,N_7750);
or U15290 (N_15290,N_9628,N_9688);
nor U15291 (N_15291,N_8438,N_11861);
nand U15292 (N_15292,N_11414,N_8173);
nand U15293 (N_15293,N_11984,N_9961);
or U15294 (N_15294,N_10597,N_7635);
nor U15295 (N_15295,N_8644,N_6836);
and U15296 (N_15296,N_10836,N_8795);
or U15297 (N_15297,N_11411,N_11906);
or U15298 (N_15298,N_11829,N_11023);
or U15299 (N_15299,N_8883,N_11714);
xnor U15300 (N_15300,N_10042,N_7362);
nand U15301 (N_15301,N_9633,N_10904);
xor U15302 (N_15302,N_12426,N_8363);
nor U15303 (N_15303,N_7544,N_11691);
nand U15304 (N_15304,N_8881,N_10080);
and U15305 (N_15305,N_8536,N_7889);
xor U15306 (N_15306,N_12436,N_7534);
nand U15307 (N_15307,N_9243,N_11768);
nor U15308 (N_15308,N_9679,N_7624);
nand U15309 (N_15309,N_9003,N_7769);
or U15310 (N_15310,N_11626,N_11849);
nor U15311 (N_15311,N_8183,N_7091);
nand U15312 (N_15312,N_7797,N_9801);
nand U15313 (N_15313,N_6791,N_11221);
nor U15314 (N_15314,N_12131,N_8171);
and U15315 (N_15315,N_7670,N_6727);
nand U15316 (N_15316,N_12413,N_8142);
nand U15317 (N_15317,N_11333,N_10684);
xor U15318 (N_15318,N_6338,N_10995);
or U15319 (N_15319,N_11290,N_7998);
nor U15320 (N_15320,N_7119,N_10193);
nand U15321 (N_15321,N_10982,N_9570);
nand U15322 (N_15322,N_7602,N_7977);
nor U15323 (N_15323,N_11348,N_12094);
xnor U15324 (N_15324,N_6381,N_9198);
xnor U15325 (N_15325,N_11049,N_9937);
nand U15326 (N_15326,N_10862,N_7961);
nand U15327 (N_15327,N_9451,N_8487);
nand U15328 (N_15328,N_12100,N_9938);
xnor U15329 (N_15329,N_11373,N_10699);
and U15330 (N_15330,N_9884,N_10385);
xor U15331 (N_15331,N_6908,N_9338);
or U15332 (N_15332,N_6328,N_6729);
xnor U15333 (N_15333,N_11644,N_7377);
or U15334 (N_15334,N_6401,N_9499);
and U15335 (N_15335,N_10446,N_10739);
nor U15336 (N_15336,N_8024,N_12326);
nor U15337 (N_15337,N_11563,N_11224);
nor U15338 (N_15338,N_8689,N_11545);
and U15339 (N_15339,N_6372,N_10192);
or U15340 (N_15340,N_6749,N_6522);
or U15341 (N_15341,N_6610,N_8506);
nor U15342 (N_15342,N_12021,N_8131);
or U15343 (N_15343,N_7934,N_8326);
nor U15344 (N_15344,N_6846,N_10459);
and U15345 (N_15345,N_7675,N_7292);
nor U15346 (N_15346,N_9983,N_8504);
nor U15347 (N_15347,N_10213,N_6510);
and U15348 (N_15348,N_10864,N_9027);
or U15349 (N_15349,N_9614,N_9344);
and U15350 (N_15350,N_10418,N_10803);
xnor U15351 (N_15351,N_6411,N_8962);
nor U15352 (N_15352,N_8272,N_6562);
and U15353 (N_15353,N_9420,N_7159);
and U15354 (N_15354,N_11452,N_6866);
or U15355 (N_15355,N_9877,N_7946);
or U15356 (N_15356,N_9271,N_7609);
and U15357 (N_15357,N_7250,N_7554);
or U15358 (N_15358,N_8042,N_10260);
and U15359 (N_15359,N_7101,N_6696);
nor U15360 (N_15360,N_10443,N_8921);
nand U15361 (N_15361,N_6607,N_9230);
and U15362 (N_15362,N_10133,N_10380);
and U15363 (N_15363,N_12025,N_9605);
and U15364 (N_15364,N_10478,N_9148);
xnor U15365 (N_15365,N_7054,N_8750);
and U15366 (N_15366,N_8524,N_7922);
and U15367 (N_15367,N_8273,N_8376);
nand U15368 (N_15368,N_8641,N_6928);
nor U15369 (N_15369,N_9845,N_9643);
and U15370 (N_15370,N_8322,N_6440);
xnor U15371 (N_15371,N_9915,N_7472);
nand U15372 (N_15372,N_12188,N_8005);
or U15373 (N_15373,N_7057,N_8167);
nand U15374 (N_15374,N_10940,N_9555);
and U15375 (N_15375,N_8000,N_7825);
nand U15376 (N_15376,N_10979,N_11425);
nand U15377 (N_15377,N_9418,N_11504);
or U15378 (N_15378,N_9787,N_6651);
and U15379 (N_15379,N_12081,N_7770);
and U15380 (N_15380,N_7206,N_10475);
or U15381 (N_15381,N_6483,N_7417);
and U15382 (N_15382,N_7913,N_8948);
or U15383 (N_15383,N_11261,N_9099);
nor U15384 (N_15384,N_10714,N_12123);
xor U15385 (N_15385,N_11726,N_11316);
nand U15386 (N_15386,N_10382,N_7073);
or U15387 (N_15387,N_6370,N_11389);
nor U15388 (N_15388,N_7899,N_11161);
or U15389 (N_15389,N_11124,N_11273);
and U15390 (N_15390,N_8492,N_11048);
or U15391 (N_15391,N_11519,N_9635);
xnor U15392 (N_15392,N_7045,N_7902);
nand U15393 (N_15393,N_8829,N_12068);
nor U15394 (N_15394,N_8343,N_6276);
nor U15395 (N_15395,N_10124,N_9510);
nor U15396 (N_15396,N_9229,N_7463);
nor U15397 (N_15397,N_10012,N_9487);
and U15398 (N_15398,N_7317,N_6842);
nor U15399 (N_15399,N_6409,N_7932);
and U15400 (N_15400,N_8636,N_6738);
and U15401 (N_15401,N_6595,N_11065);
nand U15402 (N_15402,N_8356,N_7021);
nand U15403 (N_15403,N_8243,N_10296);
or U15404 (N_15404,N_7138,N_12060);
nor U15405 (N_15405,N_7772,N_12480);
nand U15406 (N_15406,N_12279,N_9580);
nor U15407 (N_15407,N_10218,N_7183);
and U15408 (N_15408,N_10454,N_7335);
and U15409 (N_15409,N_7671,N_11404);
and U15410 (N_15410,N_6895,N_7464);
or U15411 (N_15411,N_8748,N_8949);
and U15412 (N_15412,N_7917,N_7420);
and U15413 (N_15413,N_8828,N_10726);
or U15414 (N_15414,N_10658,N_11795);
nor U15415 (N_15415,N_8289,N_8061);
nand U15416 (N_15416,N_8264,N_12278);
nand U15417 (N_15417,N_8064,N_8320);
or U15418 (N_15418,N_6790,N_7008);
and U15419 (N_15419,N_11024,N_9161);
nor U15420 (N_15420,N_12075,N_9940);
xnor U15421 (N_15421,N_9193,N_11577);
nand U15422 (N_15422,N_8091,N_7706);
nand U15423 (N_15423,N_6269,N_10541);
or U15424 (N_15424,N_11231,N_11674);
nor U15425 (N_15425,N_6300,N_8621);
nand U15426 (N_15426,N_11549,N_8527);
or U15427 (N_15427,N_12311,N_9998);
or U15428 (N_15428,N_10001,N_9325);
or U15429 (N_15429,N_7527,N_8174);
and U15430 (N_15430,N_7763,N_7585);
nor U15431 (N_15431,N_6434,N_12086);
nand U15432 (N_15432,N_10209,N_11167);
or U15433 (N_15433,N_10074,N_6877);
nor U15434 (N_15434,N_8479,N_8188);
and U15435 (N_15435,N_6489,N_11729);
nor U15436 (N_15436,N_6426,N_8128);
nor U15437 (N_15437,N_11324,N_6879);
or U15438 (N_15438,N_7911,N_11035);
nand U15439 (N_15439,N_11772,N_10574);
nor U15440 (N_15440,N_8669,N_8194);
or U15441 (N_15441,N_10137,N_10764);
nand U15442 (N_15442,N_11767,N_9444);
and U15443 (N_15443,N_6912,N_9610);
and U15444 (N_15444,N_10086,N_10056);
or U15445 (N_15445,N_6471,N_9427);
nand U15446 (N_15446,N_9797,N_8884);
or U15447 (N_15447,N_8614,N_8799);
xnor U15448 (N_15448,N_11102,N_9647);
nor U15449 (N_15449,N_8145,N_8018);
xnor U15450 (N_15450,N_9296,N_6910);
or U15451 (N_15451,N_8426,N_7943);
nand U15452 (N_15452,N_6924,N_12099);
nand U15453 (N_15453,N_11001,N_7452);
nand U15454 (N_15454,N_9760,N_9776);
nand U15455 (N_15455,N_11508,N_11410);
nand U15456 (N_15456,N_7662,N_6865);
or U15457 (N_15457,N_11036,N_11226);
or U15458 (N_15458,N_6604,N_10332);
nor U15459 (N_15459,N_9898,N_8393);
or U15460 (N_15460,N_10901,N_7015);
nand U15461 (N_15461,N_7434,N_7233);
or U15462 (N_15462,N_11169,N_7835);
xnor U15463 (N_15463,N_6825,N_11654);
nor U15464 (N_15464,N_11533,N_10637);
nor U15465 (N_15465,N_8433,N_9038);
or U15466 (N_15466,N_11237,N_11029);
or U15467 (N_15467,N_8477,N_6639);
or U15468 (N_15468,N_10155,N_9462);
or U15469 (N_15469,N_10250,N_8936);
or U15470 (N_15470,N_11482,N_8189);
and U15471 (N_15471,N_9945,N_6467);
nor U15472 (N_15472,N_7474,N_7610);
nor U15473 (N_15473,N_7975,N_7824);
nand U15474 (N_15474,N_7023,N_7332);
nor U15475 (N_15475,N_8840,N_10666);
and U15476 (N_15476,N_12145,N_8218);
nor U15477 (N_15477,N_12072,N_11470);
nor U15478 (N_15478,N_11931,N_12211);
and U15479 (N_15479,N_7827,N_9476);
or U15480 (N_15480,N_11715,N_11241);
nand U15481 (N_15481,N_11733,N_7444);
or U15482 (N_15482,N_7162,N_8709);
and U15483 (N_15483,N_7484,N_6722);
nand U15484 (N_15484,N_7746,N_9164);
or U15485 (N_15485,N_11477,N_8147);
nand U15486 (N_15486,N_9417,N_6641);
and U15487 (N_15487,N_12325,N_12007);
and U15488 (N_15488,N_8328,N_10787);
xor U15489 (N_15489,N_9777,N_9399);
and U15490 (N_15490,N_8307,N_10039);
and U15491 (N_15491,N_10808,N_7066);
and U15492 (N_15492,N_6258,N_9810);
and U15493 (N_15493,N_11296,N_11181);
xor U15494 (N_15494,N_9981,N_6819);
xor U15495 (N_15495,N_6870,N_7579);
xor U15496 (N_15496,N_9367,N_8517);
or U15497 (N_15497,N_9629,N_7788);
nor U15498 (N_15498,N_10845,N_6389);
or U15499 (N_15499,N_7978,N_11184);
nand U15500 (N_15500,N_10902,N_12235);
and U15501 (N_15501,N_6801,N_6255);
and U15502 (N_15502,N_7449,N_6809);
or U15503 (N_15503,N_8447,N_10718);
or U15504 (N_15504,N_9262,N_11926);
or U15505 (N_15505,N_6523,N_8670);
and U15506 (N_15506,N_7287,N_8692);
nand U15507 (N_15507,N_11842,N_7075);
or U15508 (N_15508,N_11091,N_10487);
xnor U15509 (N_15509,N_9413,N_6445);
xor U15510 (N_15510,N_6750,N_9764);
nand U15511 (N_15511,N_11689,N_10677);
nand U15512 (N_15512,N_12297,N_9348);
and U15513 (N_15513,N_6433,N_9082);
nor U15514 (N_15514,N_7056,N_8069);
nor U15515 (N_15515,N_7800,N_12051);
or U15516 (N_15516,N_7058,N_8827);
and U15517 (N_15517,N_8304,N_9634);
nand U15518 (N_15518,N_7278,N_6961);
xor U15519 (N_15519,N_8470,N_6375);
and U15520 (N_15520,N_10110,N_7346);
nor U15521 (N_15521,N_6774,N_7789);
or U15522 (N_15522,N_9768,N_11611);
or U15523 (N_15523,N_8707,N_7737);
nand U15524 (N_15524,N_11274,N_11934);
or U15525 (N_15525,N_6711,N_12383);
nor U15526 (N_15526,N_9879,N_12083);
nand U15527 (N_15527,N_7809,N_10470);
nand U15528 (N_15528,N_7391,N_9018);
and U15529 (N_15529,N_11007,N_9467);
and U15530 (N_15530,N_8529,N_9067);
or U15531 (N_15531,N_10844,N_7360);
nor U15532 (N_15532,N_8181,N_11461);
or U15533 (N_15533,N_8029,N_11937);
and U15534 (N_15534,N_11152,N_8130);
nor U15535 (N_15535,N_7113,N_11558);
nand U15536 (N_15536,N_8338,N_12285);
xor U15537 (N_15537,N_6517,N_8378);
xnor U15538 (N_15538,N_8654,N_6658);
nor U15539 (N_15539,N_9246,N_9863);
nand U15540 (N_15540,N_10710,N_12148);
nor U15541 (N_15541,N_12266,N_8916);
and U15542 (N_15542,N_11638,N_10805);
and U15543 (N_15543,N_9973,N_7145);
nand U15544 (N_15544,N_11437,N_12220);
nand U15545 (N_15545,N_10024,N_9607);
nand U15546 (N_15546,N_12448,N_7850);
nand U15547 (N_15547,N_6572,N_12004);
nand U15548 (N_15548,N_10938,N_9601);
nand U15549 (N_15549,N_6730,N_8563);
nor U15550 (N_15550,N_8033,N_8265);
nor U15551 (N_15551,N_7009,N_9727);
xor U15552 (N_15552,N_10520,N_8213);
or U15553 (N_15553,N_11529,N_6882);
nor U15554 (N_15554,N_11615,N_10634);
nor U15555 (N_15555,N_12212,N_10498);
nor U15556 (N_15556,N_11682,N_11602);
and U15557 (N_15557,N_7300,N_9584);
and U15558 (N_15558,N_10895,N_9929);
or U15559 (N_15559,N_7982,N_9969);
or U15560 (N_15560,N_8429,N_7202);
nor U15561 (N_15561,N_10552,N_6294);
and U15562 (N_15562,N_12287,N_11745);
xor U15563 (N_15563,N_10820,N_9461);
and U15564 (N_15564,N_10615,N_7890);
nor U15565 (N_15565,N_10381,N_10472);
nand U15566 (N_15566,N_9370,N_11276);
and U15567 (N_15567,N_8295,N_11287);
or U15568 (N_15568,N_6346,N_9548);
and U15569 (N_15569,N_10489,N_9324);
or U15570 (N_15570,N_11543,N_11407);
or U15571 (N_15571,N_6435,N_9092);
or U15572 (N_15572,N_8554,N_8857);
and U15573 (N_15573,N_7897,N_11884);
or U15574 (N_15574,N_8534,N_11575);
xor U15575 (N_15575,N_10084,N_6643);
nand U15576 (N_15576,N_7689,N_7876);
nand U15577 (N_15577,N_8955,N_7249);
and U15578 (N_15578,N_10353,N_11387);
xnor U15579 (N_15579,N_9227,N_10639);
and U15580 (N_15580,N_10310,N_9397);
and U15581 (N_15581,N_8068,N_7301);
nor U15582 (N_15582,N_11586,N_11483);
nand U15583 (N_15583,N_7268,N_6939);
nand U15584 (N_15584,N_7928,N_12465);
nand U15585 (N_15585,N_7217,N_9006);
xor U15586 (N_15586,N_8664,N_11472);
nor U15587 (N_15587,N_8785,N_9298);
xnor U15588 (N_15588,N_7637,N_6739);
nor U15589 (N_15589,N_8794,N_8475);
nand U15590 (N_15590,N_6975,N_9913);
xor U15591 (N_15591,N_11222,N_9020);
nand U15592 (N_15592,N_6492,N_11990);
or U15593 (N_15593,N_11636,N_7845);
and U15594 (N_15594,N_12352,N_8357);
or U15595 (N_15595,N_7010,N_10957);
nor U15596 (N_15596,N_10465,N_7502);
nand U15597 (N_15597,N_12360,N_11888);
and U15598 (N_15598,N_8382,N_9639);
and U15599 (N_15599,N_6768,N_6676);
and U15600 (N_15600,N_7791,N_8471);
nand U15601 (N_15601,N_10032,N_10993);
and U15602 (N_15602,N_6755,N_11303);
nand U15603 (N_15603,N_11641,N_7059);
or U15604 (N_15604,N_10659,N_6807);
nor U15605 (N_15605,N_9781,N_8481);
nand U15606 (N_15606,N_9516,N_11608);
nand U15607 (N_15607,N_11603,N_10978);
nand U15608 (N_15608,N_8531,N_7664);
and U15609 (N_15609,N_10742,N_10101);
nand U15610 (N_15610,N_9866,N_12452);
nor U15611 (N_15611,N_8150,N_11814);
nor U15612 (N_15612,N_6655,N_8386);
xor U15613 (N_15613,N_10660,N_8606);
or U15614 (N_15614,N_11185,N_11520);
and U15615 (N_15615,N_10185,N_9564);
nor U15616 (N_15616,N_10370,N_12244);
or U15617 (N_15617,N_9139,N_10438);
or U15618 (N_15618,N_8581,N_8876);
nor U15619 (N_15619,N_11335,N_9331);
and U15620 (N_15620,N_10676,N_8920);
and U15621 (N_15621,N_9439,N_6415);
nor U15622 (N_15622,N_7412,N_7701);
nor U15623 (N_15623,N_10140,N_10228);
or U15624 (N_15624,N_11857,N_10053);
nor U15625 (N_15625,N_9790,N_8928);
and U15626 (N_15626,N_9835,N_11228);
nor U15627 (N_15627,N_9934,N_10857);
and U15628 (N_15628,N_10923,N_7987);
nand U15629 (N_15629,N_8555,N_9644);
or U15630 (N_15630,N_11562,N_9905);
nand U15631 (N_15631,N_7289,N_6427);
nand U15632 (N_15632,N_9910,N_10275);
or U15633 (N_15633,N_6643,N_10211);
nand U15634 (N_15634,N_9330,N_9931);
and U15635 (N_15635,N_11077,N_6944);
and U15636 (N_15636,N_6714,N_11618);
or U15637 (N_15637,N_9350,N_9852);
nand U15638 (N_15638,N_8988,N_7513);
and U15639 (N_15639,N_9486,N_9854);
and U15640 (N_15640,N_8531,N_8957);
and U15641 (N_15641,N_7338,N_11433);
or U15642 (N_15642,N_11642,N_7369);
nand U15643 (N_15643,N_6969,N_8671);
or U15644 (N_15644,N_11873,N_10613);
nand U15645 (N_15645,N_9098,N_9231);
nor U15646 (N_15646,N_9029,N_7508);
or U15647 (N_15647,N_9043,N_6686);
nor U15648 (N_15648,N_9858,N_11851);
and U15649 (N_15649,N_10109,N_7396);
nand U15650 (N_15650,N_6910,N_7665);
or U15651 (N_15651,N_7840,N_8851);
xnor U15652 (N_15652,N_12267,N_7737);
or U15653 (N_15653,N_8575,N_6932);
nand U15654 (N_15654,N_9529,N_10759);
xor U15655 (N_15655,N_10365,N_9735);
or U15656 (N_15656,N_10327,N_9275);
and U15657 (N_15657,N_8300,N_12004);
nor U15658 (N_15658,N_11285,N_10588);
or U15659 (N_15659,N_8029,N_11647);
nand U15660 (N_15660,N_10295,N_12397);
or U15661 (N_15661,N_10441,N_6309);
nor U15662 (N_15662,N_10601,N_8513);
and U15663 (N_15663,N_11270,N_12182);
and U15664 (N_15664,N_12073,N_7289);
or U15665 (N_15665,N_11677,N_7875);
nand U15666 (N_15666,N_11019,N_8135);
or U15667 (N_15667,N_9885,N_7278);
nor U15668 (N_15668,N_6914,N_8606);
and U15669 (N_15669,N_10669,N_11124);
and U15670 (N_15670,N_8652,N_12110);
nor U15671 (N_15671,N_11048,N_9561);
nand U15672 (N_15672,N_11990,N_6830);
nor U15673 (N_15673,N_11637,N_11462);
and U15674 (N_15674,N_9828,N_8325);
and U15675 (N_15675,N_7473,N_10909);
or U15676 (N_15676,N_11578,N_12393);
xor U15677 (N_15677,N_12292,N_11340);
nor U15678 (N_15678,N_9179,N_12060);
and U15679 (N_15679,N_8757,N_8598);
nand U15680 (N_15680,N_11957,N_10482);
nand U15681 (N_15681,N_10373,N_10439);
and U15682 (N_15682,N_10914,N_8304);
nand U15683 (N_15683,N_7782,N_11519);
nand U15684 (N_15684,N_11257,N_7657);
and U15685 (N_15685,N_7938,N_12188);
nand U15686 (N_15686,N_12423,N_9669);
xor U15687 (N_15687,N_8110,N_12467);
nor U15688 (N_15688,N_10585,N_6673);
nand U15689 (N_15689,N_12154,N_9036);
nand U15690 (N_15690,N_8206,N_8631);
or U15691 (N_15691,N_9955,N_6633);
and U15692 (N_15692,N_7152,N_11294);
and U15693 (N_15693,N_9948,N_6414);
nor U15694 (N_15694,N_9671,N_6591);
and U15695 (N_15695,N_12091,N_11947);
or U15696 (N_15696,N_7882,N_7782);
or U15697 (N_15697,N_9871,N_7816);
or U15698 (N_15698,N_6614,N_6408);
nand U15699 (N_15699,N_10652,N_7747);
or U15700 (N_15700,N_6562,N_10182);
and U15701 (N_15701,N_9359,N_11876);
and U15702 (N_15702,N_8967,N_10271);
or U15703 (N_15703,N_7886,N_7603);
xor U15704 (N_15704,N_10267,N_6412);
nand U15705 (N_15705,N_7478,N_6875);
or U15706 (N_15706,N_8961,N_11408);
or U15707 (N_15707,N_12013,N_9592);
or U15708 (N_15708,N_10347,N_11478);
or U15709 (N_15709,N_8412,N_12057);
xor U15710 (N_15710,N_8144,N_8697);
or U15711 (N_15711,N_10424,N_11234);
or U15712 (N_15712,N_9588,N_9089);
nor U15713 (N_15713,N_11645,N_9813);
or U15714 (N_15714,N_7600,N_9046);
xnor U15715 (N_15715,N_10447,N_7296);
nand U15716 (N_15716,N_9166,N_10967);
and U15717 (N_15717,N_10503,N_12139);
and U15718 (N_15718,N_6805,N_6997);
or U15719 (N_15719,N_9305,N_8125);
xnor U15720 (N_15720,N_6371,N_10209);
or U15721 (N_15721,N_10303,N_8633);
xor U15722 (N_15722,N_8565,N_6813);
or U15723 (N_15723,N_8289,N_7391);
nand U15724 (N_15724,N_11290,N_10658);
or U15725 (N_15725,N_7575,N_7379);
nor U15726 (N_15726,N_6269,N_7922);
nor U15727 (N_15727,N_11965,N_9158);
xor U15728 (N_15728,N_7746,N_10111);
or U15729 (N_15729,N_9183,N_6588);
nor U15730 (N_15730,N_8934,N_10252);
nand U15731 (N_15731,N_12493,N_7327);
nand U15732 (N_15732,N_7366,N_7319);
and U15733 (N_15733,N_12402,N_10061);
or U15734 (N_15734,N_9392,N_8455);
nor U15735 (N_15735,N_10426,N_10031);
and U15736 (N_15736,N_9932,N_8723);
and U15737 (N_15737,N_8608,N_11952);
nand U15738 (N_15738,N_11593,N_6471);
or U15739 (N_15739,N_7092,N_6656);
nand U15740 (N_15740,N_6815,N_10398);
or U15741 (N_15741,N_10893,N_7817);
nor U15742 (N_15742,N_12465,N_7167);
nand U15743 (N_15743,N_7177,N_11561);
nor U15744 (N_15744,N_7559,N_11790);
or U15745 (N_15745,N_10858,N_7080);
xnor U15746 (N_15746,N_9574,N_6862);
nor U15747 (N_15747,N_7684,N_8433);
or U15748 (N_15748,N_8547,N_11177);
nand U15749 (N_15749,N_12253,N_12146);
and U15750 (N_15750,N_10682,N_10800);
nor U15751 (N_15751,N_8489,N_9126);
and U15752 (N_15752,N_8303,N_7087);
xnor U15753 (N_15753,N_7809,N_9848);
or U15754 (N_15754,N_10799,N_10740);
nand U15755 (N_15755,N_11392,N_11332);
and U15756 (N_15756,N_8787,N_8724);
nor U15757 (N_15757,N_9691,N_11120);
and U15758 (N_15758,N_11473,N_12079);
or U15759 (N_15759,N_7868,N_10133);
and U15760 (N_15760,N_9201,N_8006);
and U15761 (N_15761,N_6376,N_8111);
and U15762 (N_15762,N_6415,N_10879);
nor U15763 (N_15763,N_8168,N_10552);
and U15764 (N_15764,N_6437,N_12210);
xnor U15765 (N_15765,N_9524,N_8145);
nor U15766 (N_15766,N_10084,N_11922);
nand U15767 (N_15767,N_7376,N_12334);
xnor U15768 (N_15768,N_9140,N_11749);
and U15769 (N_15769,N_9914,N_6580);
or U15770 (N_15770,N_7303,N_8267);
and U15771 (N_15771,N_10650,N_10387);
nor U15772 (N_15772,N_10457,N_6731);
xnor U15773 (N_15773,N_7906,N_8904);
nand U15774 (N_15774,N_8236,N_10087);
or U15775 (N_15775,N_9459,N_11899);
nor U15776 (N_15776,N_8426,N_7784);
or U15777 (N_15777,N_6774,N_11177);
nand U15778 (N_15778,N_7979,N_10615);
nor U15779 (N_15779,N_8452,N_8359);
nor U15780 (N_15780,N_6280,N_9606);
nor U15781 (N_15781,N_9168,N_8318);
and U15782 (N_15782,N_12133,N_8502);
and U15783 (N_15783,N_6260,N_7939);
or U15784 (N_15784,N_10201,N_9388);
nand U15785 (N_15785,N_11964,N_6676);
nand U15786 (N_15786,N_8718,N_8764);
or U15787 (N_15787,N_12248,N_7155);
nor U15788 (N_15788,N_12361,N_11186);
or U15789 (N_15789,N_6724,N_11815);
nor U15790 (N_15790,N_12139,N_11694);
or U15791 (N_15791,N_10633,N_8127);
or U15792 (N_15792,N_12176,N_8556);
nor U15793 (N_15793,N_7049,N_11703);
or U15794 (N_15794,N_6374,N_9864);
and U15795 (N_15795,N_7546,N_7491);
and U15796 (N_15796,N_12175,N_7346);
nand U15797 (N_15797,N_8376,N_6845);
or U15798 (N_15798,N_12335,N_6434);
nor U15799 (N_15799,N_10328,N_7302);
and U15800 (N_15800,N_10476,N_8820);
nor U15801 (N_15801,N_9253,N_10444);
nor U15802 (N_15802,N_11784,N_7952);
and U15803 (N_15803,N_9909,N_7786);
nand U15804 (N_15804,N_7495,N_6947);
nand U15805 (N_15805,N_12449,N_7285);
nor U15806 (N_15806,N_8594,N_7149);
nor U15807 (N_15807,N_11647,N_6374);
and U15808 (N_15808,N_9515,N_6611);
nor U15809 (N_15809,N_6278,N_8469);
or U15810 (N_15810,N_6934,N_12374);
nor U15811 (N_15811,N_8709,N_10289);
nor U15812 (N_15812,N_8557,N_6374);
nand U15813 (N_15813,N_11756,N_9936);
nand U15814 (N_15814,N_10176,N_6591);
nor U15815 (N_15815,N_9010,N_8657);
nand U15816 (N_15816,N_8212,N_7642);
and U15817 (N_15817,N_10442,N_9176);
nor U15818 (N_15818,N_9893,N_11886);
or U15819 (N_15819,N_9322,N_6922);
or U15820 (N_15820,N_10678,N_11489);
nand U15821 (N_15821,N_9519,N_6853);
xnor U15822 (N_15822,N_8765,N_9948);
and U15823 (N_15823,N_9155,N_11039);
xor U15824 (N_15824,N_10647,N_9752);
nor U15825 (N_15825,N_10264,N_10864);
xor U15826 (N_15826,N_7943,N_11833);
or U15827 (N_15827,N_11854,N_8948);
nor U15828 (N_15828,N_8076,N_9842);
nor U15829 (N_15829,N_10014,N_11803);
and U15830 (N_15830,N_12258,N_6901);
or U15831 (N_15831,N_9007,N_10988);
or U15832 (N_15832,N_10586,N_7587);
and U15833 (N_15833,N_8534,N_8832);
nand U15834 (N_15834,N_7880,N_9144);
xor U15835 (N_15835,N_10143,N_11743);
or U15836 (N_15836,N_7788,N_11360);
nor U15837 (N_15837,N_10162,N_10205);
nand U15838 (N_15838,N_7582,N_7096);
and U15839 (N_15839,N_9382,N_9256);
and U15840 (N_15840,N_10805,N_12345);
nor U15841 (N_15841,N_7613,N_11251);
nand U15842 (N_15842,N_11717,N_8235);
or U15843 (N_15843,N_6902,N_12049);
nand U15844 (N_15844,N_10471,N_12336);
nor U15845 (N_15845,N_8909,N_8500);
nor U15846 (N_15846,N_9105,N_12049);
and U15847 (N_15847,N_9093,N_11744);
or U15848 (N_15848,N_8630,N_8550);
or U15849 (N_15849,N_10149,N_7943);
or U15850 (N_15850,N_9289,N_12372);
xnor U15851 (N_15851,N_9098,N_7784);
nor U15852 (N_15852,N_9534,N_6632);
or U15853 (N_15853,N_11273,N_8843);
or U15854 (N_15854,N_6488,N_7458);
or U15855 (N_15855,N_8158,N_8878);
nor U15856 (N_15856,N_6334,N_10847);
xor U15857 (N_15857,N_9966,N_6641);
nand U15858 (N_15858,N_11254,N_10514);
and U15859 (N_15859,N_8440,N_7693);
nand U15860 (N_15860,N_9599,N_11036);
or U15861 (N_15861,N_9857,N_7235);
and U15862 (N_15862,N_6877,N_7282);
nand U15863 (N_15863,N_10406,N_9191);
or U15864 (N_15864,N_6489,N_8243);
or U15865 (N_15865,N_8058,N_12392);
nor U15866 (N_15866,N_9797,N_11356);
nand U15867 (N_15867,N_9364,N_10465);
or U15868 (N_15868,N_12219,N_9066);
nand U15869 (N_15869,N_10119,N_10885);
nand U15870 (N_15870,N_9489,N_10276);
nand U15871 (N_15871,N_8465,N_6777);
and U15872 (N_15872,N_7177,N_6372);
nor U15873 (N_15873,N_9863,N_9320);
and U15874 (N_15874,N_12384,N_6548);
nor U15875 (N_15875,N_8996,N_6937);
xnor U15876 (N_15876,N_12205,N_10558);
or U15877 (N_15877,N_12055,N_9648);
nor U15878 (N_15878,N_11317,N_7451);
and U15879 (N_15879,N_6459,N_6508);
xnor U15880 (N_15880,N_6870,N_9035);
or U15881 (N_15881,N_9825,N_6855);
nand U15882 (N_15882,N_12236,N_10659);
nand U15883 (N_15883,N_6369,N_7770);
xor U15884 (N_15884,N_10380,N_7241);
nor U15885 (N_15885,N_9608,N_9049);
nand U15886 (N_15886,N_6857,N_9093);
and U15887 (N_15887,N_11671,N_7534);
or U15888 (N_15888,N_9139,N_8224);
and U15889 (N_15889,N_12482,N_9119);
nor U15890 (N_15890,N_10114,N_9193);
nor U15891 (N_15891,N_9335,N_11814);
nand U15892 (N_15892,N_9523,N_8401);
or U15893 (N_15893,N_8767,N_11932);
and U15894 (N_15894,N_7269,N_6686);
nand U15895 (N_15895,N_10109,N_6694);
nor U15896 (N_15896,N_9712,N_10482);
nand U15897 (N_15897,N_12165,N_10680);
or U15898 (N_15898,N_6353,N_7668);
and U15899 (N_15899,N_8328,N_12324);
nor U15900 (N_15900,N_10339,N_6852);
and U15901 (N_15901,N_9042,N_7105);
or U15902 (N_15902,N_7126,N_7311);
nand U15903 (N_15903,N_6685,N_6319);
and U15904 (N_15904,N_6533,N_9865);
nor U15905 (N_15905,N_7305,N_6918);
nor U15906 (N_15906,N_9316,N_6655);
xnor U15907 (N_15907,N_10116,N_9849);
or U15908 (N_15908,N_11658,N_8384);
and U15909 (N_15909,N_6314,N_7559);
or U15910 (N_15910,N_7996,N_7037);
nor U15911 (N_15911,N_6637,N_7313);
or U15912 (N_15912,N_9331,N_11422);
nor U15913 (N_15913,N_10166,N_10855);
nand U15914 (N_15914,N_8952,N_9350);
or U15915 (N_15915,N_7689,N_7453);
and U15916 (N_15916,N_8461,N_12372);
xor U15917 (N_15917,N_12382,N_11208);
nand U15918 (N_15918,N_7430,N_7925);
nand U15919 (N_15919,N_12311,N_9993);
nor U15920 (N_15920,N_9559,N_11761);
or U15921 (N_15921,N_11327,N_9981);
or U15922 (N_15922,N_8168,N_6696);
xor U15923 (N_15923,N_11395,N_12433);
nor U15924 (N_15924,N_8328,N_9233);
nand U15925 (N_15925,N_11056,N_8416);
nand U15926 (N_15926,N_11724,N_6369);
nor U15927 (N_15927,N_9626,N_10332);
nor U15928 (N_15928,N_8042,N_7950);
or U15929 (N_15929,N_8538,N_11181);
or U15930 (N_15930,N_10594,N_12337);
nor U15931 (N_15931,N_8839,N_7260);
nand U15932 (N_15932,N_10098,N_8387);
nand U15933 (N_15933,N_10599,N_8053);
nor U15934 (N_15934,N_11519,N_9661);
xnor U15935 (N_15935,N_9638,N_7631);
nor U15936 (N_15936,N_6682,N_10984);
or U15937 (N_15937,N_7509,N_9575);
and U15938 (N_15938,N_8822,N_10607);
xor U15939 (N_15939,N_6790,N_12168);
or U15940 (N_15940,N_10501,N_11260);
or U15941 (N_15941,N_6682,N_9567);
nand U15942 (N_15942,N_9515,N_6813);
and U15943 (N_15943,N_11649,N_11676);
or U15944 (N_15944,N_11239,N_10925);
nand U15945 (N_15945,N_11694,N_12238);
and U15946 (N_15946,N_9498,N_6840);
and U15947 (N_15947,N_10646,N_10209);
and U15948 (N_15948,N_8906,N_9239);
nor U15949 (N_15949,N_7335,N_7250);
nor U15950 (N_15950,N_7197,N_7664);
or U15951 (N_15951,N_6684,N_7499);
and U15952 (N_15952,N_9856,N_11461);
nor U15953 (N_15953,N_7958,N_7287);
nor U15954 (N_15954,N_6630,N_10234);
nor U15955 (N_15955,N_9659,N_12095);
and U15956 (N_15956,N_9525,N_9684);
nor U15957 (N_15957,N_8779,N_12051);
and U15958 (N_15958,N_11466,N_10311);
nor U15959 (N_15959,N_11434,N_8776);
or U15960 (N_15960,N_8416,N_11316);
nand U15961 (N_15961,N_10827,N_7709);
nor U15962 (N_15962,N_9120,N_10678);
or U15963 (N_15963,N_9218,N_7645);
and U15964 (N_15964,N_8061,N_9252);
or U15965 (N_15965,N_10275,N_8353);
or U15966 (N_15966,N_8673,N_10456);
and U15967 (N_15967,N_11723,N_11063);
nor U15968 (N_15968,N_9844,N_8123);
nor U15969 (N_15969,N_10530,N_8071);
or U15970 (N_15970,N_9779,N_11248);
nor U15971 (N_15971,N_11675,N_8151);
xnor U15972 (N_15972,N_8150,N_11695);
nor U15973 (N_15973,N_12189,N_11355);
and U15974 (N_15974,N_8753,N_7421);
nor U15975 (N_15975,N_12335,N_9898);
or U15976 (N_15976,N_12262,N_8620);
nand U15977 (N_15977,N_6274,N_9181);
and U15978 (N_15978,N_10584,N_9300);
nor U15979 (N_15979,N_9451,N_6344);
or U15980 (N_15980,N_7036,N_8639);
and U15981 (N_15981,N_7177,N_11111);
nand U15982 (N_15982,N_12110,N_6999);
nand U15983 (N_15983,N_8199,N_6724);
and U15984 (N_15984,N_7059,N_7394);
and U15985 (N_15985,N_9376,N_6281);
or U15986 (N_15986,N_10187,N_10674);
and U15987 (N_15987,N_9152,N_8709);
xnor U15988 (N_15988,N_10833,N_7555);
nor U15989 (N_15989,N_10573,N_11755);
nor U15990 (N_15990,N_10433,N_7677);
nor U15991 (N_15991,N_7441,N_9789);
and U15992 (N_15992,N_8512,N_10053);
nand U15993 (N_15993,N_12414,N_9718);
nand U15994 (N_15994,N_11059,N_8348);
or U15995 (N_15995,N_6298,N_8527);
nand U15996 (N_15996,N_9433,N_8676);
and U15997 (N_15997,N_7418,N_11244);
or U15998 (N_15998,N_10439,N_7000);
nor U15999 (N_15999,N_11770,N_8562);
or U16000 (N_16000,N_6726,N_7929);
nand U16001 (N_16001,N_9381,N_11073);
and U16002 (N_16002,N_7424,N_9029);
or U16003 (N_16003,N_9184,N_11311);
or U16004 (N_16004,N_6587,N_7553);
or U16005 (N_16005,N_10399,N_11261);
or U16006 (N_16006,N_11297,N_7263);
and U16007 (N_16007,N_7770,N_7057);
or U16008 (N_16008,N_8345,N_8728);
nor U16009 (N_16009,N_9729,N_7796);
and U16010 (N_16010,N_8722,N_8175);
and U16011 (N_16011,N_7825,N_9932);
nor U16012 (N_16012,N_6458,N_9354);
or U16013 (N_16013,N_10890,N_6302);
nand U16014 (N_16014,N_8624,N_8396);
or U16015 (N_16015,N_11745,N_12273);
or U16016 (N_16016,N_10796,N_7123);
and U16017 (N_16017,N_10165,N_7054);
nand U16018 (N_16018,N_9326,N_11923);
and U16019 (N_16019,N_7922,N_8209);
nand U16020 (N_16020,N_8303,N_12103);
nor U16021 (N_16021,N_8131,N_7635);
or U16022 (N_16022,N_10105,N_7137);
nor U16023 (N_16023,N_8570,N_7232);
xor U16024 (N_16024,N_11965,N_9594);
nor U16025 (N_16025,N_6641,N_12021);
xor U16026 (N_16026,N_10360,N_8788);
or U16027 (N_16027,N_8757,N_11558);
nand U16028 (N_16028,N_6547,N_11548);
nor U16029 (N_16029,N_8687,N_9895);
nand U16030 (N_16030,N_7322,N_8468);
and U16031 (N_16031,N_7880,N_6768);
and U16032 (N_16032,N_11738,N_10121);
nor U16033 (N_16033,N_11543,N_10848);
nand U16034 (N_16034,N_6438,N_7547);
xnor U16035 (N_16035,N_10317,N_10716);
or U16036 (N_16036,N_7606,N_6509);
nor U16037 (N_16037,N_8587,N_11687);
or U16038 (N_16038,N_11428,N_12298);
or U16039 (N_16039,N_8483,N_6559);
nand U16040 (N_16040,N_8107,N_7553);
and U16041 (N_16041,N_8760,N_7871);
and U16042 (N_16042,N_7842,N_6269);
nor U16043 (N_16043,N_9635,N_11779);
nor U16044 (N_16044,N_6310,N_9859);
nand U16045 (N_16045,N_6308,N_7261);
nand U16046 (N_16046,N_6742,N_7706);
and U16047 (N_16047,N_6463,N_12246);
and U16048 (N_16048,N_12103,N_9331);
nand U16049 (N_16049,N_11948,N_10059);
nor U16050 (N_16050,N_8590,N_9476);
nor U16051 (N_16051,N_11466,N_8486);
nor U16052 (N_16052,N_11582,N_7751);
nor U16053 (N_16053,N_6394,N_10414);
xnor U16054 (N_16054,N_6851,N_8992);
or U16055 (N_16055,N_12348,N_12282);
nor U16056 (N_16056,N_10009,N_9061);
and U16057 (N_16057,N_11540,N_12323);
and U16058 (N_16058,N_7180,N_9244);
or U16059 (N_16059,N_10974,N_7946);
nand U16060 (N_16060,N_11881,N_8603);
xnor U16061 (N_16061,N_12412,N_10793);
nand U16062 (N_16062,N_7286,N_11318);
or U16063 (N_16063,N_9038,N_6748);
nand U16064 (N_16064,N_10999,N_6629);
xnor U16065 (N_16065,N_6418,N_10340);
or U16066 (N_16066,N_6677,N_9954);
nor U16067 (N_16067,N_10191,N_11172);
nand U16068 (N_16068,N_8683,N_6637);
nor U16069 (N_16069,N_9535,N_11983);
nand U16070 (N_16070,N_12134,N_8618);
nor U16071 (N_16071,N_10553,N_9054);
nand U16072 (N_16072,N_9493,N_9524);
and U16073 (N_16073,N_8964,N_7396);
nor U16074 (N_16074,N_6711,N_9234);
nand U16075 (N_16075,N_6712,N_11621);
nand U16076 (N_16076,N_10179,N_11798);
or U16077 (N_16077,N_10425,N_8160);
nor U16078 (N_16078,N_11440,N_9115);
nand U16079 (N_16079,N_11834,N_12010);
nand U16080 (N_16080,N_10561,N_11820);
nor U16081 (N_16081,N_7858,N_8031);
nand U16082 (N_16082,N_10692,N_8651);
nand U16083 (N_16083,N_12059,N_11720);
or U16084 (N_16084,N_10717,N_8803);
nor U16085 (N_16085,N_7932,N_11269);
or U16086 (N_16086,N_11376,N_8855);
xor U16087 (N_16087,N_11933,N_7215);
or U16088 (N_16088,N_7716,N_7466);
nor U16089 (N_16089,N_11843,N_6690);
nand U16090 (N_16090,N_10790,N_8963);
and U16091 (N_16091,N_9970,N_10399);
and U16092 (N_16092,N_8319,N_11007);
and U16093 (N_16093,N_9080,N_7535);
or U16094 (N_16094,N_6579,N_9223);
nand U16095 (N_16095,N_11808,N_12060);
nor U16096 (N_16096,N_7477,N_6798);
nor U16097 (N_16097,N_8055,N_6543);
or U16098 (N_16098,N_11261,N_10097);
nor U16099 (N_16099,N_7942,N_10376);
or U16100 (N_16100,N_8518,N_9415);
nand U16101 (N_16101,N_11090,N_7775);
or U16102 (N_16102,N_6373,N_11430);
xnor U16103 (N_16103,N_12114,N_10569);
and U16104 (N_16104,N_6265,N_6613);
and U16105 (N_16105,N_6737,N_9479);
nand U16106 (N_16106,N_9813,N_11263);
or U16107 (N_16107,N_8823,N_12226);
or U16108 (N_16108,N_10802,N_10370);
nand U16109 (N_16109,N_9748,N_8191);
and U16110 (N_16110,N_8192,N_9616);
and U16111 (N_16111,N_10305,N_8530);
xor U16112 (N_16112,N_11099,N_9234);
and U16113 (N_16113,N_10142,N_8101);
nor U16114 (N_16114,N_7126,N_6588);
or U16115 (N_16115,N_8779,N_11734);
and U16116 (N_16116,N_8291,N_6625);
or U16117 (N_16117,N_8804,N_8451);
or U16118 (N_16118,N_7521,N_10284);
nor U16119 (N_16119,N_11882,N_6679);
nand U16120 (N_16120,N_10180,N_12069);
nor U16121 (N_16121,N_11717,N_9389);
or U16122 (N_16122,N_10803,N_10097);
nand U16123 (N_16123,N_6737,N_11962);
nor U16124 (N_16124,N_6828,N_10189);
and U16125 (N_16125,N_10914,N_9663);
or U16126 (N_16126,N_6589,N_12372);
nor U16127 (N_16127,N_8656,N_10010);
or U16128 (N_16128,N_8872,N_6742);
or U16129 (N_16129,N_8157,N_10972);
nand U16130 (N_16130,N_10589,N_9156);
nand U16131 (N_16131,N_10557,N_8116);
or U16132 (N_16132,N_10982,N_12431);
nand U16133 (N_16133,N_10289,N_7895);
or U16134 (N_16134,N_8036,N_10361);
or U16135 (N_16135,N_11255,N_11768);
nand U16136 (N_16136,N_6510,N_11179);
nor U16137 (N_16137,N_10154,N_10507);
or U16138 (N_16138,N_11716,N_11873);
xnor U16139 (N_16139,N_10893,N_11144);
xor U16140 (N_16140,N_10628,N_7546);
and U16141 (N_16141,N_12437,N_8553);
and U16142 (N_16142,N_7654,N_7304);
xor U16143 (N_16143,N_9655,N_8876);
nor U16144 (N_16144,N_7162,N_7580);
nor U16145 (N_16145,N_11137,N_8537);
or U16146 (N_16146,N_8454,N_9207);
and U16147 (N_16147,N_9523,N_7799);
nand U16148 (N_16148,N_6990,N_11159);
nor U16149 (N_16149,N_7694,N_8366);
and U16150 (N_16150,N_7876,N_10224);
and U16151 (N_16151,N_11234,N_12236);
xnor U16152 (N_16152,N_9628,N_8841);
or U16153 (N_16153,N_9352,N_10296);
xnor U16154 (N_16154,N_7925,N_11519);
xor U16155 (N_16155,N_6491,N_11097);
and U16156 (N_16156,N_6941,N_10151);
nor U16157 (N_16157,N_8011,N_6962);
or U16158 (N_16158,N_6729,N_8505);
or U16159 (N_16159,N_10187,N_7767);
nor U16160 (N_16160,N_7082,N_6999);
and U16161 (N_16161,N_10634,N_9436);
nand U16162 (N_16162,N_10686,N_8341);
nand U16163 (N_16163,N_10903,N_6653);
and U16164 (N_16164,N_10882,N_7544);
nor U16165 (N_16165,N_7603,N_7615);
and U16166 (N_16166,N_10872,N_12010);
nand U16167 (N_16167,N_7997,N_9907);
nand U16168 (N_16168,N_11507,N_8235);
and U16169 (N_16169,N_8551,N_9281);
and U16170 (N_16170,N_11655,N_10753);
or U16171 (N_16171,N_11607,N_11107);
or U16172 (N_16172,N_7676,N_8046);
or U16173 (N_16173,N_6277,N_7292);
and U16174 (N_16174,N_10640,N_8631);
nand U16175 (N_16175,N_11938,N_7396);
xnor U16176 (N_16176,N_10615,N_10216);
or U16177 (N_16177,N_11539,N_7932);
and U16178 (N_16178,N_8349,N_8155);
nor U16179 (N_16179,N_6304,N_9563);
and U16180 (N_16180,N_6791,N_11672);
nand U16181 (N_16181,N_7038,N_9833);
and U16182 (N_16182,N_12368,N_10800);
xor U16183 (N_16183,N_10572,N_6855);
and U16184 (N_16184,N_11295,N_12346);
and U16185 (N_16185,N_12334,N_7790);
nor U16186 (N_16186,N_12261,N_11517);
and U16187 (N_16187,N_11967,N_8714);
and U16188 (N_16188,N_12345,N_11155);
nand U16189 (N_16189,N_8039,N_10173);
nor U16190 (N_16190,N_7616,N_6359);
or U16191 (N_16191,N_11383,N_8044);
and U16192 (N_16192,N_7267,N_11880);
or U16193 (N_16193,N_7881,N_10572);
nor U16194 (N_16194,N_6958,N_6388);
and U16195 (N_16195,N_11064,N_6397);
nor U16196 (N_16196,N_10672,N_9058);
and U16197 (N_16197,N_9575,N_12459);
nor U16198 (N_16198,N_6773,N_8777);
or U16199 (N_16199,N_9229,N_7199);
and U16200 (N_16200,N_8631,N_10707);
nor U16201 (N_16201,N_10873,N_6638);
or U16202 (N_16202,N_11729,N_11835);
nor U16203 (N_16203,N_7119,N_8362);
nand U16204 (N_16204,N_7096,N_7968);
nor U16205 (N_16205,N_11984,N_8487);
and U16206 (N_16206,N_8033,N_10284);
or U16207 (N_16207,N_10427,N_10063);
nand U16208 (N_16208,N_8722,N_11631);
and U16209 (N_16209,N_8358,N_7528);
nor U16210 (N_16210,N_7792,N_10091);
nor U16211 (N_16211,N_9963,N_7145);
and U16212 (N_16212,N_10668,N_7792);
or U16213 (N_16213,N_8400,N_7600);
nor U16214 (N_16214,N_7407,N_9152);
and U16215 (N_16215,N_6969,N_9916);
and U16216 (N_16216,N_11714,N_8431);
or U16217 (N_16217,N_8572,N_8099);
or U16218 (N_16218,N_7747,N_10722);
or U16219 (N_16219,N_8058,N_9542);
xor U16220 (N_16220,N_11998,N_6588);
and U16221 (N_16221,N_9001,N_11805);
or U16222 (N_16222,N_8058,N_7054);
xor U16223 (N_16223,N_6375,N_6852);
xor U16224 (N_16224,N_9217,N_8289);
nand U16225 (N_16225,N_10199,N_6740);
nor U16226 (N_16226,N_9234,N_7392);
and U16227 (N_16227,N_10668,N_9390);
and U16228 (N_16228,N_8690,N_11258);
or U16229 (N_16229,N_8171,N_6951);
and U16230 (N_16230,N_10256,N_11802);
or U16231 (N_16231,N_6592,N_10612);
nor U16232 (N_16232,N_7684,N_8194);
nand U16233 (N_16233,N_7942,N_10492);
and U16234 (N_16234,N_7755,N_10580);
or U16235 (N_16235,N_10472,N_12048);
nand U16236 (N_16236,N_6776,N_9429);
or U16237 (N_16237,N_9227,N_10291);
and U16238 (N_16238,N_7207,N_8611);
nand U16239 (N_16239,N_8127,N_6998);
nand U16240 (N_16240,N_7591,N_11585);
or U16241 (N_16241,N_7401,N_10365);
nand U16242 (N_16242,N_11064,N_9369);
and U16243 (N_16243,N_9029,N_12439);
or U16244 (N_16244,N_9390,N_8997);
and U16245 (N_16245,N_11559,N_12348);
or U16246 (N_16246,N_12416,N_8979);
or U16247 (N_16247,N_9241,N_9780);
nor U16248 (N_16248,N_8308,N_6917);
xor U16249 (N_16249,N_9975,N_9184);
and U16250 (N_16250,N_7402,N_8233);
xnor U16251 (N_16251,N_10767,N_8040);
nor U16252 (N_16252,N_6433,N_10562);
or U16253 (N_16253,N_7280,N_10838);
and U16254 (N_16254,N_10249,N_7810);
nand U16255 (N_16255,N_11457,N_10031);
nor U16256 (N_16256,N_11621,N_9618);
nand U16257 (N_16257,N_10945,N_9727);
or U16258 (N_16258,N_9626,N_8017);
nand U16259 (N_16259,N_8491,N_9455);
nor U16260 (N_16260,N_12302,N_9547);
nand U16261 (N_16261,N_11155,N_8497);
and U16262 (N_16262,N_8518,N_11289);
and U16263 (N_16263,N_9266,N_12112);
and U16264 (N_16264,N_11829,N_9898);
and U16265 (N_16265,N_7713,N_11679);
or U16266 (N_16266,N_8701,N_7799);
nand U16267 (N_16267,N_12117,N_8061);
or U16268 (N_16268,N_6329,N_11971);
nand U16269 (N_16269,N_12454,N_9983);
nor U16270 (N_16270,N_9099,N_6420);
or U16271 (N_16271,N_7703,N_9371);
nand U16272 (N_16272,N_7174,N_12211);
and U16273 (N_16273,N_6317,N_8013);
or U16274 (N_16274,N_8460,N_9766);
and U16275 (N_16275,N_6534,N_8995);
or U16276 (N_16276,N_12336,N_8703);
xor U16277 (N_16277,N_9379,N_6605);
nand U16278 (N_16278,N_9518,N_6493);
and U16279 (N_16279,N_9486,N_7861);
nor U16280 (N_16280,N_9972,N_8575);
nand U16281 (N_16281,N_7911,N_12060);
nor U16282 (N_16282,N_7002,N_10232);
or U16283 (N_16283,N_9202,N_6452);
nand U16284 (N_16284,N_6453,N_11025);
and U16285 (N_16285,N_8273,N_6984);
or U16286 (N_16286,N_12129,N_7104);
or U16287 (N_16287,N_11877,N_11186);
or U16288 (N_16288,N_11158,N_12209);
nand U16289 (N_16289,N_9938,N_9939);
or U16290 (N_16290,N_7925,N_9886);
or U16291 (N_16291,N_8215,N_9009);
nor U16292 (N_16292,N_11436,N_11393);
and U16293 (N_16293,N_6846,N_7336);
and U16294 (N_16294,N_10614,N_9806);
and U16295 (N_16295,N_12134,N_11912);
or U16296 (N_16296,N_9519,N_11568);
nor U16297 (N_16297,N_8763,N_8277);
nor U16298 (N_16298,N_8233,N_9539);
and U16299 (N_16299,N_11599,N_11940);
and U16300 (N_16300,N_7568,N_8275);
or U16301 (N_16301,N_9171,N_7115);
nand U16302 (N_16302,N_7056,N_12069);
nand U16303 (N_16303,N_9135,N_8869);
nand U16304 (N_16304,N_11769,N_10213);
nor U16305 (N_16305,N_9321,N_11916);
and U16306 (N_16306,N_7636,N_10035);
nand U16307 (N_16307,N_11299,N_9363);
and U16308 (N_16308,N_7770,N_6263);
and U16309 (N_16309,N_10020,N_11640);
nor U16310 (N_16310,N_7784,N_7118);
nand U16311 (N_16311,N_9575,N_7343);
and U16312 (N_16312,N_8771,N_6620);
xor U16313 (N_16313,N_10432,N_8472);
nor U16314 (N_16314,N_6815,N_12413);
nor U16315 (N_16315,N_10108,N_6750);
nor U16316 (N_16316,N_10040,N_10251);
and U16317 (N_16317,N_6790,N_11889);
and U16318 (N_16318,N_7800,N_11327);
or U16319 (N_16319,N_7484,N_10349);
xor U16320 (N_16320,N_6545,N_7690);
and U16321 (N_16321,N_9261,N_8481);
and U16322 (N_16322,N_8027,N_11676);
nor U16323 (N_16323,N_11992,N_7538);
nand U16324 (N_16324,N_10771,N_6851);
xnor U16325 (N_16325,N_12110,N_8112);
xor U16326 (N_16326,N_9849,N_7655);
or U16327 (N_16327,N_7757,N_9790);
or U16328 (N_16328,N_8154,N_7307);
and U16329 (N_16329,N_11137,N_10738);
nand U16330 (N_16330,N_7922,N_9413);
and U16331 (N_16331,N_8842,N_7304);
nor U16332 (N_16332,N_11583,N_11890);
or U16333 (N_16333,N_8365,N_7379);
and U16334 (N_16334,N_10775,N_12117);
or U16335 (N_16335,N_10539,N_6368);
nor U16336 (N_16336,N_7546,N_7816);
or U16337 (N_16337,N_8450,N_10118);
nand U16338 (N_16338,N_8641,N_9389);
or U16339 (N_16339,N_11918,N_10692);
and U16340 (N_16340,N_9910,N_8956);
nand U16341 (N_16341,N_7811,N_9682);
nand U16342 (N_16342,N_7823,N_12010);
nand U16343 (N_16343,N_8422,N_9910);
or U16344 (N_16344,N_7218,N_9545);
nand U16345 (N_16345,N_10124,N_9650);
and U16346 (N_16346,N_8883,N_8920);
or U16347 (N_16347,N_8664,N_8778);
nand U16348 (N_16348,N_8672,N_7246);
nand U16349 (N_16349,N_9767,N_8364);
and U16350 (N_16350,N_10925,N_8786);
nand U16351 (N_16351,N_11159,N_12488);
nand U16352 (N_16352,N_9936,N_12263);
and U16353 (N_16353,N_6632,N_12061);
nand U16354 (N_16354,N_7839,N_6663);
or U16355 (N_16355,N_6970,N_7857);
and U16356 (N_16356,N_7279,N_8066);
xnor U16357 (N_16357,N_7934,N_6582);
nand U16358 (N_16358,N_7965,N_12128);
and U16359 (N_16359,N_6811,N_7061);
or U16360 (N_16360,N_7116,N_7710);
nor U16361 (N_16361,N_10737,N_12151);
nor U16362 (N_16362,N_12017,N_9162);
or U16363 (N_16363,N_6877,N_10346);
and U16364 (N_16364,N_7365,N_9350);
and U16365 (N_16365,N_8539,N_8563);
or U16366 (N_16366,N_8963,N_6925);
or U16367 (N_16367,N_10026,N_8675);
nor U16368 (N_16368,N_11305,N_7462);
or U16369 (N_16369,N_6542,N_11703);
nand U16370 (N_16370,N_12440,N_9314);
nor U16371 (N_16371,N_8350,N_7131);
xnor U16372 (N_16372,N_9652,N_6660);
or U16373 (N_16373,N_9709,N_7930);
nand U16374 (N_16374,N_11789,N_8713);
nor U16375 (N_16375,N_9551,N_10431);
and U16376 (N_16376,N_6913,N_9779);
and U16377 (N_16377,N_6882,N_8937);
or U16378 (N_16378,N_9157,N_7503);
or U16379 (N_16379,N_8366,N_8618);
and U16380 (N_16380,N_7449,N_7836);
nor U16381 (N_16381,N_9252,N_7862);
or U16382 (N_16382,N_6952,N_6833);
nand U16383 (N_16383,N_10936,N_8912);
and U16384 (N_16384,N_9345,N_12429);
nor U16385 (N_16385,N_9032,N_8788);
xnor U16386 (N_16386,N_8514,N_10324);
nor U16387 (N_16387,N_11015,N_11318);
or U16388 (N_16388,N_12206,N_10730);
nor U16389 (N_16389,N_7567,N_7463);
nand U16390 (N_16390,N_7467,N_6922);
nand U16391 (N_16391,N_11512,N_8970);
nand U16392 (N_16392,N_11870,N_7133);
xnor U16393 (N_16393,N_7431,N_8436);
nand U16394 (N_16394,N_7284,N_6330);
xnor U16395 (N_16395,N_9652,N_9150);
and U16396 (N_16396,N_7786,N_10140);
and U16397 (N_16397,N_8936,N_6730);
and U16398 (N_16398,N_11535,N_6486);
nand U16399 (N_16399,N_12233,N_9326);
nor U16400 (N_16400,N_7761,N_7013);
or U16401 (N_16401,N_9077,N_10938);
nor U16402 (N_16402,N_9048,N_12433);
or U16403 (N_16403,N_7307,N_11407);
nor U16404 (N_16404,N_6283,N_9917);
and U16405 (N_16405,N_11575,N_7396);
nand U16406 (N_16406,N_7416,N_7950);
and U16407 (N_16407,N_8480,N_9954);
xnor U16408 (N_16408,N_6366,N_10672);
or U16409 (N_16409,N_10019,N_7110);
or U16410 (N_16410,N_8778,N_7927);
or U16411 (N_16411,N_6328,N_11085);
or U16412 (N_16412,N_12479,N_11228);
and U16413 (N_16413,N_11311,N_9474);
xor U16414 (N_16414,N_10923,N_9299);
or U16415 (N_16415,N_12143,N_6669);
and U16416 (N_16416,N_9143,N_9417);
and U16417 (N_16417,N_7019,N_12412);
and U16418 (N_16418,N_12273,N_11257);
or U16419 (N_16419,N_8581,N_9817);
and U16420 (N_16420,N_9791,N_11135);
nand U16421 (N_16421,N_9771,N_8211);
nand U16422 (N_16422,N_8341,N_6749);
and U16423 (N_16423,N_8441,N_12310);
or U16424 (N_16424,N_10450,N_11047);
and U16425 (N_16425,N_6292,N_10764);
and U16426 (N_16426,N_12111,N_11706);
or U16427 (N_16427,N_7231,N_10739);
nor U16428 (N_16428,N_6348,N_11171);
nor U16429 (N_16429,N_9709,N_8253);
nand U16430 (N_16430,N_9395,N_8986);
nand U16431 (N_16431,N_11448,N_10633);
xor U16432 (N_16432,N_7531,N_11460);
nor U16433 (N_16433,N_9249,N_11345);
and U16434 (N_16434,N_7384,N_11066);
and U16435 (N_16435,N_10202,N_6927);
or U16436 (N_16436,N_9600,N_8982);
and U16437 (N_16437,N_9893,N_6846);
and U16438 (N_16438,N_10441,N_7939);
or U16439 (N_16439,N_11375,N_8830);
and U16440 (N_16440,N_8297,N_12339);
nor U16441 (N_16441,N_7417,N_8692);
xnor U16442 (N_16442,N_9257,N_8533);
and U16443 (N_16443,N_12273,N_8208);
nor U16444 (N_16444,N_11546,N_6544);
nand U16445 (N_16445,N_8880,N_7599);
or U16446 (N_16446,N_10966,N_8456);
nand U16447 (N_16447,N_9114,N_9933);
xnor U16448 (N_16448,N_9462,N_11164);
nand U16449 (N_16449,N_11811,N_8281);
or U16450 (N_16450,N_11473,N_9305);
nor U16451 (N_16451,N_7568,N_9115);
xnor U16452 (N_16452,N_11622,N_11100);
nor U16453 (N_16453,N_6521,N_9236);
or U16454 (N_16454,N_11877,N_12474);
nand U16455 (N_16455,N_8382,N_10709);
and U16456 (N_16456,N_12255,N_10075);
nand U16457 (N_16457,N_8652,N_12371);
and U16458 (N_16458,N_6932,N_7787);
nor U16459 (N_16459,N_9781,N_12170);
nor U16460 (N_16460,N_6370,N_8151);
and U16461 (N_16461,N_11937,N_10077);
or U16462 (N_16462,N_8465,N_7085);
nor U16463 (N_16463,N_6611,N_6484);
nand U16464 (N_16464,N_6941,N_9357);
nand U16465 (N_16465,N_9793,N_8574);
nand U16466 (N_16466,N_8061,N_7595);
xnor U16467 (N_16467,N_7352,N_6362);
and U16468 (N_16468,N_10779,N_6376);
nor U16469 (N_16469,N_10900,N_9768);
nor U16470 (N_16470,N_9035,N_7020);
nor U16471 (N_16471,N_6664,N_6715);
and U16472 (N_16472,N_6939,N_6325);
and U16473 (N_16473,N_9417,N_6356);
and U16474 (N_16474,N_8135,N_6481);
nand U16475 (N_16475,N_7672,N_9847);
and U16476 (N_16476,N_12298,N_10942);
nor U16477 (N_16477,N_9976,N_8349);
nor U16478 (N_16478,N_11411,N_8297);
xnor U16479 (N_16479,N_11320,N_10010);
or U16480 (N_16480,N_11713,N_8428);
or U16481 (N_16481,N_11422,N_8783);
and U16482 (N_16482,N_7594,N_7301);
or U16483 (N_16483,N_6908,N_11795);
nor U16484 (N_16484,N_6359,N_12156);
and U16485 (N_16485,N_8359,N_6885);
or U16486 (N_16486,N_9903,N_8016);
and U16487 (N_16487,N_8498,N_9254);
and U16488 (N_16488,N_10707,N_11160);
xor U16489 (N_16489,N_9438,N_7255);
and U16490 (N_16490,N_6610,N_8081);
and U16491 (N_16491,N_7329,N_7764);
nor U16492 (N_16492,N_10144,N_11581);
nor U16493 (N_16493,N_10652,N_8972);
nand U16494 (N_16494,N_7824,N_10220);
nor U16495 (N_16495,N_11952,N_11443);
or U16496 (N_16496,N_8256,N_8191);
and U16497 (N_16497,N_8371,N_11305);
and U16498 (N_16498,N_8040,N_10833);
and U16499 (N_16499,N_10039,N_12082);
nor U16500 (N_16500,N_7895,N_11050);
nor U16501 (N_16501,N_11059,N_7605);
or U16502 (N_16502,N_8489,N_8401);
and U16503 (N_16503,N_6455,N_7896);
nor U16504 (N_16504,N_11896,N_11127);
or U16505 (N_16505,N_7937,N_6288);
nor U16506 (N_16506,N_11185,N_7191);
nor U16507 (N_16507,N_6657,N_10079);
nor U16508 (N_16508,N_11650,N_10122);
or U16509 (N_16509,N_7842,N_7200);
or U16510 (N_16510,N_10752,N_11575);
nor U16511 (N_16511,N_11938,N_7454);
or U16512 (N_16512,N_10810,N_9136);
nor U16513 (N_16513,N_10494,N_9421);
xor U16514 (N_16514,N_11332,N_8766);
and U16515 (N_16515,N_8740,N_8951);
nor U16516 (N_16516,N_8459,N_8057);
xor U16517 (N_16517,N_9516,N_12433);
and U16518 (N_16518,N_6717,N_7374);
or U16519 (N_16519,N_7750,N_11752);
and U16520 (N_16520,N_6791,N_11944);
nand U16521 (N_16521,N_9074,N_7073);
nor U16522 (N_16522,N_11558,N_7170);
xnor U16523 (N_16523,N_8120,N_11282);
nor U16524 (N_16524,N_10903,N_6667);
nor U16525 (N_16525,N_9597,N_9755);
and U16526 (N_16526,N_11375,N_9960);
nand U16527 (N_16527,N_11351,N_6468);
and U16528 (N_16528,N_8754,N_11940);
nand U16529 (N_16529,N_11947,N_9998);
nand U16530 (N_16530,N_11623,N_7875);
or U16531 (N_16531,N_7180,N_11579);
and U16532 (N_16532,N_9779,N_8396);
nand U16533 (N_16533,N_10014,N_9572);
nand U16534 (N_16534,N_8087,N_6544);
and U16535 (N_16535,N_8896,N_7746);
xnor U16536 (N_16536,N_10957,N_11840);
or U16537 (N_16537,N_7438,N_7693);
nand U16538 (N_16538,N_9893,N_8392);
and U16539 (N_16539,N_6888,N_7962);
nand U16540 (N_16540,N_8357,N_9365);
or U16541 (N_16541,N_7304,N_7079);
and U16542 (N_16542,N_8770,N_8380);
nand U16543 (N_16543,N_9736,N_8952);
or U16544 (N_16544,N_8699,N_10695);
nand U16545 (N_16545,N_6888,N_8761);
nand U16546 (N_16546,N_10594,N_8724);
or U16547 (N_16547,N_10438,N_12334);
nand U16548 (N_16548,N_6647,N_10465);
or U16549 (N_16549,N_10546,N_6754);
nor U16550 (N_16550,N_12362,N_8080);
xor U16551 (N_16551,N_11870,N_11083);
or U16552 (N_16552,N_9850,N_9703);
and U16553 (N_16553,N_9887,N_7463);
and U16554 (N_16554,N_6306,N_11304);
or U16555 (N_16555,N_7621,N_10759);
nand U16556 (N_16556,N_11702,N_12278);
or U16557 (N_16557,N_6642,N_11489);
and U16558 (N_16558,N_10852,N_10077);
xnor U16559 (N_16559,N_9617,N_8007);
and U16560 (N_16560,N_7532,N_10047);
and U16561 (N_16561,N_10686,N_12293);
nand U16562 (N_16562,N_8472,N_12400);
or U16563 (N_16563,N_11892,N_9450);
nand U16564 (N_16564,N_8439,N_11096);
xnor U16565 (N_16565,N_12409,N_12360);
and U16566 (N_16566,N_8009,N_11713);
or U16567 (N_16567,N_7261,N_7863);
nand U16568 (N_16568,N_11134,N_10258);
nand U16569 (N_16569,N_11423,N_8324);
nand U16570 (N_16570,N_7425,N_11780);
or U16571 (N_16571,N_7139,N_9995);
and U16572 (N_16572,N_6701,N_8668);
nand U16573 (N_16573,N_7599,N_7247);
or U16574 (N_16574,N_7742,N_10416);
nand U16575 (N_16575,N_12177,N_7674);
or U16576 (N_16576,N_12451,N_6863);
nor U16577 (N_16577,N_10342,N_9904);
or U16578 (N_16578,N_7553,N_10975);
nor U16579 (N_16579,N_11026,N_7356);
nand U16580 (N_16580,N_8574,N_6757);
or U16581 (N_16581,N_12399,N_6680);
or U16582 (N_16582,N_8831,N_12075);
nor U16583 (N_16583,N_8768,N_12398);
and U16584 (N_16584,N_10587,N_11167);
xnor U16585 (N_16585,N_11432,N_9288);
nor U16586 (N_16586,N_10331,N_8407);
or U16587 (N_16587,N_12147,N_9702);
xnor U16588 (N_16588,N_11125,N_10982);
nor U16589 (N_16589,N_11692,N_6791);
nor U16590 (N_16590,N_8270,N_8260);
nor U16591 (N_16591,N_8554,N_9463);
or U16592 (N_16592,N_9486,N_12451);
and U16593 (N_16593,N_7224,N_8764);
nand U16594 (N_16594,N_11067,N_6495);
or U16595 (N_16595,N_7822,N_10695);
or U16596 (N_16596,N_10426,N_9248);
or U16597 (N_16597,N_10424,N_11386);
nand U16598 (N_16598,N_9358,N_7801);
nand U16599 (N_16599,N_7899,N_9654);
nand U16600 (N_16600,N_10665,N_12198);
xnor U16601 (N_16601,N_6552,N_7991);
nand U16602 (N_16602,N_11179,N_11298);
or U16603 (N_16603,N_6509,N_7942);
and U16604 (N_16604,N_7534,N_7622);
nor U16605 (N_16605,N_7813,N_9873);
xor U16606 (N_16606,N_6394,N_11925);
or U16607 (N_16607,N_9439,N_9039);
nand U16608 (N_16608,N_8519,N_7792);
and U16609 (N_16609,N_9533,N_10991);
or U16610 (N_16610,N_10293,N_6351);
xor U16611 (N_16611,N_10292,N_10484);
nor U16612 (N_16612,N_9890,N_10621);
or U16613 (N_16613,N_9558,N_7687);
and U16614 (N_16614,N_6770,N_8359);
nor U16615 (N_16615,N_6528,N_8079);
nor U16616 (N_16616,N_9900,N_8639);
or U16617 (N_16617,N_9067,N_10508);
xnor U16618 (N_16618,N_8876,N_7906);
and U16619 (N_16619,N_12213,N_10202);
or U16620 (N_16620,N_8836,N_9161);
or U16621 (N_16621,N_10572,N_6581);
or U16622 (N_16622,N_9135,N_12012);
nor U16623 (N_16623,N_11913,N_7305);
nand U16624 (N_16624,N_12098,N_6387);
and U16625 (N_16625,N_12224,N_8451);
and U16626 (N_16626,N_8324,N_7950);
nand U16627 (N_16627,N_10799,N_10861);
nand U16628 (N_16628,N_7916,N_7030);
or U16629 (N_16629,N_12195,N_12105);
and U16630 (N_16630,N_9638,N_10471);
and U16631 (N_16631,N_12269,N_11709);
or U16632 (N_16632,N_9822,N_10539);
xor U16633 (N_16633,N_6251,N_12038);
or U16634 (N_16634,N_6708,N_8260);
nand U16635 (N_16635,N_9070,N_6891);
nor U16636 (N_16636,N_11851,N_7304);
and U16637 (N_16637,N_12000,N_9543);
or U16638 (N_16638,N_11738,N_7161);
or U16639 (N_16639,N_10140,N_8058);
and U16640 (N_16640,N_11635,N_8657);
or U16641 (N_16641,N_7034,N_12360);
xor U16642 (N_16642,N_9892,N_10565);
and U16643 (N_16643,N_11962,N_9340);
or U16644 (N_16644,N_7462,N_6761);
and U16645 (N_16645,N_10716,N_7564);
nor U16646 (N_16646,N_7419,N_6360);
nand U16647 (N_16647,N_8750,N_12293);
and U16648 (N_16648,N_6318,N_7195);
or U16649 (N_16649,N_9257,N_8479);
or U16650 (N_16650,N_10537,N_7967);
xor U16651 (N_16651,N_11770,N_7413);
and U16652 (N_16652,N_11354,N_7304);
nor U16653 (N_16653,N_9755,N_9401);
and U16654 (N_16654,N_9309,N_8689);
nor U16655 (N_16655,N_11927,N_10882);
nand U16656 (N_16656,N_10733,N_9260);
and U16657 (N_16657,N_8759,N_11432);
or U16658 (N_16658,N_7052,N_7139);
nand U16659 (N_16659,N_12097,N_11317);
nand U16660 (N_16660,N_10263,N_9836);
or U16661 (N_16661,N_9573,N_9253);
nor U16662 (N_16662,N_9074,N_7424);
nand U16663 (N_16663,N_6558,N_8028);
nand U16664 (N_16664,N_9262,N_7623);
or U16665 (N_16665,N_7005,N_10265);
or U16666 (N_16666,N_11959,N_6367);
and U16667 (N_16667,N_9929,N_10075);
nor U16668 (N_16668,N_11646,N_6789);
and U16669 (N_16669,N_7175,N_6922);
nand U16670 (N_16670,N_7832,N_12255);
and U16671 (N_16671,N_10839,N_8201);
nor U16672 (N_16672,N_9291,N_10089);
nand U16673 (N_16673,N_6403,N_7478);
or U16674 (N_16674,N_10715,N_6959);
xnor U16675 (N_16675,N_10108,N_8821);
or U16676 (N_16676,N_7172,N_8926);
and U16677 (N_16677,N_11331,N_10374);
xor U16678 (N_16678,N_8751,N_10430);
or U16679 (N_16679,N_11808,N_7930);
nor U16680 (N_16680,N_8480,N_9252);
or U16681 (N_16681,N_6605,N_6731);
nor U16682 (N_16682,N_12444,N_9267);
nor U16683 (N_16683,N_11744,N_9344);
nand U16684 (N_16684,N_6560,N_10836);
xor U16685 (N_16685,N_11307,N_11007);
and U16686 (N_16686,N_6267,N_7969);
nor U16687 (N_16687,N_12042,N_6823);
or U16688 (N_16688,N_8330,N_6880);
or U16689 (N_16689,N_10529,N_9171);
or U16690 (N_16690,N_6932,N_10993);
and U16691 (N_16691,N_8054,N_7891);
nor U16692 (N_16692,N_9751,N_10453);
nor U16693 (N_16693,N_8323,N_8224);
nor U16694 (N_16694,N_9912,N_9803);
nor U16695 (N_16695,N_7954,N_6717);
or U16696 (N_16696,N_10023,N_10885);
nand U16697 (N_16697,N_9451,N_12296);
or U16698 (N_16698,N_12202,N_9488);
or U16699 (N_16699,N_7707,N_8646);
nor U16700 (N_16700,N_7166,N_7927);
nand U16701 (N_16701,N_9405,N_7778);
or U16702 (N_16702,N_10582,N_8466);
nor U16703 (N_16703,N_9181,N_9152);
nand U16704 (N_16704,N_9710,N_9440);
and U16705 (N_16705,N_10357,N_8421);
or U16706 (N_16706,N_9178,N_9985);
and U16707 (N_16707,N_10896,N_8203);
or U16708 (N_16708,N_8712,N_9490);
xnor U16709 (N_16709,N_10413,N_8485);
and U16710 (N_16710,N_9602,N_9090);
nor U16711 (N_16711,N_11806,N_6654);
nor U16712 (N_16712,N_8541,N_10366);
nand U16713 (N_16713,N_11865,N_7637);
nor U16714 (N_16714,N_10877,N_7335);
xor U16715 (N_16715,N_11936,N_8326);
nand U16716 (N_16716,N_11997,N_7345);
or U16717 (N_16717,N_10903,N_9055);
or U16718 (N_16718,N_11822,N_10804);
nor U16719 (N_16719,N_7495,N_8319);
nand U16720 (N_16720,N_8146,N_7671);
nor U16721 (N_16721,N_10111,N_8184);
or U16722 (N_16722,N_7438,N_11495);
or U16723 (N_16723,N_9305,N_7081);
and U16724 (N_16724,N_6545,N_8155);
and U16725 (N_16725,N_9090,N_8836);
or U16726 (N_16726,N_9922,N_10117);
or U16727 (N_16727,N_8611,N_7438);
and U16728 (N_16728,N_8985,N_9663);
nand U16729 (N_16729,N_7372,N_11129);
and U16730 (N_16730,N_6640,N_8010);
nand U16731 (N_16731,N_10274,N_10934);
and U16732 (N_16732,N_11038,N_8476);
nand U16733 (N_16733,N_9221,N_7523);
xor U16734 (N_16734,N_7666,N_8210);
or U16735 (N_16735,N_9068,N_10714);
nand U16736 (N_16736,N_11246,N_8893);
nor U16737 (N_16737,N_7103,N_9293);
and U16738 (N_16738,N_11241,N_7311);
or U16739 (N_16739,N_12346,N_9674);
xnor U16740 (N_16740,N_11974,N_10097);
nor U16741 (N_16741,N_11036,N_9289);
or U16742 (N_16742,N_10292,N_10127);
nand U16743 (N_16743,N_8758,N_10733);
nand U16744 (N_16744,N_12003,N_11997);
nand U16745 (N_16745,N_11213,N_12057);
nor U16746 (N_16746,N_11563,N_9970);
or U16747 (N_16747,N_12093,N_12401);
nor U16748 (N_16748,N_9540,N_6911);
and U16749 (N_16749,N_6586,N_10266);
nor U16750 (N_16750,N_6557,N_6562);
and U16751 (N_16751,N_10910,N_7197);
and U16752 (N_16752,N_7403,N_7339);
and U16753 (N_16753,N_8835,N_8432);
and U16754 (N_16754,N_7582,N_8385);
or U16755 (N_16755,N_7318,N_7811);
nor U16756 (N_16756,N_7733,N_9974);
nand U16757 (N_16757,N_10646,N_11690);
xor U16758 (N_16758,N_6370,N_7353);
xnor U16759 (N_16759,N_9419,N_6937);
nand U16760 (N_16760,N_7852,N_10477);
xor U16761 (N_16761,N_9359,N_9495);
nor U16762 (N_16762,N_7405,N_9161);
or U16763 (N_16763,N_9103,N_11193);
nand U16764 (N_16764,N_7687,N_8592);
or U16765 (N_16765,N_8288,N_10163);
and U16766 (N_16766,N_12167,N_9283);
nand U16767 (N_16767,N_7187,N_12263);
xnor U16768 (N_16768,N_9191,N_8741);
nand U16769 (N_16769,N_8548,N_9408);
nor U16770 (N_16770,N_12453,N_10836);
nor U16771 (N_16771,N_12243,N_12489);
nor U16772 (N_16772,N_9258,N_9116);
xor U16773 (N_16773,N_7037,N_6812);
xor U16774 (N_16774,N_11188,N_10580);
nor U16775 (N_16775,N_9726,N_6606);
and U16776 (N_16776,N_6736,N_12385);
or U16777 (N_16777,N_10744,N_6637);
or U16778 (N_16778,N_10553,N_11391);
or U16779 (N_16779,N_10064,N_9920);
or U16780 (N_16780,N_6863,N_9633);
nand U16781 (N_16781,N_6888,N_11415);
and U16782 (N_16782,N_7761,N_10239);
and U16783 (N_16783,N_7529,N_11534);
and U16784 (N_16784,N_8921,N_10521);
or U16785 (N_16785,N_7858,N_7162);
nor U16786 (N_16786,N_7702,N_11891);
or U16787 (N_16787,N_11422,N_7210);
nor U16788 (N_16788,N_6313,N_11498);
or U16789 (N_16789,N_10553,N_10574);
nor U16790 (N_16790,N_8523,N_9850);
or U16791 (N_16791,N_10089,N_8208);
nor U16792 (N_16792,N_11074,N_10330);
xnor U16793 (N_16793,N_10196,N_9592);
or U16794 (N_16794,N_11318,N_8229);
nor U16795 (N_16795,N_9754,N_10684);
nand U16796 (N_16796,N_10068,N_11693);
or U16797 (N_16797,N_10485,N_11729);
or U16798 (N_16798,N_6376,N_11016);
and U16799 (N_16799,N_7465,N_7990);
nand U16800 (N_16800,N_7280,N_8069);
nand U16801 (N_16801,N_6339,N_10078);
nand U16802 (N_16802,N_6914,N_12150);
and U16803 (N_16803,N_8056,N_8240);
or U16804 (N_16804,N_10061,N_11511);
nor U16805 (N_16805,N_6391,N_6513);
and U16806 (N_16806,N_11901,N_6931);
nor U16807 (N_16807,N_8894,N_8568);
xor U16808 (N_16808,N_8738,N_11357);
and U16809 (N_16809,N_11971,N_8172);
or U16810 (N_16810,N_6251,N_10626);
and U16811 (N_16811,N_10513,N_9857);
or U16812 (N_16812,N_8574,N_8880);
and U16813 (N_16813,N_7918,N_9353);
or U16814 (N_16814,N_9032,N_10614);
or U16815 (N_16815,N_8165,N_10611);
xnor U16816 (N_16816,N_6762,N_8704);
or U16817 (N_16817,N_7834,N_10887);
or U16818 (N_16818,N_6255,N_9503);
nor U16819 (N_16819,N_9110,N_10773);
nor U16820 (N_16820,N_11490,N_9368);
nand U16821 (N_16821,N_8572,N_11112);
or U16822 (N_16822,N_11691,N_9846);
and U16823 (N_16823,N_10031,N_9532);
and U16824 (N_16824,N_9781,N_10393);
nand U16825 (N_16825,N_6650,N_9604);
nand U16826 (N_16826,N_10213,N_8766);
and U16827 (N_16827,N_11585,N_9564);
nand U16828 (N_16828,N_12493,N_11963);
and U16829 (N_16829,N_8895,N_8820);
nand U16830 (N_16830,N_9210,N_9148);
or U16831 (N_16831,N_11560,N_10912);
and U16832 (N_16832,N_9792,N_10483);
nor U16833 (N_16833,N_9626,N_11108);
and U16834 (N_16834,N_7467,N_6589);
and U16835 (N_16835,N_7407,N_6659);
xnor U16836 (N_16836,N_9884,N_11748);
nor U16837 (N_16837,N_10064,N_7520);
or U16838 (N_16838,N_7852,N_6552);
nor U16839 (N_16839,N_6544,N_7266);
xor U16840 (N_16840,N_9442,N_6646);
nor U16841 (N_16841,N_8664,N_9550);
nor U16842 (N_16842,N_11200,N_11283);
and U16843 (N_16843,N_7394,N_8800);
and U16844 (N_16844,N_12020,N_9283);
or U16845 (N_16845,N_10774,N_6652);
and U16846 (N_16846,N_7725,N_11095);
or U16847 (N_16847,N_9880,N_11486);
nand U16848 (N_16848,N_11440,N_7701);
and U16849 (N_16849,N_10407,N_11136);
and U16850 (N_16850,N_9632,N_10298);
or U16851 (N_16851,N_8617,N_8074);
xor U16852 (N_16852,N_7937,N_10231);
xnor U16853 (N_16853,N_10522,N_11715);
nor U16854 (N_16854,N_10499,N_6733);
and U16855 (N_16855,N_11191,N_9655);
and U16856 (N_16856,N_10331,N_7713);
nand U16857 (N_16857,N_11228,N_7008);
nand U16858 (N_16858,N_9239,N_10059);
or U16859 (N_16859,N_11439,N_7817);
and U16860 (N_16860,N_12153,N_6950);
nand U16861 (N_16861,N_10864,N_9577);
nor U16862 (N_16862,N_9924,N_6539);
nand U16863 (N_16863,N_7200,N_7847);
xor U16864 (N_16864,N_11839,N_10676);
nand U16865 (N_16865,N_11627,N_7750);
nand U16866 (N_16866,N_6613,N_7231);
or U16867 (N_16867,N_6566,N_9983);
or U16868 (N_16868,N_8196,N_6925);
nor U16869 (N_16869,N_7427,N_7066);
nor U16870 (N_16870,N_8567,N_8139);
and U16871 (N_16871,N_8618,N_9074);
xnor U16872 (N_16872,N_6829,N_9594);
or U16873 (N_16873,N_9594,N_11448);
nor U16874 (N_16874,N_11346,N_9817);
or U16875 (N_16875,N_10920,N_7317);
nand U16876 (N_16876,N_7674,N_10583);
nand U16877 (N_16877,N_10219,N_9347);
nor U16878 (N_16878,N_10442,N_9994);
nor U16879 (N_16879,N_9543,N_8669);
nor U16880 (N_16880,N_11557,N_7166);
nor U16881 (N_16881,N_11756,N_7423);
nand U16882 (N_16882,N_10949,N_7378);
nor U16883 (N_16883,N_9596,N_11156);
or U16884 (N_16884,N_9524,N_10012);
and U16885 (N_16885,N_10504,N_10371);
and U16886 (N_16886,N_8993,N_6974);
xor U16887 (N_16887,N_10499,N_9753);
and U16888 (N_16888,N_6938,N_10864);
or U16889 (N_16889,N_7105,N_8291);
nor U16890 (N_16890,N_6349,N_8019);
nor U16891 (N_16891,N_7723,N_6641);
or U16892 (N_16892,N_11505,N_8876);
nor U16893 (N_16893,N_10314,N_9538);
nor U16894 (N_16894,N_12448,N_10183);
and U16895 (N_16895,N_11654,N_6800);
or U16896 (N_16896,N_11750,N_6559);
nor U16897 (N_16897,N_9714,N_7370);
nand U16898 (N_16898,N_8622,N_9840);
nor U16899 (N_16899,N_8824,N_10770);
and U16900 (N_16900,N_8745,N_10434);
nand U16901 (N_16901,N_9644,N_8730);
nand U16902 (N_16902,N_10558,N_6275);
nand U16903 (N_16903,N_12096,N_11173);
nand U16904 (N_16904,N_11845,N_6515);
nand U16905 (N_16905,N_10724,N_11132);
xnor U16906 (N_16906,N_8913,N_6625);
xnor U16907 (N_16907,N_10749,N_9644);
or U16908 (N_16908,N_11547,N_11003);
or U16909 (N_16909,N_10812,N_6960);
nand U16910 (N_16910,N_6270,N_7365);
and U16911 (N_16911,N_9067,N_8830);
nand U16912 (N_16912,N_10957,N_8698);
nand U16913 (N_16913,N_6764,N_10024);
nand U16914 (N_16914,N_9320,N_8113);
nand U16915 (N_16915,N_9413,N_8179);
and U16916 (N_16916,N_10870,N_11751);
and U16917 (N_16917,N_8587,N_7369);
nor U16918 (N_16918,N_8284,N_11964);
nor U16919 (N_16919,N_6889,N_7757);
nor U16920 (N_16920,N_11534,N_6517);
or U16921 (N_16921,N_11047,N_10487);
or U16922 (N_16922,N_8469,N_11527);
nand U16923 (N_16923,N_7990,N_6539);
xnor U16924 (N_16924,N_8061,N_10819);
and U16925 (N_16925,N_10558,N_8267);
or U16926 (N_16926,N_9894,N_8887);
and U16927 (N_16927,N_8206,N_11348);
xor U16928 (N_16928,N_10705,N_6365);
and U16929 (N_16929,N_10191,N_11989);
and U16930 (N_16930,N_11084,N_8388);
nor U16931 (N_16931,N_9801,N_8717);
nand U16932 (N_16932,N_6503,N_12264);
nor U16933 (N_16933,N_9533,N_10855);
nor U16934 (N_16934,N_9659,N_12397);
and U16935 (N_16935,N_10826,N_8828);
nor U16936 (N_16936,N_7166,N_9077);
nor U16937 (N_16937,N_7979,N_8725);
nand U16938 (N_16938,N_10596,N_8278);
nor U16939 (N_16939,N_7809,N_7657);
xnor U16940 (N_16940,N_7536,N_11014);
nand U16941 (N_16941,N_8840,N_7602);
or U16942 (N_16942,N_8406,N_9407);
and U16943 (N_16943,N_11434,N_10352);
and U16944 (N_16944,N_7538,N_6895);
nor U16945 (N_16945,N_12182,N_6780);
and U16946 (N_16946,N_7591,N_8737);
or U16947 (N_16947,N_9175,N_9024);
or U16948 (N_16948,N_12237,N_8253);
and U16949 (N_16949,N_7737,N_8583);
xor U16950 (N_16950,N_8154,N_11581);
nand U16951 (N_16951,N_6781,N_7835);
and U16952 (N_16952,N_6619,N_7066);
or U16953 (N_16953,N_7652,N_7390);
nor U16954 (N_16954,N_6979,N_11133);
nand U16955 (N_16955,N_11730,N_7828);
or U16956 (N_16956,N_9883,N_7581);
nor U16957 (N_16957,N_12414,N_7131);
nand U16958 (N_16958,N_7940,N_10496);
or U16959 (N_16959,N_9946,N_8734);
and U16960 (N_16960,N_10012,N_10208);
or U16961 (N_16961,N_12061,N_7581);
nand U16962 (N_16962,N_10414,N_12299);
or U16963 (N_16963,N_7386,N_9976);
nor U16964 (N_16964,N_9067,N_12402);
nand U16965 (N_16965,N_8913,N_9531);
or U16966 (N_16966,N_9909,N_8161);
or U16967 (N_16967,N_11746,N_10012);
or U16968 (N_16968,N_7070,N_10193);
nand U16969 (N_16969,N_9076,N_8040);
and U16970 (N_16970,N_7041,N_7557);
nand U16971 (N_16971,N_11362,N_8706);
nand U16972 (N_16972,N_7350,N_10964);
nand U16973 (N_16973,N_11282,N_9886);
nand U16974 (N_16974,N_7391,N_9002);
nor U16975 (N_16975,N_8745,N_10116);
or U16976 (N_16976,N_11607,N_9900);
or U16977 (N_16977,N_10385,N_7695);
and U16978 (N_16978,N_7745,N_10352);
nand U16979 (N_16979,N_11944,N_10320);
and U16980 (N_16980,N_7667,N_7294);
xnor U16981 (N_16981,N_11489,N_8940);
nor U16982 (N_16982,N_12370,N_9300);
or U16983 (N_16983,N_6375,N_10851);
nor U16984 (N_16984,N_12226,N_8520);
and U16985 (N_16985,N_6414,N_8394);
nand U16986 (N_16986,N_7618,N_12481);
or U16987 (N_16987,N_7851,N_6549);
and U16988 (N_16988,N_11309,N_7091);
nand U16989 (N_16989,N_10746,N_8720);
or U16990 (N_16990,N_11393,N_11256);
and U16991 (N_16991,N_10535,N_8123);
nand U16992 (N_16992,N_6723,N_8400);
nor U16993 (N_16993,N_8224,N_11847);
nand U16994 (N_16994,N_7070,N_8799);
nand U16995 (N_16995,N_7411,N_6986);
and U16996 (N_16996,N_7607,N_12466);
nand U16997 (N_16997,N_10487,N_8620);
or U16998 (N_16998,N_10116,N_7391);
or U16999 (N_16999,N_10219,N_7531);
nor U17000 (N_17000,N_9071,N_12014);
and U17001 (N_17001,N_9165,N_8228);
or U17002 (N_17002,N_10790,N_8083);
and U17003 (N_17003,N_8001,N_8271);
nor U17004 (N_17004,N_11969,N_10052);
or U17005 (N_17005,N_9759,N_12360);
nand U17006 (N_17006,N_7099,N_8018);
nand U17007 (N_17007,N_9141,N_7131);
nand U17008 (N_17008,N_9150,N_12390);
nand U17009 (N_17009,N_11704,N_11907);
or U17010 (N_17010,N_9867,N_10584);
and U17011 (N_17011,N_10057,N_7152);
or U17012 (N_17012,N_11264,N_10995);
xor U17013 (N_17013,N_10168,N_6630);
nand U17014 (N_17014,N_12022,N_7110);
nor U17015 (N_17015,N_6588,N_10480);
xor U17016 (N_17016,N_7415,N_10326);
nand U17017 (N_17017,N_9945,N_11443);
nor U17018 (N_17018,N_12177,N_10323);
xor U17019 (N_17019,N_8391,N_11976);
or U17020 (N_17020,N_12196,N_9338);
and U17021 (N_17021,N_9237,N_10333);
nand U17022 (N_17022,N_6702,N_11683);
and U17023 (N_17023,N_7699,N_7442);
and U17024 (N_17024,N_8281,N_10517);
and U17025 (N_17025,N_6766,N_9502);
or U17026 (N_17026,N_6979,N_6353);
nor U17027 (N_17027,N_7683,N_6271);
and U17028 (N_17028,N_12021,N_8662);
or U17029 (N_17029,N_11112,N_11472);
nor U17030 (N_17030,N_10885,N_7007);
nand U17031 (N_17031,N_9590,N_7100);
and U17032 (N_17032,N_7900,N_9721);
or U17033 (N_17033,N_6323,N_10806);
nand U17034 (N_17034,N_6600,N_9786);
nor U17035 (N_17035,N_11595,N_10504);
nor U17036 (N_17036,N_10849,N_7282);
nand U17037 (N_17037,N_10564,N_6859);
nand U17038 (N_17038,N_10610,N_11681);
nor U17039 (N_17039,N_8327,N_7751);
nand U17040 (N_17040,N_9711,N_12163);
or U17041 (N_17041,N_9496,N_9795);
nand U17042 (N_17042,N_7397,N_8894);
nand U17043 (N_17043,N_8795,N_8341);
nor U17044 (N_17044,N_11797,N_11141);
nand U17045 (N_17045,N_12394,N_10577);
and U17046 (N_17046,N_10256,N_8065);
nor U17047 (N_17047,N_12121,N_9489);
nand U17048 (N_17048,N_11418,N_6984);
nor U17049 (N_17049,N_10940,N_6269);
or U17050 (N_17050,N_11621,N_8886);
nand U17051 (N_17051,N_9106,N_12387);
and U17052 (N_17052,N_8569,N_9984);
nand U17053 (N_17053,N_11481,N_6840);
nor U17054 (N_17054,N_12287,N_7982);
and U17055 (N_17055,N_11763,N_11136);
and U17056 (N_17056,N_6450,N_9333);
and U17057 (N_17057,N_10679,N_8587);
nor U17058 (N_17058,N_12339,N_8055);
xor U17059 (N_17059,N_11856,N_9142);
nor U17060 (N_17060,N_9846,N_9571);
and U17061 (N_17061,N_7182,N_6675);
nand U17062 (N_17062,N_9162,N_9576);
xnor U17063 (N_17063,N_10358,N_11464);
nor U17064 (N_17064,N_12332,N_9305);
nand U17065 (N_17065,N_8615,N_10074);
xor U17066 (N_17066,N_9471,N_7585);
and U17067 (N_17067,N_7217,N_11162);
or U17068 (N_17068,N_9208,N_10093);
and U17069 (N_17069,N_7606,N_8333);
xor U17070 (N_17070,N_9329,N_7964);
nand U17071 (N_17071,N_8887,N_9983);
and U17072 (N_17072,N_9337,N_9799);
or U17073 (N_17073,N_10993,N_12064);
and U17074 (N_17074,N_8790,N_12099);
nand U17075 (N_17075,N_7680,N_7633);
and U17076 (N_17076,N_9190,N_10453);
nor U17077 (N_17077,N_6442,N_9493);
or U17078 (N_17078,N_8765,N_10653);
nor U17079 (N_17079,N_7207,N_7343);
nor U17080 (N_17080,N_12056,N_10580);
nor U17081 (N_17081,N_7233,N_10795);
or U17082 (N_17082,N_10815,N_11736);
or U17083 (N_17083,N_11628,N_9520);
nor U17084 (N_17084,N_8481,N_11166);
nand U17085 (N_17085,N_12098,N_11918);
xnor U17086 (N_17086,N_7625,N_6853);
nand U17087 (N_17087,N_7322,N_11928);
or U17088 (N_17088,N_12485,N_6594);
nand U17089 (N_17089,N_11277,N_12180);
or U17090 (N_17090,N_10008,N_10401);
or U17091 (N_17091,N_9903,N_10619);
nand U17092 (N_17092,N_10973,N_6778);
or U17093 (N_17093,N_8673,N_10606);
and U17094 (N_17094,N_8009,N_10230);
and U17095 (N_17095,N_11959,N_9779);
nand U17096 (N_17096,N_11183,N_6853);
nor U17097 (N_17097,N_7279,N_11916);
and U17098 (N_17098,N_11458,N_11541);
or U17099 (N_17099,N_9984,N_11605);
nand U17100 (N_17100,N_12395,N_8755);
nor U17101 (N_17101,N_8805,N_8204);
or U17102 (N_17102,N_7875,N_7961);
and U17103 (N_17103,N_11111,N_8521);
nand U17104 (N_17104,N_8054,N_11277);
and U17105 (N_17105,N_7858,N_7428);
or U17106 (N_17106,N_12486,N_10680);
nor U17107 (N_17107,N_8647,N_8951);
and U17108 (N_17108,N_9922,N_8630);
or U17109 (N_17109,N_8596,N_11476);
and U17110 (N_17110,N_6375,N_7179);
nor U17111 (N_17111,N_10479,N_12423);
nand U17112 (N_17112,N_11141,N_8871);
and U17113 (N_17113,N_6398,N_11597);
xnor U17114 (N_17114,N_11906,N_8178);
and U17115 (N_17115,N_8494,N_7014);
nor U17116 (N_17116,N_6865,N_10097);
and U17117 (N_17117,N_9365,N_10537);
xnor U17118 (N_17118,N_6308,N_6719);
and U17119 (N_17119,N_11251,N_8989);
and U17120 (N_17120,N_10514,N_6399);
nand U17121 (N_17121,N_10716,N_9186);
and U17122 (N_17122,N_8815,N_8531);
nor U17123 (N_17123,N_7457,N_11205);
or U17124 (N_17124,N_9060,N_9572);
xor U17125 (N_17125,N_7141,N_12062);
nor U17126 (N_17126,N_7319,N_9811);
nor U17127 (N_17127,N_7818,N_11352);
nand U17128 (N_17128,N_11889,N_10992);
nand U17129 (N_17129,N_7258,N_9972);
nand U17130 (N_17130,N_11978,N_12289);
and U17131 (N_17131,N_10258,N_7656);
xor U17132 (N_17132,N_12343,N_10351);
and U17133 (N_17133,N_7365,N_9243);
or U17134 (N_17134,N_6292,N_10361);
or U17135 (N_17135,N_8413,N_10372);
or U17136 (N_17136,N_10039,N_10432);
and U17137 (N_17137,N_9735,N_11321);
or U17138 (N_17138,N_9501,N_8834);
and U17139 (N_17139,N_7930,N_11856);
nand U17140 (N_17140,N_7203,N_8131);
or U17141 (N_17141,N_11412,N_6257);
nor U17142 (N_17142,N_6325,N_12474);
nor U17143 (N_17143,N_10001,N_8504);
and U17144 (N_17144,N_8716,N_8725);
nor U17145 (N_17145,N_11248,N_12465);
or U17146 (N_17146,N_7243,N_10286);
and U17147 (N_17147,N_6746,N_11865);
xnor U17148 (N_17148,N_7049,N_7211);
nor U17149 (N_17149,N_10435,N_10289);
or U17150 (N_17150,N_9495,N_6488);
or U17151 (N_17151,N_10871,N_6580);
or U17152 (N_17152,N_9095,N_8556);
xnor U17153 (N_17153,N_11100,N_9304);
xnor U17154 (N_17154,N_9823,N_7529);
nand U17155 (N_17155,N_12116,N_10918);
and U17156 (N_17156,N_9574,N_10482);
nor U17157 (N_17157,N_11010,N_10243);
nand U17158 (N_17158,N_8589,N_10625);
and U17159 (N_17159,N_9737,N_11415);
or U17160 (N_17160,N_7586,N_7443);
xnor U17161 (N_17161,N_9789,N_10110);
or U17162 (N_17162,N_9480,N_11526);
or U17163 (N_17163,N_10177,N_6419);
or U17164 (N_17164,N_8354,N_10299);
and U17165 (N_17165,N_6537,N_9083);
or U17166 (N_17166,N_8565,N_11291);
or U17167 (N_17167,N_11106,N_11815);
nand U17168 (N_17168,N_9701,N_9086);
nor U17169 (N_17169,N_7848,N_11852);
xnor U17170 (N_17170,N_7976,N_6794);
xor U17171 (N_17171,N_9543,N_12168);
and U17172 (N_17172,N_12020,N_7095);
or U17173 (N_17173,N_12067,N_6644);
and U17174 (N_17174,N_12239,N_11565);
nand U17175 (N_17175,N_12110,N_9927);
or U17176 (N_17176,N_10036,N_9414);
or U17177 (N_17177,N_6863,N_6779);
nand U17178 (N_17178,N_7237,N_8411);
nor U17179 (N_17179,N_11810,N_9403);
and U17180 (N_17180,N_10499,N_9531);
or U17181 (N_17181,N_8238,N_10407);
or U17182 (N_17182,N_11417,N_8742);
or U17183 (N_17183,N_9984,N_9545);
and U17184 (N_17184,N_6762,N_8388);
nor U17185 (N_17185,N_10394,N_7557);
nor U17186 (N_17186,N_10130,N_11952);
nand U17187 (N_17187,N_6431,N_12328);
or U17188 (N_17188,N_7838,N_7315);
nor U17189 (N_17189,N_9396,N_8373);
nor U17190 (N_17190,N_11637,N_9119);
and U17191 (N_17191,N_7286,N_11869);
or U17192 (N_17192,N_8950,N_8016);
and U17193 (N_17193,N_8996,N_11974);
nand U17194 (N_17194,N_6851,N_6524);
nand U17195 (N_17195,N_10706,N_9169);
xnor U17196 (N_17196,N_12145,N_10175);
and U17197 (N_17197,N_10924,N_10060);
or U17198 (N_17198,N_10423,N_10130);
and U17199 (N_17199,N_10889,N_10559);
or U17200 (N_17200,N_9201,N_8149);
or U17201 (N_17201,N_7280,N_9326);
and U17202 (N_17202,N_9585,N_10627);
nor U17203 (N_17203,N_7077,N_12475);
and U17204 (N_17204,N_11848,N_12388);
xnor U17205 (N_17205,N_7933,N_12329);
nor U17206 (N_17206,N_11339,N_10988);
and U17207 (N_17207,N_12289,N_11010);
or U17208 (N_17208,N_8840,N_8219);
and U17209 (N_17209,N_11654,N_8877);
nor U17210 (N_17210,N_8219,N_11439);
nor U17211 (N_17211,N_9520,N_6393);
nand U17212 (N_17212,N_11657,N_9922);
xor U17213 (N_17213,N_11742,N_11498);
nand U17214 (N_17214,N_11743,N_6635);
nand U17215 (N_17215,N_10143,N_8701);
nand U17216 (N_17216,N_8614,N_8445);
nor U17217 (N_17217,N_9271,N_6651);
and U17218 (N_17218,N_9897,N_6343);
nand U17219 (N_17219,N_8583,N_12177);
nor U17220 (N_17220,N_7882,N_7625);
xnor U17221 (N_17221,N_10631,N_9254);
nand U17222 (N_17222,N_6868,N_11855);
or U17223 (N_17223,N_9600,N_9476);
nand U17224 (N_17224,N_8273,N_10595);
xnor U17225 (N_17225,N_11706,N_10683);
xnor U17226 (N_17226,N_8070,N_7337);
nor U17227 (N_17227,N_8588,N_6372);
nand U17228 (N_17228,N_9724,N_12041);
and U17229 (N_17229,N_10541,N_11783);
or U17230 (N_17230,N_8581,N_6348);
or U17231 (N_17231,N_7518,N_10907);
or U17232 (N_17232,N_9503,N_8487);
nand U17233 (N_17233,N_10687,N_11086);
nor U17234 (N_17234,N_10871,N_6342);
and U17235 (N_17235,N_12339,N_7824);
xor U17236 (N_17236,N_8031,N_11331);
nand U17237 (N_17237,N_8166,N_11059);
xnor U17238 (N_17238,N_9745,N_7354);
nor U17239 (N_17239,N_7565,N_7867);
and U17240 (N_17240,N_11471,N_9336);
or U17241 (N_17241,N_9436,N_7290);
nor U17242 (N_17242,N_8527,N_8538);
or U17243 (N_17243,N_9438,N_8791);
or U17244 (N_17244,N_10019,N_8540);
and U17245 (N_17245,N_12035,N_10823);
and U17246 (N_17246,N_8788,N_9591);
and U17247 (N_17247,N_9802,N_6878);
xor U17248 (N_17248,N_7170,N_11345);
nor U17249 (N_17249,N_12056,N_12307);
xnor U17250 (N_17250,N_7284,N_9729);
nor U17251 (N_17251,N_11187,N_8879);
nor U17252 (N_17252,N_10537,N_9134);
or U17253 (N_17253,N_11532,N_6679);
xnor U17254 (N_17254,N_6638,N_8244);
nand U17255 (N_17255,N_10551,N_10933);
nand U17256 (N_17256,N_8628,N_11430);
nand U17257 (N_17257,N_12175,N_9955);
nand U17258 (N_17258,N_10916,N_7207);
xnor U17259 (N_17259,N_11453,N_10743);
xor U17260 (N_17260,N_8129,N_8813);
and U17261 (N_17261,N_11905,N_11038);
nand U17262 (N_17262,N_10044,N_10102);
or U17263 (N_17263,N_7440,N_9673);
and U17264 (N_17264,N_8467,N_10069);
nand U17265 (N_17265,N_11323,N_9875);
and U17266 (N_17266,N_8659,N_7216);
and U17267 (N_17267,N_9505,N_10545);
nand U17268 (N_17268,N_11907,N_10767);
nand U17269 (N_17269,N_10258,N_11374);
nor U17270 (N_17270,N_6395,N_9864);
or U17271 (N_17271,N_6442,N_7119);
xor U17272 (N_17272,N_9559,N_11892);
and U17273 (N_17273,N_8937,N_8535);
and U17274 (N_17274,N_12003,N_9524);
or U17275 (N_17275,N_12082,N_10386);
xnor U17276 (N_17276,N_9465,N_9084);
and U17277 (N_17277,N_9191,N_6533);
or U17278 (N_17278,N_9540,N_12199);
or U17279 (N_17279,N_9269,N_6300);
or U17280 (N_17280,N_8970,N_8641);
or U17281 (N_17281,N_8080,N_8143);
and U17282 (N_17282,N_7489,N_6875);
or U17283 (N_17283,N_12486,N_7324);
xor U17284 (N_17284,N_11782,N_8818);
or U17285 (N_17285,N_8171,N_9424);
nand U17286 (N_17286,N_9630,N_11391);
or U17287 (N_17287,N_9021,N_8724);
and U17288 (N_17288,N_8501,N_8438);
xnor U17289 (N_17289,N_6926,N_10545);
nor U17290 (N_17290,N_8459,N_8336);
and U17291 (N_17291,N_10211,N_11860);
nand U17292 (N_17292,N_11473,N_8280);
nor U17293 (N_17293,N_12191,N_10158);
nand U17294 (N_17294,N_7099,N_10241);
xnor U17295 (N_17295,N_12297,N_11085);
or U17296 (N_17296,N_9078,N_6929);
nand U17297 (N_17297,N_8154,N_10844);
nand U17298 (N_17298,N_10067,N_9729);
or U17299 (N_17299,N_12077,N_6962);
nand U17300 (N_17300,N_10652,N_12027);
and U17301 (N_17301,N_12264,N_8826);
and U17302 (N_17302,N_11470,N_11069);
or U17303 (N_17303,N_6450,N_10050);
or U17304 (N_17304,N_10934,N_8964);
and U17305 (N_17305,N_12261,N_9514);
and U17306 (N_17306,N_6542,N_10288);
and U17307 (N_17307,N_12446,N_8215);
nor U17308 (N_17308,N_12165,N_7416);
nor U17309 (N_17309,N_10246,N_11136);
nand U17310 (N_17310,N_8505,N_6784);
and U17311 (N_17311,N_9225,N_9164);
and U17312 (N_17312,N_12247,N_8677);
and U17313 (N_17313,N_8227,N_9740);
nor U17314 (N_17314,N_8399,N_7789);
and U17315 (N_17315,N_11254,N_11817);
xnor U17316 (N_17316,N_6823,N_8642);
and U17317 (N_17317,N_9901,N_12054);
or U17318 (N_17318,N_11796,N_8375);
and U17319 (N_17319,N_12362,N_8969);
nand U17320 (N_17320,N_6468,N_8839);
nor U17321 (N_17321,N_7851,N_11887);
and U17322 (N_17322,N_6735,N_10039);
nor U17323 (N_17323,N_9525,N_7768);
and U17324 (N_17324,N_12193,N_9982);
and U17325 (N_17325,N_9391,N_7830);
or U17326 (N_17326,N_11171,N_8540);
and U17327 (N_17327,N_11696,N_9246);
and U17328 (N_17328,N_8861,N_9486);
nand U17329 (N_17329,N_9432,N_9799);
and U17330 (N_17330,N_9813,N_11836);
or U17331 (N_17331,N_9184,N_6822);
or U17332 (N_17332,N_8160,N_7661);
nor U17333 (N_17333,N_10756,N_8282);
and U17334 (N_17334,N_8944,N_12022);
nor U17335 (N_17335,N_11186,N_8534);
nor U17336 (N_17336,N_12438,N_7641);
or U17337 (N_17337,N_7103,N_8096);
or U17338 (N_17338,N_8611,N_6596);
and U17339 (N_17339,N_11835,N_7823);
or U17340 (N_17340,N_8879,N_10135);
nor U17341 (N_17341,N_7468,N_10870);
or U17342 (N_17342,N_9647,N_6890);
nand U17343 (N_17343,N_7949,N_8282);
nand U17344 (N_17344,N_7261,N_11364);
or U17345 (N_17345,N_8139,N_6387);
or U17346 (N_17346,N_10847,N_7961);
nand U17347 (N_17347,N_9942,N_9485);
or U17348 (N_17348,N_11008,N_12072);
or U17349 (N_17349,N_11359,N_7486);
nor U17350 (N_17350,N_7940,N_6910);
or U17351 (N_17351,N_10261,N_10914);
and U17352 (N_17352,N_11759,N_6564);
and U17353 (N_17353,N_8305,N_6583);
or U17354 (N_17354,N_9253,N_7436);
or U17355 (N_17355,N_10778,N_7920);
nor U17356 (N_17356,N_6644,N_11712);
xor U17357 (N_17357,N_8848,N_10910);
nand U17358 (N_17358,N_7672,N_8575);
nand U17359 (N_17359,N_9162,N_10412);
nor U17360 (N_17360,N_11511,N_6468);
nand U17361 (N_17361,N_11227,N_11150);
nand U17362 (N_17362,N_10445,N_10163);
or U17363 (N_17363,N_7532,N_10725);
or U17364 (N_17364,N_6986,N_11000);
or U17365 (N_17365,N_7871,N_6254);
or U17366 (N_17366,N_12096,N_10432);
nor U17367 (N_17367,N_8424,N_6742);
nor U17368 (N_17368,N_10860,N_6389);
or U17369 (N_17369,N_9773,N_10544);
nand U17370 (N_17370,N_11678,N_6785);
nor U17371 (N_17371,N_10497,N_7844);
nand U17372 (N_17372,N_7616,N_9980);
and U17373 (N_17373,N_9581,N_11382);
nand U17374 (N_17374,N_9358,N_6782);
and U17375 (N_17375,N_9606,N_8889);
nor U17376 (N_17376,N_10262,N_10182);
and U17377 (N_17377,N_6295,N_9962);
or U17378 (N_17378,N_7762,N_7952);
nand U17379 (N_17379,N_8722,N_9546);
nor U17380 (N_17380,N_10095,N_9487);
nand U17381 (N_17381,N_12359,N_11503);
xnor U17382 (N_17382,N_8526,N_9325);
xnor U17383 (N_17383,N_6663,N_9732);
and U17384 (N_17384,N_9335,N_7788);
nand U17385 (N_17385,N_10433,N_10792);
or U17386 (N_17386,N_7759,N_6507);
and U17387 (N_17387,N_8200,N_7681);
or U17388 (N_17388,N_8812,N_9756);
nand U17389 (N_17389,N_9413,N_8461);
or U17390 (N_17390,N_8649,N_12147);
and U17391 (N_17391,N_11985,N_11322);
nor U17392 (N_17392,N_8803,N_6582);
xnor U17393 (N_17393,N_9806,N_10997);
nor U17394 (N_17394,N_8995,N_10215);
xor U17395 (N_17395,N_9102,N_10698);
xnor U17396 (N_17396,N_8576,N_11752);
nand U17397 (N_17397,N_8212,N_12354);
and U17398 (N_17398,N_7191,N_6835);
and U17399 (N_17399,N_8377,N_6945);
xnor U17400 (N_17400,N_9155,N_11281);
and U17401 (N_17401,N_8594,N_7665);
or U17402 (N_17402,N_7314,N_10724);
nor U17403 (N_17403,N_7893,N_9385);
or U17404 (N_17404,N_11254,N_11592);
or U17405 (N_17405,N_9919,N_10933);
xor U17406 (N_17406,N_7187,N_7906);
or U17407 (N_17407,N_7010,N_10492);
or U17408 (N_17408,N_11725,N_9532);
or U17409 (N_17409,N_9638,N_7088);
nand U17410 (N_17410,N_6868,N_9547);
nand U17411 (N_17411,N_9769,N_10119);
nand U17412 (N_17412,N_7243,N_11731);
nand U17413 (N_17413,N_8361,N_8291);
nor U17414 (N_17414,N_10186,N_11785);
or U17415 (N_17415,N_8287,N_6504);
xor U17416 (N_17416,N_10298,N_9332);
or U17417 (N_17417,N_10164,N_8658);
and U17418 (N_17418,N_8916,N_9591);
nor U17419 (N_17419,N_9996,N_6405);
or U17420 (N_17420,N_7344,N_9685);
xnor U17421 (N_17421,N_11740,N_7419);
nor U17422 (N_17422,N_11408,N_7713);
nand U17423 (N_17423,N_7665,N_9696);
nand U17424 (N_17424,N_9774,N_12319);
or U17425 (N_17425,N_10933,N_8184);
or U17426 (N_17426,N_10227,N_9370);
nor U17427 (N_17427,N_7732,N_11935);
and U17428 (N_17428,N_10014,N_9375);
nand U17429 (N_17429,N_12195,N_10958);
nor U17430 (N_17430,N_8225,N_12250);
nand U17431 (N_17431,N_9585,N_11317);
or U17432 (N_17432,N_6477,N_7936);
nand U17433 (N_17433,N_11160,N_10441);
nand U17434 (N_17434,N_9070,N_8977);
or U17435 (N_17435,N_7762,N_7820);
and U17436 (N_17436,N_11046,N_12150);
and U17437 (N_17437,N_6530,N_11420);
xor U17438 (N_17438,N_10701,N_10094);
nor U17439 (N_17439,N_6334,N_8414);
nand U17440 (N_17440,N_7183,N_11440);
and U17441 (N_17441,N_8191,N_8733);
nand U17442 (N_17442,N_9733,N_12165);
and U17443 (N_17443,N_9978,N_8597);
or U17444 (N_17444,N_9978,N_12310);
nor U17445 (N_17445,N_8528,N_7416);
nor U17446 (N_17446,N_11933,N_9485);
nor U17447 (N_17447,N_11348,N_10346);
or U17448 (N_17448,N_10418,N_9800);
and U17449 (N_17449,N_11990,N_10328);
xnor U17450 (N_17450,N_10090,N_7470);
nand U17451 (N_17451,N_9473,N_10549);
nand U17452 (N_17452,N_12490,N_9882);
nand U17453 (N_17453,N_8980,N_12109);
and U17454 (N_17454,N_8423,N_7481);
nor U17455 (N_17455,N_12060,N_8769);
and U17456 (N_17456,N_10537,N_8628);
xnor U17457 (N_17457,N_12078,N_7613);
nand U17458 (N_17458,N_11568,N_6647);
and U17459 (N_17459,N_7785,N_9893);
xor U17460 (N_17460,N_10224,N_11571);
nor U17461 (N_17461,N_9788,N_12114);
and U17462 (N_17462,N_7998,N_8687);
nor U17463 (N_17463,N_12361,N_6471);
or U17464 (N_17464,N_9971,N_8481);
or U17465 (N_17465,N_9363,N_8754);
or U17466 (N_17466,N_11196,N_7159);
and U17467 (N_17467,N_8138,N_11249);
nand U17468 (N_17468,N_8362,N_10408);
nand U17469 (N_17469,N_10508,N_9482);
xor U17470 (N_17470,N_11232,N_7168);
nor U17471 (N_17471,N_11043,N_6832);
nand U17472 (N_17472,N_7154,N_8206);
nand U17473 (N_17473,N_7273,N_10453);
and U17474 (N_17474,N_12056,N_6370);
nand U17475 (N_17475,N_9566,N_12280);
or U17476 (N_17476,N_8429,N_8419);
nor U17477 (N_17477,N_12169,N_9127);
and U17478 (N_17478,N_6390,N_6699);
nand U17479 (N_17479,N_10188,N_11338);
or U17480 (N_17480,N_6929,N_11508);
nor U17481 (N_17481,N_9848,N_10862);
and U17482 (N_17482,N_11224,N_7112);
nor U17483 (N_17483,N_10533,N_11794);
nor U17484 (N_17484,N_8938,N_8411);
nand U17485 (N_17485,N_7520,N_12486);
or U17486 (N_17486,N_11570,N_11775);
xor U17487 (N_17487,N_7848,N_6269);
nand U17488 (N_17488,N_12276,N_7414);
nor U17489 (N_17489,N_7044,N_8656);
nand U17490 (N_17490,N_8407,N_10302);
nor U17491 (N_17491,N_8011,N_11944);
nand U17492 (N_17492,N_9255,N_8105);
and U17493 (N_17493,N_10335,N_10641);
or U17494 (N_17494,N_11156,N_7380);
nor U17495 (N_17495,N_12286,N_7396);
or U17496 (N_17496,N_11347,N_6852);
xor U17497 (N_17497,N_9516,N_8854);
nor U17498 (N_17498,N_10751,N_11583);
and U17499 (N_17499,N_10439,N_9910);
or U17500 (N_17500,N_8148,N_9129);
nand U17501 (N_17501,N_9046,N_6483);
nand U17502 (N_17502,N_11373,N_12418);
nor U17503 (N_17503,N_8883,N_8429);
xor U17504 (N_17504,N_8118,N_9286);
nor U17505 (N_17505,N_10898,N_6398);
and U17506 (N_17506,N_12295,N_10322);
nand U17507 (N_17507,N_9996,N_11999);
nor U17508 (N_17508,N_9730,N_10131);
and U17509 (N_17509,N_8677,N_9402);
xnor U17510 (N_17510,N_8261,N_6836);
nand U17511 (N_17511,N_9360,N_8232);
nor U17512 (N_17512,N_11865,N_10938);
nor U17513 (N_17513,N_10738,N_10120);
nand U17514 (N_17514,N_8411,N_12307);
nand U17515 (N_17515,N_9013,N_12078);
xor U17516 (N_17516,N_11805,N_8796);
and U17517 (N_17517,N_9026,N_8448);
nor U17518 (N_17518,N_7689,N_8469);
nand U17519 (N_17519,N_11233,N_8439);
nand U17520 (N_17520,N_12471,N_6750);
or U17521 (N_17521,N_9377,N_8922);
or U17522 (N_17522,N_7761,N_6881);
and U17523 (N_17523,N_10467,N_7606);
nand U17524 (N_17524,N_12081,N_11179);
or U17525 (N_17525,N_8355,N_12358);
and U17526 (N_17526,N_11473,N_7741);
nor U17527 (N_17527,N_11013,N_9896);
or U17528 (N_17528,N_7213,N_6928);
xor U17529 (N_17529,N_9321,N_8666);
or U17530 (N_17530,N_9315,N_6713);
xor U17531 (N_17531,N_7954,N_11923);
nand U17532 (N_17532,N_10357,N_8070);
or U17533 (N_17533,N_12226,N_9987);
nand U17534 (N_17534,N_9071,N_11178);
and U17535 (N_17535,N_7524,N_7362);
nand U17536 (N_17536,N_9008,N_10574);
nand U17537 (N_17537,N_10660,N_6388);
xnor U17538 (N_17538,N_8058,N_6821);
and U17539 (N_17539,N_7669,N_8018);
nand U17540 (N_17540,N_9286,N_8031);
and U17541 (N_17541,N_11857,N_8366);
nor U17542 (N_17542,N_9722,N_8173);
nand U17543 (N_17543,N_8674,N_6631);
nand U17544 (N_17544,N_12416,N_9429);
and U17545 (N_17545,N_8683,N_9694);
or U17546 (N_17546,N_10090,N_11559);
or U17547 (N_17547,N_10160,N_9340);
and U17548 (N_17548,N_8897,N_10593);
and U17549 (N_17549,N_9729,N_7328);
nor U17550 (N_17550,N_8353,N_7994);
nor U17551 (N_17551,N_6717,N_9982);
xor U17552 (N_17552,N_9176,N_7627);
and U17553 (N_17553,N_10257,N_7306);
xor U17554 (N_17554,N_11207,N_6786);
nand U17555 (N_17555,N_10621,N_7451);
nor U17556 (N_17556,N_8181,N_11007);
and U17557 (N_17557,N_11941,N_6907);
nor U17558 (N_17558,N_11577,N_11315);
and U17559 (N_17559,N_8413,N_7606);
nor U17560 (N_17560,N_7620,N_7483);
nor U17561 (N_17561,N_9797,N_9961);
or U17562 (N_17562,N_9064,N_8223);
nor U17563 (N_17563,N_10401,N_11112);
or U17564 (N_17564,N_7654,N_8953);
nor U17565 (N_17565,N_11277,N_8722);
or U17566 (N_17566,N_6451,N_10766);
or U17567 (N_17567,N_12141,N_9140);
or U17568 (N_17568,N_8189,N_12051);
nand U17569 (N_17569,N_8573,N_10576);
and U17570 (N_17570,N_11268,N_7274);
or U17571 (N_17571,N_7209,N_10072);
and U17572 (N_17572,N_7276,N_9030);
nor U17573 (N_17573,N_6318,N_6557);
or U17574 (N_17574,N_7066,N_6843);
and U17575 (N_17575,N_6725,N_6466);
nor U17576 (N_17576,N_8755,N_6483);
nand U17577 (N_17577,N_11850,N_12114);
nor U17578 (N_17578,N_10112,N_7103);
or U17579 (N_17579,N_6654,N_11397);
or U17580 (N_17580,N_6809,N_11942);
and U17581 (N_17581,N_6854,N_11601);
nand U17582 (N_17582,N_9836,N_6782);
nand U17583 (N_17583,N_7795,N_7098);
or U17584 (N_17584,N_8368,N_11277);
xor U17585 (N_17585,N_11626,N_8675);
and U17586 (N_17586,N_10727,N_10744);
or U17587 (N_17587,N_10312,N_8583);
nor U17588 (N_17588,N_11056,N_7228);
nor U17589 (N_17589,N_11971,N_8702);
and U17590 (N_17590,N_7079,N_12026);
or U17591 (N_17591,N_8781,N_9345);
or U17592 (N_17592,N_9645,N_6579);
and U17593 (N_17593,N_9430,N_6479);
or U17594 (N_17594,N_11253,N_6408);
nor U17595 (N_17595,N_6985,N_10446);
and U17596 (N_17596,N_11993,N_7393);
and U17597 (N_17597,N_10228,N_8262);
nor U17598 (N_17598,N_11724,N_8276);
nor U17599 (N_17599,N_10050,N_6480);
nor U17600 (N_17600,N_9034,N_10779);
nand U17601 (N_17601,N_11518,N_11382);
and U17602 (N_17602,N_11106,N_7803);
or U17603 (N_17603,N_7118,N_12280);
nor U17604 (N_17604,N_9076,N_11759);
nor U17605 (N_17605,N_6252,N_8772);
or U17606 (N_17606,N_8554,N_9393);
or U17607 (N_17607,N_10154,N_7140);
or U17608 (N_17608,N_8989,N_8713);
or U17609 (N_17609,N_11221,N_12495);
nor U17610 (N_17610,N_11367,N_6759);
nor U17611 (N_17611,N_11391,N_8911);
or U17612 (N_17612,N_11885,N_8644);
nand U17613 (N_17613,N_7603,N_11923);
and U17614 (N_17614,N_7406,N_7987);
nor U17615 (N_17615,N_9118,N_7030);
nand U17616 (N_17616,N_8600,N_8588);
nor U17617 (N_17617,N_10795,N_8259);
or U17618 (N_17618,N_6257,N_9572);
xnor U17619 (N_17619,N_7272,N_6608);
or U17620 (N_17620,N_7196,N_10342);
and U17621 (N_17621,N_9140,N_6399);
and U17622 (N_17622,N_9273,N_7381);
nor U17623 (N_17623,N_12097,N_11028);
nand U17624 (N_17624,N_12004,N_8626);
and U17625 (N_17625,N_7162,N_9821);
nand U17626 (N_17626,N_7826,N_9189);
or U17627 (N_17627,N_11648,N_8345);
xor U17628 (N_17628,N_10924,N_8044);
nor U17629 (N_17629,N_7494,N_8592);
or U17630 (N_17630,N_11492,N_8511);
nand U17631 (N_17631,N_8449,N_7144);
and U17632 (N_17632,N_6968,N_11541);
nor U17633 (N_17633,N_11920,N_8544);
or U17634 (N_17634,N_11311,N_9034);
and U17635 (N_17635,N_9863,N_9608);
nor U17636 (N_17636,N_9319,N_6919);
or U17637 (N_17637,N_9976,N_6858);
or U17638 (N_17638,N_7860,N_6677);
and U17639 (N_17639,N_7566,N_7591);
or U17640 (N_17640,N_8371,N_7842);
nand U17641 (N_17641,N_7414,N_11861);
or U17642 (N_17642,N_10644,N_8338);
or U17643 (N_17643,N_10413,N_12299);
or U17644 (N_17644,N_6560,N_6447);
nor U17645 (N_17645,N_7948,N_10652);
or U17646 (N_17646,N_8978,N_8246);
nor U17647 (N_17647,N_9626,N_10650);
nand U17648 (N_17648,N_8293,N_6513);
nand U17649 (N_17649,N_9301,N_8018);
xor U17650 (N_17650,N_10605,N_10409);
and U17651 (N_17651,N_11925,N_9854);
and U17652 (N_17652,N_9015,N_12359);
nand U17653 (N_17653,N_10917,N_10458);
and U17654 (N_17654,N_8692,N_12366);
or U17655 (N_17655,N_8831,N_11227);
or U17656 (N_17656,N_11640,N_8628);
or U17657 (N_17657,N_10681,N_10443);
and U17658 (N_17658,N_9520,N_9483);
or U17659 (N_17659,N_12484,N_8623);
nor U17660 (N_17660,N_8814,N_10295);
or U17661 (N_17661,N_7013,N_11338);
nand U17662 (N_17662,N_9833,N_10873);
nand U17663 (N_17663,N_11202,N_9729);
or U17664 (N_17664,N_8890,N_11958);
nand U17665 (N_17665,N_8045,N_7191);
nand U17666 (N_17666,N_8230,N_8069);
nand U17667 (N_17667,N_10928,N_10376);
or U17668 (N_17668,N_10237,N_9701);
nor U17669 (N_17669,N_12001,N_8521);
nand U17670 (N_17670,N_11363,N_8433);
xnor U17671 (N_17671,N_10624,N_11149);
or U17672 (N_17672,N_11875,N_6500);
or U17673 (N_17673,N_7632,N_11692);
nor U17674 (N_17674,N_8379,N_11840);
or U17675 (N_17675,N_12042,N_12340);
or U17676 (N_17676,N_6665,N_11895);
and U17677 (N_17677,N_8147,N_7199);
nand U17678 (N_17678,N_10200,N_9124);
and U17679 (N_17679,N_8840,N_8205);
nor U17680 (N_17680,N_11342,N_8877);
nor U17681 (N_17681,N_10367,N_8253);
or U17682 (N_17682,N_9132,N_7625);
and U17683 (N_17683,N_9901,N_9122);
and U17684 (N_17684,N_11226,N_9682);
or U17685 (N_17685,N_10118,N_9424);
nand U17686 (N_17686,N_10787,N_7865);
xnor U17687 (N_17687,N_12150,N_11044);
or U17688 (N_17688,N_7844,N_10834);
nor U17689 (N_17689,N_11771,N_9417);
or U17690 (N_17690,N_6256,N_12427);
nor U17691 (N_17691,N_9711,N_10614);
nor U17692 (N_17692,N_7861,N_6968);
xnor U17693 (N_17693,N_10829,N_10359);
xnor U17694 (N_17694,N_12307,N_7154);
nand U17695 (N_17695,N_12202,N_12003);
nor U17696 (N_17696,N_7717,N_9540);
or U17697 (N_17697,N_6770,N_12319);
nor U17698 (N_17698,N_7523,N_12102);
or U17699 (N_17699,N_11023,N_12039);
nor U17700 (N_17700,N_10876,N_12435);
nor U17701 (N_17701,N_7474,N_9747);
or U17702 (N_17702,N_6971,N_9957);
nand U17703 (N_17703,N_7627,N_10230);
and U17704 (N_17704,N_10396,N_6535);
or U17705 (N_17705,N_11372,N_9425);
nand U17706 (N_17706,N_7682,N_11935);
or U17707 (N_17707,N_8310,N_11227);
xnor U17708 (N_17708,N_9648,N_12400);
nor U17709 (N_17709,N_11532,N_7694);
or U17710 (N_17710,N_10814,N_10305);
xor U17711 (N_17711,N_8345,N_8912);
and U17712 (N_17712,N_8790,N_11955);
nor U17713 (N_17713,N_11628,N_9023);
or U17714 (N_17714,N_11780,N_11526);
or U17715 (N_17715,N_7410,N_8265);
nor U17716 (N_17716,N_11424,N_7776);
and U17717 (N_17717,N_8933,N_8629);
or U17718 (N_17718,N_6997,N_7213);
nor U17719 (N_17719,N_11247,N_11537);
nand U17720 (N_17720,N_8903,N_6765);
and U17721 (N_17721,N_10781,N_12058);
xor U17722 (N_17722,N_6760,N_7767);
nor U17723 (N_17723,N_7352,N_11152);
and U17724 (N_17724,N_6824,N_9911);
nor U17725 (N_17725,N_6501,N_9734);
and U17726 (N_17726,N_10012,N_11135);
nor U17727 (N_17727,N_11246,N_11765);
nor U17728 (N_17728,N_10745,N_8443);
nor U17729 (N_17729,N_9449,N_10095);
nand U17730 (N_17730,N_7386,N_6940);
or U17731 (N_17731,N_11615,N_11763);
and U17732 (N_17732,N_8206,N_11430);
and U17733 (N_17733,N_10988,N_8383);
or U17734 (N_17734,N_6724,N_11704);
nor U17735 (N_17735,N_7348,N_6502);
nand U17736 (N_17736,N_11733,N_11635);
and U17737 (N_17737,N_8102,N_10213);
nor U17738 (N_17738,N_11909,N_7335);
nand U17739 (N_17739,N_11855,N_12217);
or U17740 (N_17740,N_10280,N_11504);
or U17741 (N_17741,N_8915,N_8589);
or U17742 (N_17742,N_12069,N_10364);
or U17743 (N_17743,N_9618,N_12042);
and U17744 (N_17744,N_7211,N_11350);
and U17745 (N_17745,N_8388,N_6767);
or U17746 (N_17746,N_7933,N_7486);
xor U17747 (N_17747,N_12310,N_9967);
or U17748 (N_17748,N_8694,N_10453);
and U17749 (N_17749,N_9318,N_11969);
nand U17750 (N_17750,N_9166,N_12258);
nor U17751 (N_17751,N_10561,N_9636);
nand U17752 (N_17752,N_7906,N_7165);
or U17753 (N_17753,N_9395,N_11681);
or U17754 (N_17754,N_12173,N_8819);
and U17755 (N_17755,N_11656,N_7335);
nand U17756 (N_17756,N_6955,N_8131);
nor U17757 (N_17757,N_10189,N_7409);
and U17758 (N_17758,N_8156,N_7930);
nor U17759 (N_17759,N_11718,N_8123);
nand U17760 (N_17760,N_10172,N_6804);
or U17761 (N_17761,N_10202,N_9260);
xor U17762 (N_17762,N_10593,N_10005);
or U17763 (N_17763,N_8800,N_8261);
or U17764 (N_17764,N_9481,N_8330);
and U17765 (N_17765,N_9618,N_11725);
xnor U17766 (N_17766,N_11504,N_7712);
nor U17767 (N_17767,N_8047,N_6552);
and U17768 (N_17768,N_11038,N_11071);
or U17769 (N_17769,N_6905,N_10658);
nand U17770 (N_17770,N_6578,N_10379);
xnor U17771 (N_17771,N_7448,N_7671);
nand U17772 (N_17772,N_8783,N_6819);
and U17773 (N_17773,N_10905,N_9566);
nor U17774 (N_17774,N_12431,N_7483);
nand U17775 (N_17775,N_10054,N_8489);
or U17776 (N_17776,N_9412,N_11065);
or U17777 (N_17777,N_8961,N_6432);
nor U17778 (N_17778,N_7994,N_9065);
or U17779 (N_17779,N_11734,N_9600);
or U17780 (N_17780,N_7129,N_11726);
or U17781 (N_17781,N_8576,N_12139);
xnor U17782 (N_17782,N_7665,N_8009);
and U17783 (N_17783,N_10194,N_8845);
xor U17784 (N_17784,N_11460,N_6682);
nor U17785 (N_17785,N_9383,N_11270);
nand U17786 (N_17786,N_11523,N_11694);
nand U17787 (N_17787,N_11908,N_8742);
xnor U17788 (N_17788,N_11562,N_7653);
nor U17789 (N_17789,N_10997,N_9432);
and U17790 (N_17790,N_8629,N_10785);
xnor U17791 (N_17791,N_11547,N_8076);
nand U17792 (N_17792,N_8242,N_7714);
and U17793 (N_17793,N_7369,N_8251);
and U17794 (N_17794,N_10233,N_9654);
nand U17795 (N_17795,N_7923,N_7983);
and U17796 (N_17796,N_12349,N_8665);
nor U17797 (N_17797,N_11434,N_6399);
or U17798 (N_17798,N_10141,N_11386);
nor U17799 (N_17799,N_7030,N_7745);
or U17800 (N_17800,N_8771,N_11004);
and U17801 (N_17801,N_7750,N_8268);
nor U17802 (N_17802,N_7596,N_7028);
nor U17803 (N_17803,N_9300,N_6352);
nand U17804 (N_17804,N_9207,N_7986);
nand U17805 (N_17805,N_9896,N_8912);
xnor U17806 (N_17806,N_10499,N_9606);
nand U17807 (N_17807,N_11319,N_6838);
nor U17808 (N_17808,N_10577,N_11493);
or U17809 (N_17809,N_9991,N_6577);
and U17810 (N_17810,N_6784,N_9098);
and U17811 (N_17811,N_12364,N_7656);
and U17812 (N_17812,N_9096,N_9657);
or U17813 (N_17813,N_12135,N_7969);
and U17814 (N_17814,N_8760,N_11972);
or U17815 (N_17815,N_10170,N_12406);
and U17816 (N_17816,N_9981,N_11106);
and U17817 (N_17817,N_7065,N_8696);
and U17818 (N_17818,N_12341,N_8426);
and U17819 (N_17819,N_11898,N_8577);
or U17820 (N_17820,N_8880,N_10538);
or U17821 (N_17821,N_12392,N_8895);
and U17822 (N_17822,N_12248,N_11512);
xor U17823 (N_17823,N_7561,N_6843);
or U17824 (N_17824,N_7463,N_6427);
nor U17825 (N_17825,N_7766,N_7555);
xor U17826 (N_17826,N_9448,N_11904);
and U17827 (N_17827,N_9687,N_11400);
nor U17828 (N_17828,N_11073,N_6623);
nand U17829 (N_17829,N_9412,N_6872);
nor U17830 (N_17830,N_10335,N_12294);
or U17831 (N_17831,N_6380,N_8596);
xor U17832 (N_17832,N_10551,N_6602);
or U17833 (N_17833,N_11773,N_7555);
or U17834 (N_17834,N_9124,N_7767);
nand U17835 (N_17835,N_11719,N_9060);
and U17836 (N_17836,N_11726,N_12046);
nand U17837 (N_17837,N_10181,N_10217);
or U17838 (N_17838,N_7080,N_10253);
nand U17839 (N_17839,N_11063,N_9520);
or U17840 (N_17840,N_7689,N_6462);
nor U17841 (N_17841,N_8835,N_9037);
nand U17842 (N_17842,N_10169,N_12018);
or U17843 (N_17843,N_11008,N_9116);
and U17844 (N_17844,N_11554,N_6360);
or U17845 (N_17845,N_9760,N_6555);
or U17846 (N_17846,N_7114,N_9940);
and U17847 (N_17847,N_11458,N_11510);
or U17848 (N_17848,N_6920,N_8423);
or U17849 (N_17849,N_10766,N_10265);
or U17850 (N_17850,N_9836,N_11023);
xor U17851 (N_17851,N_11698,N_11203);
and U17852 (N_17852,N_10951,N_8025);
or U17853 (N_17853,N_10928,N_9001);
or U17854 (N_17854,N_10459,N_7904);
and U17855 (N_17855,N_7400,N_6817);
and U17856 (N_17856,N_12460,N_9372);
and U17857 (N_17857,N_7019,N_11215);
nand U17858 (N_17858,N_9730,N_7175);
nand U17859 (N_17859,N_12290,N_10255);
nand U17860 (N_17860,N_7430,N_9993);
or U17861 (N_17861,N_6732,N_8607);
and U17862 (N_17862,N_6635,N_8728);
and U17863 (N_17863,N_11618,N_8873);
nor U17864 (N_17864,N_11147,N_12368);
nand U17865 (N_17865,N_9339,N_10616);
and U17866 (N_17866,N_6408,N_10124);
and U17867 (N_17867,N_7004,N_10673);
or U17868 (N_17868,N_7253,N_8381);
nor U17869 (N_17869,N_9718,N_10268);
and U17870 (N_17870,N_10914,N_11634);
or U17871 (N_17871,N_9258,N_11385);
nor U17872 (N_17872,N_12059,N_10183);
or U17873 (N_17873,N_9228,N_11131);
nand U17874 (N_17874,N_12431,N_9407);
nand U17875 (N_17875,N_6571,N_9629);
xor U17876 (N_17876,N_7442,N_10318);
nand U17877 (N_17877,N_11386,N_10942);
nor U17878 (N_17878,N_12065,N_11800);
and U17879 (N_17879,N_9130,N_7413);
nand U17880 (N_17880,N_11868,N_6450);
nor U17881 (N_17881,N_8443,N_9126);
nor U17882 (N_17882,N_11634,N_8320);
nor U17883 (N_17883,N_6596,N_8641);
and U17884 (N_17884,N_9280,N_6438);
nand U17885 (N_17885,N_9931,N_12338);
xnor U17886 (N_17886,N_12280,N_10956);
or U17887 (N_17887,N_8346,N_9121);
or U17888 (N_17888,N_6478,N_6255);
nand U17889 (N_17889,N_8635,N_10768);
and U17890 (N_17890,N_9534,N_9615);
nor U17891 (N_17891,N_10902,N_11104);
nor U17892 (N_17892,N_8771,N_10605);
nor U17893 (N_17893,N_10244,N_11423);
nand U17894 (N_17894,N_10030,N_9209);
and U17895 (N_17895,N_6394,N_10405);
nand U17896 (N_17896,N_9536,N_11551);
nor U17897 (N_17897,N_6458,N_9469);
nor U17898 (N_17898,N_7533,N_11844);
nand U17899 (N_17899,N_11129,N_11167);
or U17900 (N_17900,N_9475,N_7445);
and U17901 (N_17901,N_7329,N_6477);
and U17902 (N_17902,N_10442,N_6277);
nand U17903 (N_17903,N_9319,N_7270);
and U17904 (N_17904,N_9501,N_8021);
nor U17905 (N_17905,N_7585,N_8566);
or U17906 (N_17906,N_11512,N_10475);
and U17907 (N_17907,N_8488,N_7552);
and U17908 (N_17908,N_9514,N_8920);
and U17909 (N_17909,N_11236,N_7460);
or U17910 (N_17910,N_12386,N_9896);
or U17911 (N_17911,N_8434,N_7778);
nor U17912 (N_17912,N_6444,N_9952);
or U17913 (N_17913,N_6801,N_8132);
nand U17914 (N_17914,N_7830,N_11646);
nor U17915 (N_17915,N_10634,N_9586);
nor U17916 (N_17916,N_7146,N_7847);
and U17917 (N_17917,N_10336,N_9305);
xnor U17918 (N_17918,N_12365,N_10490);
nor U17919 (N_17919,N_11444,N_11815);
or U17920 (N_17920,N_9702,N_6571);
and U17921 (N_17921,N_7820,N_6752);
nand U17922 (N_17922,N_11653,N_12496);
or U17923 (N_17923,N_6760,N_6747);
and U17924 (N_17924,N_6861,N_9140);
and U17925 (N_17925,N_6891,N_9531);
xnor U17926 (N_17926,N_6999,N_6544);
xor U17927 (N_17927,N_11686,N_8277);
nand U17928 (N_17928,N_7997,N_8413);
nor U17929 (N_17929,N_8563,N_6563);
or U17930 (N_17930,N_10953,N_8521);
nand U17931 (N_17931,N_7918,N_8172);
nor U17932 (N_17932,N_8292,N_7356);
and U17933 (N_17933,N_11728,N_8737);
nand U17934 (N_17934,N_10061,N_9028);
nor U17935 (N_17935,N_8912,N_11161);
xor U17936 (N_17936,N_11138,N_8310);
xnor U17937 (N_17937,N_9813,N_8099);
or U17938 (N_17938,N_6319,N_7105);
and U17939 (N_17939,N_9441,N_11572);
and U17940 (N_17940,N_11868,N_9108);
and U17941 (N_17941,N_6445,N_11980);
nor U17942 (N_17942,N_10377,N_6597);
or U17943 (N_17943,N_8653,N_9172);
nand U17944 (N_17944,N_9396,N_12349);
or U17945 (N_17945,N_9767,N_11816);
or U17946 (N_17946,N_10068,N_12368);
xnor U17947 (N_17947,N_8042,N_9110);
and U17948 (N_17948,N_10655,N_7759);
xnor U17949 (N_17949,N_8132,N_11948);
or U17950 (N_17950,N_10638,N_7395);
or U17951 (N_17951,N_7976,N_9439);
or U17952 (N_17952,N_8644,N_10951);
and U17953 (N_17953,N_6342,N_10011);
nor U17954 (N_17954,N_6542,N_9695);
xnor U17955 (N_17955,N_8829,N_10288);
nand U17956 (N_17956,N_6919,N_7795);
or U17957 (N_17957,N_10770,N_10137);
nand U17958 (N_17958,N_8307,N_6667);
and U17959 (N_17959,N_8917,N_9719);
xnor U17960 (N_17960,N_10115,N_10648);
nor U17961 (N_17961,N_11406,N_10107);
nand U17962 (N_17962,N_9448,N_8909);
xnor U17963 (N_17963,N_7820,N_11927);
nor U17964 (N_17964,N_8398,N_9334);
or U17965 (N_17965,N_10390,N_11607);
nor U17966 (N_17966,N_12085,N_9621);
xor U17967 (N_17967,N_10111,N_10818);
nand U17968 (N_17968,N_11671,N_9234);
and U17969 (N_17969,N_10291,N_12153);
nand U17970 (N_17970,N_9302,N_10648);
or U17971 (N_17971,N_11948,N_8561);
nor U17972 (N_17972,N_11960,N_11740);
nand U17973 (N_17973,N_7315,N_10194);
nor U17974 (N_17974,N_8672,N_8883);
or U17975 (N_17975,N_10663,N_10420);
or U17976 (N_17976,N_7586,N_6494);
xor U17977 (N_17977,N_6429,N_9902);
or U17978 (N_17978,N_8486,N_10702);
nand U17979 (N_17979,N_6966,N_12409);
and U17980 (N_17980,N_8249,N_12112);
nand U17981 (N_17981,N_9467,N_10838);
nor U17982 (N_17982,N_9696,N_7466);
nand U17983 (N_17983,N_11557,N_7720);
xnor U17984 (N_17984,N_12402,N_11249);
or U17985 (N_17985,N_12199,N_9758);
nor U17986 (N_17986,N_9257,N_9677);
and U17987 (N_17987,N_8504,N_10120);
and U17988 (N_17988,N_11211,N_8935);
and U17989 (N_17989,N_9843,N_6466);
nand U17990 (N_17990,N_11379,N_9354);
nor U17991 (N_17991,N_6329,N_10620);
nor U17992 (N_17992,N_8898,N_11690);
nand U17993 (N_17993,N_6378,N_6866);
nor U17994 (N_17994,N_7100,N_11902);
nand U17995 (N_17995,N_8657,N_7205);
xor U17996 (N_17996,N_11386,N_6931);
xnor U17997 (N_17997,N_11813,N_9558);
nor U17998 (N_17998,N_11683,N_9180);
and U17999 (N_17999,N_11421,N_7956);
nand U18000 (N_18000,N_7899,N_6320);
nor U18001 (N_18001,N_8820,N_7458);
xor U18002 (N_18002,N_7904,N_7554);
nor U18003 (N_18003,N_9044,N_8676);
nand U18004 (N_18004,N_7945,N_7611);
nand U18005 (N_18005,N_7477,N_7995);
nand U18006 (N_18006,N_11388,N_12063);
nor U18007 (N_18007,N_11037,N_9650);
nor U18008 (N_18008,N_7200,N_9855);
nor U18009 (N_18009,N_7210,N_10994);
nor U18010 (N_18010,N_9294,N_6343);
or U18011 (N_18011,N_10718,N_7333);
nor U18012 (N_18012,N_6316,N_11047);
xnor U18013 (N_18013,N_11452,N_12263);
nand U18014 (N_18014,N_11148,N_10016);
nor U18015 (N_18015,N_12229,N_10889);
nand U18016 (N_18016,N_7741,N_7971);
xnor U18017 (N_18017,N_7150,N_11386);
and U18018 (N_18018,N_10419,N_7057);
nand U18019 (N_18019,N_7382,N_8157);
nand U18020 (N_18020,N_9392,N_7858);
and U18021 (N_18021,N_10670,N_11758);
and U18022 (N_18022,N_7217,N_7793);
nor U18023 (N_18023,N_11239,N_8696);
nor U18024 (N_18024,N_7747,N_9304);
and U18025 (N_18025,N_11010,N_7562);
nor U18026 (N_18026,N_6388,N_10890);
and U18027 (N_18027,N_11793,N_9933);
nor U18028 (N_18028,N_9691,N_8827);
or U18029 (N_18029,N_12472,N_7891);
or U18030 (N_18030,N_7980,N_8604);
and U18031 (N_18031,N_12011,N_7798);
nor U18032 (N_18032,N_11143,N_8172);
or U18033 (N_18033,N_6727,N_9382);
nand U18034 (N_18034,N_7793,N_7710);
nand U18035 (N_18035,N_6992,N_9822);
nor U18036 (N_18036,N_9558,N_10049);
and U18037 (N_18037,N_10557,N_9914);
nor U18038 (N_18038,N_7901,N_8411);
nand U18039 (N_18039,N_7142,N_9334);
and U18040 (N_18040,N_9821,N_10427);
nor U18041 (N_18041,N_8604,N_11177);
xnor U18042 (N_18042,N_6724,N_12005);
and U18043 (N_18043,N_7613,N_6388);
nand U18044 (N_18044,N_6504,N_6785);
and U18045 (N_18045,N_8976,N_7024);
and U18046 (N_18046,N_6501,N_9576);
nor U18047 (N_18047,N_10851,N_8484);
nand U18048 (N_18048,N_6386,N_7837);
nand U18049 (N_18049,N_8529,N_6986);
nand U18050 (N_18050,N_12046,N_7129);
and U18051 (N_18051,N_9904,N_8362);
and U18052 (N_18052,N_7885,N_12413);
and U18053 (N_18053,N_12155,N_9386);
or U18054 (N_18054,N_6775,N_6646);
nand U18055 (N_18055,N_9017,N_10889);
nand U18056 (N_18056,N_9024,N_10949);
and U18057 (N_18057,N_9326,N_8045);
nor U18058 (N_18058,N_12225,N_11356);
nand U18059 (N_18059,N_6358,N_12108);
nand U18060 (N_18060,N_6690,N_6896);
xor U18061 (N_18061,N_11207,N_7144);
and U18062 (N_18062,N_6273,N_10775);
nor U18063 (N_18063,N_12222,N_12076);
or U18064 (N_18064,N_8264,N_10788);
or U18065 (N_18065,N_11162,N_10909);
or U18066 (N_18066,N_9749,N_7502);
nand U18067 (N_18067,N_10800,N_6427);
nand U18068 (N_18068,N_10334,N_7391);
nand U18069 (N_18069,N_12012,N_7872);
xnor U18070 (N_18070,N_8187,N_7270);
nand U18071 (N_18071,N_11375,N_8154);
xor U18072 (N_18072,N_7740,N_8154);
and U18073 (N_18073,N_6719,N_10821);
nor U18074 (N_18074,N_7444,N_9101);
nand U18075 (N_18075,N_8029,N_7290);
and U18076 (N_18076,N_9002,N_7751);
or U18077 (N_18077,N_11632,N_9905);
and U18078 (N_18078,N_10765,N_6641);
nor U18079 (N_18079,N_6597,N_9243);
or U18080 (N_18080,N_6250,N_10982);
and U18081 (N_18081,N_6630,N_9805);
or U18082 (N_18082,N_11138,N_9857);
or U18083 (N_18083,N_6333,N_6693);
nor U18084 (N_18084,N_12056,N_10125);
nand U18085 (N_18085,N_6547,N_7041);
xnor U18086 (N_18086,N_11446,N_9212);
and U18087 (N_18087,N_9951,N_11603);
nand U18088 (N_18088,N_11887,N_10713);
xor U18089 (N_18089,N_11642,N_11897);
and U18090 (N_18090,N_9745,N_8800);
or U18091 (N_18091,N_7030,N_12467);
xnor U18092 (N_18092,N_9376,N_12071);
nand U18093 (N_18093,N_12365,N_12366);
nand U18094 (N_18094,N_7171,N_6451);
xnor U18095 (N_18095,N_9959,N_9905);
nor U18096 (N_18096,N_10249,N_8230);
nor U18097 (N_18097,N_10175,N_6510);
and U18098 (N_18098,N_8712,N_11156);
and U18099 (N_18099,N_7460,N_7389);
and U18100 (N_18100,N_9468,N_11226);
nor U18101 (N_18101,N_11131,N_10643);
or U18102 (N_18102,N_10036,N_8861);
or U18103 (N_18103,N_12035,N_7331);
nor U18104 (N_18104,N_9667,N_9518);
and U18105 (N_18105,N_10962,N_9342);
xnor U18106 (N_18106,N_8151,N_7022);
xor U18107 (N_18107,N_7629,N_7638);
xor U18108 (N_18108,N_9852,N_7543);
nor U18109 (N_18109,N_11085,N_11676);
nand U18110 (N_18110,N_7768,N_8807);
and U18111 (N_18111,N_7342,N_10617);
and U18112 (N_18112,N_8491,N_8648);
or U18113 (N_18113,N_9009,N_7547);
and U18114 (N_18114,N_12063,N_10157);
or U18115 (N_18115,N_8483,N_7512);
and U18116 (N_18116,N_7223,N_11289);
and U18117 (N_18117,N_11803,N_9508);
nor U18118 (N_18118,N_7883,N_6878);
and U18119 (N_18119,N_8111,N_11693);
nand U18120 (N_18120,N_10333,N_7737);
nor U18121 (N_18121,N_9434,N_11938);
xor U18122 (N_18122,N_7230,N_9864);
nand U18123 (N_18123,N_9556,N_9213);
or U18124 (N_18124,N_8766,N_6875);
and U18125 (N_18125,N_11166,N_9497);
and U18126 (N_18126,N_6820,N_8538);
nand U18127 (N_18127,N_10449,N_11633);
or U18128 (N_18128,N_10364,N_10688);
nand U18129 (N_18129,N_8107,N_6955);
xor U18130 (N_18130,N_7169,N_10853);
xnor U18131 (N_18131,N_12417,N_7560);
nand U18132 (N_18132,N_7667,N_6720);
and U18133 (N_18133,N_10544,N_7043);
nor U18134 (N_18134,N_6357,N_8253);
and U18135 (N_18135,N_10545,N_11689);
nor U18136 (N_18136,N_9821,N_10619);
xnor U18137 (N_18137,N_10070,N_11949);
xnor U18138 (N_18138,N_11803,N_7902);
xnor U18139 (N_18139,N_7883,N_6584);
and U18140 (N_18140,N_9367,N_8381);
or U18141 (N_18141,N_7857,N_12488);
or U18142 (N_18142,N_10022,N_9327);
and U18143 (N_18143,N_11681,N_6438);
nand U18144 (N_18144,N_9833,N_10884);
nor U18145 (N_18145,N_7590,N_8565);
nand U18146 (N_18146,N_6875,N_11185);
nor U18147 (N_18147,N_8028,N_6435);
nand U18148 (N_18148,N_6549,N_7174);
nand U18149 (N_18149,N_6985,N_6420);
nor U18150 (N_18150,N_8727,N_9850);
nor U18151 (N_18151,N_9707,N_11009);
nand U18152 (N_18152,N_9580,N_12380);
nor U18153 (N_18153,N_8972,N_11322);
or U18154 (N_18154,N_8244,N_6847);
xor U18155 (N_18155,N_8139,N_11789);
nor U18156 (N_18156,N_6488,N_8729);
and U18157 (N_18157,N_8433,N_8350);
nand U18158 (N_18158,N_10447,N_9925);
nor U18159 (N_18159,N_8159,N_10963);
or U18160 (N_18160,N_9335,N_9115);
and U18161 (N_18161,N_10975,N_9280);
and U18162 (N_18162,N_8606,N_9545);
xor U18163 (N_18163,N_6979,N_9440);
nand U18164 (N_18164,N_7157,N_11572);
nor U18165 (N_18165,N_9841,N_7099);
nand U18166 (N_18166,N_9882,N_9822);
or U18167 (N_18167,N_10877,N_11116);
nor U18168 (N_18168,N_10178,N_8611);
and U18169 (N_18169,N_11241,N_6878);
or U18170 (N_18170,N_9092,N_10908);
and U18171 (N_18171,N_9155,N_9881);
xnor U18172 (N_18172,N_10869,N_8739);
and U18173 (N_18173,N_6416,N_8586);
nand U18174 (N_18174,N_7555,N_6829);
nand U18175 (N_18175,N_11701,N_7222);
and U18176 (N_18176,N_9416,N_11537);
xor U18177 (N_18177,N_11908,N_9107);
xor U18178 (N_18178,N_7426,N_10318);
xor U18179 (N_18179,N_7207,N_12369);
and U18180 (N_18180,N_11583,N_7215);
xnor U18181 (N_18181,N_11443,N_8393);
nand U18182 (N_18182,N_7065,N_7232);
or U18183 (N_18183,N_6314,N_8327);
or U18184 (N_18184,N_11417,N_10425);
nor U18185 (N_18185,N_10465,N_11223);
xnor U18186 (N_18186,N_7004,N_10111);
nand U18187 (N_18187,N_6570,N_8945);
nand U18188 (N_18188,N_11351,N_9077);
and U18189 (N_18189,N_9559,N_6515);
nor U18190 (N_18190,N_9596,N_8054);
and U18191 (N_18191,N_9769,N_9679);
nor U18192 (N_18192,N_10466,N_7733);
or U18193 (N_18193,N_9332,N_11175);
nand U18194 (N_18194,N_9571,N_6896);
or U18195 (N_18195,N_7671,N_11655);
and U18196 (N_18196,N_11308,N_7030);
nand U18197 (N_18197,N_6543,N_10055);
xor U18198 (N_18198,N_8812,N_11703);
nor U18199 (N_18199,N_7443,N_8248);
or U18200 (N_18200,N_10930,N_10654);
nor U18201 (N_18201,N_11238,N_11796);
and U18202 (N_18202,N_11285,N_12294);
and U18203 (N_18203,N_6306,N_8189);
or U18204 (N_18204,N_6848,N_7804);
or U18205 (N_18205,N_8100,N_11129);
or U18206 (N_18206,N_12221,N_11747);
or U18207 (N_18207,N_12397,N_9439);
nor U18208 (N_18208,N_12209,N_9878);
xor U18209 (N_18209,N_11818,N_12283);
nand U18210 (N_18210,N_10626,N_8501);
nand U18211 (N_18211,N_9816,N_9802);
nor U18212 (N_18212,N_8941,N_8950);
xnor U18213 (N_18213,N_10456,N_10272);
and U18214 (N_18214,N_8916,N_10972);
or U18215 (N_18215,N_6299,N_10623);
nor U18216 (N_18216,N_7032,N_7924);
xnor U18217 (N_18217,N_8208,N_10944);
nor U18218 (N_18218,N_9932,N_11980);
nand U18219 (N_18219,N_12217,N_9564);
xor U18220 (N_18220,N_11387,N_7838);
or U18221 (N_18221,N_7343,N_8441);
nor U18222 (N_18222,N_8647,N_9919);
and U18223 (N_18223,N_9749,N_6959);
or U18224 (N_18224,N_9152,N_8894);
and U18225 (N_18225,N_11410,N_6393);
or U18226 (N_18226,N_10309,N_6983);
or U18227 (N_18227,N_7139,N_7004);
nand U18228 (N_18228,N_10387,N_7903);
nor U18229 (N_18229,N_10142,N_7422);
and U18230 (N_18230,N_7790,N_9823);
or U18231 (N_18231,N_9280,N_6323);
or U18232 (N_18232,N_10411,N_10395);
nor U18233 (N_18233,N_10235,N_7688);
and U18234 (N_18234,N_10730,N_6619);
xor U18235 (N_18235,N_9562,N_6765);
nand U18236 (N_18236,N_9908,N_9848);
or U18237 (N_18237,N_8302,N_10570);
nor U18238 (N_18238,N_8386,N_11522);
or U18239 (N_18239,N_12353,N_9874);
nor U18240 (N_18240,N_8755,N_8944);
and U18241 (N_18241,N_7078,N_6940);
and U18242 (N_18242,N_8796,N_10583);
and U18243 (N_18243,N_11649,N_9743);
or U18244 (N_18244,N_9974,N_11449);
and U18245 (N_18245,N_12391,N_9149);
or U18246 (N_18246,N_11182,N_6447);
or U18247 (N_18247,N_12065,N_9365);
xnor U18248 (N_18248,N_12387,N_9617);
or U18249 (N_18249,N_9795,N_9722);
nor U18250 (N_18250,N_11150,N_9630);
or U18251 (N_18251,N_6634,N_10867);
nand U18252 (N_18252,N_8990,N_11273);
and U18253 (N_18253,N_8357,N_12006);
xor U18254 (N_18254,N_8907,N_7780);
or U18255 (N_18255,N_7737,N_6704);
nand U18256 (N_18256,N_9693,N_7428);
nand U18257 (N_18257,N_10971,N_10581);
and U18258 (N_18258,N_7803,N_10315);
and U18259 (N_18259,N_6380,N_9890);
xor U18260 (N_18260,N_6705,N_10448);
nand U18261 (N_18261,N_8412,N_8219);
xnor U18262 (N_18262,N_11953,N_10743);
or U18263 (N_18263,N_7098,N_11928);
nor U18264 (N_18264,N_6395,N_9026);
nand U18265 (N_18265,N_8014,N_9754);
nand U18266 (N_18266,N_11456,N_7969);
nor U18267 (N_18267,N_9978,N_7792);
nand U18268 (N_18268,N_8960,N_7603);
and U18269 (N_18269,N_9769,N_10462);
nand U18270 (N_18270,N_10428,N_7174);
nor U18271 (N_18271,N_11232,N_9441);
nor U18272 (N_18272,N_9472,N_8155);
nand U18273 (N_18273,N_9485,N_12289);
or U18274 (N_18274,N_6406,N_11831);
nand U18275 (N_18275,N_8070,N_10996);
nand U18276 (N_18276,N_10836,N_12177);
nand U18277 (N_18277,N_11738,N_10574);
or U18278 (N_18278,N_9795,N_10223);
nand U18279 (N_18279,N_11326,N_11371);
and U18280 (N_18280,N_6612,N_11506);
xor U18281 (N_18281,N_7650,N_9754);
nor U18282 (N_18282,N_10872,N_9848);
and U18283 (N_18283,N_9581,N_11898);
xor U18284 (N_18284,N_6488,N_10080);
and U18285 (N_18285,N_11157,N_8438);
nor U18286 (N_18286,N_12016,N_11023);
xor U18287 (N_18287,N_9875,N_10697);
nand U18288 (N_18288,N_12173,N_8678);
nor U18289 (N_18289,N_11316,N_12387);
nand U18290 (N_18290,N_10395,N_9836);
xnor U18291 (N_18291,N_8472,N_10461);
or U18292 (N_18292,N_8505,N_10583);
nor U18293 (N_18293,N_8621,N_12437);
xnor U18294 (N_18294,N_9724,N_7084);
nand U18295 (N_18295,N_10140,N_10398);
nand U18296 (N_18296,N_10899,N_12361);
nand U18297 (N_18297,N_8614,N_7125);
xnor U18298 (N_18298,N_10868,N_7191);
nand U18299 (N_18299,N_8853,N_11569);
nor U18300 (N_18300,N_11631,N_9151);
nand U18301 (N_18301,N_11047,N_10120);
and U18302 (N_18302,N_10482,N_6290);
and U18303 (N_18303,N_12485,N_10783);
or U18304 (N_18304,N_8660,N_8328);
nor U18305 (N_18305,N_11390,N_11370);
nor U18306 (N_18306,N_12441,N_10893);
xnor U18307 (N_18307,N_7641,N_8004);
and U18308 (N_18308,N_6641,N_9090);
nand U18309 (N_18309,N_6552,N_9333);
nor U18310 (N_18310,N_8751,N_11404);
nor U18311 (N_18311,N_12264,N_6384);
or U18312 (N_18312,N_12439,N_10155);
xor U18313 (N_18313,N_12150,N_10955);
nand U18314 (N_18314,N_7361,N_10240);
nand U18315 (N_18315,N_8966,N_12163);
nor U18316 (N_18316,N_10987,N_11308);
or U18317 (N_18317,N_9359,N_12055);
and U18318 (N_18318,N_7055,N_10702);
nor U18319 (N_18319,N_6336,N_9314);
or U18320 (N_18320,N_6787,N_8680);
or U18321 (N_18321,N_6463,N_6911);
xor U18322 (N_18322,N_9441,N_9083);
nand U18323 (N_18323,N_10214,N_9407);
and U18324 (N_18324,N_7969,N_9542);
nor U18325 (N_18325,N_8183,N_6871);
nand U18326 (N_18326,N_8396,N_10934);
or U18327 (N_18327,N_6690,N_11360);
nand U18328 (N_18328,N_6406,N_8551);
nor U18329 (N_18329,N_9424,N_7129);
nor U18330 (N_18330,N_12477,N_11788);
and U18331 (N_18331,N_7123,N_6465);
nor U18332 (N_18332,N_7343,N_6970);
and U18333 (N_18333,N_6863,N_11261);
and U18334 (N_18334,N_6882,N_11503);
nand U18335 (N_18335,N_11319,N_11130);
nand U18336 (N_18336,N_7211,N_10158);
xor U18337 (N_18337,N_10198,N_8860);
or U18338 (N_18338,N_11382,N_10596);
and U18339 (N_18339,N_11411,N_7654);
nor U18340 (N_18340,N_10723,N_9122);
or U18341 (N_18341,N_8946,N_6395);
nand U18342 (N_18342,N_8254,N_6440);
and U18343 (N_18343,N_7758,N_7899);
nor U18344 (N_18344,N_8971,N_10136);
or U18345 (N_18345,N_6872,N_6672);
nor U18346 (N_18346,N_11800,N_10919);
xor U18347 (N_18347,N_12418,N_11184);
xnor U18348 (N_18348,N_10576,N_12042);
or U18349 (N_18349,N_6278,N_8874);
and U18350 (N_18350,N_9987,N_6396);
nor U18351 (N_18351,N_6597,N_6937);
or U18352 (N_18352,N_9942,N_11106);
and U18353 (N_18353,N_10937,N_11629);
nand U18354 (N_18354,N_8227,N_7362);
nand U18355 (N_18355,N_8852,N_6361);
nand U18356 (N_18356,N_9271,N_10646);
nor U18357 (N_18357,N_10237,N_12434);
and U18358 (N_18358,N_7947,N_7349);
nor U18359 (N_18359,N_11717,N_6787);
and U18360 (N_18360,N_7247,N_8307);
and U18361 (N_18361,N_6595,N_12377);
nand U18362 (N_18362,N_8525,N_6948);
or U18363 (N_18363,N_8063,N_9757);
and U18364 (N_18364,N_11405,N_7662);
nor U18365 (N_18365,N_6677,N_7725);
nor U18366 (N_18366,N_6372,N_8796);
or U18367 (N_18367,N_11479,N_10585);
nor U18368 (N_18368,N_11062,N_10089);
and U18369 (N_18369,N_9811,N_10938);
and U18370 (N_18370,N_10417,N_11495);
and U18371 (N_18371,N_6741,N_8439);
nand U18372 (N_18372,N_6250,N_10357);
nor U18373 (N_18373,N_9271,N_6801);
or U18374 (N_18374,N_7598,N_6864);
nor U18375 (N_18375,N_6363,N_11915);
and U18376 (N_18376,N_7548,N_11585);
nand U18377 (N_18377,N_10860,N_9649);
nor U18378 (N_18378,N_8893,N_9604);
nor U18379 (N_18379,N_9339,N_10914);
or U18380 (N_18380,N_8736,N_10480);
and U18381 (N_18381,N_7893,N_10018);
nor U18382 (N_18382,N_10379,N_9700);
nor U18383 (N_18383,N_10510,N_8207);
or U18384 (N_18384,N_11181,N_9072);
and U18385 (N_18385,N_12242,N_7950);
nand U18386 (N_18386,N_10768,N_8422);
or U18387 (N_18387,N_7176,N_8019);
and U18388 (N_18388,N_10848,N_10444);
or U18389 (N_18389,N_7191,N_10698);
or U18390 (N_18390,N_7720,N_10406);
and U18391 (N_18391,N_8331,N_7336);
nand U18392 (N_18392,N_7096,N_12035);
and U18393 (N_18393,N_8621,N_7065);
nor U18394 (N_18394,N_12276,N_8569);
nor U18395 (N_18395,N_7517,N_11042);
nor U18396 (N_18396,N_8268,N_8136);
or U18397 (N_18397,N_12106,N_8011);
or U18398 (N_18398,N_9935,N_7023);
nand U18399 (N_18399,N_6371,N_7368);
nand U18400 (N_18400,N_12408,N_8035);
nor U18401 (N_18401,N_7074,N_10876);
or U18402 (N_18402,N_11213,N_6564);
and U18403 (N_18403,N_8712,N_8622);
nor U18404 (N_18404,N_6969,N_6412);
or U18405 (N_18405,N_6722,N_8178);
nor U18406 (N_18406,N_7972,N_9236);
or U18407 (N_18407,N_11674,N_10388);
nand U18408 (N_18408,N_7595,N_6928);
nor U18409 (N_18409,N_10321,N_12010);
or U18410 (N_18410,N_8366,N_7327);
xnor U18411 (N_18411,N_7207,N_10624);
and U18412 (N_18412,N_8783,N_11866);
and U18413 (N_18413,N_6628,N_8837);
or U18414 (N_18414,N_7677,N_9492);
or U18415 (N_18415,N_10239,N_10689);
and U18416 (N_18416,N_9758,N_10244);
xnor U18417 (N_18417,N_10388,N_12085);
or U18418 (N_18418,N_10981,N_9737);
nand U18419 (N_18419,N_9288,N_12335);
xor U18420 (N_18420,N_11185,N_9865);
or U18421 (N_18421,N_8774,N_8495);
and U18422 (N_18422,N_11314,N_6579);
nand U18423 (N_18423,N_10829,N_7768);
and U18424 (N_18424,N_6537,N_7821);
or U18425 (N_18425,N_6801,N_10500);
nor U18426 (N_18426,N_11179,N_6563);
nor U18427 (N_18427,N_8201,N_7190);
nand U18428 (N_18428,N_10434,N_9027);
nand U18429 (N_18429,N_9119,N_10907);
nand U18430 (N_18430,N_7797,N_7660);
and U18431 (N_18431,N_8434,N_8478);
xnor U18432 (N_18432,N_11316,N_6922);
nor U18433 (N_18433,N_11101,N_8562);
xnor U18434 (N_18434,N_11861,N_12092);
and U18435 (N_18435,N_7612,N_10983);
nor U18436 (N_18436,N_9400,N_9809);
nand U18437 (N_18437,N_9029,N_7939);
or U18438 (N_18438,N_7131,N_7312);
nand U18439 (N_18439,N_11409,N_12183);
xor U18440 (N_18440,N_6373,N_7189);
xor U18441 (N_18441,N_9430,N_10192);
nor U18442 (N_18442,N_8768,N_11809);
or U18443 (N_18443,N_9861,N_9804);
nand U18444 (N_18444,N_11260,N_8830);
and U18445 (N_18445,N_10743,N_7421);
or U18446 (N_18446,N_6387,N_11590);
and U18447 (N_18447,N_10269,N_11286);
nand U18448 (N_18448,N_9103,N_7714);
nor U18449 (N_18449,N_6881,N_8104);
nor U18450 (N_18450,N_6688,N_10808);
xnor U18451 (N_18451,N_11645,N_8163);
or U18452 (N_18452,N_9714,N_8219);
and U18453 (N_18453,N_6660,N_11770);
or U18454 (N_18454,N_7658,N_10660);
or U18455 (N_18455,N_11334,N_11877);
or U18456 (N_18456,N_7544,N_6291);
nand U18457 (N_18457,N_12459,N_7365);
nor U18458 (N_18458,N_9632,N_8440);
nand U18459 (N_18459,N_11209,N_8502);
or U18460 (N_18460,N_6572,N_9144);
and U18461 (N_18461,N_10646,N_9635);
or U18462 (N_18462,N_7249,N_8694);
nor U18463 (N_18463,N_10084,N_10789);
or U18464 (N_18464,N_11409,N_11940);
or U18465 (N_18465,N_8696,N_6688);
xor U18466 (N_18466,N_8481,N_9645);
nand U18467 (N_18467,N_10164,N_8451);
nand U18468 (N_18468,N_10099,N_8366);
or U18469 (N_18469,N_11764,N_8249);
xor U18470 (N_18470,N_12083,N_10971);
or U18471 (N_18471,N_8679,N_7883);
and U18472 (N_18472,N_7214,N_9886);
and U18473 (N_18473,N_10522,N_9504);
or U18474 (N_18474,N_7044,N_7677);
or U18475 (N_18475,N_11361,N_12038);
nor U18476 (N_18476,N_9498,N_9994);
nor U18477 (N_18477,N_12300,N_8632);
and U18478 (N_18478,N_11178,N_7104);
and U18479 (N_18479,N_11536,N_7290);
or U18480 (N_18480,N_10188,N_11132);
and U18481 (N_18481,N_8464,N_9521);
nor U18482 (N_18482,N_7003,N_9622);
xor U18483 (N_18483,N_11775,N_7673);
nand U18484 (N_18484,N_8324,N_10532);
or U18485 (N_18485,N_9917,N_9692);
nor U18486 (N_18486,N_9643,N_10690);
nor U18487 (N_18487,N_10939,N_6502);
nor U18488 (N_18488,N_10115,N_6359);
xnor U18489 (N_18489,N_8932,N_12465);
and U18490 (N_18490,N_7027,N_12023);
or U18491 (N_18491,N_7019,N_9314);
and U18492 (N_18492,N_8405,N_12483);
nand U18493 (N_18493,N_10617,N_7005);
nand U18494 (N_18494,N_9717,N_11183);
nand U18495 (N_18495,N_7693,N_10679);
nor U18496 (N_18496,N_10270,N_7527);
and U18497 (N_18497,N_7181,N_8262);
and U18498 (N_18498,N_10241,N_9305);
or U18499 (N_18499,N_7961,N_9685);
nor U18500 (N_18500,N_7991,N_8702);
and U18501 (N_18501,N_10209,N_12402);
and U18502 (N_18502,N_10742,N_7106);
xor U18503 (N_18503,N_8123,N_9357);
nor U18504 (N_18504,N_9846,N_8566);
nor U18505 (N_18505,N_7418,N_12255);
nor U18506 (N_18506,N_10209,N_7009);
and U18507 (N_18507,N_7575,N_7130);
xor U18508 (N_18508,N_7036,N_6707);
nor U18509 (N_18509,N_10959,N_8306);
nor U18510 (N_18510,N_6377,N_10711);
xor U18511 (N_18511,N_10377,N_9705);
nand U18512 (N_18512,N_12283,N_8405);
and U18513 (N_18513,N_11639,N_7743);
or U18514 (N_18514,N_10429,N_9848);
nand U18515 (N_18515,N_6527,N_10371);
nand U18516 (N_18516,N_10394,N_8780);
and U18517 (N_18517,N_7443,N_11561);
nor U18518 (N_18518,N_6793,N_7089);
nand U18519 (N_18519,N_6830,N_7531);
nand U18520 (N_18520,N_6556,N_8725);
nor U18521 (N_18521,N_7240,N_10174);
and U18522 (N_18522,N_6889,N_9038);
nand U18523 (N_18523,N_9905,N_8908);
nand U18524 (N_18524,N_11550,N_9036);
nand U18525 (N_18525,N_8816,N_9565);
or U18526 (N_18526,N_10942,N_9478);
nand U18527 (N_18527,N_7111,N_6599);
and U18528 (N_18528,N_8928,N_10273);
or U18529 (N_18529,N_7529,N_7610);
or U18530 (N_18530,N_11446,N_10639);
and U18531 (N_18531,N_10265,N_10701);
nor U18532 (N_18532,N_11799,N_8872);
nor U18533 (N_18533,N_6356,N_7727);
nor U18534 (N_18534,N_12455,N_7624);
nand U18535 (N_18535,N_9580,N_12277);
or U18536 (N_18536,N_8951,N_9308);
nand U18537 (N_18537,N_12374,N_8383);
nor U18538 (N_18538,N_6342,N_8607);
or U18539 (N_18539,N_10064,N_10307);
nor U18540 (N_18540,N_6385,N_7686);
or U18541 (N_18541,N_6293,N_9606);
nand U18542 (N_18542,N_6551,N_10410);
or U18543 (N_18543,N_8052,N_11918);
nand U18544 (N_18544,N_9565,N_11401);
nand U18545 (N_18545,N_11022,N_6340);
nor U18546 (N_18546,N_10023,N_9262);
xor U18547 (N_18547,N_7069,N_10458);
xnor U18548 (N_18548,N_10828,N_7199);
nor U18549 (N_18549,N_6535,N_10339);
or U18550 (N_18550,N_7031,N_10002);
nand U18551 (N_18551,N_11503,N_9698);
nand U18552 (N_18552,N_6264,N_8516);
nand U18553 (N_18553,N_6722,N_11188);
nand U18554 (N_18554,N_9235,N_12474);
nor U18555 (N_18555,N_8936,N_12082);
nand U18556 (N_18556,N_10208,N_11263);
nor U18557 (N_18557,N_8336,N_11757);
or U18558 (N_18558,N_6605,N_8125);
nand U18559 (N_18559,N_10324,N_12024);
or U18560 (N_18560,N_6284,N_9361);
nor U18561 (N_18561,N_8402,N_6556);
nor U18562 (N_18562,N_9139,N_6361);
nand U18563 (N_18563,N_6893,N_9095);
and U18564 (N_18564,N_7818,N_8410);
and U18565 (N_18565,N_8231,N_11755);
nor U18566 (N_18566,N_11619,N_7014);
nor U18567 (N_18567,N_7090,N_8768);
nor U18568 (N_18568,N_11068,N_8883);
nand U18569 (N_18569,N_6519,N_9491);
nand U18570 (N_18570,N_10616,N_6360);
nor U18571 (N_18571,N_10606,N_6983);
nand U18572 (N_18572,N_10542,N_9621);
nor U18573 (N_18573,N_7883,N_9574);
nor U18574 (N_18574,N_10818,N_7406);
nor U18575 (N_18575,N_6317,N_7291);
nand U18576 (N_18576,N_7018,N_6525);
and U18577 (N_18577,N_9257,N_10425);
nor U18578 (N_18578,N_8633,N_7120);
nand U18579 (N_18579,N_10124,N_8064);
xnor U18580 (N_18580,N_8900,N_9343);
nor U18581 (N_18581,N_8882,N_6504);
nand U18582 (N_18582,N_6948,N_11447);
nor U18583 (N_18583,N_8977,N_11561);
and U18584 (N_18584,N_11634,N_6451);
xor U18585 (N_18585,N_12473,N_12250);
and U18586 (N_18586,N_7967,N_12345);
xor U18587 (N_18587,N_9379,N_9029);
or U18588 (N_18588,N_9204,N_10887);
and U18589 (N_18589,N_11181,N_9699);
xnor U18590 (N_18590,N_11745,N_11733);
and U18591 (N_18591,N_11363,N_12167);
or U18592 (N_18592,N_8085,N_10390);
xnor U18593 (N_18593,N_10775,N_9645);
xnor U18594 (N_18594,N_8556,N_11596);
nand U18595 (N_18595,N_9814,N_6671);
nor U18596 (N_18596,N_7337,N_10109);
nand U18597 (N_18597,N_11891,N_9911);
and U18598 (N_18598,N_9885,N_7741);
or U18599 (N_18599,N_11660,N_11821);
nor U18600 (N_18600,N_12191,N_12223);
and U18601 (N_18601,N_12287,N_9646);
and U18602 (N_18602,N_11780,N_12290);
nor U18603 (N_18603,N_8538,N_8208);
or U18604 (N_18604,N_7079,N_12485);
nand U18605 (N_18605,N_8571,N_10065);
nor U18606 (N_18606,N_9186,N_10792);
or U18607 (N_18607,N_12321,N_10897);
nand U18608 (N_18608,N_11835,N_7461);
nor U18609 (N_18609,N_9127,N_9478);
or U18610 (N_18610,N_7467,N_11908);
or U18611 (N_18611,N_9292,N_8577);
nand U18612 (N_18612,N_11837,N_6859);
nand U18613 (N_18613,N_11390,N_6942);
nor U18614 (N_18614,N_11813,N_6873);
or U18615 (N_18615,N_11084,N_10720);
and U18616 (N_18616,N_11228,N_10888);
nand U18617 (N_18617,N_12034,N_9077);
nor U18618 (N_18618,N_8605,N_7575);
and U18619 (N_18619,N_12275,N_8495);
and U18620 (N_18620,N_8487,N_7684);
or U18621 (N_18621,N_6519,N_6363);
nand U18622 (N_18622,N_8585,N_9444);
xor U18623 (N_18623,N_11604,N_6698);
and U18624 (N_18624,N_9959,N_7439);
nor U18625 (N_18625,N_8360,N_11913);
or U18626 (N_18626,N_6320,N_12130);
and U18627 (N_18627,N_10191,N_8843);
nand U18628 (N_18628,N_7807,N_6389);
and U18629 (N_18629,N_10554,N_11074);
and U18630 (N_18630,N_8410,N_8023);
or U18631 (N_18631,N_7077,N_8852);
or U18632 (N_18632,N_7232,N_12484);
nand U18633 (N_18633,N_9211,N_8453);
xnor U18634 (N_18634,N_11203,N_7305);
nor U18635 (N_18635,N_6340,N_10880);
nor U18636 (N_18636,N_10026,N_11748);
or U18637 (N_18637,N_8850,N_7929);
and U18638 (N_18638,N_10092,N_10801);
and U18639 (N_18639,N_7214,N_10350);
or U18640 (N_18640,N_8466,N_6609);
nand U18641 (N_18641,N_9983,N_12211);
or U18642 (N_18642,N_8653,N_8792);
and U18643 (N_18643,N_11555,N_7388);
and U18644 (N_18644,N_11484,N_9001);
nor U18645 (N_18645,N_10619,N_9652);
or U18646 (N_18646,N_8545,N_9953);
and U18647 (N_18647,N_8303,N_9494);
nor U18648 (N_18648,N_11537,N_7843);
or U18649 (N_18649,N_10444,N_7649);
or U18650 (N_18650,N_12216,N_8839);
or U18651 (N_18651,N_9312,N_10289);
nor U18652 (N_18652,N_12148,N_11985);
nor U18653 (N_18653,N_6457,N_11317);
nand U18654 (N_18654,N_6675,N_6614);
xnor U18655 (N_18655,N_7847,N_7795);
and U18656 (N_18656,N_11861,N_9848);
nor U18657 (N_18657,N_11723,N_6429);
nand U18658 (N_18658,N_8150,N_10162);
xor U18659 (N_18659,N_12224,N_10890);
and U18660 (N_18660,N_9951,N_8040);
nand U18661 (N_18661,N_11878,N_9468);
or U18662 (N_18662,N_7224,N_6916);
nor U18663 (N_18663,N_6671,N_6318);
or U18664 (N_18664,N_11891,N_7245);
nor U18665 (N_18665,N_9288,N_6867);
and U18666 (N_18666,N_8656,N_7619);
nor U18667 (N_18667,N_6706,N_6677);
nor U18668 (N_18668,N_10964,N_11115);
nand U18669 (N_18669,N_7846,N_6803);
xnor U18670 (N_18670,N_9774,N_7601);
or U18671 (N_18671,N_8536,N_11159);
and U18672 (N_18672,N_9167,N_11399);
xnor U18673 (N_18673,N_7551,N_8624);
xnor U18674 (N_18674,N_6883,N_11052);
or U18675 (N_18675,N_8459,N_10695);
nand U18676 (N_18676,N_12289,N_12026);
or U18677 (N_18677,N_9033,N_6533);
nand U18678 (N_18678,N_6512,N_7671);
and U18679 (N_18679,N_10135,N_9258);
or U18680 (N_18680,N_10835,N_8353);
nor U18681 (N_18681,N_7165,N_10306);
nand U18682 (N_18682,N_10804,N_9705);
and U18683 (N_18683,N_8389,N_7905);
xor U18684 (N_18684,N_11212,N_9070);
and U18685 (N_18685,N_7607,N_8653);
or U18686 (N_18686,N_7637,N_7584);
and U18687 (N_18687,N_7262,N_8821);
and U18688 (N_18688,N_7807,N_9315);
nand U18689 (N_18689,N_10483,N_9411);
or U18690 (N_18690,N_10213,N_10447);
nand U18691 (N_18691,N_11375,N_7046);
xnor U18692 (N_18692,N_6574,N_11042);
nand U18693 (N_18693,N_7897,N_11741);
and U18694 (N_18694,N_11823,N_11848);
or U18695 (N_18695,N_8893,N_6543);
and U18696 (N_18696,N_6903,N_7269);
and U18697 (N_18697,N_9189,N_12438);
and U18698 (N_18698,N_11059,N_6687);
nor U18699 (N_18699,N_8448,N_9579);
xnor U18700 (N_18700,N_9599,N_11854);
or U18701 (N_18701,N_6259,N_9772);
xor U18702 (N_18702,N_11390,N_10628);
nand U18703 (N_18703,N_6558,N_7702);
nor U18704 (N_18704,N_10024,N_10218);
xor U18705 (N_18705,N_8406,N_11459);
nand U18706 (N_18706,N_11641,N_10290);
nand U18707 (N_18707,N_8924,N_6424);
and U18708 (N_18708,N_12249,N_6513);
or U18709 (N_18709,N_11657,N_11827);
or U18710 (N_18710,N_10306,N_9420);
nand U18711 (N_18711,N_12219,N_8727);
nor U18712 (N_18712,N_6487,N_11958);
and U18713 (N_18713,N_9934,N_7938);
nor U18714 (N_18714,N_11160,N_11979);
or U18715 (N_18715,N_9521,N_12361);
nor U18716 (N_18716,N_12075,N_8927);
and U18717 (N_18717,N_7792,N_7733);
or U18718 (N_18718,N_8150,N_10124);
or U18719 (N_18719,N_6738,N_11435);
nor U18720 (N_18720,N_10351,N_11173);
and U18721 (N_18721,N_8469,N_8991);
nor U18722 (N_18722,N_9774,N_7774);
nand U18723 (N_18723,N_6751,N_12318);
xor U18724 (N_18724,N_8388,N_11461);
and U18725 (N_18725,N_11373,N_9999);
and U18726 (N_18726,N_11792,N_7272);
or U18727 (N_18727,N_10283,N_7707);
or U18728 (N_18728,N_7950,N_10345);
or U18729 (N_18729,N_10294,N_12224);
or U18730 (N_18730,N_7933,N_9647);
and U18731 (N_18731,N_9837,N_9332);
nor U18732 (N_18732,N_6257,N_7086);
nand U18733 (N_18733,N_7274,N_8217);
nor U18734 (N_18734,N_10852,N_6776);
nand U18735 (N_18735,N_7731,N_8796);
or U18736 (N_18736,N_11409,N_7867);
and U18737 (N_18737,N_12129,N_7860);
nand U18738 (N_18738,N_11335,N_12413);
or U18739 (N_18739,N_10681,N_11767);
nand U18740 (N_18740,N_9913,N_7274);
nor U18741 (N_18741,N_11610,N_8307);
nand U18742 (N_18742,N_7203,N_10296);
and U18743 (N_18743,N_7910,N_6643);
nand U18744 (N_18744,N_12481,N_8058);
nand U18745 (N_18745,N_10934,N_9903);
or U18746 (N_18746,N_9447,N_11601);
xnor U18747 (N_18747,N_11164,N_6312);
xor U18748 (N_18748,N_8695,N_10058);
nor U18749 (N_18749,N_12326,N_9137);
or U18750 (N_18750,N_13456,N_15546);
nor U18751 (N_18751,N_13671,N_18648);
nor U18752 (N_18752,N_13429,N_14135);
and U18753 (N_18753,N_13954,N_14970);
nor U18754 (N_18754,N_13739,N_16768);
nand U18755 (N_18755,N_13244,N_14964);
and U18756 (N_18756,N_12821,N_17753);
or U18757 (N_18757,N_17624,N_14297);
nand U18758 (N_18758,N_14017,N_16864);
nor U18759 (N_18759,N_17464,N_13310);
and U18760 (N_18760,N_13157,N_18181);
xor U18761 (N_18761,N_14211,N_18348);
or U18762 (N_18762,N_16850,N_15582);
nor U18763 (N_18763,N_17262,N_16669);
nor U18764 (N_18764,N_14436,N_18503);
nand U18765 (N_18765,N_16194,N_17233);
nand U18766 (N_18766,N_17076,N_18469);
or U18767 (N_18767,N_16759,N_17538);
or U18768 (N_18768,N_14468,N_15153);
or U18769 (N_18769,N_13446,N_16448);
nor U18770 (N_18770,N_14856,N_14972);
and U18771 (N_18771,N_15585,N_17007);
and U18772 (N_18772,N_16557,N_17554);
nor U18773 (N_18773,N_14294,N_16829);
or U18774 (N_18774,N_14668,N_17545);
or U18775 (N_18775,N_12730,N_17163);
nor U18776 (N_18776,N_12950,N_16090);
or U18777 (N_18777,N_13442,N_17400);
nand U18778 (N_18778,N_18679,N_18383);
nor U18779 (N_18779,N_18378,N_15513);
nand U18780 (N_18780,N_14681,N_17313);
nand U18781 (N_18781,N_15710,N_17204);
xor U18782 (N_18782,N_13598,N_13184);
nor U18783 (N_18783,N_12788,N_13772);
and U18784 (N_18784,N_16873,N_17973);
nor U18785 (N_18785,N_14346,N_13647);
nor U18786 (N_18786,N_15182,N_15680);
nor U18787 (N_18787,N_17318,N_14005);
xor U18788 (N_18788,N_13232,N_13464);
nand U18789 (N_18789,N_15438,N_13433);
nor U18790 (N_18790,N_18620,N_14612);
nor U18791 (N_18791,N_14875,N_12646);
nor U18792 (N_18792,N_13735,N_18059);
and U18793 (N_18793,N_17169,N_18668);
and U18794 (N_18794,N_17943,N_18377);
or U18795 (N_18795,N_13240,N_12806);
nand U18796 (N_18796,N_12922,N_17458);
xnor U18797 (N_18797,N_17648,N_18542);
xnor U18798 (N_18798,N_18103,N_13057);
and U18799 (N_18799,N_16795,N_18177);
and U18800 (N_18800,N_12863,N_13052);
and U18801 (N_18801,N_15681,N_14307);
and U18802 (N_18802,N_18025,N_13520);
nand U18803 (N_18803,N_12944,N_17911);
nand U18804 (N_18804,N_14826,N_16957);
nand U18805 (N_18805,N_18399,N_16776);
nor U18806 (N_18806,N_14166,N_17472);
xor U18807 (N_18807,N_13821,N_16104);
nand U18808 (N_18808,N_13907,N_18747);
nand U18809 (N_18809,N_16345,N_16322);
xnor U18810 (N_18810,N_18360,N_13952);
and U18811 (N_18811,N_15693,N_14852);
nand U18812 (N_18812,N_17328,N_17178);
nand U18813 (N_18813,N_18288,N_16545);
nand U18814 (N_18814,N_14165,N_16998);
or U18815 (N_18815,N_14953,N_14778);
nor U18816 (N_18816,N_13006,N_15008);
nor U18817 (N_18817,N_13131,N_18601);
or U18818 (N_18818,N_18621,N_15672);
xor U18819 (N_18819,N_13694,N_12770);
and U18820 (N_18820,N_15951,N_17218);
or U18821 (N_18821,N_18168,N_14072);
and U18822 (N_18822,N_15524,N_14999);
or U18823 (N_18823,N_18568,N_15066);
or U18824 (N_18824,N_17131,N_18258);
nand U18825 (N_18825,N_17798,N_13391);
and U18826 (N_18826,N_14935,N_14322);
and U18827 (N_18827,N_17626,N_17587);
nand U18828 (N_18828,N_13769,N_13067);
nand U18829 (N_18829,N_14115,N_12832);
and U18830 (N_18830,N_18211,N_12514);
nand U18831 (N_18831,N_14305,N_16696);
and U18832 (N_18832,N_15236,N_17620);
or U18833 (N_18833,N_16835,N_17424);
nor U18834 (N_18834,N_17055,N_13030);
nor U18835 (N_18835,N_13040,N_18627);
and U18836 (N_18836,N_18556,N_15692);
xor U18837 (N_18837,N_16456,N_14537);
nand U18838 (N_18838,N_12562,N_13750);
nor U18839 (N_18839,N_16547,N_16543);
and U18840 (N_18840,N_15092,N_18604);
nand U18841 (N_18841,N_13373,N_17170);
or U18842 (N_18842,N_17580,N_12621);
nand U18843 (N_18843,N_17572,N_17980);
nand U18844 (N_18844,N_13675,N_15905);
nor U18845 (N_18845,N_14960,N_16906);
nor U18846 (N_18846,N_17738,N_12535);
and U18847 (N_18847,N_18657,N_14950);
or U18848 (N_18848,N_13225,N_16130);
and U18849 (N_18849,N_15103,N_14860);
and U18850 (N_18850,N_18241,N_16180);
nor U18851 (N_18851,N_12977,N_17921);
and U18852 (N_18852,N_13210,N_16990);
nand U18853 (N_18853,N_13121,N_13970);
and U18854 (N_18854,N_12726,N_12777);
nor U18855 (N_18855,N_14541,N_17718);
nor U18856 (N_18856,N_15992,N_13602);
nor U18857 (N_18857,N_18460,N_12751);
or U18858 (N_18858,N_14576,N_13689);
nand U18859 (N_18859,N_17503,N_16184);
or U18860 (N_18860,N_16647,N_12901);
or U18861 (N_18861,N_13323,N_16117);
nor U18862 (N_18862,N_18151,N_16783);
and U18863 (N_18863,N_15673,N_18057);
or U18864 (N_18864,N_16828,N_18479);
xor U18865 (N_18865,N_13020,N_18401);
nand U18866 (N_18866,N_17286,N_12874);
xnor U18867 (N_18867,N_16955,N_15645);
and U18868 (N_18868,N_13820,N_17792);
nand U18869 (N_18869,N_17008,N_14223);
nand U18870 (N_18870,N_13175,N_17717);
xor U18871 (N_18871,N_15306,N_14405);
nor U18872 (N_18872,N_16763,N_14507);
nand U18873 (N_18873,N_18036,N_18087);
nand U18874 (N_18874,N_17110,N_15535);
or U18875 (N_18875,N_15715,N_18565);
and U18876 (N_18876,N_16132,N_16659);
or U18877 (N_18877,N_17404,N_12866);
nand U18878 (N_18878,N_14736,N_16211);
or U18879 (N_18879,N_12787,N_12558);
and U18880 (N_18880,N_13214,N_16351);
or U18881 (N_18881,N_18131,N_13793);
or U18882 (N_18882,N_13130,N_17579);
nand U18883 (N_18883,N_15572,N_14470);
nand U18884 (N_18884,N_14367,N_17230);
or U18885 (N_18885,N_17202,N_16907);
and U18886 (N_18886,N_16409,N_16642);
nor U18887 (N_18887,N_18016,N_15067);
and U18888 (N_18888,N_16625,N_18563);
nor U18889 (N_18889,N_13123,N_12830);
or U18890 (N_18890,N_12500,N_17302);
nor U18891 (N_18891,N_16773,N_12639);
or U18892 (N_18892,N_14989,N_16366);
or U18893 (N_18893,N_13438,N_16931);
and U18894 (N_18894,N_13742,N_13036);
and U18895 (N_18895,N_14800,N_17126);
or U18896 (N_18896,N_13447,N_15938);
xnor U18897 (N_18897,N_16865,N_13218);
nand U18898 (N_18898,N_14861,N_14694);
and U18899 (N_18899,N_16526,N_17461);
nand U18900 (N_18900,N_13805,N_15638);
or U18901 (N_18901,N_13008,N_17395);
and U18902 (N_18902,N_15144,N_15317);
and U18903 (N_18903,N_15140,N_18380);
nor U18904 (N_18904,N_14228,N_16400);
and U18905 (N_18905,N_16886,N_15360);
nor U18906 (N_18906,N_17097,N_13297);
nand U18907 (N_18907,N_15191,N_14256);
or U18908 (N_18908,N_15525,N_17460);
nand U18909 (N_18909,N_16534,N_14081);
and U18910 (N_18910,N_15705,N_16286);
and U18911 (N_18911,N_14476,N_14579);
xnor U18912 (N_18912,N_16633,N_17242);
nand U18913 (N_18913,N_15800,N_15313);
nand U18914 (N_18914,N_16247,N_18375);
nand U18915 (N_18915,N_18649,N_12587);
or U18916 (N_18916,N_17037,N_12900);
nand U18917 (N_18917,N_15217,N_16272);
or U18918 (N_18918,N_17432,N_18420);
or U18919 (N_18919,N_17625,N_13001);
nor U18920 (N_18920,N_15735,N_12841);
nor U18921 (N_18921,N_14233,N_13737);
or U18922 (N_18922,N_15012,N_14885);
and U18923 (N_18923,N_15519,N_17933);
or U18924 (N_18924,N_13824,N_18743);
and U18925 (N_18925,N_15377,N_17951);
nand U18926 (N_18926,N_17031,N_15965);
and U18927 (N_18927,N_16606,N_12610);
nand U18928 (N_18928,N_17952,N_14142);
nand U18929 (N_18929,N_16772,N_16672);
nand U18930 (N_18930,N_12843,N_12810);
nand U18931 (N_18931,N_15199,N_16922);
or U18932 (N_18932,N_13510,N_15979);
or U18933 (N_18933,N_16600,N_13029);
nor U18934 (N_18934,N_13435,N_14685);
and U18935 (N_18935,N_13364,N_14383);
and U18936 (N_18936,N_18163,N_15192);
nand U18937 (N_18937,N_15070,N_13181);
and U18938 (N_18938,N_17357,N_14409);
nand U18939 (N_18939,N_13807,N_18736);
nand U18940 (N_18940,N_15810,N_13081);
and U18941 (N_18941,N_13691,N_12741);
nor U18942 (N_18942,N_17489,N_16452);
and U18943 (N_18943,N_16686,N_15826);
nand U18944 (N_18944,N_18090,N_13745);
or U18945 (N_18945,N_13738,N_15210);
nand U18946 (N_18946,N_16649,N_18662);
or U18947 (N_18947,N_17713,N_14869);
or U18948 (N_18948,N_13579,N_14615);
nand U18949 (N_18949,N_12601,N_17253);
nand U18950 (N_18950,N_17012,N_13055);
nor U18951 (N_18951,N_18693,N_18699);
nor U18952 (N_18952,N_16479,N_14190);
or U18953 (N_18953,N_17750,N_14114);
and U18954 (N_18954,N_15508,N_15180);
and U18955 (N_18955,N_13427,N_16116);
and U18956 (N_18956,N_16439,N_17878);
or U18957 (N_18957,N_12973,N_13555);
nor U18958 (N_18958,N_14969,N_17695);
and U18959 (N_18959,N_16435,N_13904);
nand U18960 (N_18960,N_18523,N_18101);
nand U18961 (N_18961,N_16170,N_14345);
nand U18962 (N_18962,N_18382,N_14203);
or U18963 (N_18963,N_17238,N_13116);
nand U18964 (N_18964,N_16142,N_15606);
xor U18965 (N_18965,N_14168,N_17142);
nor U18966 (N_18966,N_14111,N_12573);
nand U18967 (N_18967,N_13448,N_14110);
nand U18968 (N_18968,N_16205,N_14762);
nand U18969 (N_18969,N_16831,N_17497);
or U18970 (N_18970,N_14557,N_15728);
and U18971 (N_18971,N_15036,N_15166);
or U18972 (N_18972,N_15806,N_16332);
and U18973 (N_18973,N_16958,N_12755);
and U18974 (N_18974,N_17824,N_15427);
or U18975 (N_18975,N_14451,N_12765);
and U18976 (N_18976,N_15514,N_18157);
nor U18977 (N_18977,N_14770,N_13919);
and U18978 (N_18978,N_12820,N_18226);
xor U18979 (N_18979,N_13961,N_17985);
nand U18980 (N_18980,N_16294,N_15481);
and U18981 (N_18981,N_14318,N_12749);
or U18982 (N_18982,N_18642,N_17562);
or U18983 (N_18983,N_14855,N_14899);
or U18984 (N_18984,N_12642,N_15075);
nand U18985 (N_18985,N_14439,N_16326);
and U18986 (N_18986,N_13000,N_14518);
or U18987 (N_18987,N_18189,N_14487);
nand U18988 (N_18988,N_16623,N_16089);
and U18989 (N_18989,N_18314,N_14026);
nor U18990 (N_18990,N_16373,N_13329);
and U18991 (N_18991,N_14289,N_16268);
or U18992 (N_18992,N_15696,N_12694);
and U18993 (N_18993,N_17616,N_17035);
nor U18994 (N_18994,N_15338,N_13632);
xor U18995 (N_18995,N_17439,N_18456);
and U18996 (N_18996,N_15471,N_14582);
and U18997 (N_18997,N_17449,N_12551);
or U18998 (N_18998,N_14455,N_15505);
nand U18999 (N_18999,N_15213,N_14786);
nor U19000 (N_19000,N_17108,N_16925);
xnor U19001 (N_19001,N_15386,N_14123);
nand U19002 (N_19002,N_16058,N_12933);
nand U19003 (N_19003,N_13636,N_18242);
nand U19004 (N_19004,N_15613,N_17231);
xnor U19005 (N_19005,N_13452,N_17467);
or U19006 (N_19006,N_16393,N_12989);
and U19007 (N_19007,N_13193,N_15867);
or U19008 (N_19008,N_17276,N_18345);
and U19009 (N_19009,N_16472,N_14335);
xor U19010 (N_19010,N_15850,N_15375);
or U19011 (N_19011,N_14535,N_14325);
nand U19012 (N_19012,N_15296,N_14659);
and U19013 (N_19013,N_18678,N_17285);
or U19014 (N_19014,N_15455,N_14027);
nand U19015 (N_19015,N_17950,N_15456);
nand U19016 (N_19016,N_16960,N_13279);
nand U19017 (N_19017,N_13562,N_17398);
nand U19018 (N_19018,N_17466,N_17329);
and U19019 (N_19019,N_16410,N_14914);
or U19020 (N_19020,N_15972,N_13440);
nor U19021 (N_19021,N_13237,N_15004);
nor U19022 (N_19022,N_18472,N_14750);
and U19023 (N_19023,N_13565,N_16640);
and U19024 (N_19024,N_15077,N_16370);
and U19025 (N_19025,N_17589,N_14365);
nand U19026 (N_19026,N_14236,N_16348);
nand U19027 (N_19027,N_15526,N_14699);
or U19028 (N_19028,N_16018,N_14744);
and U19029 (N_19029,N_17160,N_16317);
nand U19030 (N_19030,N_18173,N_12555);
and U19031 (N_19031,N_14174,N_14978);
and U19032 (N_19032,N_15350,N_17038);
nand U19033 (N_19033,N_16022,N_13744);
nor U19034 (N_19034,N_16983,N_15176);
nand U19035 (N_19035,N_12892,N_13226);
and U19036 (N_19036,N_14196,N_15043);
nand U19037 (N_19037,N_17528,N_13953);
and U19038 (N_19038,N_13450,N_16807);
and U19039 (N_19039,N_14908,N_18712);
nand U19040 (N_19040,N_16114,N_18525);
nand U19041 (N_19041,N_14632,N_15409);
and U19042 (N_19042,N_15579,N_13345);
or U19043 (N_19043,N_15968,N_12699);
nand U19044 (N_19044,N_16401,N_17598);
or U19045 (N_19045,N_16385,N_18408);
and U19046 (N_19046,N_15532,N_13019);
nor U19047 (N_19047,N_17105,N_13665);
or U19048 (N_19048,N_18133,N_14814);
or U19049 (N_19049,N_17984,N_14783);
and U19050 (N_19050,N_18144,N_15963);
xnor U19051 (N_19051,N_18078,N_13731);
or U19052 (N_19052,N_16542,N_13822);
nor U19053 (N_19053,N_14520,N_13037);
or U19054 (N_19054,N_13120,N_14274);
and U19055 (N_19055,N_17557,N_16398);
nand U19056 (N_19056,N_16597,N_16586);
nor U19057 (N_19057,N_16263,N_16487);
nor U19058 (N_19058,N_14387,N_18441);
or U19059 (N_19059,N_13944,N_14946);
or U19060 (N_19060,N_17189,N_13327);
or U19061 (N_19061,N_16668,N_12630);
nor U19062 (N_19062,N_16037,N_14245);
and U19063 (N_19063,N_16858,N_12873);
or U19064 (N_19064,N_14868,N_17474);
nand U19065 (N_19065,N_16863,N_13563);
nor U19066 (N_19066,N_18310,N_17867);
nand U19067 (N_19067,N_13927,N_13467);
and U19068 (N_19068,N_18160,N_17061);
nand U19069 (N_19069,N_18607,N_18582);
nand U19070 (N_19070,N_14059,N_18710);
xor U19071 (N_19071,N_14572,N_14639);
nor U19072 (N_19072,N_17645,N_17471);
or U19073 (N_19073,N_18416,N_16650);
nor U19074 (N_19074,N_13716,N_13615);
nand U19075 (N_19075,N_16391,N_18511);
nor U19076 (N_19076,N_13150,N_17124);
and U19077 (N_19077,N_16518,N_17021);
or U19078 (N_19078,N_13233,N_16723);
nand U19079 (N_19079,N_13153,N_12693);
nor U19080 (N_19080,N_16742,N_14870);
nor U19081 (N_19081,N_14737,N_17348);
nor U19082 (N_19082,N_15602,N_15847);
and U19083 (N_19083,N_14392,N_14317);
xnor U19084 (N_19084,N_18120,N_18319);
nor U19085 (N_19085,N_18706,N_17327);
or U19086 (N_19086,N_17307,N_12522);
or U19087 (N_19087,N_13287,N_16025);
or U19088 (N_19088,N_16760,N_14850);
or U19089 (N_19089,N_14082,N_12794);
nor U19090 (N_19090,N_14377,N_17200);
and U19091 (N_19091,N_15405,N_14272);
nor U19092 (N_19092,N_17090,N_15171);
or U19093 (N_19093,N_13867,N_16564);
or U19094 (N_19094,N_13347,N_16706);
nor U19095 (N_19095,N_15124,N_16971);
and U19096 (N_19096,N_13227,N_17071);
and U19097 (N_19097,N_15913,N_15614);
or U19098 (N_19098,N_13418,N_17212);
nor U19099 (N_19099,N_15742,N_15984);
nor U19100 (N_19100,N_17425,N_18749);
and U19101 (N_19101,N_16530,N_18577);
xor U19102 (N_19102,N_16793,N_18448);
and U19103 (N_19103,N_12860,N_16525);
or U19104 (N_19104,N_14382,N_16019);
xnor U19105 (N_19105,N_14074,N_17185);
nand U19106 (N_19106,N_14430,N_15644);
xnor U19107 (N_19107,N_17759,N_13158);
or U19108 (N_19108,N_16897,N_17550);
nand U19109 (N_19109,N_17801,N_16368);
or U19110 (N_19110,N_14492,N_16535);
and U19111 (N_19111,N_16929,N_13882);
or U19112 (N_19112,N_15621,N_14633);
and U19113 (N_19113,N_18427,N_14255);
or U19114 (N_19114,N_16698,N_14480);
and U19115 (N_19115,N_17455,N_14414);
and U19116 (N_19116,N_18017,N_17186);
nor U19117 (N_19117,N_14253,N_15442);
and U19118 (N_19118,N_18450,N_15899);
nor U19119 (N_19119,N_12739,N_12967);
or U19120 (N_19120,N_13207,N_17855);
nor U19121 (N_19121,N_14846,N_16364);
and U19122 (N_19122,N_17889,N_15906);
nand U19123 (N_19123,N_15113,N_16881);
nor U19124 (N_19124,N_15443,N_18721);
and U19125 (N_19125,N_16411,N_12512);
and U19126 (N_19126,N_14254,N_18682);
and U19127 (N_19127,N_14882,N_13618);
xnor U19128 (N_19128,N_16193,N_13729);
nor U19129 (N_19129,N_15612,N_15904);
xnor U19130 (N_19130,N_17143,N_14120);
nor U19131 (N_19131,N_18652,N_16033);
or U19132 (N_19132,N_15868,N_14299);
or U19133 (N_19133,N_15059,N_16430);
nor U19134 (N_19134,N_18022,N_13965);
nor U19135 (N_19135,N_14441,N_14058);
or U19136 (N_19136,N_15679,N_15559);
nand U19137 (N_19137,N_18088,N_12778);
or U19138 (N_19138,N_17870,N_14333);
and U19139 (N_19139,N_15274,N_12965);
or U19140 (N_19140,N_15385,N_16841);
nor U19141 (N_19141,N_13727,N_12527);
or U19142 (N_19142,N_18728,N_17087);
xnor U19143 (N_19143,N_15599,N_15252);
or U19144 (N_19144,N_16000,N_15511);
nand U19145 (N_19145,N_17125,N_13049);
nand U19146 (N_19146,N_14817,N_15898);
nor U19147 (N_19147,N_13692,N_14929);
and U19148 (N_19148,N_18066,N_13568);
nand U19149 (N_19149,N_14743,N_16168);
nor U19150 (N_19150,N_13222,N_16165);
and U19151 (N_19151,N_15743,N_17248);
xnor U19152 (N_19152,N_15139,N_13298);
and U19153 (N_19153,N_16914,N_14771);
and U19154 (N_19154,N_14684,N_16273);
nor U19155 (N_19155,N_17256,N_18050);
nor U19156 (N_19156,N_16297,N_15566);
nor U19157 (N_19157,N_13360,N_14774);
nand U19158 (N_19158,N_15190,N_15448);
nand U19159 (N_19159,N_16762,N_12556);
nor U19160 (N_19160,N_15620,N_14936);
nand U19161 (N_19161,N_14543,N_15724);
or U19162 (N_19162,N_16813,N_15859);
nor U19163 (N_19163,N_14832,N_14944);
nor U19164 (N_19164,N_14401,N_17931);
or U19165 (N_19165,N_17896,N_16766);
and U19166 (N_19166,N_14652,N_12793);
and U19167 (N_19167,N_17465,N_14550);
nand U19168 (N_19168,N_16316,N_17848);
nor U19169 (N_19169,N_17049,N_17499);
nor U19170 (N_19170,N_16751,N_15974);
and U19171 (N_19171,N_16655,N_18094);
and U19172 (N_19172,N_13264,N_14608);
nand U19173 (N_19173,N_14079,N_13685);
nor U19174 (N_19174,N_13110,N_18461);
and U19175 (N_19175,N_14623,N_14140);
nor U19176 (N_19176,N_17162,N_16475);
xnor U19177 (N_19177,N_16639,N_16810);
xnor U19178 (N_19178,N_16678,N_16310);
and U19179 (N_19179,N_13290,N_14995);
and U19180 (N_19180,N_18518,N_18075);
and U19181 (N_19181,N_17287,N_18392);
xor U19182 (N_19182,N_14278,N_15381);
nand U19183 (N_19183,N_13484,N_14465);
or U19184 (N_19184,N_13143,N_12593);
or U19185 (N_19185,N_15186,N_14679);
and U19186 (N_19186,N_18367,N_17222);
nand U19187 (N_19187,N_13414,N_14113);
and U19188 (N_19188,N_13540,N_18396);
nor U19189 (N_19189,N_17808,N_12896);
xnor U19190 (N_19190,N_17634,N_18521);
or U19191 (N_19191,N_17082,N_17775);
and U19192 (N_19192,N_13413,N_16199);
nor U19193 (N_19193,N_16467,N_18562);
or U19194 (N_19194,N_17910,N_16377);
nand U19195 (N_19195,N_15098,N_13724);
and U19196 (N_19196,N_16556,N_15382);
and U19197 (N_19197,N_17849,N_13500);
and U19198 (N_19198,N_17188,N_17098);
xor U19199 (N_19199,N_15307,N_15569);
or U19200 (N_19200,N_17026,N_14805);
nand U19201 (N_19201,N_13794,N_17877);
nor U19202 (N_19202,N_12920,N_13838);
and U19203 (N_19203,N_13905,N_12827);
nor U19204 (N_19204,N_15121,N_15441);
nand U19205 (N_19205,N_14285,N_13726);
or U19206 (N_19206,N_12822,N_17257);
and U19207 (N_19207,N_13886,N_17258);
nor U19208 (N_19208,N_15771,N_14107);
nor U19209 (N_19209,N_14246,N_13677);
nor U19210 (N_19210,N_13659,N_18379);
nand U19211 (N_19211,N_17776,N_18298);
or U19212 (N_19212,N_13419,N_13890);
and U19213 (N_19213,N_12924,N_15099);
nor U19214 (N_19214,N_14719,N_13176);
nor U19215 (N_19215,N_16569,N_13703);
nand U19216 (N_19216,N_18655,N_13092);
or U19217 (N_19217,N_15878,N_16460);
nor U19218 (N_19218,N_14522,N_14157);
nor U19219 (N_19219,N_17698,N_12768);
and U19220 (N_19220,N_17869,N_15809);
nand U19221 (N_19221,N_15808,N_13514);
and U19222 (N_19222,N_17681,N_14516);
and U19223 (N_19223,N_12651,N_16024);
nor U19224 (N_19224,N_12854,N_13900);
nor U19225 (N_19225,N_16651,N_14619);
nor U19226 (N_19226,N_17807,N_16519);
or U19227 (N_19227,N_17661,N_12627);
nor U19228 (N_19228,N_13761,N_17380);
nor U19229 (N_19229,N_13234,N_18656);
nand U19230 (N_19230,N_17516,N_16476);
and U19231 (N_19231,N_15339,N_15081);
nand U19232 (N_19232,N_18217,N_16283);
xor U19233 (N_19233,N_18186,N_15894);
and U19234 (N_19234,N_13702,N_18554);
or U19235 (N_19235,N_14583,N_13725);
or U19236 (N_19236,N_13245,N_14338);
nand U19237 (N_19237,N_15198,N_14812);
nor U19238 (N_19238,N_17114,N_15895);
and U19239 (N_19239,N_18030,N_17803);
nand U19240 (N_19240,N_17442,N_17161);
nor U19241 (N_19241,N_18697,N_17408);
and U19242 (N_19242,N_15491,N_17029);
xor U19243 (N_19243,N_17168,N_12771);
nand U19244 (N_19244,N_17350,N_15215);
and U19245 (N_19245,N_15311,N_15760);
or U19246 (N_19246,N_13015,N_13983);
xor U19247 (N_19247,N_18669,N_15840);
or U19248 (N_19248,N_17385,N_16054);
or U19249 (N_19249,N_12575,N_16604);
or U19250 (N_19250,N_17868,N_15541);
xnor U19251 (N_19251,N_18414,N_15285);
and U19252 (N_19252,N_18372,N_13135);
xnor U19253 (N_19253,N_16528,N_12576);
or U19254 (N_19254,N_16048,N_16796);
and U19255 (N_19255,N_12814,N_12842);
nor U19256 (N_19256,N_13757,N_15393);
xnor U19257 (N_19257,N_18272,N_18128);
and U19258 (N_19258,N_18143,N_17043);
nor U19259 (N_19259,N_16269,N_13169);
or U19260 (N_19260,N_18606,N_16573);
nor U19261 (N_19261,N_14311,N_13064);
or U19262 (N_19262,N_16750,N_16913);
and U19263 (N_19263,N_15723,N_16945);
nand U19264 (N_19264,N_13178,N_14494);
xor U19265 (N_19265,N_18340,N_13425);
and U19266 (N_19266,N_15189,N_15320);
nand U19267 (N_19267,N_15440,N_12907);
or U19268 (N_19268,N_15013,N_15688);
nand U19269 (N_19269,N_17482,N_14523);
and U19270 (N_19270,N_17755,N_14450);
or U19271 (N_19271,N_17779,N_17128);
and U19272 (N_19272,N_12962,N_16031);
nand U19273 (N_19273,N_15828,N_13711);
nand U19274 (N_19274,N_16360,N_16361);
nor U19275 (N_19275,N_16118,N_18457);
nor U19276 (N_19276,N_14039,N_15889);
or U19277 (N_19277,N_16438,N_13270);
or U19278 (N_19278,N_12742,N_15232);
xor U19279 (N_19279,N_17790,N_14965);
nand U19280 (N_19280,N_15562,N_12680);
and U19281 (N_19281,N_18193,N_17736);
or U19282 (N_19282,N_14791,N_12937);
nor U19283 (N_19283,N_13436,N_16330);
or U19284 (N_19284,N_12951,N_12623);
or U19285 (N_19285,N_17403,N_16092);
and U19286 (N_19286,N_13931,N_13066);
or U19287 (N_19287,N_12574,N_18107);
or U19288 (N_19288,N_13097,N_13635);
nand U19289 (N_19289,N_13385,N_17336);
and U19290 (N_19290,N_12783,N_13192);
nand U19291 (N_19291,N_13912,N_16173);
nor U19292 (N_19292,N_14656,N_13941);
or U19293 (N_19293,N_16675,N_18139);
nor U19294 (N_19294,N_13809,N_15838);
and U19295 (N_19295,N_18342,N_15574);
or U19296 (N_19296,N_12523,N_16708);
nand U19297 (N_19297,N_13094,N_13841);
nor U19298 (N_19298,N_18454,N_17700);
or U19299 (N_19299,N_16266,N_15061);
or U19300 (N_19300,N_14471,N_15029);
or U19301 (N_19301,N_12604,N_13586);
nor U19302 (N_19302,N_15988,N_15365);
nor U19303 (N_19303,N_14620,N_15719);
or U19304 (N_19304,N_15045,N_17372);
nor U19305 (N_19305,N_14966,N_14725);
and U19306 (N_19306,N_18393,N_18497);
nor U19307 (N_19307,N_15212,N_13048);
nor U19308 (N_19308,N_13172,N_18261);
or U19309 (N_19309,N_18164,N_17605);
nand U19310 (N_19310,N_13106,N_14491);
nor U19311 (N_19311,N_13852,N_14224);
xnor U19312 (N_19312,N_17524,N_17937);
or U19313 (N_19313,N_17093,N_18082);
or U19314 (N_19314,N_13208,N_12583);
and U19315 (N_19315,N_17271,N_14421);
nor U19316 (N_19316,N_17641,N_14796);
and U19317 (N_19317,N_13167,N_16710);
and U19318 (N_19318,N_16507,N_15053);
xor U19319 (N_19319,N_18593,N_17410);
xor U19320 (N_19320,N_17614,N_17426);
or U19321 (N_19321,N_17969,N_14066);
or U19322 (N_19322,N_15194,N_18038);
and U19323 (N_19323,N_16246,N_17249);
nand U19324 (N_19324,N_16029,N_15125);
nor U19325 (N_19325,N_16223,N_16085);
and U19326 (N_19326,N_14473,N_16874);
nand U19327 (N_19327,N_16271,N_14277);
or U19328 (N_19328,N_16309,N_13539);
and U19329 (N_19329,N_18527,N_15286);
nand U19330 (N_19330,N_18418,N_14469);
nand U19331 (N_19331,N_15222,N_15362);
nor U19332 (N_19332,N_14903,N_14347);
or U19333 (N_19333,N_16821,N_18136);
xnor U19334 (N_19334,N_12994,N_17486);
or U19335 (N_19335,N_15702,N_16663);
and U19336 (N_19336,N_13068,N_12879);
nand U19337 (N_19337,N_16485,N_17512);
nand U19338 (N_19338,N_15003,N_18599);
and U19339 (N_19339,N_18114,N_17819);
nand U19340 (N_19340,N_15909,N_17763);
nand U19341 (N_19341,N_12910,N_18486);
nand U19342 (N_19342,N_14308,N_14024);
and U19343 (N_19343,N_12577,N_14009);
xnor U19344 (N_19344,N_13828,N_15466);
nand U19345 (N_19345,N_16561,N_14546);
nor U19346 (N_19346,N_13278,N_12502);
or U19347 (N_19347,N_14564,N_15499);
nor U19348 (N_19348,N_17631,N_14043);
and U19349 (N_19349,N_12804,N_14874);
or U19350 (N_19350,N_17356,N_17818);
nor U19351 (N_19351,N_15678,N_15046);
nand U19352 (N_19352,N_15105,N_12688);
or U19353 (N_19353,N_13212,N_13376);
xnor U19354 (N_19354,N_14563,N_13099);
nor U19355 (N_19355,N_14023,N_12586);
nor U19356 (N_19356,N_14754,N_14891);
and U19357 (N_19357,N_14849,N_18112);
or U19358 (N_19358,N_12505,N_15544);
or U19359 (N_19359,N_17412,N_18292);
nand U19360 (N_19360,N_16167,N_15298);
or U19361 (N_19361,N_18321,N_13543);
and U19362 (N_19362,N_12585,N_13595);
nand U19363 (N_19363,N_13499,N_14806);
nand U19364 (N_19364,N_18572,N_16095);
nand U19365 (N_19365,N_17595,N_12689);
xnor U19366 (N_19366,N_13782,N_15279);
nor U19367 (N_19367,N_13404,N_17772);
or U19368 (N_19368,N_13050,N_12743);
or U19369 (N_19369,N_17002,N_18584);
and U19370 (N_19370,N_14219,N_17938);
nor U19371 (N_19371,N_14987,N_16711);
nand U19372 (N_19372,N_16933,N_13363);
and U19373 (N_19373,N_18462,N_16036);
nor U19374 (N_19374,N_16335,N_13215);
xor U19375 (N_19375,N_13074,N_17993);
or U19376 (N_19376,N_15112,N_17184);
xnor U19377 (N_19377,N_14955,N_13787);
xor U19378 (N_19378,N_15251,N_17051);
nor U19379 (N_19379,N_14069,N_18701);
or U19380 (N_19380,N_15647,N_17553);
nor U19381 (N_19381,N_18650,N_15280);
nand U19382 (N_19382,N_12548,N_16061);
and U19383 (N_19383,N_14189,N_15604);
and U19384 (N_19384,N_16825,N_15801);
nand U19385 (N_19385,N_15221,N_14763);
or U19386 (N_19386,N_13394,N_15581);
nor U19387 (N_19387,N_13028,N_14979);
or U19388 (N_19388,N_14423,N_16347);
nand U19389 (N_19389,N_15407,N_16832);
and U19390 (N_19390,N_13490,N_12719);
or U19391 (N_19391,N_15908,N_17362);
or U19392 (N_19392,N_13498,N_16068);
nand U19393 (N_19393,N_12976,N_12732);
xor U19394 (N_19394,N_15312,N_13183);
or U19395 (N_19395,N_14235,N_15785);
nand U19396 (N_19396,N_18306,N_16028);
and U19397 (N_19397,N_12766,N_13406);
and U19398 (N_19398,N_15355,N_15711);
and U19399 (N_19399,N_13117,N_17793);
nand U19400 (N_19400,N_16397,N_17521);
nor U19401 (N_19401,N_17941,N_18023);
nand U19402 (N_19402,N_16190,N_17558);
nor U19403 (N_19403,N_13459,N_17828);
and U19404 (N_19404,N_18476,N_15954);
or U19405 (N_19405,N_17133,N_14328);
nor U19406 (N_19406,N_18708,N_13554);
or U19407 (N_19407,N_15825,N_16860);
or U19408 (N_19408,N_13246,N_16256);
nor U19409 (N_19409,N_14186,N_15796);
xnor U19410 (N_19410,N_18350,N_18464);
nand U19411 (N_19411,N_17582,N_17069);
or U19412 (N_19412,N_16902,N_18534);
nor U19413 (N_19413,N_15932,N_17887);
and U19414 (N_19414,N_16253,N_16337);
nor U19415 (N_19415,N_12539,N_13061);
nand U19416 (N_19416,N_15492,N_16073);
and U19417 (N_19417,N_18332,N_17227);
and U19418 (N_19418,N_16080,N_13259);
xor U19419 (N_19419,N_18070,N_16578);
or U19420 (N_19420,N_12913,N_16171);
nor U19421 (N_19421,N_17963,N_14130);
nor U19422 (N_19422,N_15143,N_13004);
and U19423 (N_19423,N_14864,N_12660);
nor U19424 (N_19424,N_12996,N_15248);
xor U19425 (N_19425,N_17965,N_17809);
nor U19426 (N_19426,N_18257,N_13331);
nand U19427 (N_19427,N_14268,N_17908);
and U19428 (N_19428,N_18110,N_14054);
and U19429 (N_19429,N_18666,N_16732);
xnor U19430 (N_19430,N_13656,N_18552);
xnor U19431 (N_19431,N_16306,N_14638);
nor U19432 (N_19432,N_18702,N_18443);
nor U19433 (N_19433,N_14688,N_14984);
or U19434 (N_19434,N_12533,N_17827);
and U19435 (N_19435,N_12880,N_12745);
xnor U19436 (N_19436,N_14907,N_14881);
nor U19437 (N_19437,N_16941,N_17209);
and U19438 (N_19438,N_15607,N_15618);
nor U19439 (N_19439,N_17765,N_12618);
or U19440 (N_19440,N_13070,N_17714);
and U19441 (N_19441,N_14597,N_14605);
or U19442 (N_19442,N_16357,N_14259);
and U19443 (N_19443,N_17643,N_13471);
and U19444 (N_19444,N_13883,N_13211);
xor U19445 (N_19445,N_12645,N_14415);
and U19446 (N_19446,N_13198,N_16694);
and U19447 (N_19447,N_14109,N_18644);
or U19448 (N_19448,N_15486,N_18688);
xor U19449 (N_19449,N_16027,N_16144);
or U19450 (N_19450,N_14241,N_13981);
nand U19451 (N_19451,N_14209,N_14670);
xor U19452 (N_19452,N_14693,N_14094);
and U19453 (N_19453,N_13434,N_14068);
and U19454 (N_19454,N_12947,N_13680);
nand U19455 (N_19455,N_14721,N_13752);
and U19456 (N_19456,N_17729,N_17067);
or U19457 (N_19457,N_16229,N_16106);
xnor U19458 (N_19458,N_12953,N_17858);
nand U19459 (N_19459,N_18600,N_18505);
xor U19460 (N_19460,N_18191,N_14065);
and U19461 (N_19461,N_15671,N_15734);
xnor U19462 (N_19462,N_14780,N_16544);
nor U19463 (N_19463,N_12931,N_15687);
nand U19464 (N_19464,N_13239,N_15230);
nor U19465 (N_19465,N_16295,N_17526);
xor U19466 (N_19466,N_13087,N_13749);
or U19467 (N_19467,N_13840,N_13709);
nor U19468 (N_19468,N_15503,N_15162);
and U19469 (N_19469,N_14118,N_17346);
nand U19470 (N_19470,N_15211,N_15055);
nor U19471 (N_19471,N_16172,N_17979);
nand U19472 (N_19472,N_13380,N_15554);
nand U19473 (N_19473,N_15435,N_17094);
nor U19474 (N_19474,N_18513,N_18097);
nand U19475 (N_19475,N_12868,N_17284);
nand U19476 (N_19476,N_17906,N_16697);
and U19477 (N_19477,N_13478,N_14313);
and U19478 (N_19478,N_18533,N_18675);
nor U19479 (N_19479,N_15869,N_17376);
or U19480 (N_19480,N_13564,N_17633);
or U19481 (N_19481,N_13548,N_13791);
nand U19482 (N_19482,N_18263,N_17243);
nand U19483 (N_19483,N_13492,N_18585);
or U19484 (N_19484,N_16491,N_14594);
nor U19485 (N_19485,N_14666,N_13445);
xor U19486 (N_19486,N_15369,N_15449);
nor U19487 (N_19487,N_16904,N_15865);
nor U19488 (N_19488,N_15964,N_17915);
nand U19489 (N_19489,N_15730,N_13274);
or U19490 (N_19490,N_17800,N_15022);
and U19491 (N_19491,N_18081,N_15424);
nor U19492 (N_19492,N_18098,N_13877);
nor U19493 (N_19493,N_14590,N_16548);
or U19494 (N_19494,N_16204,N_16208);
and U19495 (N_19495,N_16580,N_16378);
nand U19496 (N_19496,N_12615,N_12638);
xnor U19497 (N_19497,N_13903,N_15955);
nor U19498 (N_19498,N_12513,N_14265);
nand U19499 (N_19499,N_17283,N_18575);
or U19500 (N_19500,N_17304,N_12869);
nor U19501 (N_19501,N_13926,N_15646);
nor U19502 (N_19502,N_13221,N_13773);
nand U19503 (N_19503,N_13580,N_13876);
and U19504 (N_19504,N_18297,N_15106);
nor U19505 (N_19505,N_13678,N_17612);
or U19506 (N_19506,N_13666,N_15858);
nor U19507 (N_19507,N_15950,N_15476);
nand U19508 (N_19508,N_15578,N_12812);
nand U19509 (N_19509,N_18729,N_13646);
nor U19510 (N_19510,N_18313,N_13114);
nand U19511 (N_19511,N_15933,N_13513);
nand U19512 (N_19512,N_15804,N_15587);
nand U19513 (N_19513,N_17991,N_17207);
nor U19514 (N_19514,N_13269,N_13353);
nor U19515 (N_19515,N_18528,N_16016);
nor U19516 (N_19516,N_17054,N_12993);
or U19517 (N_19517,N_16992,N_16124);
xnor U19518 (N_19518,N_15118,N_17371);
and U19519 (N_19519,N_17767,N_14675);
nand U19520 (N_19520,N_16918,N_13166);
and U19521 (N_19521,N_16927,N_17017);
and U19522 (N_19522,N_17216,N_16060);
nor U19523 (N_19523,N_17315,N_13639);
and U19524 (N_19524,N_15042,N_18251);
nor U19525 (N_19525,N_15358,N_18431);
and U19526 (N_19526,N_17543,N_16392);
nand U19527 (N_19527,N_14394,N_15631);
nor U19528 (N_19528,N_12853,N_18588);
or U19529 (N_19529,N_13249,N_14003);
nor U19530 (N_19530,N_18570,N_18236);
or U19531 (N_19531,N_13916,N_18033);
or U19532 (N_19532,N_12547,N_14909);
nand U19533 (N_19533,N_17703,N_18155);
and U19534 (N_19534,N_12567,N_14216);
nand U19535 (N_19535,N_16355,N_15085);
nand U19536 (N_19536,N_14601,N_15436);
nor U19537 (N_19537,N_13963,N_18536);
nor U19538 (N_19538,N_18072,N_14613);
nor U19539 (N_19539,N_14099,N_16975);
nor U19540 (N_19540,N_14432,N_12560);
nand U19541 (N_19541,N_16838,N_16139);
nor U19542 (N_19542,N_14442,N_15034);
nand U19543 (N_19543,N_18658,N_15203);
and U19544 (N_19544,N_17618,N_17757);
and U19545 (N_19545,N_18714,N_18004);
or U19546 (N_19546,N_12652,N_17654);
nand U19547 (N_19547,N_16277,N_18694);
nand U19548 (N_19548,N_12762,N_17441);
and U19549 (N_19549,N_15842,N_15147);
or U19550 (N_19550,N_15071,N_13021);
nand U19551 (N_19551,N_17191,N_13164);
or U19552 (N_19552,N_13179,N_16242);
or U19553 (N_19553,N_13383,N_18547);
nor U19554 (N_19554,N_16720,N_15376);
or U19555 (N_19555,N_18021,N_14449);
nand U19556 (N_19556,N_12622,N_16540);
nor U19557 (N_19557,N_18137,N_15091);
nor U19558 (N_19558,N_17144,N_16126);
or U19559 (N_19559,N_17606,N_15718);
nand U19560 (N_19560,N_17364,N_18720);
or U19561 (N_19561,N_17546,N_13163);
and U19562 (N_19562,N_17182,N_17873);
or U19563 (N_19563,N_12952,N_15656);
nand U19564 (N_19564,N_14243,N_18596);
nor U19565 (N_19565,N_18742,N_14366);
nor U19566 (N_19566,N_15543,N_14919);
nand U19567 (N_19567,N_14985,N_14403);
nand U19568 (N_19568,N_13267,N_13417);
or U19569 (N_19569,N_14373,N_14038);
nor U19570 (N_19570,N_15321,N_16722);
and U19571 (N_19571,N_17747,N_17171);
and U19572 (N_19572,N_14599,N_18522);
nand U19573 (N_19573,N_15291,N_15990);
nand U19574 (N_19574,N_15090,N_12946);
and U19575 (N_19575,N_18254,N_17468);
and U19576 (N_19576,N_18119,N_18180);
nand U19577 (N_19577,N_16875,N_15374);
or U19578 (N_19578,N_14201,N_15542);
and U19579 (N_19579,N_13260,N_17036);
nand U19580 (N_19580,N_12826,N_18395);
and U19581 (N_19581,N_15304,N_16436);
nor U19582 (N_19582,N_13411,N_14775);
nor U19583 (N_19583,N_15952,N_14859);
nor U19584 (N_19584,N_17530,N_18412);
nand U19585 (N_19585,N_15717,N_13832);
nor U19586 (N_19586,N_17289,N_14398);
and U19587 (N_19587,N_17484,N_13453);
and U19588 (N_19588,N_18055,N_14357);
xor U19589 (N_19589,N_15721,N_14603);
nand U19590 (N_19590,N_16889,N_13043);
nor U19591 (N_19591,N_17871,N_13651);
nor U19592 (N_19592,N_13908,N_13693);
or U19593 (N_19593,N_17493,N_16787);
nor U19594 (N_19594,N_15073,N_16611);
nand U19595 (N_19595,N_13096,N_17627);
and U19596 (N_19596,N_15737,N_17323);
nand U19597 (N_19597,N_16206,N_15068);
nor U19598 (N_19598,N_18684,N_12926);
or U19599 (N_19599,N_12847,N_17913);
or U19600 (N_19600,N_14512,N_12985);
or U19601 (N_19601,N_16944,N_17141);
or U19602 (N_19602,N_15794,N_14758);
or U19603 (N_19603,N_15333,N_13768);
or U19604 (N_19604,N_17821,N_12754);
nand U19605 (N_19605,N_13875,N_13872);
and U19606 (N_19606,N_16406,N_15799);
and U19607 (N_19607,N_16299,N_15969);
or U19608 (N_19608,N_16169,N_17157);
and U19609 (N_19609,N_14747,N_15439);
nand U19610 (N_19610,N_14949,N_13679);
nor U19611 (N_19611,N_16496,N_16338);
or U19612 (N_19612,N_18300,N_15131);
and U19613 (N_19613,N_16072,N_17317);
or U19614 (N_19614,N_17693,N_16920);
and U19615 (N_19615,N_16940,N_12669);
or U19616 (N_19616,N_16816,N_14343);
and U19617 (N_19617,N_14749,N_17690);
nand U19618 (N_19618,N_18317,N_14049);
or U19619 (N_19619,N_14757,N_12640);
nor U19620 (N_19620,N_17298,N_13171);
or U19621 (N_19621,N_15394,N_16414);
and U19622 (N_19622,N_12702,N_16429);
nor U19623 (N_19623,N_15610,N_13974);
xor U19624 (N_19624,N_15664,N_18449);
nand U19625 (N_19625,N_17617,N_15596);
or U19626 (N_19626,N_15770,N_18111);
and U19627 (N_19627,N_18741,N_17127);
or U19628 (N_19628,N_14628,N_13525);
or U19629 (N_19629,N_18210,N_18619);
nand U19630 (N_19630,N_15141,N_14020);
nor U19631 (N_19631,N_15278,N_17540);
xor U19632 (N_19632,N_13161,N_16145);
and U19633 (N_19633,N_16854,N_16178);
nand U19634 (N_19634,N_16101,N_17373);
or U19635 (N_19635,N_17596,N_14141);
and U19636 (N_19636,N_14927,N_14044);
nand U19637 (N_19637,N_18006,N_18202);
or U19638 (N_19638,N_17205,N_15271);
and U19639 (N_19639,N_17085,N_14283);
nor U19640 (N_19640,N_14706,N_14941);
xor U19641 (N_19641,N_17875,N_15380);
nor U19642 (N_19642,N_14819,N_13818);
or U19643 (N_19643,N_15890,N_14380);
nand U19644 (N_19644,N_13885,N_18012);
xor U19645 (N_19645,N_17725,N_17623);
and U19646 (N_19646,N_16001,N_17679);
and U19647 (N_19647,N_15408,N_17705);
nor U19648 (N_19648,N_12666,N_18475);
nor U19649 (N_19649,N_17213,N_13869);
nor U19650 (N_19650,N_17886,N_13857);
or U19651 (N_19651,N_17366,N_12991);
or U19652 (N_19652,N_18303,N_15316);
nand U19653 (N_19653,N_13755,N_14359);
or U19654 (N_19654,N_17367,N_15021);
and U19655 (N_19655,N_17786,N_16553);
nor U19656 (N_19656,N_14208,N_18685);
or U19657 (N_19657,N_12908,N_16109);
nor U19658 (N_19658,N_15611,N_18031);
or U19659 (N_19659,N_15866,N_17577);
nor U19660 (N_19660,N_17028,N_13642);
or U19661 (N_19661,N_16107,N_15882);
nand U19662 (N_19662,N_14994,N_13468);
or U19663 (N_19663,N_18252,N_13764);
nor U19664 (N_19664,N_13937,N_14410);
or U19665 (N_19665,N_15184,N_15253);
nand U19666 (N_19666,N_17390,N_13552);
nor U19667 (N_19667,N_14239,N_16764);
and U19668 (N_19668,N_13272,N_14511);
or U19669 (N_19669,N_13149,N_17628);
nor U19670 (N_19670,N_15461,N_13457);
xnor U19671 (N_19671,N_13343,N_17444);
nor U19672 (N_19672,N_18571,N_14504);
nor U19673 (N_19673,N_12606,N_15371);
nor U19674 (N_19674,N_13115,N_12597);
nand U19675 (N_19675,N_14298,N_14087);
or U19676 (N_19676,N_16500,N_16780);
nor U19677 (N_19677,N_13475,N_14575);
nand U19678 (N_19678,N_14876,N_18388);
or U19679 (N_19679,N_17437,N_18341);
or U19680 (N_19680,N_13546,N_16589);
and U19681 (N_19681,N_17180,N_17303);
nand U19682 (N_19682,N_17311,N_16372);
and U19683 (N_19683,N_17397,N_17095);
and U19684 (N_19684,N_17758,N_15841);
or U19685 (N_19685,N_13550,N_12721);
or U19686 (N_19686,N_13884,N_15698);
nand U19687 (N_19687,N_16325,N_12653);
nand U19688 (N_19688,N_18355,N_12981);
xor U19689 (N_19689,N_13124,N_14183);
or U19690 (N_19690,N_17476,N_16617);
nor U19691 (N_19691,N_17571,N_15976);
nand U19692 (N_19692,N_15914,N_14717);
and U19693 (N_19693,N_17264,N_15403);
or U19694 (N_19694,N_13196,N_13722);
nor U19695 (N_19695,N_13951,N_14710);
nand U19696 (N_19696,N_17003,N_12982);
nand U19697 (N_19697,N_18123,N_14445);
or U19698 (N_19698,N_15269,N_18491);
and U19699 (N_19699,N_13451,N_17134);
and U19700 (N_19700,N_16440,N_17387);
nand U19701 (N_19701,N_16350,N_14712);
nor U19702 (N_19702,N_16674,N_12509);
nor U19703 (N_19703,N_16181,N_16778);
nand U19704 (N_19704,N_15445,N_17192);
or U19705 (N_19705,N_13915,N_16554);
and U19706 (N_19706,N_14281,N_13495);
and U19707 (N_19707,N_14019,N_14915);
or U19708 (N_19708,N_16570,N_12884);
or U19709 (N_19709,N_13355,N_15002);
or U19710 (N_19710,N_17568,N_18002);
nand U19711 (N_19711,N_13921,N_16683);
or U19712 (N_19712,N_15639,N_16822);
and U19713 (N_19713,N_15772,N_17917);
or U19714 (N_19714,N_15173,N_17384);
nand U19715 (N_19715,N_13302,N_18506);
and U19716 (N_19716,N_15206,N_13922);
and U19717 (N_19717,N_16799,N_12571);
nand U19718 (N_19718,N_12797,N_17354);
nand U19719 (N_19719,N_18683,N_14695);
nand U19720 (N_19720,N_18580,N_14506);
nor U19721 (N_19721,N_13825,N_16484);
or U19722 (N_19722,N_15767,N_13080);
and U19723 (N_19723,N_13942,N_18433);
and U19724 (N_19724,N_13047,N_12635);
or U19725 (N_19725,N_17473,N_13300);
xnor U19726 (N_19726,N_17680,N_14606);
nor U19727 (N_19727,N_18727,N_15467);
nor U19728 (N_19728,N_13789,N_13151);
nor U19729 (N_19729,N_13662,N_18008);
and U19730 (N_19730,N_15301,N_12705);
nor U19731 (N_19731,N_16575,N_14000);
or U19732 (N_19732,N_17232,N_17459);
nor U19733 (N_19733,N_18102,N_16585);
and U19734 (N_19734,N_18178,N_14156);
nor U19735 (N_19735,N_18290,N_16417);
nand U19736 (N_19736,N_17428,N_15892);
nor U19737 (N_19737,N_12554,N_15512);
nor U19738 (N_19738,N_13734,N_14290);
nand U19739 (N_19739,N_18598,N_17724);
xor U19740 (N_19740,N_17101,N_12603);
xnor U19741 (N_19741,N_14922,N_17064);
and U19742 (N_19742,N_16135,N_16624);
nor U19743 (N_19743,N_15773,N_13913);
nor U19744 (N_19744,N_17662,N_16343);
nand U19745 (N_19745,N_15746,N_13311);
nand U19746 (N_19746,N_16747,N_16482);
and U19747 (N_19747,N_12781,N_15329);
or U19748 (N_19748,N_17542,N_15343);
and U19749 (N_19749,N_18538,N_13241);
and U19750 (N_19750,N_14982,N_16631);
or U19751 (N_19751,N_18725,N_18744);
nor U19752 (N_19752,N_16677,N_18249);
or U19753 (N_19753,N_12939,N_13814);
or U19754 (N_19754,N_13285,N_15823);
or U19755 (N_19755,N_16098,N_14974);
or U19756 (N_19756,N_17742,N_15142);
nor U19757 (N_19757,N_13788,N_15910);
nor U19758 (N_19758,N_13133,N_17925);
xor U19759 (N_19759,N_15877,N_17592);
nand U19760 (N_19760,N_14399,N_12584);
and U19761 (N_19761,N_15856,N_18322);
nor U19762 (N_19762,N_17183,N_16924);
nand U19763 (N_19763,N_14755,N_18634);
and U19764 (N_19764,N_18026,N_13704);
nor U19765 (N_19765,N_14701,N_16510);
nand U19766 (N_19766,N_17121,N_13948);
or U19767 (N_19767,N_18301,N_17024);
or U19768 (N_19768,N_17519,N_18482);
nand U19769 (N_19769,N_15086,N_12708);
nand U19770 (N_19770,N_12625,N_14646);
nor U19771 (N_19771,N_16055,N_17394);
nand U19772 (N_19772,N_17102,N_15255);
or U19773 (N_19773,N_15336,N_13410);
nand U19774 (N_19774,N_14084,N_14568);
or U19775 (N_19775,N_15916,N_17752);
xnor U19776 (N_19776,N_17660,N_18077);
nor U19777 (N_19777,N_16287,N_13968);
xor U19778 (N_19778,N_18344,N_12819);
and U19779 (N_19779,N_17859,N_18287);
nand U19780 (N_19780,N_16673,N_18560);
or U19781 (N_19781,N_17522,N_15634);
xnor U19782 (N_19782,N_18320,N_13339);
and U19783 (N_19783,N_17632,N_17443);
and U19784 (N_19784,N_13661,N_17563);
nor U19785 (N_19785,N_12643,N_16644);
xnor U19786 (N_19786,N_12711,N_13705);
and U19787 (N_19787,N_18735,N_16969);
and U19788 (N_19788,N_13524,N_13573);
nand U19789 (N_19789,N_14014,N_13938);
or U19790 (N_19790,N_15762,N_18040);
nand U19791 (N_19791,N_14558,N_15547);
nand U19792 (N_19792,N_16730,N_17088);
and U19793 (N_19793,N_17130,N_13802);
and U19794 (N_19794,N_16513,N_12882);
or U19795 (N_19795,N_15084,N_14997);
nor U19796 (N_19796,N_17560,N_17237);
or U19797 (N_19797,N_13868,N_17960);
and U19798 (N_19798,N_12563,N_16892);
or U19799 (N_19799,N_17063,N_17335);
nand U19800 (N_19800,N_14591,N_14865);
or U19801 (N_19801,N_18576,N_17597);
nand U19802 (N_19802,N_17139,N_15887);
nor U19803 (N_19803,N_13480,N_17649);
or U19804 (N_19804,N_13076,N_16610);
and U19805 (N_19805,N_16973,N_16291);
xor U19806 (N_19806,N_14207,N_18277);
nand U19807 (N_19807,N_14643,N_14830);
and U19808 (N_19808,N_17047,N_17942);
and U19809 (N_19809,N_18289,N_17865);
and U19810 (N_19810,N_14514,N_13377);
and U19811 (N_19811,N_15778,N_16856);
or U19812 (N_19812,N_18167,N_13634);
nand U19813 (N_19813,N_14937,N_17923);
and U19814 (N_19814,N_14735,N_12696);
or U19815 (N_19815,N_15233,N_17065);
and U19816 (N_19816,N_14053,N_16846);
nand U19817 (N_19817,N_17072,N_14419);
nand U19818 (N_19818,N_15295,N_16616);
or U19819 (N_19819,N_16725,N_12521);
nor U19820 (N_19820,N_13091,N_16943);
or U19821 (N_19821,N_17997,N_15530);
nor U19822 (N_19822,N_15420,N_13136);
nand U19823 (N_19823,N_18692,N_16094);
nor U19824 (N_19824,N_18268,N_13616);
nor U19825 (N_19825,N_17355,N_13082);
or U19826 (N_19826,N_17020,N_17850);
nor U19827 (N_19827,N_14878,N_15060);
nand U19828 (N_19828,N_18722,N_17214);
xnor U19829 (N_19829,N_15149,N_12849);
nor U19830 (N_19830,N_13102,N_16367);
and U19831 (N_19831,N_13930,N_13617);
and U19832 (N_19832,N_18463,N_17578);
nand U19833 (N_19833,N_13627,N_16505);
nand U19834 (N_19834,N_15666,N_13532);
and U19835 (N_19835,N_13681,N_15676);
and U19836 (N_19836,N_14400,N_13370);
and U19837 (N_19837,N_16481,N_17201);
and U19838 (N_19838,N_12964,N_14336);
and U19839 (N_19839,N_18368,N_12893);
and U19840 (N_19840,N_14916,N_18260);
or U19841 (N_19841,N_15318,N_16627);
and U19842 (N_19842,N_13031,N_14342);
nor U19843 (N_19843,N_13538,N_14155);
and U19844 (N_19844,N_16840,N_16198);
or U19845 (N_19845,N_18228,N_18238);
and U19846 (N_19846,N_15897,N_13042);
and U19847 (N_19847,N_16756,N_13710);
or U19848 (N_19848,N_17830,N_18624);
nand U19849 (N_19849,N_12629,N_18039);
nor U19850 (N_19850,N_18085,N_18623);
or U19851 (N_19851,N_14301,N_13217);
or U19852 (N_19852,N_14835,N_16739);
xor U19853 (N_19853,N_17456,N_13594);
nor U19854 (N_19854,N_14968,N_18273);
or U19855 (N_19855,N_13713,N_12559);
nor U19856 (N_19856,N_18222,N_14034);
or U19857 (N_19857,N_17536,N_14022);
nand U19858 (N_19858,N_16174,N_13182);
nand U19859 (N_19859,N_12930,N_17375);
xnor U19860 (N_19860,N_15277,N_14871);
and U19861 (N_19861,N_16989,N_16081);
or U19862 (N_19862,N_16777,N_16681);
and U19863 (N_19863,N_16314,N_14407);
and U19864 (N_19864,N_16153,N_18643);
or U19865 (N_19865,N_12534,N_17196);
and U19866 (N_19866,N_15425,N_16634);
nand U19867 (N_19867,N_18219,N_16962);
xor U19868 (N_19868,N_16082,N_12531);
or U19869 (N_19869,N_13736,N_15164);
and U19870 (N_19870,N_14577,N_18680);
nor U19871 (N_19871,N_16851,N_18541);
or U19872 (N_19872,N_16735,N_17591);
nor U19873 (N_19873,N_17559,N_13007);
nor U19874 (N_19874,N_13859,N_17025);
and U19875 (N_19875,N_15145,N_18557);
nor U19876 (N_19876,N_14724,N_15970);
nor U19877 (N_19877,N_18364,N_13523);
or U19878 (N_19878,N_14901,N_17699);
or U19879 (N_19879,N_14258,N_12698);
nand U19880 (N_19880,N_15341,N_13412);
and U19881 (N_19881,N_15774,N_18361);
or U19882 (N_19882,N_17172,N_13865);
or U19883 (N_19883,N_12510,N_15402);
and U19884 (N_19884,N_16078,N_15814);
or U19885 (N_19885,N_17135,N_15359);
nand U19886 (N_19886,N_12803,N_18618);
nor U19887 (N_19887,N_15845,N_15695);
and U19888 (N_19888,N_12565,N_13708);
nor U19889 (N_19889,N_13177,N_14355);
xor U19890 (N_19890,N_14958,N_17234);
or U19891 (N_19891,N_15120,N_13925);
and U19892 (N_19892,N_15356,N_18629);
and U19893 (N_19893,N_16645,N_15941);
xnor U19894 (N_19894,N_13849,N_12582);
xnor U19895 (N_19895,N_13851,N_14282);
nand U19896 (N_19896,N_17939,N_16520);
or U19897 (N_19897,N_13119,N_17861);
or U19898 (N_19898,N_15395,N_16968);
or U19899 (N_19899,N_13733,N_14760);
nor U19900 (N_19900,N_15815,N_15051);
nand U19901 (N_19901,N_16872,N_15683);
and U19902 (N_19902,N_12674,N_15372);
nand U19903 (N_19903,N_15303,N_18325);
or U19904 (N_19904,N_15925,N_18019);
and U19905 (N_19905,N_15110,N_14554);
nor U19906 (N_19906,N_14368,N_18504);
and U19907 (N_19907,N_13624,N_14654);
nor U19908 (N_19908,N_18558,N_15789);
and U19909 (N_19909,N_18127,N_13699);
nor U19910 (N_19910,N_13597,N_18062);
or U19911 (N_19911,N_18060,N_12809);
nor U19912 (N_19912,N_13767,N_17711);
and U19913 (N_19913,N_18530,N_13075);
nand U19914 (N_19914,N_16817,N_15833);
and U19915 (N_19915,N_17992,N_13431);
nor U19916 (N_19916,N_14479,N_17229);
nor U19917 (N_19917,N_17341,N_16809);
nand U19918 (N_19918,N_17140,N_13319);
or U19919 (N_19919,N_14683,N_16067);
and U19920 (N_19920,N_16026,N_16052);
and U19921 (N_19921,N_15739,N_16166);
nor U19922 (N_19922,N_13084,N_17041);
nor U19923 (N_19923,N_12722,N_18221);
xnor U19924 (N_19924,N_18665,N_18492);
and U19925 (N_19925,N_13316,N_12733);
xnor U19926 (N_19926,N_17566,N_17296);
nor U19927 (N_19927,N_15094,N_15783);
nand U19928 (N_19928,N_17446,N_17096);
nand U19929 (N_19929,N_18718,N_15982);
or U19930 (N_19930,N_13776,N_14808);
or U19931 (N_19931,N_18027,N_17739);
nand U19932 (N_19932,N_17653,N_16449);
or U19933 (N_19933,N_16282,N_16919);
nand U19934 (N_19934,N_14918,N_17586);
or U19935 (N_19935,N_12649,N_16836);
and U19936 (N_19936,N_15947,N_15244);
and U19937 (N_19937,N_16562,N_13461);
nand U19938 (N_19938,N_16463,N_13328);
and U19939 (N_19939,N_12867,N_14062);
or U19940 (N_19940,N_17111,N_15881);
nand U19941 (N_19941,N_15433,N_14586);
nand U19942 (N_19942,N_15290,N_14569);
nor U19943 (N_19943,N_14902,N_17198);
nor U19944 (N_19944,N_14602,N_15861);
xnor U19945 (N_19945,N_17494,N_15039);
nor U19946 (N_19946,N_16582,N_18076);
or U19947 (N_19947,N_14509,N_17805);
or U19948 (N_19948,N_14973,N_17475);
and U19949 (N_19949,N_14988,N_12975);
and U19950 (N_19950,N_14566,N_18671);
xnor U19951 (N_19951,N_14702,N_15709);
or U19952 (N_19952,N_15626,N_14225);
nor U19953 (N_19953,N_18365,N_16842);
nand U19954 (N_19954,N_17206,N_17891);
nor U19955 (N_19955,N_13591,N_17179);
or U19956 (N_19956,N_18271,N_14073);
and U19957 (N_19957,N_17383,N_16789);
and U19958 (N_19958,N_16421,N_12724);
or U19959 (N_19959,N_17706,N_17436);
nor U19960 (N_19960,N_15764,N_17874);
and U19961 (N_19961,N_18308,N_15837);
or U19962 (N_19962,N_17275,N_12617);
or U19963 (N_19963,N_13989,N_12641);
xor U19964 (N_19964,N_15662,N_13476);
nand U19965 (N_19965,N_14898,N_16953);
nand U19966 (N_19966,N_14637,N_18686);
and U19967 (N_19967,N_12670,N_15903);
nor U19968 (N_19968,N_18116,N_15048);
nand U19969 (N_19969,N_15600,N_12683);
and U19970 (N_19970,N_13566,N_13695);
and U19971 (N_19971,N_17255,N_13203);
nand U19972 (N_19972,N_12712,N_13188);
and U19973 (N_19973,N_14270,N_14928);
nor U19974 (N_19974,N_16131,N_14242);
nand U19975 (N_19975,N_17083,N_17109);
or U19976 (N_19976,N_12515,N_13655);
and U19977 (N_19977,N_13839,N_15790);
or U19978 (N_19978,N_15050,N_13407);
or U19979 (N_19979,N_12506,N_18421);
nand U19980 (N_19980,N_14332,N_15447);
nor U19981 (N_19981,N_16344,N_15167);
nor U19982 (N_19982,N_13988,N_14845);
nor U19983 (N_19983,N_15087,N_17491);
or U19984 (N_19984,N_15761,N_15337);
and U19985 (N_19985,N_14273,N_16758);
nor U19986 (N_19986,N_14692,N_14237);
xnor U19987 (N_19987,N_13723,N_14370);
or U19988 (N_19988,N_17048,N_16855);
nand U19989 (N_19989,N_17297,N_18602);
nand U19990 (N_19990,N_16895,N_17673);
and U19991 (N_19991,N_14840,N_18451);
and U19992 (N_19992,N_15658,N_14621);
xor U19993 (N_19993,N_17990,N_15097);
xnor U19994 (N_19994,N_17477,N_17590);
xor U19995 (N_19995,N_15249,N_13493);
nor U19996 (N_19996,N_15896,N_12546);
nor U19997 (N_19997,N_12813,N_13527);
or U19998 (N_19998,N_17392,N_13432);
nor U19999 (N_19999,N_14128,N_17956);
or U20000 (N_20000,N_13187,N_15668);
or U20001 (N_20001,N_14939,N_18270);
or U20002 (N_20002,N_14772,N_17034);
nand U20003 (N_20003,N_14625,N_13263);
nand U20004 (N_20004,N_15011,N_15082);
or U20005 (N_20005,N_13073,N_14287);
nor U20006 (N_20006,N_16857,N_17719);
and U20007 (N_20007,N_15254,N_17112);
nor U20008 (N_20008,N_16121,N_18197);
nand U20009 (N_20009,N_14674,N_14841);
or U20010 (N_20010,N_17381,N_16648);
or U20011 (N_20011,N_13779,N_18651);
nor U20012 (N_20012,N_13902,N_13760);
or U20013 (N_20013,N_18407,N_16408);
or U20014 (N_20014,N_16323,N_13976);
xor U20015 (N_20015,N_16819,N_13497);
or U20016 (N_20016,N_13334,N_17946);
or U20017 (N_20017,N_15388,N_12955);
nor U20018 (N_20018,N_14472,N_13235);
nand U20019 (N_20019,N_14350,N_15404);
xor U20020 (N_20020,N_13536,N_16761);
nor U20021 (N_20021,N_14658,N_14477);
nor U20022 (N_20022,N_12753,N_16608);
or U20023 (N_20023,N_12960,N_18543);
nor U20024 (N_20024,N_17534,N_18502);
and U20025 (N_20025,N_15625,N_15923);
nor U20026 (N_20026,N_16469,N_17716);
and U20027 (N_20027,N_13401,N_17610);
and U20028 (N_20028,N_14356,N_15017);
and U20029 (N_20029,N_15281,N_13397);
nand U20030 (N_20030,N_14948,N_16566);
or U20031 (N_20031,N_14418,N_16105);
xor U20032 (N_20032,N_13238,N_13199);
and U20033 (N_20033,N_16252,N_18467);
nand U20034 (N_20034,N_16459,N_16833);
nand U20035 (N_20035,N_17155,N_13250);
nor U20036 (N_20036,N_17841,N_17585);
nor U20037 (N_20037,N_12792,N_17966);
nand U20038 (N_20038,N_15603,N_18073);
xor U20039 (N_20039,N_17040,N_14080);
and U20040 (N_20040,N_17438,N_13730);
and U20041 (N_20041,N_14312,N_16622);
and U20042 (N_20042,N_15685,N_15766);
nor U20043 (N_20043,N_15803,N_15653);
and U20044 (N_20044,N_13018,N_13910);
nor U20045 (N_20045,N_15047,N_13650);
or U20046 (N_20046,N_12791,N_15065);
nor U20047 (N_20047,N_17005,N_14291);
and U20048 (N_20048,N_17795,N_13648);
and U20049 (N_20049,N_13085,N_16737);
nor U20050 (N_20050,N_14292,N_15712);
and U20051 (N_20051,N_18480,N_17211);
and U20052 (N_20052,N_16729,N_12681);
and U20053 (N_20053,N_15942,N_13392);
nand U20054 (N_20054,N_16490,N_15390);
nand U20055 (N_20055,N_16473,N_14376);
or U20056 (N_20056,N_12909,N_16431);
nand U20057 (N_20057,N_13489,N_14556);
nand U20058 (N_20058,N_16380,N_13786);
and U20059 (N_20059,N_15235,N_15294);
nand U20060 (N_20060,N_18140,N_15127);
or U20061 (N_20061,N_14393,N_17263);
and U20062 (N_20062,N_17015,N_18495);
or U20063 (N_20063,N_18531,N_14797);
nor U20064 (N_20064,N_15401,N_13095);
and U20065 (N_20065,N_16056,N_18428);
nand U20066 (N_20066,N_14417,N_13545);
nand U20067 (N_20067,N_17901,N_14438);
nand U20068 (N_20068,N_13874,N_18705);
nand U20069 (N_20069,N_13299,N_14607);
nand U20070 (N_20070,N_14462,N_16186);
xor U20071 (N_20071,N_14279,N_18390);
or U20072 (N_20072,N_15259,N_13388);
nor U20073 (N_20073,N_14818,N_14645);
or U20074 (N_20074,N_18018,N_16363);
and U20075 (N_20075,N_14716,N_17982);
or U20076 (N_20076,N_12856,N_14434);
or U20077 (N_20077,N_17769,N_14204);
nand U20078 (N_20078,N_12748,N_14154);
nand U20079 (N_20079,N_15935,N_14464);
or U20080 (N_20080,N_17269,N_14452);
nand U20081 (N_20081,N_15088,N_12611);
and U20082 (N_20082,N_12564,N_17817);
and U20083 (N_20083,N_16847,N_17527);
nor U20084 (N_20084,N_17529,N_14498);
nor U20085 (N_20085,N_13415,N_18458);
nand U20086 (N_20086,N_14467,N_18166);
and U20087 (N_20087,N_16493,N_13674);
nand U20088 (N_20088,N_16119,N_16010);
nand U20089 (N_20089,N_15114,N_18622);
or U20090 (N_20090,N_12972,N_17515);
nor U20091 (N_20091,N_15487,N_12773);
and U20092 (N_20092,N_15834,N_14175);
and U20093 (N_20093,N_12897,N_17322);
nor U20094 (N_20094,N_16216,N_18381);
or U20095 (N_20095,N_18192,N_17462);
and U20096 (N_20096,N_14897,N_13252);
or U20097 (N_20097,N_15028,N_18385);
nor U20098 (N_20098,N_13946,N_14879);
nand U20099 (N_20099,N_16915,N_15994);
xnor U20100 (N_20100,N_15056,N_16581);
and U20101 (N_20101,N_17675,N_13314);
and U20102 (N_20102,N_13798,N_18093);
xor U20103 (N_20103,N_16432,N_16976);
or U20104 (N_20104,N_18426,N_13368);
nor U20105 (N_20105,N_14151,N_13879);
xor U20106 (N_20106,N_16532,N_18429);
nor U20107 (N_20107,N_18489,N_18096);
nand U20108 (N_20108,N_13086,N_14159);
nand U20109 (N_20109,N_16797,N_15411);
and U20110 (N_20110,N_18231,N_14329);
nand U20111 (N_20111,N_13454,N_15288);
or U20112 (N_20112,N_17360,N_18386);
nand U20113 (N_20113,N_17488,N_15675);
nand U20114 (N_20114,N_14931,N_17940);
nand U20115 (N_20115,N_17033,N_16527);
nor U20116 (N_20116,N_14642,N_18213);
xor U20117 (N_20117,N_17898,N_15361);
or U20118 (N_20118,N_18237,N_14618);
xor U20119 (N_20119,N_15769,N_17305);
and U20120 (N_20120,N_18564,N_17260);
or U20121 (N_20121,N_14257,N_18335);
or U20122 (N_20122,N_13891,N_14185);
nor U20123 (N_20123,N_13262,N_16839);
and U20124 (N_20124,N_17683,N_16192);
nor U20125 (N_20125,N_18432,N_12569);
or U20126 (N_20126,N_16200,N_14302);
nand U20127 (N_20127,N_17574,N_16240);
nor U20128 (N_20128,N_15515,N_16689);
and U20129 (N_20129,N_17454,N_18726);
and U20130 (N_20130,N_15537,N_17864);
xor U20131 (N_20131,N_16883,N_15156);
nand U20132 (N_20132,N_14742,N_18146);
nor U20133 (N_20133,N_13613,N_14528);
nand U20134 (N_20134,N_18138,N_17583);
or U20135 (N_20135,N_17288,N_14631);
xnor U20136 (N_20136,N_13281,N_17989);
nand U20137 (N_20137,N_13054,N_17411);
nand U20138 (N_20138,N_13979,N_12579);
and U20139 (N_20139,N_14932,N_12661);
and U20140 (N_20140,N_14021,N_15262);
nand U20141 (N_20141,N_18285,N_13289);
nand U20142 (N_20142,N_18264,N_12588);
nor U20143 (N_20143,N_17983,N_12544);
nor U20144 (N_20144,N_16917,N_16043);
nor U20145 (N_20145,N_18653,N_15782);
nor U20146 (N_20146,N_17430,N_15701);
nand U20147 (N_20147,N_16103,N_14525);
xnor U20148 (N_20148,N_13335,N_15911);
and U20149 (N_20149,N_14127,N_15020);
nor U20150 (N_20150,N_15119,N_14040);
nand U20151 (N_20151,N_14954,N_13972);
nand U20152 (N_20152,N_15822,N_17783);
and U20153 (N_20153,N_16100,N_18034);
nand U20154 (N_20154,N_14715,N_14751);
and U20155 (N_20155,N_12818,N_16389);
nor U20156 (N_20156,N_15392,N_16584);
xnor U20157 (N_20157,N_13600,N_13687);
nor U20158 (N_20158,N_14810,N_13698);
nor U20159 (N_20159,N_15169,N_17885);
or U20160 (N_20160,N_18639,N_18519);
and U20161 (N_20161,N_16212,N_13005);
and U20162 (N_20162,N_14229,N_12507);
nor U20163 (N_20163,N_15651,N_14288);
and U20164 (N_20164,N_13200,N_17106);
xnor U20165 (N_20165,N_15005,N_13720);
nand U20166 (N_20166,N_12591,N_13118);
nor U20167 (N_20167,N_15931,N_18010);
or U20168 (N_20168,N_17268,N_16853);
and U20169 (N_20169,N_14991,N_13462);
and U20170 (N_20170,N_16679,N_14663);
nand U20171 (N_20171,N_17838,N_13236);
nor U20172 (N_20172,N_13605,N_12825);
and U20173 (N_20173,N_15722,N_14889);
and U20174 (N_20174,N_13984,N_12895);
or U20175 (N_20175,N_16305,N_15025);
nand U20176 (N_20176,N_15751,N_17646);
or U20177 (N_20177,N_15727,N_14956);
nand U20178 (N_20178,N_15567,N_13561);
or U20179 (N_20179,N_12706,N_15948);
or U20180 (N_20180,N_16986,N_15200);
nor U20181 (N_20181,N_15247,N_16603);
nor U20182 (N_20182,N_15753,N_16442);
or U20183 (N_20183,N_17883,N_15736);
or U20184 (N_20184,N_13474,N_17159);
or U20185 (N_20185,N_16163,N_17787);
and U20186 (N_20186,N_15226,N_16352);
xnor U20187 (N_20187,N_15915,N_15208);
nor U20188 (N_20188,N_13487,N_16278);
or U20189 (N_20189,N_13491,N_18069);
and U20190 (N_20190,N_16587,N_13386);
and U20191 (N_20191,N_17294,N_13132);
nand U20192 (N_20192,N_15780,N_16741);
nor U20193 (N_20193,N_16896,N_14976);
and U20194 (N_20194,N_13439,N_17832);
xnor U20195 (N_20195,N_16023,N_16952);
or U20196 (N_20196,N_18389,N_17549);
and U20197 (N_20197,N_15623,N_13185);
nand U20198 (N_20198,N_15888,N_14624);
and U20199 (N_20199,N_15573,N_13542);
nand U20200 (N_20200,N_15843,N_13957);
and U20201 (N_20201,N_12936,N_12767);
and U20202 (N_20202,N_16108,N_14429);
nand U20203 (N_20203,N_15927,N_16477);
nor U20204 (N_20204,N_18715,N_15009);
nand U20205 (N_20205,N_15493,N_18305);
or U20206 (N_20206,N_13273,N_18208);
nor U20207 (N_20207,N_18394,N_16514);
nand U20208 (N_20208,N_15136,N_13673);
and U20209 (N_20209,N_16963,N_16399);
and U20210 (N_20210,N_14804,N_17342);
nor U20211 (N_20211,N_18501,N_12650);
xnor U20212 (N_20212,N_15482,N_13098);
xnor U20213 (N_20213,N_18330,N_14148);
and U20214 (N_20214,N_13190,N_14904);
nand U20215 (N_20215,N_15754,N_17059);
nand U20216 (N_20216,N_15999,N_13186);
and U20217 (N_20217,N_15483,N_15201);
xor U20218 (N_20218,N_13934,N_13369);
nor U20219 (N_20219,N_16422,N_15366);
or U20220 (N_20220,N_17658,N_15556);
xnor U20221 (N_20221,N_13077,N_15686);
or U20222 (N_20222,N_16034,N_13810);
nor U20223 (N_20223,N_14220,N_16798);
and U20224 (N_20224,N_13356,N_14894);
nor U20225 (N_20225,N_13804,N_16237);
nor U20226 (N_20226,N_16529,N_15713);
nor U20227 (N_20227,N_15590,N_12942);
or U20228 (N_20228,N_14986,N_17823);
or U20229 (N_20229,N_17636,N_16978);
and U20230 (N_20230,N_14779,N_16868);
nor U20231 (N_20231,N_14205,N_13399);
nor U20232 (N_20232,N_13113,N_16928);
and U20233 (N_20233,N_13228,N_15652);
nor U20234 (N_20234,N_13672,N_14527);
nand U20235 (N_20235,N_17080,N_14192);
nor U20236 (N_20236,N_12520,N_15250);
nand U20237 (N_20237,N_17333,N_18339);
or U20238 (N_20238,N_16251,N_14075);
nand U20239 (N_20239,N_18328,N_16731);
nor U20240 (N_20240,N_15517,N_12659);
and U20241 (N_20241,N_16137,N_16690);
or U20242 (N_20242,N_17525,N_18280);
nand U20243 (N_20243,N_12862,N_15475);
xor U20244 (N_20244,N_15608,N_15876);
or U20245 (N_20245,N_17281,N_13288);
nor U20246 (N_20246,N_17450,N_16740);
nor U20247 (N_20247,N_17748,N_15677);
nor U20248 (N_20248,N_18074,N_18555);
nand U20249 (N_20249,N_14505,N_16012);
or U20250 (N_20250,N_18052,N_13589);
or U20251 (N_20251,N_18091,N_17847);
or U20252 (N_20252,N_18470,N_14813);
nor U20253 (N_20253,N_17754,N_17894);
and U20254 (N_20254,N_16775,N_18745);
and U20255 (N_20255,N_14173,N_13923);
or U20256 (N_20256,N_17447,N_17167);
and U20257 (N_20257,N_15907,N_18020);
or U20258 (N_20258,N_12906,N_13294);
and U20259 (N_20259,N_17860,N_12700);
xor U20260 (N_20260,N_14108,N_13558);
nor U20261 (N_20261,N_17655,N_16233);
xor U20262 (N_20262,N_15726,N_16215);
or U20263 (N_20263,N_17378,N_12729);
and U20264 (N_20264,N_17581,N_15414);
nand U20265 (N_20265,N_14532,N_15151);
or U20266 (N_20266,N_16619,N_14160);
and U20267 (N_20267,N_15458,N_15174);
or U20268 (N_20268,N_13126,N_15030);
xor U20269 (N_20269,N_18553,N_14337);
nand U20270 (N_20270,N_18063,N_18194);
nand U20271 (N_20271,N_15550,N_16826);
and U20272 (N_20272,N_12715,N_13521);
nor U20273 (N_20273,N_17235,N_15863);
or U20274 (N_20274,N_17115,N_16996);
or U20275 (N_20275,N_16824,N_16972);
nor U20276 (N_20276,N_16568,N_16757);
or U20277 (N_20277,N_15539,N_17670);
or U20278 (N_20278,N_13125,N_14653);
nand U20279 (N_20279,N_16267,N_14718);
nand U20280 (N_20280,N_17893,N_14194);
and U20281 (N_20281,N_17842,N_13089);
or U20282 (N_20282,N_15981,N_16013);
or U20283 (N_20283,N_16320,N_16769);
nor U20284 (N_20284,N_16588,N_13567);
nand U20285 (N_20285,N_15839,N_17900);
and U20286 (N_20286,N_15368,N_15738);
xnor U20287 (N_20287,N_12914,N_17944);
and U20288 (N_20288,N_17483,N_14872);
nor U20289 (N_20289,N_17014,N_18001);
and U20290 (N_20290,N_16458,N_15836);
nand U20291 (N_20291,N_17564,N_17409);
nand U20292 (N_20292,N_13357,N_12903);
nand U20293 (N_20293,N_17239,N_14815);
nor U20294 (N_20294,N_15591,N_17602);
nand U20295 (N_20295,N_14910,N_16148);
nand U20296 (N_20296,N_12501,N_14006);
or U20297 (N_20297,N_15798,N_14728);
and U20298 (N_20298,N_13777,N_18165);
or U20299 (N_20299,N_16412,N_17704);
nand U20300 (N_20300,N_15502,N_16844);
or U20301 (N_20301,N_15619,N_17349);
nor U20302 (N_20302,N_13162,N_16112);
nand U20303 (N_20303,N_12723,N_16386);
and U20304 (N_20304,N_12530,N_15792);
nor U20305 (N_20305,N_14100,N_18362);
or U20306 (N_20306,N_14457,N_12561);
and U20307 (N_20307,N_14286,N_17413);
or U20308 (N_20308,N_14143,N_17009);
or U20309 (N_20309,N_18498,N_12695);
or U20310 (N_20310,N_17949,N_13382);
and U20311 (N_20311,N_16296,N_18079);
or U20312 (N_20312,N_14547,N_14425);
nor U20313 (N_20313,N_16993,N_12752);
or U20314 (N_20314,N_14048,N_16339);
and U20315 (N_20315,N_17644,N_14240);
nor U20316 (N_20316,N_12572,N_15079);
or U20317 (N_20317,N_17295,N_12545);
and U20318 (N_20318,N_17509,N_12529);
or U20319 (N_20319,N_17537,N_13372);
nor U20320 (N_20320,N_14406,N_18130);
nor U20321 (N_20321,N_14176,N_17507);
nand U20322 (N_20322,N_14010,N_13301);
or U20323 (N_20323,N_15985,N_12961);
nor U20324 (N_20324,N_13359,N_15570);
nand U20325 (N_20325,N_14862,N_15642);
and U20326 (N_20326,N_16494,N_17422);
xor U20327 (N_20327,N_16577,N_13516);
nand U20328 (N_20328,N_14626,N_16903);
or U20329 (N_20329,N_16143,N_17451);
and U20330 (N_20330,N_16618,N_14773);
or U20331 (N_20331,N_16800,N_15795);
nor U20332 (N_20332,N_15635,N_13400);
xor U20333 (N_20333,N_16728,N_15240);
nand U20334 (N_20334,N_14938,N_12728);
nor U20335 (N_20335,N_12612,N_15276);
xnor U20336 (N_20336,N_15787,N_12600);
nor U20337 (N_20337,N_14217,N_17988);
and U20338 (N_20338,N_16416,N_14705);
or U20339 (N_20339,N_14007,N_12958);
xnor U20340 (N_20340,N_18224,N_15568);
and U20341 (N_20341,N_13670,N_12526);
and U20342 (N_20342,N_16805,N_16788);
and U20343 (N_20343,N_16660,N_14264);
or U20344 (N_20344,N_14320,N_13626);
or U20345 (N_20345,N_17187,N_12848);
or U20346 (N_20346,N_17062,N_16070);
or U20347 (N_20347,N_15627,N_14521);
and U20348 (N_20348,N_16053,N_15057);
nor U20349 (N_20349,N_16203,N_16784);
nand U20350 (N_20350,N_17501,N_17219);
xnor U20351 (N_20351,N_13045,N_15133);
xnor U20352 (N_20352,N_15406,N_12971);
nor U20353 (N_20353,N_14402,N_18080);
nand U20354 (N_20354,N_18359,N_14276);
nand U20355 (N_20355,N_16333,N_18374);
nor U20356 (N_20356,N_17332,N_13023);
and U20357 (N_20357,N_15891,N_13139);
and U20358 (N_20358,N_17300,N_13254);
nand U20359 (N_20359,N_16704,N_12744);
and U20360 (N_20360,N_13741,N_16714);
nor U20361 (N_20361,N_13599,N_12657);
xor U20362 (N_20362,N_15669,N_16921);
or U20363 (N_20363,N_15966,N_14404);
nand U20364 (N_20364,N_13109,N_16076);
and U20365 (N_20365,N_14647,N_16632);
and U20366 (N_20366,N_12553,N_15667);
and U20367 (N_20367,N_13366,N_18267);
or U20368 (N_20368,N_17567,N_13463);
and U20369 (N_20369,N_14181,N_17247);
or U20370 (N_20370,N_17324,N_15930);
or U20371 (N_20371,N_18265,N_13144);
or U20372 (N_20372,N_13231,N_14222);
nand U20373 (N_20373,N_15348,N_12844);
and U20374 (N_20374,N_17919,N_13284);
nor U20375 (N_20375,N_16113,N_14630);
or U20376 (N_20376,N_12543,N_13996);
xnor U20377 (N_20377,N_13295,N_12727);
nand U20378 (N_20378,N_13894,N_17647);
xor U20379 (N_20379,N_16327,N_16792);
or U20380 (N_20380,N_14923,N_16177);
nor U20381 (N_20381,N_14129,N_15459);
nor U20382 (N_20382,N_14249,N_14696);
nor U20383 (N_20383,N_16084,N_15234);
or U20384 (N_20384,N_13313,N_16691);
nor U20385 (N_20385,N_18516,N_15820);
nor U20386 (N_20386,N_18248,N_17674);
and U20387 (N_20387,N_17056,N_13895);
nor U20388 (N_20388,N_12974,N_13608);
nand U20389 (N_20389,N_15418,N_13887);
xor U20390 (N_20390,N_18635,N_13759);
nor U20391 (N_20391,N_14018,N_18632);
nor U20392 (N_20392,N_12978,N_17073);
nand U20393 (N_20393,N_17370,N_17916);
or U20394 (N_20394,N_15159,N_15101);
nand U20395 (N_20395,N_15454,N_15924);
nor U20396 (N_20396,N_14990,N_17414);
xnor U20397 (N_20397,N_13112,N_15659);
and U20398 (N_20398,N_16395,N_17604);
and U20399 (N_20399,N_16898,N_17788);
or U20400 (N_20400,N_13936,N_16558);
nor U20401 (N_20401,N_17351,N_17081);
or U20402 (N_20402,N_16302,N_18583);
nand U20403 (N_20403,N_18333,N_13628);
nand U20404 (N_20404,N_16046,N_12648);
and U20405 (N_20405,N_16220,N_13093);
nand U20406 (N_20406,N_15919,N_14047);
nand U20407 (N_20407,N_15227,N_14446);
nand U20408 (N_20408,N_16179,N_13812);
nor U20409 (N_20409,N_12968,N_17052);
and U20410 (N_20410,N_18647,N_14740);
and U20411 (N_20411,N_12875,N_16091);
and U20412 (N_20412,N_17152,N_17709);
nand U20413 (N_20413,N_17510,N_13991);
or U20414 (N_20414,N_16935,N_16869);
nand U20415 (N_20415,N_13059,N_13762);
nor U20416 (N_20416,N_16006,N_13265);
or U20417 (N_20417,N_16002,N_16123);
or U20418 (N_20418,N_14443,N_15175);
nor U20419 (N_20419,N_15520,N_17217);
or U20420 (N_20420,N_14733,N_14182);
nand U20421 (N_20421,N_18548,N_13129);
and U20422 (N_20422,N_13630,N_18135);
nor U20423 (N_20423,N_13588,N_18284);
and U20424 (N_20424,N_17732,N_18589);
nor U20425 (N_20425,N_12704,N_15322);
and U20426 (N_20426,N_13389,N_13629);
xor U20427 (N_20427,N_12979,N_16893);
or U20428 (N_20428,N_13079,N_12517);
nand U20429 (N_20429,N_14221,N_13831);
nand U20430 (N_20430,N_18126,N_17976);
and U20431 (N_20431,N_12935,N_16451);
or U20432 (N_20432,N_13612,N_17535);
nand U20433 (N_20433,N_16334,N_17784);
nor U20434 (N_20434,N_18406,N_18141);
or U20435 (N_20435,N_18083,N_15451);
or U20436 (N_20436,N_12631,N_15154);
and U20437 (N_20437,N_17266,N_18357);
nand U20438 (N_20438,N_17651,N_13220);
nand U20439 (N_20439,N_13652,N_17967);
nor U20440 (N_20440,N_16987,N_18283);
nand U20441 (N_20441,N_17084,N_17639);
nor U20442 (N_20442,N_18316,N_14117);
or U20443 (N_20443,N_15126,N_17978);
or U20444 (N_20444,N_13549,N_14482);
or U20445 (N_20445,N_15367,N_15699);
or U20446 (N_20446,N_16083,N_18592);
xor U20447 (N_20447,N_15155,N_13575);
and U20448 (N_20448,N_13531,N_16785);
and U20449 (N_20449,N_18508,N_13390);
nor U20450 (N_20450,N_12779,N_15759);
or U20451 (N_20451,N_14041,N_15229);
nor U20452 (N_20452,N_15063,N_17435);
or U20453 (N_20453,N_15516,N_17487);
or U20454 (N_20454,N_14012,N_15007);
nor U20455 (N_20455,N_17888,N_17023);
nand U20456 (N_20456,N_16285,N_16870);
and U20457 (N_20457,N_18490,N_15315);
or U20458 (N_20458,N_13352,N_17731);
nor U20459 (N_20459,N_12790,N_13864);
and U20460 (N_20460,N_13721,N_16746);
or U20461 (N_20461,N_17688,N_15160);
nand U20462 (N_20462,N_15855,N_15917);
or U20463 (N_20463,N_16612,N_12757);
nor U20464 (N_20464,N_17321,N_14851);
or U20465 (N_20465,N_14212,N_14184);
nand U20466 (N_20466,N_17773,N_13853);
or U20467 (N_20467,N_12654,N_16591);
and U20468 (N_20468,N_16008,N_14759);
and U20469 (N_20469,N_15123,N_14158);
or U20470 (N_20470,N_13858,N_16538);
and U20471 (N_20471,N_16021,N_16702);
xor U20472 (N_20472,N_15324,N_13898);
nand U20473 (N_20473,N_15707,N_13140);
xor U20474 (N_20474,N_16524,N_17347);
nand U20475 (N_20475,N_17265,N_18610);
nor U20476 (N_20476,N_12833,N_15824);
nand U20477 (N_20477,N_13534,N_18358);
nand U20478 (N_20478,N_14132,N_12858);
or U20479 (N_20479,N_13758,N_12859);
nor U20480 (N_20480,N_12717,N_17820);
nand U20481 (N_20481,N_16270,N_12746);
nor U20482 (N_20482,N_18282,N_15246);
xor U20483 (N_20483,N_13873,N_17576);
nand U20484 (N_20484,N_17934,N_14363);
and U20485 (N_20485,N_16415,N_13625);
nor U20486 (N_20486,N_18286,N_15557);
nor U20487 (N_20487,N_14627,N_18731);
xor U20488 (N_20488,N_15326,N_12785);
nand U20489 (N_20489,N_17145,N_18616);
xnor U20490 (N_20490,N_17174,N_12672);
and U20491 (N_20491,N_16767,N_14390);
nand U20492 (N_20492,N_17981,N_18011);
and U20493 (N_20493,N_16040,N_14261);
and U20494 (N_20494,N_16362,N_13977);
and U20495 (N_20495,N_13684,N_15545);
nand U20496 (N_20496,N_15428,N_16665);
nor U20497 (N_20497,N_14678,N_13896);
and U20498 (N_20498,N_15300,N_18311);
nand U20499 (N_20499,N_15549,N_14562);
or U20500 (N_20500,N_16891,N_16733);
nor U20501 (N_20501,N_13307,N_13283);
or U20502 (N_20502,N_16402,N_18067);
and U20503 (N_20503,N_14592,N_16226);
and U20504 (N_20504,N_13013,N_13165);
nand U20505 (N_20505,N_15354,N_16911);
and U20506 (N_20506,N_14001,N_18545);
or U20507 (N_20507,N_17928,N_17132);
nand U20508 (N_20508,N_16574,N_16232);
nand U20509 (N_20509,N_17079,N_17301);
nor U20510 (N_20510,N_16274,N_14798);
nor U20511 (N_20511,N_17846,N_18425);
nand U20512 (N_20512,N_17707,N_15282);
and U20513 (N_20513,N_12798,N_16942);
and U20514 (N_20514,N_17701,N_17480);
nor U20515 (N_20515,N_16715,N_18493);
nor U20516 (N_20516,N_13398,N_17010);
nor U20517 (N_20517,N_15245,N_17334);
or U20518 (N_20518,N_16038,N_15423);
and U20519 (N_20519,N_17331,N_14210);
nand U20520 (N_20520,N_17722,N_12872);
nand U20521 (N_20521,N_16183,N_13195);
nand U20522 (N_20522,N_14501,N_18343);
or U20523 (N_20523,N_15284,N_17608);
nand U20524 (N_20524,N_13649,N_13987);
or U20525 (N_20525,N_18687,N_17531);
and U20526 (N_20526,N_13309,N_16900);
nand U20527 (N_20527,N_16474,N_13958);
nand U20528 (N_20528,N_18185,N_18405);
and U20529 (N_20529,N_15893,N_14057);
nand U20530 (N_20530,N_13488,N_18740);
or U20531 (N_20531,N_16977,N_16495);
or U20532 (N_20532,N_16820,N_15504);
or U20533 (N_20533,N_18099,N_15629);
and U20534 (N_20534,N_16818,N_15870);
and U20535 (N_20535,N_16596,N_15605);
or U20536 (N_20536,N_17030,N_14193);
or U20537 (N_20537,N_12878,N_17419);
or U20538 (N_20538,N_15400,N_13303);
nand U20539 (N_20539,N_17814,N_14839);
and U20540 (N_20540,N_18748,N_15485);
nand U20541 (N_20541,N_12938,N_17594);
or U20542 (N_20542,N_18674,N_17621);
nand U20543 (N_20543,N_17987,N_17292);
nand U20544 (N_20544,N_18371,N_16453);
or U20545 (N_20545,N_16752,N_17190);
or U20546 (N_20546,N_18214,N_17694);
nor U20547 (N_20547,N_13256,N_14340);
nor U20548 (N_20548,N_13494,N_15962);
nand U20549 (N_20549,N_16899,N_18259);
nor U20550 (N_20550,N_13660,N_12915);
nand U20551 (N_20551,N_16265,N_15729);
or U20552 (N_20552,N_14263,N_17388);
nand U20553 (N_20553,N_15181,N_17954);
xor U20554 (N_20554,N_16563,N_15457);
or U20555 (N_20555,N_14088,N_14306);
nand U20556 (N_20556,N_13421,N_17829);
or U20557 (N_20557,N_15138,N_15548);
xnor U20558 (N_20558,N_14857,N_17836);
nand U20559 (N_20559,N_17273,N_12772);
nand U20560 (N_20560,N_17905,N_15563);
nand U20561 (N_20561,N_15918,N_16646);
and U20562 (N_20562,N_17947,N_18170);
and U20563 (N_20563,N_16466,N_14664);
and U20564 (N_20564,N_14147,N_16051);
or U20565 (N_20565,N_14384,N_15643);
and U20566 (N_20566,N_13009,N_16806);
nor U20567 (N_20567,N_15237,N_15577);
nand U20568 (N_20568,N_14354,N_16959);
nand U20569 (N_20569,N_17221,N_13866);
and U20570 (N_20570,N_14016,N_18058);
and U20571 (N_20571,N_17764,N_13104);
nor U20572 (N_20572,N_16261,N_14660);
xnor U20573 (N_20573,N_13771,N_17668);
nand U20574 (N_20574,N_14617,N_17330);
nand U20575 (N_20575,N_16680,N_18529);
nand U20576 (N_20576,N_15397,N_15462);
nand U20577 (N_20577,N_16719,N_16909);
nor U20578 (N_20578,N_12557,N_14727);
xor U20579 (N_20579,N_18245,N_14364);
or U20580 (N_20580,N_13189,N_15260);
nor U20581 (N_20581,N_14896,N_13994);
and U20582 (N_20582,N_15786,N_17374);
and U20583 (N_20583,N_17999,N_16947);
nand U20584 (N_20584,N_15387,N_17203);
or U20585 (N_20585,N_16238,N_12855);
or U20586 (N_20586,N_12857,N_18124);
nand U20587 (N_20587,N_16236,N_18132);
nor U20588 (N_20588,N_17044,N_17697);
or U20589 (N_20589,N_14567,N_14495);
or U20590 (N_20590,N_16667,N_13945);
or U20591 (N_20591,N_13026,N_14598);
or U20592 (N_20592,N_14483,N_13053);
nand U20593 (N_20593,N_16652,N_16565);
or U20594 (N_20594,N_18000,N_16281);
and U20595 (N_20595,N_13275,N_15172);
xor U20596 (N_20596,N_13795,N_18403);
nor U20597 (N_20597,N_14816,N_15731);
or U20598 (N_20598,N_13145,N_15588);
and U20599 (N_20599,N_16770,N_17862);
and U20600 (N_20600,N_16946,N_13341);
or U20601 (N_20601,N_18439,N_14883);
and U20602 (N_20602,N_16576,N_18129);
or U20603 (N_20603,N_14499,N_17421);
and U20604 (N_20604,N_16465,N_18691);
nand U20605 (N_20605,N_13959,N_13645);
or U20606 (N_20606,N_18724,N_12834);
and U20607 (N_20607,N_15332,N_13906);
and U20608 (N_20608,N_16991,N_16288);
and U20609 (N_20609,N_17175,N_15031);
and U20610 (N_20610,N_15756,N_16602);
or U20611 (N_20611,N_15488,N_15996);
nor U20612 (N_20612,N_18474,N_14051);
xnor U20613 (N_20613,N_17278,N_15748);
xor U20614 (N_20614,N_14459,N_18255);
nor U20615 (N_20615,N_14195,N_15018);
or U20616 (N_20616,N_17158,N_17353);
and U20617 (N_20617,N_17822,N_14803);
nor U20618 (N_20618,N_14787,N_12917);
nand U20619 (N_20619,N_16307,N_17826);
nand U20620 (N_20620,N_13784,N_17099);
or U20621 (N_20621,N_17514,N_16444);
and U20622 (N_20622,N_13473,N_15864);
xnor U20623 (N_20623,N_16499,N_18278);
nand U20624 (N_20624,N_14453,N_14671);
or U20625 (N_20625,N_15980,N_16468);
and U20626 (N_20626,N_15857,N_18452);
and U20627 (N_20627,N_12829,N_15763);
and U20628 (N_20628,N_12871,N_13044);
xnor U20629 (N_20629,N_12888,N_14900);
and U20630 (N_20630,N_17359,N_16289);
nand U20631 (N_20631,N_16523,N_14980);
nor U20632 (N_20632,N_16753,N_14266);
and U20633 (N_20633,N_15014,N_18149);
nor U20634 (N_20634,N_13578,N_13519);
or U20635 (N_20635,N_13668,N_14199);
nor U20636 (N_20636,N_14745,N_15875);
or U20637 (N_20637,N_18645,N_17856);
or U20638 (N_20638,N_15694,N_15654);
or U20639 (N_20639,N_17226,N_14959);
nor U20640 (N_20640,N_15058,N_17053);
nand U20641 (N_20641,N_16134,N_17691);
nor U20642 (N_20642,N_17463,N_14655);
or U20643 (N_20643,N_18225,N_14873);
and U20644 (N_20644,N_18659,N_13088);
and U20645 (N_20645,N_17727,N_13041);
nor U20646 (N_20646,N_16599,N_16552);
xnor U20647 (N_20647,N_15598,N_17338);
nor U20648 (N_20648,N_12690,N_16202);
and U20649 (N_20649,N_16088,N_12887);
nor U20650 (N_20650,N_16221,N_17866);
xor U20651 (N_20651,N_18121,N_16341);
or U20652 (N_20652,N_16064,N_16292);
xor U20653 (N_20653,N_17195,N_13993);
xnor U20654 (N_20654,N_14351,N_12845);
and U20655 (N_20655,N_15470,N_17279);
and U20656 (N_20656,N_13590,N_14649);
or U20657 (N_20657,N_13947,N_13127);
nand U20658 (N_20658,N_14833,N_16151);
nand U20659 (N_20659,N_15689,N_18232);
nand U20660 (N_20660,N_17042,N_12687);
nand U20661 (N_20661,N_13669,N_15929);
and U20662 (N_20662,N_15615,N_14105);
nor U20663 (N_20663,N_14529,N_15207);
or U20664 (N_20664,N_15831,N_18294);
nand U20665 (N_20665,N_14634,N_12775);
xor U20666 (N_20666,N_16125,N_18169);
and U20667 (N_20667,N_17851,N_13803);
or U20668 (N_20668,N_12990,N_18064);
nor U20669 (N_20669,N_13918,N_12807);
nor U20670 (N_20670,N_16879,N_17876);
nor U20671 (N_20671,N_18158,N_13477);
xnor U20672 (N_20672,N_15489,N_13870);
nand U20673 (N_20673,N_17743,N_15902);
nor U20674 (N_20674,N_14339,N_17151);
and U20675 (N_20675,N_14799,N_16765);
and U20676 (N_20676,N_13258,N_16140);
or U20677 (N_20677,N_18417,N_13701);
nor U20678 (N_20678,N_16713,N_13325);
nor U20679 (N_20679,N_13638,N_14713);
nor U20680 (N_20680,N_18279,N_14488);
nor U20681 (N_20681,N_14247,N_14629);
or U20682 (N_20682,N_18028,N_16222);
nand U20683 (N_20683,N_14440,N_14795);
nor U20684 (N_20684,N_14531,N_12988);
and U20685 (N_20685,N_17309,N_14395);
nand U20686 (N_20686,N_15920,N_17245);
nor U20687 (N_20687,N_14144,N_16517);
xor U20688 (N_20688,N_16197,N_12578);
nand U20689 (N_20689,N_12984,N_13835);
nor U20690 (N_20690,N_14191,N_17326);
and U20691 (N_20691,N_13148,N_14981);
and U20692 (N_20692,N_13479,N_13174);
and U20693 (N_20693,N_14824,N_14540);
nor U20694 (N_20694,N_12956,N_17685);
xnor U20695 (N_20695,N_16867,N_13100);
nand U20696 (N_20696,N_16011,N_18615);
nor U20697 (N_20697,N_17994,N_14411);
xor U20698 (N_20698,N_15064,N_16951);
and U20699 (N_20699,N_17389,N_14063);
nor U20700 (N_20700,N_17039,N_18089);
nor U20701 (N_20701,N_18373,N_13783);
nand U20702 (N_20702,N_15188,N_12802);
xnor U20703 (N_20703,N_15901,N_15330);
and U20704 (N_20704,N_18227,N_18218);
and U20705 (N_20705,N_17733,N_13682);
or U20706 (N_20706,N_13790,N_18459);
nand U20707 (N_20707,N_18546,N_13667);
xnor U20708 (N_20708,N_18677,N_14167);
or U20709 (N_20709,N_18239,N_12966);
xor U20710 (N_20710,N_15971,N_16965);
and U20711 (N_20711,N_13990,N_12504);
and U20712 (N_20712,N_17199,N_13155);
nor U20713 (N_20713,N_17236,N_14963);
and U20714 (N_20714,N_16661,N_17986);
xnor U20715 (N_20715,N_18356,N_13743);
nor U20716 (N_20716,N_15310,N_15432);
or U20717 (N_20717,N_18337,N_14843);
or U20718 (N_20718,N_16717,N_16662);
nand U20719 (N_20719,N_14524,N_15871);
and U20720 (N_20720,N_18045,N_12983);
nor U20721 (N_20721,N_13033,N_17066);
nor U20722 (N_20722,N_16497,N_16994);
and U20723 (N_20723,N_17393,N_14046);
and U20724 (N_20724,N_15347,N_16185);
nand U20725 (N_20725,N_14061,N_17927);
or U20726 (N_20726,N_14609,N_16418);
or U20727 (N_20727,N_17244,N_17166);
nand U20728 (N_20728,N_14271,N_16884);
nor U20729 (N_20729,N_16057,N_16207);
nand U20730 (N_20730,N_18086,N_14536);
or U20731 (N_20731,N_16433,N_15775);
and U20732 (N_20732,N_14435,N_16549);
and U20733 (N_20733,N_16506,N_14055);
nor U20734 (N_20734,N_12580,N_13732);
or U20735 (N_20735,N_14500,N_16866);
nor U20736 (N_20736,N_13878,N_17959);
and U20737 (N_20737,N_16262,N_18717);
nor U20738 (N_20738,N_16384,N_13156);
xor U20739 (N_20739,N_13778,N_18281);
nor U20740 (N_20740,N_12943,N_15936);
nor U20741 (N_20741,N_15805,N_15096);
xnor U20742 (N_20742,N_17588,N_16555);
nor U20743 (N_20743,N_12786,N_13529);
nor U20744 (N_20744,N_14967,N_16700);
nor U20745 (N_20745,N_16284,N_15287);
nor U20746 (N_20746,N_15419,N_15334);
and U20747 (N_20747,N_15416,N_13173);
nor U20748 (N_20748,N_15522,N_13318);
nor U20749 (N_20749,N_13956,N_13718);
nand U20750 (N_20750,N_15500,N_17721);
nor U20751 (N_20751,N_12619,N_17405);
nor U20752 (N_20752,N_13103,N_17831);
or U20753 (N_20753,N_15755,N_15069);
nor U20754 (N_20754,N_15072,N_12644);
nand U20755 (N_20755,N_15967,N_16727);
and U20756 (N_20756,N_16136,N_13282);
nor U20757 (N_20757,N_14102,N_14983);
xnor U20758 (N_20758,N_13010,N_16848);
nor U20759 (N_20759,N_12963,N_13842);
nand U20760 (N_20760,N_12883,N_14474);
nand U20761 (N_20761,N_16462,N_13191);
or U20762 (N_20762,N_16890,N_14930);
and U20763 (N_20763,N_12916,N_13663);
xor U20764 (N_20764,N_16235,N_18269);
or U20765 (N_20765,N_15218,N_17259);
and U20766 (N_20766,N_13349,N_16804);
nand U20767 (N_20767,N_15214,N_12816);
or U20768 (N_20768,N_16441,N_18150);
nand U20769 (N_20769,N_15268,N_18512);
nand U20770 (N_20770,N_17164,N_12620);
nor U20771 (N_20771,N_13371,N_12898);
nor U20772 (N_20772,N_17872,N_14037);
nand U20773 (N_20773,N_13016,N_17573);
xnor U20774 (N_20774,N_15819,N_17046);
xnor U20775 (N_20775,N_16701,N_12685);
xor U20776 (N_20776,N_17570,N_16533);
nand U20777 (N_20777,N_12835,N_13083);
nand U20778 (N_20778,N_15765,N_16321);
or U20779 (N_20779,N_15862,N_18631);
or U20780 (N_20780,N_14269,N_15292);
nor U20781 (N_20781,N_15956,N_13572);
and U20782 (N_20782,N_15714,N_14489);
nand U20783 (N_20783,N_17728,N_15498);
or U20784 (N_20784,N_16592,N_14854);
or U20785 (N_20785,N_14837,N_14752);
or U20786 (N_20786,N_13306,N_15076);
nor U20787 (N_20787,N_14831,N_17696);
nand U20788 (N_20788,N_15417,N_14998);
and U20789 (N_20789,N_16365,N_16814);
and U20790 (N_20790,N_16213,N_12828);
nand U20791 (N_20791,N_15655,N_15364);
nand U20792 (N_20792,N_13603,N_14456);
or U20793 (N_20793,N_17379,N_16111);
and U20794 (N_20794,N_14996,N_15219);
nor U20795 (N_20795,N_14729,N_16086);
nand U20796 (N_20796,N_13204,N_18569);
nor U20797 (N_20797,N_17749,N_17825);
or U20798 (N_20798,N_15001,N_15168);
or U20799 (N_20799,N_13785,N_13022);
or U20800 (N_20800,N_18477,N_18510);
nor U20801 (N_20801,N_13396,N_14035);
xor U20802 (N_20802,N_15684,N_13933);
nand U20803 (N_20803,N_15997,N_18152);
nor U20804 (N_20804,N_13266,N_13637);
or U20805 (N_20805,N_16536,N_15273);
or U20806 (N_20806,N_13154,N_15531);
and U20807 (N_20807,N_15565,N_17806);
or U20808 (N_20808,N_14251,N_18400);
or U20809 (N_20809,N_16425,N_15437);
or U20810 (N_20810,N_15216,N_14587);
or U20811 (N_20811,N_14788,N_18387);
and U20812 (N_20812,N_17149,N_13604);
xor U20813 (N_20813,N_13056,N_15265);
nor U20814 (N_20814,N_18595,N_13690);
or U20815 (N_20815,N_15640,N_15346);
nor U20816 (N_20816,N_16999,N_13308);
and U20817 (N_20817,N_18603,N_14497);
nor U20818 (N_20818,N_13999,N_17197);
or U20819 (N_20819,N_17210,N_17730);
or U20820 (N_20820,N_15507,N_13515);
and U20821 (N_20821,N_18625,N_15116);
nor U20822 (N_20822,N_15886,N_16279);
or U20823 (N_20823,N_16790,N_13065);
or U20824 (N_20824,N_18250,N_15628);
nor U20825 (N_20825,N_13465,N_14641);
xor U20826 (N_20826,N_16676,N_13268);
nand U20827 (N_20827,N_15937,N_17310);
and U20828 (N_20828,N_16353,N_15293);
and U20829 (N_20829,N_18044,N_14293);
nor U20830 (N_20830,N_13924,N_18029);
and U20831 (N_20831,N_17520,N_13893);
and U20832 (N_20832,N_12995,N_14866);
nand U20833 (N_20833,N_14180,N_13815);
nand U20834 (N_20834,N_13881,N_17240);
nand U20835 (N_20835,N_14104,N_17513);
xor U20836 (N_20836,N_15816,N_12607);
xnor U20837 (N_20837,N_13017,N_17686);
or U20838 (N_20838,N_14188,N_18187);
or U20839 (N_20839,N_16087,N_14707);
or U20840 (N_20840,N_15509,N_17684);
nor U20841 (N_20841,N_18690,N_15044);
and U20842 (N_20842,N_18409,N_17027);
and U20843 (N_20843,N_17156,N_18594);
and U20844 (N_20844,N_18716,N_18608);
nor U20845 (N_20845,N_15258,N_15430);
nand U20846 (N_20846,N_15165,N_17246);
or U20847 (N_20847,N_14496,N_12780);
nand U20848 (N_20848,N_13470,N_12764);
nand U20849 (N_20849,N_15912,N_13847);
or U20850 (N_20850,N_13748,N_16707);
nand U20851 (N_20851,N_17964,N_17453);
nand U20852 (N_20852,N_15283,N_14580);
and U20853 (N_20853,N_14682,N_12667);
or U20854 (N_20854,N_15299,N_16961);
nor U20855 (N_20855,N_14444,N_17050);
nor U20856 (N_20856,N_18161,N_17854);
nor U20857 (N_20857,N_16241,N_18483);
or U20858 (N_20858,N_18434,N_13338);
and U20859 (N_20859,N_17936,N_13641);
nand U20860 (N_20860,N_13502,N_16455);
nor U20861 (N_20861,N_16311,N_13537);
xor U20862 (N_20862,N_16744,N_13511);
nand U20863 (N_20863,N_18065,N_17495);
nor U20864 (N_20864,N_16189,N_18349);
nor U20865 (N_20865,N_12921,N_18134);
nor U20866 (N_20866,N_13522,N_15032);
or U20867 (N_20867,N_15089,N_18207);
nand U20868 (N_20868,N_14884,N_13330);
nor U20869 (N_20869,N_18440,N_15469);
and U20870 (N_20870,N_17469,N_12632);
and U20871 (N_20871,N_16934,N_15345);
nor U20872 (N_20872,N_17741,N_13128);
xnor U20873 (N_20873,N_12633,N_17843);
or U20874 (N_20874,N_17682,N_16017);
nand U20875 (N_20875,N_18696,N_13142);
nor U20876 (N_20876,N_18397,N_14163);
xnor U20877 (N_20877,N_16598,N_16318);
and U20878 (N_20878,N_15130,N_15148);
or U20879 (N_20879,N_15661,N_17479);
nand U20880 (N_20880,N_12980,N_13766);
and U20881 (N_20881,N_17401,N_14284);
nand U20882 (N_20882,N_14552,N_17224);
or U20883 (N_20883,N_15370,N_13576);
or U20884 (N_20884,N_16066,N_17740);
nand U20885 (N_20885,N_15093,N_13686);
or U20886 (N_20886,N_17282,N_13326);
xor U20887 (N_20887,N_16567,N_15708);
xor U20888 (N_20888,N_16537,N_14324);
nand U20889 (N_20889,N_18201,N_14067);
or U20890 (N_20890,N_14433,N_14917);
or U20891 (N_20891,N_15314,N_16849);
and U20892 (N_20892,N_14149,N_16621);
nor U20893 (N_20893,N_18609,N_12886);
or U20894 (N_20894,N_13409,N_14372);
or U20895 (N_20895,N_14131,N_14397);
nor U20896 (N_20896,N_18315,N_16894);
or U20897 (N_20897,N_12536,N_12714);
and U20898 (N_20898,N_15495,N_16219);
nand U20899 (N_20899,N_18145,N_15305);
nand U20900 (N_20900,N_17970,N_13105);
nand U20901 (N_20901,N_15575,N_13379);
or U20902 (N_20902,N_18670,N_16551);
or U20903 (N_20903,N_18015,N_14730);
nand U20904 (N_20904,N_13978,N_15389);
or U20905 (N_20905,N_13830,N_14820);
xor U20906 (N_20906,N_12912,N_18363);
nor U20907 (N_20907,N_14661,N_13897);
nand U20908 (N_20908,N_18351,N_16045);
and U20909 (N_20909,N_14677,N_14604);
nor U20910 (N_20910,N_13035,N_17502);
and U20911 (N_20911,N_17723,N_13712);
nand U20912 (N_20912,N_14690,N_15609);
and U20913 (N_20913,N_17377,N_13813);
nand U20914 (N_20914,N_12928,N_16077);
and U20915 (N_20915,N_15023,N_13526);
nor U20916 (N_20916,N_14611,N_15006);
nor U20917 (N_20917,N_14714,N_12647);
nand U20918 (N_20918,N_16464,N_13224);
nand U20919 (N_20919,N_17815,N_12668);
or U20920 (N_20920,N_14315,N_16342);
or U20921 (N_20921,N_18007,N_16653);
nor U20922 (N_20922,N_17600,N_13530);
and U20923 (N_20923,N_13291,N_12997);
nor U20924 (N_20924,N_18713,N_13248);
xnor U20925 (N_20925,N_12655,N_15412);
and U20926 (N_20926,N_17974,N_15552);
nand U20927 (N_20927,N_12969,N_14083);
nand U20928 (N_20928,N_13607,N_17666);
nand U20929 (N_20929,N_14248,N_14262);
nand U20930 (N_20930,N_15195,N_12594);
nor U20931 (N_20931,N_16319,N_13402);
nor U20932 (N_20932,N_18591,N_14486);
nand U20933 (N_20933,N_12679,N_13774);
nand U20934 (N_20934,N_13837,N_18035);
nor U20935 (N_20935,N_16954,N_14215);
nand U20936 (N_20936,N_17058,N_17745);
nand U20937 (N_20937,N_16349,N_16250);
or U20938 (N_20938,N_15528,N_14056);
nor U20939 (N_20939,N_18711,N_12852);
nand U20940 (N_20940,N_15601,N_15740);
xnor U20941 (N_20941,N_14036,N_16150);
and U20942 (N_20942,N_15884,N_18309);
xor U20943 (N_20943,N_15943,N_15270);
nand U20944 (N_20944,N_15928,N_14858);
or U20945 (N_20945,N_16483,N_16379);
or U20946 (N_20946,N_15410,N_17490);
and U20947 (N_20947,N_13819,N_17306);
nor U20948 (N_20948,N_17812,N_16015);
nand U20949 (N_20949,N_17406,N_13610);
nand U20950 (N_20950,N_16383,N_16120);
xor U20951 (N_20951,N_16666,N_17440);
or U20952 (N_20952,N_16802,N_12589);
and U20953 (N_20953,N_17272,N_15564);
xnor U20954 (N_20954,N_16239,N_14076);
and U20955 (N_20955,N_12665,N_13374);
and U20956 (N_20956,N_14170,N_12737);
or U20957 (N_20957,N_18719,N_12636);
nand U20958 (N_20958,N_18524,N_17552);
nor U20959 (N_20959,N_12581,N_12861);
xnor U20960 (N_20960,N_15379,N_17399);
and U20961 (N_20961,N_18455,N_15589);
xor U20962 (N_20962,N_18106,N_12608);
and U20963 (N_20963,N_12678,N_13395);
nor U20964 (N_20964,N_14358,N_14139);
nor U20965 (N_20965,N_14230,N_15538);
nand U20966 (N_20966,N_16097,N_14648);
nor U20967 (N_20967,N_17737,N_14137);
nand U20968 (N_20968,N_16938,N_18336);
and U20969 (N_20969,N_13939,N_18500);
and U20970 (N_20970,N_18411,N_13032);
or U20971 (N_20971,N_16794,N_12734);
nor U20972 (N_20972,N_13152,N_16712);
xnor U20973 (N_20973,N_18532,N_17270);
xor U20974 (N_20974,N_15239,N_12616);
and U20975 (N_20975,N_18215,N_15853);
xor U20976 (N_20976,N_14323,N_13929);
or U20977 (N_20977,N_16313,N_13829);
and U20978 (N_20978,N_18661,N_18422);
xnor U20979 (N_20979,N_14951,N_13337);
or U20980 (N_20980,N_17407,N_14697);
nand U20981 (N_20981,N_18636,N_12720);
or U20982 (N_20982,N_14667,N_12637);
nor U20983 (N_20983,N_13982,N_14704);
nand U20984 (N_20984,N_18703,N_13700);
and U20985 (N_20985,N_17420,N_14867);
xnor U20986 (N_20986,N_17136,N_16486);
or U20987 (N_20987,N_18100,N_16146);
and U20988 (N_20988,N_18203,N_17892);
xor U20989 (N_20989,N_17555,N_12590);
and U20990 (N_20990,N_13146,N_14947);
or U20991 (N_20991,N_13219,N_14096);
nand U20992 (N_20992,N_14934,N_13455);
nor U20993 (N_20993,N_13025,N_18573);
xnor U20994 (N_20994,N_13387,N_15758);
or U20995 (N_20995,N_14244,N_15797);
nor U20996 (N_20996,N_18605,N_12769);
and U20997 (N_20997,N_15633,N_18014);
xnor U20998 (N_20998,N_12703,N_13011);
and U20999 (N_20999,N_15973,N_12684);
nor U21000 (N_21000,N_17715,N_13775);
nand U21001 (N_21001,N_14539,N_15725);
or U21002 (N_21002,N_14836,N_14792);
nor U21003 (N_21003,N_18295,N_12902);
and U21004 (N_21004,N_14700,N_16248);
nor U21005 (N_21005,N_16069,N_17735);
nor U21006 (N_21006,N_14565,N_14584);
and U21007 (N_21007,N_16304,N_14303);
nand U21008 (N_21008,N_15716,N_15238);
or U21009 (N_21009,N_18423,N_15583);
or U21010 (N_21010,N_17091,N_14825);
xor U21011 (N_21011,N_18544,N_17671);
nand U21012 (N_21012,N_17345,N_14971);
or U21013 (N_21013,N_17478,N_16771);
xor U21014 (N_21014,N_16298,N_15080);
nor U21015 (N_21015,N_14893,N_14741);
nor U21016 (N_21016,N_18205,N_14686);
and U21017 (N_21017,N_12609,N_18051);
and U21018 (N_21018,N_14822,N_16626);
or U21019 (N_21019,N_13763,N_14756);
and U21020 (N_21020,N_17181,N_15630);
or U21021 (N_21021,N_15323,N_18009);
nand U21022 (N_21022,N_15926,N_14732);
nand U21023 (N_21023,N_16560,N_13547);
nor U21024 (N_21024,N_18517,N_15781);
nand U21025 (N_21025,N_14829,N_18654);
and U21026 (N_21026,N_16515,N_13780);
nand U21027 (N_21027,N_12676,N_14739);
and U21028 (N_21028,N_14635,N_17452);
or U21029 (N_21029,N_14280,N_13253);
and U21030 (N_21030,N_13321,N_13861);
or U21031 (N_21031,N_13350,N_12934);
and U21032 (N_21032,N_16948,N_15860);
and U21033 (N_21033,N_18318,N_13715);
and U21034 (N_21034,N_12658,N_17751);
nand U21035 (N_21035,N_17687,N_12805);
nand U21036 (N_21036,N_13101,N_16716);
or U21037 (N_21037,N_18274,N_16830);
and U21038 (N_21038,N_15220,N_16880);
nor U21039 (N_21039,N_17802,N_15453);
or U21040 (N_21040,N_14420,N_17016);
or U21041 (N_21041,N_16748,N_15015);
xor U21042 (N_21042,N_13168,N_14025);
nor U21043 (N_21043,N_17386,N_14321);
nand U21044 (N_21044,N_16227,N_16930);
xor U21045 (N_21045,N_17251,N_18487);
xor U21046 (N_21046,N_17308,N_17777);
nand U21047 (N_21047,N_16276,N_14454);
or U21048 (N_21048,N_15793,N_13633);
xnor U21049 (N_21049,N_17565,N_18481);
nand U21050 (N_21050,N_15107,N_13483);
and U21051 (N_21051,N_13512,N_14781);
nor U21052 (N_21052,N_15494,N_15813);
nor U21053 (N_21053,N_12987,N_12850);
or U21054 (N_21054,N_14091,N_14150);
and U21055 (N_21055,N_15832,N_14753);
nor U21056 (N_21056,N_14145,N_18419);
nand U21057 (N_21057,N_15257,N_17996);
nand U21058 (N_21058,N_12756,N_13180);
xor U21059 (N_21059,N_14657,N_17470);
or U21060 (N_21060,N_14794,N_17652);
or U21061 (N_21061,N_16375,N_13601);
nand U21062 (N_21062,N_16234,N_12795);
nor U21063 (N_21063,N_12919,N_18509);
or U21064 (N_21064,N_13631,N_14169);
nand U21065 (N_21065,N_14206,N_17086);
nor U21066 (N_21066,N_14171,N_13034);
nor U21067 (N_21067,N_14600,N_18118);
or U21068 (N_21068,N_17929,N_16050);
xor U21069 (N_21069,N_18539,N_12701);
nor U21070 (N_21070,N_14060,N_12918);
nand U21071 (N_21071,N_14766,N_17337);
and U21072 (N_21072,N_17638,N_16195);
or U21073 (N_21073,N_14502,N_14460);
and U21074 (N_21074,N_12664,N_18494);
nor U21075 (N_21075,N_14226,N_18200);
or U21076 (N_21076,N_17019,N_17068);
nor U21077 (N_21077,N_16044,N_14004);
nor U21078 (N_21078,N_15383,N_18056);
xor U21079 (N_21079,N_18520,N_15527);
and U21080 (N_21080,N_14515,N_12682);
xor U21081 (N_21081,N_13223,N_15473);
nor U21082 (N_21082,N_17018,N_13826);
nor U21083 (N_21083,N_18147,N_14790);
or U21084 (N_21084,N_17609,N_18468);
and U21085 (N_21085,N_15193,N_12697);
or U21086 (N_21086,N_16340,N_13756);
and U21087 (N_21087,N_13472,N_15536);
nand U21088 (N_21088,N_16390,N_17000);
nand U21089 (N_21089,N_16358,N_15228);
or U21090 (N_21090,N_18223,N_12840);
nor U21091 (N_21091,N_14352,N_14748);
nor U21092 (N_21092,N_12598,N_17958);
nand U21093 (N_21093,N_15049,N_18707);
nand U21094 (N_21094,N_17998,N_13754);
or U21095 (N_21095,N_18041,N_16559);
and U21096 (N_21096,N_17635,N_16885);
nand U21097 (N_21097,N_16671,N_15267);
nand U21098 (N_21098,N_14802,N_16152);
nand U21099 (N_21099,N_15426,N_14975);
nor U21100 (N_21100,N_12542,N_12508);
and U21101 (N_21101,N_14090,N_15848);
or U21102 (N_21102,N_15170,N_16424);
xnor U21103 (N_21103,N_15490,N_16912);
and U21104 (N_21104,N_13856,N_13134);
nor U21105 (N_21105,N_18437,N_12932);
xor U21106 (N_21106,N_16394,N_13986);
nand U21107 (N_21107,N_12877,N_12801);
nand U21108 (N_21108,N_14672,N_16801);
xnor U21109 (N_21109,N_13553,N_17280);
or U21110 (N_21110,N_18590,N_16359);
xnor U21111 (N_21111,N_15452,N_17363);
and U21112 (N_21112,N_16628,N_18156);
or U21113 (N_21113,N_13460,N_18175);
nor U21114 (N_21114,N_12671,N_17325);
and U21115 (N_21115,N_15691,N_15934);
and U21116 (N_21116,N_15062,N_17541);
or U21117 (N_21117,N_17845,N_18587);
nand U21118 (N_21118,N_12540,N_16541);
and U21119 (N_21119,N_13574,N_15117);
or U21120 (N_21120,N_16231,N_13243);
xor U21121 (N_21121,N_16910,N_17650);
nand U21122 (N_21122,N_13426,N_13571);
nand U21123 (N_21123,N_15134,N_12911);
and U21124 (N_21124,N_15468,N_18171);
or U21125 (N_21125,N_14933,N_16071);
nor U21126 (N_21126,N_14437,N_14519);
or U21127 (N_21127,N_15741,N_13403);
xor U21128 (N_21128,N_15597,N_12959);
nor U21129 (N_21129,N_15496,N_13508);
nand U21130 (N_21130,N_18612,N_14475);
nand U21131 (N_21131,N_14834,N_13640);
and U21132 (N_21132,N_13276,N_14560);
or U21133 (N_21133,N_16405,N_18637);
nor U21134 (N_21134,N_17903,N_15584);
and U21135 (N_21135,N_13201,N_15478);
and U21136 (N_21136,N_14341,N_18413);
nand U21137 (N_21137,N_13344,N_16695);
xor U21138 (N_21138,N_18734,N_16705);
nor U21139 (N_21139,N_18689,N_18404);
and U21140 (N_21140,N_12999,N_16437);
nor U21141 (N_21141,N_16664,N_16982);
nand U21142 (N_21142,N_17599,N_14412);
nand U21143 (N_21143,N_13997,N_15529);
nand U21144 (N_21144,N_14353,N_15811);
and U21145 (N_21145,N_16188,N_15146);
nand U21146 (N_21146,N_15019,N_13393);
or U21147 (N_21147,N_18737,N_18660);
nor U21148 (N_21148,N_14589,N_14913);
or U21149 (N_21149,N_16354,N_12789);
or U21150 (N_21150,N_14581,N_16595);
nand U21151 (N_21151,N_14008,N_14961);
or U21152 (N_21152,N_16614,N_15649);
and U21153 (N_21153,N_14510,N_16882);
nor U21154 (N_21154,N_18551,N_15852);
and U21155 (N_21155,N_12613,N_14571);
or U21156 (N_21156,N_16736,N_13975);
nand U21157 (N_21157,N_18376,N_13871);
or U21158 (N_21158,N_15421,N_16745);
and U21159 (N_21159,N_13159,N_15384);
or U21160 (N_21160,N_15523,N_14326);
and U21161 (N_21161,N_14764,N_16147);
nand U21162 (N_21162,N_16786,N_15571);
nand U21163 (N_21163,N_18698,N_13375);
nand U21164 (N_21164,N_13060,N_16791);
or U21165 (N_21165,N_18188,N_17391);
nor U21166 (N_21166,N_17619,N_13046);
and U21167 (N_21167,N_16489,N_17434);
nand U21168 (N_21168,N_13507,N_16336);
nand U21169 (N_21169,N_18068,N_12750);
nand U21170 (N_21170,N_12673,N_14784);
or U21171 (N_21171,N_18398,N_15506);
nand U21172 (N_21172,N_13194,N_14890);
nor U21173 (N_21173,N_15415,N_16258);
or U21174 (N_21174,N_18488,N_17961);
nand U21175 (N_21175,N_16209,N_13420);
xnor U21176 (N_21176,N_16703,N_18229);
nand U21177 (N_21177,N_17250,N_17150);
and U21178 (N_21178,N_16827,N_12799);
nor U21179 (N_21179,N_15821,N_18496);
and U21180 (N_21180,N_17622,N_17962);
or U21181 (N_21181,N_15327,N_16593);
nand U21182 (N_21182,N_15026,N_12925);
nand U21183 (N_21183,N_16346,N_16149);
nand U21184 (N_21184,N_14877,N_16396);
and U21185 (N_21185,N_14077,N_17881);
or U21186 (N_21186,N_13707,N_13559);
or U21187 (N_21187,N_18061,N_18369);
nand U21188 (N_21188,N_13315,N_17882);
nand U21189 (N_21189,N_17863,N_12865);
and U21190 (N_21190,N_17930,N_13593);
nand U21191 (N_21191,N_16387,N_17176);
nand U21192 (N_21192,N_17935,N_17971);
and U21193 (N_21193,N_14578,N_15977);
and U21194 (N_21194,N_14045,N_14940);
or U21195 (N_21195,N_14555,N_14234);
nor U21196 (N_21196,N_14545,N_17498);
xnor U21197 (N_21197,N_14738,N_14993);
nand U21198 (N_21198,N_18184,N_13430);
xnor U21199 (N_21199,N_14426,N_16654);
nor U21200 (N_21200,N_12731,N_13506);
or U21201 (N_21201,N_14466,N_13746);
and U21202 (N_21202,N_13740,N_15373);
nor U21203 (N_21203,N_18115,N_13138);
or U21204 (N_21204,N_17708,N_18581);
nor U21205 (N_21205,N_14097,N_17448);
nor U21206 (N_21206,N_15413,N_14463);
xnor U21207 (N_21207,N_14920,N_18162);
or U21208 (N_21208,N_16376,N_17778);
xnor U21209 (N_21209,N_15959,N_18410);
and U21210 (N_21210,N_16970,N_13765);
and U21211 (N_21211,N_15161,N_17433);
and U21212 (N_21212,N_16388,N_18549);
nor U21213 (N_21213,N_12776,N_15157);
and U21214 (N_21214,N_16369,N_15752);
and U21215 (N_21215,N_17107,N_17129);
and U21216 (N_21216,N_13932,N_13855);
or U21217 (N_21217,N_17640,N_17771);
and U21218 (N_21218,N_15953,N_16877);
and U21219 (N_21219,N_16329,N_18154);
nand U21220 (N_21220,N_18095,N_15788);
nand U21221 (N_21221,N_16413,N_14614);
or U21222 (N_21222,N_14827,N_16754);
or U21223 (N_21223,N_15135,N_14379);
nand U21224 (N_21224,N_12537,N_17504);
or U21225 (N_21225,N_16550,N_17551);
nor U21226 (N_21226,N_17228,N_14316);
nand U21227 (N_21227,N_17907,N_12782);
nand U21228 (N_21228,N_13354,N_18108);
nor U21229 (N_21229,N_17556,N_15960);
nand U21230 (N_21230,N_16932,N_17902);
nor U21231 (N_21231,N_17659,N_17569);
nand U21232 (N_21232,N_12998,N_13003);
nor U21233 (N_21233,N_15624,N_16579);
nand U21234 (N_21234,N_15179,N_18646);
or U21235 (N_21235,N_18262,N_18032);
nor U21236 (N_21236,N_15351,N_15340);
xnor U21237 (N_21237,N_14726,N_15854);
nor U21238 (N_21238,N_17500,N_15308);
or U21239 (N_21239,N_15518,N_17104);
and U21240 (N_21240,N_15802,N_17791);
nand U21241 (N_21241,N_13985,N_17637);
and U21242 (N_21242,N_13570,N_16974);
or U21243 (N_21243,N_13071,N_13848);
or U21244 (N_21244,N_13108,N_16156);
or U21245 (N_21245,N_15463,N_17153);
nand U21246 (N_21246,N_16492,N_15944);
and U21247 (N_21247,N_15989,N_16009);
or U21248 (N_21248,N_17418,N_13322);
nand U21249 (N_21249,N_18104,N_13644);
and U21250 (N_21250,N_13351,N_13966);
or U21251 (N_21251,N_16264,N_18550);
and U21252 (N_21252,N_14906,N_15791);
nand U21253 (N_21253,N_12735,N_16096);
nand U21254 (N_21254,N_15744,N_14888);
nand U21255 (N_21255,N_17890,N_15378);
nor U21256 (N_21256,N_18176,N_17117);
nor U21257 (N_21257,N_13535,N_17584);
and U21258 (N_21258,N_16047,N_15592);
nor U21259 (N_21259,N_15690,N_16949);
nor U21260 (N_21260,N_15616,N_15434);
nor U21261 (N_21261,N_18484,N_17154);
or U21262 (N_21262,N_17261,N_13611);
nand U21263 (N_21263,N_12986,N_17122);
nor U21264 (N_21264,N_16249,N_13797);
and U21265 (N_21265,N_17533,N_17760);
and U21266 (N_21266,N_17629,N_14644);
nor U21267 (N_21267,N_15949,N_13969);
xnor U21268 (N_21268,N_15391,N_12957);
or U21269 (N_21269,N_17485,N_18182);
or U21270 (N_21270,N_16637,N_15150);
or U21271 (N_21271,N_14842,N_15263);
and U21272 (N_21272,N_13038,N_13336);
and U21273 (N_21273,N_17518,N_12677);
and U21274 (N_21274,N_14388,N_18352);
nor U21275 (N_21275,N_16175,N_15873);
or U21276 (N_21276,N_13292,N_14197);
and U21277 (N_21277,N_14880,N_18196);
nand U21278 (N_21278,N_13728,N_15095);
or U21279 (N_21279,N_15540,N_14977);
and U21280 (N_21280,N_12718,N_16162);
or U21281 (N_21281,N_14785,N_17678);
and U21282 (N_21282,N_17948,N_15835);
nor U21283 (N_21283,N_17879,N_12626);
or U21284 (N_21284,N_17013,N_18566);
and U21285 (N_21285,N_12602,N_14295);
xnor U21286 (N_21286,N_17100,N_13293);
or U21287 (N_21287,N_15256,N_15975);
nand U21288 (N_21288,N_13014,N_17593);
xnor U21289 (N_21289,N_18730,N_16133);
xor U21290 (N_21290,N_14689,N_17782);
nor U21291 (N_21291,N_14122,N_17835);
or U21292 (N_21292,N_17734,N_15872);
nor U21293 (N_21293,N_15446,N_17173);
or U21294 (N_21294,N_15558,N_18013);
nand U21295 (N_21295,N_14665,N_17057);
or U21296 (N_21296,N_12710,N_18638);
nor U21297 (N_21297,N_13811,N_15777);
and U21298 (N_21298,N_15035,N_12592);
nor U21299 (N_21299,N_14844,N_16905);
xor U21300 (N_21300,N_17924,N_15586);
nand U21301 (N_21301,N_17561,N_13205);
or U21302 (N_21302,N_18466,N_16670);
nor U21303 (N_21303,N_15289,N_17977);
and U21304 (N_21304,N_15052,N_14416);
nand U21305 (N_21305,N_18535,N_16110);
nor U21306 (N_21306,N_15553,N_16937);
or U21307 (N_21307,N_14912,N_14029);
and U21308 (N_21308,N_15108,N_16607);
and U21309 (N_21309,N_12817,N_17252);
and U21310 (N_21310,N_15054,N_17955);
and U21311 (N_21311,N_16774,N_15534);
or U21312 (N_21312,N_13381,N_15501);
xor U21313 (N_21313,N_14386,N_16726);
nand U21314 (N_21314,N_13583,N_16062);
or U21315 (N_21315,N_15555,N_14098);
xnor U21316 (N_21316,N_12716,N_16629);
and U21317 (N_21317,N_16075,N_17241);
and U21318 (N_21318,N_17909,N_16985);
xor U21319 (N_21319,N_12941,N_17532);
nand U21320 (N_21320,N_13706,N_16887);
and U21321 (N_21321,N_18471,N_15115);
nand U21322 (N_21322,N_12881,N_14734);
xor U21323 (N_21323,N_14992,N_16428);
nand U21324 (N_21324,N_13719,N_16059);
xnor U21325 (N_21325,N_13863,N_13899);
nand U21326 (N_21326,N_18424,N_14789);
and U21327 (N_21327,N_15460,N_14369);
and U21328 (N_21328,N_15663,N_16984);
xor U21329 (N_21329,N_13664,N_14782);
nand U21330 (N_21330,N_14769,N_12528);
nor U21331 (N_21331,N_14548,N_15998);
and U21332 (N_21332,N_15617,N_13582);
nand U21333 (N_21333,N_12923,N_12824);
and U21334 (N_21334,N_18117,N_15266);
and U21335 (N_21335,N_18054,N_14448);
or U21336 (N_21336,N_15187,N_16315);
or U21337 (N_21337,N_17352,N_14911);
nor U21338 (N_21338,N_12516,N_16404);
and U21339 (N_21339,N_14349,N_14709);
or U21340 (N_21340,N_13581,N_13405);
and U21341 (N_21341,N_18681,N_13643);
and U21342 (N_21342,N_17517,N_13949);
and U21343 (N_21343,N_14595,N_15325);
nand U21344 (N_21344,N_12889,N_17811);
nor U21345 (N_21345,N_14231,N_18042);
or U21346 (N_21346,N_14895,N_16443);
nor U21347 (N_21347,N_12851,N_13443);
and U21348 (N_21348,N_16480,N_18630);
nand U21349 (N_21349,N_18046,N_16129);
nor U21350 (N_21350,N_15129,N_15010);
and U21351 (N_21351,N_16328,N_16682);
nand U21352 (N_21352,N_14703,N_18700);
nor U21353 (N_21353,N_15674,N_18220);
and U21354 (N_21354,N_15041,N_16638);
and U21355 (N_21355,N_18478,N_15261);
nor U21356 (N_21356,N_15202,N_12992);
or U21357 (N_21357,N_16039,N_15480);
or U21358 (N_21358,N_13843,N_13846);
and U21359 (N_21359,N_16876,N_15987);
nand U21360 (N_21360,N_12954,N_16244);
or U21361 (N_21361,N_17922,N_15078);
and U21362 (N_21362,N_16699,N_15275);
or U21363 (N_21363,N_13928,N_13255);
and U21364 (N_21364,N_18537,N_12815);
nor U21365 (N_21365,N_13995,N_17006);
or U21366 (N_21366,N_14396,N_13935);
nand U21367 (N_21367,N_16964,N_16504);
nand U21368 (N_21368,N_17215,N_14478);
and U21369 (N_21369,N_18092,N_14360);
nor U21370 (N_21370,N_18327,N_15102);
xor U21371 (N_21371,N_14330,N_15328);
xnor U21372 (N_21372,N_15818,N_17314);
or U21373 (N_21373,N_15885,N_12759);
and U21374 (N_21374,N_18005,N_17613);
nor U21375 (N_21375,N_13251,N_15632);
and U21376 (N_21376,N_17677,N_16980);
nor U21377 (N_21377,N_15510,N_14549);
and U21378 (N_21378,N_15650,N_14103);
or U21379 (N_21379,N_13533,N_12948);
xnor U21380 (N_21380,N_15109,N_17427);
and U21381 (N_21381,N_13423,N_14553);
xor U21382 (N_21382,N_12738,N_14886);
nor U21383 (N_21383,N_12758,N_13621);
nand U21384 (N_21384,N_15946,N_17402);
nor U21385 (N_21385,N_17932,N_13486);
and U21386 (N_21386,N_15309,N_13569);
and U21387 (N_21387,N_13428,N_13496);
nor U21388 (N_21388,N_14086,N_17746);
xor U21389 (N_21389,N_17667,N_15940);
xnor U21390 (N_21390,N_14200,N_12532);
and U21391 (N_21391,N_16079,N_18047);
nand U21392 (N_21392,N_12663,N_16643);
and U21393 (N_21393,N_13424,N_18640);
or U21394 (N_21394,N_12784,N_16447);
nor U21395 (N_21395,N_13799,N_18447);
nand U21396 (N_21396,N_16217,N_16501);
and U21397 (N_21397,N_14943,N_16888);
or U21398 (N_21398,N_17669,N_15593);
xor U21399 (N_21399,N_16605,N_13261);
or U21400 (N_21400,N_15648,N_15431);
or U21401 (N_21401,N_15817,N_18291);
and U21402 (N_21402,N_16201,N_14708);
nand U21403 (N_21403,N_14561,N_18613);
nand U21404 (N_21404,N_16005,N_12550);
nand U21405 (N_21405,N_15682,N_16157);
nor U21406 (N_21406,N_15670,N_18672);
nand U21407 (N_21407,N_15185,N_16502);
nor U21408 (N_21408,N_18053,N_14622);
and U21409 (N_21409,N_13892,N_18485);
nand U21410 (N_21410,N_14493,N_14640);
xnor U21411 (N_21411,N_15396,N_17511);
nand U21412 (N_21412,N_12675,N_18304);
nand U21413 (N_21413,N_12831,N_13973);
nor U21414 (N_21414,N_18366,N_13658);
nand U21415 (N_21415,N_16997,N_16511);
nor U21416 (N_21416,N_15880,N_14267);
or U21417 (N_21417,N_14385,N_17804);
and U21418 (N_21418,N_15660,N_18234);
or U21419 (N_21419,N_12927,N_15700);
nand U21420 (N_21420,N_12890,N_14596);
or U21421 (N_21421,N_17796,N_17539);
and U21422 (N_21422,N_16823,N_16035);
and U21423 (N_21423,N_15993,N_12774);
xnor U21424 (N_21424,N_12891,N_17123);
xnor U21425 (N_21425,N_15521,N_13845);
or U21426 (N_21426,N_13280,N_18084);
and U21427 (N_21427,N_17904,N_14484);
nand U21428 (N_21428,N_17220,N_17423);
and U21429 (N_21429,N_18199,N_17194);
or U21430 (N_21430,N_17118,N_14669);
nand U21431 (N_21431,N_12870,N_17692);
nand U21432 (N_21432,N_14344,N_16749);
or U21433 (N_21433,N_13967,N_15083);
or U21434 (N_21434,N_18695,N_18465);
or U21435 (N_21435,N_14768,N_15465);
nand U21436 (N_21436,N_15958,N_17770);
xnor U21437 (N_21437,N_16155,N_17630);
and U21438 (N_21438,N_16571,N_13517);
nand U21439 (N_21439,N_13714,N_14119);
nor U21440 (N_21440,N_14042,N_13416);
xnor U21441 (N_21441,N_13441,N_14327);
nor U21442 (N_21442,N_17837,N_18473);
or U21443 (N_21443,N_16457,N_15983);
nor U21444 (N_21444,N_14260,N_13481);
xnor U21445 (N_21445,N_18709,N_15703);
or U21446 (N_21446,N_17193,N_17254);
nand U21447 (N_21447,N_18540,N_18296);
nand U21448 (N_21448,N_14942,N_14413);
and U21449 (N_21449,N_16516,N_16738);
and U21450 (N_21450,N_15874,N_15037);
or U21451 (N_21451,N_14408,N_14793);
and U21452 (N_21452,N_18347,N_17208);
and U21453 (N_21453,N_13964,N_14152);
nand U21454 (N_21454,N_14348,N_13556);
or U21455 (N_21455,N_14673,N_16245);
xnor U21456 (N_21456,N_16693,N_14687);
and U21457 (N_21457,N_18430,N_15827);
nor U21458 (N_21458,N_13827,N_16779);
and U21459 (N_21459,N_16049,N_16030);
nand U21460 (N_21460,N_13063,N_15225);
nor U21461 (N_21461,N_16601,N_18247);
and U21462 (N_21462,N_13482,N_16224);
or U21463 (N_21463,N_14945,N_14892);
nor U21464 (N_21464,N_18195,N_17797);
and U21465 (N_21465,N_18514,N_13147);
xor U21466 (N_21466,N_13683,N_13676);
xnor U21467 (N_21467,N_15560,N_13654);
nand U21468 (N_21468,N_16381,N_17926);
and U21469 (N_21469,N_16259,N_14458);
xnor U21470 (N_21470,N_12525,N_15883);
and U21471 (N_21471,N_14238,N_14422);
and U21472 (N_21472,N_18663,N_13090);
nand U21473 (N_21473,N_12808,N_15027);
nand U21474 (N_21474,N_17972,N_18723);
nand U21475 (N_21475,N_14314,N_14485);
nand U21476 (N_21476,N_17165,N_13296);
or U21477 (N_21477,N_18586,N_18559);
and U21478 (N_21478,N_18071,N_14588);
nand U21479 (N_21479,N_17544,N_18738);
or U21480 (N_21480,N_12518,N_14133);
nor U21481 (N_21481,N_15784,N_12596);
or U21482 (N_21482,N_17092,N_12549);
nand U21483 (N_21483,N_14136,N_16403);
nor U21484 (N_21484,N_14610,N_16539);
nor U21485 (N_21485,N_14124,N_17945);
nor U21486 (N_21486,N_15665,N_16187);
nand U21487 (N_21487,N_12503,N_14691);
or U21488 (N_21488,N_17853,N_13466);
or U21489 (N_21489,N_14924,N_14777);
nand U21490 (N_21490,N_17001,N_13027);
nor U21491 (N_21491,N_16275,N_18253);
nand U21492 (N_21492,N_18334,N_15576);
nand U21493 (N_21493,N_13346,N_16427);
or U21494 (N_21494,N_16837,N_14187);
nor U21495 (N_21495,N_18628,N_18153);
nor U21496 (N_21496,N_14085,N_17225);
nand U21497 (N_21497,N_18402,N_15357);
and U21498 (N_21498,N_14013,N_13458);
and U21499 (N_21499,N_14028,N_14093);
nor U21500 (N_21500,N_16685,N_12899);
and U21501 (N_21501,N_13911,N_14177);
and U21502 (N_21502,N_13408,N_16228);
nand U21503 (N_21503,N_16161,N_16280);
nand U21504 (N_21504,N_14481,N_15768);
and U21505 (N_21505,N_13518,N_13696);
and U21506 (N_21506,N_17897,N_13242);
xnor U21507 (N_21507,N_13806,N_15464);
and U21508 (N_21508,N_17774,N_18574);
and U21509 (N_21509,N_13823,N_13962);
or U21510 (N_21510,N_15152,N_12839);
nand U21511 (N_21511,N_13160,N_14823);
nor U21512 (N_21512,N_12541,N_17022);
nand U21513 (N_21513,N_14378,N_17120);
xnor U21514 (N_21514,N_15399,N_18206);
and U21515 (N_21515,N_14052,N_15986);
nand U21516 (N_21516,N_15477,N_14526);
nand U21517 (N_21517,N_14202,N_18391);
and U21518 (N_21518,N_17119,N_14952);
or U21519 (N_21519,N_18445,N_16450);
nor U21520 (N_21520,N_17744,N_13889);
nor U21521 (N_21521,N_15939,N_12725);
xnor U21522 (N_21522,N_13833,N_12605);
nor U21523 (N_21523,N_18037,N_17505);
nor U21524 (N_21524,N_17768,N_17789);
xor U21525 (N_21525,N_15450,N_16901);
nor U21526 (N_21526,N_17607,N_16546);
or U21527 (N_21527,N_16434,N_16781);
nor U21528 (N_21528,N_16225,N_13230);
and U21529 (N_21529,N_15474,N_17957);
xor U21530 (N_21530,N_14767,N_16721);
nand U21531 (N_21531,N_18209,N_12713);
nand U21532 (N_21532,N_18307,N_16636);
nand U21533 (N_21533,N_18435,N_18329);
and U21534 (N_21534,N_15335,N_14962);
nand U21535 (N_21535,N_15922,N_17075);
and U21536 (N_21536,N_18198,N_18105);
nor U21537 (N_21537,N_14490,N_14232);
xnor U21538 (N_21538,N_15812,N_18526);
or U21539 (N_21539,N_13901,N_17547);
xor U21540 (N_21540,N_17710,N_14616);
nand U21541 (N_21541,N_14162,N_13365);
or U21542 (N_21542,N_14078,N_18125);
and U21543 (N_21543,N_14887,N_14031);
or U21544 (N_21544,N_15561,N_16014);
nor U21545 (N_21545,N_13247,N_15830);
xor U21546 (N_21546,N_14116,N_13980);
nor U21547 (N_21547,N_12568,N_18673);
nor U21548 (N_21548,N_14559,N_18043);
nand U21549 (N_21549,N_18346,N_17603);
nor U21550 (N_21550,N_13505,N_13361);
nor U21551 (N_21551,N_13213,N_16214);
and U21552 (N_21552,N_13069,N_16254);
nor U21553 (N_21553,N_14542,N_18122);
nor U21554 (N_21554,N_13197,N_16158);
or U21555 (N_21555,N_17361,N_12763);
nor U21556 (N_21556,N_16382,N_16521);
nor U21557 (N_21557,N_16407,N_15331);
and U21558 (N_21558,N_16032,N_17223);
and U21559 (N_21559,N_14731,N_17726);
nand U21560 (N_21560,N_12709,N_12811);
nor U21561 (N_21561,N_16641,N_12760);
nor U21562 (N_21562,N_16243,N_14811);
nor U21563 (N_21563,N_15851,N_13469);
or U21564 (N_21564,N_15846,N_16862);
and U21565 (N_21565,N_14765,N_14071);
nand U21566 (N_21566,N_16293,N_17548);
nor U21567 (N_21567,N_16454,N_12552);
nor U21568 (N_21568,N_17340,N_15641);
xor U21569 (N_21569,N_17011,N_17702);
xor U21570 (N_21570,N_14125,N_16160);
nor U21571 (N_21571,N_18746,N_15024);
nor U21572 (N_21572,N_16755,N_15732);
nor U21573 (N_21573,N_15132,N_14838);
nand U21574 (N_21574,N_17844,N_17492);
or U21575 (N_21575,N_13688,N_12599);
and U21576 (N_21576,N_13362,N_16260);
or U21577 (N_21577,N_17293,N_13862);
nand U21578 (N_21578,N_16956,N_14146);
and U21579 (N_21579,N_14033,N_16290);
or U21580 (N_21580,N_16815,N_17481);
nand U21581 (N_21581,N_15352,N_17369);
nor U21582 (N_21582,N_14275,N_15704);
nor U21583 (N_21583,N_13992,N_16301);
nor U21584 (N_21584,N_12949,N_14503);
xnor U21585 (N_21585,N_12904,N_14585);
and U21586 (N_21586,N_15921,N_18597);
xor U21587 (N_21587,N_18370,N_15429);
nor U21588 (N_21588,N_16127,N_16312);
nor U21589 (N_21589,N_16812,N_16461);
nor U21590 (N_21590,N_18617,N_17103);
or U21591 (N_21591,N_14636,N_15776);
nand U21592 (N_21592,N_15349,N_13792);
nand U21593 (N_21593,N_14905,N_16939);
nand U21594 (N_21594,N_16445,N_17920);
and U21595 (N_21595,N_17523,N_12836);
or U21596 (N_21596,N_18733,N_16859);
and U21597 (N_21597,N_15747,N_16138);
nor U21598 (N_21598,N_16255,N_12519);
nor U21599 (N_21599,N_16210,N_16020);
and U21600 (N_21600,N_18578,N_13834);
and U21601 (N_21601,N_13592,N_16718);
and U21602 (N_21602,N_13653,N_12929);
or U21603 (N_21603,N_12761,N_18172);
and U21604 (N_21604,N_18438,N_16590);
nand U21605 (N_21605,N_17077,N_17676);
or U21606 (N_21606,N_13137,N_15353);
nor U21607 (N_21607,N_13509,N_18174);
or U21608 (N_21608,N_13614,N_16154);
nor U21609 (N_21609,N_16308,N_14534);
nand U21610 (N_21610,N_16159,N_15594);
nor U21611 (N_21611,N_14533,N_13606);
and U21612 (N_21612,N_18444,N_16803);
nand U21613 (N_21613,N_17657,N_15706);
or U21614 (N_21614,N_14361,N_18216);
and U21615 (N_21615,N_17147,N_14089);
nor U21616 (N_21616,N_15040,N_13503);
and U21617 (N_21617,N_17813,N_17116);
nor U21618 (N_21618,N_18567,N_17756);
and U21619 (N_21619,N_16684,N_17895);
xor U21620 (N_21620,N_14172,N_16995);
or U21621 (N_21621,N_13622,N_15183);
or U21622 (N_21622,N_15241,N_17912);
nand U21623 (N_21623,N_16981,N_13585);
and U21624 (N_21624,N_17601,N_13012);
nand U21625 (N_21625,N_18275,N_14447);
nor U21626 (N_21626,N_16176,N_15991);
and U21627 (N_21627,N_16191,N_13623);
nand U21628 (N_21628,N_15829,N_13449);
nand U21629 (N_21629,N_13551,N_14680);
xor U21630 (N_21630,N_14925,N_17312);
or U21631 (N_21631,N_15551,N_17299);
and U21632 (N_21632,N_13541,N_14112);
nor U21633 (N_21633,N_16041,N_15074);
or U21634 (N_21634,N_12740,N_16782);
xor U21635 (N_21635,N_17316,N_17799);
xnor U21636 (N_21636,N_14134,N_14761);
and U21637 (N_21637,N_13444,N_16508);
and U21638 (N_21638,N_13808,N_13960);
or U21639 (N_21639,N_13920,N_17506);
nor U21640 (N_21640,N_17138,N_13317);
nand U21641 (N_21641,N_17089,N_18003);
or U21642 (N_21642,N_17611,N_16420);
nand U21643 (N_21643,N_15580,N_18324);
or U21644 (N_21644,N_15595,N_17953);
xor U21645 (N_21645,N_14517,N_12940);
and U21646 (N_21646,N_15900,N_16594);
nor U21647 (N_21647,N_16979,N_15750);
nor U21648 (N_21648,N_14179,N_15128);
or U21649 (N_21649,N_14011,N_15844);
and U21650 (N_21650,N_16498,N_13141);
or U21651 (N_21651,N_17344,N_17839);
nand U21652 (N_21652,N_17642,N_14070);
nand U21653 (N_21653,N_15484,N_14227);
or U21654 (N_21654,N_14250,N_13422);
and U21655 (N_21655,N_15033,N_16658);
or U21656 (N_21656,N_17720,N_15807);
and U21657 (N_21657,N_14218,N_14300);
and U21658 (N_21658,N_17833,N_17834);
or U21659 (N_21659,N_14711,N_13697);
or U21660 (N_21660,N_18633,N_17496);
nor U21661 (N_21661,N_18664,N_16916);
xor U21662 (N_21662,N_14304,N_16724);
nor U21663 (N_21663,N_15197,N_16811);
nor U21664 (N_21664,N_13039,N_18142);
and U21665 (N_21665,N_18266,N_15757);
nand U21666 (N_21666,N_17816,N_15243);
and U21667 (N_21667,N_18246,N_14508);
xor U21668 (N_21668,N_14015,N_14296);
or U21669 (N_21669,N_18353,N_17780);
or U21670 (N_21670,N_17785,N_13111);
and U21671 (N_21671,N_14863,N_13051);
xor U21672 (N_21672,N_16478,N_18159);
nand U21673 (N_21673,N_12570,N_12511);
and U21674 (N_21674,N_12823,N_13305);
or U21675 (N_21675,N_17665,N_12837);
xnor U21676 (N_21676,N_15344,N_15264);
xor U21677 (N_21677,N_17320,N_16692);
nor U21678 (N_21678,N_16908,N_15749);
nand U21679 (N_21679,N_15472,N_17880);
nor U21680 (N_21680,N_14573,N_16923);
and U21681 (N_21681,N_15398,N_15479);
nor U21682 (N_21682,N_14252,N_18667);
nand U21683 (N_21683,N_16141,N_13854);
and U21684 (N_21684,N_15720,N_14720);
and U21685 (N_21685,N_13312,N_17445);
and U21686 (N_21686,N_13122,N_13340);
nor U21687 (N_21687,N_13107,N_12970);
xnor U21688 (N_21688,N_17290,N_13304);
or U21689 (N_21689,N_14126,N_17968);
xor U21690 (N_21690,N_16099,N_18446);
or U21691 (N_21691,N_16065,N_14921);
nand U21692 (N_21692,N_18331,N_14544);
and U21693 (N_21693,N_18024,N_14374);
nor U21694 (N_21694,N_16630,N_13747);
xnor U21695 (N_21695,N_15622,N_15957);
or U21696 (N_21696,N_16522,N_18312);
nand U21697 (N_21697,N_14926,N_12838);
or U21698 (N_21698,N_14530,N_14178);
nor U21699 (N_21699,N_13358,N_14092);
and U21700 (N_21700,N_17148,N_14389);
xor U21701 (N_21701,N_17615,N_15319);
xnor U21702 (N_21702,N_15779,N_16446);
nand U21703 (N_21703,N_13577,N_17852);
nand U21704 (N_21704,N_13544,N_15209);
nor U21705 (N_21705,N_15163,N_13880);
and U21706 (N_21706,N_17267,N_14375);
nand U21707 (N_21707,N_18626,N_15497);
or U21708 (N_21708,N_15122,N_17995);
xor U21709 (N_21709,N_14153,N_14722);
nand U21710 (N_21710,N_13058,N_18579);
nand U21711 (N_21711,N_13801,N_15636);
and U21712 (N_21712,N_14310,N_15879);
xnor U21713 (N_21713,N_14957,N_12538);
xnor U21714 (N_21714,N_15204,N_13587);
nand U21715 (N_21715,N_17761,N_14828);
nor U21716 (N_21716,N_13584,N_13333);
and U21717 (N_21717,N_17672,N_14431);
nand U21718 (N_21718,N_17177,N_18109);
nand U21719 (N_21719,N_16852,N_16845);
xnor U21720 (N_21720,N_12524,N_16861);
nor U21721 (N_21721,N_15038,N_15104);
or U21722 (N_21722,N_18293,N_16042);
and U21723 (N_21723,N_13072,N_18323);
or U21724 (N_21724,N_15444,N_13367);
nand U21725 (N_21725,N_14198,N_12876);
xnor U21726 (N_21726,N_13229,N_16687);
and U21727 (N_21727,N_12736,N_16871);
nand U21728 (N_21728,N_17762,N_17429);
and U21729 (N_21729,N_13943,N_12885);
and U21730 (N_21730,N_13717,N_13940);
nand U21731 (N_21731,N_15111,N_13384);
nor U21732 (N_21732,N_17291,N_18049);
and U21733 (N_21733,N_17417,N_13657);
nor U21734 (N_21734,N_13342,N_16324);
xor U21735 (N_21735,N_17060,N_16834);
nand U21736 (N_21736,N_12614,N_13971);
nand U21737 (N_21737,N_18276,N_14002);
and U21738 (N_21738,N_15745,N_15223);
nor U21739 (N_21739,N_16426,N_15297);
or U21740 (N_21740,N_16115,N_17975);
nor U21741 (N_21741,N_13751,N_18113);
or U21742 (N_21742,N_18190,N_18436);
and U21743 (N_21743,N_12595,N_16936);
and U21744 (N_21744,N_13216,N_18326);
nor U21745 (N_21745,N_13619,N_13078);
or U21746 (N_21746,N_17137,N_18240);
nand U21747 (N_21747,N_14362,N_14847);
nor U21748 (N_21748,N_14030,N_16531);
nor U21749 (N_21749,N_18233,N_17343);
xnor U21750 (N_21750,N_13170,N_17508);
nand U21751 (N_21751,N_18561,N_14723);
nand U21752 (N_21752,N_13998,N_18507);
and U21753 (N_21753,N_16635,N_13378);
nor U21754 (N_21754,N_14651,N_17918);
or U21755 (N_21755,N_12864,N_14213);
and U21756 (N_21756,N_13485,N_17840);
nand U21757 (N_21757,N_16331,N_16688);
nor U21758 (N_21758,N_14853,N_16230);
and U21759 (N_21759,N_14776,N_13950);
and U21760 (N_21760,N_13348,N_16003);
nor U21761 (N_21761,N_17689,N_14461);
xnor U21762 (N_21762,N_15533,N_18338);
nor U21763 (N_21763,N_13504,N_16656);
and U21764 (N_21764,N_12905,N_14428);
or U21765 (N_21765,N_14848,N_14551);
nand U21766 (N_21766,N_13062,N_16218);
nor U21767 (N_21767,N_18739,N_13206);
nand U21768 (N_21768,N_13202,N_16709);
nand U21769 (N_21769,N_16615,N_17365);
nor U21770 (N_21770,N_12894,N_16196);
and U21771 (N_21771,N_13620,N_13917);
or U21772 (N_21772,N_18179,N_13770);
and U21773 (N_21773,N_17070,N_16374);
nand U21774 (N_21774,N_16613,N_15302);
or U21775 (N_21775,N_17113,N_18299);
nand U21776 (N_21776,N_17794,N_18204);
or U21777 (N_21777,N_12800,N_16583);
or U21778 (N_21778,N_14650,N_14570);
nand U21779 (N_21779,N_13271,N_15945);
nor U21780 (N_21780,N_18183,N_13596);
nor U21781 (N_21781,N_16657,N_18676);
and U21782 (N_21782,N_13320,N_14214);
nand U21783 (N_21783,N_13955,N_17032);
and U21784 (N_21784,N_16843,N_15342);
nor U21785 (N_21785,N_15016,N_13888);
nand U21786 (N_21786,N_17656,N_14676);
nand U21787 (N_21787,N_13850,N_15272);
nand U21788 (N_21788,N_13609,N_16102);
or U21789 (N_21789,N_18442,N_13257);
or U21790 (N_21790,N_16988,N_14807);
or U21791 (N_21791,N_14427,N_18235);
xor U21792 (N_21792,N_16007,N_15961);
nand U21793 (N_21793,N_17277,N_16182);
nand U21794 (N_21794,N_13836,N_16878);
nand U21795 (N_21795,N_14164,N_18244);
nor U21796 (N_21796,N_17415,N_14334);
nor U21797 (N_21797,N_14121,N_17914);
nor U21798 (N_21798,N_12624,N_17457);
nor U21799 (N_21799,N_16257,N_16503);
nor U21800 (N_21800,N_16572,N_13860);
xnor U21801 (N_21801,N_15697,N_15231);
or U21802 (N_21802,N_18614,N_15100);
xnor U21803 (N_21803,N_15224,N_17416);
or U21804 (N_21804,N_13286,N_15363);
nor U21805 (N_21805,N_12686,N_16063);
xor U21806 (N_21806,N_14371,N_12634);
or U21807 (N_21807,N_18302,N_15137);
xnor U21808 (N_21808,N_14101,N_16926);
nor U21809 (N_21809,N_13557,N_12691);
or U21810 (N_21810,N_18515,N_16303);
or U21811 (N_21811,N_13024,N_13909);
nor U21812 (N_21812,N_15178,N_13332);
nor U21813 (N_21813,N_15422,N_15995);
nand U21814 (N_21814,N_13796,N_13781);
and U21815 (N_21815,N_16509,N_16967);
xor U21816 (N_21816,N_15242,N_18243);
xnor U21817 (N_21817,N_18704,N_15000);
nor U21818 (N_21818,N_18641,N_12747);
nor U21819 (N_21819,N_14809,N_14574);
nand U21820 (N_21820,N_13324,N_15657);
and U21821 (N_21821,N_17319,N_16734);
or U21822 (N_21822,N_17712,N_18415);
nand U21823 (N_21823,N_16470,N_17004);
or U21824 (N_21824,N_13753,N_16471);
or U21825 (N_21825,N_17368,N_17146);
nand U21826 (N_21826,N_12566,N_13437);
nand U21827 (N_21827,N_14424,N_18384);
nor U21828 (N_21828,N_18499,N_16128);
nand U21829 (N_21829,N_14064,N_17575);
nor U21830 (N_21830,N_18732,N_18148);
or U21831 (N_21831,N_17663,N_14050);
and U21832 (N_21832,N_12628,N_16808);
xor U21833 (N_21833,N_13528,N_16512);
nand U21834 (N_21834,N_15158,N_14331);
nor U21835 (N_21835,N_17664,N_17884);
nor U21836 (N_21836,N_16356,N_16093);
nand U21837 (N_21837,N_17045,N_18230);
or U21838 (N_21838,N_14538,N_16371);
nor U21839 (N_21839,N_17358,N_16488);
and U21840 (N_21840,N_12796,N_12945);
and U21841 (N_21841,N_14391,N_14513);
nand U21842 (N_21842,N_18048,N_16004);
or U21843 (N_21843,N_13002,N_13914);
or U21844 (N_21844,N_17431,N_18453);
nor U21845 (N_21845,N_15177,N_17396);
or U21846 (N_21846,N_13277,N_18354);
nand U21847 (N_21847,N_14161,N_16743);
xor U21848 (N_21848,N_12846,N_13560);
nand U21849 (N_21849,N_18256,N_17078);
xnor U21850 (N_21850,N_14319,N_13501);
or U21851 (N_21851,N_15637,N_14032);
xor U21852 (N_21852,N_15733,N_15205);
xor U21853 (N_21853,N_14801,N_14095);
or U21854 (N_21854,N_12656,N_16950);
and U21855 (N_21855,N_17274,N_17781);
nand U21856 (N_21856,N_12707,N_13816);
nor U21857 (N_21857,N_14106,N_14662);
or U21858 (N_21858,N_17766,N_18611);
nor U21859 (N_21859,N_17857,N_17339);
nand U21860 (N_21860,N_13209,N_16966);
or U21861 (N_21861,N_14821,N_16300);
or U21862 (N_21862,N_14593,N_12692);
nor U21863 (N_21863,N_15978,N_18212);
nor U21864 (N_21864,N_16074,N_13817);
nand U21865 (N_21865,N_16419,N_14381);
or U21866 (N_21866,N_14746,N_17382);
and U21867 (N_21867,N_16122,N_14698);
and U21868 (N_21868,N_16423,N_15849);
nand U21869 (N_21869,N_13844,N_16164);
nor U21870 (N_21870,N_16609,N_16620);
and U21871 (N_21871,N_17810,N_14138);
and U21872 (N_21872,N_13800,N_12662);
or U21873 (N_21873,N_15196,N_17899);
nor U21874 (N_21874,N_17074,N_14309);
nor U21875 (N_21875,N_17362,N_13958);
or U21876 (N_21876,N_15738,N_17162);
or U21877 (N_21877,N_15314,N_17618);
and U21878 (N_21878,N_15022,N_16268);
xnor U21879 (N_21879,N_13642,N_16990);
and U21880 (N_21880,N_16851,N_15476);
nor U21881 (N_21881,N_14764,N_18649);
or U21882 (N_21882,N_15797,N_12806);
nand U21883 (N_21883,N_15586,N_18238);
nand U21884 (N_21884,N_15917,N_12954);
nor U21885 (N_21885,N_16090,N_17695);
nor U21886 (N_21886,N_18220,N_13182);
nand U21887 (N_21887,N_18621,N_14258);
nand U21888 (N_21888,N_12807,N_14522);
and U21889 (N_21889,N_12631,N_14425);
and U21890 (N_21890,N_14856,N_16553);
nand U21891 (N_21891,N_12597,N_13808);
nor U21892 (N_21892,N_14122,N_13015);
or U21893 (N_21893,N_12673,N_18314);
nand U21894 (N_21894,N_15661,N_16375);
xnor U21895 (N_21895,N_13422,N_15513);
or U21896 (N_21896,N_16701,N_15665);
nand U21897 (N_21897,N_15322,N_15958);
or U21898 (N_21898,N_14285,N_17399);
nor U21899 (N_21899,N_13239,N_17001);
or U21900 (N_21900,N_15189,N_14979);
and U21901 (N_21901,N_16491,N_15928);
or U21902 (N_21902,N_16474,N_13940);
nor U21903 (N_21903,N_14308,N_13615);
xnor U21904 (N_21904,N_14737,N_14065);
and U21905 (N_21905,N_18167,N_16978);
or U21906 (N_21906,N_18435,N_15296);
and U21907 (N_21907,N_15488,N_14766);
nand U21908 (N_21908,N_18239,N_18721);
nor U21909 (N_21909,N_15655,N_18537);
and U21910 (N_21910,N_18262,N_18036);
nor U21911 (N_21911,N_13602,N_17845);
and U21912 (N_21912,N_13133,N_13763);
nor U21913 (N_21913,N_17075,N_12758);
nor U21914 (N_21914,N_17937,N_14915);
nand U21915 (N_21915,N_16075,N_15910);
nor U21916 (N_21916,N_13028,N_18124);
xor U21917 (N_21917,N_13677,N_16533);
or U21918 (N_21918,N_13621,N_17981);
and U21919 (N_21919,N_13973,N_13674);
or U21920 (N_21920,N_17875,N_18369);
nor U21921 (N_21921,N_15123,N_16497);
and U21922 (N_21922,N_17052,N_15033);
nor U21923 (N_21923,N_12952,N_17189);
nand U21924 (N_21924,N_13132,N_17975);
or U21925 (N_21925,N_16403,N_17823);
xor U21926 (N_21926,N_17829,N_14771);
nor U21927 (N_21927,N_12795,N_13019);
and U21928 (N_21928,N_16927,N_17093);
or U21929 (N_21929,N_14133,N_17162);
nand U21930 (N_21930,N_18111,N_18347);
xnor U21931 (N_21931,N_17296,N_18605);
nand U21932 (N_21932,N_17055,N_14029);
and U21933 (N_21933,N_16548,N_13486);
or U21934 (N_21934,N_15417,N_12595);
nand U21935 (N_21935,N_16771,N_16680);
and U21936 (N_21936,N_15516,N_18608);
xnor U21937 (N_21937,N_15081,N_13669);
nand U21938 (N_21938,N_12847,N_13185);
xnor U21939 (N_21939,N_14619,N_17637);
nand U21940 (N_21940,N_18450,N_14317);
and U21941 (N_21941,N_13862,N_14072);
or U21942 (N_21942,N_16821,N_14011);
nand U21943 (N_21943,N_13291,N_13762);
or U21944 (N_21944,N_18291,N_13345);
and U21945 (N_21945,N_16276,N_17830);
and U21946 (N_21946,N_14056,N_16161);
or U21947 (N_21947,N_13092,N_16421);
nand U21948 (N_21948,N_16523,N_14356);
nor U21949 (N_21949,N_18350,N_18145);
nor U21950 (N_21950,N_17440,N_15944);
nor U21951 (N_21951,N_13430,N_17314);
and U21952 (N_21952,N_15995,N_18355);
or U21953 (N_21953,N_13230,N_13324);
nand U21954 (N_21954,N_15851,N_18150);
nand U21955 (N_21955,N_14805,N_14356);
or U21956 (N_21956,N_15573,N_18610);
nand U21957 (N_21957,N_15941,N_14803);
or U21958 (N_21958,N_12602,N_17566);
and U21959 (N_21959,N_15074,N_18083);
and U21960 (N_21960,N_13662,N_16552);
nor U21961 (N_21961,N_16445,N_14018);
or U21962 (N_21962,N_14836,N_16578);
nand U21963 (N_21963,N_13080,N_18739);
nand U21964 (N_21964,N_14795,N_15810);
and U21965 (N_21965,N_17209,N_15982);
and U21966 (N_21966,N_17053,N_14958);
nor U21967 (N_21967,N_14677,N_18610);
nor U21968 (N_21968,N_13210,N_18588);
nand U21969 (N_21969,N_14077,N_18357);
nand U21970 (N_21970,N_18272,N_14737);
nand U21971 (N_21971,N_13420,N_17300);
or U21972 (N_21972,N_12656,N_13654);
nor U21973 (N_21973,N_12655,N_18657);
or U21974 (N_21974,N_14190,N_13734);
nor U21975 (N_21975,N_18412,N_17242);
or U21976 (N_21976,N_13413,N_14118);
or U21977 (N_21977,N_14416,N_13724);
xor U21978 (N_21978,N_17906,N_13257);
or U21979 (N_21979,N_14632,N_14830);
nand U21980 (N_21980,N_14593,N_16856);
nor U21981 (N_21981,N_15042,N_18430);
nand U21982 (N_21982,N_15818,N_17703);
nand U21983 (N_21983,N_18393,N_14958);
nor U21984 (N_21984,N_15523,N_13049);
nor U21985 (N_21985,N_16364,N_15242);
nor U21986 (N_21986,N_16805,N_15666);
nor U21987 (N_21987,N_16413,N_17891);
and U21988 (N_21988,N_15760,N_13109);
nand U21989 (N_21989,N_13315,N_16073);
nand U21990 (N_21990,N_14002,N_18387);
nor U21991 (N_21991,N_13714,N_13378);
nor U21992 (N_21992,N_16417,N_17932);
and U21993 (N_21993,N_16182,N_12947);
nor U21994 (N_21994,N_12972,N_14162);
nand U21995 (N_21995,N_18029,N_16217);
nor U21996 (N_21996,N_18152,N_16017);
nand U21997 (N_21997,N_17332,N_14008);
and U21998 (N_21998,N_17704,N_13435);
xnor U21999 (N_21999,N_18356,N_16877);
or U22000 (N_22000,N_14597,N_14356);
and U22001 (N_22001,N_17491,N_15842);
and U22002 (N_22002,N_16121,N_18157);
or U22003 (N_22003,N_18695,N_13603);
and U22004 (N_22004,N_16326,N_16912);
or U22005 (N_22005,N_15380,N_13665);
or U22006 (N_22006,N_15407,N_16263);
nor U22007 (N_22007,N_14342,N_18257);
or U22008 (N_22008,N_13756,N_18069);
nor U22009 (N_22009,N_13410,N_18291);
nor U22010 (N_22010,N_15002,N_15557);
and U22011 (N_22011,N_18222,N_14353);
nor U22012 (N_22012,N_15148,N_16816);
and U22013 (N_22013,N_16030,N_15177);
nand U22014 (N_22014,N_16296,N_17444);
or U22015 (N_22015,N_14204,N_17275);
or U22016 (N_22016,N_15974,N_15742);
nand U22017 (N_22017,N_13628,N_17725);
nand U22018 (N_22018,N_13690,N_15270);
or U22019 (N_22019,N_16475,N_16101);
and U22020 (N_22020,N_15084,N_14545);
nor U22021 (N_22021,N_12871,N_13183);
nand U22022 (N_22022,N_18685,N_15887);
and U22023 (N_22023,N_14091,N_15975);
xnor U22024 (N_22024,N_13409,N_15359);
or U22025 (N_22025,N_14627,N_16999);
or U22026 (N_22026,N_14689,N_15976);
nor U22027 (N_22027,N_18268,N_14252);
nor U22028 (N_22028,N_17298,N_16187);
and U22029 (N_22029,N_14783,N_15977);
nor U22030 (N_22030,N_17048,N_13395);
nor U22031 (N_22031,N_13878,N_14415);
and U22032 (N_22032,N_17288,N_12867);
nand U22033 (N_22033,N_17335,N_17388);
nor U22034 (N_22034,N_18360,N_12693);
nand U22035 (N_22035,N_16121,N_14894);
or U22036 (N_22036,N_16270,N_15456);
nor U22037 (N_22037,N_13767,N_17864);
nand U22038 (N_22038,N_15889,N_15620);
nand U22039 (N_22039,N_15788,N_14877);
nor U22040 (N_22040,N_12952,N_16269);
nand U22041 (N_22041,N_17947,N_16466);
nand U22042 (N_22042,N_16850,N_15819);
nor U22043 (N_22043,N_13822,N_12975);
or U22044 (N_22044,N_14400,N_16984);
nand U22045 (N_22045,N_15750,N_17966);
or U22046 (N_22046,N_17081,N_17068);
or U22047 (N_22047,N_13019,N_13386);
or U22048 (N_22048,N_18664,N_18669);
or U22049 (N_22049,N_13489,N_13432);
or U22050 (N_22050,N_17173,N_15673);
nor U22051 (N_22051,N_14919,N_16066);
nor U22052 (N_22052,N_16457,N_13369);
nand U22053 (N_22053,N_14778,N_13238);
nor U22054 (N_22054,N_13306,N_18414);
or U22055 (N_22055,N_15646,N_12962);
nand U22056 (N_22056,N_15715,N_13885);
nand U22057 (N_22057,N_15225,N_17678);
nor U22058 (N_22058,N_13307,N_14198);
nor U22059 (N_22059,N_13977,N_14893);
nor U22060 (N_22060,N_13684,N_16444);
or U22061 (N_22061,N_15488,N_17869);
nor U22062 (N_22062,N_16486,N_18529);
or U22063 (N_22063,N_14885,N_15601);
and U22064 (N_22064,N_16615,N_18195);
and U22065 (N_22065,N_17719,N_13826);
nor U22066 (N_22066,N_12778,N_13961);
xnor U22067 (N_22067,N_17886,N_18665);
and U22068 (N_22068,N_13290,N_14364);
and U22069 (N_22069,N_18552,N_13833);
and U22070 (N_22070,N_12529,N_15175);
or U22071 (N_22071,N_13629,N_16155);
and U22072 (N_22072,N_15709,N_12757);
nor U22073 (N_22073,N_16753,N_12847);
nor U22074 (N_22074,N_16839,N_17541);
and U22075 (N_22075,N_15440,N_18351);
or U22076 (N_22076,N_14654,N_15354);
or U22077 (N_22077,N_16283,N_16140);
xor U22078 (N_22078,N_13012,N_14699);
or U22079 (N_22079,N_15906,N_12899);
or U22080 (N_22080,N_15925,N_18076);
nor U22081 (N_22081,N_17859,N_14328);
nor U22082 (N_22082,N_17095,N_13855);
nor U22083 (N_22083,N_13885,N_14210);
nand U22084 (N_22084,N_17829,N_15988);
nor U22085 (N_22085,N_14788,N_16070);
and U22086 (N_22086,N_15029,N_17672);
xor U22087 (N_22087,N_17968,N_16795);
nor U22088 (N_22088,N_15109,N_12775);
nor U22089 (N_22089,N_16577,N_13493);
and U22090 (N_22090,N_15142,N_13900);
xnor U22091 (N_22091,N_17684,N_16769);
nand U22092 (N_22092,N_14910,N_12676);
and U22093 (N_22093,N_14225,N_18642);
or U22094 (N_22094,N_14039,N_13469);
nor U22095 (N_22095,N_15824,N_16792);
and U22096 (N_22096,N_15553,N_17414);
and U22097 (N_22097,N_17795,N_17631);
nor U22098 (N_22098,N_15137,N_14186);
or U22099 (N_22099,N_18387,N_17468);
xnor U22100 (N_22100,N_16665,N_15052);
or U22101 (N_22101,N_18073,N_12564);
or U22102 (N_22102,N_15652,N_13400);
or U22103 (N_22103,N_13188,N_13500);
or U22104 (N_22104,N_12804,N_15486);
and U22105 (N_22105,N_15742,N_16715);
nand U22106 (N_22106,N_16307,N_14822);
nand U22107 (N_22107,N_12567,N_12848);
nor U22108 (N_22108,N_15883,N_12703);
and U22109 (N_22109,N_16373,N_15899);
nand U22110 (N_22110,N_13854,N_17064);
nand U22111 (N_22111,N_13358,N_12520);
nand U22112 (N_22112,N_15907,N_15774);
nand U22113 (N_22113,N_16365,N_12644);
and U22114 (N_22114,N_15168,N_15625);
xnor U22115 (N_22115,N_17870,N_13933);
xor U22116 (N_22116,N_16353,N_17799);
and U22117 (N_22117,N_13600,N_15534);
nor U22118 (N_22118,N_13305,N_17617);
and U22119 (N_22119,N_12965,N_14003);
xnor U22120 (N_22120,N_14513,N_14737);
nand U22121 (N_22121,N_14851,N_12883);
or U22122 (N_22122,N_17547,N_16055);
nand U22123 (N_22123,N_14362,N_18395);
nand U22124 (N_22124,N_18621,N_12825);
or U22125 (N_22125,N_16265,N_18457);
nand U22126 (N_22126,N_14866,N_17675);
nor U22127 (N_22127,N_16154,N_17386);
nand U22128 (N_22128,N_15360,N_15031);
nor U22129 (N_22129,N_16678,N_16778);
nand U22130 (N_22130,N_16330,N_16472);
nor U22131 (N_22131,N_17136,N_14936);
nand U22132 (N_22132,N_12580,N_18030);
nand U22133 (N_22133,N_16439,N_18701);
and U22134 (N_22134,N_13519,N_13304);
xor U22135 (N_22135,N_17582,N_16157);
nor U22136 (N_22136,N_16879,N_13449);
nor U22137 (N_22137,N_14645,N_14579);
nand U22138 (N_22138,N_16472,N_17039);
or U22139 (N_22139,N_13180,N_13244);
xor U22140 (N_22140,N_14965,N_16896);
and U22141 (N_22141,N_16895,N_17300);
and U22142 (N_22142,N_15841,N_15374);
or U22143 (N_22143,N_15201,N_17974);
nand U22144 (N_22144,N_17302,N_15331);
nor U22145 (N_22145,N_13976,N_17247);
or U22146 (N_22146,N_14935,N_14883);
nor U22147 (N_22147,N_13142,N_17520);
or U22148 (N_22148,N_16419,N_15994);
nand U22149 (N_22149,N_13725,N_17202);
nor U22150 (N_22150,N_13735,N_14719);
and U22151 (N_22151,N_12920,N_15821);
xnor U22152 (N_22152,N_12846,N_13375);
nand U22153 (N_22153,N_16905,N_15659);
nand U22154 (N_22154,N_18742,N_16696);
and U22155 (N_22155,N_15793,N_17880);
and U22156 (N_22156,N_15264,N_14009);
nor U22157 (N_22157,N_16110,N_15578);
nand U22158 (N_22158,N_13270,N_13204);
or U22159 (N_22159,N_17494,N_15733);
nand U22160 (N_22160,N_18085,N_16883);
nand U22161 (N_22161,N_13532,N_12713);
xnor U22162 (N_22162,N_13901,N_16026);
nor U22163 (N_22163,N_14724,N_14020);
and U22164 (N_22164,N_16410,N_17580);
nand U22165 (N_22165,N_15528,N_12930);
xor U22166 (N_22166,N_17756,N_15696);
nand U22167 (N_22167,N_16825,N_18466);
or U22168 (N_22168,N_15024,N_14467);
nand U22169 (N_22169,N_17783,N_12887);
xor U22170 (N_22170,N_18453,N_14061);
and U22171 (N_22171,N_14798,N_18332);
xnor U22172 (N_22172,N_14797,N_17926);
and U22173 (N_22173,N_15378,N_15063);
nand U22174 (N_22174,N_13194,N_17367);
nor U22175 (N_22175,N_16076,N_18170);
nand U22176 (N_22176,N_14937,N_15811);
nor U22177 (N_22177,N_16634,N_16991);
nor U22178 (N_22178,N_13568,N_18536);
nor U22179 (N_22179,N_13074,N_13195);
nor U22180 (N_22180,N_13749,N_15241);
xor U22181 (N_22181,N_18305,N_15819);
and U22182 (N_22182,N_14988,N_17721);
nand U22183 (N_22183,N_17638,N_16783);
or U22184 (N_22184,N_17506,N_16670);
or U22185 (N_22185,N_15011,N_15566);
nand U22186 (N_22186,N_13400,N_18540);
and U22187 (N_22187,N_17360,N_15735);
xnor U22188 (N_22188,N_12573,N_15210);
or U22189 (N_22189,N_12848,N_16846);
or U22190 (N_22190,N_16053,N_18475);
nor U22191 (N_22191,N_13625,N_15031);
or U22192 (N_22192,N_15850,N_13620);
nor U22193 (N_22193,N_16019,N_18357);
nor U22194 (N_22194,N_14862,N_15777);
and U22195 (N_22195,N_17350,N_17968);
nand U22196 (N_22196,N_18220,N_15544);
nand U22197 (N_22197,N_15663,N_17431);
nor U22198 (N_22198,N_17795,N_13191);
xor U22199 (N_22199,N_17820,N_14328);
or U22200 (N_22200,N_15706,N_17922);
nor U22201 (N_22201,N_18009,N_14475);
and U22202 (N_22202,N_18429,N_15662);
and U22203 (N_22203,N_18013,N_17612);
xnor U22204 (N_22204,N_13943,N_16004);
xnor U22205 (N_22205,N_15711,N_16210);
or U22206 (N_22206,N_13720,N_12649);
and U22207 (N_22207,N_16878,N_16522);
and U22208 (N_22208,N_18728,N_16998);
or U22209 (N_22209,N_15426,N_15939);
or U22210 (N_22210,N_16355,N_17154);
nand U22211 (N_22211,N_12938,N_17958);
or U22212 (N_22212,N_14384,N_18062);
nor U22213 (N_22213,N_17313,N_16482);
nand U22214 (N_22214,N_12925,N_15605);
xor U22215 (N_22215,N_16462,N_18593);
nand U22216 (N_22216,N_13015,N_17532);
nand U22217 (N_22217,N_16811,N_17290);
nand U22218 (N_22218,N_16127,N_18110);
and U22219 (N_22219,N_16887,N_15128);
and U22220 (N_22220,N_15516,N_14695);
xnor U22221 (N_22221,N_13591,N_16324);
nor U22222 (N_22222,N_14676,N_13293);
nor U22223 (N_22223,N_16053,N_13147);
and U22224 (N_22224,N_18707,N_15136);
and U22225 (N_22225,N_14962,N_12762);
nand U22226 (N_22226,N_18629,N_13355);
nor U22227 (N_22227,N_16319,N_15869);
or U22228 (N_22228,N_13680,N_16371);
or U22229 (N_22229,N_17481,N_17892);
nor U22230 (N_22230,N_13495,N_16717);
and U22231 (N_22231,N_16360,N_12789);
nor U22232 (N_22232,N_17660,N_17107);
or U22233 (N_22233,N_18351,N_13124);
nor U22234 (N_22234,N_12791,N_14458);
nor U22235 (N_22235,N_18536,N_12913);
or U22236 (N_22236,N_17976,N_15037);
xnor U22237 (N_22237,N_12536,N_17774);
xor U22238 (N_22238,N_12571,N_13403);
xor U22239 (N_22239,N_17587,N_14011);
and U22240 (N_22240,N_16023,N_16210);
nor U22241 (N_22241,N_18599,N_16814);
nand U22242 (N_22242,N_16901,N_12542);
nand U22243 (N_22243,N_15209,N_18211);
nand U22244 (N_22244,N_13524,N_18700);
and U22245 (N_22245,N_15164,N_15076);
or U22246 (N_22246,N_13071,N_12879);
nor U22247 (N_22247,N_15809,N_13758);
nand U22248 (N_22248,N_13631,N_13226);
nor U22249 (N_22249,N_16178,N_13274);
nor U22250 (N_22250,N_15427,N_13136);
nor U22251 (N_22251,N_13751,N_15768);
nor U22252 (N_22252,N_13817,N_15106);
nand U22253 (N_22253,N_14615,N_18569);
nor U22254 (N_22254,N_13763,N_13968);
or U22255 (N_22255,N_13593,N_15249);
nor U22256 (N_22256,N_18688,N_17675);
nor U22257 (N_22257,N_13122,N_14545);
nand U22258 (N_22258,N_16897,N_15466);
nand U22259 (N_22259,N_17934,N_14281);
and U22260 (N_22260,N_16719,N_15459);
nor U22261 (N_22261,N_14859,N_13996);
nor U22262 (N_22262,N_17097,N_14824);
nor U22263 (N_22263,N_14743,N_14801);
and U22264 (N_22264,N_18464,N_13657);
nand U22265 (N_22265,N_14487,N_15823);
nand U22266 (N_22266,N_16249,N_15967);
nor U22267 (N_22267,N_15068,N_13792);
nand U22268 (N_22268,N_16874,N_14042);
and U22269 (N_22269,N_13064,N_14541);
nand U22270 (N_22270,N_15099,N_14451);
nor U22271 (N_22271,N_12864,N_13550);
xor U22272 (N_22272,N_18701,N_14085);
nand U22273 (N_22273,N_18682,N_18718);
xor U22274 (N_22274,N_17414,N_12521);
and U22275 (N_22275,N_14971,N_13064);
nand U22276 (N_22276,N_13931,N_13051);
and U22277 (N_22277,N_18154,N_13910);
and U22278 (N_22278,N_14828,N_12863);
nor U22279 (N_22279,N_12796,N_16552);
nor U22280 (N_22280,N_16233,N_15856);
nand U22281 (N_22281,N_15703,N_17829);
nand U22282 (N_22282,N_13313,N_16556);
and U22283 (N_22283,N_13779,N_12990);
or U22284 (N_22284,N_17944,N_14256);
or U22285 (N_22285,N_12918,N_16895);
or U22286 (N_22286,N_16937,N_16346);
and U22287 (N_22287,N_16067,N_15313);
nand U22288 (N_22288,N_16415,N_18711);
nor U22289 (N_22289,N_18140,N_15712);
nor U22290 (N_22290,N_12921,N_16147);
or U22291 (N_22291,N_14522,N_13957);
and U22292 (N_22292,N_15028,N_15821);
nand U22293 (N_22293,N_15688,N_17260);
and U22294 (N_22294,N_12700,N_14381);
or U22295 (N_22295,N_13225,N_15639);
or U22296 (N_22296,N_15297,N_17426);
and U22297 (N_22297,N_17759,N_12855);
or U22298 (N_22298,N_16194,N_18045);
or U22299 (N_22299,N_18572,N_12660);
and U22300 (N_22300,N_18563,N_14646);
and U22301 (N_22301,N_14109,N_14029);
nand U22302 (N_22302,N_16919,N_16166);
nor U22303 (N_22303,N_13902,N_13408);
nand U22304 (N_22304,N_15979,N_16868);
nand U22305 (N_22305,N_14813,N_13901);
nor U22306 (N_22306,N_15040,N_18616);
or U22307 (N_22307,N_16576,N_14141);
or U22308 (N_22308,N_18596,N_14076);
and U22309 (N_22309,N_16773,N_18512);
nor U22310 (N_22310,N_14216,N_16470);
xor U22311 (N_22311,N_17529,N_18453);
nand U22312 (N_22312,N_17356,N_12615);
nor U22313 (N_22313,N_18422,N_14540);
nor U22314 (N_22314,N_14848,N_16139);
nand U22315 (N_22315,N_15433,N_14268);
nor U22316 (N_22316,N_13898,N_18358);
nand U22317 (N_22317,N_17074,N_14089);
or U22318 (N_22318,N_17275,N_15969);
nor U22319 (N_22319,N_14396,N_15565);
xor U22320 (N_22320,N_18496,N_14615);
nor U22321 (N_22321,N_13139,N_17276);
nand U22322 (N_22322,N_14368,N_15961);
or U22323 (N_22323,N_16296,N_14650);
nand U22324 (N_22324,N_18512,N_13723);
nor U22325 (N_22325,N_17560,N_16184);
nor U22326 (N_22326,N_12535,N_15923);
and U22327 (N_22327,N_14125,N_12898);
xnor U22328 (N_22328,N_15799,N_16744);
nand U22329 (N_22329,N_16044,N_16800);
or U22330 (N_22330,N_17246,N_13078);
nor U22331 (N_22331,N_17508,N_16320);
or U22332 (N_22332,N_15853,N_17035);
or U22333 (N_22333,N_18419,N_15783);
nand U22334 (N_22334,N_13233,N_13340);
and U22335 (N_22335,N_17596,N_12579);
or U22336 (N_22336,N_16688,N_16151);
nor U22337 (N_22337,N_15572,N_16881);
nand U22338 (N_22338,N_17306,N_14253);
nand U22339 (N_22339,N_18707,N_13050);
nand U22340 (N_22340,N_16935,N_18290);
nand U22341 (N_22341,N_15930,N_13693);
or U22342 (N_22342,N_13148,N_16184);
nor U22343 (N_22343,N_14509,N_18054);
nor U22344 (N_22344,N_14228,N_16087);
and U22345 (N_22345,N_14206,N_17854);
and U22346 (N_22346,N_16831,N_15007);
nand U22347 (N_22347,N_16779,N_17925);
nor U22348 (N_22348,N_17400,N_13719);
and U22349 (N_22349,N_14043,N_16158);
and U22350 (N_22350,N_15036,N_12785);
xnor U22351 (N_22351,N_15212,N_15671);
or U22352 (N_22352,N_16831,N_13846);
or U22353 (N_22353,N_15208,N_14411);
nor U22354 (N_22354,N_17536,N_15466);
xnor U22355 (N_22355,N_15841,N_17506);
nor U22356 (N_22356,N_16762,N_15056);
or U22357 (N_22357,N_15611,N_13917);
nand U22358 (N_22358,N_18104,N_16675);
nor U22359 (N_22359,N_16493,N_13472);
nand U22360 (N_22360,N_16040,N_15795);
nor U22361 (N_22361,N_13660,N_13853);
or U22362 (N_22362,N_16192,N_18365);
nor U22363 (N_22363,N_17921,N_12814);
nor U22364 (N_22364,N_12861,N_14009);
nor U22365 (N_22365,N_13679,N_15605);
nand U22366 (N_22366,N_14554,N_13964);
nor U22367 (N_22367,N_18496,N_15031);
or U22368 (N_22368,N_14802,N_16062);
and U22369 (N_22369,N_13923,N_15423);
nand U22370 (N_22370,N_13359,N_16198);
nand U22371 (N_22371,N_14301,N_17535);
xor U22372 (N_22372,N_14627,N_16728);
and U22373 (N_22373,N_17796,N_14865);
nor U22374 (N_22374,N_17770,N_12724);
nor U22375 (N_22375,N_12550,N_14228);
nand U22376 (N_22376,N_18069,N_13877);
nor U22377 (N_22377,N_13912,N_12637);
nand U22378 (N_22378,N_16290,N_18276);
nand U22379 (N_22379,N_13407,N_14007);
and U22380 (N_22380,N_14467,N_13107);
xnor U22381 (N_22381,N_16574,N_18403);
nor U22382 (N_22382,N_17272,N_12846);
nor U22383 (N_22383,N_12700,N_13074);
or U22384 (N_22384,N_14332,N_17747);
nand U22385 (N_22385,N_12587,N_14309);
nor U22386 (N_22386,N_14438,N_17727);
nand U22387 (N_22387,N_13238,N_16355);
nand U22388 (N_22388,N_13843,N_18246);
and U22389 (N_22389,N_13462,N_15470);
or U22390 (N_22390,N_14592,N_13823);
nor U22391 (N_22391,N_13787,N_13345);
or U22392 (N_22392,N_18016,N_16424);
and U22393 (N_22393,N_13277,N_13220);
or U22394 (N_22394,N_14801,N_13703);
xor U22395 (N_22395,N_14456,N_13101);
xnor U22396 (N_22396,N_17216,N_15875);
and U22397 (N_22397,N_13341,N_13157);
and U22398 (N_22398,N_15863,N_13065);
and U22399 (N_22399,N_16284,N_15685);
xnor U22400 (N_22400,N_14619,N_17265);
xnor U22401 (N_22401,N_14860,N_17202);
and U22402 (N_22402,N_12949,N_18461);
and U22403 (N_22403,N_13440,N_14158);
nand U22404 (N_22404,N_14587,N_15165);
nor U22405 (N_22405,N_15952,N_18724);
or U22406 (N_22406,N_14462,N_15423);
and U22407 (N_22407,N_15564,N_16408);
nand U22408 (N_22408,N_13361,N_13265);
and U22409 (N_22409,N_18508,N_18033);
nor U22410 (N_22410,N_13863,N_16796);
nor U22411 (N_22411,N_14234,N_18123);
or U22412 (N_22412,N_18176,N_18019);
or U22413 (N_22413,N_16321,N_13798);
nand U22414 (N_22414,N_13251,N_16310);
or U22415 (N_22415,N_14659,N_18324);
nor U22416 (N_22416,N_14254,N_13029);
and U22417 (N_22417,N_12835,N_12597);
and U22418 (N_22418,N_17649,N_13974);
nand U22419 (N_22419,N_15930,N_16125);
nand U22420 (N_22420,N_16985,N_17856);
or U22421 (N_22421,N_18280,N_18265);
or U22422 (N_22422,N_17284,N_17932);
xnor U22423 (N_22423,N_15742,N_13719);
nor U22424 (N_22424,N_15184,N_17983);
and U22425 (N_22425,N_18689,N_14862);
or U22426 (N_22426,N_13175,N_18555);
and U22427 (N_22427,N_13664,N_13596);
or U22428 (N_22428,N_13242,N_15641);
and U22429 (N_22429,N_16788,N_17034);
or U22430 (N_22430,N_16199,N_17859);
and U22431 (N_22431,N_12992,N_13066);
and U22432 (N_22432,N_16664,N_12652);
nand U22433 (N_22433,N_12916,N_16222);
and U22434 (N_22434,N_13787,N_18397);
or U22435 (N_22435,N_16325,N_17562);
nand U22436 (N_22436,N_17837,N_15005);
nand U22437 (N_22437,N_18726,N_13014);
or U22438 (N_22438,N_15343,N_12857);
nand U22439 (N_22439,N_13223,N_14594);
nor U22440 (N_22440,N_14786,N_14684);
nand U22441 (N_22441,N_18401,N_13194);
nand U22442 (N_22442,N_15330,N_16029);
and U22443 (N_22443,N_14983,N_13792);
nand U22444 (N_22444,N_13731,N_12603);
and U22445 (N_22445,N_18598,N_15681);
nand U22446 (N_22446,N_13773,N_13466);
and U22447 (N_22447,N_14780,N_16861);
and U22448 (N_22448,N_17656,N_14238);
nand U22449 (N_22449,N_16852,N_16461);
or U22450 (N_22450,N_14750,N_15012);
and U22451 (N_22451,N_14864,N_16609);
and U22452 (N_22452,N_13947,N_16902);
nand U22453 (N_22453,N_15727,N_17743);
or U22454 (N_22454,N_18417,N_17436);
and U22455 (N_22455,N_15113,N_12897);
nand U22456 (N_22456,N_12936,N_13918);
and U22457 (N_22457,N_17589,N_13689);
or U22458 (N_22458,N_12911,N_16326);
nor U22459 (N_22459,N_16282,N_17486);
xor U22460 (N_22460,N_15343,N_14690);
and U22461 (N_22461,N_17737,N_17114);
nand U22462 (N_22462,N_18226,N_14250);
nor U22463 (N_22463,N_15585,N_15765);
and U22464 (N_22464,N_15056,N_13740);
nor U22465 (N_22465,N_13061,N_15636);
nor U22466 (N_22466,N_15339,N_18343);
and U22467 (N_22467,N_16396,N_13594);
or U22468 (N_22468,N_17749,N_15943);
and U22469 (N_22469,N_13990,N_14287);
and U22470 (N_22470,N_13281,N_14543);
or U22471 (N_22471,N_15885,N_18467);
nand U22472 (N_22472,N_12629,N_16260);
nand U22473 (N_22473,N_15061,N_16408);
and U22474 (N_22474,N_15264,N_12933);
nand U22475 (N_22475,N_17969,N_13940);
or U22476 (N_22476,N_18629,N_17773);
nor U22477 (N_22477,N_12956,N_16727);
nand U22478 (N_22478,N_18421,N_18066);
nand U22479 (N_22479,N_16981,N_13630);
nor U22480 (N_22480,N_13157,N_15501);
xor U22481 (N_22481,N_16694,N_15049);
nor U22482 (N_22482,N_14238,N_15761);
nor U22483 (N_22483,N_15409,N_16299);
nor U22484 (N_22484,N_14092,N_13237);
or U22485 (N_22485,N_14261,N_18561);
or U22486 (N_22486,N_16296,N_16981);
nor U22487 (N_22487,N_14624,N_15180);
nor U22488 (N_22488,N_12991,N_18599);
xor U22489 (N_22489,N_13224,N_13960);
and U22490 (N_22490,N_16698,N_14794);
nor U22491 (N_22491,N_14978,N_13002);
and U22492 (N_22492,N_13984,N_15412);
and U22493 (N_22493,N_13026,N_12961);
nor U22494 (N_22494,N_16623,N_17268);
xor U22495 (N_22495,N_13981,N_17974);
or U22496 (N_22496,N_15797,N_14787);
nand U22497 (N_22497,N_16152,N_13927);
and U22498 (N_22498,N_14611,N_14777);
nor U22499 (N_22499,N_18645,N_17444);
nor U22500 (N_22500,N_16628,N_18023);
nand U22501 (N_22501,N_12652,N_17080);
xnor U22502 (N_22502,N_14539,N_17952);
or U22503 (N_22503,N_17892,N_13232);
nor U22504 (N_22504,N_15809,N_15057);
or U22505 (N_22505,N_15035,N_17013);
nor U22506 (N_22506,N_15770,N_18036);
or U22507 (N_22507,N_15964,N_16264);
or U22508 (N_22508,N_18598,N_16177);
nand U22509 (N_22509,N_13245,N_14275);
nor U22510 (N_22510,N_17947,N_15069);
xnor U22511 (N_22511,N_12809,N_17369);
nand U22512 (N_22512,N_15796,N_16781);
and U22513 (N_22513,N_18647,N_16541);
and U22514 (N_22514,N_17041,N_17514);
nor U22515 (N_22515,N_12961,N_17404);
nor U22516 (N_22516,N_17800,N_18612);
and U22517 (N_22517,N_18117,N_15382);
nand U22518 (N_22518,N_13436,N_18447);
nand U22519 (N_22519,N_15845,N_14095);
or U22520 (N_22520,N_16456,N_18512);
nor U22521 (N_22521,N_18071,N_16387);
xnor U22522 (N_22522,N_12766,N_12571);
and U22523 (N_22523,N_13731,N_14310);
nand U22524 (N_22524,N_18662,N_17741);
or U22525 (N_22525,N_14933,N_14626);
and U22526 (N_22526,N_17055,N_17888);
or U22527 (N_22527,N_12590,N_13657);
and U22528 (N_22528,N_16919,N_13325);
or U22529 (N_22529,N_14536,N_17586);
nor U22530 (N_22530,N_12597,N_13120);
or U22531 (N_22531,N_14010,N_12873);
xor U22532 (N_22532,N_16875,N_17285);
and U22533 (N_22533,N_13160,N_18377);
or U22534 (N_22534,N_18494,N_18302);
nor U22535 (N_22535,N_14811,N_18042);
and U22536 (N_22536,N_12922,N_18408);
nor U22537 (N_22537,N_15758,N_14100);
nand U22538 (N_22538,N_18673,N_17535);
nand U22539 (N_22539,N_12583,N_17085);
or U22540 (N_22540,N_14648,N_18718);
nor U22541 (N_22541,N_16518,N_17264);
nor U22542 (N_22542,N_16245,N_15700);
or U22543 (N_22543,N_12900,N_17806);
nor U22544 (N_22544,N_15462,N_16848);
and U22545 (N_22545,N_15851,N_14487);
nor U22546 (N_22546,N_13614,N_18046);
nor U22547 (N_22547,N_12983,N_15670);
and U22548 (N_22548,N_18601,N_14897);
nor U22549 (N_22549,N_16538,N_16742);
and U22550 (N_22550,N_13138,N_14289);
or U22551 (N_22551,N_14449,N_13015);
and U22552 (N_22552,N_14562,N_15663);
nand U22553 (N_22553,N_15487,N_13512);
nand U22554 (N_22554,N_15547,N_12686);
nor U22555 (N_22555,N_12683,N_17959);
nand U22556 (N_22556,N_18436,N_16462);
and U22557 (N_22557,N_16530,N_14616);
nand U22558 (N_22558,N_15666,N_16111);
xor U22559 (N_22559,N_17690,N_16539);
xnor U22560 (N_22560,N_18049,N_12875);
and U22561 (N_22561,N_18221,N_13600);
and U22562 (N_22562,N_17647,N_18550);
or U22563 (N_22563,N_15336,N_13404);
or U22564 (N_22564,N_18234,N_17105);
or U22565 (N_22565,N_16957,N_14618);
or U22566 (N_22566,N_15048,N_15709);
and U22567 (N_22567,N_16323,N_12881);
and U22568 (N_22568,N_14930,N_18364);
nor U22569 (N_22569,N_16110,N_15991);
nand U22570 (N_22570,N_16109,N_18606);
or U22571 (N_22571,N_16238,N_13109);
or U22572 (N_22572,N_17893,N_15235);
nor U22573 (N_22573,N_16798,N_14181);
nor U22574 (N_22574,N_15684,N_18721);
nand U22575 (N_22575,N_15792,N_18232);
nand U22576 (N_22576,N_12927,N_18265);
nor U22577 (N_22577,N_17335,N_17492);
xnor U22578 (N_22578,N_12511,N_14635);
or U22579 (N_22579,N_17973,N_18445);
nand U22580 (N_22580,N_17038,N_13748);
nor U22581 (N_22581,N_16978,N_18625);
nor U22582 (N_22582,N_15324,N_17653);
nor U22583 (N_22583,N_18188,N_14676);
nand U22584 (N_22584,N_13843,N_13951);
and U22585 (N_22585,N_17155,N_14696);
nand U22586 (N_22586,N_16290,N_15230);
nand U22587 (N_22587,N_12981,N_13618);
nor U22588 (N_22588,N_17420,N_15168);
or U22589 (N_22589,N_17265,N_15915);
and U22590 (N_22590,N_16657,N_13823);
or U22591 (N_22591,N_17301,N_15047);
nor U22592 (N_22592,N_17553,N_18544);
and U22593 (N_22593,N_14085,N_18322);
nor U22594 (N_22594,N_14604,N_18234);
or U22595 (N_22595,N_13716,N_15327);
xor U22596 (N_22596,N_16278,N_16943);
xor U22597 (N_22597,N_13001,N_15148);
or U22598 (N_22598,N_13994,N_17914);
or U22599 (N_22599,N_15421,N_13573);
or U22600 (N_22600,N_14553,N_15585);
and U22601 (N_22601,N_17064,N_17774);
nand U22602 (N_22602,N_12955,N_16636);
and U22603 (N_22603,N_18290,N_13926);
nor U22604 (N_22604,N_15699,N_12868);
and U22605 (N_22605,N_15156,N_14083);
or U22606 (N_22606,N_14700,N_16214);
nor U22607 (N_22607,N_14787,N_12594);
nand U22608 (N_22608,N_14984,N_17029);
nand U22609 (N_22609,N_14011,N_14264);
nand U22610 (N_22610,N_12675,N_17603);
nand U22611 (N_22611,N_18048,N_13161);
and U22612 (N_22612,N_15251,N_18393);
or U22613 (N_22613,N_13600,N_18484);
and U22614 (N_22614,N_16626,N_16130);
nor U22615 (N_22615,N_17223,N_17543);
nor U22616 (N_22616,N_12708,N_18214);
nand U22617 (N_22617,N_15428,N_13255);
or U22618 (N_22618,N_17753,N_17527);
nand U22619 (N_22619,N_15026,N_13625);
nor U22620 (N_22620,N_14893,N_13071);
and U22621 (N_22621,N_16539,N_14310);
nand U22622 (N_22622,N_16440,N_17923);
nor U22623 (N_22623,N_17890,N_16520);
xnor U22624 (N_22624,N_14704,N_15091);
nor U22625 (N_22625,N_15380,N_18277);
and U22626 (N_22626,N_17338,N_12844);
nor U22627 (N_22627,N_14606,N_13604);
nand U22628 (N_22628,N_14828,N_18326);
xor U22629 (N_22629,N_14626,N_16493);
and U22630 (N_22630,N_13779,N_12676);
or U22631 (N_22631,N_15387,N_15705);
and U22632 (N_22632,N_14797,N_14346);
or U22633 (N_22633,N_16524,N_18188);
and U22634 (N_22634,N_16965,N_13689);
nor U22635 (N_22635,N_12838,N_18712);
nand U22636 (N_22636,N_15569,N_15615);
or U22637 (N_22637,N_14023,N_16482);
or U22638 (N_22638,N_15529,N_13058);
nand U22639 (N_22639,N_17008,N_12773);
and U22640 (N_22640,N_15697,N_14068);
nand U22641 (N_22641,N_14924,N_12862);
and U22642 (N_22642,N_15482,N_17403);
xor U22643 (N_22643,N_13387,N_14520);
nand U22644 (N_22644,N_16862,N_13996);
xor U22645 (N_22645,N_18505,N_18301);
xor U22646 (N_22646,N_15721,N_14416);
xor U22647 (N_22647,N_14525,N_15613);
or U22648 (N_22648,N_13944,N_14905);
and U22649 (N_22649,N_14119,N_15873);
nand U22650 (N_22650,N_13833,N_13262);
or U22651 (N_22651,N_14758,N_15437);
and U22652 (N_22652,N_14066,N_14715);
nand U22653 (N_22653,N_18311,N_15549);
nand U22654 (N_22654,N_16474,N_17817);
nor U22655 (N_22655,N_14041,N_13369);
nand U22656 (N_22656,N_12588,N_12613);
or U22657 (N_22657,N_16556,N_12514);
xor U22658 (N_22658,N_13468,N_17556);
nor U22659 (N_22659,N_12601,N_16392);
and U22660 (N_22660,N_17497,N_13117);
and U22661 (N_22661,N_16290,N_14627);
nand U22662 (N_22662,N_16018,N_13850);
and U22663 (N_22663,N_17496,N_17328);
and U22664 (N_22664,N_18246,N_13599);
nand U22665 (N_22665,N_17557,N_17825);
xnor U22666 (N_22666,N_12540,N_15797);
nand U22667 (N_22667,N_14663,N_18725);
or U22668 (N_22668,N_14180,N_17461);
nand U22669 (N_22669,N_16966,N_15410);
nor U22670 (N_22670,N_15527,N_15822);
xor U22671 (N_22671,N_17418,N_17975);
xor U22672 (N_22672,N_18201,N_15415);
or U22673 (N_22673,N_15778,N_14144);
or U22674 (N_22674,N_18304,N_13896);
nand U22675 (N_22675,N_15825,N_17720);
nor U22676 (N_22676,N_15374,N_15595);
and U22677 (N_22677,N_13463,N_15927);
or U22678 (N_22678,N_15904,N_14305);
nand U22679 (N_22679,N_14314,N_16477);
nor U22680 (N_22680,N_14725,N_18202);
nor U22681 (N_22681,N_16392,N_17869);
nand U22682 (N_22682,N_14810,N_18605);
or U22683 (N_22683,N_15680,N_14250);
nor U22684 (N_22684,N_15498,N_16200);
and U22685 (N_22685,N_15435,N_16952);
or U22686 (N_22686,N_13661,N_15515);
nand U22687 (N_22687,N_12647,N_14429);
or U22688 (N_22688,N_17575,N_12783);
and U22689 (N_22689,N_14004,N_12899);
nor U22690 (N_22690,N_18724,N_16413);
and U22691 (N_22691,N_16182,N_14018);
and U22692 (N_22692,N_13299,N_13507);
nand U22693 (N_22693,N_18508,N_15275);
or U22694 (N_22694,N_15317,N_16498);
nor U22695 (N_22695,N_12875,N_14318);
nand U22696 (N_22696,N_18043,N_16687);
nand U22697 (N_22697,N_18095,N_14428);
and U22698 (N_22698,N_15093,N_13224);
or U22699 (N_22699,N_18409,N_14179);
and U22700 (N_22700,N_17405,N_12724);
nor U22701 (N_22701,N_16657,N_15891);
nor U22702 (N_22702,N_18378,N_18068);
nand U22703 (N_22703,N_18330,N_17665);
or U22704 (N_22704,N_15141,N_16016);
nand U22705 (N_22705,N_15296,N_13520);
or U22706 (N_22706,N_16925,N_12896);
nor U22707 (N_22707,N_17184,N_16211);
and U22708 (N_22708,N_13108,N_14425);
and U22709 (N_22709,N_15549,N_13531);
and U22710 (N_22710,N_13584,N_12698);
nand U22711 (N_22711,N_13745,N_17353);
or U22712 (N_22712,N_16515,N_16269);
nor U22713 (N_22713,N_15256,N_16967);
or U22714 (N_22714,N_17377,N_16515);
and U22715 (N_22715,N_15168,N_17304);
and U22716 (N_22716,N_14448,N_16739);
and U22717 (N_22717,N_18393,N_18372);
nor U22718 (N_22718,N_17433,N_16987);
nand U22719 (N_22719,N_16686,N_14207);
or U22720 (N_22720,N_18440,N_13123);
nand U22721 (N_22721,N_17646,N_12707);
or U22722 (N_22722,N_14158,N_17905);
nor U22723 (N_22723,N_15681,N_13128);
or U22724 (N_22724,N_13617,N_13678);
nand U22725 (N_22725,N_16558,N_14064);
or U22726 (N_22726,N_13170,N_15618);
or U22727 (N_22727,N_13003,N_17902);
nand U22728 (N_22728,N_13175,N_16573);
xnor U22729 (N_22729,N_14854,N_17564);
or U22730 (N_22730,N_15827,N_18611);
and U22731 (N_22731,N_12544,N_15930);
and U22732 (N_22732,N_13634,N_18424);
xor U22733 (N_22733,N_16697,N_15996);
or U22734 (N_22734,N_17215,N_16951);
nor U22735 (N_22735,N_12686,N_13557);
xor U22736 (N_22736,N_16005,N_14666);
nor U22737 (N_22737,N_14458,N_18053);
xnor U22738 (N_22738,N_12734,N_18103);
nor U22739 (N_22739,N_13025,N_15090);
nor U22740 (N_22740,N_17347,N_17227);
or U22741 (N_22741,N_16157,N_17922);
nor U22742 (N_22742,N_14959,N_16260);
or U22743 (N_22743,N_14782,N_15249);
xnor U22744 (N_22744,N_16818,N_14179);
nor U22745 (N_22745,N_17085,N_14141);
or U22746 (N_22746,N_14127,N_15740);
and U22747 (N_22747,N_15934,N_16789);
and U22748 (N_22748,N_17197,N_15016);
xnor U22749 (N_22749,N_13016,N_13867);
nand U22750 (N_22750,N_14878,N_16450);
or U22751 (N_22751,N_15306,N_13936);
nand U22752 (N_22752,N_17165,N_16011);
and U22753 (N_22753,N_15925,N_14215);
or U22754 (N_22754,N_18332,N_14076);
and U22755 (N_22755,N_12566,N_18307);
and U22756 (N_22756,N_14769,N_18636);
and U22757 (N_22757,N_17188,N_13457);
nand U22758 (N_22758,N_13082,N_18413);
or U22759 (N_22759,N_13055,N_14445);
nor U22760 (N_22760,N_15440,N_18454);
xnor U22761 (N_22761,N_14650,N_18277);
and U22762 (N_22762,N_14967,N_16873);
nor U22763 (N_22763,N_16399,N_15440);
xor U22764 (N_22764,N_18738,N_18499);
or U22765 (N_22765,N_15025,N_13076);
nand U22766 (N_22766,N_17682,N_13924);
nand U22767 (N_22767,N_18302,N_15551);
or U22768 (N_22768,N_16292,N_13866);
nor U22769 (N_22769,N_14421,N_13162);
nand U22770 (N_22770,N_14997,N_14662);
nand U22771 (N_22771,N_14851,N_14122);
or U22772 (N_22772,N_12525,N_17246);
and U22773 (N_22773,N_12659,N_15543);
and U22774 (N_22774,N_18183,N_12625);
nor U22775 (N_22775,N_18589,N_15581);
and U22776 (N_22776,N_16396,N_14741);
nand U22777 (N_22777,N_17347,N_18007);
xnor U22778 (N_22778,N_13176,N_16957);
and U22779 (N_22779,N_17709,N_12858);
nor U22780 (N_22780,N_17589,N_16091);
nor U22781 (N_22781,N_13000,N_13240);
or U22782 (N_22782,N_14121,N_13168);
xor U22783 (N_22783,N_13727,N_14526);
nand U22784 (N_22784,N_16606,N_14113);
xor U22785 (N_22785,N_16957,N_15431);
and U22786 (N_22786,N_12568,N_18429);
and U22787 (N_22787,N_16610,N_17157);
and U22788 (N_22788,N_13549,N_12696);
or U22789 (N_22789,N_18027,N_16821);
nand U22790 (N_22790,N_18146,N_13757);
nand U22791 (N_22791,N_17437,N_12761);
and U22792 (N_22792,N_14017,N_14893);
nor U22793 (N_22793,N_17224,N_18202);
and U22794 (N_22794,N_13645,N_16585);
nor U22795 (N_22795,N_18076,N_15515);
nor U22796 (N_22796,N_12835,N_15953);
nor U22797 (N_22797,N_13739,N_14310);
nand U22798 (N_22798,N_15719,N_14733);
xor U22799 (N_22799,N_13953,N_14187);
nand U22800 (N_22800,N_16925,N_17885);
or U22801 (N_22801,N_15211,N_14652);
and U22802 (N_22802,N_16063,N_17425);
or U22803 (N_22803,N_15720,N_14903);
or U22804 (N_22804,N_16964,N_17753);
xor U22805 (N_22805,N_17581,N_14708);
and U22806 (N_22806,N_18556,N_16886);
or U22807 (N_22807,N_14072,N_17475);
or U22808 (N_22808,N_16756,N_15565);
or U22809 (N_22809,N_13871,N_14621);
xnor U22810 (N_22810,N_18100,N_16560);
or U22811 (N_22811,N_16688,N_15668);
or U22812 (N_22812,N_14611,N_16278);
nand U22813 (N_22813,N_12580,N_18583);
nand U22814 (N_22814,N_13984,N_14735);
or U22815 (N_22815,N_16704,N_17754);
xnor U22816 (N_22816,N_14663,N_15950);
nand U22817 (N_22817,N_15020,N_17640);
or U22818 (N_22818,N_18307,N_13892);
nand U22819 (N_22819,N_16418,N_17503);
or U22820 (N_22820,N_14940,N_16275);
and U22821 (N_22821,N_17277,N_16315);
and U22822 (N_22822,N_15005,N_15003);
nor U22823 (N_22823,N_15549,N_18490);
or U22824 (N_22824,N_14937,N_12974);
nand U22825 (N_22825,N_17189,N_16102);
and U22826 (N_22826,N_14158,N_18076);
xor U22827 (N_22827,N_17677,N_14108);
and U22828 (N_22828,N_15731,N_18077);
nor U22829 (N_22829,N_12753,N_18251);
or U22830 (N_22830,N_18188,N_17007);
or U22831 (N_22831,N_15885,N_15789);
nand U22832 (N_22832,N_16277,N_17417);
nor U22833 (N_22833,N_18420,N_15542);
nor U22834 (N_22834,N_16987,N_12681);
or U22835 (N_22835,N_17693,N_14931);
nor U22836 (N_22836,N_14010,N_15321);
nor U22837 (N_22837,N_15098,N_17041);
nor U22838 (N_22838,N_12583,N_14644);
nor U22839 (N_22839,N_17278,N_14776);
and U22840 (N_22840,N_13126,N_17478);
or U22841 (N_22841,N_14577,N_16269);
and U22842 (N_22842,N_12860,N_16452);
or U22843 (N_22843,N_14030,N_17161);
and U22844 (N_22844,N_13359,N_17382);
nor U22845 (N_22845,N_14547,N_17908);
and U22846 (N_22846,N_18538,N_14582);
nor U22847 (N_22847,N_17953,N_18373);
nand U22848 (N_22848,N_16945,N_18446);
or U22849 (N_22849,N_13306,N_15758);
nor U22850 (N_22850,N_14083,N_18673);
and U22851 (N_22851,N_17872,N_18707);
nand U22852 (N_22852,N_13925,N_14061);
or U22853 (N_22853,N_16201,N_15486);
or U22854 (N_22854,N_14469,N_16959);
nor U22855 (N_22855,N_12897,N_18172);
nand U22856 (N_22856,N_14686,N_14618);
or U22857 (N_22857,N_17890,N_13322);
and U22858 (N_22858,N_15088,N_16645);
xnor U22859 (N_22859,N_17993,N_14673);
and U22860 (N_22860,N_14232,N_14073);
or U22861 (N_22861,N_13692,N_14908);
or U22862 (N_22862,N_16445,N_15114);
nand U22863 (N_22863,N_18090,N_17307);
nor U22864 (N_22864,N_16448,N_17814);
nand U22865 (N_22865,N_12967,N_14036);
nand U22866 (N_22866,N_13598,N_14145);
xor U22867 (N_22867,N_13846,N_15206);
or U22868 (N_22868,N_13083,N_13226);
or U22869 (N_22869,N_12800,N_15956);
xor U22870 (N_22870,N_14096,N_17176);
and U22871 (N_22871,N_16346,N_15897);
or U22872 (N_22872,N_13389,N_16306);
nor U22873 (N_22873,N_13648,N_13178);
or U22874 (N_22874,N_12507,N_13664);
and U22875 (N_22875,N_13508,N_14253);
and U22876 (N_22876,N_14240,N_16796);
and U22877 (N_22877,N_16523,N_15534);
nor U22878 (N_22878,N_14860,N_12557);
xor U22879 (N_22879,N_15678,N_12947);
nand U22880 (N_22880,N_18125,N_16319);
nand U22881 (N_22881,N_16253,N_13875);
nor U22882 (N_22882,N_17844,N_15033);
or U22883 (N_22883,N_14417,N_13177);
nor U22884 (N_22884,N_14420,N_13274);
nand U22885 (N_22885,N_17628,N_13858);
xor U22886 (N_22886,N_15775,N_12827);
and U22887 (N_22887,N_12705,N_13296);
nor U22888 (N_22888,N_18063,N_16053);
and U22889 (N_22889,N_16924,N_15248);
nor U22890 (N_22890,N_12985,N_17202);
nor U22891 (N_22891,N_15256,N_12836);
nor U22892 (N_22892,N_15901,N_13737);
nor U22893 (N_22893,N_15011,N_16716);
or U22894 (N_22894,N_17137,N_12757);
nor U22895 (N_22895,N_14320,N_16303);
nand U22896 (N_22896,N_17431,N_17415);
nor U22897 (N_22897,N_17288,N_13126);
xnor U22898 (N_22898,N_18185,N_13228);
or U22899 (N_22899,N_13694,N_12500);
and U22900 (N_22900,N_16266,N_12805);
xnor U22901 (N_22901,N_18031,N_16362);
nand U22902 (N_22902,N_14088,N_12528);
or U22903 (N_22903,N_17075,N_13567);
nand U22904 (N_22904,N_13326,N_17736);
nor U22905 (N_22905,N_16827,N_12986);
nor U22906 (N_22906,N_13091,N_17870);
or U22907 (N_22907,N_16244,N_18689);
or U22908 (N_22908,N_18224,N_18550);
or U22909 (N_22909,N_13827,N_16869);
nor U22910 (N_22910,N_18741,N_15538);
nor U22911 (N_22911,N_18282,N_13385);
nand U22912 (N_22912,N_14022,N_12626);
nand U22913 (N_22913,N_16992,N_12688);
nor U22914 (N_22914,N_17023,N_16399);
or U22915 (N_22915,N_12861,N_13619);
nand U22916 (N_22916,N_14778,N_14187);
and U22917 (N_22917,N_14244,N_14002);
nor U22918 (N_22918,N_17643,N_15257);
or U22919 (N_22919,N_17057,N_14995);
or U22920 (N_22920,N_16381,N_14206);
or U22921 (N_22921,N_17290,N_15533);
nor U22922 (N_22922,N_14498,N_13512);
nand U22923 (N_22923,N_15476,N_16242);
or U22924 (N_22924,N_14917,N_14799);
or U22925 (N_22925,N_18149,N_12612);
and U22926 (N_22926,N_18105,N_12838);
nand U22927 (N_22927,N_16526,N_12891);
and U22928 (N_22928,N_16216,N_17264);
and U22929 (N_22929,N_14525,N_16825);
nor U22930 (N_22930,N_17844,N_16943);
nor U22931 (N_22931,N_16532,N_16589);
and U22932 (N_22932,N_18419,N_15222);
nor U22933 (N_22933,N_15008,N_16742);
nand U22934 (N_22934,N_18660,N_16678);
or U22935 (N_22935,N_15123,N_15772);
and U22936 (N_22936,N_18638,N_16457);
and U22937 (N_22937,N_13617,N_15562);
nor U22938 (N_22938,N_16872,N_16893);
nor U22939 (N_22939,N_16533,N_17259);
nor U22940 (N_22940,N_16017,N_16060);
nor U22941 (N_22941,N_18433,N_17425);
and U22942 (N_22942,N_15589,N_12904);
or U22943 (N_22943,N_14093,N_17303);
nor U22944 (N_22944,N_16099,N_16077);
nand U22945 (N_22945,N_18694,N_14151);
nor U22946 (N_22946,N_13000,N_16430);
nand U22947 (N_22947,N_17336,N_13281);
and U22948 (N_22948,N_14681,N_17591);
nor U22949 (N_22949,N_13934,N_13858);
and U22950 (N_22950,N_15212,N_14988);
xnor U22951 (N_22951,N_18268,N_13720);
or U22952 (N_22952,N_17660,N_17479);
or U22953 (N_22953,N_14548,N_16771);
nor U22954 (N_22954,N_12817,N_13705);
nand U22955 (N_22955,N_12629,N_18290);
and U22956 (N_22956,N_15897,N_14430);
or U22957 (N_22957,N_18453,N_17414);
nand U22958 (N_22958,N_12859,N_15560);
nor U22959 (N_22959,N_15933,N_17182);
nand U22960 (N_22960,N_15572,N_18483);
or U22961 (N_22961,N_15699,N_13484);
nand U22962 (N_22962,N_13833,N_18162);
and U22963 (N_22963,N_16226,N_15530);
nand U22964 (N_22964,N_15106,N_12874);
or U22965 (N_22965,N_13289,N_12854);
nand U22966 (N_22966,N_13042,N_16463);
or U22967 (N_22967,N_17441,N_16100);
nor U22968 (N_22968,N_13164,N_18534);
or U22969 (N_22969,N_18400,N_13005);
nand U22970 (N_22970,N_17949,N_18489);
nor U22971 (N_22971,N_13409,N_14076);
or U22972 (N_22972,N_16370,N_14593);
or U22973 (N_22973,N_16910,N_15580);
or U22974 (N_22974,N_16673,N_14523);
and U22975 (N_22975,N_13113,N_16687);
nor U22976 (N_22976,N_13778,N_15530);
nand U22977 (N_22977,N_14274,N_18037);
nor U22978 (N_22978,N_15341,N_14242);
xnor U22979 (N_22979,N_18097,N_14386);
and U22980 (N_22980,N_17336,N_17569);
nor U22981 (N_22981,N_16922,N_17266);
and U22982 (N_22982,N_17843,N_18189);
or U22983 (N_22983,N_18558,N_18377);
and U22984 (N_22984,N_13338,N_14388);
nand U22985 (N_22985,N_12629,N_14896);
xnor U22986 (N_22986,N_14029,N_13204);
or U22987 (N_22987,N_17540,N_12724);
or U22988 (N_22988,N_17322,N_14411);
or U22989 (N_22989,N_17192,N_17895);
or U22990 (N_22990,N_18695,N_18690);
nand U22991 (N_22991,N_13110,N_12815);
nor U22992 (N_22992,N_14106,N_16890);
nor U22993 (N_22993,N_13315,N_16225);
or U22994 (N_22994,N_12647,N_15765);
nand U22995 (N_22995,N_18155,N_14609);
nand U22996 (N_22996,N_16876,N_14603);
nor U22997 (N_22997,N_15004,N_16358);
nand U22998 (N_22998,N_18475,N_17364);
xnor U22999 (N_22999,N_15520,N_13344);
nand U23000 (N_23000,N_15798,N_16899);
nand U23001 (N_23001,N_12772,N_14576);
nand U23002 (N_23002,N_17852,N_14896);
nand U23003 (N_23003,N_16325,N_17924);
nand U23004 (N_23004,N_14985,N_12732);
xnor U23005 (N_23005,N_16535,N_18600);
and U23006 (N_23006,N_14681,N_16507);
xnor U23007 (N_23007,N_17329,N_18450);
nand U23008 (N_23008,N_13707,N_18400);
nor U23009 (N_23009,N_13999,N_13470);
and U23010 (N_23010,N_14502,N_18642);
nand U23011 (N_23011,N_13042,N_18494);
or U23012 (N_23012,N_18331,N_17678);
nand U23013 (N_23013,N_12925,N_17730);
or U23014 (N_23014,N_15346,N_17162);
and U23015 (N_23015,N_15326,N_18416);
nand U23016 (N_23016,N_14408,N_14136);
xnor U23017 (N_23017,N_17655,N_14961);
or U23018 (N_23018,N_17158,N_15020);
and U23019 (N_23019,N_15438,N_17225);
nor U23020 (N_23020,N_14670,N_17637);
nor U23021 (N_23021,N_17795,N_14587);
and U23022 (N_23022,N_17283,N_17944);
nor U23023 (N_23023,N_17953,N_13827);
nand U23024 (N_23024,N_12508,N_18699);
nor U23025 (N_23025,N_13551,N_15826);
nor U23026 (N_23026,N_15882,N_13738);
xnor U23027 (N_23027,N_17652,N_16910);
or U23028 (N_23028,N_18481,N_13972);
or U23029 (N_23029,N_14450,N_18030);
or U23030 (N_23030,N_15387,N_16123);
xor U23031 (N_23031,N_12577,N_13694);
and U23032 (N_23032,N_13813,N_18672);
or U23033 (N_23033,N_17366,N_17630);
nor U23034 (N_23034,N_16435,N_16064);
and U23035 (N_23035,N_18146,N_15665);
or U23036 (N_23036,N_13711,N_17590);
and U23037 (N_23037,N_15972,N_14988);
nand U23038 (N_23038,N_15869,N_14721);
nand U23039 (N_23039,N_12967,N_17461);
nor U23040 (N_23040,N_15938,N_16489);
nand U23041 (N_23041,N_13807,N_14342);
or U23042 (N_23042,N_18575,N_15547);
nand U23043 (N_23043,N_16035,N_13268);
or U23044 (N_23044,N_15006,N_15308);
nand U23045 (N_23045,N_13547,N_15797);
or U23046 (N_23046,N_16949,N_15937);
xnor U23047 (N_23047,N_18289,N_17110);
or U23048 (N_23048,N_17473,N_18368);
and U23049 (N_23049,N_17659,N_15001);
xnor U23050 (N_23050,N_13419,N_18516);
or U23051 (N_23051,N_14332,N_17739);
or U23052 (N_23052,N_13676,N_14216);
nand U23053 (N_23053,N_13057,N_16818);
nor U23054 (N_23054,N_17425,N_18568);
and U23055 (N_23055,N_17873,N_15772);
or U23056 (N_23056,N_13309,N_12641);
or U23057 (N_23057,N_16007,N_18241);
nand U23058 (N_23058,N_17551,N_15033);
xnor U23059 (N_23059,N_13805,N_13303);
nand U23060 (N_23060,N_18105,N_16034);
and U23061 (N_23061,N_13760,N_16478);
and U23062 (N_23062,N_16470,N_15898);
or U23063 (N_23063,N_12692,N_16487);
or U23064 (N_23064,N_16177,N_15855);
and U23065 (N_23065,N_13741,N_17045);
or U23066 (N_23066,N_17484,N_12903);
nor U23067 (N_23067,N_13409,N_14581);
nand U23068 (N_23068,N_17184,N_13637);
nor U23069 (N_23069,N_17161,N_15663);
xor U23070 (N_23070,N_17892,N_14058);
and U23071 (N_23071,N_16508,N_13300);
nand U23072 (N_23072,N_12600,N_12695);
nand U23073 (N_23073,N_13478,N_18051);
or U23074 (N_23074,N_15066,N_14909);
nand U23075 (N_23075,N_17092,N_17490);
or U23076 (N_23076,N_18172,N_14322);
nand U23077 (N_23077,N_14468,N_13225);
nand U23078 (N_23078,N_18674,N_14380);
and U23079 (N_23079,N_16123,N_17213);
or U23080 (N_23080,N_14383,N_18088);
or U23081 (N_23081,N_14088,N_15288);
nor U23082 (N_23082,N_17899,N_18121);
nand U23083 (N_23083,N_14226,N_16926);
or U23084 (N_23084,N_17033,N_13064);
and U23085 (N_23085,N_12510,N_17642);
or U23086 (N_23086,N_14734,N_16664);
xnor U23087 (N_23087,N_15461,N_14440);
nand U23088 (N_23088,N_13704,N_14343);
nand U23089 (N_23089,N_16662,N_18472);
or U23090 (N_23090,N_17974,N_17042);
nand U23091 (N_23091,N_15555,N_13847);
nand U23092 (N_23092,N_13026,N_17128);
nor U23093 (N_23093,N_14402,N_17004);
xnor U23094 (N_23094,N_14550,N_15509);
nand U23095 (N_23095,N_14781,N_14579);
nor U23096 (N_23096,N_15671,N_15915);
nor U23097 (N_23097,N_15226,N_14421);
and U23098 (N_23098,N_15417,N_12896);
nand U23099 (N_23099,N_17594,N_16065);
and U23100 (N_23100,N_17205,N_14845);
or U23101 (N_23101,N_15464,N_14442);
and U23102 (N_23102,N_14060,N_13018);
nor U23103 (N_23103,N_14869,N_14656);
nand U23104 (N_23104,N_17846,N_16159);
nor U23105 (N_23105,N_13858,N_15659);
nor U23106 (N_23106,N_17012,N_17321);
nor U23107 (N_23107,N_16278,N_14240);
or U23108 (N_23108,N_16124,N_15698);
nand U23109 (N_23109,N_13013,N_13508);
nand U23110 (N_23110,N_13428,N_16027);
and U23111 (N_23111,N_13725,N_18671);
xor U23112 (N_23112,N_14599,N_18720);
nand U23113 (N_23113,N_16847,N_14221);
nand U23114 (N_23114,N_16271,N_13835);
nor U23115 (N_23115,N_16624,N_12637);
and U23116 (N_23116,N_16731,N_14393);
and U23117 (N_23117,N_16961,N_12615);
nor U23118 (N_23118,N_15725,N_14080);
nand U23119 (N_23119,N_13172,N_15070);
nor U23120 (N_23120,N_15518,N_14836);
xnor U23121 (N_23121,N_12679,N_18366);
or U23122 (N_23122,N_12692,N_14978);
nor U23123 (N_23123,N_14195,N_18737);
and U23124 (N_23124,N_14081,N_14619);
or U23125 (N_23125,N_16890,N_14004);
xnor U23126 (N_23126,N_17441,N_13192);
and U23127 (N_23127,N_16040,N_17435);
nand U23128 (N_23128,N_13255,N_15328);
nor U23129 (N_23129,N_16430,N_13758);
or U23130 (N_23130,N_18219,N_16969);
nor U23131 (N_23131,N_14548,N_14726);
nand U23132 (N_23132,N_13569,N_17867);
nand U23133 (N_23133,N_16408,N_13324);
and U23134 (N_23134,N_15786,N_17134);
nor U23135 (N_23135,N_13186,N_16621);
nor U23136 (N_23136,N_13002,N_14795);
nor U23137 (N_23137,N_17034,N_18280);
and U23138 (N_23138,N_13477,N_17657);
nor U23139 (N_23139,N_18028,N_13947);
and U23140 (N_23140,N_14314,N_16427);
and U23141 (N_23141,N_13574,N_16375);
or U23142 (N_23142,N_13665,N_17369);
and U23143 (N_23143,N_15453,N_17815);
nand U23144 (N_23144,N_18730,N_12777);
nand U23145 (N_23145,N_13956,N_16814);
and U23146 (N_23146,N_17539,N_13008);
nor U23147 (N_23147,N_13732,N_15612);
nand U23148 (N_23148,N_17345,N_18208);
nor U23149 (N_23149,N_16817,N_18617);
or U23150 (N_23150,N_17623,N_17171);
nor U23151 (N_23151,N_16572,N_13293);
nor U23152 (N_23152,N_14834,N_15678);
nand U23153 (N_23153,N_15591,N_15966);
nor U23154 (N_23154,N_12508,N_18636);
or U23155 (N_23155,N_18713,N_12514);
or U23156 (N_23156,N_13970,N_13575);
or U23157 (N_23157,N_12573,N_16972);
nand U23158 (N_23158,N_17836,N_17757);
or U23159 (N_23159,N_15018,N_16452);
and U23160 (N_23160,N_18352,N_16329);
nor U23161 (N_23161,N_15178,N_15036);
and U23162 (N_23162,N_18403,N_12568);
nand U23163 (N_23163,N_14293,N_16866);
and U23164 (N_23164,N_14930,N_17851);
nor U23165 (N_23165,N_18487,N_17462);
or U23166 (N_23166,N_18090,N_16826);
nor U23167 (N_23167,N_16800,N_13284);
and U23168 (N_23168,N_18564,N_12777);
or U23169 (N_23169,N_16960,N_13556);
nand U23170 (N_23170,N_14264,N_14999);
and U23171 (N_23171,N_12590,N_12657);
nand U23172 (N_23172,N_18264,N_13179);
and U23173 (N_23173,N_14041,N_16777);
nor U23174 (N_23174,N_17478,N_14351);
and U23175 (N_23175,N_13276,N_17110);
nand U23176 (N_23176,N_15624,N_16843);
nand U23177 (N_23177,N_13086,N_18066);
and U23178 (N_23178,N_12947,N_17531);
nand U23179 (N_23179,N_17243,N_17542);
nor U23180 (N_23180,N_14087,N_17213);
nor U23181 (N_23181,N_18738,N_16918);
nand U23182 (N_23182,N_17976,N_14735);
and U23183 (N_23183,N_13129,N_17205);
and U23184 (N_23184,N_14090,N_15214);
nor U23185 (N_23185,N_14796,N_12708);
nor U23186 (N_23186,N_16465,N_15534);
xnor U23187 (N_23187,N_17368,N_18515);
xnor U23188 (N_23188,N_14025,N_14973);
and U23189 (N_23189,N_14532,N_14451);
nor U23190 (N_23190,N_16481,N_14215);
and U23191 (N_23191,N_13597,N_15295);
and U23192 (N_23192,N_17644,N_13345);
nand U23193 (N_23193,N_13333,N_18339);
or U23194 (N_23194,N_18120,N_13470);
nand U23195 (N_23195,N_15398,N_14274);
nand U23196 (N_23196,N_15898,N_18598);
and U23197 (N_23197,N_13072,N_18396);
nor U23198 (N_23198,N_13135,N_12617);
and U23199 (N_23199,N_18533,N_13443);
or U23200 (N_23200,N_14021,N_14905);
or U23201 (N_23201,N_13347,N_14731);
or U23202 (N_23202,N_17850,N_17345);
nor U23203 (N_23203,N_16946,N_12739);
or U23204 (N_23204,N_17656,N_14103);
nand U23205 (N_23205,N_15648,N_15970);
xnor U23206 (N_23206,N_13780,N_16453);
or U23207 (N_23207,N_15400,N_15580);
xor U23208 (N_23208,N_16567,N_16541);
or U23209 (N_23209,N_12840,N_15913);
or U23210 (N_23210,N_18096,N_12762);
nor U23211 (N_23211,N_18226,N_17970);
nor U23212 (N_23212,N_12676,N_14183);
or U23213 (N_23213,N_14379,N_16176);
xnor U23214 (N_23214,N_18035,N_17727);
nand U23215 (N_23215,N_18725,N_17811);
nor U23216 (N_23216,N_13592,N_16222);
and U23217 (N_23217,N_18115,N_16076);
nor U23218 (N_23218,N_17412,N_17791);
nor U23219 (N_23219,N_18202,N_16890);
xnor U23220 (N_23220,N_17152,N_16643);
and U23221 (N_23221,N_15448,N_17452);
nor U23222 (N_23222,N_12868,N_13178);
xor U23223 (N_23223,N_16237,N_18206);
and U23224 (N_23224,N_15253,N_14887);
nand U23225 (N_23225,N_13089,N_17153);
or U23226 (N_23226,N_18389,N_16669);
and U23227 (N_23227,N_15895,N_13954);
and U23228 (N_23228,N_15849,N_17717);
xnor U23229 (N_23229,N_12615,N_16166);
nand U23230 (N_23230,N_12705,N_17149);
or U23231 (N_23231,N_14729,N_15127);
or U23232 (N_23232,N_13801,N_17100);
and U23233 (N_23233,N_13864,N_18631);
nor U23234 (N_23234,N_16863,N_13637);
nor U23235 (N_23235,N_13785,N_16791);
nand U23236 (N_23236,N_14736,N_16598);
and U23237 (N_23237,N_13917,N_16415);
or U23238 (N_23238,N_18153,N_15096);
nand U23239 (N_23239,N_13447,N_15570);
nand U23240 (N_23240,N_15584,N_15053);
nand U23241 (N_23241,N_14204,N_13794);
and U23242 (N_23242,N_17403,N_15717);
nand U23243 (N_23243,N_16263,N_13473);
nor U23244 (N_23244,N_14072,N_18698);
or U23245 (N_23245,N_17342,N_15960);
xnor U23246 (N_23246,N_16262,N_16416);
or U23247 (N_23247,N_17430,N_17219);
xor U23248 (N_23248,N_16370,N_18616);
xor U23249 (N_23249,N_12800,N_16858);
nor U23250 (N_23250,N_18334,N_16582);
or U23251 (N_23251,N_14925,N_18732);
nand U23252 (N_23252,N_15475,N_15723);
nor U23253 (N_23253,N_15979,N_17620);
nand U23254 (N_23254,N_16520,N_18671);
and U23255 (N_23255,N_15230,N_12942);
nor U23256 (N_23256,N_13248,N_15712);
and U23257 (N_23257,N_15315,N_16598);
or U23258 (N_23258,N_17191,N_15594);
and U23259 (N_23259,N_18537,N_13923);
nand U23260 (N_23260,N_12995,N_14669);
and U23261 (N_23261,N_16508,N_18254);
or U23262 (N_23262,N_18655,N_16069);
nor U23263 (N_23263,N_14787,N_14821);
nor U23264 (N_23264,N_17927,N_12853);
or U23265 (N_23265,N_13857,N_16488);
nor U23266 (N_23266,N_14110,N_17939);
nand U23267 (N_23267,N_17756,N_13908);
nand U23268 (N_23268,N_14241,N_12973);
nor U23269 (N_23269,N_15363,N_17207);
or U23270 (N_23270,N_15895,N_13142);
and U23271 (N_23271,N_15667,N_16541);
nor U23272 (N_23272,N_12606,N_18217);
or U23273 (N_23273,N_16370,N_13911);
and U23274 (N_23274,N_18164,N_13761);
or U23275 (N_23275,N_14932,N_18541);
nor U23276 (N_23276,N_18013,N_18724);
xnor U23277 (N_23277,N_17406,N_14848);
or U23278 (N_23278,N_15997,N_18674);
nand U23279 (N_23279,N_12693,N_14789);
or U23280 (N_23280,N_13441,N_16127);
nor U23281 (N_23281,N_13587,N_17916);
nand U23282 (N_23282,N_16624,N_17517);
nand U23283 (N_23283,N_17344,N_16450);
nor U23284 (N_23284,N_15708,N_13448);
nand U23285 (N_23285,N_13670,N_18292);
nor U23286 (N_23286,N_17342,N_16873);
and U23287 (N_23287,N_17871,N_17726);
or U23288 (N_23288,N_15731,N_18167);
or U23289 (N_23289,N_13426,N_17282);
nor U23290 (N_23290,N_16893,N_15644);
xor U23291 (N_23291,N_17368,N_12559);
xnor U23292 (N_23292,N_15742,N_16295);
or U23293 (N_23293,N_13972,N_15756);
nand U23294 (N_23294,N_15123,N_16092);
nor U23295 (N_23295,N_17324,N_14737);
or U23296 (N_23296,N_17442,N_17632);
or U23297 (N_23297,N_13988,N_14920);
nand U23298 (N_23298,N_18053,N_15113);
or U23299 (N_23299,N_15815,N_15024);
and U23300 (N_23300,N_14139,N_15815);
or U23301 (N_23301,N_13098,N_13379);
and U23302 (N_23302,N_14427,N_18598);
nand U23303 (N_23303,N_13540,N_18419);
or U23304 (N_23304,N_17123,N_16703);
and U23305 (N_23305,N_15247,N_17530);
nand U23306 (N_23306,N_14623,N_16089);
or U23307 (N_23307,N_13048,N_15372);
nor U23308 (N_23308,N_12852,N_16239);
or U23309 (N_23309,N_16582,N_13080);
nor U23310 (N_23310,N_15962,N_15982);
and U23311 (N_23311,N_17325,N_15553);
nor U23312 (N_23312,N_16956,N_18064);
and U23313 (N_23313,N_14692,N_17884);
nand U23314 (N_23314,N_16564,N_13124);
nor U23315 (N_23315,N_13483,N_17124);
and U23316 (N_23316,N_16907,N_15785);
or U23317 (N_23317,N_12766,N_15567);
nor U23318 (N_23318,N_14993,N_13787);
nand U23319 (N_23319,N_14166,N_17026);
nand U23320 (N_23320,N_15714,N_18377);
nand U23321 (N_23321,N_14217,N_12752);
and U23322 (N_23322,N_13065,N_17818);
and U23323 (N_23323,N_13001,N_13724);
nand U23324 (N_23324,N_14450,N_13447);
nand U23325 (N_23325,N_15847,N_13095);
or U23326 (N_23326,N_16747,N_17166);
nand U23327 (N_23327,N_15540,N_13320);
and U23328 (N_23328,N_18729,N_17660);
nor U23329 (N_23329,N_18253,N_16537);
and U23330 (N_23330,N_16928,N_17725);
nor U23331 (N_23331,N_15599,N_16833);
nor U23332 (N_23332,N_16479,N_14904);
xnor U23333 (N_23333,N_18621,N_16742);
and U23334 (N_23334,N_14445,N_17316);
nor U23335 (N_23335,N_12959,N_17477);
nand U23336 (N_23336,N_13916,N_15286);
nand U23337 (N_23337,N_15153,N_12502);
nor U23338 (N_23338,N_18631,N_12774);
xor U23339 (N_23339,N_14456,N_15527);
and U23340 (N_23340,N_13384,N_12892);
nand U23341 (N_23341,N_17217,N_18687);
or U23342 (N_23342,N_12833,N_15368);
nand U23343 (N_23343,N_16526,N_14539);
or U23344 (N_23344,N_16581,N_12851);
or U23345 (N_23345,N_13089,N_15183);
nand U23346 (N_23346,N_13992,N_18749);
nand U23347 (N_23347,N_18549,N_12574);
or U23348 (N_23348,N_16759,N_14514);
and U23349 (N_23349,N_16560,N_15796);
or U23350 (N_23350,N_13472,N_13064);
nor U23351 (N_23351,N_17642,N_15049);
nand U23352 (N_23352,N_13360,N_15488);
and U23353 (N_23353,N_17454,N_16031);
nand U23354 (N_23354,N_13607,N_12628);
nor U23355 (N_23355,N_17773,N_18740);
nand U23356 (N_23356,N_16883,N_12612);
nand U23357 (N_23357,N_16154,N_15596);
xnor U23358 (N_23358,N_18495,N_13762);
nand U23359 (N_23359,N_14405,N_18608);
and U23360 (N_23360,N_14107,N_12927);
nand U23361 (N_23361,N_14672,N_13257);
nand U23362 (N_23362,N_15650,N_17835);
or U23363 (N_23363,N_14784,N_15896);
or U23364 (N_23364,N_18136,N_14062);
nand U23365 (N_23365,N_15853,N_16050);
and U23366 (N_23366,N_13392,N_15373);
nand U23367 (N_23367,N_18681,N_16393);
nor U23368 (N_23368,N_14274,N_13166);
nand U23369 (N_23369,N_15172,N_15037);
nor U23370 (N_23370,N_14229,N_15662);
or U23371 (N_23371,N_16799,N_16324);
nand U23372 (N_23372,N_14062,N_14735);
nand U23373 (N_23373,N_13142,N_16310);
nand U23374 (N_23374,N_18325,N_18045);
and U23375 (N_23375,N_14714,N_13751);
or U23376 (N_23376,N_13294,N_15787);
and U23377 (N_23377,N_17279,N_13738);
nand U23378 (N_23378,N_17052,N_16280);
nand U23379 (N_23379,N_18459,N_14790);
or U23380 (N_23380,N_12661,N_14593);
xnor U23381 (N_23381,N_13157,N_17476);
or U23382 (N_23382,N_15343,N_16412);
or U23383 (N_23383,N_17555,N_14634);
nor U23384 (N_23384,N_17818,N_14983);
nor U23385 (N_23385,N_17742,N_18636);
nor U23386 (N_23386,N_14629,N_17749);
and U23387 (N_23387,N_15108,N_17308);
and U23388 (N_23388,N_18602,N_17811);
nand U23389 (N_23389,N_12751,N_15509);
and U23390 (N_23390,N_14262,N_17267);
nand U23391 (N_23391,N_15585,N_15382);
nor U23392 (N_23392,N_18500,N_13628);
and U23393 (N_23393,N_17701,N_13989);
nor U23394 (N_23394,N_17219,N_17738);
and U23395 (N_23395,N_14896,N_14455);
or U23396 (N_23396,N_18389,N_12591);
nand U23397 (N_23397,N_17198,N_14054);
and U23398 (N_23398,N_17118,N_15220);
or U23399 (N_23399,N_18313,N_16262);
nand U23400 (N_23400,N_13153,N_17670);
or U23401 (N_23401,N_13861,N_18155);
or U23402 (N_23402,N_13664,N_15975);
nor U23403 (N_23403,N_15448,N_15936);
nand U23404 (N_23404,N_16409,N_13833);
and U23405 (N_23405,N_14564,N_13650);
and U23406 (N_23406,N_12767,N_13299);
nand U23407 (N_23407,N_16030,N_15226);
nor U23408 (N_23408,N_18658,N_15444);
or U23409 (N_23409,N_14531,N_17440);
or U23410 (N_23410,N_16010,N_13474);
or U23411 (N_23411,N_14056,N_18261);
or U23412 (N_23412,N_15455,N_13770);
and U23413 (N_23413,N_15671,N_15040);
and U23414 (N_23414,N_12848,N_16734);
and U23415 (N_23415,N_16650,N_14702);
or U23416 (N_23416,N_18256,N_15329);
or U23417 (N_23417,N_13144,N_13282);
nand U23418 (N_23418,N_12708,N_15609);
nand U23419 (N_23419,N_12835,N_17863);
nand U23420 (N_23420,N_14683,N_15593);
nor U23421 (N_23421,N_16606,N_15936);
xor U23422 (N_23422,N_12948,N_14079);
nor U23423 (N_23423,N_17314,N_17379);
or U23424 (N_23424,N_17268,N_14117);
nor U23425 (N_23425,N_14819,N_15304);
or U23426 (N_23426,N_15966,N_12736);
or U23427 (N_23427,N_14919,N_14290);
nor U23428 (N_23428,N_16128,N_13660);
nand U23429 (N_23429,N_16633,N_17391);
nand U23430 (N_23430,N_13213,N_15849);
nand U23431 (N_23431,N_14129,N_16747);
nand U23432 (N_23432,N_12593,N_15884);
and U23433 (N_23433,N_16224,N_18697);
nor U23434 (N_23434,N_16187,N_13095);
nor U23435 (N_23435,N_13348,N_15583);
and U23436 (N_23436,N_15798,N_15196);
nand U23437 (N_23437,N_15968,N_14838);
and U23438 (N_23438,N_16049,N_15345);
nand U23439 (N_23439,N_13022,N_13196);
or U23440 (N_23440,N_15850,N_17839);
or U23441 (N_23441,N_17200,N_14432);
nand U23442 (N_23442,N_15525,N_17815);
and U23443 (N_23443,N_18164,N_14306);
nand U23444 (N_23444,N_17342,N_14993);
or U23445 (N_23445,N_16350,N_13299);
or U23446 (N_23446,N_15779,N_16160);
or U23447 (N_23447,N_12649,N_17809);
or U23448 (N_23448,N_14528,N_17548);
or U23449 (N_23449,N_15331,N_18031);
or U23450 (N_23450,N_14829,N_16201);
nand U23451 (N_23451,N_16650,N_18273);
and U23452 (N_23452,N_13203,N_15836);
or U23453 (N_23453,N_18657,N_17747);
xnor U23454 (N_23454,N_13591,N_15308);
nor U23455 (N_23455,N_17632,N_17848);
or U23456 (N_23456,N_17392,N_15876);
and U23457 (N_23457,N_12927,N_12899);
nand U23458 (N_23458,N_16765,N_13448);
and U23459 (N_23459,N_12713,N_17406);
nand U23460 (N_23460,N_18225,N_15412);
nand U23461 (N_23461,N_14801,N_13513);
nand U23462 (N_23462,N_17345,N_17386);
nand U23463 (N_23463,N_14709,N_15668);
or U23464 (N_23464,N_15448,N_13451);
nand U23465 (N_23465,N_12751,N_16873);
or U23466 (N_23466,N_16967,N_13148);
nor U23467 (N_23467,N_17216,N_13047);
and U23468 (N_23468,N_17624,N_14226);
xnor U23469 (N_23469,N_15796,N_13178);
nor U23470 (N_23470,N_14806,N_18206);
nand U23471 (N_23471,N_13306,N_17833);
nand U23472 (N_23472,N_17476,N_16674);
and U23473 (N_23473,N_15384,N_16807);
xor U23474 (N_23474,N_17133,N_17939);
or U23475 (N_23475,N_16582,N_13403);
and U23476 (N_23476,N_17239,N_13976);
or U23477 (N_23477,N_13010,N_17032);
or U23478 (N_23478,N_12711,N_15120);
nand U23479 (N_23479,N_17904,N_12860);
nand U23480 (N_23480,N_14732,N_16924);
xor U23481 (N_23481,N_16830,N_16952);
nand U23482 (N_23482,N_16669,N_15663);
nand U23483 (N_23483,N_17551,N_18458);
or U23484 (N_23484,N_14334,N_18523);
and U23485 (N_23485,N_14922,N_16419);
nand U23486 (N_23486,N_15158,N_17238);
nand U23487 (N_23487,N_14506,N_13087);
nand U23488 (N_23488,N_14692,N_15984);
or U23489 (N_23489,N_12767,N_17253);
or U23490 (N_23490,N_15834,N_12555);
and U23491 (N_23491,N_18326,N_13535);
xnor U23492 (N_23492,N_12535,N_17852);
nand U23493 (N_23493,N_14905,N_18163);
or U23494 (N_23494,N_16265,N_13123);
nor U23495 (N_23495,N_14971,N_12908);
and U23496 (N_23496,N_14216,N_13605);
or U23497 (N_23497,N_16664,N_17969);
and U23498 (N_23498,N_13084,N_17988);
nor U23499 (N_23499,N_13787,N_16688);
nand U23500 (N_23500,N_17891,N_18493);
nor U23501 (N_23501,N_16020,N_16361);
and U23502 (N_23502,N_14626,N_12692);
xnor U23503 (N_23503,N_15714,N_13883);
nand U23504 (N_23504,N_15583,N_14037);
nand U23505 (N_23505,N_15965,N_16930);
nand U23506 (N_23506,N_14545,N_16128);
and U23507 (N_23507,N_15392,N_12524);
or U23508 (N_23508,N_15561,N_16750);
and U23509 (N_23509,N_14575,N_16497);
and U23510 (N_23510,N_14044,N_15391);
or U23511 (N_23511,N_13612,N_14330);
nor U23512 (N_23512,N_15118,N_17457);
nor U23513 (N_23513,N_16052,N_18719);
nor U23514 (N_23514,N_15166,N_13945);
or U23515 (N_23515,N_14591,N_14262);
or U23516 (N_23516,N_13797,N_18429);
xnor U23517 (N_23517,N_15621,N_15466);
and U23518 (N_23518,N_16215,N_13011);
and U23519 (N_23519,N_16804,N_13176);
and U23520 (N_23520,N_17243,N_12569);
nor U23521 (N_23521,N_12747,N_13713);
and U23522 (N_23522,N_17620,N_14927);
or U23523 (N_23523,N_14675,N_17493);
nor U23524 (N_23524,N_14985,N_16566);
or U23525 (N_23525,N_15056,N_18686);
and U23526 (N_23526,N_14252,N_14583);
nand U23527 (N_23527,N_13650,N_18470);
and U23528 (N_23528,N_17058,N_16294);
or U23529 (N_23529,N_14296,N_13865);
nand U23530 (N_23530,N_12975,N_17848);
and U23531 (N_23531,N_15636,N_17034);
or U23532 (N_23532,N_15926,N_14060);
and U23533 (N_23533,N_18080,N_17844);
or U23534 (N_23534,N_15836,N_17753);
nor U23535 (N_23535,N_17287,N_15917);
and U23536 (N_23536,N_14693,N_12622);
nand U23537 (N_23537,N_15379,N_13541);
nand U23538 (N_23538,N_18725,N_14381);
and U23539 (N_23539,N_13769,N_15435);
or U23540 (N_23540,N_15399,N_13295);
nor U23541 (N_23541,N_13639,N_15188);
nor U23542 (N_23542,N_16610,N_15135);
and U23543 (N_23543,N_13492,N_13572);
nand U23544 (N_23544,N_13359,N_14141);
and U23545 (N_23545,N_18165,N_18132);
and U23546 (N_23546,N_18614,N_16680);
or U23547 (N_23547,N_14985,N_16254);
nor U23548 (N_23548,N_14527,N_18016);
nor U23549 (N_23549,N_15814,N_18396);
nor U23550 (N_23550,N_16394,N_16038);
or U23551 (N_23551,N_18679,N_15071);
and U23552 (N_23552,N_13145,N_16431);
and U23553 (N_23553,N_13655,N_18388);
or U23554 (N_23554,N_16227,N_13740);
nor U23555 (N_23555,N_15027,N_12590);
nor U23556 (N_23556,N_13379,N_18573);
nand U23557 (N_23557,N_18510,N_17569);
and U23558 (N_23558,N_14926,N_13406);
nor U23559 (N_23559,N_15750,N_13804);
nand U23560 (N_23560,N_17363,N_16131);
nand U23561 (N_23561,N_13475,N_16483);
and U23562 (N_23562,N_16295,N_14160);
and U23563 (N_23563,N_14594,N_17490);
xnor U23564 (N_23564,N_18138,N_18632);
nor U23565 (N_23565,N_12520,N_14861);
nand U23566 (N_23566,N_17282,N_16793);
or U23567 (N_23567,N_14643,N_17617);
or U23568 (N_23568,N_17087,N_15630);
nor U23569 (N_23569,N_14388,N_16663);
or U23570 (N_23570,N_14785,N_13867);
nor U23571 (N_23571,N_16720,N_18327);
xor U23572 (N_23572,N_18480,N_18713);
or U23573 (N_23573,N_16712,N_16259);
xnor U23574 (N_23574,N_15832,N_18404);
nor U23575 (N_23575,N_13574,N_14438);
nor U23576 (N_23576,N_18129,N_16746);
and U23577 (N_23577,N_14077,N_13490);
and U23578 (N_23578,N_17997,N_17456);
or U23579 (N_23579,N_17835,N_17895);
or U23580 (N_23580,N_13649,N_17009);
xor U23581 (N_23581,N_15659,N_17143);
and U23582 (N_23582,N_15028,N_13250);
nor U23583 (N_23583,N_14030,N_15817);
nor U23584 (N_23584,N_14226,N_15605);
nand U23585 (N_23585,N_15622,N_14952);
nand U23586 (N_23586,N_15931,N_17453);
nand U23587 (N_23587,N_13881,N_15135);
nand U23588 (N_23588,N_16386,N_14771);
nand U23589 (N_23589,N_15193,N_18056);
or U23590 (N_23590,N_18732,N_13521);
nand U23591 (N_23591,N_17644,N_18064);
nor U23592 (N_23592,N_18540,N_14825);
nand U23593 (N_23593,N_17535,N_13753);
and U23594 (N_23594,N_17051,N_17189);
xnor U23595 (N_23595,N_13122,N_18404);
xor U23596 (N_23596,N_15200,N_18161);
or U23597 (N_23597,N_16648,N_18087);
and U23598 (N_23598,N_14693,N_16927);
nor U23599 (N_23599,N_13558,N_15380);
and U23600 (N_23600,N_17052,N_17452);
or U23601 (N_23601,N_14074,N_14130);
and U23602 (N_23602,N_18537,N_13754);
nand U23603 (N_23603,N_18648,N_14317);
and U23604 (N_23604,N_15477,N_15178);
nor U23605 (N_23605,N_13996,N_16044);
and U23606 (N_23606,N_13404,N_17599);
xor U23607 (N_23607,N_14365,N_15957);
nor U23608 (N_23608,N_15075,N_18181);
or U23609 (N_23609,N_18012,N_17973);
or U23610 (N_23610,N_13607,N_18312);
nor U23611 (N_23611,N_16155,N_17061);
or U23612 (N_23612,N_14252,N_14501);
or U23613 (N_23613,N_16208,N_17993);
and U23614 (N_23614,N_13601,N_17028);
and U23615 (N_23615,N_18194,N_13763);
or U23616 (N_23616,N_17972,N_15107);
and U23617 (N_23617,N_14205,N_15282);
nand U23618 (N_23618,N_17805,N_17652);
and U23619 (N_23619,N_16492,N_17215);
or U23620 (N_23620,N_15098,N_16565);
or U23621 (N_23621,N_12804,N_13853);
or U23622 (N_23622,N_18327,N_17229);
nand U23623 (N_23623,N_15945,N_13530);
or U23624 (N_23624,N_12875,N_16831);
or U23625 (N_23625,N_17915,N_12671);
nor U23626 (N_23626,N_15925,N_18056);
xor U23627 (N_23627,N_17877,N_14106);
nor U23628 (N_23628,N_15277,N_12994);
nand U23629 (N_23629,N_16149,N_16570);
or U23630 (N_23630,N_13066,N_16492);
nand U23631 (N_23631,N_14648,N_14223);
nor U23632 (N_23632,N_14342,N_16443);
nand U23633 (N_23633,N_16975,N_16250);
and U23634 (N_23634,N_15666,N_14459);
nand U23635 (N_23635,N_15828,N_14153);
or U23636 (N_23636,N_16691,N_13861);
or U23637 (N_23637,N_18313,N_14143);
or U23638 (N_23638,N_12922,N_16013);
or U23639 (N_23639,N_14742,N_15977);
nand U23640 (N_23640,N_15131,N_15775);
nor U23641 (N_23641,N_14180,N_14544);
nand U23642 (N_23642,N_18427,N_15684);
nand U23643 (N_23643,N_16263,N_17990);
nand U23644 (N_23644,N_12602,N_15856);
xnor U23645 (N_23645,N_17271,N_16705);
xor U23646 (N_23646,N_18157,N_12799);
and U23647 (N_23647,N_17828,N_15825);
nor U23648 (N_23648,N_16177,N_17543);
or U23649 (N_23649,N_16335,N_13322);
or U23650 (N_23650,N_14951,N_18195);
nor U23651 (N_23651,N_17779,N_14200);
and U23652 (N_23652,N_16900,N_15795);
nor U23653 (N_23653,N_14067,N_14721);
or U23654 (N_23654,N_15460,N_13781);
nor U23655 (N_23655,N_12930,N_15718);
and U23656 (N_23656,N_16810,N_17656);
nand U23657 (N_23657,N_16824,N_15901);
nand U23658 (N_23658,N_15607,N_14582);
or U23659 (N_23659,N_18114,N_14306);
nor U23660 (N_23660,N_16505,N_14988);
nand U23661 (N_23661,N_18664,N_14307);
or U23662 (N_23662,N_14495,N_15671);
nand U23663 (N_23663,N_17678,N_16571);
and U23664 (N_23664,N_14856,N_15363);
or U23665 (N_23665,N_18358,N_15415);
nand U23666 (N_23666,N_17028,N_13047);
nor U23667 (N_23667,N_15703,N_17094);
nand U23668 (N_23668,N_17973,N_16827);
nor U23669 (N_23669,N_18266,N_18102);
nor U23670 (N_23670,N_17252,N_15311);
or U23671 (N_23671,N_17578,N_18733);
and U23672 (N_23672,N_18614,N_12843);
xor U23673 (N_23673,N_14804,N_15694);
nand U23674 (N_23674,N_15969,N_17576);
or U23675 (N_23675,N_15225,N_14583);
and U23676 (N_23676,N_16144,N_17779);
nand U23677 (N_23677,N_18292,N_18084);
nand U23678 (N_23678,N_15678,N_16428);
nand U23679 (N_23679,N_13390,N_17444);
or U23680 (N_23680,N_16555,N_13196);
and U23681 (N_23681,N_17295,N_17035);
and U23682 (N_23682,N_16552,N_17758);
nor U23683 (N_23683,N_14697,N_16218);
or U23684 (N_23684,N_14919,N_12877);
or U23685 (N_23685,N_12783,N_15533);
and U23686 (N_23686,N_12934,N_16948);
and U23687 (N_23687,N_16614,N_14152);
or U23688 (N_23688,N_13427,N_15267);
or U23689 (N_23689,N_14530,N_18094);
or U23690 (N_23690,N_18177,N_14451);
nor U23691 (N_23691,N_16370,N_14805);
nor U23692 (N_23692,N_17936,N_14304);
or U23693 (N_23693,N_12984,N_13393);
nor U23694 (N_23694,N_16024,N_17473);
and U23695 (N_23695,N_17651,N_15906);
nor U23696 (N_23696,N_13659,N_14812);
or U23697 (N_23697,N_13073,N_14002);
nor U23698 (N_23698,N_17470,N_14907);
and U23699 (N_23699,N_16250,N_13491);
nand U23700 (N_23700,N_13895,N_15802);
and U23701 (N_23701,N_14494,N_12943);
nand U23702 (N_23702,N_17093,N_18201);
nor U23703 (N_23703,N_13394,N_14600);
xnor U23704 (N_23704,N_18123,N_17360);
and U23705 (N_23705,N_16506,N_13009);
nor U23706 (N_23706,N_14281,N_17210);
and U23707 (N_23707,N_17526,N_13569);
nand U23708 (N_23708,N_17164,N_14569);
nor U23709 (N_23709,N_14877,N_14737);
nand U23710 (N_23710,N_18385,N_12964);
nor U23711 (N_23711,N_15766,N_14342);
and U23712 (N_23712,N_18538,N_17619);
nor U23713 (N_23713,N_17292,N_18389);
nor U23714 (N_23714,N_15487,N_12519);
nand U23715 (N_23715,N_16538,N_18576);
nand U23716 (N_23716,N_13099,N_16286);
nand U23717 (N_23717,N_14267,N_17501);
and U23718 (N_23718,N_15122,N_12741);
and U23719 (N_23719,N_17914,N_15844);
and U23720 (N_23720,N_12602,N_14888);
nor U23721 (N_23721,N_15068,N_18692);
or U23722 (N_23722,N_17354,N_17329);
and U23723 (N_23723,N_18693,N_15607);
or U23724 (N_23724,N_18492,N_17361);
nor U23725 (N_23725,N_13877,N_17368);
and U23726 (N_23726,N_15326,N_16012);
nand U23727 (N_23727,N_16116,N_13874);
nand U23728 (N_23728,N_12572,N_13579);
or U23729 (N_23729,N_12812,N_14456);
nor U23730 (N_23730,N_17507,N_17921);
and U23731 (N_23731,N_17632,N_15385);
or U23732 (N_23732,N_13427,N_13968);
and U23733 (N_23733,N_16114,N_17886);
xor U23734 (N_23734,N_17442,N_14963);
nand U23735 (N_23735,N_16636,N_15156);
nor U23736 (N_23736,N_16841,N_18253);
or U23737 (N_23737,N_15269,N_13125);
and U23738 (N_23738,N_17969,N_17017);
xor U23739 (N_23739,N_14256,N_14529);
and U23740 (N_23740,N_16671,N_14993);
and U23741 (N_23741,N_15855,N_12525);
nand U23742 (N_23742,N_13488,N_15052);
xnor U23743 (N_23743,N_14084,N_14716);
nand U23744 (N_23744,N_17369,N_16567);
nor U23745 (N_23745,N_15862,N_18127);
and U23746 (N_23746,N_16268,N_13605);
nor U23747 (N_23747,N_14331,N_14082);
xnor U23748 (N_23748,N_16796,N_14933);
nor U23749 (N_23749,N_15388,N_18200);
nor U23750 (N_23750,N_13221,N_14667);
nand U23751 (N_23751,N_17181,N_12987);
nand U23752 (N_23752,N_14420,N_13407);
and U23753 (N_23753,N_17723,N_18475);
nand U23754 (N_23754,N_15370,N_15978);
and U23755 (N_23755,N_16920,N_17070);
nand U23756 (N_23756,N_13158,N_12782);
or U23757 (N_23757,N_18186,N_16554);
nand U23758 (N_23758,N_16461,N_16735);
and U23759 (N_23759,N_13037,N_14374);
nand U23760 (N_23760,N_14740,N_15089);
nor U23761 (N_23761,N_18035,N_12930);
or U23762 (N_23762,N_14197,N_12951);
nand U23763 (N_23763,N_14090,N_15295);
and U23764 (N_23764,N_13674,N_18002);
nor U23765 (N_23765,N_14745,N_15961);
nand U23766 (N_23766,N_16516,N_16857);
nor U23767 (N_23767,N_14222,N_13339);
nand U23768 (N_23768,N_13745,N_14299);
or U23769 (N_23769,N_17271,N_15882);
and U23770 (N_23770,N_12632,N_15287);
xnor U23771 (N_23771,N_18362,N_18709);
nand U23772 (N_23772,N_15201,N_16027);
nor U23773 (N_23773,N_13986,N_17943);
or U23774 (N_23774,N_16046,N_15816);
xor U23775 (N_23775,N_14874,N_14650);
and U23776 (N_23776,N_18222,N_18536);
nand U23777 (N_23777,N_17100,N_12994);
or U23778 (N_23778,N_18107,N_17969);
nor U23779 (N_23779,N_14708,N_12831);
and U23780 (N_23780,N_15854,N_15734);
nor U23781 (N_23781,N_13591,N_16058);
and U23782 (N_23782,N_15046,N_16024);
or U23783 (N_23783,N_17521,N_16114);
and U23784 (N_23784,N_17567,N_14217);
or U23785 (N_23785,N_15079,N_12926);
nand U23786 (N_23786,N_18061,N_16574);
nand U23787 (N_23787,N_16621,N_16264);
and U23788 (N_23788,N_18623,N_17094);
or U23789 (N_23789,N_18380,N_14587);
and U23790 (N_23790,N_15194,N_15986);
xor U23791 (N_23791,N_15847,N_16202);
nand U23792 (N_23792,N_14279,N_16171);
and U23793 (N_23793,N_13782,N_16773);
and U23794 (N_23794,N_15921,N_17237);
xnor U23795 (N_23795,N_13549,N_18637);
nand U23796 (N_23796,N_12791,N_17725);
and U23797 (N_23797,N_14040,N_17578);
xnor U23798 (N_23798,N_15483,N_17891);
nor U23799 (N_23799,N_13570,N_12886);
nand U23800 (N_23800,N_15697,N_12636);
xor U23801 (N_23801,N_17724,N_13486);
nand U23802 (N_23802,N_13919,N_13359);
and U23803 (N_23803,N_12854,N_17714);
nor U23804 (N_23804,N_14121,N_17306);
or U23805 (N_23805,N_14055,N_15307);
or U23806 (N_23806,N_12738,N_14443);
nand U23807 (N_23807,N_12963,N_12875);
nand U23808 (N_23808,N_15510,N_16327);
or U23809 (N_23809,N_18384,N_13663);
or U23810 (N_23810,N_13354,N_16546);
or U23811 (N_23811,N_13576,N_18500);
nand U23812 (N_23812,N_16007,N_14137);
or U23813 (N_23813,N_18282,N_18631);
and U23814 (N_23814,N_17775,N_15423);
nor U23815 (N_23815,N_15321,N_18319);
and U23816 (N_23816,N_15744,N_18525);
and U23817 (N_23817,N_16908,N_15768);
or U23818 (N_23818,N_14538,N_13649);
and U23819 (N_23819,N_14828,N_15273);
or U23820 (N_23820,N_17291,N_13863);
and U23821 (N_23821,N_13354,N_14680);
nor U23822 (N_23822,N_16964,N_18707);
nor U23823 (N_23823,N_17632,N_18664);
and U23824 (N_23824,N_17301,N_17610);
and U23825 (N_23825,N_14338,N_13649);
nand U23826 (N_23826,N_13927,N_16077);
nand U23827 (N_23827,N_17342,N_17133);
or U23828 (N_23828,N_18744,N_18096);
xnor U23829 (N_23829,N_14390,N_18207);
or U23830 (N_23830,N_13862,N_16941);
and U23831 (N_23831,N_14871,N_13120);
and U23832 (N_23832,N_12884,N_15774);
nand U23833 (N_23833,N_17728,N_18726);
nand U23834 (N_23834,N_17304,N_17486);
and U23835 (N_23835,N_17678,N_13099);
and U23836 (N_23836,N_14887,N_12762);
nand U23837 (N_23837,N_12634,N_14813);
nor U23838 (N_23838,N_16270,N_18124);
xnor U23839 (N_23839,N_13811,N_16779);
nor U23840 (N_23840,N_13759,N_18097);
nor U23841 (N_23841,N_17219,N_15891);
and U23842 (N_23842,N_14050,N_16192);
nand U23843 (N_23843,N_15119,N_12552);
and U23844 (N_23844,N_18327,N_14690);
and U23845 (N_23845,N_14324,N_18335);
or U23846 (N_23846,N_16824,N_14948);
and U23847 (N_23847,N_12807,N_16082);
nor U23848 (N_23848,N_14490,N_13664);
and U23849 (N_23849,N_13320,N_13170);
nor U23850 (N_23850,N_18379,N_16781);
and U23851 (N_23851,N_16074,N_18173);
xor U23852 (N_23852,N_18005,N_12800);
or U23853 (N_23853,N_14274,N_14053);
and U23854 (N_23854,N_15232,N_15784);
and U23855 (N_23855,N_14273,N_18522);
xor U23856 (N_23856,N_14033,N_16569);
and U23857 (N_23857,N_15403,N_12800);
xnor U23858 (N_23858,N_17264,N_13175);
nand U23859 (N_23859,N_13966,N_15814);
nor U23860 (N_23860,N_18322,N_14940);
nand U23861 (N_23861,N_16634,N_16544);
and U23862 (N_23862,N_15768,N_12675);
nor U23863 (N_23863,N_17923,N_14016);
nor U23864 (N_23864,N_17116,N_18242);
nand U23865 (N_23865,N_16000,N_17232);
and U23866 (N_23866,N_13787,N_14727);
and U23867 (N_23867,N_15059,N_16242);
nand U23868 (N_23868,N_18041,N_15880);
and U23869 (N_23869,N_15114,N_15549);
or U23870 (N_23870,N_16081,N_14571);
nor U23871 (N_23871,N_17168,N_15289);
or U23872 (N_23872,N_13372,N_18517);
nand U23873 (N_23873,N_15634,N_16263);
or U23874 (N_23874,N_17882,N_17333);
or U23875 (N_23875,N_16443,N_18558);
or U23876 (N_23876,N_17531,N_16697);
or U23877 (N_23877,N_14704,N_17772);
nand U23878 (N_23878,N_14847,N_16034);
or U23879 (N_23879,N_17466,N_12591);
and U23880 (N_23880,N_17890,N_15899);
and U23881 (N_23881,N_13854,N_15400);
nor U23882 (N_23882,N_16060,N_14120);
and U23883 (N_23883,N_18168,N_17072);
xor U23884 (N_23884,N_15820,N_16749);
nand U23885 (N_23885,N_18605,N_16653);
nor U23886 (N_23886,N_17692,N_18586);
nand U23887 (N_23887,N_12558,N_18420);
or U23888 (N_23888,N_13812,N_13386);
and U23889 (N_23889,N_13017,N_14158);
nand U23890 (N_23890,N_15340,N_12645);
and U23891 (N_23891,N_14454,N_16287);
nor U23892 (N_23892,N_18053,N_14175);
xnor U23893 (N_23893,N_15604,N_18282);
and U23894 (N_23894,N_16076,N_18538);
nor U23895 (N_23895,N_18609,N_15773);
nand U23896 (N_23896,N_12834,N_15603);
nand U23897 (N_23897,N_17341,N_16288);
nor U23898 (N_23898,N_17942,N_15603);
nor U23899 (N_23899,N_15551,N_16529);
and U23900 (N_23900,N_14352,N_16669);
nand U23901 (N_23901,N_17881,N_14071);
and U23902 (N_23902,N_16700,N_14100);
nand U23903 (N_23903,N_18357,N_14266);
nand U23904 (N_23904,N_15754,N_16086);
or U23905 (N_23905,N_13974,N_17591);
nor U23906 (N_23906,N_13031,N_17636);
and U23907 (N_23907,N_15683,N_14236);
or U23908 (N_23908,N_17432,N_15897);
nand U23909 (N_23909,N_18718,N_16774);
nor U23910 (N_23910,N_12508,N_14743);
and U23911 (N_23911,N_14755,N_17023);
nand U23912 (N_23912,N_17878,N_12855);
nor U23913 (N_23913,N_17046,N_14811);
nand U23914 (N_23914,N_17706,N_15256);
nor U23915 (N_23915,N_17795,N_14324);
and U23916 (N_23916,N_16750,N_18358);
and U23917 (N_23917,N_15503,N_17786);
xnor U23918 (N_23918,N_17140,N_16147);
or U23919 (N_23919,N_14683,N_18156);
and U23920 (N_23920,N_16963,N_13891);
or U23921 (N_23921,N_12871,N_14935);
nor U23922 (N_23922,N_18439,N_15702);
xnor U23923 (N_23923,N_15254,N_14968);
nor U23924 (N_23924,N_14221,N_14463);
xnor U23925 (N_23925,N_14291,N_12943);
nand U23926 (N_23926,N_14711,N_18320);
and U23927 (N_23927,N_18098,N_17613);
and U23928 (N_23928,N_17999,N_17706);
or U23929 (N_23929,N_16239,N_14063);
nor U23930 (N_23930,N_15114,N_13364);
nand U23931 (N_23931,N_18001,N_17122);
and U23932 (N_23932,N_16382,N_14587);
and U23933 (N_23933,N_16344,N_14479);
or U23934 (N_23934,N_14532,N_14805);
and U23935 (N_23935,N_15464,N_18673);
nand U23936 (N_23936,N_17399,N_12817);
nand U23937 (N_23937,N_18067,N_12683);
nand U23938 (N_23938,N_14721,N_18271);
xnor U23939 (N_23939,N_17830,N_15870);
nor U23940 (N_23940,N_14094,N_14805);
nor U23941 (N_23941,N_14373,N_16951);
nor U23942 (N_23942,N_12820,N_13752);
or U23943 (N_23943,N_14065,N_12798);
and U23944 (N_23944,N_17607,N_13218);
xor U23945 (N_23945,N_12672,N_18231);
nand U23946 (N_23946,N_12654,N_14800);
nand U23947 (N_23947,N_16567,N_17266);
xnor U23948 (N_23948,N_17013,N_16098);
and U23949 (N_23949,N_15459,N_17298);
xor U23950 (N_23950,N_12633,N_18460);
nand U23951 (N_23951,N_14546,N_15575);
nor U23952 (N_23952,N_13694,N_16788);
nor U23953 (N_23953,N_17848,N_14796);
nor U23954 (N_23954,N_14278,N_14797);
and U23955 (N_23955,N_16222,N_17343);
or U23956 (N_23956,N_13673,N_16217);
nor U23957 (N_23957,N_18237,N_15675);
xor U23958 (N_23958,N_18227,N_13628);
and U23959 (N_23959,N_13454,N_17772);
nor U23960 (N_23960,N_13560,N_16502);
nand U23961 (N_23961,N_18505,N_13808);
nor U23962 (N_23962,N_12532,N_14749);
nand U23963 (N_23963,N_13714,N_16468);
nor U23964 (N_23964,N_18467,N_18552);
xnor U23965 (N_23965,N_16152,N_14768);
or U23966 (N_23966,N_16809,N_17934);
xnor U23967 (N_23967,N_16685,N_15199);
nor U23968 (N_23968,N_13130,N_16517);
nor U23969 (N_23969,N_18048,N_12611);
and U23970 (N_23970,N_12524,N_17138);
and U23971 (N_23971,N_18321,N_17498);
nand U23972 (N_23972,N_14959,N_15636);
nand U23973 (N_23973,N_14237,N_12580);
and U23974 (N_23974,N_16310,N_16043);
and U23975 (N_23975,N_14869,N_17623);
nor U23976 (N_23976,N_12520,N_13065);
or U23977 (N_23977,N_17501,N_14352);
nand U23978 (N_23978,N_13908,N_13822);
or U23979 (N_23979,N_13429,N_18498);
and U23980 (N_23980,N_17770,N_16475);
xnor U23981 (N_23981,N_15363,N_15370);
and U23982 (N_23982,N_15959,N_18562);
nand U23983 (N_23983,N_15293,N_16969);
and U23984 (N_23984,N_18298,N_17821);
or U23985 (N_23985,N_12552,N_18163);
or U23986 (N_23986,N_13260,N_17024);
xor U23987 (N_23987,N_16036,N_16144);
nor U23988 (N_23988,N_14894,N_15122);
and U23989 (N_23989,N_15036,N_16870);
and U23990 (N_23990,N_16248,N_18109);
nand U23991 (N_23991,N_14956,N_17275);
nand U23992 (N_23992,N_16997,N_14867);
and U23993 (N_23993,N_17709,N_12641);
nand U23994 (N_23994,N_17191,N_12762);
or U23995 (N_23995,N_13437,N_12957);
and U23996 (N_23996,N_18693,N_16547);
nor U23997 (N_23997,N_15606,N_18428);
or U23998 (N_23998,N_16581,N_16779);
nand U23999 (N_23999,N_18564,N_16708);
or U24000 (N_24000,N_14384,N_17068);
nand U24001 (N_24001,N_13615,N_14526);
or U24002 (N_24002,N_18428,N_13931);
nand U24003 (N_24003,N_18584,N_18722);
nor U24004 (N_24004,N_15270,N_17386);
and U24005 (N_24005,N_15738,N_18077);
nand U24006 (N_24006,N_13561,N_16788);
and U24007 (N_24007,N_14088,N_13843);
nand U24008 (N_24008,N_16420,N_17470);
nor U24009 (N_24009,N_14372,N_13597);
nor U24010 (N_24010,N_18232,N_18661);
nor U24011 (N_24011,N_13010,N_16483);
and U24012 (N_24012,N_16216,N_13939);
nor U24013 (N_24013,N_14532,N_14011);
nor U24014 (N_24014,N_17857,N_13767);
xnor U24015 (N_24015,N_16456,N_14161);
and U24016 (N_24016,N_12724,N_13598);
or U24017 (N_24017,N_13552,N_16970);
xor U24018 (N_24018,N_13127,N_13414);
or U24019 (N_24019,N_14881,N_16585);
or U24020 (N_24020,N_18328,N_16204);
nand U24021 (N_24021,N_15803,N_13234);
nor U24022 (N_24022,N_13772,N_13300);
nand U24023 (N_24023,N_17716,N_16994);
nand U24024 (N_24024,N_14232,N_13454);
nor U24025 (N_24025,N_16019,N_18499);
or U24026 (N_24026,N_14608,N_12796);
nand U24027 (N_24027,N_13193,N_18469);
nor U24028 (N_24028,N_15702,N_12633);
nor U24029 (N_24029,N_13345,N_17895);
nor U24030 (N_24030,N_14683,N_18511);
nor U24031 (N_24031,N_15362,N_17814);
nor U24032 (N_24032,N_13559,N_15356);
nand U24033 (N_24033,N_17508,N_13123);
nand U24034 (N_24034,N_14103,N_13245);
and U24035 (N_24035,N_17220,N_13181);
nor U24036 (N_24036,N_12577,N_13941);
nand U24037 (N_24037,N_13802,N_18696);
or U24038 (N_24038,N_13671,N_18210);
xnor U24039 (N_24039,N_13519,N_12689);
nor U24040 (N_24040,N_16831,N_13056);
and U24041 (N_24041,N_15049,N_17482);
or U24042 (N_24042,N_14937,N_15149);
nor U24043 (N_24043,N_16860,N_15374);
or U24044 (N_24044,N_14885,N_16361);
and U24045 (N_24045,N_16037,N_16764);
or U24046 (N_24046,N_18517,N_15688);
nand U24047 (N_24047,N_12540,N_17907);
nand U24048 (N_24048,N_16692,N_13591);
or U24049 (N_24049,N_18296,N_13578);
nand U24050 (N_24050,N_13763,N_18024);
and U24051 (N_24051,N_15880,N_17269);
nand U24052 (N_24052,N_18461,N_14296);
and U24053 (N_24053,N_17145,N_12971);
nor U24054 (N_24054,N_14136,N_14784);
nand U24055 (N_24055,N_16665,N_13391);
and U24056 (N_24056,N_16352,N_17045);
nor U24057 (N_24057,N_14811,N_13023);
nand U24058 (N_24058,N_15096,N_16367);
or U24059 (N_24059,N_18295,N_17796);
nand U24060 (N_24060,N_15958,N_15241);
nand U24061 (N_24061,N_16781,N_13264);
nor U24062 (N_24062,N_17636,N_13301);
nor U24063 (N_24063,N_14346,N_16357);
or U24064 (N_24064,N_12560,N_16629);
nand U24065 (N_24065,N_15500,N_16820);
xor U24066 (N_24066,N_15031,N_16943);
nand U24067 (N_24067,N_14313,N_12918);
and U24068 (N_24068,N_14911,N_16397);
or U24069 (N_24069,N_14752,N_14009);
nor U24070 (N_24070,N_17187,N_17114);
and U24071 (N_24071,N_14644,N_13884);
or U24072 (N_24072,N_14601,N_13128);
and U24073 (N_24073,N_18615,N_16326);
nor U24074 (N_24074,N_18018,N_17120);
nor U24075 (N_24075,N_15635,N_15759);
and U24076 (N_24076,N_14809,N_17590);
and U24077 (N_24077,N_17283,N_16257);
nor U24078 (N_24078,N_14116,N_13583);
nor U24079 (N_24079,N_15226,N_13469);
and U24080 (N_24080,N_16074,N_15481);
and U24081 (N_24081,N_17227,N_14379);
xnor U24082 (N_24082,N_14125,N_17443);
xor U24083 (N_24083,N_12975,N_16652);
and U24084 (N_24084,N_15876,N_15566);
or U24085 (N_24085,N_16217,N_13452);
nand U24086 (N_24086,N_15691,N_15494);
or U24087 (N_24087,N_18285,N_18527);
xor U24088 (N_24088,N_17432,N_12551);
or U24089 (N_24089,N_14900,N_17489);
nor U24090 (N_24090,N_13117,N_18597);
xor U24091 (N_24091,N_16835,N_13164);
or U24092 (N_24092,N_13852,N_15008);
nor U24093 (N_24093,N_15372,N_14424);
nor U24094 (N_24094,N_16401,N_18743);
nand U24095 (N_24095,N_15020,N_17763);
nor U24096 (N_24096,N_16877,N_14825);
xnor U24097 (N_24097,N_16239,N_16803);
or U24098 (N_24098,N_16991,N_16524);
and U24099 (N_24099,N_17235,N_14839);
and U24100 (N_24100,N_12739,N_16123);
and U24101 (N_24101,N_17924,N_16519);
nor U24102 (N_24102,N_13575,N_17593);
and U24103 (N_24103,N_15705,N_12714);
nand U24104 (N_24104,N_17246,N_12598);
or U24105 (N_24105,N_15068,N_18391);
nand U24106 (N_24106,N_12585,N_12645);
nand U24107 (N_24107,N_18729,N_13321);
or U24108 (N_24108,N_12705,N_13329);
or U24109 (N_24109,N_12519,N_17447);
and U24110 (N_24110,N_13422,N_13457);
or U24111 (N_24111,N_17396,N_16304);
and U24112 (N_24112,N_17986,N_12938);
nor U24113 (N_24113,N_12899,N_18258);
and U24114 (N_24114,N_18025,N_16537);
xnor U24115 (N_24115,N_16127,N_16109);
nand U24116 (N_24116,N_14303,N_16258);
and U24117 (N_24117,N_18098,N_15040);
xor U24118 (N_24118,N_16087,N_14233);
and U24119 (N_24119,N_18452,N_15664);
nand U24120 (N_24120,N_12682,N_14567);
nor U24121 (N_24121,N_15510,N_16347);
nand U24122 (N_24122,N_13232,N_12514);
and U24123 (N_24123,N_18219,N_13127);
and U24124 (N_24124,N_16266,N_17372);
nand U24125 (N_24125,N_16591,N_17283);
and U24126 (N_24126,N_14193,N_18410);
and U24127 (N_24127,N_14340,N_16441);
xnor U24128 (N_24128,N_17148,N_14302);
or U24129 (N_24129,N_13149,N_16907);
nand U24130 (N_24130,N_14823,N_17322);
or U24131 (N_24131,N_14397,N_15887);
nand U24132 (N_24132,N_15459,N_15890);
nand U24133 (N_24133,N_13122,N_18698);
nand U24134 (N_24134,N_15680,N_12883);
nor U24135 (N_24135,N_17789,N_14183);
or U24136 (N_24136,N_17823,N_12665);
nor U24137 (N_24137,N_12904,N_16856);
and U24138 (N_24138,N_16010,N_18581);
nand U24139 (N_24139,N_16864,N_18677);
or U24140 (N_24140,N_15735,N_15040);
xnor U24141 (N_24141,N_12523,N_13362);
or U24142 (N_24142,N_15815,N_18452);
nand U24143 (N_24143,N_16724,N_18162);
or U24144 (N_24144,N_16911,N_16647);
and U24145 (N_24145,N_17735,N_17953);
xnor U24146 (N_24146,N_17584,N_14229);
or U24147 (N_24147,N_16804,N_14129);
nor U24148 (N_24148,N_16232,N_13520);
or U24149 (N_24149,N_13168,N_16090);
or U24150 (N_24150,N_12798,N_15241);
nor U24151 (N_24151,N_12552,N_16932);
and U24152 (N_24152,N_18497,N_16954);
nand U24153 (N_24153,N_18036,N_17023);
nand U24154 (N_24154,N_16784,N_17730);
and U24155 (N_24155,N_17228,N_14668);
or U24156 (N_24156,N_16042,N_16453);
and U24157 (N_24157,N_17674,N_13097);
and U24158 (N_24158,N_14478,N_16813);
and U24159 (N_24159,N_17811,N_14007);
nor U24160 (N_24160,N_12891,N_18099);
and U24161 (N_24161,N_18642,N_13685);
nand U24162 (N_24162,N_14604,N_16054);
xnor U24163 (N_24163,N_13210,N_17764);
or U24164 (N_24164,N_15177,N_16329);
nand U24165 (N_24165,N_16471,N_17201);
or U24166 (N_24166,N_14847,N_16275);
nor U24167 (N_24167,N_17868,N_17944);
and U24168 (N_24168,N_14285,N_16310);
and U24169 (N_24169,N_16496,N_16723);
nor U24170 (N_24170,N_14516,N_15021);
nor U24171 (N_24171,N_16940,N_15679);
nand U24172 (N_24172,N_13403,N_17200);
or U24173 (N_24173,N_15779,N_14915);
and U24174 (N_24174,N_15520,N_18488);
or U24175 (N_24175,N_13949,N_12772);
nor U24176 (N_24176,N_14517,N_16613);
and U24177 (N_24177,N_14706,N_14779);
and U24178 (N_24178,N_17151,N_17578);
nor U24179 (N_24179,N_13565,N_18482);
nor U24180 (N_24180,N_14796,N_14061);
nand U24181 (N_24181,N_16512,N_15609);
or U24182 (N_24182,N_17826,N_15318);
xor U24183 (N_24183,N_12639,N_12627);
xor U24184 (N_24184,N_16606,N_18664);
or U24185 (N_24185,N_17561,N_17973);
and U24186 (N_24186,N_16298,N_13567);
nor U24187 (N_24187,N_18481,N_17631);
nor U24188 (N_24188,N_17064,N_15293);
nor U24189 (N_24189,N_17394,N_12517);
or U24190 (N_24190,N_15692,N_14364);
or U24191 (N_24191,N_18526,N_14531);
and U24192 (N_24192,N_18035,N_13698);
xnor U24193 (N_24193,N_16276,N_13265);
and U24194 (N_24194,N_13114,N_18124);
and U24195 (N_24195,N_13883,N_16145);
nor U24196 (N_24196,N_16433,N_12631);
and U24197 (N_24197,N_12529,N_18425);
and U24198 (N_24198,N_15607,N_14424);
nand U24199 (N_24199,N_18526,N_17058);
or U24200 (N_24200,N_13899,N_14121);
and U24201 (N_24201,N_16138,N_15381);
and U24202 (N_24202,N_15662,N_12664);
nor U24203 (N_24203,N_13942,N_17458);
and U24204 (N_24204,N_17242,N_17194);
and U24205 (N_24205,N_16921,N_16595);
and U24206 (N_24206,N_13957,N_15285);
and U24207 (N_24207,N_14206,N_18014);
nor U24208 (N_24208,N_12888,N_12908);
xor U24209 (N_24209,N_16048,N_12983);
nor U24210 (N_24210,N_13288,N_15514);
nand U24211 (N_24211,N_18028,N_15135);
and U24212 (N_24212,N_16452,N_17933);
or U24213 (N_24213,N_14154,N_15709);
or U24214 (N_24214,N_15520,N_12836);
nor U24215 (N_24215,N_16219,N_15601);
nand U24216 (N_24216,N_16541,N_14528);
and U24217 (N_24217,N_14128,N_15899);
and U24218 (N_24218,N_17473,N_16898);
and U24219 (N_24219,N_18387,N_15200);
nand U24220 (N_24220,N_18345,N_13861);
nor U24221 (N_24221,N_12911,N_18071);
nand U24222 (N_24222,N_13552,N_16228);
nand U24223 (N_24223,N_12890,N_14019);
and U24224 (N_24224,N_13523,N_15932);
nor U24225 (N_24225,N_15289,N_16648);
nor U24226 (N_24226,N_16150,N_14548);
and U24227 (N_24227,N_15257,N_14508);
or U24228 (N_24228,N_14652,N_18306);
or U24229 (N_24229,N_18229,N_15022);
nor U24230 (N_24230,N_15485,N_16359);
xor U24231 (N_24231,N_17440,N_16000);
nand U24232 (N_24232,N_15702,N_16882);
nand U24233 (N_24233,N_16052,N_16944);
nand U24234 (N_24234,N_17572,N_18227);
nor U24235 (N_24235,N_15801,N_12502);
nand U24236 (N_24236,N_14331,N_18272);
and U24237 (N_24237,N_17207,N_18625);
or U24238 (N_24238,N_16756,N_15024);
nand U24239 (N_24239,N_13675,N_14272);
or U24240 (N_24240,N_18139,N_18021);
or U24241 (N_24241,N_17697,N_16495);
or U24242 (N_24242,N_16265,N_13054);
and U24243 (N_24243,N_13546,N_13952);
or U24244 (N_24244,N_18017,N_14993);
nor U24245 (N_24245,N_18208,N_15166);
and U24246 (N_24246,N_15274,N_15363);
nor U24247 (N_24247,N_12527,N_16375);
nand U24248 (N_24248,N_17857,N_18359);
nand U24249 (N_24249,N_17220,N_17765);
nand U24250 (N_24250,N_17841,N_15249);
nand U24251 (N_24251,N_15609,N_15919);
nor U24252 (N_24252,N_16824,N_14708);
and U24253 (N_24253,N_18737,N_17968);
xnor U24254 (N_24254,N_16868,N_16442);
or U24255 (N_24255,N_17436,N_14072);
xnor U24256 (N_24256,N_13814,N_13108);
nand U24257 (N_24257,N_17352,N_13544);
xor U24258 (N_24258,N_14427,N_17680);
nor U24259 (N_24259,N_13768,N_17190);
nor U24260 (N_24260,N_15969,N_17458);
or U24261 (N_24261,N_16248,N_17050);
or U24262 (N_24262,N_15736,N_15997);
and U24263 (N_24263,N_16564,N_16591);
nor U24264 (N_24264,N_13079,N_13333);
nor U24265 (N_24265,N_13484,N_14148);
or U24266 (N_24266,N_15540,N_15372);
or U24267 (N_24267,N_13592,N_14432);
xor U24268 (N_24268,N_16778,N_14464);
and U24269 (N_24269,N_14689,N_14142);
or U24270 (N_24270,N_18242,N_15771);
or U24271 (N_24271,N_14957,N_13617);
or U24272 (N_24272,N_18456,N_16997);
nand U24273 (N_24273,N_15044,N_14886);
nor U24274 (N_24274,N_14482,N_14764);
xnor U24275 (N_24275,N_14714,N_18127);
or U24276 (N_24276,N_15302,N_15828);
nand U24277 (N_24277,N_17056,N_16614);
nand U24278 (N_24278,N_17994,N_14861);
and U24279 (N_24279,N_14558,N_17329);
nor U24280 (N_24280,N_16234,N_16476);
nand U24281 (N_24281,N_16608,N_15482);
nor U24282 (N_24282,N_13562,N_15663);
nand U24283 (N_24283,N_13329,N_16571);
and U24284 (N_24284,N_17609,N_13744);
and U24285 (N_24285,N_15724,N_14760);
or U24286 (N_24286,N_16759,N_18435);
nor U24287 (N_24287,N_14617,N_14193);
nor U24288 (N_24288,N_14787,N_18008);
nand U24289 (N_24289,N_17302,N_14774);
xor U24290 (N_24290,N_18331,N_13861);
or U24291 (N_24291,N_15540,N_15598);
or U24292 (N_24292,N_18689,N_14691);
or U24293 (N_24293,N_13833,N_18131);
and U24294 (N_24294,N_15008,N_17415);
or U24295 (N_24295,N_17332,N_17352);
or U24296 (N_24296,N_14099,N_16748);
nand U24297 (N_24297,N_16096,N_12592);
nand U24298 (N_24298,N_16671,N_18694);
nand U24299 (N_24299,N_16064,N_18738);
nor U24300 (N_24300,N_13729,N_17120);
nand U24301 (N_24301,N_16742,N_16462);
and U24302 (N_24302,N_13360,N_16611);
nor U24303 (N_24303,N_13547,N_16920);
nand U24304 (N_24304,N_17103,N_13786);
nand U24305 (N_24305,N_18423,N_17896);
nor U24306 (N_24306,N_14210,N_18192);
or U24307 (N_24307,N_13287,N_17753);
nand U24308 (N_24308,N_15106,N_13520);
nor U24309 (N_24309,N_16775,N_14812);
nand U24310 (N_24310,N_15564,N_16550);
nand U24311 (N_24311,N_14249,N_15510);
xor U24312 (N_24312,N_18128,N_15351);
and U24313 (N_24313,N_16320,N_16776);
or U24314 (N_24314,N_14416,N_16883);
and U24315 (N_24315,N_16039,N_12584);
nor U24316 (N_24316,N_15179,N_13365);
nor U24317 (N_24317,N_13714,N_13384);
nor U24318 (N_24318,N_16263,N_14313);
nand U24319 (N_24319,N_15622,N_12711);
nor U24320 (N_24320,N_15672,N_13268);
or U24321 (N_24321,N_12684,N_17735);
and U24322 (N_24322,N_16901,N_14607);
nand U24323 (N_24323,N_15464,N_14015);
or U24324 (N_24324,N_12824,N_17232);
nor U24325 (N_24325,N_15246,N_17597);
nand U24326 (N_24326,N_15356,N_15709);
or U24327 (N_24327,N_13442,N_14818);
nor U24328 (N_24328,N_17658,N_14367);
nand U24329 (N_24329,N_16222,N_14966);
nand U24330 (N_24330,N_14454,N_17879);
nand U24331 (N_24331,N_12972,N_18508);
nand U24332 (N_24332,N_18278,N_17289);
nand U24333 (N_24333,N_14359,N_12916);
nand U24334 (N_24334,N_14968,N_17914);
or U24335 (N_24335,N_17670,N_16287);
and U24336 (N_24336,N_16114,N_15438);
or U24337 (N_24337,N_12630,N_16804);
nand U24338 (N_24338,N_17996,N_13170);
xnor U24339 (N_24339,N_16240,N_18451);
nor U24340 (N_24340,N_18147,N_15288);
or U24341 (N_24341,N_15221,N_17158);
or U24342 (N_24342,N_14429,N_16941);
or U24343 (N_24343,N_17098,N_14727);
or U24344 (N_24344,N_17924,N_14218);
or U24345 (N_24345,N_18743,N_15682);
and U24346 (N_24346,N_15561,N_12940);
and U24347 (N_24347,N_16218,N_12833);
and U24348 (N_24348,N_17825,N_15012);
nand U24349 (N_24349,N_17274,N_14754);
or U24350 (N_24350,N_14877,N_17827);
nor U24351 (N_24351,N_18692,N_17683);
nand U24352 (N_24352,N_18212,N_14159);
nand U24353 (N_24353,N_14236,N_14723);
and U24354 (N_24354,N_15297,N_12975);
or U24355 (N_24355,N_13738,N_16676);
nand U24356 (N_24356,N_13067,N_15064);
nand U24357 (N_24357,N_14988,N_12609);
nor U24358 (N_24358,N_13690,N_14219);
nand U24359 (N_24359,N_13905,N_18465);
nor U24360 (N_24360,N_18701,N_16524);
or U24361 (N_24361,N_17992,N_15261);
or U24362 (N_24362,N_16366,N_13975);
or U24363 (N_24363,N_17183,N_17258);
or U24364 (N_24364,N_12729,N_12585);
or U24365 (N_24365,N_18634,N_15135);
nand U24366 (N_24366,N_12841,N_13390);
nor U24367 (N_24367,N_17563,N_14545);
or U24368 (N_24368,N_16631,N_14172);
nand U24369 (N_24369,N_14972,N_17570);
or U24370 (N_24370,N_14137,N_17727);
nor U24371 (N_24371,N_13535,N_18277);
nor U24372 (N_24372,N_13644,N_12614);
nand U24373 (N_24373,N_14039,N_14737);
nand U24374 (N_24374,N_13024,N_17032);
or U24375 (N_24375,N_12688,N_17379);
nand U24376 (N_24376,N_13890,N_17791);
nor U24377 (N_24377,N_18181,N_18257);
nor U24378 (N_24378,N_13578,N_13666);
nor U24379 (N_24379,N_12680,N_18660);
nor U24380 (N_24380,N_14263,N_15220);
and U24381 (N_24381,N_14945,N_16563);
and U24382 (N_24382,N_13182,N_14230);
and U24383 (N_24383,N_14029,N_15847);
and U24384 (N_24384,N_13415,N_15499);
and U24385 (N_24385,N_15007,N_16978);
nand U24386 (N_24386,N_17499,N_16480);
and U24387 (N_24387,N_17391,N_15313);
and U24388 (N_24388,N_17622,N_14666);
and U24389 (N_24389,N_16153,N_17025);
or U24390 (N_24390,N_13732,N_16977);
nand U24391 (N_24391,N_16113,N_15098);
or U24392 (N_24392,N_12868,N_13715);
or U24393 (N_24393,N_18067,N_17898);
nor U24394 (N_24394,N_17379,N_13677);
nand U24395 (N_24395,N_13133,N_13636);
or U24396 (N_24396,N_14427,N_15478);
nand U24397 (N_24397,N_18616,N_14693);
and U24398 (N_24398,N_14228,N_18381);
or U24399 (N_24399,N_13547,N_12650);
nor U24400 (N_24400,N_16822,N_13846);
nand U24401 (N_24401,N_13102,N_16966);
nand U24402 (N_24402,N_16254,N_17335);
nor U24403 (N_24403,N_17881,N_13028);
or U24404 (N_24404,N_16010,N_15178);
or U24405 (N_24405,N_18308,N_18615);
nand U24406 (N_24406,N_14919,N_14994);
or U24407 (N_24407,N_15548,N_14016);
nor U24408 (N_24408,N_15059,N_13087);
nor U24409 (N_24409,N_18078,N_14617);
or U24410 (N_24410,N_14363,N_18581);
nand U24411 (N_24411,N_17191,N_18682);
nand U24412 (N_24412,N_14004,N_16914);
and U24413 (N_24413,N_13849,N_13072);
nor U24414 (N_24414,N_14221,N_13286);
nand U24415 (N_24415,N_17627,N_15113);
or U24416 (N_24416,N_17586,N_14827);
and U24417 (N_24417,N_17337,N_14700);
nand U24418 (N_24418,N_17546,N_16375);
xor U24419 (N_24419,N_13933,N_14210);
nor U24420 (N_24420,N_15605,N_15553);
or U24421 (N_24421,N_18202,N_15830);
xnor U24422 (N_24422,N_18256,N_15696);
and U24423 (N_24423,N_15044,N_17222);
nand U24424 (N_24424,N_17585,N_15650);
nor U24425 (N_24425,N_15462,N_18434);
and U24426 (N_24426,N_17118,N_15261);
nor U24427 (N_24427,N_16663,N_15869);
nor U24428 (N_24428,N_12541,N_18449);
and U24429 (N_24429,N_15449,N_16776);
nand U24430 (N_24430,N_17646,N_14696);
nor U24431 (N_24431,N_15258,N_13775);
nand U24432 (N_24432,N_17176,N_14856);
or U24433 (N_24433,N_15891,N_14407);
nor U24434 (N_24434,N_13733,N_14783);
or U24435 (N_24435,N_17655,N_13237);
nand U24436 (N_24436,N_17138,N_15431);
and U24437 (N_24437,N_17022,N_16575);
nor U24438 (N_24438,N_13530,N_16289);
nand U24439 (N_24439,N_13260,N_16130);
or U24440 (N_24440,N_14862,N_18088);
nor U24441 (N_24441,N_13636,N_15811);
and U24442 (N_24442,N_17775,N_13904);
nand U24443 (N_24443,N_17849,N_17063);
or U24444 (N_24444,N_16458,N_16228);
nand U24445 (N_24445,N_14572,N_14952);
nand U24446 (N_24446,N_17758,N_14104);
or U24447 (N_24447,N_13615,N_14890);
and U24448 (N_24448,N_17251,N_13980);
nand U24449 (N_24449,N_15240,N_14127);
nor U24450 (N_24450,N_15050,N_13882);
or U24451 (N_24451,N_14159,N_17205);
and U24452 (N_24452,N_15045,N_15006);
nand U24453 (N_24453,N_13575,N_16748);
xor U24454 (N_24454,N_18282,N_15649);
nor U24455 (N_24455,N_15598,N_15440);
xnor U24456 (N_24456,N_12503,N_14682);
nand U24457 (N_24457,N_15714,N_14497);
xnor U24458 (N_24458,N_15106,N_16318);
nor U24459 (N_24459,N_12827,N_18036);
and U24460 (N_24460,N_14144,N_16460);
and U24461 (N_24461,N_15840,N_14812);
nand U24462 (N_24462,N_13166,N_14177);
nand U24463 (N_24463,N_16214,N_17830);
nand U24464 (N_24464,N_15822,N_15773);
xor U24465 (N_24465,N_14083,N_16476);
nor U24466 (N_24466,N_17867,N_16654);
and U24467 (N_24467,N_16307,N_13790);
and U24468 (N_24468,N_18045,N_17760);
or U24469 (N_24469,N_18054,N_17922);
and U24470 (N_24470,N_13994,N_15063);
and U24471 (N_24471,N_16709,N_17766);
or U24472 (N_24472,N_18546,N_16502);
nand U24473 (N_24473,N_14007,N_18047);
nand U24474 (N_24474,N_14968,N_12558);
or U24475 (N_24475,N_13584,N_17822);
nor U24476 (N_24476,N_14800,N_17846);
nand U24477 (N_24477,N_18471,N_16563);
nand U24478 (N_24478,N_15230,N_18583);
or U24479 (N_24479,N_18108,N_12789);
and U24480 (N_24480,N_14946,N_17571);
nor U24481 (N_24481,N_16864,N_18742);
nor U24482 (N_24482,N_18476,N_14633);
nand U24483 (N_24483,N_17455,N_15236);
nand U24484 (N_24484,N_15084,N_16898);
and U24485 (N_24485,N_14543,N_18536);
and U24486 (N_24486,N_12617,N_14658);
xnor U24487 (N_24487,N_16549,N_18649);
xnor U24488 (N_24488,N_18402,N_17029);
nand U24489 (N_24489,N_12940,N_18335);
or U24490 (N_24490,N_18686,N_16863);
nand U24491 (N_24491,N_14296,N_12511);
nand U24492 (N_24492,N_15367,N_18140);
or U24493 (N_24493,N_16861,N_14189);
nor U24494 (N_24494,N_17035,N_13919);
and U24495 (N_24495,N_14044,N_12999);
nor U24496 (N_24496,N_15836,N_14992);
and U24497 (N_24497,N_18559,N_18172);
xor U24498 (N_24498,N_16474,N_18224);
nand U24499 (N_24499,N_13082,N_12910);
or U24500 (N_24500,N_14731,N_15383);
nand U24501 (N_24501,N_18710,N_14073);
nand U24502 (N_24502,N_13167,N_12976);
and U24503 (N_24503,N_12815,N_13210);
nor U24504 (N_24504,N_16430,N_16099);
or U24505 (N_24505,N_16423,N_17293);
nor U24506 (N_24506,N_16543,N_17009);
or U24507 (N_24507,N_18458,N_12770);
nand U24508 (N_24508,N_16944,N_13738);
nor U24509 (N_24509,N_14435,N_16815);
nor U24510 (N_24510,N_12727,N_18344);
xor U24511 (N_24511,N_15856,N_14294);
nand U24512 (N_24512,N_17983,N_16471);
and U24513 (N_24513,N_12794,N_14937);
nor U24514 (N_24514,N_18061,N_16745);
nand U24515 (N_24515,N_15135,N_13068);
nor U24516 (N_24516,N_14070,N_15689);
or U24517 (N_24517,N_17265,N_13696);
and U24518 (N_24518,N_13615,N_12747);
xnor U24519 (N_24519,N_16425,N_18073);
nor U24520 (N_24520,N_12522,N_14159);
nand U24521 (N_24521,N_15182,N_17399);
and U24522 (N_24522,N_16357,N_18425);
nor U24523 (N_24523,N_14530,N_17440);
nand U24524 (N_24524,N_13961,N_17192);
xor U24525 (N_24525,N_17041,N_16740);
xnor U24526 (N_24526,N_14035,N_12747);
and U24527 (N_24527,N_12902,N_13312);
or U24528 (N_24528,N_14101,N_17193);
and U24529 (N_24529,N_12535,N_15973);
nand U24530 (N_24530,N_13789,N_13297);
nand U24531 (N_24531,N_17389,N_15099);
and U24532 (N_24532,N_17322,N_12863);
or U24533 (N_24533,N_18577,N_14294);
and U24534 (N_24534,N_12912,N_18391);
xor U24535 (N_24535,N_16925,N_17487);
or U24536 (N_24536,N_12517,N_13370);
or U24537 (N_24537,N_15009,N_17807);
nand U24538 (N_24538,N_17042,N_13082);
nand U24539 (N_24539,N_12843,N_14185);
and U24540 (N_24540,N_16953,N_15893);
nand U24541 (N_24541,N_18143,N_14607);
and U24542 (N_24542,N_18296,N_17057);
nand U24543 (N_24543,N_17905,N_13720);
or U24544 (N_24544,N_15123,N_12808);
xor U24545 (N_24545,N_18095,N_18711);
or U24546 (N_24546,N_14153,N_16656);
or U24547 (N_24547,N_15280,N_14572);
and U24548 (N_24548,N_12930,N_18221);
nand U24549 (N_24549,N_18579,N_12962);
and U24550 (N_24550,N_14762,N_13965);
or U24551 (N_24551,N_17890,N_16139);
or U24552 (N_24552,N_18509,N_15597);
xor U24553 (N_24553,N_15254,N_18359);
xor U24554 (N_24554,N_15958,N_16650);
nand U24555 (N_24555,N_14559,N_16885);
and U24556 (N_24556,N_13797,N_15315);
nand U24557 (N_24557,N_15760,N_15620);
and U24558 (N_24558,N_16037,N_18169);
nor U24559 (N_24559,N_13855,N_14360);
and U24560 (N_24560,N_13098,N_16688);
and U24561 (N_24561,N_15558,N_16972);
nand U24562 (N_24562,N_17444,N_17510);
or U24563 (N_24563,N_14344,N_16179);
or U24564 (N_24564,N_16234,N_14314);
nor U24565 (N_24565,N_14643,N_13795);
xor U24566 (N_24566,N_13737,N_16679);
and U24567 (N_24567,N_17185,N_16329);
or U24568 (N_24568,N_17874,N_16835);
and U24569 (N_24569,N_14578,N_12612);
or U24570 (N_24570,N_15404,N_18021);
and U24571 (N_24571,N_18341,N_15722);
nor U24572 (N_24572,N_18331,N_13172);
nand U24573 (N_24573,N_14096,N_18365);
xnor U24574 (N_24574,N_17700,N_18112);
or U24575 (N_24575,N_15601,N_15406);
nor U24576 (N_24576,N_16392,N_13675);
nor U24577 (N_24577,N_12563,N_13011);
xnor U24578 (N_24578,N_14538,N_16434);
nand U24579 (N_24579,N_15378,N_14335);
nor U24580 (N_24580,N_14029,N_14707);
nand U24581 (N_24581,N_14584,N_17051);
nand U24582 (N_24582,N_16407,N_13466);
or U24583 (N_24583,N_16245,N_13142);
nand U24584 (N_24584,N_18441,N_15845);
xnor U24585 (N_24585,N_12986,N_14160);
nand U24586 (N_24586,N_18324,N_18584);
and U24587 (N_24587,N_16881,N_16797);
and U24588 (N_24588,N_16760,N_13327);
nor U24589 (N_24589,N_13016,N_15889);
and U24590 (N_24590,N_14813,N_16833);
nand U24591 (N_24591,N_14434,N_18472);
nor U24592 (N_24592,N_18035,N_17851);
or U24593 (N_24593,N_17937,N_12995);
and U24594 (N_24594,N_14528,N_17633);
or U24595 (N_24595,N_15465,N_16621);
nand U24596 (N_24596,N_13265,N_16948);
or U24597 (N_24597,N_12745,N_14077);
xor U24598 (N_24598,N_17110,N_14661);
nor U24599 (N_24599,N_18662,N_12849);
nor U24600 (N_24600,N_17632,N_16548);
nand U24601 (N_24601,N_15901,N_16832);
or U24602 (N_24602,N_14332,N_14435);
nand U24603 (N_24603,N_15583,N_15569);
nand U24604 (N_24604,N_18018,N_14268);
or U24605 (N_24605,N_14001,N_14364);
or U24606 (N_24606,N_14446,N_12737);
xnor U24607 (N_24607,N_17235,N_13317);
or U24608 (N_24608,N_16087,N_18149);
or U24609 (N_24609,N_17648,N_14573);
nand U24610 (N_24610,N_12643,N_17560);
nand U24611 (N_24611,N_14950,N_13657);
or U24612 (N_24612,N_14531,N_18261);
nand U24613 (N_24613,N_16869,N_15203);
or U24614 (N_24614,N_12952,N_13111);
and U24615 (N_24615,N_13670,N_16201);
nor U24616 (N_24616,N_18137,N_15510);
or U24617 (N_24617,N_14737,N_17502);
and U24618 (N_24618,N_17770,N_17120);
xnor U24619 (N_24619,N_12576,N_18050);
and U24620 (N_24620,N_13712,N_13807);
nand U24621 (N_24621,N_12790,N_14061);
or U24622 (N_24622,N_18152,N_13010);
and U24623 (N_24623,N_17524,N_17029);
and U24624 (N_24624,N_18537,N_17870);
and U24625 (N_24625,N_14314,N_15763);
xor U24626 (N_24626,N_17055,N_17825);
and U24627 (N_24627,N_14751,N_13714);
nand U24628 (N_24628,N_18733,N_15710);
and U24629 (N_24629,N_17218,N_18491);
and U24630 (N_24630,N_14314,N_17662);
nor U24631 (N_24631,N_16675,N_16049);
xnor U24632 (N_24632,N_18597,N_13154);
xnor U24633 (N_24633,N_17965,N_17011);
and U24634 (N_24634,N_13028,N_13631);
and U24635 (N_24635,N_13349,N_15860);
and U24636 (N_24636,N_14682,N_17954);
xor U24637 (N_24637,N_13291,N_13584);
nand U24638 (N_24638,N_17672,N_17660);
xor U24639 (N_24639,N_16436,N_16211);
nand U24640 (N_24640,N_15849,N_13835);
and U24641 (N_24641,N_15366,N_16438);
and U24642 (N_24642,N_16002,N_15405);
nand U24643 (N_24643,N_18638,N_18734);
nand U24644 (N_24644,N_17544,N_16165);
nor U24645 (N_24645,N_14868,N_18645);
nand U24646 (N_24646,N_17780,N_17371);
nand U24647 (N_24647,N_17620,N_12586);
and U24648 (N_24648,N_17521,N_15039);
or U24649 (N_24649,N_13848,N_13618);
nand U24650 (N_24650,N_17091,N_14810);
xor U24651 (N_24651,N_16974,N_14206);
nand U24652 (N_24652,N_16461,N_17715);
or U24653 (N_24653,N_17332,N_13778);
nand U24654 (N_24654,N_17845,N_16928);
xor U24655 (N_24655,N_14030,N_16908);
or U24656 (N_24656,N_18122,N_15441);
nor U24657 (N_24657,N_17262,N_16308);
or U24658 (N_24658,N_14782,N_16548);
and U24659 (N_24659,N_12887,N_18554);
nand U24660 (N_24660,N_14446,N_17099);
nand U24661 (N_24661,N_13427,N_13277);
nor U24662 (N_24662,N_17863,N_14085);
nor U24663 (N_24663,N_15909,N_15907);
xor U24664 (N_24664,N_16027,N_13288);
nor U24665 (N_24665,N_14668,N_16069);
nand U24666 (N_24666,N_17968,N_16236);
or U24667 (N_24667,N_17592,N_13315);
and U24668 (N_24668,N_18162,N_18242);
and U24669 (N_24669,N_16725,N_16618);
xor U24670 (N_24670,N_18324,N_18745);
and U24671 (N_24671,N_16382,N_16636);
nand U24672 (N_24672,N_16176,N_16006);
xnor U24673 (N_24673,N_17786,N_18015);
and U24674 (N_24674,N_14138,N_13408);
nand U24675 (N_24675,N_13701,N_16624);
nand U24676 (N_24676,N_14863,N_13788);
nand U24677 (N_24677,N_18414,N_17322);
and U24678 (N_24678,N_17116,N_18531);
and U24679 (N_24679,N_17277,N_16730);
nand U24680 (N_24680,N_17635,N_16152);
and U24681 (N_24681,N_13382,N_16465);
nor U24682 (N_24682,N_12994,N_13851);
nor U24683 (N_24683,N_14267,N_13548);
and U24684 (N_24684,N_14665,N_14286);
nand U24685 (N_24685,N_15584,N_15631);
and U24686 (N_24686,N_13574,N_16605);
nor U24687 (N_24687,N_18161,N_15759);
nand U24688 (N_24688,N_16110,N_12650);
xor U24689 (N_24689,N_18722,N_14235);
nand U24690 (N_24690,N_14889,N_13520);
nand U24691 (N_24691,N_17558,N_18676);
or U24692 (N_24692,N_17957,N_13161);
nand U24693 (N_24693,N_18536,N_16480);
nor U24694 (N_24694,N_14832,N_16886);
nor U24695 (N_24695,N_13031,N_14790);
nand U24696 (N_24696,N_15359,N_12845);
nor U24697 (N_24697,N_13346,N_17054);
nor U24698 (N_24698,N_15788,N_14662);
xor U24699 (N_24699,N_18127,N_12746);
and U24700 (N_24700,N_13860,N_13671);
nand U24701 (N_24701,N_15900,N_18025);
xnor U24702 (N_24702,N_12633,N_13551);
and U24703 (N_24703,N_17190,N_18351);
nand U24704 (N_24704,N_18199,N_18003);
nand U24705 (N_24705,N_14496,N_12876);
and U24706 (N_24706,N_17542,N_14640);
and U24707 (N_24707,N_17363,N_14668);
xnor U24708 (N_24708,N_18687,N_17265);
xnor U24709 (N_24709,N_13673,N_12851);
and U24710 (N_24710,N_14303,N_15350);
and U24711 (N_24711,N_12821,N_17849);
nand U24712 (N_24712,N_18451,N_12839);
xnor U24713 (N_24713,N_14649,N_17244);
nor U24714 (N_24714,N_13476,N_15215);
nand U24715 (N_24715,N_13215,N_16703);
nor U24716 (N_24716,N_17710,N_16668);
nand U24717 (N_24717,N_12551,N_17011);
or U24718 (N_24718,N_12931,N_16929);
or U24719 (N_24719,N_16429,N_17220);
nand U24720 (N_24720,N_13108,N_17687);
and U24721 (N_24721,N_16655,N_13221);
nand U24722 (N_24722,N_12596,N_14786);
and U24723 (N_24723,N_15843,N_16770);
or U24724 (N_24724,N_15820,N_17293);
nand U24725 (N_24725,N_16989,N_18693);
xor U24726 (N_24726,N_16115,N_13317);
nand U24727 (N_24727,N_13733,N_16643);
nor U24728 (N_24728,N_16433,N_14318);
nand U24729 (N_24729,N_17099,N_15860);
nand U24730 (N_24730,N_13244,N_17206);
nor U24731 (N_24731,N_13228,N_18228);
and U24732 (N_24732,N_15714,N_14010);
and U24733 (N_24733,N_16638,N_13953);
or U24734 (N_24734,N_18193,N_14944);
or U24735 (N_24735,N_14052,N_14956);
nand U24736 (N_24736,N_15340,N_18542);
nor U24737 (N_24737,N_14249,N_13157);
xnor U24738 (N_24738,N_16700,N_13291);
or U24739 (N_24739,N_13204,N_18388);
or U24740 (N_24740,N_14492,N_14227);
nand U24741 (N_24741,N_15094,N_18253);
and U24742 (N_24742,N_17629,N_18520);
and U24743 (N_24743,N_13666,N_18240);
nand U24744 (N_24744,N_18481,N_12700);
or U24745 (N_24745,N_17207,N_13278);
nor U24746 (N_24746,N_14829,N_14716);
nand U24747 (N_24747,N_12852,N_18422);
or U24748 (N_24748,N_14501,N_15362);
nor U24749 (N_24749,N_13307,N_18274);
nand U24750 (N_24750,N_13079,N_18474);
xnor U24751 (N_24751,N_15936,N_16821);
nand U24752 (N_24752,N_12656,N_13683);
nor U24753 (N_24753,N_15070,N_14194);
nor U24754 (N_24754,N_12706,N_17806);
and U24755 (N_24755,N_18015,N_16582);
nand U24756 (N_24756,N_18588,N_16696);
and U24757 (N_24757,N_14858,N_16092);
and U24758 (N_24758,N_17718,N_16039);
or U24759 (N_24759,N_14756,N_17789);
or U24760 (N_24760,N_13694,N_14782);
and U24761 (N_24761,N_16125,N_18503);
nor U24762 (N_24762,N_17564,N_12687);
and U24763 (N_24763,N_13081,N_14151);
and U24764 (N_24764,N_14542,N_18567);
nand U24765 (N_24765,N_18056,N_18310);
nand U24766 (N_24766,N_13893,N_13915);
xnor U24767 (N_24767,N_13400,N_15199);
nand U24768 (N_24768,N_17968,N_13862);
and U24769 (N_24769,N_12742,N_18717);
nor U24770 (N_24770,N_17355,N_17948);
and U24771 (N_24771,N_14852,N_13844);
or U24772 (N_24772,N_18378,N_17515);
nor U24773 (N_24773,N_15561,N_15775);
nor U24774 (N_24774,N_17586,N_14863);
xnor U24775 (N_24775,N_16287,N_18009);
and U24776 (N_24776,N_15117,N_18365);
nand U24777 (N_24777,N_14551,N_16073);
nand U24778 (N_24778,N_18365,N_13981);
nor U24779 (N_24779,N_15635,N_18374);
and U24780 (N_24780,N_17912,N_15338);
nor U24781 (N_24781,N_14933,N_17930);
nand U24782 (N_24782,N_15657,N_16655);
xor U24783 (N_24783,N_17889,N_15839);
or U24784 (N_24784,N_16393,N_12915);
or U24785 (N_24785,N_14087,N_17310);
xor U24786 (N_24786,N_14948,N_16253);
nand U24787 (N_24787,N_15829,N_14679);
and U24788 (N_24788,N_13276,N_17224);
nor U24789 (N_24789,N_13657,N_17667);
and U24790 (N_24790,N_16355,N_18410);
or U24791 (N_24791,N_17636,N_16903);
or U24792 (N_24792,N_16726,N_12697);
xor U24793 (N_24793,N_13379,N_13822);
nor U24794 (N_24794,N_18505,N_17288);
and U24795 (N_24795,N_13805,N_17996);
and U24796 (N_24796,N_16489,N_13301);
xnor U24797 (N_24797,N_13519,N_18440);
and U24798 (N_24798,N_12805,N_13335);
xor U24799 (N_24799,N_13781,N_17775);
nor U24800 (N_24800,N_18581,N_15326);
xor U24801 (N_24801,N_16977,N_18268);
or U24802 (N_24802,N_17480,N_15304);
or U24803 (N_24803,N_14375,N_18572);
xnor U24804 (N_24804,N_13237,N_14091);
and U24805 (N_24805,N_18609,N_17755);
or U24806 (N_24806,N_15273,N_14879);
nand U24807 (N_24807,N_17585,N_14838);
nand U24808 (N_24808,N_15888,N_18547);
and U24809 (N_24809,N_18125,N_12550);
or U24810 (N_24810,N_16766,N_14406);
nor U24811 (N_24811,N_17733,N_14554);
nand U24812 (N_24812,N_13059,N_18180);
xor U24813 (N_24813,N_15834,N_15783);
and U24814 (N_24814,N_18399,N_12938);
nor U24815 (N_24815,N_15119,N_14973);
xor U24816 (N_24816,N_14630,N_16683);
nand U24817 (N_24817,N_15210,N_16301);
nor U24818 (N_24818,N_14107,N_14504);
and U24819 (N_24819,N_17762,N_18026);
or U24820 (N_24820,N_17933,N_14320);
or U24821 (N_24821,N_14794,N_17821);
and U24822 (N_24822,N_18029,N_13348);
nand U24823 (N_24823,N_14955,N_18288);
xnor U24824 (N_24824,N_18635,N_14181);
and U24825 (N_24825,N_13713,N_14595);
or U24826 (N_24826,N_16002,N_16621);
nor U24827 (N_24827,N_12823,N_13076);
xor U24828 (N_24828,N_17388,N_17021);
and U24829 (N_24829,N_14938,N_18179);
nand U24830 (N_24830,N_17863,N_17701);
and U24831 (N_24831,N_14788,N_14624);
nand U24832 (N_24832,N_16759,N_14181);
xnor U24833 (N_24833,N_15337,N_16117);
nand U24834 (N_24834,N_17828,N_14287);
and U24835 (N_24835,N_12968,N_18091);
xor U24836 (N_24836,N_17386,N_13454);
nor U24837 (N_24837,N_16780,N_12675);
nor U24838 (N_24838,N_18458,N_14091);
nor U24839 (N_24839,N_13567,N_16699);
and U24840 (N_24840,N_14641,N_16686);
and U24841 (N_24841,N_14108,N_13364);
or U24842 (N_24842,N_14537,N_13501);
nor U24843 (N_24843,N_16958,N_14514);
and U24844 (N_24844,N_16384,N_12538);
xor U24845 (N_24845,N_17786,N_16317);
and U24846 (N_24846,N_15290,N_17058);
xor U24847 (N_24847,N_15159,N_13139);
and U24848 (N_24848,N_12562,N_13626);
nor U24849 (N_24849,N_13600,N_15144);
or U24850 (N_24850,N_18254,N_14111);
nand U24851 (N_24851,N_13105,N_13061);
and U24852 (N_24852,N_17749,N_12978);
and U24853 (N_24853,N_15020,N_16247);
or U24854 (N_24854,N_18604,N_15633);
nor U24855 (N_24855,N_13891,N_17316);
nand U24856 (N_24856,N_16611,N_13706);
xor U24857 (N_24857,N_18558,N_16051);
and U24858 (N_24858,N_16564,N_13114);
or U24859 (N_24859,N_13753,N_16990);
nor U24860 (N_24860,N_17086,N_18071);
or U24861 (N_24861,N_18198,N_13409);
nor U24862 (N_24862,N_13210,N_15288);
and U24863 (N_24863,N_17481,N_13136);
and U24864 (N_24864,N_13361,N_13220);
nor U24865 (N_24865,N_15165,N_16907);
and U24866 (N_24866,N_15315,N_13008);
or U24867 (N_24867,N_13778,N_16839);
nand U24868 (N_24868,N_13562,N_12801);
and U24869 (N_24869,N_13037,N_18550);
and U24870 (N_24870,N_17870,N_14269);
nor U24871 (N_24871,N_14491,N_16402);
and U24872 (N_24872,N_16680,N_18116);
nand U24873 (N_24873,N_17045,N_18377);
and U24874 (N_24874,N_15471,N_16407);
nand U24875 (N_24875,N_16616,N_16593);
and U24876 (N_24876,N_17936,N_16039);
or U24877 (N_24877,N_14411,N_17786);
nand U24878 (N_24878,N_17482,N_18482);
xor U24879 (N_24879,N_12899,N_18474);
xor U24880 (N_24880,N_14531,N_18015);
or U24881 (N_24881,N_13093,N_17205);
nand U24882 (N_24882,N_15292,N_17982);
and U24883 (N_24883,N_16521,N_18305);
and U24884 (N_24884,N_12736,N_14544);
nor U24885 (N_24885,N_16849,N_16135);
or U24886 (N_24886,N_17026,N_17547);
and U24887 (N_24887,N_17918,N_15294);
or U24888 (N_24888,N_17518,N_15618);
or U24889 (N_24889,N_18454,N_14191);
nor U24890 (N_24890,N_18740,N_15337);
or U24891 (N_24891,N_17957,N_14323);
xor U24892 (N_24892,N_18201,N_17248);
or U24893 (N_24893,N_13446,N_15974);
nand U24894 (N_24894,N_14770,N_14749);
and U24895 (N_24895,N_18465,N_16774);
and U24896 (N_24896,N_12725,N_18744);
nand U24897 (N_24897,N_13002,N_17433);
and U24898 (N_24898,N_15921,N_16137);
and U24899 (N_24899,N_13929,N_18441);
nor U24900 (N_24900,N_13871,N_15687);
or U24901 (N_24901,N_17042,N_16667);
or U24902 (N_24902,N_14471,N_18296);
nand U24903 (N_24903,N_12702,N_14146);
and U24904 (N_24904,N_17416,N_14272);
nand U24905 (N_24905,N_16263,N_17867);
nor U24906 (N_24906,N_14687,N_14657);
nor U24907 (N_24907,N_18013,N_14276);
xor U24908 (N_24908,N_15664,N_15615);
or U24909 (N_24909,N_13035,N_13353);
nand U24910 (N_24910,N_13236,N_17600);
and U24911 (N_24911,N_13890,N_13411);
nand U24912 (N_24912,N_17246,N_16653);
nor U24913 (N_24913,N_17789,N_13035);
nor U24914 (N_24914,N_16250,N_13507);
or U24915 (N_24915,N_13705,N_16292);
nand U24916 (N_24916,N_15442,N_16845);
xnor U24917 (N_24917,N_14366,N_15369);
nand U24918 (N_24918,N_16148,N_18587);
nand U24919 (N_24919,N_16197,N_17699);
or U24920 (N_24920,N_18421,N_13055);
or U24921 (N_24921,N_16623,N_14881);
xor U24922 (N_24922,N_16106,N_15782);
nor U24923 (N_24923,N_16864,N_15234);
nand U24924 (N_24924,N_13898,N_14793);
nand U24925 (N_24925,N_14361,N_17775);
nor U24926 (N_24926,N_17300,N_18544);
nor U24927 (N_24927,N_16899,N_17145);
xor U24928 (N_24928,N_13087,N_16229);
nor U24929 (N_24929,N_14856,N_14791);
or U24930 (N_24930,N_12778,N_16306);
nor U24931 (N_24931,N_13522,N_15692);
or U24932 (N_24932,N_15310,N_17220);
xor U24933 (N_24933,N_15500,N_14031);
and U24934 (N_24934,N_12676,N_18670);
nand U24935 (N_24935,N_12748,N_18563);
or U24936 (N_24936,N_17741,N_16955);
nand U24937 (N_24937,N_18432,N_13417);
nor U24938 (N_24938,N_13602,N_13151);
xor U24939 (N_24939,N_14690,N_14602);
or U24940 (N_24940,N_14597,N_14810);
nor U24941 (N_24941,N_18012,N_12521);
and U24942 (N_24942,N_13395,N_17985);
and U24943 (N_24943,N_18348,N_15082);
and U24944 (N_24944,N_15599,N_13345);
or U24945 (N_24945,N_12849,N_13143);
nand U24946 (N_24946,N_16970,N_14875);
nand U24947 (N_24947,N_16821,N_14437);
and U24948 (N_24948,N_15421,N_17073);
and U24949 (N_24949,N_12857,N_16142);
nor U24950 (N_24950,N_15915,N_17166);
and U24951 (N_24951,N_15517,N_14020);
nand U24952 (N_24952,N_16818,N_18339);
and U24953 (N_24953,N_13739,N_16317);
nand U24954 (N_24954,N_12572,N_18112);
nor U24955 (N_24955,N_18201,N_16804);
and U24956 (N_24956,N_17060,N_15558);
or U24957 (N_24957,N_12924,N_18639);
nor U24958 (N_24958,N_18234,N_14845);
and U24959 (N_24959,N_18640,N_13385);
or U24960 (N_24960,N_18075,N_16136);
nor U24961 (N_24961,N_12814,N_13441);
or U24962 (N_24962,N_15456,N_12714);
or U24963 (N_24963,N_15202,N_13226);
nor U24964 (N_24964,N_15224,N_16561);
xnor U24965 (N_24965,N_14339,N_14123);
nor U24966 (N_24966,N_15495,N_17813);
nor U24967 (N_24967,N_15244,N_16653);
and U24968 (N_24968,N_17731,N_15420);
or U24969 (N_24969,N_12787,N_16379);
or U24970 (N_24970,N_17664,N_17917);
nand U24971 (N_24971,N_14837,N_13210);
nor U24972 (N_24972,N_17271,N_13064);
nor U24973 (N_24973,N_17538,N_18519);
and U24974 (N_24974,N_17748,N_15154);
nor U24975 (N_24975,N_18450,N_17039);
or U24976 (N_24976,N_15818,N_16865);
xor U24977 (N_24977,N_15583,N_13835);
nor U24978 (N_24978,N_13383,N_18523);
nand U24979 (N_24979,N_16508,N_16867);
nand U24980 (N_24980,N_18008,N_14451);
or U24981 (N_24981,N_14291,N_16935);
nor U24982 (N_24982,N_16615,N_16953);
nor U24983 (N_24983,N_18294,N_17547);
or U24984 (N_24984,N_18579,N_18327);
and U24985 (N_24985,N_18157,N_13513);
and U24986 (N_24986,N_18043,N_16358);
or U24987 (N_24987,N_15226,N_18174);
or U24988 (N_24988,N_16198,N_15644);
nand U24989 (N_24989,N_17449,N_15813);
nand U24990 (N_24990,N_14452,N_14684);
and U24991 (N_24991,N_15647,N_17338);
nor U24992 (N_24992,N_14344,N_17974);
xor U24993 (N_24993,N_15010,N_16846);
nor U24994 (N_24994,N_14115,N_16869);
nor U24995 (N_24995,N_15709,N_17194);
nor U24996 (N_24996,N_18010,N_15683);
or U24997 (N_24997,N_17328,N_14011);
nor U24998 (N_24998,N_14883,N_13002);
and U24999 (N_24999,N_15086,N_13899);
or UO_0 (O_0,N_20714,N_19752);
or UO_1 (O_1,N_24204,N_20112);
and UO_2 (O_2,N_19746,N_20487);
or UO_3 (O_3,N_19683,N_23069);
nor UO_4 (O_4,N_23075,N_23730);
and UO_5 (O_5,N_18917,N_20069);
or UO_6 (O_6,N_22200,N_18923);
nand UO_7 (O_7,N_22057,N_22343);
nand UO_8 (O_8,N_18817,N_21971);
or UO_9 (O_9,N_21191,N_22601);
and UO_10 (O_10,N_21727,N_20799);
nor UO_11 (O_11,N_21333,N_21217);
or UO_12 (O_12,N_20052,N_23007);
nor UO_13 (O_13,N_20746,N_23156);
nor UO_14 (O_14,N_22403,N_23027);
or UO_15 (O_15,N_18919,N_21065);
and UO_16 (O_16,N_19736,N_23187);
or UO_17 (O_17,N_24621,N_19930);
and UO_18 (O_18,N_19399,N_23408);
or UO_19 (O_19,N_22292,N_21218);
or UO_20 (O_20,N_24208,N_21583);
xor UO_21 (O_21,N_20968,N_23029);
nand UO_22 (O_22,N_19065,N_24757);
nor UO_23 (O_23,N_24414,N_20607);
and UO_24 (O_24,N_19138,N_20536);
and UO_25 (O_25,N_24037,N_23948);
nand UO_26 (O_26,N_18865,N_20914);
nand UO_27 (O_27,N_21664,N_20299);
nor UO_28 (O_28,N_19115,N_21617);
or UO_29 (O_29,N_24876,N_23748);
nand UO_30 (O_30,N_20077,N_18932);
nor UO_31 (O_31,N_22071,N_24012);
nor UO_32 (O_32,N_19780,N_23595);
nor UO_33 (O_33,N_20308,N_19617);
nand UO_34 (O_34,N_20220,N_21627);
nand UO_35 (O_35,N_21759,N_23777);
and UO_36 (O_36,N_19969,N_20380);
nand UO_37 (O_37,N_21426,N_21523);
xor UO_38 (O_38,N_23284,N_22198);
or UO_39 (O_39,N_21320,N_23419);
nand UO_40 (O_40,N_19188,N_20849);
nor UO_41 (O_41,N_24633,N_19601);
or UO_42 (O_42,N_24662,N_21927);
nand UO_43 (O_43,N_23165,N_23736);
nor UO_44 (O_44,N_22822,N_22813);
nor UO_45 (O_45,N_19511,N_19095);
and UO_46 (O_46,N_24669,N_23118);
or UO_47 (O_47,N_19184,N_24148);
nand UO_48 (O_48,N_21745,N_23635);
and UO_49 (O_49,N_22969,N_21750);
nor UO_50 (O_50,N_24460,N_24896);
nand UO_51 (O_51,N_21965,N_24030);
nand UO_52 (O_52,N_21298,N_19951);
and UO_53 (O_53,N_20305,N_24438);
nand UO_54 (O_54,N_21033,N_23528);
and UO_55 (O_55,N_21317,N_23105);
nand UO_56 (O_56,N_21060,N_20066);
nand UO_57 (O_57,N_22862,N_20794);
and UO_58 (O_58,N_23906,N_19869);
nand UO_59 (O_59,N_22475,N_19647);
nor UO_60 (O_60,N_21593,N_18765);
and UO_61 (O_61,N_21176,N_21407);
nand UO_62 (O_62,N_21355,N_22283);
nand UO_63 (O_63,N_22157,N_24390);
and UO_64 (O_64,N_22344,N_24888);
or UO_65 (O_65,N_20547,N_22917);
nor UO_66 (O_66,N_22927,N_23471);
nand UO_67 (O_67,N_23117,N_23776);
and UO_68 (O_68,N_22385,N_24128);
and UO_69 (O_69,N_19712,N_24894);
nand UO_70 (O_70,N_22105,N_21113);
nand UO_71 (O_71,N_23751,N_19959);
and UO_72 (O_72,N_19850,N_23895);
nand UO_73 (O_73,N_22471,N_19463);
xor UO_74 (O_74,N_19534,N_20832);
and UO_75 (O_75,N_23110,N_22731);
and UO_76 (O_76,N_20773,N_20784);
and UO_77 (O_77,N_24606,N_23283);
or UO_78 (O_78,N_24651,N_19225);
and UO_79 (O_79,N_23141,N_23641);
nand UO_80 (O_80,N_20336,N_22875);
nor UO_81 (O_81,N_22247,N_22762);
nand UO_82 (O_82,N_19989,N_22237);
or UO_83 (O_83,N_24683,N_21173);
nor UO_84 (O_84,N_24476,N_22557);
nor UO_85 (O_85,N_23220,N_23583);
nand UO_86 (O_86,N_23737,N_23056);
nor UO_87 (O_87,N_23609,N_23098);
nor UO_88 (O_88,N_23249,N_19892);
and UO_89 (O_89,N_19475,N_20423);
or UO_90 (O_90,N_20053,N_21710);
nand UO_91 (O_91,N_24219,N_21536);
or UO_92 (O_92,N_21830,N_21517);
or UO_93 (O_93,N_24825,N_20814);
xor UO_94 (O_94,N_20043,N_23678);
and UO_95 (O_95,N_19057,N_22548);
or UO_96 (O_96,N_21327,N_19323);
and UO_97 (O_97,N_23424,N_20479);
and UO_98 (O_98,N_21474,N_24758);
nand UO_99 (O_99,N_23394,N_22315);
and UO_100 (O_100,N_24268,N_24556);
and UO_101 (O_101,N_21575,N_22698);
and UO_102 (O_102,N_19744,N_19690);
and UO_103 (O_103,N_23959,N_20433);
and UO_104 (O_104,N_19276,N_20242);
xor UO_105 (O_105,N_22400,N_21243);
or UO_106 (O_106,N_24631,N_21085);
and UO_107 (O_107,N_20939,N_19902);
or UO_108 (O_108,N_21364,N_23778);
and UO_109 (O_109,N_22324,N_22345);
nor UO_110 (O_110,N_20218,N_19564);
nor UO_111 (O_111,N_18750,N_19049);
or UO_112 (O_112,N_21799,N_20994);
and UO_113 (O_113,N_19351,N_24347);
nor UO_114 (O_114,N_19470,N_24277);
xor UO_115 (O_115,N_22778,N_24750);
nor UO_116 (O_116,N_19460,N_21852);
and UO_117 (O_117,N_24361,N_22236);
nor UO_118 (O_118,N_24023,N_23236);
and UO_119 (O_119,N_23252,N_21313);
or UO_120 (O_120,N_21335,N_23083);
nor UO_121 (O_121,N_19195,N_22387);
nand UO_122 (O_122,N_24906,N_23649);
nor UO_123 (O_123,N_19749,N_23209);
and UO_124 (O_124,N_19753,N_22188);
nand UO_125 (O_125,N_21239,N_23500);
or UO_126 (O_126,N_21299,N_20734);
and UO_127 (O_127,N_19334,N_24930);
nor UO_128 (O_128,N_21270,N_19888);
nand UO_129 (O_129,N_20504,N_20241);
and UO_130 (O_130,N_22162,N_22456);
and UO_131 (O_131,N_22826,N_21637);
nand UO_132 (O_132,N_21418,N_22679);
nor UO_133 (O_133,N_22375,N_19603);
and UO_134 (O_134,N_19200,N_21214);
nand UO_135 (O_135,N_21509,N_24063);
or UO_136 (O_136,N_24837,N_19354);
nor UO_137 (O_137,N_22141,N_22242);
nor UO_138 (O_138,N_24922,N_19359);
or UO_139 (O_139,N_22608,N_18853);
or UO_140 (O_140,N_20376,N_19238);
or UO_141 (O_141,N_20127,N_24742);
and UO_142 (O_142,N_23967,N_18790);
nand UO_143 (O_143,N_23227,N_21230);
and UO_144 (O_144,N_22795,N_20749);
and UO_145 (O_145,N_23484,N_19838);
nand UO_146 (O_146,N_22463,N_21223);
nand UO_147 (O_147,N_22244,N_19536);
nor UO_148 (O_148,N_20712,N_22876);
and UO_149 (O_149,N_21700,N_19010);
or UO_150 (O_150,N_24514,N_19980);
and UO_151 (O_151,N_23046,N_22542);
or UO_152 (O_152,N_24425,N_23816);
and UO_153 (O_153,N_20475,N_21045);
nor UO_154 (O_154,N_20330,N_19222);
nor UO_155 (O_155,N_22058,N_24415);
nand UO_156 (O_156,N_21224,N_22089);
nand UO_157 (O_157,N_20103,N_22154);
nand UO_158 (O_158,N_23501,N_22765);
or UO_159 (O_159,N_23675,N_22081);
nor UO_160 (O_160,N_18757,N_20196);
nor UO_161 (O_161,N_21374,N_24617);
or UO_162 (O_162,N_19551,N_19061);
nand UO_163 (O_163,N_21978,N_23302);
and UO_164 (O_164,N_19429,N_20611);
or UO_165 (O_165,N_19447,N_20012);
nor UO_166 (O_166,N_21932,N_20016);
and UO_167 (O_167,N_20115,N_21164);
and UO_168 (O_168,N_22352,N_20454);
or UO_169 (O_169,N_24459,N_21018);
or UO_170 (O_170,N_21434,N_20055);
xor UO_171 (O_171,N_23604,N_18986);
nor UO_172 (O_172,N_20206,N_20616);
xnor UO_173 (O_173,N_21987,N_20544);
nand UO_174 (O_174,N_21263,N_21849);
nand UO_175 (O_175,N_23971,N_23341);
nand UO_176 (O_176,N_21135,N_23093);
or UO_177 (O_177,N_22570,N_18949);
xor UO_178 (O_178,N_22147,N_23329);
and UO_179 (O_179,N_19609,N_22069);
and UO_180 (O_180,N_22335,N_23063);
nand UO_181 (O_181,N_22026,N_22811);
or UO_182 (O_182,N_23181,N_20062);
nand UO_183 (O_183,N_24871,N_24777);
and UO_184 (O_184,N_21545,N_24635);
xnor UO_185 (O_185,N_23089,N_21560);
nand UO_186 (O_186,N_22368,N_24049);
nor UO_187 (O_187,N_23290,N_23812);
nand UO_188 (O_188,N_21826,N_22912);
nand UO_189 (O_189,N_21737,N_19881);
nand UO_190 (O_190,N_22593,N_22836);
nor UO_191 (O_191,N_24565,N_20645);
or UO_192 (O_192,N_21543,N_20343);
xor UO_193 (O_193,N_19678,N_22134);
nand UO_194 (O_194,N_23418,N_24566);
nor UO_195 (O_195,N_23712,N_21010);
and UO_196 (O_196,N_21557,N_23799);
nor UO_197 (O_197,N_19730,N_19080);
or UO_198 (O_198,N_23710,N_23946);
nand UO_199 (O_199,N_20687,N_22202);
and UO_200 (O_200,N_23828,N_21151);
nand UO_201 (O_201,N_22043,N_19866);
nor UO_202 (O_202,N_24103,N_18925);
xnor UO_203 (O_203,N_22156,N_20233);
nor UO_204 (O_204,N_20576,N_21579);
and UO_205 (O_205,N_19229,N_21207);
and UO_206 (O_206,N_19374,N_23880);
xor UO_207 (O_207,N_23041,N_21665);
nor UO_208 (O_208,N_20665,N_24122);
xnor UO_209 (O_209,N_19607,N_18997);
nand UO_210 (O_210,N_22587,N_20523);
or UO_211 (O_211,N_23771,N_24674);
nand UO_212 (O_212,N_24144,N_20800);
nor UO_213 (O_213,N_23877,N_21953);
nor UO_214 (O_214,N_20011,N_24769);
or UO_215 (O_215,N_23718,N_22068);
nor UO_216 (O_216,N_20867,N_19788);
nor UO_217 (O_217,N_24601,N_24223);
nor UO_218 (O_218,N_22524,N_19649);
or UO_219 (O_219,N_19360,N_24948);
and UO_220 (O_220,N_22700,N_19885);
and UO_221 (O_221,N_21741,N_22351);
nand UO_222 (O_222,N_21205,N_24504);
xnor UO_223 (O_223,N_22021,N_20182);
or UO_224 (O_224,N_22295,N_19908);
and UO_225 (O_225,N_20561,N_22824);
nor UO_226 (O_226,N_21316,N_23904);
nand UO_227 (O_227,N_24340,N_21247);
or UO_228 (O_228,N_23147,N_22361);
nor UO_229 (O_229,N_18764,N_20930);
nand UO_230 (O_230,N_24630,N_23783);
and UO_231 (O_231,N_23891,N_22753);
nor UO_232 (O_232,N_23473,N_24234);
nor UO_233 (O_233,N_19365,N_19146);
nand UO_234 (O_234,N_20642,N_23930);
or UO_235 (O_235,N_20880,N_22033);
or UO_236 (O_236,N_24105,N_20562);
nand UO_237 (O_237,N_21376,N_22281);
or UO_238 (O_238,N_20201,N_20435);
or UO_239 (O_239,N_20093,N_24279);
and UO_240 (O_240,N_21213,N_24066);
nand UO_241 (O_241,N_19269,N_24790);
or UO_242 (O_242,N_20097,N_19471);
nor UO_243 (O_243,N_22533,N_24952);
nor UO_244 (O_244,N_20662,N_20686);
nand UO_245 (O_245,N_23305,N_24690);
and UO_246 (O_246,N_20884,N_23177);
nor UO_247 (O_247,N_23740,N_19362);
nand UO_248 (O_248,N_24907,N_21489);
and UO_249 (O_249,N_20728,N_20168);
nor UO_250 (O_250,N_23131,N_23317);
or UO_251 (O_251,N_23690,N_23988);
and UO_252 (O_252,N_18948,N_24130);
and UO_253 (O_253,N_21469,N_22946);
or UO_254 (O_254,N_22092,N_20854);
nor UO_255 (O_255,N_20322,N_22558);
nor UO_256 (O_256,N_19762,N_20946);
and UO_257 (O_257,N_22590,N_23049);
or UO_258 (O_258,N_21133,N_20223);
xor UO_259 (O_259,N_21793,N_22279);
and UO_260 (O_260,N_23065,N_20422);
or UO_261 (O_261,N_22660,N_23493);
and UO_262 (O_262,N_21834,N_22851);
nand UO_263 (O_263,N_21858,N_23239);
and UO_264 (O_264,N_23703,N_21656);
and UO_265 (O_265,N_19427,N_20643);
nor UO_266 (O_266,N_21502,N_24508);
and UO_267 (O_267,N_21901,N_23092);
nand UO_268 (O_268,N_23003,N_23100);
and UO_269 (O_269,N_19262,N_21859);
and UO_270 (O_270,N_24549,N_24588);
xor UO_271 (O_271,N_24868,N_24120);
xor UO_272 (O_272,N_19003,N_23786);
nand UO_273 (O_273,N_21920,N_23992);
xor UO_274 (O_274,N_20264,N_22887);
nand UO_275 (O_275,N_21780,N_20154);
or UO_276 (O_276,N_22234,N_20222);
xnor UO_277 (O_277,N_22790,N_23307);
or UO_278 (O_278,N_22757,N_19940);
or UO_279 (O_279,N_19986,N_19270);
and UO_280 (O_280,N_24110,N_24127);
and UO_281 (O_281,N_23143,N_22665);
and UO_282 (O_282,N_20042,N_21492);
or UO_283 (O_283,N_21401,N_20989);
nor UO_284 (O_284,N_21014,N_20636);
nor UO_285 (O_285,N_22829,N_22846);
or UO_286 (O_286,N_20882,N_18892);
nand UO_287 (O_287,N_20088,N_24131);
and UO_288 (O_288,N_22818,N_24041);
xnor UO_289 (O_289,N_23939,N_24681);
nand UO_290 (O_290,N_21857,N_21928);
nand UO_291 (O_291,N_22952,N_19757);
and UO_292 (O_292,N_21378,N_24248);
xor UO_293 (O_293,N_20948,N_21605);
and UO_294 (O_294,N_19593,N_19535);
or UO_295 (O_295,N_20837,N_19805);
nand UO_296 (O_296,N_20270,N_23689);
nor UO_297 (O_297,N_22775,N_24736);
nand UO_298 (O_298,N_19274,N_21459);
xnor UO_299 (O_299,N_20740,N_20213);
and UO_300 (O_300,N_19512,N_21360);
or UO_301 (O_301,N_21359,N_22699);
xnor UO_302 (O_302,N_23983,N_24691);
and UO_303 (O_303,N_24490,N_22615);
and UO_304 (O_304,N_20683,N_20952);
nand UO_305 (O_305,N_24119,N_22366);
or UO_306 (O_306,N_18784,N_19926);
nand UO_307 (O_307,N_19679,N_24335);
nand UO_308 (O_308,N_24656,N_24387);
and UO_309 (O_309,N_19209,N_21069);
nand UO_310 (O_310,N_20742,N_23134);
or UO_311 (O_311,N_20410,N_22937);
nor UO_312 (O_312,N_19106,N_20263);
nand UO_313 (O_313,N_20278,N_23374);
and UO_314 (O_314,N_23403,N_20160);
nand UO_315 (O_315,N_19456,N_19178);
xnor UO_316 (O_316,N_24336,N_19469);
and UO_317 (O_317,N_21311,N_20731);
xnor UO_318 (O_318,N_18929,N_20887);
nor UO_319 (O_319,N_19112,N_24190);
nor UO_320 (O_320,N_22730,N_22951);
nor UO_321 (O_321,N_19592,N_23504);
and UO_322 (O_322,N_19978,N_23232);
nand UO_323 (O_323,N_24174,N_22987);
or UO_324 (O_324,N_22502,N_21382);
or UO_325 (O_325,N_22310,N_20889);
nor UO_326 (O_326,N_23045,N_20477);
and UO_327 (O_327,N_19473,N_20426);
and UO_328 (O_328,N_19711,N_19819);
and UO_329 (O_329,N_22497,N_19890);
nand UO_330 (O_330,N_24269,N_21292);
or UO_331 (O_331,N_21400,N_20723);
or UO_332 (O_332,N_23381,N_22055);
and UO_333 (O_333,N_22493,N_22461);
nand UO_334 (O_334,N_24618,N_22773);
nand UO_335 (O_335,N_19085,N_24975);
or UO_336 (O_336,N_23086,N_21094);
xor UO_337 (O_337,N_23468,N_23598);
xor UO_338 (O_338,N_20720,N_19030);
xnor UO_339 (O_339,N_22135,N_19402);
nand UO_340 (O_340,N_22374,N_21861);
nor UO_341 (O_341,N_19719,N_24983);
nand UO_342 (O_342,N_19656,N_19944);
nand UO_343 (O_343,N_21450,N_20176);
and UO_344 (O_344,N_20214,N_23763);
nand UO_345 (O_345,N_20071,N_24233);
or UO_346 (O_346,N_21647,N_22733);
xor UO_347 (O_347,N_24530,N_22285);
nor UO_348 (O_348,N_23565,N_20653);
and UO_349 (O_349,N_24467,N_21676);
and UO_350 (O_350,N_20092,N_24480);
nand UO_351 (O_351,N_24659,N_20838);
nor UO_352 (O_352,N_22563,N_23330);
xnor UO_353 (O_353,N_24173,N_22238);
nor UO_354 (O_354,N_21451,N_23995);
and UO_355 (O_355,N_23961,N_23130);
xnor UO_356 (O_356,N_23132,N_21200);
and UO_357 (O_357,N_19221,N_21597);
nor UO_358 (O_358,N_22776,N_23261);
nand UO_359 (O_359,N_22977,N_21673);
and UO_360 (O_360,N_24774,N_18804);
or UO_361 (O_361,N_21332,N_24360);
and UO_362 (O_362,N_18874,N_20638);
nand UO_363 (O_363,N_23673,N_20979);
and UO_364 (O_364,N_24011,N_24661);
or UO_365 (O_365,N_24892,N_19130);
and UO_366 (O_366,N_23052,N_21309);
nand UO_367 (O_367,N_21357,N_18939);
nor UO_368 (O_368,N_19194,N_19499);
or UO_369 (O_369,N_21348,N_21833);
or UO_370 (O_370,N_22627,N_21630);
nor UO_371 (O_371,N_21267,N_20312);
and UO_372 (O_372,N_20896,N_23681);
and UO_373 (O_373,N_21611,N_19828);
and UO_374 (O_374,N_19979,N_23701);
and UO_375 (O_375,N_19637,N_21437);
or UO_376 (O_376,N_24596,N_24872);
nand UO_377 (O_377,N_20186,N_24629);
nor UO_378 (O_378,N_23300,N_24961);
or UO_379 (O_379,N_22536,N_19038);
nor UO_380 (O_380,N_20462,N_19949);
nor UO_381 (O_381,N_19830,N_20424);
nor UO_382 (O_382,N_23004,N_24838);
nand UO_383 (O_383,N_23514,N_20689);
nand UO_384 (O_384,N_20370,N_22713);
nand UO_385 (O_385,N_24881,N_21513);
xnor UO_386 (O_386,N_19801,N_20598);
and UO_387 (O_387,N_24400,N_20879);
and UO_388 (O_388,N_24735,N_24739);
nor UO_389 (O_389,N_19661,N_21943);
and UO_390 (O_390,N_23533,N_24473);
and UO_391 (O_391,N_21421,N_19345);
or UO_392 (O_392,N_19305,N_20126);
nor UO_393 (O_393,N_21913,N_21758);
and UO_394 (O_394,N_22488,N_23759);
xnor UO_395 (O_395,N_22327,N_18773);
nor UO_396 (O_396,N_22769,N_21508);
and UO_397 (O_397,N_24314,N_21442);
nand UO_398 (O_398,N_24007,N_23670);
or UO_399 (O_399,N_22933,N_24501);
or UO_400 (O_400,N_23125,N_19741);
nor UO_401 (O_401,N_22926,N_20904);
and UO_402 (O_402,N_20005,N_22803);
or UO_403 (O_403,N_20592,N_22208);
nand UO_404 (O_404,N_19822,N_21540);
nor UO_405 (O_405,N_24727,N_20812);
or UO_406 (O_406,N_24502,N_20828);
nor UO_407 (O_407,N_23372,N_23756);
nand UO_408 (O_408,N_19862,N_20783);
xnor UO_409 (O_409,N_21340,N_23588);
nor UO_410 (O_410,N_23270,N_22985);
or UO_411 (O_411,N_19646,N_18852);
nor UO_412 (O_412,N_22336,N_20219);
nand UO_413 (O_413,N_19787,N_21417);
or UO_414 (O_414,N_21137,N_24577);
nand UO_415 (O_415,N_20709,N_22175);
and UO_416 (O_416,N_20318,N_21763);
nand UO_417 (O_417,N_19074,N_21628);
and UO_418 (O_418,N_21643,N_22353);
or UO_419 (O_419,N_20418,N_19379);
nand UO_420 (O_420,N_20587,N_22392);
and UO_421 (O_421,N_19504,N_18943);
or UO_422 (O_422,N_24116,N_19595);
and UO_423 (O_423,N_21271,N_19616);
nor UO_424 (O_424,N_20679,N_23656);
nor UO_425 (O_425,N_21169,N_19439);
nor UO_426 (O_426,N_23121,N_21550);
and UO_427 (O_427,N_19383,N_22280);
or UO_428 (O_428,N_23162,N_19449);
or UO_429 (O_429,N_24334,N_21435);
and UO_430 (O_430,N_23507,N_23070);
and UO_431 (O_431,N_19956,N_20132);
nand UO_432 (O_432,N_20770,N_19925);
or UO_433 (O_433,N_20265,N_20624);
and UO_434 (O_434,N_24230,N_24099);
nor UO_435 (O_435,N_20191,N_24937);
nor UO_436 (O_436,N_24442,N_19966);
nor UO_437 (O_437,N_24283,N_24404);
nor UO_438 (O_438,N_19059,N_24026);
nand UO_439 (O_439,N_22265,N_19281);
xor UO_440 (O_440,N_21306,N_22715);
and UO_441 (O_441,N_20341,N_20925);
nand UO_442 (O_442,N_20399,N_19101);
nand UO_443 (O_443,N_23022,N_19489);
and UO_444 (O_444,N_20471,N_23139);
nor UO_445 (O_445,N_19620,N_20409);
or UO_446 (O_446,N_21093,N_18785);
or UO_447 (O_447,N_24734,N_20025);
nand UO_448 (O_448,N_19555,N_23426);
or UO_449 (O_449,N_20951,N_24005);
nor UO_450 (O_450,N_19437,N_22095);
and UO_451 (O_451,N_24196,N_24798);
xnor UO_452 (O_452,N_19322,N_21925);
nand UO_453 (O_453,N_19834,N_21968);
and UO_454 (O_454,N_21206,N_24959);
xnor UO_455 (O_455,N_20795,N_23957);
nor UO_456 (O_456,N_22203,N_23950);
or UO_457 (O_457,N_23437,N_19955);
and UO_458 (O_458,N_21918,N_21527);
and UO_459 (O_459,N_20374,N_20569);
and UO_460 (O_460,N_24216,N_23286);
or UO_461 (O_461,N_22342,N_19910);
and UO_462 (O_462,N_19267,N_19199);
nor UO_463 (O_463,N_23519,N_22300);
nand UO_464 (O_464,N_18944,N_19053);
nor UO_465 (O_465,N_20648,N_20021);
nor UO_466 (O_466,N_23407,N_22477);
and UO_467 (O_467,N_24600,N_20497);
or UO_468 (O_468,N_24371,N_19675);
nor UO_469 (O_469,N_22535,N_23151);
nor UO_470 (O_470,N_21037,N_19018);
and UO_471 (O_471,N_20086,N_19035);
and UO_472 (O_472,N_24315,N_19825);
and UO_473 (O_473,N_24698,N_24285);
or UO_474 (O_474,N_21017,N_22064);
nand UO_475 (O_475,N_20906,N_23862);
nand UO_476 (O_476,N_19230,N_21368);
nor UO_477 (O_477,N_19696,N_19873);
nor UO_478 (O_478,N_23900,N_19538);
and UO_479 (O_479,N_24579,N_21095);
or UO_480 (O_480,N_22381,N_22696);
nor UO_481 (O_481,N_22891,N_23886);
nand UO_482 (O_482,N_21850,N_18837);
and UO_483 (O_483,N_21250,N_21251);
nand UO_484 (O_484,N_22522,N_24312);
nor UO_485 (O_485,N_18862,N_24582);
or UO_486 (O_486,N_19159,N_21020);
or UO_487 (O_487,N_22894,N_23927);
nand UO_488 (O_488,N_24036,N_23137);
and UO_489 (O_489,N_21244,N_23590);
nor UO_490 (O_490,N_24353,N_19062);
nor UO_491 (O_491,N_24499,N_22636);
and UO_492 (O_492,N_20581,N_21089);
nand UO_493 (O_493,N_20164,N_19371);
xnor UO_494 (O_494,N_20572,N_21580);
nand UO_495 (O_495,N_24008,N_20626);
nor UO_496 (O_496,N_19915,N_24465);
or UO_497 (O_497,N_19490,N_21854);
or UO_498 (O_498,N_22308,N_23911);
or UO_499 (O_499,N_21929,N_24278);
xor UO_500 (O_500,N_19196,N_20987);
and UO_501 (O_501,N_21687,N_21013);
nor UO_502 (O_502,N_18876,N_18888);
or UO_503 (O_503,N_19911,N_19933);
nand UO_504 (O_504,N_22323,N_21672);
and UO_505 (O_505,N_21875,N_19135);
xnor UO_506 (O_506,N_22272,N_19275);
or UO_507 (O_507,N_20524,N_23765);
nor UO_508 (O_508,N_24187,N_22859);
and UO_509 (O_509,N_19476,N_24802);
and UO_510 (O_510,N_20649,N_22847);
nand UO_511 (O_511,N_21003,N_23617);
nor UO_512 (O_512,N_23191,N_21369);
nand UO_513 (O_513,N_18971,N_24432);
nor UO_514 (O_514,N_19895,N_19558);
nor UO_515 (O_515,N_19879,N_22277);
nor UO_516 (O_516,N_24725,N_24967);
nand UO_517 (O_517,N_18793,N_23859);
nand UO_518 (O_518,N_24455,N_19000);
nor UO_519 (O_519,N_19820,N_22519);
nand UO_520 (O_520,N_22594,N_21996);
and UO_521 (O_521,N_21118,N_21768);
and UO_522 (O_522,N_24383,N_22761);
xor UO_523 (O_523,N_19265,N_21428);
and UO_524 (O_524,N_20815,N_23970);
nand UO_525 (O_525,N_23242,N_21804);
nor UO_526 (O_526,N_24358,N_24226);
or UO_527 (O_527,N_19303,N_22384);
and UO_528 (O_528,N_22298,N_18845);
xor UO_529 (O_529,N_20185,N_23033);
nand UO_530 (O_530,N_24391,N_20027);
or UO_531 (O_531,N_24274,N_21386);
nand UO_532 (O_532,N_18782,N_23592);
and UO_533 (O_533,N_19798,N_23578);
or UO_534 (O_534,N_20589,N_20333);
xor UO_535 (O_535,N_19293,N_21797);
nand UO_536 (O_536,N_19784,N_23219);
nor UO_537 (O_537,N_20175,N_23016);
nor UO_538 (O_538,N_24960,N_20873);
or UO_539 (O_539,N_22348,N_20140);
or UO_540 (O_540,N_20963,N_19457);
and UO_541 (O_541,N_22890,N_19483);
nor UO_542 (O_542,N_24028,N_24109);
nor UO_543 (O_543,N_21577,N_19356);
nand UO_544 (O_544,N_23572,N_23485);
nor UO_545 (O_545,N_20997,N_20375);
or UO_546 (O_546,N_22334,N_21939);
nand UO_547 (O_547,N_21002,N_22802);
and UO_548 (O_548,N_19190,N_20104);
or UO_549 (O_549,N_22062,N_21454);
nor UO_550 (O_550,N_22693,N_20358);
or UO_551 (O_551,N_22127,N_19168);
or UO_552 (O_552,N_24828,N_24150);
or UO_553 (O_553,N_20959,N_23258);
or UO_554 (O_554,N_20284,N_19211);
nand UO_555 (O_555,N_23265,N_22578);
nor UO_556 (O_556,N_20384,N_19676);
or UO_557 (O_557,N_19508,N_23923);
and UO_558 (O_558,N_20147,N_24949);
or UO_559 (O_559,N_20517,N_20179);
or UO_560 (O_560,N_23412,N_24715);
xor UO_561 (O_561,N_21977,N_21096);
or UO_562 (O_562,N_20508,N_22740);
or UO_563 (O_563,N_23082,N_23753);
nor UO_564 (O_564,N_21189,N_20252);
nor UO_565 (O_565,N_19170,N_24550);
or UO_566 (O_566,N_24847,N_22856);
and UO_567 (O_567,N_21680,N_21049);
or UO_568 (O_568,N_22426,N_24981);
or UO_569 (O_569,N_23179,N_21234);
or UO_570 (O_570,N_20216,N_18870);
or UO_571 (O_571,N_22562,N_21078);
or UO_572 (O_572,N_21044,N_24970);
and UO_573 (O_573,N_24914,N_18755);
nor UO_574 (O_574,N_22148,N_22137);
nor UO_575 (O_575,N_21805,N_22701);
or UO_576 (O_576,N_22122,N_24700);
and UO_577 (O_577,N_22464,N_23400);
nor UO_578 (O_578,N_20037,N_21246);
or UO_579 (O_579,N_21088,N_24319);
nor UO_580 (O_580,N_24220,N_21958);
nand UO_581 (O_581,N_24263,N_24421);
or UO_582 (O_582,N_21116,N_20516);
or UO_583 (O_583,N_19430,N_23491);
nor UO_584 (O_584,N_20232,N_19081);
or UO_585 (O_585,N_22663,N_22642);
nor UO_586 (O_586,N_22404,N_18936);
and UO_587 (O_587,N_21381,N_19765);
nand UO_588 (O_588,N_23685,N_22339);
and UO_589 (O_589,N_19405,N_24147);
and UO_590 (O_590,N_23199,N_23411);
xnor UO_591 (O_591,N_22868,N_18947);
nor UO_592 (O_592,N_19991,N_24607);
or UO_593 (O_593,N_20688,N_20067);
xor UO_594 (O_594,N_19677,N_22666);
nand UO_595 (O_595,N_19826,N_19549);
or UO_596 (O_596,N_24295,N_22409);
nand UO_597 (O_597,N_24747,N_23858);
nor UO_598 (O_598,N_22899,N_22632);
and UO_599 (O_599,N_20594,N_20548);
or UO_600 (O_600,N_24273,N_21114);
and UO_601 (O_601,N_18995,N_21934);
and UO_602 (O_602,N_19810,N_21423);
nand UO_603 (O_603,N_24932,N_22936);
and UO_604 (O_604,N_19735,N_23230);
or UO_605 (O_605,N_23054,N_18752);
and UO_606 (O_606,N_22329,N_19527);
nand UO_607 (O_607,N_23116,N_22395);
and UO_608 (O_608,N_22910,N_21101);
or UO_609 (O_609,N_23650,N_21649);
and UO_610 (O_610,N_20924,N_18957);
xnor UO_611 (O_611,N_22180,N_18871);
nand UO_612 (O_612,N_21329,N_22433);
xor UO_613 (O_613,N_21501,N_21608);
or UO_614 (O_614,N_23969,N_24753);
or UO_615 (O_615,N_22844,N_20448);
and UO_616 (O_616,N_21194,N_21068);
nor UO_617 (O_617,N_20796,N_23562);
xor UO_618 (O_618,N_21353,N_24716);
or UO_619 (O_619,N_22144,N_23413);
nand UO_620 (O_620,N_19468,N_23809);
and UO_621 (O_621,N_22585,N_23461);
nand UO_622 (O_622,N_18859,N_21462);
nand UO_623 (O_623,N_24010,N_23463);
and UO_624 (O_624,N_21457,N_21827);
and UO_625 (O_625,N_24664,N_21757);
and UO_626 (O_626,N_22121,N_20116);
nand UO_627 (O_627,N_21781,N_22087);
nand UO_628 (O_628,N_21526,N_21258);
nor UO_629 (O_629,N_20353,N_19698);
nand UO_630 (O_630,N_22831,N_19836);
nor UO_631 (O_631,N_24841,N_19342);
nand UO_632 (O_632,N_22223,N_21890);
or UO_633 (O_633,N_23289,N_22160);
or UO_634 (O_634,N_18907,N_23154);
and UO_635 (O_635,N_20009,N_22512);
nor UO_636 (O_636,N_19248,N_23316);
xor UO_637 (O_637,N_24589,N_19353);
xor UO_638 (O_638,N_20273,N_21008);
and UO_639 (O_639,N_24627,N_24991);
nand UO_640 (O_640,N_19854,N_19807);
and UO_641 (O_641,N_22388,N_22569);
nor UO_642 (O_642,N_21648,N_23306);
and UO_643 (O_643,N_19522,N_19939);
nor UO_644 (O_644,N_20455,N_22618);
nand UO_645 (O_645,N_23795,N_23457);
and UO_646 (O_646,N_19425,N_23944);
nor UO_647 (O_647,N_20184,N_24832);
nand UO_648 (O_648,N_24343,N_21175);
nand UO_649 (O_649,N_22186,N_22798);
and UO_650 (O_650,N_20654,N_19177);
or UO_651 (O_651,N_18920,N_22800);
nor UO_652 (O_652,N_21172,N_18826);
nand UO_653 (O_653,N_19660,N_19546);
nand UO_654 (O_654,N_20427,N_21475);
or UO_655 (O_655,N_19068,N_22495);
or UO_656 (O_656,N_19414,N_19935);
nor UO_657 (O_657,N_20839,N_22346);
or UO_658 (O_658,N_22107,N_19576);
nand UO_659 (O_659,N_23466,N_24197);
or UO_660 (O_660,N_24489,N_18847);
and UO_661 (O_661,N_24377,N_21227);
nor UO_662 (O_662,N_20236,N_20151);
nor UO_663 (O_663,N_22136,N_20923);
xnor UO_664 (O_664,N_22637,N_24094);
nor UO_665 (O_665,N_21158,N_23356);
xnor UO_666 (O_666,N_19153,N_20927);
xnor UO_667 (O_667,N_18946,N_22001);
nor UO_668 (O_668,N_20802,N_24016);
and UO_669 (O_669,N_24513,N_22881);
or UO_670 (O_670,N_19385,N_20338);
and UO_671 (O_671,N_20733,N_21744);
or UO_672 (O_672,N_23871,N_19604);
and UO_673 (O_673,N_19307,N_20543);
or UO_674 (O_674,N_20910,N_21219);
xor UO_675 (O_675,N_22934,N_23280);
xnor UO_676 (O_676,N_19396,N_23563);
or UO_677 (O_677,N_19495,N_19662);
and UO_678 (O_678,N_24644,N_22720);
or UO_679 (O_679,N_22705,N_22918);
nor UO_680 (O_680,N_23028,N_19975);
nor UO_681 (O_681,N_24839,N_19545);
nor UO_682 (O_682,N_22580,N_20897);
nand UO_683 (O_683,N_23920,N_22340);
nor UO_684 (O_684,N_19540,N_24142);
and UO_685 (O_685,N_22774,N_22786);
or UO_686 (O_686,N_24982,N_22362);
nor UO_687 (O_687,N_20736,N_19277);
nor UO_688 (O_688,N_23477,N_22997);
xnor UO_689 (O_689,N_19117,N_19710);
xor UO_690 (O_690,N_23531,N_21035);
or UO_691 (O_691,N_21504,N_19845);
or UO_692 (O_692,N_24305,N_20443);
nor UO_693 (O_693,N_21099,N_23148);
or UO_694 (O_694,N_23326,N_23106);
nand UO_695 (O_695,N_21872,N_22956);
nor UO_696 (O_696,N_22165,N_22904);
and UO_697 (O_697,N_21180,N_22419);
and UO_698 (O_698,N_19621,N_18879);
and UO_699 (O_699,N_19723,N_19652);
or UO_700 (O_700,N_24355,N_22613);
or UO_701 (O_701,N_23585,N_20459);
xnor UO_702 (O_702,N_22290,N_21422);
and UO_703 (O_703,N_22142,N_22022);
and UO_704 (O_704,N_22976,N_19877);
and UO_705 (O_705,N_21772,N_22586);
nor UO_706 (O_706,N_19121,N_23766);
nor UO_707 (O_707,N_20018,N_22664);
xor UO_708 (O_708,N_19441,N_21149);
and UO_709 (O_709,N_19290,N_19648);
and UO_710 (O_710,N_23527,N_22116);
nor UO_711 (O_711,N_22301,N_20875);
nand UO_712 (O_712,N_21392,N_24272);
nor UO_713 (O_713,N_20248,N_20442);
nand UO_714 (O_714,N_19250,N_22755);
nand UO_715 (O_715,N_21375,N_24412);
or UO_716 (O_716,N_21699,N_21873);
or UO_717 (O_717,N_20325,N_20657);
or UO_718 (O_718,N_22504,N_24449);
nor UO_719 (O_719,N_21638,N_22044);
nand UO_720 (O_720,N_22897,N_20342);
xor UO_721 (O_721,N_19800,N_21592);
and UO_722 (O_722,N_22779,N_22115);
nand UO_723 (O_723,N_24924,N_21838);
and UO_724 (O_724,N_22743,N_22226);
nand UO_725 (O_725,N_22748,N_22595);
or UO_726 (O_726,N_21245,N_19972);
nor UO_727 (O_727,N_22389,N_19321);
or UO_728 (O_728,N_23094,N_20710);
nor UO_729 (O_729,N_24240,N_24297);
nor UO_730 (O_730,N_23818,N_24349);
nor UO_731 (O_731,N_23439,N_20143);
nor UO_732 (O_732,N_21097,N_19131);
nand UO_733 (O_733,N_20673,N_22791);
xnor UO_734 (O_734,N_22643,N_19169);
and UO_735 (O_735,N_23813,N_23299);
nand UO_736 (O_736,N_23580,N_21521);
and UO_737 (O_737,N_23523,N_23458);
or UO_738 (O_738,N_20357,N_22688);
or UO_739 (O_739,N_24214,N_24956);
nand UO_740 (O_740,N_20274,N_21972);
or UO_741 (O_741,N_19006,N_21198);
nand UO_742 (O_742,N_24517,N_23746);
or UO_743 (O_743,N_23126,N_23168);
nand UO_744 (O_744,N_19500,N_24702);
and UO_745 (O_745,N_23570,N_20056);
xor UO_746 (O_746,N_20489,N_22870);
nand UO_747 (O_747,N_21066,N_21651);
and UO_748 (O_748,N_23925,N_19843);
nor UO_749 (O_749,N_21921,N_23719);
and UO_750 (O_750,N_24902,N_23826);
nand UO_751 (O_751,N_19938,N_21455);
nand UO_752 (O_752,N_23073,N_22113);
or UO_753 (O_753,N_24649,N_19289);
nor UO_754 (O_754,N_20340,N_22161);
and UO_755 (O_755,N_20888,N_24800);
nor UO_756 (O_756,N_18976,N_19804);
or UO_757 (O_757,N_19105,N_19586);
nand UO_758 (O_758,N_24027,N_23707);
and UO_759 (O_759,N_20114,N_22287);
and UO_760 (O_760,N_22721,N_18802);
and UO_761 (O_761,N_21050,N_19389);
nor UO_762 (O_762,N_19532,N_22054);
xnor UO_763 (O_763,N_18900,N_22975);
xnor UO_764 (O_764,N_24406,N_20751);
or UO_765 (O_765,N_19347,N_21966);
nor UO_766 (O_766,N_22211,N_20612);
and UO_767 (O_767,N_21845,N_19839);
and UO_768 (O_768,N_22416,N_22048);
xor UO_769 (O_769,N_22964,N_24696);
nand UO_770 (O_770,N_24898,N_23291);
and UO_771 (O_771,N_18855,N_22559);
or UO_772 (O_772,N_24962,N_20001);
nor UO_773 (O_773,N_23492,N_21562);
nand UO_774 (O_774,N_22038,N_19770);
nand UO_775 (O_775,N_21122,N_23176);
nand UO_776 (O_776,N_18980,N_23645);
nand UO_777 (O_777,N_20609,N_20584);
xor UO_778 (O_778,N_20782,N_22484);
or UO_779 (O_779,N_20320,N_20950);
and UO_780 (O_780,N_19119,N_23427);
xnor UO_781 (O_781,N_20335,N_23274);
and UO_782 (O_782,N_24855,N_22396);
xnor UO_783 (O_783,N_23658,N_21624);
and UO_784 (O_784,N_23614,N_24752);
or UO_785 (O_785,N_23916,N_23520);
or UO_786 (O_786,N_24299,N_23887);
nor UO_787 (O_787,N_20706,N_23788);
nor UO_788 (O_788,N_23951,N_22832);
xnor UO_789 (O_789,N_21468,N_22889);
nand UO_790 (O_790,N_22230,N_23741);
nor UO_791 (O_791,N_19832,N_20999);
and UO_792 (O_792,N_23222,N_19497);
and UO_793 (O_793,N_20618,N_21403);
or UO_794 (O_794,N_23535,N_22712);
nand UO_795 (O_795,N_19686,N_18820);
nor UO_796 (O_796,N_19946,N_24578);
xnor UO_797 (O_797,N_22126,N_22645);
nor UO_798 (O_798,N_21030,N_20313);
and UO_799 (O_799,N_24765,N_23436);
nor UO_800 (O_800,N_24281,N_24882);
nand UO_801 (O_801,N_21121,N_22393);
nor UO_802 (O_802,N_19452,N_24859);
and UO_803 (O_803,N_19050,N_20148);
nor UO_804 (O_804,N_24788,N_21693);
or UO_805 (O_805,N_18960,N_19745);
or UO_806 (O_806,N_20577,N_24134);
or UO_807 (O_807,N_24978,N_21367);
nor UO_808 (O_808,N_20139,N_22443);
nand UO_809 (O_809,N_20610,N_23135);
nand UO_810 (O_810,N_22994,N_23359);
nand UO_811 (O_811,N_23217,N_20641);
or UO_812 (O_812,N_22756,N_20327);
xnor UO_813 (O_813,N_23250,N_20975);
or UO_814 (O_814,N_24682,N_22489);
or UO_815 (O_815,N_21025,N_22710);
and UO_816 (O_816,N_20659,N_22325);
and UO_817 (O_817,N_23225,N_23345);
and UO_818 (O_818,N_21995,N_21801);
nor UO_819 (O_819,N_23893,N_19077);
nand UO_820 (O_820,N_22459,N_19341);
nor UO_821 (O_821,N_19433,N_24031);
or UO_822 (O_822,N_23267,N_23987);
and UO_823 (O_823,N_19874,N_22622);
nand UO_824 (O_824,N_19369,N_24926);
and UO_825 (O_825,N_24829,N_22529);
nor UO_826 (O_826,N_22943,N_21749);
nor UO_827 (O_827,N_18950,N_19233);
and UO_828 (O_828,N_21650,N_23700);
and UO_829 (O_829,N_24373,N_23346);
or UO_830 (O_830,N_21167,N_20121);
nand UO_831 (O_831,N_22961,N_18967);
nor UO_832 (O_832,N_19894,N_20553);
and UO_833 (O_833,N_21564,N_21396);
or UO_834 (O_834,N_20501,N_19298);
or UO_835 (O_835,N_19103,N_21716);
nand UO_836 (O_836,N_19140,N_23373);
nand UO_837 (O_837,N_24471,N_22672);
and UO_838 (O_838,N_22349,N_20844);
and UO_839 (O_839,N_23158,N_18787);
or UO_840 (O_840,N_23683,N_21603);
nor UO_841 (O_841,N_19633,N_19751);
nand UO_842 (O_842,N_18758,N_24171);
nor UO_843 (O_843,N_23091,N_22574);
or UO_844 (O_844,N_24184,N_19263);
xnor UO_845 (O_845,N_22467,N_24714);
and UO_846 (O_846,N_23367,N_19840);
and UO_847 (O_847,N_24492,N_18886);
and UO_848 (O_848,N_23529,N_21924);
and UO_849 (O_849,N_22163,N_24836);
nand UO_850 (O_850,N_19013,N_20901);
and UO_851 (O_851,N_23061,N_24300);
and UO_852 (O_852,N_22682,N_24671);
or UO_853 (O_853,N_22785,N_21907);
nand UO_854 (O_854,N_20328,N_21126);
nand UO_855 (O_855,N_19108,N_20482);
xor UO_856 (O_856,N_19769,N_20905);
nand UO_857 (O_857,N_24860,N_19976);
nand UO_858 (O_858,N_22018,N_19004);
nand UO_859 (O_859,N_21988,N_20029);
nor UO_860 (O_860,N_19821,N_22341);
or UO_861 (O_861,N_24282,N_19766);
nand UO_862 (O_862,N_22452,N_24206);
and UO_863 (O_863,N_22531,N_23287);
and UO_864 (O_864,N_21842,N_23540);
nand UO_865 (O_865,N_23019,N_21936);
or UO_866 (O_866,N_22794,N_19718);
and UO_867 (O_867,N_21983,N_18970);
or UO_868 (O_868,N_23076,N_20613);
or UO_869 (O_869,N_24221,N_23048);
xnor UO_870 (O_870,N_20360,N_23431);
nor UO_871 (O_871,N_21280,N_20693);
or UO_872 (O_872,N_19713,N_21714);
or UO_873 (O_873,N_22278,N_21751);
or UO_874 (O_874,N_23042,N_19672);
or UO_875 (O_875,N_20347,N_20964);
or UO_876 (O_876,N_21584,N_20476);
or UO_877 (O_877,N_19543,N_22090);
and UO_878 (O_878,N_21438,N_19240);
and UO_879 (O_879,N_21102,N_21430);
or UO_880 (O_880,N_23803,N_23888);
xor UO_881 (O_881,N_24773,N_19525);
nor UO_882 (O_882,N_21039,N_22900);
nand UO_883 (O_883,N_21882,N_24006);
nand UO_884 (O_884,N_24628,N_23146);
xor UO_885 (O_885,N_20199,N_21273);
nor UO_886 (O_886,N_22199,N_22179);
and UO_887 (O_887,N_20834,N_23835);
or UO_888 (O_888,N_19781,N_21998);
nor UO_889 (O_889,N_21946,N_21707);
or UO_890 (O_890,N_22649,N_21556);
nor UO_891 (O_891,N_21823,N_20614);
and UO_892 (O_892,N_21503,N_24409);
and UO_893 (O_893,N_19411,N_19145);
or UO_894 (O_894,N_19936,N_18868);
and UO_895 (O_895,N_23376,N_24721);
and UO_896 (O_896,N_23676,N_19191);
and UO_897 (O_897,N_20122,N_18854);
and UO_898 (O_898,N_19167,N_19688);
nand UO_899 (O_899,N_20664,N_22714);
and UO_900 (O_900,N_19373,N_18930);
and UO_901 (O_901,N_22949,N_24571);
xnor UO_902 (O_902,N_19867,N_19358);
xor UO_903 (O_903,N_21209,N_19961);
or UO_904 (O_904,N_24337,N_21344);
or UO_905 (O_905,N_20703,N_21646);
or UO_906 (O_906,N_19280,N_23962);
nand UO_907 (O_907,N_20349,N_20972);
nand UO_908 (O_908,N_24893,N_22540);
nand UO_909 (O_909,N_24227,N_21110);
or UO_910 (O_910,N_21301,N_24885);
nand UO_911 (O_911,N_24942,N_23339);
and UO_912 (O_912,N_19375,N_20058);
and UO_913 (O_913,N_22959,N_20848);
or UO_914 (O_914,N_21303,N_19084);
and UO_915 (O_915,N_24560,N_20292);
nand UO_916 (O_916,N_22114,N_24161);
nor UO_917 (O_917,N_22706,N_21788);
xnor UO_918 (O_918,N_20494,N_23447);
nor UO_919 (O_919,N_19086,N_19756);
and UO_920 (O_920,N_22539,N_21967);
nor UO_921 (O_921,N_20100,N_19792);
and UO_922 (O_922,N_23850,N_20000);
or UO_923 (O_923,N_21449,N_20245);
and UO_924 (O_924,N_19134,N_23537);
nand UO_925 (O_925,N_19697,N_18890);
and UO_926 (O_926,N_19205,N_21753);
and UO_927 (O_927,N_24494,N_20416);
or UO_928 (O_928,N_24013,N_19198);
nor UO_929 (O_929,N_20600,N_23210);
or UO_930 (O_930,N_20762,N_20549);
and UO_931 (O_931,N_22566,N_23513);
and UO_932 (O_932,N_24257,N_21690);
xor UO_933 (O_933,N_23958,N_23470);
nor UO_934 (O_934,N_23919,N_21981);
or UO_935 (O_935,N_21215,N_24611);
and UO_936 (O_936,N_22898,N_20129);
xor UO_937 (O_937,N_20259,N_18867);
or UO_938 (O_938,N_20464,N_24813);
and UO_939 (O_939,N_24450,N_21910);
nor UO_940 (O_940,N_24535,N_19842);
or UO_941 (O_941,N_23539,N_24359);
nor UO_942 (O_942,N_24889,N_20297);
and UO_943 (O_943,N_20809,N_22821);
or UO_944 (O_944,N_22079,N_22658);
nand UO_945 (O_945,N_24580,N_22332);
nand UO_946 (O_946,N_24976,N_21563);
nor UO_947 (O_947,N_19514,N_23416);
nand UO_948 (O_948,N_23978,N_23112);
nor UO_949 (O_949,N_20102,N_22874);
nor UO_950 (O_950,N_21571,N_24093);
nand UO_951 (O_951,N_21448,N_24911);
nor UO_952 (O_952,N_23797,N_22181);
or UO_953 (O_953,N_24920,N_23972);
nand UO_954 (O_954,N_22448,N_19264);
nor UO_955 (O_955,N_23621,N_24657);
or UO_956 (O_956,N_24551,N_21846);
nor UO_957 (O_957,N_23240,N_19998);
nor UO_958 (O_958,N_21546,N_21472);
nand UO_959 (O_959,N_22727,N_24599);
nand UO_960 (O_960,N_22254,N_23940);
nand UO_961 (O_961,N_20597,N_22801);
and UO_962 (O_962,N_19097,N_23902);
or UO_963 (O_963,N_24316,N_23541);
nor UO_964 (O_964,N_20928,N_21594);
and UO_965 (O_965,N_24692,N_22219);
nand UO_966 (O_966,N_19075,N_23342);
nor UO_967 (O_967,N_24256,N_22248);
nand UO_968 (O_968,N_24078,N_23066);
and UO_969 (O_969,N_19635,N_20984);
nor UO_970 (O_970,N_18751,N_24770);
nor UO_971 (O_971,N_20215,N_23361);
and UO_972 (O_972,N_23371,N_20918);
and UO_973 (O_973,N_24198,N_20378);
nand UO_974 (O_974,N_23684,N_21341);
xor UO_975 (O_975,N_21444,N_21802);
and UO_976 (O_976,N_23554,N_20048);
nor UO_977 (O_977,N_22852,N_21071);
nand UO_978 (O_978,N_24251,N_24075);
or UO_979 (O_979,N_21460,N_19995);
nand UO_980 (O_980,N_24532,N_23273);
and UO_981 (O_981,N_21657,N_23750);
or UO_982 (O_982,N_23605,N_24151);
or UO_983 (O_983,N_24479,N_20933);
nor UO_984 (O_984,N_20729,N_19451);
or UO_985 (O_985,N_23336,N_20172);
xor UO_986 (O_986,N_24772,N_19575);
nor UO_987 (O_987,N_18969,N_19045);
and UO_988 (O_988,N_24834,N_22702);
nand UO_989 (O_989,N_20221,N_23863);
and UO_990 (O_990,N_20237,N_22195);
nor UO_991 (O_991,N_23494,N_21465);
or UO_992 (O_992,N_20329,N_23058);
nor UO_993 (O_993,N_19294,N_24516);
nor UO_994 (O_994,N_21840,N_23599);
nor UO_995 (O_995,N_23846,N_22629);
xnor UO_996 (O_996,N_23698,N_24957);
or UO_997 (O_997,N_24745,N_24792);
or UO_998 (O_998,N_19249,N_22472);
nor UO_999 (O_999,N_23949,N_24135);
nor UO_1000 (O_1000,N_18988,N_22942);
and UO_1001 (O_1001,N_22421,N_21761);
and UO_1002 (O_1002,N_23624,N_23264);
nand UO_1003 (O_1003,N_22652,N_19761);
or UO_1004 (O_1004,N_24822,N_23095);
nor UO_1005 (O_1005,N_20851,N_24250);
and UO_1006 (O_1006,N_24994,N_23364);
nor UO_1007 (O_1007,N_23186,N_23749);
nor UO_1008 (O_1008,N_24378,N_24603);
xnor UO_1009 (O_1009,N_23576,N_20467);
nand UO_1010 (O_1010,N_22781,N_19639);
or UO_1011 (O_1011,N_24779,N_21105);
nand UO_1012 (O_1012,N_20420,N_18815);
nand UO_1013 (O_1013,N_21841,N_24679);
nor UO_1014 (O_1014,N_24807,N_20361);
and UO_1015 (O_1015,N_23884,N_21961);
and UO_1016 (O_1016,N_21906,N_19217);
xor UO_1017 (O_1017,N_21704,N_20671);
nand UO_1018 (O_1018,N_19663,N_20257);
and UO_1019 (O_1019,N_21432,N_23184);
nor UO_1020 (O_1020,N_24413,N_23488);
and UO_1021 (O_1021,N_19727,N_24927);
nor UO_1022 (O_1022,N_22554,N_18777);
and UO_1023 (O_1023,N_22695,N_21653);
xnor UO_1024 (O_1024,N_18799,N_21941);
and UO_1025 (O_1025,N_20793,N_21922);
or UO_1026 (O_1026,N_23102,N_22690);
nand UO_1027 (O_1027,N_20603,N_23693);
or UO_1028 (O_1028,N_20119,N_19036);
nor UO_1029 (O_1029,N_19814,N_20858);
nand UO_1030 (O_1030,N_20249,N_24520);
nand UO_1031 (O_1031,N_24708,N_19436);
nand UO_1032 (O_1032,N_22967,N_23295);
nand UO_1033 (O_1033,N_20836,N_22049);
or UO_1034 (O_1034,N_18831,N_24537);
xor UO_1035 (O_1035,N_24989,N_20023);
xor UO_1036 (O_1036,N_22420,N_19102);
nor UO_1037 (O_1037,N_20463,N_19550);
and UO_1038 (O_1038,N_19372,N_20282);
nand UO_1039 (O_1039,N_23760,N_23729);
xor UO_1040 (O_1040,N_22750,N_21070);
nor UO_1041 (O_1041,N_20054,N_20737);
nand UO_1042 (O_1042,N_24811,N_20862);
or UO_1043 (O_1043,N_22112,N_20760);
nand UO_1044 (O_1044,N_21466,N_19378);
and UO_1045 (O_1045,N_19423,N_22450);
or UO_1046 (O_1046,N_24574,N_19308);
nor UO_1047 (O_1047,N_22470,N_19120);
or UO_1048 (O_1048,N_23792,N_20546);
or UO_1049 (O_1049,N_24020,N_20806);
nand UO_1050 (O_1050,N_22013,N_21576);
nor UO_1051 (O_1051,N_24043,N_20872);
or UO_1052 (O_1052,N_23084,N_19201);
or UO_1053 (O_1053,N_21703,N_21855);
or UO_1054 (O_1054,N_21909,N_24703);
nand UO_1055 (O_1055,N_18952,N_21445);
nand UO_1056 (O_1056,N_21602,N_20030);
or UO_1057 (O_1057,N_20935,N_19459);
nand UO_1058 (O_1058,N_20078,N_24040);
and UO_1059 (O_1059,N_21145,N_24382);
nand UO_1060 (O_1060,N_22436,N_19227);
nand UO_1061 (O_1061,N_21568,N_18883);
and UO_1062 (O_1062,N_21520,N_20075);
and UO_1063 (O_1063,N_22412,N_22073);
nor UO_1064 (O_1064,N_20387,N_22410);
or UO_1065 (O_1065,N_20371,N_22610);
or UO_1066 (O_1066,N_23839,N_22583);
nand UO_1067 (O_1067,N_19462,N_24433);
or UO_1068 (O_1068,N_21082,N_21144);
nand UO_1069 (O_1069,N_20593,N_24640);
or UO_1070 (O_1070,N_24643,N_24352);
and UO_1071 (O_1071,N_24029,N_21136);
xor UO_1072 (O_1072,N_24645,N_21876);
and UO_1073 (O_1073,N_18989,N_20436);
nor UO_1074 (O_1074,N_23830,N_20535);
nor UO_1075 (O_1075,N_24766,N_21724);
nor UO_1076 (O_1076,N_22076,N_23872);
xnor UO_1077 (O_1077,N_23415,N_20368);
xor UO_1078 (O_1078,N_22950,N_20189);
and UO_1079 (O_1079,N_22173,N_20388);
and UO_1080 (O_1080,N_21621,N_19509);
and UO_1081 (O_1081,N_23646,N_19340);
and UO_1082 (O_1082,N_22655,N_22444);
nor UO_1083 (O_1083,N_21377,N_22921);
or UO_1084 (O_1084,N_20492,N_20908);
xnor UO_1085 (O_1085,N_23246,N_23739);
nand UO_1086 (O_1086,N_22617,N_19073);
or UO_1087 (O_1087,N_20020,N_24469);
and UO_1088 (O_1088,N_19408,N_24484);
nand UO_1089 (O_1089,N_24534,N_24817);
nor UO_1090 (O_1090,N_24818,N_23285);
and UO_1091 (O_1091,N_19056,N_24781);
nand UO_1092 (O_1092,N_20695,N_19185);
nand UO_1093 (O_1093,N_21275,N_19071);
xor UO_1094 (O_1094,N_21130,N_21295);
or UO_1095 (O_1095,N_19314,N_22184);
xnor UO_1096 (O_1096,N_22726,N_21463);
xor UO_1097 (O_1097,N_20392,N_20496);
or UO_1098 (O_1098,N_20076,N_23213);
and UO_1099 (O_1099,N_21997,N_21669);
or UO_1100 (O_1100,N_20690,N_19802);
or UO_1101 (O_1101,N_22296,N_22468);
and UO_1102 (O_1102,N_21645,N_19777);
nand UO_1103 (O_1103,N_22953,N_19029);
nor UO_1104 (O_1104,N_21177,N_21994);
nand UO_1105 (O_1105,N_23384,N_19645);
nor UO_1106 (O_1106,N_23564,N_19815);
nor UO_1107 (O_1107,N_19789,N_23347);
nor UO_1108 (O_1108,N_21515,N_22357);
xor UO_1109 (O_1109,N_18956,N_20118);
nor UO_1110 (O_1110,N_24756,N_21986);
nand UO_1111 (O_1111,N_22514,N_21210);
and UO_1112 (O_1112,N_21480,N_21038);
nor UO_1113 (O_1113,N_20606,N_19636);
and UO_1114 (O_1114,N_23228,N_21253);
or UO_1115 (O_1115,N_23550,N_19632);
nand UO_1116 (O_1116,N_21383,N_19613);
nand UO_1117 (O_1117,N_19728,N_22958);
xnor UO_1118 (O_1118,N_23122,N_22810);
and UO_1119 (O_1119,N_22837,N_23755);
or UO_1120 (O_1120,N_19629,N_18864);
and UO_1121 (O_1121,N_21291,N_23282);
nor UO_1122 (O_1122,N_18972,N_19450);
nor UO_1123 (O_1123,N_20661,N_23206);
or UO_1124 (O_1124,N_18941,N_21847);
xor UO_1125 (O_1125,N_21813,N_22611);
nor UO_1126 (O_1126,N_19952,N_23138);
nand UO_1127 (O_1127,N_20251,N_19715);
or UO_1128 (O_1128,N_24320,N_23836);
xor UO_1129 (O_1129,N_20205,N_20545);
and UO_1130 (O_1130,N_23603,N_21277);
nor UO_1131 (O_1131,N_23142,N_23078);
nand UO_1132 (O_1132,N_20538,N_24375);
nor UO_1133 (O_1133,N_22623,N_22011);
nand UO_1134 (O_1134,N_24287,N_22650);
nor UO_1135 (O_1135,N_23772,N_19631);
nand UO_1136 (O_1136,N_20650,N_22681);
nand UO_1137 (O_1137,N_24687,N_23973);
and UO_1138 (O_1138,N_19481,N_21349);
or UO_1139 (O_1139,N_20540,N_24934);
nand UO_1140 (O_1140,N_21225,N_23833);
nor UO_1141 (O_1141,N_22598,N_23397);
nor UO_1142 (O_1142,N_24462,N_22189);
nor UO_1143 (O_1143,N_22842,N_23023);
xor UO_1144 (O_1144,N_19228,N_24243);
and UO_1145 (O_1145,N_24396,N_19566);
nand UO_1146 (O_1146,N_19181,N_21723);
or UO_1147 (O_1147,N_24115,N_20101);
nand UO_1148 (O_1148,N_20256,N_24673);
nor UO_1149 (O_1149,N_22040,N_23686);
nand UO_1150 (O_1150,N_23716,N_20769);
and UO_1151 (O_1151,N_23097,N_23183);
nor UO_1152 (O_1152,N_18996,N_24096);
and UO_1153 (O_1153,N_21056,N_21425);
nor UO_1154 (O_1154,N_23975,N_23050);
or UO_1155 (O_1155,N_19901,N_19440);
nand UO_1156 (O_1156,N_19333,N_24207);
or UO_1157 (O_1157,N_22225,N_19858);
nor UO_1158 (O_1158,N_19132,N_19638);
nand UO_1159 (O_1159,N_24236,N_22397);
and UO_1160 (O_1160,N_20180,N_21524);
nor UO_1161 (O_1161,N_21810,N_19640);
nand UO_1162 (O_1162,N_22111,N_22257);
xor UO_1163 (O_1163,N_23680,N_24945);
nand UO_1164 (O_1164,N_23981,N_20502);
nand UO_1165 (O_1165,N_22509,N_22582);
and UO_1166 (O_1166,N_21077,N_21944);
xnor UO_1167 (O_1167,N_21817,N_19919);
xor UO_1168 (O_1168,N_21411,N_24987);
nor UO_1169 (O_1169,N_24487,N_23085);
nor UO_1170 (O_1170,N_24192,N_19602);
and UO_1171 (O_1171,N_22439,N_23417);
nor UO_1172 (O_1172,N_24483,N_20469);
or UO_1173 (O_1173,N_21266,N_23525);
nand UO_1174 (O_1174,N_20289,N_20899);
and UO_1175 (O_1175,N_23747,N_21203);
nand UO_1176 (O_1176,N_24827,N_24875);
nand UO_1177 (O_1177,N_24389,N_21337);
and UO_1178 (O_1178,N_21912,N_20229);
nor UO_1179 (O_1179,N_19401,N_22739);
nand UO_1180 (O_1180,N_22194,N_24044);
nand UO_1181 (O_1181,N_19253,N_19526);
or UO_1182 (O_1182,N_21590,N_22091);
or UO_1183 (O_1183,N_24912,N_21461);
nor UO_1184 (O_1184,N_22204,N_23642);
nand UO_1185 (O_1185,N_21803,N_21338);
nor UO_1186 (O_1186,N_23638,N_20089);
nand UO_1187 (O_1187,N_24228,N_21187);
nor UO_1188 (O_1188,N_20678,N_18848);
and UO_1189 (O_1189,N_23047,N_24594);
or UO_1190 (O_1190,N_21497,N_23620);
and UO_1191 (O_1191,N_20108,N_21006);
or UO_1192 (O_1192,N_24085,N_20453);
and UO_1193 (O_1193,N_19278,N_18953);
and UO_1194 (O_1194,N_22358,N_23214);
nand UO_1195 (O_1195,N_22854,N_19041);
and UO_1196 (O_1196,N_19288,N_24485);
and UO_1197 (O_1197,N_23532,N_19835);
nand UO_1198 (O_1198,N_19070,N_19357);
nor UO_1199 (O_1199,N_20017,N_23352);
or UO_1200 (O_1200,N_18789,N_24114);
nor UO_1201 (O_1201,N_21290,N_20817);
or UO_1202 (O_1202,N_24575,N_20623);
or UO_1203 (O_1203,N_22545,N_21160);
nor UO_1204 (O_1204,N_21323,N_22139);
nor UO_1205 (O_1205,N_22217,N_22999);
or UO_1206 (O_1206,N_19503,N_20311);
nor UO_1207 (O_1207,N_23874,N_23674);
nand UO_1208 (O_1208,N_22787,N_21574);
nor UO_1209 (O_1209,N_22106,N_22820);
or UO_1210 (O_1210,N_19404,N_23221);
nor UO_1211 (O_1211,N_20957,N_24497);
nor UO_1212 (O_1212,N_18819,N_21279);
nor UO_1213 (O_1213,N_19891,N_22441);
or UO_1214 (O_1214,N_23947,N_21980);
and UO_1215 (O_1215,N_20821,N_18909);
or UO_1216 (O_1216,N_20393,N_20886);
nor UO_1217 (O_1217,N_22304,N_18835);
xor UO_1218 (O_1218,N_22723,N_24905);
nand UO_1219 (O_1219,N_24768,N_22783);
xnor UO_1220 (O_1220,N_21319,N_21240);
and UO_1221 (O_1221,N_24886,N_19226);
or UO_1222 (O_1222,N_20810,N_20321);
or UO_1223 (O_1223,N_20601,N_23321);
nand UO_1224 (O_1224,N_21894,N_20405);
xnor UO_1225 (O_1225,N_22641,N_22427);
or UO_1226 (O_1226,N_21895,N_22766);
or UO_1227 (O_1227,N_24345,N_20713);
nand UO_1228 (O_1228,N_21640,N_21618);
and UO_1229 (O_1229,N_24732,N_18781);
nor UO_1230 (O_1230,N_20499,N_24426);
or UO_1231 (O_1231,N_21496,N_24035);
and UO_1232 (O_1232,N_24165,N_24009);
nand UO_1233 (O_1233,N_22429,N_21581);
and UO_1234 (O_1234,N_21346,N_24819);
and UO_1235 (O_1235,N_19693,N_22925);
nand UO_1236 (O_1236,N_19608,N_22919);
and UO_1237 (O_1237,N_22576,N_23103);
nand UO_1238 (O_1238,N_20019,N_22913);
nor UO_1239 (O_1239,N_20522,N_22408);
nand UO_1240 (O_1240,N_20138,N_22651);
nand UO_1241 (O_1241,N_24943,N_23014);
or UO_1242 (O_1242,N_23402,N_21233);
or UO_1243 (O_1243,N_19848,N_23350);
or UO_1244 (O_1244,N_20771,N_19156);
nor UO_1245 (O_1245,N_23607,N_19665);
or UO_1246 (O_1246,N_19523,N_24451);
or UO_1247 (O_1247,N_19161,N_20565);
and UO_1248 (O_1248,N_24154,N_24339);
nor UO_1249 (O_1249,N_20381,N_22550);
and UO_1250 (O_1250,N_24466,N_24079);
xor UO_1251 (O_1251,N_23409,N_21237);
and UO_1252 (O_1252,N_22834,N_20940);
and UO_1253 (O_1253,N_20870,N_22527);
or UO_1254 (O_1254,N_24980,N_19896);
and UO_1255 (O_1255,N_24646,N_22644);
nand UO_1256 (O_1256,N_24953,N_22036);
or UO_1257 (O_1257,N_22984,N_24731);
and UO_1258 (O_1258,N_23486,N_23506);
nand UO_1259 (O_1259,N_21326,N_23865);
nor UO_1260 (O_1260,N_22873,N_19960);
nand UO_1261 (O_1261,N_19763,N_24422);
xor UO_1262 (O_1262,N_19983,N_24619);
xnor UO_1263 (O_1263,N_23794,N_23932);
or UO_1264 (O_1264,N_23615,N_20190);
nand UO_1265 (O_1265,N_24289,N_21558);
or UO_1266 (O_1266,N_24055,N_20355);
and UO_1267 (O_1267,N_22074,N_22380);
xnor UO_1268 (O_1268,N_23432,N_20345);
nand UO_1269 (O_1269,N_22520,N_23965);
or UO_1270 (O_1270,N_21388,N_21746);
nand UO_1271 (O_1271,N_20224,N_21402);
and UO_1272 (O_1272,N_24437,N_20781);
nor UO_1273 (O_1273,N_19026,N_20630);
nand UO_1274 (O_1274,N_20419,N_18770);
xnor UO_1275 (O_1275,N_20319,N_20787);
or UO_1276 (O_1276,N_19040,N_20439);
nand UO_1277 (O_1277,N_24883,N_21081);
and UO_1278 (O_1278,N_21436,N_23163);
nor UO_1279 (O_1279,N_20738,N_24705);
nand UO_1280 (O_1280,N_20165,N_18786);
nand UO_1281 (O_1281,N_21778,N_22425);
nand UO_1282 (O_1282,N_18857,N_21278);
nor UO_1283 (O_1283,N_24474,N_18882);
nor UO_1284 (O_1284,N_22747,N_21930);
nor UO_1285 (O_1285,N_22228,N_24794);
or UO_1286 (O_1286,N_22648,N_21863);
and UO_1287 (O_1287,N_21923,N_24515);
and UO_1288 (O_1288,N_22023,N_24218);
or UO_1289 (O_1289,N_23262,N_20208);
or UO_1290 (O_1290,N_20111,N_23358);
and UO_1291 (O_1291,N_20488,N_24614);
nor UO_1292 (O_1292,N_22528,N_20302);
xnor UO_1293 (O_1293,N_19568,N_19311);
xor UO_1294 (O_1294,N_20203,N_24341);
nor UO_1295 (O_1295,N_24276,N_21076);
or UO_1296 (O_1296,N_18977,N_20758);
xnor UO_1297 (O_1297,N_21685,N_23059);
and UO_1298 (O_1298,N_23968,N_23120);
or UO_1299 (O_1299,N_24521,N_24854);
nor UO_1300 (O_1300,N_21153,N_23153);
xnor UO_1301 (O_1301,N_21570,N_19630);
xor UO_1302 (O_1302,N_22302,N_18866);
or UO_1303 (O_1303,N_24057,N_23038);
and UO_1304 (O_1304,N_20198,N_24763);
nand UO_1305 (O_1305,N_23630,N_20326);
nand UO_1306 (O_1306,N_20556,N_23542);
nor UO_1307 (O_1307,N_22500,N_24801);
or UO_1308 (O_1308,N_18913,N_19355);
or UO_1309 (O_1309,N_19912,N_24175);
nand UO_1310 (O_1310,N_21061,N_23841);
and UO_1311 (O_1311,N_20842,N_24977);
xnor UO_1312 (O_1312,N_24331,N_23834);
or UO_1313 (O_1313,N_22526,N_21706);
and UO_1314 (O_1314,N_20383,N_23666);
nor UO_1315 (O_1315,N_21942,N_23960);
and UO_1316 (O_1316,N_19005,N_19223);
xor UO_1317 (O_1317,N_24348,N_22506);
and UO_1318 (O_1318,N_22169,N_22972);
nand UO_1319 (O_1319,N_22383,N_22877);
and UO_1320 (O_1320,N_20166,N_20856);
nand UO_1321 (O_1321,N_19619,N_22515);
nand UO_1322 (O_1322,N_20646,N_22763);
nand UO_1323 (O_1323,N_22125,N_20801);
and UO_1324 (O_1324,N_23446,N_18940);
or UO_1325 (O_1325,N_20633,N_19897);
nand UO_1326 (O_1326,N_24125,N_24354);
and UO_1327 (O_1327,N_21962,N_23829);
nand UO_1328 (O_1328,N_21879,N_23175);
nor UO_1329 (O_1329,N_23174,N_23569);
nor UO_1330 (O_1330,N_20373,N_23655);
and UO_1331 (O_1331,N_22738,N_23170);
and UO_1332 (O_1332,N_24897,N_19064);
nand UO_1333 (O_1333,N_21046,N_20395);
nor UO_1334 (O_1334,N_21181,N_19687);
nor UO_1335 (O_1335,N_22019,N_21881);
nor UO_1336 (O_1336,N_21975,N_22382);
or UO_1337 (O_1337,N_20449,N_23860);
and UO_1338 (O_1338,N_20937,N_23293);
nand UO_1339 (O_1339,N_19022,N_21620);
and UO_1340 (O_1340,N_19024,N_22654);
nand UO_1341 (O_1341,N_19114,N_21127);
nor UO_1342 (O_1342,N_21074,N_24053);
or UO_1343 (O_1343,N_19856,N_22729);
nor UO_1344 (O_1344,N_24840,N_23854);
nor UO_1345 (O_1345,N_22039,N_23338);
or UO_1346 (O_1346,N_22498,N_21908);
nand UO_1347 (O_1347,N_24229,N_19498);
nor UO_1348 (O_1348,N_19705,N_22584);
and UO_1349 (O_1349,N_22451,N_20512);
and UO_1350 (O_1350,N_19513,N_18828);
nand UO_1351 (O_1351,N_21779,N_19083);
or UO_1352 (O_1352,N_18860,N_22691);
and UO_1353 (O_1353,N_20210,N_20110);
or UO_1354 (O_1354,N_20084,N_22944);
nand UO_1355 (O_1355,N_21433,N_21610);
nand UO_1356 (O_1356,N_23150,N_24658);
and UO_1357 (O_1357,N_20750,N_21022);
nand UO_1358 (O_1358,N_20652,N_18812);
and UO_1359 (O_1359,N_24999,N_24431);
and UO_1360 (O_1360,N_24324,N_20792);
nor UO_1361 (O_1361,N_24186,N_24874);
or UO_1362 (O_1362,N_20468,N_21334);
or UO_1363 (O_1363,N_20470,N_21512);
nand UO_1364 (O_1364,N_23982,N_22589);
xor UO_1365 (O_1365,N_22394,N_24554);
and UO_1366 (O_1366,N_24472,N_20900);
nor UO_1367 (O_1367,N_23610,N_20668);
nor UO_1368 (O_1368,N_24160,N_21957);
nand UO_1369 (O_1369,N_21108,N_20669);
nand UO_1370 (O_1370,N_23189,N_23723);
or UO_1371 (O_1371,N_23044,N_20334);
nor UO_1372 (O_1372,N_20881,N_24202);
nand UO_1373 (O_1373,N_22143,N_23099);
nor UO_1374 (O_1374,N_24330,N_19898);
and UO_1375 (O_1375,N_21394,N_24408);
or UO_1376 (O_1376,N_20428,N_24199);
and UO_1377 (O_1377,N_20980,N_18754);
nor UO_1378 (O_1378,N_23980,N_20261);
and UO_1379 (O_1379,N_23732,N_23319);
nor UO_1380 (O_1380,N_23804,N_23303);
and UO_1381 (O_1381,N_22814,N_24852);
nand UO_1382 (O_1382,N_21976,N_24688);
or UO_1383 (O_1383,N_24625,N_23021);
or UO_1384 (O_1384,N_23315,N_22288);
and UO_1385 (O_1385,N_22251,N_20926);
or UO_1386 (O_1386,N_24327,N_23448);
or UO_1387 (O_1387,N_21395,N_24191);
xnor UO_1388 (O_1388,N_23717,N_18794);
nand UO_1389 (O_1389,N_24947,N_22965);
nor UO_1390 (O_1390,N_22192,N_21947);
or UO_1391 (O_1391,N_24533,N_22907);
nor UO_1392 (O_1392,N_20767,N_23789);
nand UO_1393 (O_1393,N_23406,N_18937);
or UO_1394 (O_1394,N_22806,N_22728);
nor UO_1395 (O_1395,N_21679,N_24672);
xor UO_1396 (O_1396,N_20934,N_20351);
and UO_1397 (O_1397,N_23013,N_23873);
nand UO_1398 (O_1398,N_22631,N_22045);
xnor UO_1399 (O_1399,N_20608,N_23422);
xor UO_1400 (O_1400,N_20916,N_19857);
and UO_1401 (O_1401,N_20953,N_22108);
nor UO_1402 (O_1402,N_22008,N_20629);
nand UO_1403 (O_1403,N_19171,N_22668);
nor UO_1404 (O_1404,N_24593,N_21709);
xnor UO_1405 (O_1405,N_20871,N_22210);
and UO_1406 (O_1406,N_19445,N_22286);
nor UO_1407 (O_1407,N_22892,N_24946);
and UO_1408 (O_1408,N_19556,N_19096);
and UO_1409 (O_1409,N_20316,N_23606);
nor UO_1410 (O_1410,N_21166,N_24780);
and UO_1411 (O_1411,N_24367,N_23410);
xor UO_1412 (O_1412,N_24054,N_21530);
and UO_1413 (O_1413,N_19963,N_21080);
xor UO_1414 (O_1414,N_20412,N_24675);
nor UO_1415 (O_1415,N_24365,N_24019);
nand UO_1416 (O_1416,N_20239,N_23370);
or UO_1417 (O_1417,N_22708,N_23208);
and UO_1418 (O_1418,N_19795,N_18962);
nand UO_1419 (O_1419,N_24993,N_23281);
xnor UO_1420 (O_1420,N_23955,N_20402);
nand UO_1421 (O_1421,N_24729,N_21782);
or UO_1422 (O_1422,N_23037,N_19377);
or UO_1423 (O_1423,N_21667,N_21862);
nand UO_1424 (O_1424,N_20057,N_22960);
or UO_1425 (O_1425,N_19579,N_22297);
and UO_1426 (O_1426,N_24288,N_24787);
or UO_1427 (O_1427,N_22751,N_24608);
and UO_1428 (O_1428,N_19058,N_23064);
and UO_1429 (O_1429,N_21342,N_21697);
nor UO_1430 (O_1430,N_24531,N_21264);
or UO_1431 (O_1431,N_19326,N_23764);
nor UO_1432 (O_1432,N_19443,N_21034);
and UO_1433 (O_1433,N_23498,N_21168);
xnor UO_1434 (O_1434,N_23985,N_24265);
nor UO_1435 (O_1435,N_20698,N_20293);
nor UO_1436 (O_1436,N_23711,N_24232);
or UO_1437 (O_1437,N_23966,N_23546);
nor UO_1438 (O_1438,N_19701,N_23754);
or UO_1439 (O_1439,N_23320,N_20344);
nor UO_1440 (O_1440,N_23724,N_19299);
xor UO_1441 (O_1441,N_20967,N_24615);
or UO_1442 (O_1442,N_19435,N_22187);
and UO_1443 (O_1443,N_22671,N_19432);
or UO_1444 (O_1444,N_24581,N_21495);
nand UO_1445 (O_1445,N_20663,N_21212);
nor UO_1446 (O_1446,N_18910,N_19431);
nand UO_1447 (O_1447,N_24634,N_18869);
nor UO_1448 (O_1448,N_20672,N_21809);
nor UO_1449 (O_1449,N_23481,N_21312);
and UO_1450 (O_1450,N_23192,N_23380);
and UO_1451 (O_1451,N_22390,N_23223);
and UO_1452 (O_1452,N_20307,N_21286);
nand UO_1453 (O_1453,N_20869,N_22697);
or UO_1454 (O_1454,N_22078,N_21023);
or UO_1455 (O_1455,N_21420,N_22307);
nor UO_1456 (O_1456,N_23144,N_23697);
or UO_1457 (O_1457,N_19129,N_22002);
xnor UO_1458 (O_1458,N_19370,N_21938);
nor UO_1459 (O_1459,N_19884,N_24047);
nor UO_1460 (O_1460,N_23894,N_22371);
or UO_1461 (O_1461,N_19242,N_22995);
nand UO_1462 (O_1462,N_19009,N_24723);
or UO_1463 (O_1463,N_18762,N_20615);
or UO_1464 (O_1464,N_20032,N_23822);
and UO_1465 (O_1465,N_24444,N_21067);
nand UO_1466 (O_1466,N_19147,N_21005);
or UO_1467 (O_1467,N_19123,N_20805);
and UO_1468 (O_1468,N_20700,N_22414);
or UO_1469 (O_1469,N_22066,N_22005);
xor UO_1470 (O_1470,N_21117,N_21505);
nand UO_1471 (O_1471,N_23612,N_20080);
nand UO_1472 (O_1472,N_20162,N_22845);
nand UO_1473 (O_1473,N_19574,N_24260);
and UO_1474 (O_1474,N_21284,N_22293);
and UO_1475 (O_1475,N_19587,N_20200);
nand UO_1476 (O_1476,N_20133,N_24086);
nand UO_1477 (O_1477,N_19914,N_22085);
nor UO_1478 (O_1478,N_20098,N_20573);
nor UO_1479 (O_1479,N_22945,N_18912);
nor UO_1480 (O_1480,N_19444,N_23999);
nand UO_1481 (O_1481,N_19624,N_24022);
or UO_1482 (O_1482,N_20831,N_23815);
nor UO_1483 (O_1483,N_22176,N_23459);
and UO_1484 (O_1484,N_24895,N_20015);
and UO_1485 (O_1485,N_20035,N_22725);
nand UO_1486 (O_1486,N_19571,N_21717);
xor UO_1487 (O_1487,N_20893,N_22037);
nor UO_1488 (O_1488,N_19173,N_23665);
or UO_1489 (O_1489,N_24188,N_18921);
xor UO_1490 (O_1490,N_22455,N_22676);
nand UO_1491 (O_1491,N_24686,N_21728);
or UO_1492 (O_1492,N_23040,N_22647);
xor UO_1493 (O_1493,N_22030,N_24454);
or UO_1494 (O_1494,N_18756,N_23266);
or UO_1495 (O_1495,N_22320,N_24815);
nand UO_1496 (O_1496,N_22214,N_19573);
nor UO_1497 (O_1497,N_24865,N_24694);
and UO_1498 (O_1498,N_22151,N_22263);
and UO_1499 (O_1499,N_21598,N_20919);
and UO_1500 (O_1500,N_21539,N_24064);
nand UO_1501 (O_1501,N_24936,N_21493);
or UO_1502 (O_1502,N_20513,N_19219);
and UO_1503 (O_1503,N_19797,N_19732);
and UO_1504 (O_1504,N_24605,N_20411);
nor UO_1505 (O_1505,N_19548,N_19182);
or UO_1506 (O_1506,N_19553,N_23005);
and UO_1507 (O_1507,N_20244,N_23691);
nor UO_1508 (O_1508,N_20846,N_18772);
nand UO_1509 (O_1509,N_21380,N_23396);
and UO_1510 (O_1510,N_20588,N_23335);
xor UO_1511 (O_1511,N_19865,N_21795);
nand UO_1512 (O_1512,N_23898,N_21595);
nand UO_1513 (O_1513,N_24724,N_20574);
and UO_1514 (O_1514,N_23200,N_24741);
nand UO_1515 (O_1515,N_24117,N_24238);
nand UO_1516 (O_1516,N_24877,N_22505);
and UO_1517 (O_1517,N_19324,N_24403);
nand UO_1518 (O_1518,N_18778,N_18851);
or UO_1519 (O_1519,N_21642,N_21528);
and UO_1520 (O_1520,N_19709,N_22138);
nand UO_1521 (O_1521,N_20024,N_21807);
nor UO_1522 (O_1522,N_20575,N_21047);
nor UO_1523 (O_1523,N_22850,N_18763);
or UO_1524 (O_1524,N_18842,N_21677);
nor UO_1525 (O_1525,N_21541,N_19028);
and UO_1526 (O_1526,N_22920,N_22255);
nor UO_1527 (O_1527,N_22635,N_21409);
or UO_1528 (O_1528,N_23080,N_24524);
nand UO_1529 (O_1529,N_21686,N_23907);
nand UO_1530 (O_1530,N_24394,N_22885);
and UO_1531 (O_1531,N_22369,N_21865);
nor UO_1532 (O_1532,N_21347,N_23926);
nand UO_1533 (O_1533,N_20145,N_20070);
nor UO_1534 (O_1534,N_23390,N_21949);
nand UO_1535 (O_1535,N_21868,N_20707);
and UO_1536 (O_1536,N_19899,N_23976);
and UO_1537 (O_1537,N_22129,N_23659);
and UO_1538 (O_1538,N_23455,N_19245);
xnor UO_1539 (O_1539,N_19778,N_24405);
nand UO_1540 (O_1540,N_21729,N_23560);
or UO_1541 (O_1541,N_22938,N_23428);
or UO_1542 (O_1542,N_23480,N_23123);
nand UO_1543 (O_1543,N_24862,N_23587);
nand UO_1544 (O_1544,N_20789,N_19817);
nand UO_1545 (O_1545,N_22133,N_24294);
and UO_1546 (O_1546,N_18753,N_20500);
and UO_1547 (O_1547,N_19755,N_24042);
nor UO_1548 (O_1548,N_21790,N_18813);
nor UO_1549 (O_1549,N_20666,N_24880);
nand UO_1550 (O_1550,N_19007,N_21507);
or UO_1551 (O_1551,N_19529,N_19562);
or UO_1552 (O_1552,N_19706,N_21659);
nor UO_1553 (O_1553,N_20681,N_22438);
and UO_1554 (O_1554,N_24782,N_22772);
nor UO_1555 (O_1555,N_21582,N_24323);
nor UO_1556 (O_1556,N_22833,N_24717);
and UO_1557 (O_1557,N_23404,N_22271);
nor UO_1558 (O_1558,N_21655,N_20421);
nor UO_1559 (O_1559,N_24503,N_22457);
nand UO_1560 (O_1560,N_23688,N_22931);
or UO_1561 (O_1561,N_23036,N_18832);
nor UO_1562 (O_1562,N_22086,N_18959);
or UO_1563 (O_1563,N_18825,N_21825);
or UO_1564 (O_1564,N_22817,N_23922);
nor UO_1565 (O_1565,N_22507,N_21903);
and UO_1566 (O_1566,N_24971,N_21681);
nand UO_1567 (O_1567,N_22258,N_24900);
nand UO_1568 (O_1568,N_23012,N_23728);
nor UO_1569 (O_1569,N_21000,N_19740);
nor UO_1570 (O_1570,N_22434,N_22923);
or UO_1571 (O_1571,N_24522,N_22848);
xor UO_1572 (O_1572,N_21171,N_19704);
xor UO_1573 (O_1573,N_22575,N_24495);
or UO_1574 (O_1574,N_22261,N_23140);
and UO_1575 (O_1575,N_23226,N_24376);
and UO_1576 (O_1576,N_21052,N_22530);
nand UO_1577 (O_1577,N_21743,N_21152);
or UO_1578 (O_1578,N_21453,N_20578);
nor UO_1579 (O_1579,N_23941,N_20087);
or UO_1580 (O_1580,N_24795,N_24328);
or UO_1581 (O_1581,N_22573,N_19658);
and UO_1582 (O_1582,N_20493,N_21960);
or UO_1583 (O_1583,N_20735,N_24104);
and UO_1584 (O_1584,N_22674,N_19142);
nor UO_1585 (O_1585,N_21300,N_19987);
nor UO_1586 (O_1586,N_22640,N_23034);
xnor UO_1587 (O_1587,N_21725,N_24850);
nor UO_1588 (O_1588,N_22680,N_22347);
nand UO_1589 (O_1589,N_24749,N_20976);
and UO_1590 (O_1590,N_24254,N_21740);
xnor UO_1591 (O_1591,N_22224,N_23864);
nand UO_1592 (O_1592,N_19472,N_19397);
xor UO_1593 (O_1593,N_24457,N_22673);
nor UO_1594 (O_1594,N_22555,N_23497);
nor UO_1595 (O_1595,N_23890,N_21609);
nor UO_1596 (O_1596,N_23994,N_21937);
and UO_1597 (O_1597,N_22423,N_19971);
and UO_1598 (O_1598,N_24972,N_24126);
nand UO_1599 (O_1599,N_22805,N_20860);
nor UO_1600 (O_1600,N_22849,N_22212);
nor UO_1601 (O_1601,N_22638,N_18994);
or UO_1602 (O_1602,N_20348,N_23593);
or UO_1603 (O_1603,N_22843,N_21486);
nor UO_1604 (O_1604,N_23702,N_21336);
nor UO_1605 (O_1605,N_22440,N_20692);
nor UO_1606 (O_1606,N_24653,N_24163);
or UO_1607 (O_1607,N_23136,N_21208);
and UO_1608 (O_1608,N_22903,N_21735);
xor UO_1609 (O_1609,N_23008,N_21851);
xor UO_1610 (O_1610,N_22572,N_24689);
or UO_1611 (O_1611,N_21891,N_24808);
xor UO_1612 (O_1612,N_22350,N_21674);
or UO_1613 (O_1613,N_24830,N_18806);
nor UO_1614 (O_1614,N_23194,N_24201);
or UO_1615 (O_1615,N_19409,N_23399);
and UO_1616 (O_1616,N_24713,N_19302);
or UO_1617 (O_1617,N_24293,N_22046);
and UO_1618 (O_1618,N_22140,N_22552);
nor UO_1619 (O_1619,N_22963,N_22377);
and UO_1620 (O_1620,N_23636,N_24814);
and UO_1621 (O_1621,N_20958,N_23518);
xor UO_1622 (O_1622,N_20859,N_23616);
nor UO_1623 (O_1623,N_22612,N_23738);
and UO_1624 (O_1624,N_24222,N_18824);
and UO_1625 (O_1625,N_19737,N_24298);
or UO_1626 (O_1626,N_23855,N_20036);
nor UO_1627 (O_1627,N_23899,N_19104);
nand UO_1628 (O_1628,N_19628,N_20651);
and UO_1629 (O_1629,N_21202,N_23251);
nor UO_1630 (O_1630,N_20260,N_21184);
and UO_1631 (O_1631,N_23810,N_23622);
nor UO_1632 (O_1632,N_19089,N_24812);
nor UO_1633 (O_1633,N_21064,N_18914);
nor UO_1634 (O_1634,N_24082,N_23018);
and UO_1635 (O_1635,N_20764,N_22737);
nor UO_1636 (O_1636,N_20986,N_20438);
and UO_1637 (O_1637,N_21586,N_20560);
nor UO_1638 (O_1638,N_24939,N_20684);
xnor UO_1639 (O_1639,N_19287,N_21054);
and UO_1640 (O_1640,N_18798,N_24587);
xor UO_1641 (O_1641,N_23882,N_23905);
and UO_1642 (O_1642,N_19126,N_24693);
or UO_1643 (O_1643,N_22979,N_24564);
xor UO_1644 (O_1644,N_22216,N_21720);
or UO_1645 (O_1645,N_19011,N_20281);
nand UO_1646 (O_1646,N_24783,N_19133);
nor UO_1647 (O_1647,N_23161,N_21702);
and UO_1648 (O_1648,N_22088,N_20807);
nor UO_1649 (O_1649,N_23109,N_20890);
nand UO_1650 (O_1650,N_23260,N_24820);
nand UO_1651 (O_1651,N_21343,N_23212);
and UO_1652 (O_1652,N_23440,N_20113);
nor UO_1653 (O_1653,N_19716,N_23591);
or UO_1654 (O_1654,N_19878,N_24784);
nor UO_1655 (O_1655,N_18931,N_19889);
nor UO_1656 (O_1656,N_21282,N_24050);
nand UO_1657 (O_1657,N_20527,N_22197);
nand UO_1658 (O_1658,N_23842,N_21963);
nor UO_1659 (O_1659,N_23653,N_22973);
nand UO_1660 (O_1660,N_23912,N_19994);
and UO_1661 (O_1661,N_19208,N_22865);
nor UO_1662 (O_1662,N_19560,N_23977);
and UO_1663 (O_1663,N_21991,N_22458);
xnor UO_1664 (O_1664,N_22201,N_19349);
or UO_1665 (O_1665,N_21204,N_18928);
nand UO_1666 (O_1666,N_23438,N_23111);
nor UO_1667 (O_1667,N_24973,N_20533);
and UO_1668 (O_1668,N_21477,N_20961);
and UO_1669 (O_1669,N_19283,N_19224);
xor UO_1670 (O_1670,N_24746,N_20519);
xnor UO_1671 (O_1671,N_22906,N_19100);
or UO_1672 (O_1672,N_22252,N_24003);
and UO_1673 (O_1673,N_23253,N_19047);
nand UO_1674 (O_1674,N_20346,N_19659);
nand UO_1675 (O_1675,N_20167,N_19318);
nor UO_1676 (O_1676,N_21260,N_20150);
or UO_1677 (O_1677,N_23757,N_22717);
nand UO_1678 (O_1678,N_23557,N_21886);
or UO_1679 (O_1679,N_22406,N_21473);
or UO_1680 (O_1680,N_18902,N_19782);
nand UO_1681 (O_1681,N_21866,N_19859);
or UO_1682 (O_1682,N_19714,N_20331);
nand UO_1683 (O_1683,N_23734,N_19521);
nor UO_1684 (O_1684,N_22684,N_19179);
nor UO_1685 (O_1685,N_21053,N_19954);
nor UO_1686 (O_1686,N_24857,N_19410);
and UO_1687 (O_1687,N_23079,N_24443);
xnor UO_1688 (O_1688,N_24155,N_19320);
and UO_1689 (O_1689,N_24604,N_24797);
and UO_1690 (O_1690,N_20480,N_21888);
or UO_1691 (O_1691,N_22742,N_24482);
nor UO_1692 (O_1692,N_24113,N_21019);
nand UO_1693 (O_1693,N_20756,N_22915);
nand UO_1694 (O_1694,N_20877,N_24224);
nand UO_1695 (O_1695,N_19099,N_20786);
nand UO_1696 (O_1696,N_19806,N_23292);
nand UO_1697 (O_1697,N_24821,N_22646);
nor UO_1698 (O_1698,N_20211,N_23775);
or UO_1699 (O_1699,N_24021,N_20675);
and UO_1700 (O_1700,N_19997,N_22231);
nor UO_1701 (O_1701,N_23515,N_22006);
and UO_1702 (O_1702,N_24568,N_18918);
or UO_1703 (O_1703,N_22971,N_24899);
nand UO_1704 (O_1704,N_19474,N_22373);
and UO_1705 (O_1705,N_24525,N_20570);
and UO_1706 (O_1706,N_23935,N_24740);
or UO_1707 (O_1707,N_19176,N_18780);
nor UO_1708 (O_1708,N_23451,N_22386);
and UO_1709 (O_1709,N_21482,N_22893);
nor UO_1710 (O_1710,N_18769,N_20079);
nand UO_1711 (O_1711,N_20682,N_21458);
nor UO_1712 (O_1712,N_20161,N_21391);
nand UO_1713 (O_1713,N_18899,N_19501);
or UO_1714 (O_1714,N_20866,N_21483);
or UO_1715 (O_1715,N_20811,N_21331);
or UO_1716 (O_1716,N_24344,N_21516);
nor UO_1717 (O_1717,N_19231,N_20498);
and UO_1718 (O_1718,N_20394,N_22218);
and UO_1719 (O_1719,N_22544,N_23444);
nand UO_1720 (O_1720,N_24558,N_20829);
xor UO_1721 (O_1721,N_22888,N_20511);
nand UO_1722 (O_1722,N_19861,N_21534);
or UO_1723 (O_1723,N_21192,N_19860);
or UO_1724 (O_1724,N_22056,N_21048);
and UO_1725 (O_1725,N_20868,N_24231);
or UO_1726 (O_1726,N_21896,N_24156);
and UO_1727 (O_1727,N_21408,N_23475);
and UO_1728 (O_1728,N_24275,N_24569);
nand UO_1729 (O_1729,N_24699,N_19174);
and UO_1730 (O_1730,N_23964,N_22177);
and UO_1731 (O_1731,N_19282,N_19957);
and UO_1732 (O_1732,N_20528,N_21140);
nor UO_1733 (O_1733,N_18844,N_19945);
nand UO_1734 (O_1734,N_19799,N_23057);
xor UO_1735 (O_1735,N_20038,N_24211);
xor UO_1736 (O_1736,N_23805,N_20382);
nor UO_1737 (O_1737,N_24901,N_22330);
or UO_1738 (O_1738,N_22796,N_20857);
xnor UO_1739 (O_1739,N_24058,N_22686);
nor UO_1740 (O_1740,N_24963,N_19528);
and UO_1741 (O_1741,N_19943,N_21688);
nand UO_1742 (O_1742,N_19791,N_19893);
nor UO_1743 (O_1743,N_19213,N_21742);
and UO_1744 (O_1744,N_19692,N_24923);
xnor UO_1745 (O_1745,N_24067,N_20039);
and UO_1746 (O_1746,N_24887,N_24346);
nor UO_1747 (O_1747,N_21514,N_23496);
nand UO_1748 (O_1748,N_19612,N_22990);
xor UO_1749 (O_1749,N_19480,N_19654);
or UO_1750 (O_1750,N_19037,N_21427);
nand UO_1751 (O_1751,N_24239,N_22957);
and UO_1752 (O_1752,N_20745,N_18961);
nor UO_1753 (O_1753,N_22337,N_22607);
or UO_1754 (O_1754,N_19014,N_24427);
nor UO_1755 (O_1755,N_20209,N_20177);
xor UO_1756 (O_1756,N_19950,N_21255);
and UO_1757 (O_1757,N_23172,N_21350);
nand UO_1758 (O_1758,N_22185,N_20202);
nand UO_1759 (O_1759,N_20876,N_21984);
and UO_1760 (O_1760,N_18916,N_18884);
and UO_1761 (O_1761,N_20271,N_22250);
or UO_1762 (O_1762,N_20253,N_19052);
nor UO_1763 (O_1763,N_19496,N_19775);
nand UO_1764 (O_1764,N_22269,N_24143);
nand UO_1765 (O_1765,N_22909,N_23155);
or UO_1766 (O_1766,N_21789,N_21820);
xor UO_1767 (O_1767,N_24831,N_20719);
nand UO_1768 (O_1768,N_23547,N_21588);
xnor UO_1769 (O_1769,N_23938,N_19833);
or UO_1770 (O_1770,N_22687,N_20855);
or UO_1771 (O_1771,N_18838,N_20644);
and UO_1772 (O_1772,N_19689,N_19988);
and UO_1773 (O_1773,N_22496,N_22486);
and UO_1774 (O_1774,N_20291,N_21658);
and UO_1775 (O_1775,N_24410,N_21773);
nand UO_1776 (O_1776,N_20363,N_23727);
nor UO_1777 (O_1777,N_22213,N_24180);
nand UO_1778 (O_1778,N_23113,N_18809);
and UO_1779 (O_1779,N_23914,N_23722);
or UO_1780 (O_1780,N_21732,N_24624);
xnor UO_1781 (O_1781,N_24280,N_21914);
and UO_1782 (O_1782,N_22864,N_24002);
nor UO_1783 (O_1783,N_24878,N_24284);
or UO_1784 (O_1784,N_19547,N_22839);
nor UO_1785 (O_1785,N_19273,N_20365);
or UO_1786 (O_1786,N_23586,N_20288);
nand UO_1787 (O_1787,N_23071,N_20073);
nand UO_1788 (O_1788,N_22483,N_24245);
nand UO_1789 (O_1789,N_23840,N_23735);
or UO_1790 (O_1790,N_24660,N_19076);
nand UO_1791 (O_1791,N_22262,N_20230);
or UO_1792 (O_1792,N_20566,N_20596);
or UO_1793 (O_1793,N_22537,N_24542);
or UO_1794 (O_1794,N_22609,N_19974);
and UO_1795 (O_1795,N_20945,N_23584);
nor UO_1796 (O_1796,N_23931,N_22284);
or UO_1797 (O_1797,N_21689,N_21860);
and UO_1798 (O_1798,N_23953,N_19315);
xnor UO_1799 (O_1799,N_20949,N_21578);
nand UO_1800 (O_1800,N_19642,N_23257);
and UO_1801 (O_1801,N_22597,N_19268);
or UO_1802 (O_1802,N_22460,N_22015);
nand UO_1803 (O_1803,N_23188,N_21032);
nand UO_1804 (O_1804,N_24870,N_19087);
and UO_1805 (O_1805,N_20791,N_20583);
nor UO_1806 (O_1806,N_18843,N_19491);
nand UO_1807 (O_1807,N_21806,N_19507);
or UO_1808 (O_1808,N_20721,N_22360);
nand UO_1809 (O_1809,N_22435,N_23984);
and UO_1810 (O_1810,N_23053,N_22494);
or UO_1811 (O_1811,N_21366,N_22096);
nor UO_1812 (O_1812,N_24470,N_24478);
nand UO_1813 (O_1813,N_19413,N_18822);
nand UO_1814 (O_1814,N_19590,N_21001);
or UO_1815 (O_1815,N_19487,N_21635);
nor UO_1816 (O_1816,N_22474,N_24938);
and UO_1817 (O_1817,N_21567,N_23577);
and UO_1818 (O_1818,N_21274,N_23119);
or UO_1819 (O_1819,N_23009,N_19066);
nand UO_1820 (O_1820,N_23503,N_24052);
nor UO_1821 (O_1821,N_23333,N_20677);
or UO_1822 (O_1822,N_19870,N_24107);
nor UO_1823 (O_1823,N_22431,N_19286);
nand UO_1824 (O_1824,N_24998,N_21372);
or UO_1825 (O_1825,N_21042,N_23870);
nand UO_1826 (O_1826,N_23811,N_20892);
or UO_1827 (O_1827,N_20970,N_23395);
and UO_1828 (O_1828,N_22626,N_24225);
nand UO_1829 (O_1829,N_22908,N_20192);
nor UO_1830 (O_1830,N_24941,N_21226);
or UO_1831 (O_1831,N_22861,N_22619);
xor UO_1832 (O_1832,N_22503,N_21310);
nand UO_1833 (O_1833,N_22678,N_24091);
and UO_1834 (O_1834,N_24585,N_24849);
or UO_1835 (O_1835,N_21954,N_21304);
nor UO_1836 (O_1836,N_20072,N_21870);
nor UO_1837 (O_1837,N_18924,N_23856);
or UO_1838 (O_1838,N_20085,N_22882);
or UO_1839 (O_1839,N_19942,N_24951);
nand UO_1840 (O_1840,N_20050,N_22616);
nor UO_1841 (O_1841,N_23903,N_23178);
or UO_1842 (O_1842,N_19872,N_19767);
xor UO_1843 (O_1843,N_22928,N_24332);
nor UO_1844 (O_1844,N_21631,N_22326);
and UO_1845 (O_1845,N_21760,N_20258);
and UO_1846 (O_1846,N_24261,N_18861);
and UO_1847 (O_1847,N_22782,N_21952);
and UO_1848 (O_1848,N_21024,N_22027);
and UO_1849 (O_1849,N_22398,N_20931);
nand UO_1850 (O_1850,N_21787,N_20506);
or UO_1851 (O_1851,N_19301,N_23495);
nor UO_1852 (O_1852,N_22104,N_19668);
and UO_1853 (O_1853,N_21705,N_19494);
nor UO_1854 (O_1854,N_22060,N_19524);
and UO_1855 (O_1855,N_21877,N_22167);
or UO_1856 (O_1856,N_23344,N_20429);
or UO_1857 (O_1857,N_24290,N_19520);
or UO_1858 (O_1858,N_20747,N_19317);
nor UO_1859 (O_1859,N_24925,N_22080);
and UO_1860 (O_1860,N_24555,N_23679);
nand UO_1861 (O_1861,N_22661,N_23483);
nand UO_1862 (O_1862,N_22819,N_23713);
nor UO_1863 (O_1863,N_24764,N_19907);
or UO_1864 (O_1864,N_24908,N_19048);
nand UO_1865 (O_1865,N_19384,N_24015);
or UO_1866 (O_1866,N_20188,N_24321);
or UO_1867 (O_1867,N_20280,N_21297);
and UO_1868 (O_1868,N_21792,N_24071);
nand UO_1869 (O_1869,N_22042,N_20061);
or UO_1870 (O_1870,N_22454,N_21990);
nand UO_1871 (O_1871,N_19479,N_24655);
nor UO_1872 (O_1872,N_21832,N_20982);
nor UO_1873 (O_1873,N_23996,N_20226);
or UO_1874 (O_1874,N_24418,N_20822);
xnor UO_1875 (O_1875,N_22517,N_18942);
or UO_1876 (O_1876,N_23171,N_24397);
and UO_1877 (O_1877,N_23632,N_19094);
xnor UO_1878 (O_1878,N_24884,N_24098);
nand UO_1879 (O_1879,N_22735,N_18974);
xnor UO_1880 (O_1880,N_19506,N_23309);
nand UO_1881 (O_1881,N_21248,N_23530);
nor UO_1882 (O_1882,N_21370,N_21424);
or UO_1883 (O_1883,N_20620,N_24616);
or UO_1884 (O_1884,N_20580,N_20474);
nor UO_1885 (O_1885,N_24001,N_19419);
or UO_1886 (O_1886,N_22812,N_24620);
nand UO_1887 (O_1887,N_22465,N_23695);
nand UO_1888 (O_1888,N_19726,N_20128);
nand UO_1889 (O_1889,N_23357,N_21776);
or UO_1890 (O_1890,N_21276,N_20255);
nor UO_1891 (O_1891,N_24544,N_19016);
and UO_1892 (O_1892,N_21765,N_21762);
and UO_1893 (O_1893,N_18938,N_19685);
or UO_1894 (O_1894,N_22479,N_18978);
or UO_1895 (O_1895,N_24511,N_24759);
nor UO_1896 (O_1896,N_23773,N_24488);
nand UO_1897 (O_1897,N_19088,N_19247);
nand UO_1898 (O_1898,N_22758,N_18818);
or UO_1899 (O_1899,N_21798,N_24241);
nand UO_1900 (O_1900,N_23791,N_22871);
xor UO_1901 (O_1901,N_19681,N_21626);
nand UO_1902 (O_1902,N_22982,N_23796);
or UO_1903 (O_1903,N_22840,N_22159);
and UO_1904 (O_1904,N_19412,N_24244);
xnor UO_1905 (O_1905,N_20820,N_24638);
nand UO_1906 (O_1906,N_23790,N_21447);
nor UO_1907 (O_1907,N_23963,N_21471);
and UO_1908 (O_1908,N_21293,N_22789);
nor UO_1909 (O_1909,N_21294,N_19482);
nor UO_1910 (O_1910,N_18791,N_20034);
or UO_1911 (O_1911,N_21075,N_22716);
or UO_1912 (O_1912,N_21087,N_23324);
nor UO_1913 (O_1913,N_19809,N_23516);
and UO_1914 (O_1914,N_22232,N_19565);
and UO_1915 (O_1915,N_19381,N_21544);
nor UO_1916 (O_1916,N_21084,N_20571);
and UO_1917 (O_1917,N_21604,N_21452);
nand UO_1918 (O_1918,N_22469,N_20631);
nor UO_1919 (O_1919,N_21150,N_20379);
nor UO_1920 (O_1920,N_23654,N_20234);
and UO_1921 (O_1921,N_19160,N_20295);
nand UO_1922 (O_1922,N_23231,N_24654);
nor UO_1923 (O_1923,N_20621,N_20212);
and UO_1924 (O_1924,N_21404,N_19446);
nor UO_1925 (O_1925,N_23378,N_18878);
nor UO_1926 (O_1926,N_19279,N_21155);
nor UO_1927 (O_1927,N_22770,N_19851);
and UO_1928 (O_1928,N_23561,N_23937);
and UO_1929 (O_1929,N_20705,N_19127);
nand UO_1930 (O_1930,N_23897,N_21739);
and UO_1931 (O_1931,N_19019,N_21196);
nand UO_1932 (O_1932,N_19853,N_19582);
and UO_1933 (O_1933,N_22476,N_24141);
or UO_1934 (O_1934,N_18951,N_21031);
and UO_1935 (O_1935,N_22863,N_24500);
nand UO_1936 (O_1936,N_19025,N_24785);
and UO_1937 (O_1937,N_24969,N_24726);
nand UO_1938 (O_1938,N_20920,N_22614);
nor UO_1939 (O_1939,N_22014,N_24853);
nand UO_1940 (O_1940,N_24958,N_19255);
nand UO_1941 (O_1941,N_21288,N_20094);
nand UO_1942 (O_1942,N_24602,N_20579);
nor UO_1943 (O_1943,N_23876,N_19312);
and UO_1944 (O_1944,N_20701,N_19136);
or UO_1945 (O_1945,N_19561,N_19477);
and UO_1946 (O_1946,N_23936,N_19578);
nor UO_1947 (O_1947,N_19210,N_20804);
or UO_1948 (O_1948,N_22513,N_24851);
nor UO_1949 (O_1949,N_24933,N_19827);
nor UO_1950 (O_1950,N_23639,N_21869);
nor UO_1951 (O_1951,N_24424,N_19852);
and UO_1952 (O_1952,N_23512,N_21900);
xor UO_1953 (O_1953,N_21831,N_24966);
and UO_1954 (O_1954,N_19733,N_23544);
nand UO_1955 (O_1955,N_19694,N_21446);
xnor UO_1956 (O_1956,N_22276,N_20903);
nand UO_1957 (O_1957,N_20446,N_19257);
or UO_1958 (O_1958,N_23032,N_19552);
nor UO_1959 (O_1959,N_20003,N_19151);
nor UO_1960 (O_1960,N_23062,N_22880);
xor UO_1961 (O_1961,N_22473,N_22266);
nand UO_1962 (O_1962,N_23211,N_20044);
and UO_1963 (O_1963,N_20082,N_22745);
nor UO_1964 (O_1964,N_24306,N_23677);
or UO_1965 (O_1965,N_19948,N_20711);
and UO_1966 (O_1966,N_24145,N_21257);
nand UO_1967 (O_1967,N_21722,N_22482);
xnor UO_1968 (O_1968,N_18796,N_20715);
nand UO_1969 (O_1969,N_19599,N_23435);
nand UO_1970 (O_1970,N_24258,N_20991);
or UO_1971 (O_1971,N_23720,N_21533);
and UO_1972 (O_1972,N_22858,N_20157);
xnor UO_1973 (O_1973,N_21170,N_22415);
nand UO_1974 (O_1974,N_20240,N_20995);
xnor UO_1975 (O_1975,N_24665,N_24372);
nor UO_1976 (O_1976,N_23889,N_21661);
and UO_1977 (O_1977,N_20207,N_20909);
nand UO_1978 (O_1978,N_20385,N_22492);
nor UO_1979 (O_1979,N_22150,N_24493);
nor UO_1980 (O_1980,N_20902,N_20515);
nand UO_1981 (O_1981,N_24712,N_24931);
nor UO_1982 (O_1982,N_23425,N_24842);
and UO_1983 (O_1983,N_19670,N_21051);
nor UO_1984 (O_1984,N_22378,N_24567);
nor UO_1985 (O_1985,N_22117,N_24445);
nand UO_1986 (O_1986,N_20247,N_24386);
nand UO_1987 (O_1987,N_22128,N_20634);
and UO_1988 (O_1988,N_19486,N_23325);
and UO_1989 (O_1989,N_20617,N_20913);
nand UO_1990 (O_1990,N_23838,N_24526);
nor UO_1991 (O_1991,N_24610,N_24728);
nand UO_1992 (O_1992,N_23502,N_24754);
and UO_1993 (O_1993,N_21999,N_22929);
nand UO_1994 (O_1994,N_23256,N_19021);
or UO_1995 (O_1995,N_20450,N_22992);
or UO_1996 (O_1996,N_23660,N_20047);
nor UO_1997 (O_1997,N_19734,N_24954);
and UO_1998 (O_1998,N_19243,N_19162);
nand UO_1999 (O_1999,N_23989,N_20403);
nor UO_2000 (O_2000,N_23304,N_24678);
xnor UO_2001 (O_2001,N_23233,N_18792);
or UO_2002 (O_2002,N_21721,N_21439);
and UO_2003 (O_2003,N_20992,N_19996);
nand UO_2004 (O_2004,N_24129,N_21179);
nor UO_2005 (O_2005,N_21098,N_21666);
xor UO_2006 (O_2006,N_20907,N_22896);
or UO_2007 (O_2007,N_24668,N_23288);
or UO_2008 (O_2008,N_19682,N_20774);
nand UO_2009 (O_2009,N_22744,N_19216);
and UO_2010 (O_2010,N_21252,N_18816);
nand UO_2011 (O_2011,N_22249,N_24663);
nor UO_2012 (O_2012,N_19417,N_19554);
nand UO_2013 (O_2013,N_19152,N_21139);
nand UO_2014 (O_2014,N_21389,N_24102);
or UO_2015 (O_2015,N_24212,N_22318);
nor UO_2016 (O_2016,N_22178,N_20704);
and UO_2017 (O_2017,N_22124,N_23331);
nor UO_2018 (O_2018,N_19164,N_21718);
and UO_2019 (O_2019,N_23277,N_19292);
and UO_2020 (O_2020,N_20134,N_23442);
nand UO_2021 (O_2021,N_22317,N_20277);
and UO_2022 (O_2022,N_18850,N_19729);
and UO_2023 (O_2023,N_22948,N_23752);
or UO_2024 (O_2024,N_23087,N_19964);
nand UO_2025 (O_2025,N_23479,N_21499);
xor UO_2026 (O_2026,N_21004,N_22449);
or UO_2027 (O_2027,N_23462,N_22553);
nand UO_2028 (O_2028,N_20680,N_22041);
and UO_2029 (O_2029,N_21644,N_24069);
nand UO_2030 (O_2030,N_22525,N_21281);
nor UO_2031 (O_2031,N_22191,N_23986);
nor UO_2032 (O_2032,N_20040,N_21884);
nand UO_2033 (O_2033,N_23201,N_24760);
nand UO_2034 (O_2034,N_18836,N_20304);
or UO_2035 (O_2035,N_18768,N_20389);
or UO_2036 (O_2036,N_24738,N_22596);
nor UO_2037 (O_2037,N_20372,N_22703);
or UO_2038 (O_2038,N_21091,N_21190);
and UO_2039 (O_2039,N_23559,N_24350);
nor UO_2040 (O_2040,N_18810,N_23867);
and UO_2041 (O_2041,N_23383,N_24622);
and UO_2042 (O_2042,N_24178,N_19344);
or UO_2043 (O_2043,N_19403,N_19577);
or UO_2044 (O_2044,N_24253,N_21839);
nand UO_2045 (O_2045,N_20722,N_20243);
and UO_2046 (O_2046,N_21848,N_23296);
or UO_2047 (O_2047,N_20310,N_24507);
or UO_2048 (O_2048,N_20173,N_19256);
and UO_2049 (O_2049,N_19393,N_23241);
nand UO_2050 (O_2050,N_23423,N_22206);
and UO_2051 (O_2051,N_19285,N_18795);
and UO_2052 (O_2052,N_24181,N_23566);
or UO_2053 (O_2053,N_23051,N_21131);
nand UO_2054 (O_2054,N_24304,N_22243);
nor UO_2055 (O_2055,N_23318,N_20996);
nor UO_2056 (O_2056,N_24592,N_20993);
or UO_2057 (O_2057,N_19272,N_19442);
or UO_2058 (O_2058,N_20194,N_22131);
nand UO_2059 (O_2059,N_22518,N_24112);
and UO_2060 (O_2060,N_24536,N_20339);
nand UO_2061 (O_2061,N_24491,N_21385);
and UO_2062 (O_2062,N_19563,N_19382);
or UO_2063 (O_2063,N_22017,N_24072);
and UO_2064 (O_2064,N_20969,N_24235);
nand UO_2065 (O_2065,N_23031,N_21682);
nand UO_2066 (O_2066,N_22916,N_22399);
nand UO_2067 (O_2067,N_22625,N_19051);
and UO_2068 (O_2068,N_21011,N_21639);
nand UO_2069 (O_2069,N_23204,N_22275);
nor UO_2070 (O_2070,N_20400,N_23597);
or UO_2071 (O_2071,N_24910,N_20458);
and UO_2072 (O_2072,N_22485,N_19193);
nor UO_2073 (O_2073,N_23362,N_23913);
xor UO_2074 (O_2074,N_19415,N_19258);
nand UO_2075 (O_2075,N_23934,N_22205);
and UO_2076 (O_2076,N_19069,N_23340);
nand UO_2077 (O_2077,N_22677,N_19720);
nand UO_2078 (O_2078,N_23910,N_19111);
nor UO_2079 (O_2079,N_22010,N_20558);
nand UO_2080 (O_2080,N_22970,N_20605);
nand UO_2081 (O_2081,N_20559,N_21339);
nor UO_2082 (O_2082,N_22809,N_23817);
nand UO_2083 (O_2083,N_22767,N_19831);
and UO_2084 (O_2084,N_20779,N_20465);
or UO_2085 (O_2085,N_20568,N_23108);
nand UO_2086 (O_2086,N_22860,N_23692);
or UO_2087 (O_2087,N_19667,N_24955);
xnor UO_2088 (O_2088,N_23524,N_24264);
nor UO_2089 (O_2089,N_20557,N_19849);
or UO_2090 (O_2090,N_22634,N_23090);
and UO_2091 (O_2091,N_20170,N_19618);
or UO_2092 (O_2092,N_21412,N_20434);
nand UO_2093 (O_2093,N_21057,N_22491);
xnor UO_2094 (O_2094,N_19680,N_23917);
and UO_2095 (O_2095,N_23096,N_21786);
or UO_2096 (O_2096,N_20430,N_23802);
and UO_2097 (O_2097,N_24097,N_20622);
or UO_2098 (O_2098,N_19823,N_20637);
or UO_2099 (O_2099,N_20083,N_20109);
or UO_2100 (O_2100,N_20398,N_18887);
nand UO_2101 (O_2101,N_22966,N_24059);
nand UO_2102 (O_2102,N_20155,N_24557);
nor UO_2103 (O_2103,N_22099,N_21974);
or UO_2104 (O_2104,N_19012,N_19239);
or UO_2105 (O_2105,N_23298,N_19584);
and UO_2106 (O_2106,N_24873,N_23568);
or UO_2107 (O_2107,N_23389,N_23745);
and UO_2108 (O_2108,N_23180,N_23640);
nor UO_2109 (O_2109,N_19139,N_24720);
nand UO_2110 (O_2110,N_24038,N_21490);
or UO_2111 (O_2111,N_21456,N_23193);
and UO_2112 (O_2112,N_19149,N_20445);
xnor UO_2113 (O_2113,N_21898,N_22012);
and UO_2114 (O_2114,N_20377,N_19644);
and UO_2115 (O_2115,N_20702,N_21698);
and UO_2116 (O_2116,N_23824,N_23445);
and UO_2117 (O_2117,N_18774,N_23268);
and UO_2118 (O_2118,N_23375,N_24162);
nand UO_2119 (O_2119,N_20146,N_21510);
or UO_2120 (O_2120,N_23269,N_22331);
nor UO_2121 (O_2121,N_24100,N_19428);
nand UO_2122 (O_2122,N_22233,N_19871);
or UO_2123 (O_2123,N_24170,N_19557);
and UO_2124 (O_2124,N_19252,N_21027);
or UO_2125 (O_2125,N_21188,N_20303);
and UO_2126 (O_2126,N_21111,N_22207);
and UO_2127 (O_2127,N_22508,N_19306);
or UO_2128 (O_2128,N_19758,N_19916);
nor UO_2129 (O_2129,N_23476,N_20768);
and UO_2130 (O_2130,N_18999,N_19776);
nand UO_2131 (O_2131,N_20141,N_21775);
nor UO_2132 (O_2132,N_21993,N_24448);
and UO_2133 (O_2133,N_23456,N_21410);
or UO_2134 (O_2134,N_22268,N_24523);
nor UO_2135 (O_2135,N_21785,N_18814);
nand UO_2136 (O_2136,N_20965,N_21351);
nand UO_2137 (O_2137,N_20850,N_19968);
and UO_2138 (O_2138,N_20827,N_22273);
or UO_2139 (O_2139,N_22988,N_22523);
nand UO_2140 (O_2140,N_22930,N_23343);
nand UO_2141 (O_2141,N_24083,N_18856);
nand UO_2142 (O_2142,N_22118,N_22962);
nand UO_2143 (O_2143,N_22741,N_21079);
and UO_2144 (O_2144,N_18846,N_19542);
or UO_2145 (O_2145,N_18776,N_21363);
and UO_2146 (O_2146,N_24869,N_21143);
nor UO_2147 (O_2147,N_20404,N_21345);
xor UO_2148 (O_2148,N_23160,N_22032);
and UO_2149 (O_2149,N_19116,N_21794);
nor UO_2150 (O_2150,N_21694,N_24626);
nand UO_2151 (O_2151,N_21632,N_24215);
nor UO_2152 (O_2152,N_22447,N_23663);
and UO_2153 (O_2153,N_21814,N_23510);
nor UO_2154 (O_2154,N_22624,N_24392);
nand UO_2155 (O_2155,N_19725,N_18908);
and UO_2156 (O_2156,N_24512,N_24737);
and UO_2157 (O_2157,N_19962,N_23575);
nand UO_2158 (O_2158,N_19165,N_19197);
nand UO_2159 (O_2159,N_22633,N_20159);
nand UO_2160 (O_2160,N_24475,N_20537);
and UO_2161 (O_2161,N_20531,N_23393);
xor UO_2162 (O_2162,N_22996,N_19875);
and UO_2163 (O_2163,N_19611,N_23896);
and UO_2164 (O_2164,N_19421,N_22227);
nand UO_2165 (O_2165,N_21174,N_20599);
and UO_2166 (O_2166,N_22565,N_24676);
nand UO_2167 (O_2167,N_22866,N_20741);
or UO_2168 (O_2168,N_23714,N_18904);
or UO_2169 (O_2169,N_21828,N_21484);
xor UO_2170 (O_2170,N_23243,N_22879);
nor UO_2171 (O_2171,N_19388,N_19904);
nor UO_2172 (O_2172,N_21916,N_20204);
or UO_2173 (O_2173,N_20944,N_19118);
and UO_2174 (O_2174,N_20898,N_24101);
xnor UO_2175 (O_2175,N_19488,N_21547);
nor UO_2176 (O_2176,N_24464,N_19390);
nor UO_2177 (O_2177,N_22532,N_20830);
nand UO_2178 (O_2178,N_18903,N_24928);
nor UO_2179 (O_2179,N_24139,N_23255);
nand UO_2180 (O_2180,N_23312,N_21261);
and UO_2181 (O_2181,N_22193,N_19157);
nor UO_2182 (O_2182,N_24486,N_23699);
nand UO_2183 (O_2183,N_20283,N_23787);
or UO_2184 (O_2184,N_20332,N_24988);
nor UO_2185 (O_2185,N_21414,N_18821);
xnor UO_2186 (O_2186,N_23196,N_22437);
nor UO_2187 (O_2187,N_20947,N_24793);
xnor UO_2188 (O_2188,N_19214,N_24950);
and UO_2189 (O_2189,N_19350,N_20550);
and UO_2190 (O_2190,N_18807,N_24650);
and UO_2191 (O_2191,N_19760,N_20915);
nand UO_2192 (O_2192,N_20998,N_20227);
and UO_2193 (O_2193,N_19541,N_24992);
and UO_2194 (O_2194,N_18801,N_20131);
nand UO_2195 (O_2195,N_21554,N_24357);
nor UO_2196 (O_2196,N_24313,N_24374);
and UO_2197 (O_2197,N_20865,N_19934);
nor UO_2198 (O_2198,N_21182,N_24762);
nor UO_2199 (O_2199,N_23780,N_23465);
nand UO_2200 (O_2200,N_23182,N_18955);
or UO_2201 (O_2201,N_20973,N_19406);
nor UO_2202 (O_2202,N_23460,N_22883);
nand UO_2203 (O_2203,N_21819,N_21752);
or UO_2204 (O_2204,N_20478,N_24292);
or UO_2205 (O_2205,N_23861,N_24351);
nor UO_2206 (O_2206,N_22501,N_24407);
nand UO_2207 (O_2207,N_19380,N_24666);
nand UO_2208 (O_2208,N_19864,N_22063);
nand UO_2209 (O_2209,N_19438,N_19600);
nor UO_2210 (O_2210,N_20932,N_21864);
or UO_2211 (O_2211,N_23901,N_20408);
nor UO_2212 (O_2212,N_23954,N_24461);
xnor UO_2213 (O_2213,N_24084,N_19063);
nand UO_2214 (O_2214,N_19033,N_23581);
nor UO_2215 (O_2215,N_22947,N_22311);
xor UO_2216 (O_2216,N_20639,N_24325);
or UO_2217 (O_2217,N_23414,N_19054);
nor UO_2218 (O_2218,N_20724,N_20396);
nand UO_2219 (O_2219,N_19352,N_24917);
and UO_2220 (O_2220,N_24004,N_24179);
and UO_2221 (O_2221,N_23793,N_19015);
nor UO_2222 (O_2222,N_23311,N_19078);
nand UO_2223 (O_2223,N_20658,N_22364);
or UO_2224 (O_2224,N_20732,N_22149);
or UO_2225 (O_2225,N_23555,N_23881);
nand UO_2226 (O_2226,N_23704,N_19502);
nand UO_2227 (O_2227,N_24062,N_23237);
nand UO_2228 (O_2228,N_19519,N_23869);
or UO_2229 (O_2229,N_20840,N_23026);
or UO_2230 (O_2230,N_23386,N_24158);
nand UO_2231 (O_2231,N_20106,N_24667);
nor UO_2232 (O_2232,N_19747,N_24074);
or UO_2233 (O_2233,N_21362,N_19695);
nor UO_2234 (O_2234,N_21713,N_18891);
or UO_2235 (O_2235,N_21296,N_20685);
nor UO_2236 (O_2236,N_19837,N_24573);
nand UO_2237 (O_2237,N_20520,N_19673);
nand UO_2238 (O_2238,N_21636,N_19091);
nor UO_2239 (O_2239,N_21911,N_21015);
and UO_2240 (O_2240,N_23521,N_22282);
nand UO_2241 (O_2241,N_19722,N_20534);
or UO_2242 (O_2242,N_22605,N_21072);
and UO_2243 (O_2243,N_23002,N_22989);
and UO_2244 (O_2244,N_24595,N_24428);
nand UO_2245 (O_2245,N_20748,N_19530);
nor UO_2246 (O_2246,N_22190,N_22379);
and UO_2247 (O_2247,N_23449,N_24203);
and UO_2248 (O_2248,N_24856,N_24791);
nand UO_2249 (O_2249,N_21016,N_23633);
and UO_2250 (O_2250,N_24106,N_22174);
or UO_2251 (O_2251,N_24776,N_20262);
nor UO_2252 (O_2252,N_21791,N_21589);
or UO_2253 (O_2253,N_20491,N_24048);
xor UO_2254 (O_2254,N_18863,N_21325);
or UO_2255 (O_2255,N_20788,N_23553);
nand UO_2256 (O_2256,N_19031,N_22028);
and UO_2257 (O_2257,N_21970,N_21232);
nand UO_2258 (O_2258,N_22872,N_21106);
or UO_2259 (O_2259,N_24111,N_19163);
nor UO_2260 (O_2260,N_22119,N_24379);
nand UO_2261 (O_2261,N_20301,N_20235);
nor UO_2262 (O_2262,N_21241,N_24308);
nand UO_2263 (O_2263,N_21945,N_23368);
nor UO_2264 (O_2264,N_23991,N_19155);
nand UO_2265 (O_2265,N_23848,N_24903);
xor UO_2266 (O_2266,N_23814,N_23505);
nor UO_2267 (O_2267,N_24598,N_21555);
nand UO_2268 (O_2268,N_18873,N_21413);
nor UO_2269 (O_2269,N_19664,N_19020);
nor UO_2270 (O_2270,N_23323,N_20530);
and UO_2271 (O_2271,N_20582,N_24302);
nand UO_2272 (O_2272,N_21384,N_22291);
nor UO_2273 (O_2273,N_20852,N_23216);
and UO_2274 (O_2274,N_21747,N_22591);
xor UO_2275 (O_2275,N_24458,N_21601);
nand UO_2276 (O_2276,N_19569,N_21328);
nor UO_2277 (O_2277,N_20656,N_24430);
nand UO_2278 (O_2278,N_22094,N_23245);
and UO_2279 (O_2279,N_23010,N_22168);
nand UO_2280 (O_2280,N_19589,N_22240);
nand UO_2281 (O_2281,N_18829,N_19454);
or UO_2282 (O_2282,N_19572,N_19346);
and UO_2283 (O_2283,N_19570,N_21641);
or UO_2284 (O_2284,N_23149,N_21272);
xor UO_2285 (O_2285,N_21178,N_19990);
and UO_2286 (O_2286,N_20406,N_21163);
or UO_2287 (O_2287,N_22516,N_23742);
xor UO_2288 (O_2288,N_24548,N_19855);
or UO_2289 (O_2289,N_18808,N_23908);
or UO_2290 (O_2290,N_20074,N_24561);
and UO_2291 (O_2291,N_20144,N_22000);
or UO_2292 (O_2292,N_21818,N_19387);
nand UO_2293 (O_2293,N_22130,N_24014);
and UO_2294 (O_2294,N_20647,N_19207);
nand UO_2295 (O_2295,N_24637,N_24848);
nand UO_2296 (O_2296,N_22792,N_18760);
and UO_2297 (O_2297,N_20059,N_21522);
and UO_2298 (O_2298,N_19448,N_20413);
nand UO_2299 (O_2299,N_22422,N_21893);
and UO_2300 (O_2300,N_24563,N_21964);
and UO_2301 (O_2301,N_24326,N_21733);
nand UO_2302 (O_2302,N_20051,N_20238);
xnor UO_2303 (O_2303,N_23626,N_19291);
nand UO_2304 (O_2304,N_20978,N_20938);
nor UO_2305 (O_2305,N_23152,N_22007);
nand UO_2306 (O_2306,N_21324,N_20275);
and UO_2307 (O_2307,N_20473,N_23387);
or UO_2308 (O_2308,N_19032,N_20300);
and UO_2309 (O_2309,N_23351,N_24417);
and UO_2310 (O_2310,N_19641,N_20306);
nand UO_2311 (O_2311,N_21148,N_22823);
nor UO_2312 (O_2312,N_23545,N_19717);
or UO_2313 (O_2313,N_19721,N_22543);
or UO_2314 (O_2314,N_19043,N_24529);
xor UO_2315 (O_2315,N_24730,N_22808);
xor UO_2316 (O_2316,N_22418,N_20181);
xor UO_2317 (O_2317,N_21671,N_22229);
and UO_2318 (O_2318,N_21748,N_22220);
and UO_2319 (O_2319,N_24748,N_20362);
nor UO_2320 (O_2320,N_23104,N_19643);
and UO_2321 (O_2321,N_20081,N_24159);
nor UO_2322 (O_2322,N_20863,N_23696);
and UO_2323 (O_2323,N_19461,N_22914);
nand UO_2324 (O_2324,N_21100,N_23558);
nor UO_2325 (O_2325,N_21915,N_24816);
xnor UO_2326 (O_2326,N_23758,N_20484);
nand UO_2327 (O_2327,N_23453,N_24061);
nor UO_2328 (O_2328,N_24916,N_21289);
nand UO_2329 (O_2329,N_19137,N_20007);
or UO_2330 (O_2330,N_24311,N_22788);
nor UO_2331 (O_2331,N_23823,N_22401);
xnor UO_2332 (O_2332,N_19967,N_19992);
or UO_2333 (O_2333,N_20285,N_24539);
and UO_2334 (O_2334,N_21712,N_22376);
nand UO_2335 (O_2335,N_20225,N_19691);
xnor UO_2336 (O_2336,N_24423,N_22466);
and UO_2337 (O_2337,N_19905,N_23365);
or UO_2338 (O_2338,N_22816,N_21519);
nor UO_2339 (O_2339,N_20941,N_20415);
nand UO_2340 (O_2340,N_20635,N_22413);
or UO_2341 (O_2341,N_22417,N_22675);
or UO_2342 (O_2342,N_20156,N_19189);
and UO_2343 (O_2343,N_20585,N_22804);
nor UO_2344 (O_2344,N_20125,N_24453);
or UO_2345 (O_2345,N_20356,N_21373);
xor UO_2346 (O_2346,N_21662,N_24168);
and UO_2347 (O_2347,N_19657,N_19928);
or UO_2348 (O_2348,N_24045,N_20743);
xnor UO_2349 (O_2349,N_21406,N_19531);
or UO_2350 (O_2350,N_23276,N_23806);
nand UO_2351 (O_2351,N_21467,N_23452);
and UO_2352 (O_2352,N_21734,N_20004);
and UO_2353 (O_2353,N_24398,N_22053);
or UO_2354 (O_2354,N_24017,N_20541);
or UO_2355 (O_2355,N_21142,N_22902);
and UO_2356 (O_2356,N_18911,N_22538);
and UO_2357 (O_2357,N_24775,N_22132);
and UO_2358 (O_2358,N_24652,N_22825);
nor UO_2359 (O_2359,N_21904,N_23205);
nand UO_2360 (O_2360,N_23921,N_21305);
xor UO_2361 (O_2361,N_18775,N_22719);
nor UO_2362 (O_2362,N_21591,N_19882);
nand UO_2363 (O_2363,N_20444,N_20254);
xor UO_2364 (O_2364,N_22935,N_24584);
and UO_2365 (O_2365,N_21811,N_19591);
or UO_2366 (O_2366,N_22462,N_22955);
and UO_2367 (O_2367,N_23164,N_19464);
and UO_2368 (O_2368,N_18841,N_24639);
nor UO_2369 (O_2369,N_23543,N_21756);
xor UO_2370 (O_2370,N_24436,N_21551);
and UO_2371 (O_2371,N_24149,N_20990);
and UO_2372 (O_2372,N_23800,N_19913);
or UO_2373 (O_2373,N_20660,N_23669);
nand UO_2374 (O_2374,N_20041,N_22103);
nor UO_2375 (O_2375,N_20885,N_22171);
nor UO_2376 (O_2376,N_20352,N_21186);
and UO_2377 (O_2377,N_22322,N_21736);
nor UO_2378 (O_2378,N_24965,N_21058);
nand UO_2379 (O_2379,N_22588,N_22878);
nor UO_2380 (O_2380,N_19386,N_20246);
or UO_2381 (O_2381,N_23770,N_23254);
nor UO_2382 (O_2382,N_23853,N_19493);
and UO_2383 (O_2383,N_21771,N_21321);
and UO_2384 (O_2384,N_19090,N_22993);
or UO_2385 (O_2385,N_21696,N_21538);
nor UO_2386 (O_2386,N_20765,N_21236);
nand UO_2387 (O_2387,N_22807,N_18830);
nand UO_2388 (O_2388,N_19917,N_20825);
and UO_2389 (O_2389,N_23405,N_20853);
and UO_2390 (O_2390,N_22689,N_22752);
nand UO_2391 (O_2391,N_21531,N_23821);
nor UO_2392 (O_2392,N_20891,N_23785);
and UO_2393 (O_2393,N_21537,N_20510);
nor UO_2394 (O_2394,N_22487,N_23589);
nand UO_2395 (O_2395,N_20314,N_22534);
xor UO_2396 (O_2396,N_19329,N_23379);
nor UO_2397 (O_2397,N_20354,N_21885);
nor UO_2398 (O_2398,N_23077,N_21356);
or UO_2399 (O_2399,N_24366,N_24193);
xnor UO_2400 (O_2400,N_21844,N_22024);
and UO_2401 (O_2401,N_24172,N_21822);
xnor UO_2402 (O_2402,N_21726,N_22941);
nor UO_2403 (O_2403,N_21112,N_23744);
or UO_2404 (O_2404,N_21487,N_20591);
and UO_2405 (O_2405,N_20727,N_23602);
or UO_2406 (O_2406,N_18954,N_20753);
and UO_2407 (O_2407,N_24553,N_24065);
or UO_2408 (O_2408,N_24200,N_24879);
nor UO_2409 (O_2409,N_21041,N_23055);
nand UO_2410 (O_2410,N_24194,N_21488);
and UO_2411 (O_2411,N_23924,N_18823);
and UO_2412 (O_2412,N_24249,N_23043);
nor UO_2413 (O_2413,N_24623,N_24796);
xor UO_2414 (O_2414,N_24722,N_23015);
and UO_2415 (O_2415,N_24185,N_21147);
and UO_2416 (O_2416,N_21399,N_22453);
nand UO_2417 (O_2417,N_24167,N_23360);
or UO_2418 (O_2418,N_23687,N_24301);
and UO_2419 (O_2419,N_24209,N_21138);
or UO_2420 (O_2420,N_24092,N_19122);
nand UO_2421 (O_2421,N_24964,N_21678);
xor UO_2422 (O_2422,N_18945,N_22662);
and UO_2423 (O_2423,N_19158,N_21481);
nor UO_2424 (O_2424,N_23388,N_22481);
nand UO_2425 (O_2425,N_21028,N_23706);
nand UO_2426 (O_2426,N_23385,N_20717);
and UO_2427 (O_2427,N_21216,N_23369);
xnor UO_2428 (O_2428,N_20739,N_24997);
nor UO_2429 (O_2429,N_20483,N_22303);
xor UO_2430 (O_2430,N_22734,N_20063);
nor UO_2431 (O_2431,N_19394,N_18905);
nand UO_2432 (O_2432,N_20691,N_21933);
and UO_2433 (O_2433,N_19296,N_21670);
nor UO_2434 (O_2434,N_24496,N_23278);
or UO_2435 (O_2435,N_23159,N_20604);
or UO_2436 (O_2436,N_24806,N_24844);
xnor UO_2437 (O_2437,N_22754,N_21708);
or UO_2438 (O_2438,N_24363,N_23039);
and UO_2439 (O_2439,N_19172,N_24380);
or UO_2440 (O_2440,N_21625,N_23997);
and UO_2441 (O_2441,N_23721,N_22549);
xor UO_2442 (O_2442,N_24684,N_19932);
xor UO_2443 (O_2443,N_24641,N_19310);
xor UO_2444 (O_2444,N_19113,N_19391);
nor UO_2445 (O_2445,N_19537,N_18906);
and UO_2446 (O_2446,N_24271,N_21464);
or UO_2447 (O_2447,N_23631,N_23202);
or UO_2448 (O_2448,N_20726,N_20563);
and UO_2449 (O_2449,N_21322,N_19702);
xor UO_2450 (O_2450,N_19376,N_20090);
and UO_2451 (O_2451,N_22402,N_24056);
nor UO_2452 (O_2452,N_22639,N_19300);
nand UO_2453 (O_2453,N_21161,N_21265);
nor UO_2454 (O_2454,N_24317,N_19953);
and UO_2455 (O_2455,N_22407,N_18922);
nand UO_2456 (O_2456,N_19336,N_20105);
or UO_2457 (O_2457,N_24743,N_21767);
and UO_2458 (O_2458,N_21379,N_22102);
nand UO_2459 (O_2459,N_19906,N_23781);
xnor UO_2460 (O_2460,N_20552,N_23929);
or UO_2461 (O_2461,N_18979,N_20718);
nand UO_2462 (O_2462,N_22314,N_19539);
nor UO_2463 (O_2463,N_19338,N_24518);
and UO_2464 (O_2464,N_24318,N_19017);
nand UO_2465 (O_2465,N_21959,N_20013);
or UO_2466 (O_2466,N_22428,N_21361);
or UO_2467 (O_2467,N_24979,N_22146);
nor UO_2468 (O_2468,N_19203,N_21352);
or UO_2469 (O_2469,N_19625,N_19581);
nor UO_2470 (O_2470,N_24247,N_18875);
nor UO_2471 (O_2471,N_19544,N_19596);
nand UO_2472 (O_2472,N_19993,N_21559);
nand UO_2473 (O_2473,N_19883,N_24303);
nand UO_2474 (O_2474,N_24591,N_24540);
or UO_2475 (O_2475,N_24051,N_22793);
or UO_2476 (O_2476,N_23068,N_23743);
nand UO_2477 (O_2477,N_19466,N_18966);
nor UO_2478 (O_2478,N_22711,N_24824);
nor UO_2479 (O_2479,N_20819,N_19671);
or UO_2480 (O_2480,N_19634,N_23644);
nand UO_2481 (O_2481,N_21905,N_24452);
and UO_2482 (O_2482,N_22600,N_20495);
and UO_2483 (O_2483,N_21419,N_19034);
nand UO_2484 (O_2484,N_24370,N_23443);
or UO_2485 (O_2485,N_20286,N_18915);
nor UO_2486 (O_2486,N_24246,N_20883);
nand UO_2487 (O_2487,N_19465,N_18893);
and UO_2488 (O_2488,N_24590,N_24510);
nand UO_2489 (O_2489,N_20431,N_19110);
nand UO_2490 (O_2490,N_24996,N_23354);
and UO_2491 (O_2491,N_22556,N_20674);
xor UO_2492 (O_2492,N_24843,N_21985);
or UO_2493 (O_2493,N_23392,N_23694);
nand UO_2494 (O_2494,N_19982,N_22857);
and UO_2495 (O_2495,N_20461,N_22604);
and UO_2496 (O_2496,N_20178,N_20759);
nand UO_2497 (O_2497,N_22061,N_19674);
and UO_2498 (O_2498,N_24706,N_22372);
nor UO_2499 (O_2499,N_23998,N_21600);
nor UO_2500 (O_2500,N_21919,N_21249);
and UO_2501 (O_2501,N_20153,N_21197);
nor UO_2502 (O_2502,N_19304,N_21897);
nor UO_2503 (O_2503,N_18993,N_23198);
or UO_2504 (O_2504,N_23355,N_19331);
or UO_2505 (O_2505,N_23421,N_21663);
nand UO_2506 (O_2506,N_20554,N_19327);
and UO_2507 (O_2507,N_20833,N_20567);
nor UO_2508 (O_2508,N_24546,N_20026);
xnor UO_2509 (O_2509,N_18987,N_20099);
xor UO_2510 (O_2510,N_22424,N_23001);
nor UO_2511 (O_2511,N_19187,N_23420);
or UO_2512 (O_2512,N_19922,N_19141);
and UO_2513 (O_2513,N_22867,N_24761);
and UO_2514 (O_2514,N_24778,N_23124);
or UO_2515 (O_2515,N_20472,N_19361);
nand UO_2516 (O_2516,N_21254,N_23715);
or UO_2517 (O_2517,N_20757,N_18834);
or UO_2518 (O_2518,N_21269,N_21587);
xor UO_2519 (O_2519,N_20397,N_21940);
nor UO_2520 (O_2520,N_24095,N_19398);
and UO_2521 (O_2521,N_20425,N_19707);
and UO_2522 (O_2522,N_23000,N_23081);
and UO_2523 (O_2523,N_20841,N_21616);
and UO_2524 (O_2524,N_21498,N_22567);
nor UO_2525 (O_2525,N_24944,N_22158);
nor UO_2526 (O_2526,N_18872,N_24919);
xnor UO_2527 (O_2527,N_21675,N_22299);
nor UO_2528 (O_2528,N_20505,N_23885);
nor UO_2529 (O_2529,N_18800,N_23845);
or UO_2530 (O_2530,N_18797,N_24505);
xnor UO_2531 (O_2531,N_19605,N_18827);
or UO_2532 (O_2532,N_22446,N_18958);
and UO_2533 (O_2533,N_19773,N_20296);
and UO_2534 (O_2534,N_20667,N_23454);
or UO_2535 (O_2535,N_24420,N_22209);
xor UO_2536 (O_2536,N_21730,N_24270);
nor UO_2537 (O_2537,N_24904,N_24242);
nand UO_2538 (O_2538,N_20490,N_23279);
and UO_2539 (O_2539,N_19923,N_23807);
nor UO_2540 (O_2540,N_20725,N_19458);
nor UO_2541 (O_2541,N_23820,N_22239);
nor UO_2542 (O_2542,N_21073,N_19724);
or UO_2543 (O_2543,N_21552,N_19001);
xor UO_2544 (O_2544,N_21307,N_19072);
and UO_2545 (O_2545,N_19965,N_19610);
nand UO_2546 (O_2546,N_21777,N_21969);
and UO_2547 (O_2547,N_24586,N_24087);
and UO_2548 (O_2548,N_21992,N_23798);
nor UO_2549 (O_2549,N_20985,N_24077);
nand UO_2550 (O_2550,N_23551,N_19416);
xor UO_2551 (O_2551,N_21634,N_22182);
xnor UO_2552 (O_2552,N_23235,N_20971);
nand UO_2553 (O_2553,N_19796,N_23637);
nor UO_2554 (O_2554,N_20874,N_21812);
nor UO_2555 (O_2555,N_20826,N_24310);
nor UO_2556 (O_2556,N_20917,N_22602);
or UO_2557 (O_2557,N_24309,N_20060);
and UO_2558 (O_2558,N_23762,N_20174);
nand UO_2559 (O_2559,N_24913,N_22780);
nand UO_2560 (O_2560,N_23332,N_22480);
nor UO_2561 (O_2561,N_21623,N_20983);
and UO_2562 (O_2562,N_19754,N_23979);
nor UO_2563 (O_2563,N_23552,N_21764);
or UO_2564 (O_2564,N_19366,N_19332);
and UO_2565 (O_2565,N_22016,N_19319);
xnor UO_2566 (O_2566,N_22101,N_24833);
and UO_2567 (O_2567,N_20845,N_24541);
nor UO_2568 (O_2568,N_20981,N_22722);
nor UO_2569 (O_2569,N_20046,N_23628);
and UO_2570 (O_2570,N_19790,N_19615);
and UO_2571 (O_2571,N_24680,N_18771);
nor UO_2572 (O_2572,N_23623,N_20539);
nor UO_2573 (O_2573,N_19783,N_21242);
and UO_2574 (O_2574,N_23579,N_19929);
and UO_2575 (O_2575,N_20014,N_22445);
and UO_2576 (O_2576,N_21476,N_23157);
or UO_2577 (O_2577,N_21569,N_20266);
xnor UO_2578 (O_2578,N_21853,N_20942);
or UO_2579 (O_2579,N_23101,N_20977);
nand UO_2580 (O_2580,N_23619,N_23613);
nand UO_2581 (O_2581,N_23611,N_23114);
and UO_2582 (O_2582,N_24718,N_22034);
xor UO_2583 (O_2583,N_19772,N_21429);
nand UO_2584 (O_2584,N_23313,N_19669);
xor UO_2585 (O_2585,N_19868,N_22083);
xnor UO_2586 (O_2586,N_21622,N_21231);
and UO_2587 (O_2587,N_23167,N_20010);
or UO_2588 (O_2588,N_21318,N_19295);
or UO_2589 (O_2589,N_21683,N_22797);
and UO_2590 (O_2590,N_23348,N_21134);
nor UO_2591 (O_2591,N_23875,N_24477);
or UO_2592 (O_2592,N_24867,N_24805);
or UO_2593 (O_2593,N_20542,N_19259);
nand UO_2594 (O_2594,N_19128,N_19981);
nor UO_2595 (O_2595,N_20171,N_24986);
and UO_2596 (O_2596,N_22764,N_19748);
and UO_2597 (O_2597,N_18998,N_21146);
xor UO_2598 (O_2598,N_24333,N_19580);
or UO_2599 (O_2599,N_21220,N_23128);
or UO_2600 (O_2600,N_23549,N_23441);
or UO_2601 (O_2601,N_19337,N_20217);
and UO_2602 (O_2602,N_24940,N_19759);
and UO_2603 (O_2603,N_21354,N_24388);
nor UO_2604 (O_2604,N_22241,N_21104);
nand UO_2605 (O_2605,N_20761,N_19703);
and UO_2606 (O_2606,N_20193,N_20390);
nor UO_2607 (O_2607,N_22050,N_21026);
nor UO_2608 (O_2608,N_18982,N_22954);
nand UO_2609 (O_2609,N_19824,N_19900);
nand UO_2610 (O_2610,N_22093,N_23173);
nand UO_2611 (O_2611,N_23536,N_24068);
nor UO_2612 (O_2612,N_23060,N_18898);
and UO_2613 (O_2613,N_19144,N_20149);
nor UO_2614 (O_2614,N_23382,N_20279);
and UO_2615 (O_2615,N_24583,N_18933);
nand UO_2616 (O_2616,N_18788,N_21692);
nor UO_2617 (O_2617,N_20507,N_19921);
or UO_2618 (O_2618,N_19559,N_20676);
and UO_2619 (O_2619,N_24846,N_23878);
and UO_2620 (O_2620,N_23843,N_23832);
xor UO_2621 (O_2621,N_22070,N_22656);
nand UO_2622 (O_2622,N_23115,N_21315);
nor UO_2623 (O_2623,N_20142,N_20847);
nor UO_2624 (O_2624,N_23918,N_20790);
or UO_2625 (O_2625,N_19588,N_24441);
and UO_2626 (O_2626,N_21107,N_19335);
nor UO_2627 (O_2627,N_21195,N_22328);
and UO_2628 (O_2628,N_24771,N_20120);
or UO_2629 (O_2629,N_21103,N_19977);
nor UO_2630 (O_2630,N_22784,N_22222);
or UO_2631 (O_2631,N_20744,N_21007);
or UO_2632 (O_2632,N_22749,N_23857);
nand UO_2633 (O_2633,N_20699,N_21397);
nor UO_2634 (O_2634,N_22359,N_19023);
nor UO_2635 (O_2635,N_24562,N_22560);
nor UO_2636 (O_2636,N_20386,N_21441);
xor UO_2637 (O_2637,N_19750,N_20943);
and UO_2638 (O_2638,N_23594,N_20350);
and UO_2639 (O_2639,N_23883,N_20091);
xnor UO_2640 (O_2640,N_23993,N_20287);
and UO_2641 (O_2641,N_22110,N_23482);
xnor UO_2642 (O_2642,N_18896,N_19082);
and UO_2643 (O_2643,N_23705,N_23517);
and UO_2644 (O_2644,N_19368,N_19186);
and UO_2645 (O_2645,N_21157,N_23297);
nor UO_2646 (O_2646,N_22411,N_18811);
nor UO_2647 (O_2647,N_24755,N_24891);
and UO_2648 (O_2648,N_19060,N_21951);
or UO_2649 (O_2649,N_20816,N_19846);
nor UO_2650 (O_2650,N_24189,N_22363);
xor UO_2651 (O_2651,N_19313,N_24076);
nor UO_2652 (O_2652,N_19771,N_21808);
xnor UO_2653 (O_2653,N_23801,N_23634);
nand UO_2654 (O_2654,N_24835,N_19844);
nand UO_2655 (O_2655,N_23849,N_20778);
or UO_2656 (O_2656,N_21470,N_20195);
nand UO_2657 (O_2657,N_22830,N_22370);
or UO_2658 (O_2658,N_21494,N_21931);
or UO_2659 (O_2659,N_22581,N_20532);
nand UO_2660 (O_2660,N_18895,N_24826);
and UO_2661 (O_2661,N_21491,N_19505);
or UO_2662 (O_2662,N_22215,N_19585);
nor UO_2663 (O_2663,N_19363,N_23107);
nor UO_2664 (O_2664,N_20447,N_24018);
nor UO_2665 (O_2665,N_20955,N_23892);
xor UO_2666 (O_2666,N_19261,N_23915);
nor UO_2667 (O_2667,N_24362,N_22120);
nor UO_2668 (O_2668,N_21285,N_19434);
nand UO_2669 (O_2669,N_24845,N_24447);
nor UO_2670 (O_2670,N_19785,N_22981);
or UO_2671 (O_2671,N_20921,N_24081);
xnor UO_2672 (O_2672,N_22405,N_21633);
nor UO_2673 (O_2673,N_24369,N_20169);
or UO_2674 (O_2674,N_22077,N_20124);
or UO_2675 (O_2675,N_20290,N_19180);
or UO_2676 (O_2676,N_20564,N_23429);
or UO_2677 (O_2677,N_21009,N_23567);
nand UO_2678 (O_2678,N_21431,N_22289);
nor UO_2679 (O_2679,N_22510,N_24205);
and UO_2680 (O_2680,N_21063,N_22653);
or UO_2681 (O_2681,N_21613,N_23207);
nand UO_2682 (O_2682,N_18779,N_23314);
or UO_2683 (O_2683,N_23035,N_22911);
xor UO_2684 (O_2684,N_19598,N_24915);
nand UO_2685 (O_2685,N_19863,N_23430);
xnor UO_2686 (O_2686,N_19958,N_21549);
or UO_2687 (O_2687,N_21440,N_24381);
nor UO_2688 (O_2688,N_22442,N_22155);
xor UO_2689 (O_2689,N_19651,N_19042);
nand UO_2690 (O_2690,N_24909,N_22004);
xnor UO_2691 (O_2691,N_21229,N_22196);
and UO_2692 (O_2692,N_20752,N_19422);
or UO_2693 (O_2693,N_21596,N_23224);
or UO_2694 (O_2694,N_19813,N_21926);
or UO_2695 (O_2695,N_19786,N_23945);
or UO_2696 (O_2696,N_24368,N_20267);
or UO_2697 (O_2697,N_19234,N_20619);
or UO_2698 (O_2698,N_24024,N_18985);
or UO_2699 (O_2699,N_20008,N_24632);
and UO_2700 (O_2700,N_20697,N_23709);
nor UO_2701 (O_2701,N_24342,N_24039);
and UO_2702 (O_2702,N_20694,N_20049);
or UO_2703 (O_2703,N_19606,N_19215);
nor UO_2704 (O_2704,N_18885,N_19794);
nor UO_2705 (O_2705,N_24648,N_23990);
and UO_2706 (O_2706,N_19937,N_19039);
nor UO_2707 (O_2707,N_21856,N_23310);
or UO_2708 (O_2708,N_22551,N_24559);
nor UO_2709 (O_2709,N_23847,N_24411);
nand UO_2710 (O_2710,N_22059,N_19192);
nand UO_2711 (O_2711,N_24195,N_23731);
and UO_2712 (O_2712,N_19699,N_20526);
or UO_2713 (O_2713,N_20095,N_24481);
and UO_2714 (O_2714,N_18901,N_19220);
nand UO_2715 (O_2715,N_18964,N_24140);
xor UO_2716 (O_2716,N_20407,N_23487);
nand UO_2717 (O_2717,N_19467,N_18926);
nor UO_2718 (O_2718,N_22100,N_23248);
and UO_2719 (O_2719,N_24552,N_19453);
nor UO_2720 (O_2720,N_19742,N_22172);
and UO_2721 (O_2721,N_20777,N_20861);
xor UO_2722 (O_2722,N_24429,N_24789);
nand UO_2723 (O_2723,N_22974,N_18840);
and UO_2724 (O_2724,N_24439,N_20966);
nor UO_2725 (O_2725,N_23166,N_18767);
or UO_2726 (O_2726,N_24132,N_24255);
or UO_2727 (O_2727,N_24701,N_24858);
or UO_2728 (O_2728,N_23229,N_23779);
and UO_2729 (O_2729,N_21766,N_24034);
xor UO_2730 (O_2730,N_22980,N_22356);
nand UO_2731 (O_2731,N_20988,N_23499);
nand UO_2732 (O_2732,N_19092,N_21125);
and UO_2733 (O_2733,N_18975,N_23651);
or UO_2734 (O_2734,N_24528,N_21529);
nand UO_2735 (O_2735,N_24744,N_21774);
or UO_2736 (O_2736,N_22321,N_23337);
nand UO_2737 (O_2737,N_21615,N_24509);
nand UO_2738 (O_2738,N_22354,N_19204);
and UO_2739 (O_2739,N_20503,N_20823);
nor UO_2740 (O_2740,N_18935,N_18783);
and UO_2741 (O_2741,N_23625,N_22152);
nand UO_2742 (O_2742,N_24677,N_22621);
nor UO_2743 (O_2743,N_23974,N_22603);
and UO_2744 (O_2744,N_21955,N_22768);
nor UO_2745 (O_2745,N_23401,N_19941);
nand UO_2746 (O_2746,N_19829,N_23928);
nor UO_2747 (O_2747,N_23825,N_23349);
and UO_2748 (O_2748,N_23652,N_23556);
nand UO_2749 (O_2749,N_19244,N_20775);
nand UO_2750 (O_2750,N_20298,N_24527);
or UO_2751 (O_2751,N_21754,N_24576);
or UO_2752 (O_2752,N_23582,N_19027);
nor UO_2753 (O_2753,N_21262,N_20911);
nor UO_2754 (O_2754,N_18991,N_21040);
or UO_2755 (O_2755,N_21398,N_19774);
or UO_2756 (O_2756,N_21518,N_19046);
xor UO_2757 (O_2757,N_22704,N_24545);
and UO_2758 (O_2758,N_22009,N_24176);
or UO_2759 (O_2759,N_20625,N_24890);
and UO_2760 (O_2760,N_20602,N_22707);
and UO_2761 (O_2761,N_19418,N_19517);
nor UO_2762 (O_2762,N_23952,N_19876);
xor UO_2763 (O_2763,N_24803,N_22683);
or UO_2764 (O_2764,N_20294,N_24137);
and UO_2765 (O_2765,N_22901,N_21183);
nand UO_2766 (O_2766,N_23203,N_23708);
and UO_2767 (O_2767,N_24609,N_20158);
nor UO_2768 (O_2768,N_23574,N_19124);
nor UO_2769 (O_2769,N_23837,N_23129);
or UO_2770 (O_2770,N_22571,N_20763);
xnor UO_2771 (O_2771,N_19154,N_23215);
nor UO_2772 (O_2772,N_23434,N_23030);
nor UO_2773 (O_2773,N_20755,N_23327);
or UO_2774 (O_2774,N_19175,N_24572);
xor UO_2775 (O_2775,N_24704,N_24799);
or UO_2776 (O_2776,N_18965,N_21887);
nor UO_2777 (O_2777,N_20033,N_22264);
nor UO_2778 (O_2778,N_19597,N_23474);
and UO_2779 (O_2779,N_19738,N_19235);
nand UO_2780 (O_2780,N_22606,N_21059);
and UO_2781 (O_2781,N_19254,N_20391);
nor UO_2782 (O_2782,N_21415,N_21090);
nand UO_2783 (O_2783,N_20529,N_20954);
or UO_2784 (O_2784,N_24861,N_22511);
or UO_2785 (O_2785,N_19515,N_21479);
nor UO_2786 (O_2786,N_19339,N_19622);
nor UO_2787 (O_2787,N_22035,N_23363);
and UO_2788 (O_2788,N_20772,N_21629);
and UO_2789 (O_2789,N_20272,N_23322);
or UO_2790 (O_2790,N_19150,N_24435);
nor UO_2791 (O_2791,N_20440,N_24133);
and UO_2792 (O_2792,N_21443,N_21511);
and UO_2793 (O_2793,N_19246,N_24356);
nand UO_2794 (O_2794,N_22561,N_22667);
and UO_2795 (O_2795,N_19768,N_21302);
or UO_2796 (O_2796,N_20068,N_24033);
nor UO_2797 (O_2797,N_23668,N_20364);
or UO_2798 (O_2798,N_22736,N_19424);
nor UO_2799 (O_2799,N_19166,N_21874);
nor UO_2800 (O_2800,N_22256,N_19044);
nand UO_2801 (O_2801,N_21141,N_19803);
nand UO_2802 (O_2802,N_23596,N_23398);
and UO_2803 (O_2803,N_21695,N_19067);
nand UO_2804 (O_2804,N_22260,N_24108);
and UO_2805 (O_2805,N_22694,N_22592);
nor UO_2806 (O_2806,N_20509,N_21283);
xnor UO_2807 (O_2807,N_20317,N_21719);
or UO_2808 (O_2808,N_24307,N_19984);
nor UO_2809 (O_2809,N_22855,N_23271);
nand UO_2810 (O_2810,N_23774,N_23601);
nand UO_2811 (O_2811,N_23238,N_24710);
nor UO_2812 (O_2812,N_24138,N_24751);
nand UO_2813 (O_2813,N_19266,N_23195);
nand UO_2814 (O_2814,N_24070,N_22577);
nor UO_2815 (O_2815,N_20798,N_19407);
and UO_2816 (O_2816,N_18880,N_19492);
nor UO_2817 (O_2817,N_23667,N_21935);
nor UO_2818 (O_2818,N_22430,N_23647);
and UO_2819 (O_2819,N_20551,N_20324);
or UO_2820 (O_2820,N_21086,N_21165);
nor UO_2821 (O_2821,N_19684,N_22670);
nor UO_2822 (O_2822,N_18983,N_23733);
nand UO_2823 (O_2823,N_19309,N_21585);
nand UO_2824 (O_2824,N_24146,N_21815);
nor UO_2825 (O_2825,N_19485,N_23088);
or UO_2826 (O_2826,N_21566,N_22183);
and UO_2827 (O_2827,N_24974,N_20670);
nand UO_2828 (O_2828,N_22338,N_20456);
and UO_2829 (O_2829,N_22884,N_23879);
and UO_2830 (O_2830,N_24506,N_23489);
and UO_2831 (O_2831,N_20627,N_19764);
or UO_2832 (O_2832,N_23259,N_23391);
nor UO_2833 (O_2833,N_21124,N_24570);
and UO_2834 (O_2834,N_19909,N_20064);
and UO_2835 (O_2835,N_23956,N_22669);
xor UO_2836 (O_2836,N_21228,N_23664);
nor UO_2837 (O_2837,N_24697,N_20813);
nand UO_2838 (O_2838,N_22029,N_24709);
nor UO_2839 (O_2839,N_23782,N_23522);
or UO_2840 (O_2840,N_22391,N_21478);
or UO_2841 (O_2841,N_19055,N_24080);
and UO_2842 (O_2842,N_23508,N_22986);
xor UO_2843 (O_2843,N_19918,N_24252);
nand UO_2844 (O_2844,N_23866,N_21867);
and UO_2845 (O_2845,N_19109,N_22499);
or UO_2846 (O_2846,N_23648,N_20337);
nor UO_2847 (O_2847,N_24121,N_22771);
nand UO_2848 (O_2848,N_20486,N_23819);
or UO_2849 (O_2849,N_22869,N_18973);
and UO_2850 (O_2850,N_20518,N_21256);
nand UO_2851 (O_2851,N_24025,N_21119);
and UO_2852 (O_2852,N_20250,N_20187);
or UO_2853 (O_2853,N_23074,N_22274);
and UO_2854 (O_2854,N_23328,N_23353);
or UO_2855 (O_2855,N_18805,N_23472);
nor UO_2856 (O_2856,N_19478,N_21535);
nor UO_2857 (O_2857,N_21573,N_22221);
nand UO_2858 (O_2858,N_24719,N_21796);
nand UO_2859 (O_2859,N_21668,N_18833);
or UO_2860 (O_2860,N_22692,N_22886);
and UO_2861 (O_2861,N_24968,N_22685);
nor UO_2862 (O_2862,N_18803,N_24262);
xor UO_2863 (O_2863,N_19237,N_21769);
nand UO_2864 (O_2864,N_21973,N_22367);
or UO_2865 (O_2865,N_23263,N_21660);
nand UO_2866 (O_2866,N_18858,N_24088);
nor UO_2867 (O_2867,N_19325,N_23190);
nand UO_2868 (O_2868,N_20367,N_21387);
and UO_2869 (O_2869,N_21871,N_24364);
or UO_2870 (O_2870,N_23218,N_19811);
and UO_2871 (O_2871,N_20460,N_18894);
and UO_2872 (O_2872,N_20716,N_21083);
xnor UO_2873 (O_2873,N_19516,N_20776);
nor UO_2874 (O_2874,N_23020,N_20417);
nand UO_2875 (O_2875,N_23433,N_19297);
and UO_2876 (O_2876,N_23662,N_24123);
nand UO_2877 (O_2877,N_19999,N_18766);
nand UO_2878 (O_2878,N_20808,N_24177);
nor UO_2879 (O_2879,N_20152,N_23301);
nor UO_2880 (O_2880,N_23909,N_21956);
nor UO_2881 (O_2881,N_22895,N_22025);
or UO_2882 (O_2882,N_24809,N_20766);
nand UO_2883 (O_2883,N_21654,N_24985);
nor UO_2884 (O_2884,N_21899,N_22815);
or UO_2885 (O_2885,N_18981,N_24338);
and UO_2886 (O_2886,N_22170,N_24182);
or UO_2887 (O_2887,N_22312,N_21092);
nor UO_2888 (O_2888,N_21565,N_23169);
nor UO_2889 (O_2889,N_20315,N_22333);
and UO_2890 (O_2890,N_21783,N_23234);
xor UO_2891 (O_2891,N_24152,N_22546);
or UO_2892 (O_2892,N_22098,N_24456);
and UO_2893 (O_2893,N_22838,N_22841);
xor UO_2894 (O_2894,N_21115,N_23726);
and UO_2895 (O_2895,N_19627,N_23294);
nand UO_2896 (O_2896,N_24073,N_24434);
or UO_2897 (O_2897,N_22835,N_22905);
nor UO_2898 (O_2898,N_21548,N_22659);
and UO_2899 (O_2899,N_24810,N_19367);
nor UO_2900 (O_2900,N_24685,N_21800);
and UO_2901 (O_2901,N_24384,N_20894);
nor UO_2902 (O_2902,N_20441,N_20912);
nand UO_2903 (O_2903,N_19232,N_20452);
and UO_2904 (O_2904,N_24921,N_21612);
and UO_2905 (O_2905,N_23671,N_20640);
or UO_2906 (O_2906,N_23534,N_22145);
nand UO_2907 (O_2907,N_24440,N_23868);
or UO_2908 (O_2908,N_23067,N_24935);
nor UO_2909 (O_2909,N_20922,N_19739);
and UO_2910 (O_2910,N_23808,N_21599);
nor UO_2911 (O_2911,N_18934,N_21238);
xor UO_2912 (O_2912,N_23464,N_23133);
nand UO_2913 (O_2913,N_24468,N_19426);
or UO_2914 (O_2914,N_21055,N_21506);
nand UO_2915 (O_2915,N_20803,N_19093);
nor UO_2916 (O_2916,N_23511,N_22072);
or UO_2917 (O_2917,N_21731,N_19779);
or UO_2918 (O_2918,N_24032,N_23334);
xor UO_2919 (O_2919,N_18881,N_24786);
nand UO_2920 (O_2920,N_23478,N_22541);
and UO_2921 (O_2921,N_23469,N_20366);
nor UO_2922 (O_2922,N_18927,N_18963);
and UO_2923 (O_2923,N_21123,N_22760);
xnor UO_2924 (O_2924,N_24322,N_19818);
or UO_2925 (O_2925,N_21892,N_19107);
nand UO_2926 (O_2926,N_20632,N_18849);
or UO_2927 (O_2927,N_21691,N_24393);
nor UO_2928 (O_2928,N_24157,N_21287);
xnor UO_2929 (O_2929,N_20432,N_20895);
and UO_2930 (O_2930,N_23852,N_22568);
xnor UO_2931 (O_2931,N_21837,N_24060);
and UO_2932 (O_2932,N_23197,N_24153);
or UO_2933 (O_2933,N_19518,N_20309);
and UO_2934 (O_2934,N_21824,N_24767);
and UO_2935 (O_2935,N_18839,N_20269);
nor UO_2936 (O_2936,N_20708,N_20785);
nand UO_2937 (O_2937,N_20137,N_23017);
nand UO_2938 (O_2938,N_21784,N_20359);
nor UO_2939 (O_2939,N_19700,N_22968);
xnor UO_2940 (O_2940,N_20437,N_20031);
or UO_2941 (O_2941,N_24090,N_22724);
or UO_2942 (O_2942,N_19241,N_18889);
nor UO_2943 (O_2943,N_22166,N_22983);
nor UO_2944 (O_2944,N_20163,N_21029);
nor UO_2945 (O_2945,N_20466,N_21036);
and UO_2946 (O_2946,N_22305,N_21561);
or UO_2947 (O_2947,N_23608,N_19079);
and UO_2948 (O_2948,N_19316,N_21606);
or UO_2949 (O_2949,N_21221,N_19143);
or UO_2950 (O_2950,N_24399,N_19148);
nor UO_2951 (O_2951,N_24647,N_20451);
xnor UO_2952 (O_2952,N_22084,N_20369);
and UO_2953 (O_2953,N_18897,N_19847);
or UO_2954 (O_2954,N_21416,N_20555);
and UO_2955 (O_2955,N_19655,N_21259);
nand UO_2956 (O_2956,N_20276,N_23006);
and UO_2957 (O_2957,N_23600,N_24636);
and UO_2958 (O_2958,N_19330,N_24286);
nor UO_2959 (O_2959,N_22164,N_20818);
nand UO_2960 (O_2960,N_21835,N_21950);
and UO_2961 (O_2961,N_24395,N_22924);
or UO_2962 (O_2962,N_24929,N_20655);
and UO_2963 (O_2963,N_24124,N_21979);
nand UO_2964 (O_2964,N_22246,N_23272);
and UO_2965 (O_2965,N_21701,N_23571);
or UO_2966 (O_2966,N_24296,N_22759);
nand UO_2967 (O_2967,N_22047,N_24498);
nand UO_2968 (O_2968,N_22630,N_24210);
nand UO_2969 (O_2969,N_24695,N_23025);
xnor UO_2970 (O_2970,N_19927,N_21109);
xnor UO_2971 (O_2971,N_23784,N_22067);
nor UO_2972 (O_2972,N_21917,N_21129);
or UO_2973 (O_2973,N_19614,N_23450);
nand UO_2974 (O_2974,N_21652,N_19364);
and UO_2975 (O_2975,N_19002,N_23827);
xnor UO_2976 (O_2976,N_22940,N_22294);
nand UO_2977 (O_2977,N_24863,N_19931);
and UO_2978 (O_2978,N_22564,N_20521);
and UO_2979 (O_2979,N_21199,N_23127);
or UO_2980 (O_2980,N_23244,N_20514);
or UO_2981 (O_2981,N_22245,N_19533);
nand UO_2982 (O_2982,N_24089,N_20525);
nand UO_2983 (O_2983,N_19887,N_19395);
or UO_2984 (O_2984,N_21365,N_20135);
nor UO_2985 (O_2985,N_22978,N_19970);
nand UO_2986 (O_2986,N_24402,N_24213);
xor UO_2987 (O_2987,N_19510,N_22432);
and UO_2988 (O_2988,N_19880,N_21393);
nor UO_2989 (O_2989,N_22355,N_24990);
or UO_2990 (O_2990,N_20231,N_19008);
nand UO_2991 (O_2991,N_23024,N_22031);
and UO_2992 (O_2992,N_19392,N_22922);
or UO_2993 (O_2993,N_21159,N_22939);
nand UO_2994 (O_2994,N_21222,N_19400);
nand UO_2995 (O_2995,N_19567,N_23072);
or UO_2996 (O_2996,N_22521,N_23767);
nor UO_2997 (O_2997,N_20843,N_24519);
and UO_2998 (O_2998,N_21268,N_22628);
or UO_2999 (O_2999,N_19808,N_23145);
endmodule