module basic_500_3000_500_4_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_406,In_453);
nor U1 (N_1,In_308,In_87);
or U2 (N_2,In_284,In_184);
xnor U3 (N_3,In_246,In_195);
nor U4 (N_4,In_28,In_319);
and U5 (N_5,In_289,In_89);
and U6 (N_6,In_107,In_4);
nor U7 (N_7,In_128,In_463);
nand U8 (N_8,In_467,In_133);
or U9 (N_9,In_456,In_254);
or U10 (N_10,In_143,In_188);
xnor U11 (N_11,In_193,In_174);
or U12 (N_12,In_199,In_340);
nand U13 (N_13,In_230,In_124);
or U14 (N_14,In_106,In_435);
or U15 (N_15,In_335,In_355);
xor U16 (N_16,In_419,In_213);
nor U17 (N_17,In_446,In_336);
or U18 (N_18,In_102,In_327);
xor U19 (N_19,In_339,In_430);
and U20 (N_20,In_383,In_163);
nor U21 (N_21,In_411,In_329);
or U22 (N_22,In_484,In_236);
or U23 (N_23,In_30,In_61);
nor U24 (N_24,In_408,In_167);
or U25 (N_25,In_460,In_196);
or U26 (N_26,In_19,In_239);
and U27 (N_27,In_292,In_423);
nand U28 (N_28,In_377,In_137);
nand U29 (N_29,In_363,In_316);
and U30 (N_30,In_200,In_470);
nor U31 (N_31,In_180,In_114);
or U32 (N_32,In_5,In_313);
xor U33 (N_33,In_439,In_68);
and U34 (N_34,In_277,In_131);
nand U35 (N_35,In_354,In_225);
nand U36 (N_36,In_333,In_175);
or U37 (N_37,In_20,In_479);
and U38 (N_38,In_495,In_165);
nor U39 (N_39,In_219,In_110);
and U40 (N_40,In_265,In_25);
nand U41 (N_41,In_132,In_347);
and U42 (N_42,In_181,In_237);
or U43 (N_43,In_381,In_99);
xnor U44 (N_44,In_357,In_86);
nand U45 (N_45,In_158,In_32);
or U46 (N_46,In_95,In_40);
nor U47 (N_47,In_171,In_371);
nand U48 (N_48,In_125,In_490);
and U49 (N_49,In_187,In_358);
xor U50 (N_50,In_296,In_94);
nor U51 (N_51,In_334,In_288);
nand U52 (N_52,In_191,In_164);
and U53 (N_53,In_396,In_272);
and U54 (N_54,In_303,In_197);
and U55 (N_55,In_461,In_209);
nand U56 (N_56,In_315,In_417);
nor U57 (N_57,In_211,In_192);
or U58 (N_58,In_161,In_389);
and U59 (N_59,In_190,In_444);
nor U60 (N_60,In_27,In_310);
nor U61 (N_61,In_245,In_182);
nand U62 (N_62,In_76,In_370);
xor U63 (N_63,In_449,In_448);
and U64 (N_64,In_320,In_12);
xor U65 (N_65,In_451,In_445);
or U66 (N_66,In_42,In_44);
or U67 (N_67,In_388,In_179);
xnor U68 (N_68,In_323,In_283);
nand U69 (N_69,In_3,In_202);
nand U70 (N_70,In_499,In_255);
xnor U71 (N_71,In_14,In_241);
xnor U72 (N_72,In_261,In_485);
and U73 (N_73,In_465,In_273);
and U74 (N_74,In_349,In_328);
and U75 (N_75,In_356,In_177);
xor U76 (N_76,In_212,In_425);
nand U77 (N_77,In_491,In_100);
or U78 (N_78,In_152,In_198);
xnor U79 (N_79,In_300,In_324);
nand U80 (N_80,In_221,In_475);
and U81 (N_81,In_47,In_274);
xnor U82 (N_82,In_222,In_39);
xnor U83 (N_83,In_437,In_75);
or U84 (N_84,In_157,In_252);
nor U85 (N_85,In_287,In_204);
nor U86 (N_86,In_240,In_194);
and U87 (N_87,In_218,In_380);
nand U88 (N_88,In_186,In_142);
nand U89 (N_89,In_498,In_271);
and U90 (N_90,In_293,In_268);
or U91 (N_91,In_420,In_447);
nor U92 (N_92,In_369,In_264);
nand U93 (N_93,In_97,In_321);
or U94 (N_94,In_96,In_306);
nor U95 (N_95,In_464,In_11);
nand U96 (N_96,In_397,In_140);
nor U97 (N_97,In_80,In_312);
nor U98 (N_98,In_92,In_263);
and U99 (N_99,In_403,In_101);
or U100 (N_100,In_488,In_82);
xnor U101 (N_101,In_353,In_215);
xnor U102 (N_102,In_458,In_122);
xor U103 (N_103,In_432,In_276);
nand U104 (N_104,In_121,In_72);
xor U105 (N_105,In_382,In_496);
xor U106 (N_106,In_466,In_148);
nand U107 (N_107,In_257,In_156);
nand U108 (N_108,In_83,In_427);
or U109 (N_109,In_455,In_112);
nor U110 (N_110,In_441,In_45);
xor U111 (N_111,In_93,In_338);
or U112 (N_112,In_318,In_220);
and U113 (N_113,In_330,In_43);
or U114 (N_114,In_214,In_387);
nand U115 (N_115,In_90,In_88);
nand U116 (N_116,In_375,In_248);
nand U117 (N_117,In_373,In_66);
xnor U118 (N_118,In_365,In_457);
and U119 (N_119,In_251,In_346);
nand U120 (N_120,In_290,In_170);
and U121 (N_121,In_436,In_304);
xor U122 (N_122,In_431,In_325);
or U123 (N_123,In_185,In_150);
nor U124 (N_124,In_36,In_489);
and U125 (N_125,In_376,In_50);
or U126 (N_126,In_281,In_205);
nand U127 (N_127,In_15,In_285);
nor U128 (N_128,In_216,In_149);
nand U129 (N_129,In_41,In_84);
nor U130 (N_130,In_115,In_35);
xnor U131 (N_131,In_414,In_337);
nand U132 (N_132,In_421,In_317);
nor U133 (N_133,In_6,In_2);
nor U134 (N_134,In_223,In_81);
and U135 (N_135,In_483,In_350);
and U136 (N_136,In_208,In_37);
and U137 (N_137,In_123,In_22);
nor U138 (N_138,In_341,In_297);
nor U139 (N_139,In_60,In_229);
nand U140 (N_140,In_279,In_256);
and U141 (N_141,In_393,In_116);
or U142 (N_142,In_429,In_104);
nand U143 (N_143,In_282,In_294);
nor U144 (N_144,In_151,In_78);
nor U145 (N_145,In_24,In_207);
or U146 (N_146,In_138,In_481);
and U147 (N_147,In_259,In_392);
nor U148 (N_148,In_117,In_286);
xor U149 (N_149,In_29,In_31);
and U150 (N_150,In_79,In_10);
or U151 (N_151,In_476,In_309);
xnor U152 (N_152,In_98,In_85);
xnor U153 (N_153,In_352,In_366);
and U154 (N_154,In_53,In_57);
or U155 (N_155,In_301,In_224);
nor U156 (N_156,In_0,In_462);
nand U157 (N_157,In_494,In_409);
nand U158 (N_158,In_343,In_59);
nand U159 (N_159,In_471,In_244);
nor U160 (N_160,In_275,In_127);
and U161 (N_161,In_247,In_233);
xnor U162 (N_162,In_141,In_302);
nor U163 (N_163,In_360,In_326);
xnor U164 (N_164,In_391,In_402);
or U165 (N_165,In_7,In_159);
nand U166 (N_166,In_51,In_332);
nand U167 (N_167,In_270,In_298);
and U168 (N_168,In_487,In_203);
nor U169 (N_169,In_368,In_172);
nor U170 (N_170,In_9,In_242);
nor U171 (N_171,In_52,In_153);
nor U172 (N_172,In_351,In_146);
xor U173 (N_173,In_385,In_226);
and U174 (N_174,In_1,In_109);
xor U175 (N_175,In_443,In_422);
xnor U176 (N_176,In_46,In_413);
nor U177 (N_177,In_56,In_472);
and U178 (N_178,In_16,In_33);
nand U179 (N_179,In_278,In_386);
nand U180 (N_180,In_134,In_348);
nor U181 (N_181,In_394,In_206);
nor U182 (N_182,In_69,In_260);
or U183 (N_183,In_299,In_367);
nand U184 (N_184,In_73,In_361);
nor U185 (N_185,In_452,In_111);
and U186 (N_186,In_17,In_227);
nor U187 (N_187,In_231,In_311);
xnor U188 (N_188,In_201,In_399);
nand U189 (N_189,In_401,In_478);
nor U190 (N_190,In_249,In_65);
xnor U191 (N_191,In_407,In_307);
and U192 (N_192,In_493,In_48);
or U193 (N_193,In_482,In_295);
nand U194 (N_194,In_280,In_364);
xor U195 (N_195,In_468,In_416);
xor U196 (N_196,In_342,In_238);
or U197 (N_197,In_77,In_440);
or U198 (N_198,In_405,In_38);
or U199 (N_199,In_258,In_492);
and U200 (N_200,In_374,In_433);
or U201 (N_201,In_147,In_497);
or U202 (N_202,In_71,In_345);
and U203 (N_203,In_262,In_410);
nand U204 (N_204,In_155,In_145);
or U205 (N_205,In_486,In_176);
xor U206 (N_206,In_129,In_162);
xnor U207 (N_207,In_442,In_438);
nand U208 (N_208,In_217,In_426);
or U209 (N_209,In_395,In_243);
and U210 (N_210,In_210,In_108);
nor U211 (N_211,In_160,In_183);
nand U212 (N_212,In_459,In_34);
or U213 (N_213,In_120,In_154);
xnor U214 (N_214,In_418,In_450);
nand U215 (N_215,In_362,In_266);
nor U216 (N_216,In_378,In_434);
and U217 (N_217,In_267,In_228);
nor U218 (N_218,In_168,In_173);
nand U219 (N_219,In_253,In_269);
or U220 (N_220,In_322,In_62);
nor U221 (N_221,In_135,In_379);
nor U222 (N_222,In_8,In_454);
xnor U223 (N_223,In_344,In_359);
or U224 (N_224,In_314,In_58);
nor U225 (N_225,In_250,In_305);
nor U226 (N_226,In_404,In_113);
nand U227 (N_227,In_130,In_166);
xor U228 (N_228,In_26,In_70);
or U229 (N_229,In_54,In_126);
xor U230 (N_230,In_18,In_412);
nor U231 (N_231,In_477,In_234);
xnor U232 (N_232,In_473,In_372);
and U233 (N_233,In_169,In_67);
nand U234 (N_234,In_49,In_400);
or U235 (N_235,In_415,In_398);
and U236 (N_236,In_331,In_390);
nand U237 (N_237,In_118,In_232);
xor U238 (N_238,In_480,In_291);
xor U239 (N_239,In_13,In_63);
nand U240 (N_240,In_189,In_235);
xor U241 (N_241,In_55,In_23);
nor U242 (N_242,In_469,In_474);
xnor U243 (N_243,In_103,In_91);
xor U244 (N_244,In_136,In_144);
or U245 (N_245,In_178,In_74);
and U246 (N_246,In_105,In_139);
xor U247 (N_247,In_21,In_428);
nor U248 (N_248,In_64,In_384);
nor U249 (N_249,In_119,In_424);
xor U250 (N_250,In_235,In_230);
and U251 (N_251,In_478,In_242);
or U252 (N_252,In_345,In_7);
and U253 (N_253,In_263,In_127);
xor U254 (N_254,In_84,In_492);
nor U255 (N_255,In_247,In_158);
nor U256 (N_256,In_434,In_408);
or U257 (N_257,In_498,In_329);
xnor U258 (N_258,In_137,In_20);
and U259 (N_259,In_387,In_371);
nand U260 (N_260,In_140,In_248);
xor U261 (N_261,In_475,In_282);
nand U262 (N_262,In_15,In_153);
nor U263 (N_263,In_8,In_61);
or U264 (N_264,In_34,In_13);
nor U265 (N_265,In_392,In_401);
nor U266 (N_266,In_475,In_488);
or U267 (N_267,In_286,In_378);
nor U268 (N_268,In_215,In_361);
xnor U269 (N_269,In_389,In_340);
and U270 (N_270,In_450,In_260);
nor U271 (N_271,In_269,In_82);
and U272 (N_272,In_319,In_56);
or U273 (N_273,In_212,In_19);
and U274 (N_274,In_343,In_261);
and U275 (N_275,In_38,In_448);
nand U276 (N_276,In_460,In_313);
nand U277 (N_277,In_298,In_62);
and U278 (N_278,In_228,In_139);
and U279 (N_279,In_398,In_286);
and U280 (N_280,In_25,In_159);
xnor U281 (N_281,In_228,In_190);
and U282 (N_282,In_377,In_356);
and U283 (N_283,In_15,In_281);
and U284 (N_284,In_89,In_249);
and U285 (N_285,In_356,In_447);
xor U286 (N_286,In_141,In_439);
and U287 (N_287,In_378,In_273);
and U288 (N_288,In_379,In_467);
xnor U289 (N_289,In_171,In_414);
xnor U290 (N_290,In_466,In_480);
nand U291 (N_291,In_42,In_188);
xnor U292 (N_292,In_327,In_370);
xor U293 (N_293,In_230,In_301);
nand U294 (N_294,In_360,In_449);
or U295 (N_295,In_481,In_4);
nand U296 (N_296,In_456,In_219);
and U297 (N_297,In_34,In_361);
nor U298 (N_298,In_242,In_221);
or U299 (N_299,In_140,In_498);
xnor U300 (N_300,In_373,In_58);
nand U301 (N_301,In_463,In_57);
or U302 (N_302,In_369,In_116);
and U303 (N_303,In_252,In_204);
nor U304 (N_304,In_220,In_340);
nand U305 (N_305,In_437,In_52);
nor U306 (N_306,In_189,In_344);
nor U307 (N_307,In_342,In_3);
and U308 (N_308,In_164,In_146);
nand U309 (N_309,In_325,In_217);
xnor U310 (N_310,In_350,In_242);
nor U311 (N_311,In_358,In_55);
nor U312 (N_312,In_444,In_293);
nor U313 (N_313,In_445,In_299);
or U314 (N_314,In_313,In_33);
nor U315 (N_315,In_289,In_396);
and U316 (N_316,In_491,In_78);
xnor U317 (N_317,In_284,In_215);
xor U318 (N_318,In_160,In_328);
nand U319 (N_319,In_375,In_363);
xor U320 (N_320,In_8,In_79);
xor U321 (N_321,In_125,In_194);
or U322 (N_322,In_209,In_214);
nor U323 (N_323,In_99,In_248);
xnor U324 (N_324,In_9,In_399);
and U325 (N_325,In_185,In_26);
or U326 (N_326,In_10,In_277);
and U327 (N_327,In_17,In_110);
xor U328 (N_328,In_302,In_115);
or U329 (N_329,In_195,In_39);
or U330 (N_330,In_381,In_126);
xnor U331 (N_331,In_257,In_170);
nand U332 (N_332,In_272,In_31);
nor U333 (N_333,In_38,In_206);
xor U334 (N_334,In_234,In_324);
or U335 (N_335,In_58,In_498);
nor U336 (N_336,In_322,In_451);
nand U337 (N_337,In_167,In_25);
xor U338 (N_338,In_85,In_302);
and U339 (N_339,In_147,In_322);
or U340 (N_340,In_389,In_193);
nor U341 (N_341,In_465,In_36);
or U342 (N_342,In_96,In_339);
and U343 (N_343,In_407,In_195);
xor U344 (N_344,In_301,In_465);
nand U345 (N_345,In_293,In_51);
nor U346 (N_346,In_188,In_88);
nor U347 (N_347,In_327,In_174);
and U348 (N_348,In_109,In_225);
nor U349 (N_349,In_18,In_447);
and U350 (N_350,In_178,In_346);
or U351 (N_351,In_359,In_486);
nor U352 (N_352,In_339,In_115);
xor U353 (N_353,In_201,In_96);
xor U354 (N_354,In_31,In_318);
nor U355 (N_355,In_42,In_261);
nand U356 (N_356,In_53,In_497);
nand U357 (N_357,In_184,In_354);
xnor U358 (N_358,In_301,In_249);
xnor U359 (N_359,In_163,In_294);
nor U360 (N_360,In_441,In_321);
xnor U361 (N_361,In_416,In_33);
and U362 (N_362,In_167,In_350);
xnor U363 (N_363,In_29,In_182);
nand U364 (N_364,In_201,In_2);
nor U365 (N_365,In_140,In_469);
nor U366 (N_366,In_2,In_415);
nor U367 (N_367,In_281,In_34);
or U368 (N_368,In_347,In_76);
nor U369 (N_369,In_58,In_309);
and U370 (N_370,In_251,In_57);
xnor U371 (N_371,In_367,In_387);
or U372 (N_372,In_26,In_476);
xor U373 (N_373,In_179,In_329);
or U374 (N_374,In_27,In_293);
xnor U375 (N_375,In_463,In_423);
and U376 (N_376,In_484,In_12);
nand U377 (N_377,In_107,In_161);
and U378 (N_378,In_459,In_409);
or U379 (N_379,In_44,In_321);
xor U380 (N_380,In_345,In_394);
nand U381 (N_381,In_299,In_323);
nor U382 (N_382,In_443,In_45);
xnor U383 (N_383,In_52,In_347);
or U384 (N_384,In_457,In_318);
nand U385 (N_385,In_144,In_132);
xor U386 (N_386,In_477,In_413);
nor U387 (N_387,In_39,In_409);
or U388 (N_388,In_80,In_414);
xor U389 (N_389,In_288,In_350);
nand U390 (N_390,In_95,In_449);
and U391 (N_391,In_408,In_358);
nor U392 (N_392,In_429,In_110);
or U393 (N_393,In_133,In_264);
xor U394 (N_394,In_272,In_366);
nand U395 (N_395,In_48,In_260);
xor U396 (N_396,In_238,In_327);
nand U397 (N_397,In_46,In_118);
xor U398 (N_398,In_391,In_467);
nor U399 (N_399,In_293,In_484);
or U400 (N_400,In_154,In_57);
and U401 (N_401,In_220,In_451);
nor U402 (N_402,In_339,In_324);
nand U403 (N_403,In_257,In_496);
or U404 (N_404,In_139,In_30);
nor U405 (N_405,In_384,In_473);
or U406 (N_406,In_78,In_155);
and U407 (N_407,In_37,In_118);
nand U408 (N_408,In_265,In_484);
and U409 (N_409,In_149,In_197);
and U410 (N_410,In_51,In_225);
or U411 (N_411,In_122,In_146);
and U412 (N_412,In_57,In_410);
nand U413 (N_413,In_308,In_255);
or U414 (N_414,In_144,In_260);
nor U415 (N_415,In_298,In_491);
or U416 (N_416,In_301,In_15);
xnor U417 (N_417,In_475,In_422);
nand U418 (N_418,In_354,In_16);
nor U419 (N_419,In_151,In_164);
and U420 (N_420,In_340,In_3);
nand U421 (N_421,In_88,In_267);
nor U422 (N_422,In_356,In_400);
nor U423 (N_423,In_65,In_490);
and U424 (N_424,In_253,In_360);
nor U425 (N_425,In_240,In_422);
and U426 (N_426,In_192,In_7);
nor U427 (N_427,In_183,In_17);
and U428 (N_428,In_221,In_325);
or U429 (N_429,In_307,In_214);
nand U430 (N_430,In_68,In_309);
or U431 (N_431,In_91,In_462);
or U432 (N_432,In_19,In_217);
xor U433 (N_433,In_63,In_359);
xnor U434 (N_434,In_77,In_222);
and U435 (N_435,In_263,In_99);
nand U436 (N_436,In_59,In_17);
nand U437 (N_437,In_482,In_241);
nand U438 (N_438,In_366,In_438);
xnor U439 (N_439,In_14,In_23);
nor U440 (N_440,In_237,In_294);
or U441 (N_441,In_42,In_57);
nor U442 (N_442,In_192,In_65);
or U443 (N_443,In_61,In_289);
and U444 (N_444,In_410,In_151);
and U445 (N_445,In_222,In_150);
and U446 (N_446,In_210,In_78);
xnor U447 (N_447,In_134,In_478);
and U448 (N_448,In_408,In_82);
or U449 (N_449,In_308,In_387);
or U450 (N_450,In_135,In_279);
nand U451 (N_451,In_275,In_55);
nand U452 (N_452,In_92,In_65);
or U453 (N_453,In_283,In_395);
xnor U454 (N_454,In_233,In_111);
xor U455 (N_455,In_5,In_221);
nor U456 (N_456,In_240,In_110);
or U457 (N_457,In_354,In_275);
nand U458 (N_458,In_358,In_134);
xor U459 (N_459,In_401,In_166);
and U460 (N_460,In_97,In_123);
and U461 (N_461,In_469,In_342);
nand U462 (N_462,In_206,In_90);
nor U463 (N_463,In_197,In_442);
nand U464 (N_464,In_443,In_188);
nand U465 (N_465,In_255,In_465);
nor U466 (N_466,In_417,In_253);
nand U467 (N_467,In_108,In_12);
or U468 (N_468,In_489,In_24);
nand U469 (N_469,In_380,In_56);
xor U470 (N_470,In_61,In_75);
nor U471 (N_471,In_494,In_407);
or U472 (N_472,In_87,In_58);
or U473 (N_473,In_60,In_233);
or U474 (N_474,In_421,In_55);
nand U475 (N_475,In_267,In_203);
and U476 (N_476,In_327,In_472);
or U477 (N_477,In_246,In_92);
and U478 (N_478,In_105,In_301);
or U479 (N_479,In_21,In_469);
nor U480 (N_480,In_266,In_371);
xnor U481 (N_481,In_265,In_453);
and U482 (N_482,In_309,In_150);
xor U483 (N_483,In_369,In_281);
or U484 (N_484,In_109,In_92);
and U485 (N_485,In_125,In_374);
and U486 (N_486,In_366,In_132);
nor U487 (N_487,In_109,In_293);
and U488 (N_488,In_414,In_35);
nand U489 (N_489,In_364,In_182);
xor U490 (N_490,In_158,In_483);
or U491 (N_491,In_422,In_193);
nand U492 (N_492,In_316,In_311);
nand U493 (N_493,In_479,In_283);
or U494 (N_494,In_202,In_324);
and U495 (N_495,In_135,In_6);
or U496 (N_496,In_99,In_2);
nand U497 (N_497,In_485,In_78);
and U498 (N_498,In_327,In_382);
nor U499 (N_499,In_415,In_59);
nand U500 (N_500,In_288,In_496);
and U501 (N_501,In_387,In_460);
nor U502 (N_502,In_32,In_137);
or U503 (N_503,In_40,In_244);
or U504 (N_504,In_417,In_101);
nand U505 (N_505,In_305,In_195);
and U506 (N_506,In_78,In_393);
xnor U507 (N_507,In_206,In_47);
and U508 (N_508,In_306,In_117);
or U509 (N_509,In_62,In_194);
and U510 (N_510,In_207,In_97);
nor U511 (N_511,In_17,In_252);
and U512 (N_512,In_237,In_224);
or U513 (N_513,In_291,In_225);
and U514 (N_514,In_90,In_331);
or U515 (N_515,In_370,In_292);
nor U516 (N_516,In_456,In_425);
xnor U517 (N_517,In_433,In_38);
or U518 (N_518,In_428,In_94);
nand U519 (N_519,In_335,In_81);
or U520 (N_520,In_158,In_322);
and U521 (N_521,In_193,In_383);
nor U522 (N_522,In_361,In_296);
xor U523 (N_523,In_327,In_152);
nor U524 (N_524,In_302,In_338);
xor U525 (N_525,In_208,In_357);
and U526 (N_526,In_201,In_383);
xnor U527 (N_527,In_98,In_427);
xor U528 (N_528,In_454,In_330);
nor U529 (N_529,In_100,In_244);
nand U530 (N_530,In_418,In_422);
or U531 (N_531,In_300,In_432);
nand U532 (N_532,In_174,In_452);
nor U533 (N_533,In_168,In_103);
xnor U534 (N_534,In_496,In_203);
nand U535 (N_535,In_353,In_404);
xnor U536 (N_536,In_281,In_184);
xnor U537 (N_537,In_101,In_323);
or U538 (N_538,In_253,In_215);
nand U539 (N_539,In_169,In_32);
nand U540 (N_540,In_469,In_282);
nand U541 (N_541,In_309,In_230);
xnor U542 (N_542,In_418,In_263);
nor U543 (N_543,In_487,In_116);
or U544 (N_544,In_444,In_366);
and U545 (N_545,In_140,In_82);
nand U546 (N_546,In_450,In_195);
xor U547 (N_547,In_396,In_246);
and U548 (N_548,In_347,In_202);
and U549 (N_549,In_188,In_228);
and U550 (N_550,In_296,In_151);
nand U551 (N_551,In_127,In_237);
xor U552 (N_552,In_114,In_359);
or U553 (N_553,In_230,In_326);
nor U554 (N_554,In_229,In_142);
nand U555 (N_555,In_46,In_42);
nand U556 (N_556,In_482,In_8);
nor U557 (N_557,In_273,In_293);
and U558 (N_558,In_271,In_403);
and U559 (N_559,In_14,In_149);
or U560 (N_560,In_275,In_323);
or U561 (N_561,In_400,In_80);
and U562 (N_562,In_408,In_9);
or U563 (N_563,In_166,In_449);
nor U564 (N_564,In_45,In_230);
nand U565 (N_565,In_330,In_151);
nor U566 (N_566,In_103,In_498);
or U567 (N_567,In_419,In_306);
nor U568 (N_568,In_218,In_164);
and U569 (N_569,In_78,In_103);
nand U570 (N_570,In_310,In_427);
or U571 (N_571,In_448,In_16);
or U572 (N_572,In_463,In_44);
and U573 (N_573,In_238,In_67);
nor U574 (N_574,In_482,In_71);
nor U575 (N_575,In_139,In_307);
or U576 (N_576,In_411,In_374);
and U577 (N_577,In_67,In_213);
and U578 (N_578,In_228,In_57);
or U579 (N_579,In_180,In_49);
xnor U580 (N_580,In_266,In_230);
or U581 (N_581,In_58,In_464);
or U582 (N_582,In_83,In_375);
nand U583 (N_583,In_373,In_274);
and U584 (N_584,In_371,In_174);
xor U585 (N_585,In_34,In_481);
xor U586 (N_586,In_368,In_124);
xor U587 (N_587,In_239,In_41);
and U588 (N_588,In_353,In_299);
nand U589 (N_589,In_55,In_308);
or U590 (N_590,In_160,In_391);
nand U591 (N_591,In_400,In_18);
xor U592 (N_592,In_438,In_239);
nor U593 (N_593,In_269,In_302);
nand U594 (N_594,In_46,In_496);
nor U595 (N_595,In_65,In_352);
nor U596 (N_596,In_496,In_333);
or U597 (N_597,In_331,In_479);
nor U598 (N_598,In_278,In_173);
or U599 (N_599,In_414,In_256);
or U600 (N_600,In_396,In_314);
nand U601 (N_601,In_63,In_439);
and U602 (N_602,In_67,In_194);
or U603 (N_603,In_140,In_22);
nand U604 (N_604,In_204,In_173);
nor U605 (N_605,In_5,In_22);
and U606 (N_606,In_270,In_320);
nor U607 (N_607,In_149,In_30);
xor U608 (N_608,In_444,In_202);
or U609 (N_609,In_357,In_267);
nand U610 (N_610,In_152,In_80);
or U611 (N_611,In_128,In_467);
and U612 (N_612,In_268,In_336);
nand U613 (N_613,In_394,In_53);
nor U614 (N_614,In_382,In_499);
and U615 (N_615,In_395,In_372);
and U616 (N_616,In_178,In_120);
or U617 (N_617,In_234,In_250);
nor U618 (N_618,In_410,In_22);
xnor U619 (N_619,In_495,In_169);
nor U620 (N_620,In_325,In_378);
nor U621 (N_621,In_135,In_311);
nand U622 (N_622,In_160,In_87);
nand U623 (N_623,In_268,In_426);
nand U624 (N_624,In_291,In_413);
or U625 (N_625,In_344,In_421);
or U626 (N_626,In_84,In_489);
and U627 (N_627,In_156,In_78);
and U628 (N_628,In_335,In_177);
nand U629 (N_629,In_434,In_396);
and U630 (N_630,In_198,In_281);
or U631 (N_631,In_14,In_311);
xnor U632 (N_632,In_198,In_99);
xnor U633 (N_633,In_355,In_386);
and U634 (N_634,In_264,In_345);
and U635 (N_635,In_408,In_63);
xnor U636 (N_636,In_456,In_252);
or U637 (N_637,In_281,In_457);
xor U638 (N_638,In_62,In_457);
xnor U639 (N_639,In_472,In_317);
or U640 (N_640,In_431,In_130);
and U641 (N_641,In_209,In_435);
and U642 (N_642,In_217,In_449);
nor U643 (N_643,In_196,In_63);
or U644 (N_644,In_312,In_368);
nand U645 (N_645,In_206,In_240);
and U646 (N_646,In_176,In_204);
xor U647 (N_647,In_5,In_155);
and U648 (N_648,In_81,In_26);
and U649 (N_649,In_423,In_119);
nand U650 (N_650,In_292,In_188);
nand U651 (N_651,In_231,In_114);
nand U652 (N_652,In_238,In_379);
nor U653 (N_653,In_385,In_187);
xor U654 (N_654,In_394,In_356);
or U655 (N_655,In_476,In_7);
or U656 (N_656,In_159,In_41);
or U657 (N_657,In_217,In_327);
nand U658 (N_658,In_333,In_104);
or U659 (N_659,In_68,In_217);
nand U660 (N_660,In_57,In_489);
and U661 (N_661,In_293,In_262);
nor U662 (N_662,In_197,In_140);
and U663 (N_663,In_395,In_363);
xnor U664 (N_664,In_44,In_97);
or U665 (N_665,In_192,In_162);
nand U666 (N_666,In_70,In_181);
nor U667 (N_667,In_94,In_449);
nand U668 (N_668,In_211,In_448);
or U669 (N_669,In_472,In_366);
or U670 (N_670,In_103,In_410);
nor U671 (N_671,In_411,In_284);
and U672 (N_672,In_486,In_131);
xor U673 (N_673,In_80,In_350);
or U674 (N_674,In_277,In_1);
xor U675 (N_675,In_6,In_317);
xnor U676 (N_676,In_171,In_295);
nor U677 (N_677,In_483,In_225);
nand U678 (N_678,In_416,In_48);
or U679 (N_679,In_14,In_462);
xnor U680 (N_680,In_358,In_208);
xor U681 (N_681,In_288,In_404);
nand U682 (N_682,In_241,In_396);
and U683 (N_683,In_476,In_130);
xnor U684 (N_684,In_139,In_8);
nor U685 (N_685,In_20,In_443);
nand U686 (N_686,In_97,In_235);
and U687 (N_687,In_343,In_166);
or U688 (N_688,In_334,In_315);
nor U689 (N_689,In_457,In_353);
or U690 (N_690,In_223,In_22);
or U691 (N_691,In_313,In_352);
or U692 (N_692,In_491,In_215);
and U693 (N_693,In_104,In_222);
and U694 (N_694,In_115,In_491);
xor U695 (N_695,In_127,In_309);
or U696 (N_696,In_431,In_51);
nand U697 (N_697,In_49,In_374);
or U698 (N_698,In_487,In_215);
nand U699 (N_699,In_355,In_398);
or U700 (N_700,In_71,In_208);
nor U701 (N_701,In_395,In_397);
or U702 (N_702,In_425,In_375);
or U703 (N_703,In_306,In_471);
or U704 (N_704,In_334,In_111);
and U705 (N_705,In_336,In_450);
nor U706 (N_706,In_176,In_56);
or U707 (N_707,In_303,In_375);
xnor U708 (N_708,In_436,In_225);
or U709 (N_709,In_54,In_340);
xnor U710 (N_710,In_275,In_434);
or U711 (N_711,In_327,In_359);
nor U712 (N_712,In_356,In_436);
nand U713 (N_713,In_455,In_391);
and U714 (N_714,In_321,In_55);
nor U715 (N_715,In_481,In_315);
nor U716 (N_716,In_354,In_128);
and U717 (N_717,In_237,In_222);
and U718 (N_718,In_160,In_126);
or U719 (N_719,In_385,In_486);
or U720 (N_720,In_453,In_499);
or U721 (N_721,In_460,In_493);
or U722 (N_722,In_105,In_220);
or U723 (N_723,In_460,In_314);
xnor U724 (N_724,In_433,In_287);
nand U725 (N_725,In_474,In_212);
nand U726 (N_726,In_309,In_18);
xnor U727 (N_727,In_456,In_420);
or U728 (N_728,In_54,In_28);
nand U729 (N_729,In_165,In_264);
xor U730 (N_730,In_233,In_288);
nand U731 (N_731,In_396,In_162);
nand U732 (N_732,In_439,In_186);
and U733 (N_733,In_22,In_116);
or U734 (N_734,In_209,In_221);
and U735 (N_735,In_41,In_185);
and U736 (N_736,In_487,In_200);
and U737 (N_737,In_460,In_224);
or U738 (N_738,In_18,In_213);
or U739 (N_739,In_206,In_179);
nand U740 (N_740,In_402,In_436);
nor U741 (N_741,In_404,In_264);
and U742 (N_742,In_495,In_217);
nor U743 (N_743,In_233,In_354);
nor U744 (N_744,In_89,In_428);
xnor U745 (N_745,In_11,In_324);
nor U746 (N_746,In_340,In_440);
nand U747 (N_747,In_322,In_164);
nand U748 (N_748,In_235,In_137);
nand U749 (N_749,In_420,In_54);
nor U750 (N_750,N_96,N_70);
or U751 (N_751,N_283,N_166);
or U752 (N_752,N_130,N_374);
nand U753 (N_753,N_12,N_602);
and U754 (N_754,N_304,N_69);
or U755 (N_755,N_94,N_587);
xnor U756 (N_756,N_343,N_267);
xnor U757 (N_757,N_68,N_254);
nand U758 (N_758,N_487,N_352);
or U759 (N_759,N_97,N_102);
xor U760 (N_760,N_411,N_442);
or U761 (N_761,N_468,N_675);
nor U762 (N_762,N_523,N_500);
xor U763 (N_763,N_211,N_430);
nor U764 (N_764,N_435,N_537);
xnor U765 (N_765,N_46,N_335);
nand U766 (N_766,N_456,N_49);
nor U767 (N_767,N_93,N_167);
nor U768 (N_768,N_426,N_672);
xor U769 (N_769,N_638,N_106);
or U770 (N_770,N_698,N_649);
nor U771 (N_771,N_192,N_148);
or U772 (N_772,N_339,N_629);
nor U773 (N_773,N_382,N_364);
or U774 (N_774,N_577,N_735);
and U775 (N_775,N_729,N_481);
xor U776 (N_776,N_741,N_613);
and U777 (N_777,N_718,N_677);
nor U778 (N_778,N_184,N_666);
xor U779 (N_779,N_200,N_409);
nand U780 (N_780,N_471,N_306);
nand U781 (N_781,N_333,N_476);
and U782 (N_782,N_67,N_201);
and U783 (N_783,N_312,N_278);
xor U784 (N_784,N_433,N_535);
nor U785 (N_785,N_488,N_226);
and U786 (N_786,N_238,N_30);
and U787 (N_787,N_562,N_414);
nand U788 (N_788,N_141,N_363);
nor U789 (N_789,N_318,N_216);
and U790 (N_790,N_520,N_214);
and U791 (N_791,N_38,N_708);
nand U792 (N_792,N_154,N_176);
and U793 (N_793,N_747,N_135);
xnor U794 (N_794,N_743,N_149);
xnor U795 (N_795,N_654,N_270);
xnor U796 (N_796,N_659,N_27);
and U797 (N_797,N_177,N_76);
nand U798 (N_798,N_618,N_632);
or U799 (N_799,N_244,N_515);
nand U800 (N_800,N_115,N_645);
or U801 (N_801,N_35,N_459);
or U802 (N_802,N_316,N_350);
nor U803 (N_803,N_533,N_421);
nand U804 (N_804,N_534,N_548);
nor U805 (N_805,N_678,N_39);
nor U806 (N_806,N_574,N_277);
and U807 (N_807,N_248,N_10);
or U808 (N_808,N_703,N_336);
and U809 (N_809,N_549,N_16);
or U810 (N_810,N_85,N_358);
and U811 (N_811,N_0,N_495);
and U812 (N_812,N_297,N_644);
nor U813 (N_813,N_348,N_369);
nand U814 (N_814,N_731,N_87);
xor U815 (N_815,N_491,N_9);
nor U816 (N_816,N_32,N_212);
or U817 (N_817,N_132,N_519);
or U818 (N_818,N_607,N_506);
and U819 (N_819,N_258,N_671);
nand U820 (N_820,N_257,N_377);
or U821 (N_821,N_53,N_714);
xor U822 (N_822,N_376,N_158);
xnor U823 (N_823,N_494,N_448);
nand U824 (N_824,N_619,N_172);
xor U825 (N_825,N_676,N_609);
or U826 (N_826,N_472,N_56);
nand U827 (N_827,N_740,N_474);
xnor U828 (N_828,N_58,N_662);
xor U829 (N_829,N_379,N_206);
nand U830 (N_830,N_229,N_23);
xnor U831 (N_831,N_569,N_725);
and U832 (N_832,N_664,N_564);
nor U833 (N_833,N_496,N_44);
or U834 (N_834,N_284,N_193);
and U835 (N_835,N_357,N_502);
xor U836 (N_836,N_140,N_145);
nand U837 (N_837,N_556,N_134);
nor U838 (N_838,N_41,N_40);
xnor U839 (N_839,N_593,N_247);
or U840 (N_840,N_110,N_726);
or U841 (N_841,N_422,N_103);
and U842 (N_842,N_272,N_315);
or U843 (N_843,N_510,N_608);
nand U844 (N_844,N_237,N_117);
nor U845 (N_845,N_555,N_626);
xor U846 (N_846,N_688,N_401);
nor U847 (N_847,N_462,N_341);
nand U848 (N_848,N_340,N_525);
nand U849 (N_849,N_596,N_386);
and U850 (N_850,N_100,N_710);
xor U851 (N_851,N_518,N_540);
and U852 (N_852,N_157,N_326);
xnor U853 (N_853,N_14,N_504);
nor U854 (N_854,N_338,N_559);
or U855 (N_855,N_658,N_394);
and U856 (N_856,N_291,N_657);
or U857 (N_857,N_187,N_446);
and U858 (N_858,N_427,N_734);
or U859 (N_859,N_656,N_526);
or U860 (N_860,N_13,N_451);
and U861 (N_861,N_98,N_225);
nor U862 (N_862,N_543,N_436);
xnor U863 (N_863,N_160,N_245);
nor U864 (N_864,N_371,N_652);
xor U865 (N_865,N_573,N_689);
or U866 (N_866,N_567,N_20);
nand U867 (N_867,N_292,N_286);
nor U868 (N_868,N_57,N_242);
nor U869 (N_869,N_604,N_440);
or U870 (N_870,N_388,N_499);
xor U871 (N_871,N_281,N_293);
nor U872 (N_872,N_190,N_294);
and U873 (N_873,N_538,N_365);
nand U874 (N_874,N_584,N_367);
and U875 (N_875,N_717,N_213);
nor U876 (N_876,N_22,N_696);
or U877 (N_877,N_397,N_610);
and U878 (N_878,N_156,N_113);
nand U879 (N_879,N_17,N_547);
and U880 (N_880,N_591,N_362);
nand U881 (N_881,N_334,N_739);
xnor U882 (N_882,N_640,N_480);
xnor U883 (N_883,N_528,N_551);
xnor U884 (N_884,N_660,N_265);
and U885 (N_885,N_81,N_8);
xor U886 (N_886,N_282,N_133);
nor U887 (N_887,N_307,N_709);
or U888 (N_888,N_693,N_588);
and U889 (N_889,N_152,N_178);
or U890 (N_890,N_15,N_322);
nor U891 (N_891,N_477,N_123);
nor U892 (N_892,N_712,N_461);
and U893 (N_893,N_723,N_641);
nand U894 (N_894,N_438,N_399);
nor U895 (N_895,N_196,N_31);
or U896 (N_896,N_384,N_623);
nor U897 (N_897,N_637,N_131);
nor U898 (N_898,N_509,N_575);
xor U899 (N_899,N_1,N_233);
xnor U900 (N_900,N_264,N_410);
and U901 (N_901,N_697,N_92);
xor U902 (N_902,N_303,N_521);
nand U903 (N_903,N_742,N_612);
nand U904 (N_904,N_625,N_420);
nor U905 (N_905,N_601,N_375);
nor U906 (N_906,N_126,N_473);
or U907 (N_907,N_109,N_234);
and U908 (N_908,N_568,N_191);
and U909 (N_909,N_589,N_513);
xor U910 (N_910,N_501,N_655);
or U911 (N_911,N_627,N_615);
nand U912 (N_912,N_185,N_634);
and U913 (N_913,N_252,N_391);
xnor U914 (N_914,N_570,N_143);
or U915 (N_915,N_230,N_26);
nand U916 (N_916,N_670,N_597);
nand U917 (N_917,N_482,N_255);
xnor U918 (N_918,N_301,N_415);
and U919 (N_919,N_406,N_581);
xor U920 (N_920,N_360,N_579);
and U921 (N_921,N_279,N_479);
xnor U922 (N_922,N_505,N_249);
xnor U923 (N_923,N_635,N_289);
or U924 (N_924,N_144,N_458);
or U925 (N_925,N_628,N_546);
xor U926 (N_926,N_37,N_497);
xor U927 (N_927,N_542,N_319);
xor U928 (N_928,N_437,N_180);
nand U929 (N_929,N_86,N_631);
nor U930 (N_930,N_241,N_127);
and U931 (N_931,N_380,N_353);
xnor U932 (N_932,N_606,N_125);
and U933 (N_933,N_195,N_28);
or U934 (N_934,N_309,N_616);
nand U935 (N_935,N_310,N_327);
nand U936 (N_936,N_240,N_349);
nand U937 (N_937,N_124,N_392);
and U938 (N_938,N_220,N_209);
xnor U939 (N_939,N_412,N_259);
and U940 (N_940,N_605,N_266);
xnor U941 (N_941,N_105,N_686);
xor U942 (N_942,N_373,N_48);
or U943 (N_943,N_314,N_287);
nand U944 (N_944,N_311,N_585);
nor U945 (N_945,N_337,N_661);
nor U946 (N_946,N_189,N_73);
nor U947 (N_947,N_561,N_550);
or U948 (N_948,N_91,N_381);
xor U949 (N_949,N_64,N_78);
nand U950 (N_950,N_669,N_598);
nor U951 (N_951,N_51,N_208);
nor U952 (N_952,N_478,N_325);
and U953 (N_953,N_368,N_332);
nor U954 (N_954,N_151,N_417);
and U955 (N_955,N_305,N_429);
xnor U956 (N_956,N_407,N_595);
nand U957 (N_957,N_42,N_692);
and U958 (N_958,N_159,N_227);
or U959 (N_959,N_413,N_398);
or U960 (N_960,N_285,N_682);
nor U961 (N_961,N_256,N_733);
xor U962 (N_962,N_432,N_586);
and U963 (N_963,N_330,N_385);
nor U964 (N_964,N_687,N_24);
nor U965 (N_965,N_82,N_99);
nand U966 (N_966,N_396,N_663);
or U967 (N_967,N_11,N_83);
nor U968 (N_968,N_34,N_485);
nand U969 (N_969,N_490,N_280);
and U970 (N_970,N_36,N_727);
nor U971 (N_971,N_453,N_566);
or U972 (N_972,N_439,N_444);
nor U973 (N_973,N_592,N_45);
nand U974 (N_974,N_359,N_33);
and U975 (N_975,N_320,N_389);
or U976 (N_976,N_700,N_450);
xor U977 (N_977,N_557,N_236);
nor U978 (N_978,N_695,N_18);
and U979 (N_979,N_74,N_366);
nor U980 (N_980,N_25,N_275);
or U981 (N_981,N_683,N_434);
and U982 (N_982,N_646,N_679);
or U983 (N_983,N_475,N_745);
nor U984 (N_984,N_215,N_202);
and U985 (N_985,N_722,N_173);
or U986 (N_986,N_29,N_578);
nor U987 (N_987,N_65,N_531);
or U988 (N_988,N_617,N_492);
xnor U989 (N_989,N_716,N_383);
xnor U990 (N_990,N_217,N_445);
and U991 (N_991,N_467,N_527);
nand U992 (N_992,N_514,N_54);
and U993 (N_993,N_511,N_624);
nor U994 (N_994,N_268,N_308);
and U995 (N_995,N_137,N_715);
nand U996 (N_996,N_572,N_324);
or U997 (N_997,N_121,N_503);
nor U998 (N_998,N_580,N_464);
and U999 (N_999,N_738,N_271);
or U1000 (N_1000,N_522,N_104);
xnor U1001 (N_1001,N_146,N_650);
or U1002 (N_1002,N_6,N_404);
xnor U1003 (N_1003,N_620,N_243);
nand U1004 (N_1004,N_681,N_203);
and U1005 (N_1005,N_347,N_465);
and U1006 (N_1006,N_7,N_390);
nand U1007 (N_1007,N_205,N_724);
or U1008 (N_1008,N_730,N_290);
nand U1009 (N_1009,N_484,N_351);
xor U1010 (N_1010,N_680,N_119);
or U1011 (N_1011,N_667,N_261);
and U1012 (N_1012,N_395,N_582);
nand U1013 (N_1013,N_138,N_483);
nor U1014 (N_1014,N_108,N_199);
nor U1015 (N_1015,N_170,N_639);
nand U1016 (N_1016,N_684,N_43);
nand U1017 (N_1017,N_431,N_372);
nor U1018 (N_1018,N_4,N_246);
or U1019 (N_1019,N_155,N_447);
and U1020 (N_1020,N_346,N_685);
or U1021 (N_1021,N_594,N_746);
or U1022 (N_1022,N_508,N_232);
nand U1023 (N_1023,N_165,N_253);
and U1024 (N_1024,N_52,N_512);
and U1025 (N_1025,N_198,N_393);
and U1026 (N_1026,N_553,N_183);
and U1027 (N_1027,N_95,N_370);
and U1028 (N_1028,N_179,N_603);
and U1029 (N_1029,N_642,N_75);
nor U1030 (N_1030,N_558,N_418);
xnor U1031 (N_1031,N_288,N_674);
nor U1032 (N_1032,N_162,N_188);
xor U1033 (N_1033,N_345,N_600);
and U1034 (N_1034,N_3,N_651);
xor U1035 (N_1035,N_89,N_599);
nand U1036 (N_1036,N_405,N_354);
and U1037 (N_1037,N_194,N_295);
and U1038 (N_1038,N_673,N_171);
nand U1039 (N_1039,N_90,N_704);
or U1040 (N_1040,N_120,N_62);
nand U1041 (N_1041,N_736,N_463);
xnor U1042 (N_1042,N_222,N_705);
xnor U1043 (N_1043,N_636,N_560);
or U1044 (N_1044,N_5,N_219);
and U1045 (N_1045,N_300,N_460);
xor U1046 (N_1046,N_529,N_197);
and U1047 (N_1047,N_648,N_79);
nand U1048 (N_1048,N_169,N_223);
and U1049 (N_1049,N_224,N_59);
nand U1050 (N_1050,N_61,N_118);
xor U1051 (N_1051,N_150,N_139);
xor U1052 (N_1052,N_454,N_387);
or U1053 (N_1053,N_614,N_728);
xor U1054 (N_1054,N_400,N_690);
xnor U1055 (N_1055,N_441,N_653);
or U1056 (N_1056,N_565,N_302);
nor U1057 (N_1057,N_486,N_416);
nor U1058 (N_1058,N_299,N_507);
and U1059 (N_1059,N_331,N_50);
xor U1060 (N_1060,N_524,N_80);
or U1061 (N_1061,N_47,N_60);
xnor U1062 (N_1062,N_403,N_516);
nor U1063 (N_1063,N_111,N_147);
and U1064 (N_1064,N_563,N_164);
nand U1065 (N_1065,N_274,N_536);
or U1066 (N_1066,N_544,N_298);
nor U1067 (N_1067,N_101,N_107);
xor U1068 (N_1068,N_378,N_539);
nor U1069 (N_1069,N_263,N_88);
nand U1070 (N_1070,N_114,N_153);
or U1071 (N_1071,N_744,N_112);
nor U1072 (N_1072,N_665,N_699);
nor U1073 (N_1073,N_721,N_273);
nand U1074 (N_1074,N_469,N_77);
xnor U1075 (N_1075,N_342,N_424);
and U1076 (N_1076,N_711,N_129);
or U1077 (N_1077,N_719,N_276);
xor U1078 (N_1078,N_116,N_590);
and U1079 (N_1079,N_749,N_269);
or U1080 (N_1080,N_72,N_720);
xor U1081 (N_1081,N_706,N_251);
nand U1082 (N_1082,N_423,N_181);
xnor U1083 (N_1083,N_402,N_532);
nor U1084 (N_1084,N_713,N_571);
and U1085 (N_1085,N_122,N_493);
nand U1086 (N_1086,N_313,N_470);
xor U1087 (N_1087,N_262,N_701);
and U1088 (N_1088,N_541,N_218);
or U1089 (N_1089,N_329,N_321);
xor U1090 (N_1090,N_317,N_694);
xor U1091 (N_1091,N_239,N_552);
nand U1092 (N_1092,N_702,N_182);
xor U1093 (N_1093,N_66,N_296);
or U1094 (N_1094,N_530,N_161);
nand U1095 (N_1095,N_235,N_425);
or U1096 (N_1096,N_210,N_207);
or U1097 (N_1097,N_576,N_221);
and U1098 (N_1098,N_128,N_583);
xor U1099 (N_1099,N_621,N_63);
nor U1100 (N_1100,N_455,N_163);
or U1101 (N_1101,N_457,N_668);
and U1102 (N_1102,N_428,N_449);
nand U1103 (N_1103,N_231,N_84);
nand U1104 (N_1104,N_737,N_2);
nand U1105 (N_1105,N_323,N_71);
or U1106 (N_1106,N_344,N_452);
nor U1107 (N_1107,N_21,N_443);
nor U1108 (N_1108,N_691,N_748);
or U1109 (N_1109,N_328,N_633);
xor U1110 (N_1110,N_55,N_142);
xor U1111 (N_1111,N_498,N_545);
or U1112 (N_1112,N_168,N_408);
or U1113 (N_1113,N_517,N_136);
xor U1114 (N_1114,N_643,N_186);
nor U1115 (N_1115,N_622,N_228);
nor U1116 (N_1116,N_250,N_554);
and U1117 (N_1117,N_260,N_419);
nand U1118 (N_1118,N_356,N_174);
and U1119 (N_1119,N_630,N_732);
or U1120 (N_1120,N_611,N_19);
nor U1121 (N_1121,N_355,N_489);
and U1122 (N_1122,N_466,N_707);
and U1123 (N_1123,N_647,N_361);
or U1124 (N_1124,N_204,N_175);
nor U1125 (N_1125,N_577,N_596);
or U1126 (N_1126,N_529,N_155);
or U1127 (N_1127,N_665,N_331);
xnor U1128 (N_1128,N_144,N_496);
and U1129 (N_1129,N_230,N_314);
xnor U1130 (N_1130,N_714,N_12);
xor U1131 (N_1131,N_634,N_352);
xnor U1132 (N_1132,N_595,N_154);
and U1133 (N_1133,N_210,N_535);
nor U1134 (N_1134,N_265,N_392);
nor U1135 (N_1135,N_228,N_128);
nand U1136 (N_1136,N_183,N_640);
and U1137 (N_1137,N_488,N_432);
nand U1138 (N_1138,N_79,N_551);
or U1139 (N_1139,N_252,N_708);
nor U1140 (N_1140,N_12,N_272);
nand U1141 (N_1141,N_311,N_497);
xor U1142 (N_1142,N_158,N_315);
nand U1143 (N_1143,N_374,N_34);
xor U1144 (N_1144,N_389,N_111);
and U1145 (N_1145,N_185,N_461);
and U1146 (N_1146,N_511,N_680);
nand U1147 (N_1147,N_34,N_5);
xnor U1148 (N_1148,N_707,N_366);
nand U1149 (N_1149,N_144,N_113);
or U1150 (N_1150,N_546,N_59);
or U1151 (N_1151,N_310,N_16);
nor U1152 (N_1152,N_518,N_714);
nand U1153 (N_1153,N_520,N_465);
nand U1154 (N_1154,N_584,N_399);
nor U1155 (N_1155,N_324,N_695);
nor U1156 (N_1156,N_42,N_641);
nor U1157 (N_1157,N_380,N_566);
or U1158 (N_1158,N_413,N_403);
nand U1159 (N_1159,N_197,N_42);
nand U1160 (N_1160,N_63,N_589);
nand U1161 (N_1161,N_240,N_193);
and U1162 (N_1162,N_328,N_414);
and U1163 (N_1163,N_426,N_300);
and U1164 (N_1164,N_538,N_240);
and U1165 (N_1165,N_401,N_702);
nand U1166 (N_1166,N_475,N_386);
nand U1167 (N_1167,N_586,N_743);
xnor U1168 (N_1168,N_575,N_547);
xor U1169 (N_1169,N_287,N_631);
nor U1170 (N_1170,N_699,N_430);
or U1171 (N_1171,N_268,N_561);
and U1172 (N_1172,N_679,N_85);
or U1173 (N_1173,N_631,N_129);
nand U1174 (N_1174,N_587,N_360);
or U1175 (N_1175,N_400,N_572);
and U1176 (N_1176,N_208,N_254);
xor U1177 (N_1177,N_380,N_339);
or U1178 (N_1178,N_240,N_350);
nor U1179 (N_1179,N_157,N_365);
and U1180 (N_1180,N_618,N_697);
nor U1181 (N_1181,N_30,N_226);
and U1182 (N_1182,N_449,N_191);
nor U1183 (N_1183,N_8,N_121);
and U1184 (N_1184,N_519,N_421);
nand U1185 (N_1185,N_172,N_80);
or U1186 (N_1186,N_409,N_435);
nor U1187 (N_1187,N_722,N_638);
and U1188 (N_1188,N_567,N_55);
nor U1189 (N_1189,N_605,N_324);
or U1190 (N_1190,N_624,N_285);
or U1191 (N_1191,N_328,N_612);
nand U1192 (N_1192,N_204,N_206);
nand U1193 (N_1193,N_338,N_617);
xor U1194 (N_1194,N_539,N_429);
xor U1195 (N_1195,N_409,N_247);
nand U1196 (N_1196,N_526,N_727);
and U1197 (N_1197,N_123,N_284);
xor U1198 (N_1198,N_65,N_250);
or U1199 (N_1199,N_574,N_659);
or U1200 (N_1200,N_309,N_37);
or U1201 (N_1201,N_140,N_395);
or U1202 (N_1202,N_505,N_597);
and U1203 (N_1203,N_530,N_278);
nor U1204 (N_1204,N_469,N_562);
nand U1205 (N_1205,N_613,N_357);
nor U1206 (N_1206,N_684,N_118);
xnor U1207 (N_1207,N_493,N_296);
and U1208 (N_1208,N_257,N_734);
or U1209 (N_1209,N_594,N_348);
or U1210 (N_1210,N_658,N_401);
or U1211 (N_1211,N_434,N_110);
or U1212 (N_1212,N_307,N_342);
and U1213 (N_1213,N_368,N_20);
and U1214 (N_1214,N_625,N_335);
nor U1215 (N_1215,N_53,N_363);
or U1216 (N_1216,N_507,N_314);
or U1217 (N_1217,N_645,N_710);
xnor U1218 (N_1218,N_341,N_294);
and U1219 (N_1219,N_37,N_289);
nand U1220 (N_1220,N_659,N_388);
or U1221 (N_1221,N_297,N_175);
or U1222 (N_1222,N_319,N_161);
and U1223 (N_1223,N_116,N_595);
xor U1224 (N_1224,N_60,N_631);
or U1225 (N_1225,N_315,N_121);
and U1226 (N_1226,N_127,N_121);
nand U1227 (N_1227,N_247,N_236);
or U1228 (N_1228,N_125,N_600);
nand U1229 (N_1229,N_209,N_335);
and U1230 (N_1230,N_320,N_589);
nand U1231 (N_1231,N_545,N_427);
or U1232 (N_1232,N_28,N_607);
or U1233 (N_1233,N_650,N_407);
nand U1234 (N_1234,N_78,N_570);
and U1235 (N_1235,N_705,N_742);
nand U1236 (N_1236,N_212,N_622);
nor U1237 (N_1237,N_253,N_616);
or U1238 (N_1238,N_568,N_719);
nor U1239 (N_1239,N_205,N_221);
xor U1240 (N_1240,N_749,N_355);
and U1241 (N_1241,N_449,N_25);
or U1242 (N_1242,N_256,N_394);
xnor U1243 (N_1243,N_68,N_374);
nand U1244 (N_1244,N_577,N_632);
nand U1245 (N_1245,N_728,N_405);
and U1246 (N_1246,N_199,N_740);
nor U1247 (N_1247,N_524,N_459);
xor U1248 (N_1248,N_734,N_147);
nor U1249 (N_1249,N_17,N_73);
nor U1250 (N_1250,N_226,N_505);
nor U1251 (N_1251,N_376,N_437);
or U1252 (N_1252,N_488,N_520);
xnor U1253 (N_1253,N_439,N_635);
or U1254 (N_1254,N_506,N_348);
xnor U1255 (N_1255,N_529,N_18);
nand U1256 (N_1256,N_122,N_126);
nor U1257 (N_1257,N_406,N_592);
xnor U1258 (N_1258,N_79,N_105);
or U1259 (N_1259,N_398,N_556);
or U1260 (N_1260,N_248,N_418);
nand U1261 (N_1261,N_660,N_485);
and U1262 (N_1262,N_268,N_163);
nand U1263 (N_1263,N_667,N_373);
xor U1264 (N_1264,N_40,N_683);
nor U1265 (N_1265,N_90,N_245);
nor U1266 (N_1266,N_668,N_649);
or U1267 (N_1267,N_580,N_61);
nor U1268 (N_1268,N_694,N_501);
and U1269 (N_1269,N_560,N_716);
and U1270 (N_1270,N_268,N_673);
nor U1271 (N_1271,N_540,N_72);
or U1272 (N_1272,N_730,N_417);
nor U1273 (N_1273,N_746,N_459);
and U1274 (N_1274,N_2,N_435);
xnor U1275 (N_1275,N_303,N_212);
nand U1276 (N_1276,N_65,N_42);
nor U1277 (N_1277,N_166,N_68);
nand U1278 (N_1278,N_301,N_738);
nor U1279 (N_1279,N_134,N_701);
or U1280 (N_1280,N_268,N_650);
nand U1281 (N_1281,N_525,N_54);
xnor U1282 (N_1282,N_167,N_705);
nand U1283 (N_1283,N_454,N_734);
xnor U1284 (N_1284,N_167,N_478);
nand U1285 (N_1285,N_296,N_160);
nand U1286 (N_1286,N_379,N_90);
nor U1287 (N_1287,N_391,N_736);
and U1288 (N_1288,N_166,N_469);
nor U1289 (N_1289,N_371,N_643);
and U1290 (N_1290,N_454,N_359);
nand U1291 (N_1291,N_467,N_210);
xnor U1292 (N_1292,N_531,N_100);
or U1293 (N_1293,N_596,N_498);
nand U1294 (N_1294,N_519,N_495);
nor U1295 (N_1295,N_181,N_378);
xor U1296 (N_1296,N_66,N_733);
nand U1297 (N_1297,N_237,N_330);
and U1298 (N_1298,N_27,N_87);
nor U1299 (N_1299,N_227,N_466);
and U1300 (N_1300,N_243,N_444);
or U1301 (N_1301,N_321,N_562);
or U1302 (N_1302,N_623,N_579);
nand U1303 (N_1303,N_258,N_459);
xnor U1304 (N_1304,N_641,N_337);
and U1305 (N_1305,N_453,N_284);
or U1306 (N_1306,N_243,N_170);
nor U1307 (N_1307,N_160,N_107);
and U1308 (N_1308,N_344,N_209);
nor U1309 (N_1309,N_513,N_324);
and U1310 (N_1310,N_699,N_96);
and U1311 (N_1311,N_568,N_669);
or U1312 (N_1312,N_721,N_413);
and U1313 (N_1313,N_708,N_477);
xnor U1314 (N_1314,N_706,N_230);
or U1315 (N_1315,N_301,N_73);
nor U1316 (N_1316,N_389,N_78);
and U1317 (N_1317,N_439,N_655);
and U1318 (N_1318,N_90,N_741);
nor U1319 (N_1319,N_213,N_665);
nand U1320 (N_1320,N_610,N_79);
xnor U1321 (N_1321,N_573,N_52);
xnor U1322 (N_1322,N_308,N_76);
nand U1323 (N_1323,N_650,N_599);
and U1324 (N_1324,N_642,N_495);
nor U1325 (N_1325,N_371,N_669);
xnor U1326 (N_1326,N_263,N_704);
or U1327 (N_1327,N_583,N_351);
nand U1328 (N_1328,N_374,N_610);
nor U1329 (N_1329,N_725,N_564);
or U1330 (N_1330,N_710,N_536);
and U1331 (N_1331,N_582,N_587);
nand U1332 (N_1332,N_184,N_185);
xor U1333 (N_1333,N_606,N_179);
nor U1334 (N_1334,N_529,N_668);
or U1335 (N_1335,N_432,N_123);
or U1336 (N_1336,N_510,N_226);
nor U1337 (N_1337,N_414,N_80);
or U1338 (N_1338,N_82,N_89);
nor U1339 (N_1339,N_701,N_4);
nor U1340 (N_1340,N_347,N_263);
nand U1341 (N_1341,N_169,N_5);
nor U1342 (N_1342,N_416,N_519);
xor U1343 (N_1343,N_556,N_268);
nand U1344 (N_1344,N_261,N_503);
or U1345 (N_1345,N_496,N_36);
or U1346 (N_1346,N_740,N_482);
nand U1347 (N_1347,N_450,N_523);
and U1348 (N_1348,N_100,N_342);
nor U1349 (N_1349,N_531,N_734);
xor U1350 (N_1350,N_326,N_52);
nor U1351 (N_1351,N_286,N_502);
nand U1352 (N_1352,N_174,N_583);
xor U1353 (N_1353,N_505,N_272);
nor U1354 (N_1354,N_738,N_287);
xnor U1355 (N_1355,N_23,N_488);
or U1356 (N_1356,N_721,N_287);
or U1357 (N_1357,N_396,N_181);
nand U1358 (N_1358,N_360,N_20);
xor U1359 (N_1359,N_250,N_149);
xor U1360 (N_1360,N_719,N_216);
or U1361 (N_1361,N_257,N_22);
or U1362 (N_1362,N_132,N_409);
nand U1363 (N_1363,N_124,N_317);
or U1364 (N_1364,N_725,N_165);
nor U1365 (N_1365,N_391,N_128);
nand U1366 (N_1366,N_105,N_451);
nor U1367 (N_1367,N_314,N_709);
and U1368 (N_1368,N_173,N_24);
xor U1369 (N_1369,N_277,N_206);
xnor U1370 (N_1370,N_88,N_562);
xor U1371 (N_1371,N_427,N_362);
or U1372 (N_1372,N_309,N_220);
and U1373 (N_1373,N_362,N_443);
nand U1374 (N_1374,N_89,N_746);
or U1375 (N_1375,N_364,N_490);
or U1376 (N_1376,N_460,N_211);
xnor U1377 (N_1377,N_13,N_115);
nand U1378 (N_1378,N_285,N_47);
xor U1379 (N_1379,N_256,N_554);
and U1380 (N_1380,N_180,N_441);
or U1381 (N_1381,N_234,N_153);
and U1382 (N_1382,N_208,N_348);
nor U1383 (N_1383,N_124,N_444);
xor U1384 (N_1384,N_666,N_373);
nor U1385 (N_1385,N_290,N_686);
or U1386 (N_1386,N_126,N_715);
nor U1387 (N_1387,N_92,N_252);
xor U1388 (N_1388,N_92,N_732);
nor U1389 (N_1389,N_565,N_410);
nand U1390 (N_1390,N_555,N_256);
or U1391 (N_1391,N_576,N_716);
and U1392 (N_1392,N_734,N_536);
nand U1393 (N_1393,N_47,N_327);
and U1394 (N_1394,N_496,N_156);
nor U1395 (N_1395,N_276,N_690);
or U1396 (N_1396,N_631,N_109);
nand U1397 (N_1397,N_519,N_262);
and U1398 (N_1398,N_653,N_197);
nand U1399 (N_1399,N_279,N_266);
and U1400 (N_1400,N_140,N_229);
and U1401 (N_1401,N_121,N_271);
and U1402 (N_1402,N_170,N_78);
or U1403 (N_1403,N_242,N_391);
nand U1404 (N_1404,N_440,N_99);
nor U1405 (N_1405,N_23,N_704);
nor U1406 (N_1406,N_553,N_122);
and U1407 (N_1407,N_29,N_509);
xnor U1408 (N_1408,N_445,N_224);
nor U1409 (N_1409,N_484,N_274);
nor U1410 (N_1410,N_195,N_232);
xor U1411 (N_1411,N_292,N_172);
or U1412 (N_1412,N_188,N_479);
nor U1413 (N_1413,N_548,N_268);
nor U1414 (N_1414,N_609,N_160);
nand U1415 (N_1415,N_499,N_126);
nor U1416 (N_1416,N_717,N_611);
nand U1417 (N_1417,N_588,N_572);
and U1418 (N_1418,N_289,N_675);
and U1419 (N_1419,N_262,N_366);
or U1420 (N_1420,N_401,N_596);
nor U1421 (N_1421,N_507,N_578);
nand U1422 (N_1422,N_18,N_174);
and U1423 (N_1423,N_145,N_2);
nor U1424 (N_1424,N_602,N_136);
and U1425 (N_1425,N_610,N_681);
and U1426 (N_1426,N_59,N_94);
or U1427 (N_1427,N_596,N_176);
xnor U1428 (N_1428,N_14,N_710);
and U1429 (N_1429,N_242,N_362);
nor U1430 (N_1430,N_345,N_399);
nor U1431 (N_1431,N_748,N_728);
nor U1432 (N_1432,N_207,N_688);
nand U1433 (N_1433,N_604,N_445);
nor U1434 (N_1434,N_321,N_190);
or U1435 (N_1435,N_514,N_272);
and U1436 (N_1436,N_542,N_13);
nor U1437 (N_1437,N_375,N_114);
or U1438 (N_1438,N_137,N_432);
nand U1439 (N_1439,N_646,N_698);
xor U1440 (N_1440,N_486,N_744);
nand U1441 (N_1441,N_539,N_506);
and U1442 (N_1442,N_367,N_156);
nand U1443 (N_1443,N_51,N_243);
nor U1444 (N_1444,N_319,N_491);
nand U1445 (N_1445,N_237,N_323);
nand U1446 (N_1446,N_489,N_45);
nand U1447 (N_1447,N_58,N_668);
nand U1448 (N_1448,N_382,N_537);
nor U1449 (N_1449,N_87,N_348);
xor U1450 (N_1450,N_664,N_669);
xor U1451 (N_1451,N_116,N_516);
or U1452 (N_1452,N_579,N_739);
or U1453 (N_1453,N_476,N_221);
or U1454 (N_1454,N_232,N_688);
or U1455 (N_1455,N_542,N_42);
or U1456 (N_1456,N_703,N_720);
and U1457 (N_1457,N_141,N_216);
or U1458 (N_1458,N_223,N_573);
nand U1459 (N_1459,N_34,N_177);
or U1460 (N_1460,N_684,N_620);
xnor U1461 (N_1461,N_463,N_458);
or U1462 (N_1462,N_666,N_536);
nand U1463 (N_1463,N_38,N_696);
nand U1464 (N_1464,N_84,N_329);
and U1465 (N_1465,N_666,N_258);
and U1466 (N_1466,N_460,N_278);
nand U1467 (N_1467,N_421,N_247);
and U1468 (N_1468,N_102,N_303);
nor U1469 (N_1469,N_524,N_748);
nand U1470 (N_1470,N_35,N_235);
and U1471 (N_1471,N_672,N_686);
xor U1472 (N_1472,N_66,N_93);
nand U1473 (N_1473,N_428,N_232);
nand U1474 (N_1474,N_418,N_678);
nor U1475 (N_1475,N_517,N_230);
and U1476 (N_1476,N_274,N_687);
nand U1477 (N_1477,N_749,N_306);
or U1478 (N_1478,N_720,N_467);
and U1479 (N_1479,N_622,N_564);
and U1480 (N_1480,N_218,N_327);
nand U1481 (N_1481,N_156,N_120);
nor U1482 (N_1482,N_18,N_386);
or U1483 (N_1483,N_62,N_180);
or U1484 (N_1484,N_607,N_187);
or U1485 (N_1485,N_355,N_392);
or U1486 (N_1486,N_431,N_741);
and U1487 (N_1487,N_584,N_53);
nor U1488 (N_1488,N_137,N_494);
nor U1489 (N_1489,N_465,N_648);
and U1490 (N_1490,N_141,N_292);
xnor U1491 (N_1491,N_465,N_197);
or U1492 (N_1492,N_310,N_186);
nand U1493 (N_1493,N_198,N_558);
xor U1494 (N_1494,N_716,N_55);
and U1495 (N_1495,N_529,N_713);
xor U1496 (N_1496,N_318,N_494);
and U1497 (N_1497,N_77,N_231);
xor U1498 (N_1498,N_299,N_663);
or U1499 (N_1499,N_545,N_422);
nand U1500 (N_1500,N_965,N_1165);
nand U1501 (N_1501,N_1357,N_1106);
or U1502 (N_1502,N_1051,N_809);
xnor U1503 (N_1503,N_991,N_911);
or U1504 (N_1504,N_1241,N_917);
or U1505 (N_1505,N_1240,N_1231);
xnor U1506 (N_1506,N_823,N_1353);
xnor U1507 (N_1507,N_1496,N_1274);
and U1508 (N_1508,N_768,N_1430);
and U1509 (N_1509,N_1145,N_1325);
nor U1510 (N_1510,N_1100,N_866);
nand U1511 (N_1511,N_1320,N_895);
or U1512 (N_1512,N_1227,N_1276);
and U1513 (N_1513,N_821,N_791);
nand U1514 (N_1514,N_916,N_1432);
xor U1515 (N_1515,N_832,N_1177);
nand U1516 (N_1516,N_936,N_779);
or U1517 (N_1517,N_1483,N_1207);
and U1518 (N_1518,N_1200,N_1449);
xnor U1519 (N_1519,N_928,N_1042);
xnor U1520 (N_1520,N_1013,N_776);
xor U1521 (N_1521,N_1370,N_926);
xor U1522 (N_1522,N_827,N_1262);
nand U1523 (N_1523,N_953,N_1067);
nor U1524 (N_1524,N_1162,N_1193);
xor U1525 (N_1525,N_1005,N_1028);
nor U1526 (N_1526,N_1210,N_781);
nor U1527 (N_1527,N_1123,N_909);
nor U1528 (N_1528,N_1480,N_1078);
nor U1529 (N_1529,N_1349,N_1406);
and U1530 (N_1530,N_763,N_908);
nor U1531 (N_1531,N_1378,N_1478);
nand U1532 (N_1532,N_1056,N_1220);
xor U1533 (N_1533,N_1255,N_1286);
and U1534 (N_1534,N_1239,N_1499);
nor U1535 (N_1535,N_945,N_881);
or U1536 (N_1536,N_811,N_1159);
nand U1537 (N_1537,N_1148,N_1367);
or U1538 (N_1538,N_1141,N_854);
and U1539 (N_1539,N_1484,N_1054);
or U1540 (N_1540,N_1172,N_830);
nor U1541 (N_1541,N_1047,N_1436);
nor U1542 (N_1542,N_1246,N_1282);
or U1543 (N_1543,N_884,N_990);
xnor U1544 (N_1544,N_1356,N_1365);
and U1545 (N_1545,N_1431,N_886);
nor U1546 (N_1546,N_1423,N_943);
or U1547 (N_1547,N_980,N_1296);
or U1548 (N_1548,N_1104,N_1040);
or U1549 (N_1549,N_864,N_793);
xnor U1550 (N_1550,N_970,N_865);
and U1551 (N_1551,N_921,N_1069);
nor U1552 (N_1552,N_1105,N_1301);
xnor U1553 (N_1553,N_1397,N_1329);
and U1554 (N_1554,N_1198,N_1342);
or U1555 (N_1555,N_923,N_1212);
and U1556 (N_1556,N_1147,N_798);
or U1557 (N_1557,N_1023,N_1394);
nand U1558 (N_1558,N_1179,N_974);
nor U1559 (N_1559,N_1487,N_1073);
nor U1560 (N_1560,N_1155,N_903);
and U1561 (N_1561,N_1359,N_1188);
nand U1562 (N_1562,N_1292,N_888);
or U1563 (N_1563,N_1345,N_1171);
nand U1564 (N_1564,N_952,N_996);
nor U1565 (N_1565,N_1091,N_887);
nand U1566 (N_1566,N_1303,N_754);
xnor U1567 (N_1567,N_1464,N_1333);
xnor U1568 (N_1568,N_1376,N_858);
or U1569 (N_1569,N_1335,N_859);
and U1570 (N_1570,N_1295,N_1205);
or U1571 (N_1571,N_1379,N_880);
xor U1572 (N_1572,N_848,N_1383);
or U1573 (N_1573,N_1445,N_1229);
xnor U1574 (N_1574,N_876,N_1347);
and U1575 (N_1575,N_764,N_964);
and U1576 (N_1576,N_1362,N_870);
or U1577 (N_1577,N_961,N_1124);
xnor U1578 (N_1578,N_1390,N_1313);
nor U1579 (N_1579,N_988,N_1021);
nor U1580 (N_1580,N_1052,N_1242);
nand U1581 (N_1581,N_1457,N_1417);
and U1582 (N_1582,N_1369,N_1076);
nor U1583 (N_1583,N_1354,N_1451);
or U1584 (N_1584,N_1194,N_892);
nor U1585 (N_1585,N_820,N_983);
nand U1586 (N_1586,N_987,N_1455);
and U1587 (N_1587,N_808,N_800);
nand U1588 (N_1588,N_1377,N_963);
xor U1589 (N_1589,N_1217,N_968);
or U1590 (N_1590,N_939,N_1253);
and U1591 (N_1591,N_792,N_756);
nand U1592 (N_1592,N_1248,N_1036);
or U1593 (N_1593,N_1245,N_1143);
nor U1594 (N_1594,N_824,N_816);
and U1595 (N_1595,N_753,N_1048);
nand U1596 (N_1596,N_1173,N_1183);
nor U1597 (N_1597,N_1465,N_1190);
nor U1598 (N_1598,N_1355,N_769);
or U1599 (N_1599,N_1453,N_1053);
xnor U1600 (N_1600,N_1031,N_1132);
or U1601 (N_1601,N_878,N_841);
xnor U1602 (N_1602,N_1226,N_818);
and U1603 (N_1603,N_804,N_1402);
nand U1604 (N_1604,N_861,N_1469);
nor U1605 (N_1605,N_1090,N_1059);
xnor U1606 (N_1606,N_998,N_1395);
xor U1607 (N_1607,N_1189,N_1346);
and U1608 (N_1608,N_1434,N_1482);
xnor U1609 (N_1609,N_977,N_762);
nand U1610 (N_1610,N_1294,N_1452);
nor U1611 (N_1611,N_761,N_1348);
and U1612 (N_1612,N_1087,N_1267);
xor U1613 (N_1613,N_1291,N_1236);
xnor U1614 (N_1614,N_1187,N_941);
nand U1615 (N_1615,N_1486,N_1114);
xnor U1616 (N_1616,N_1283,N_1458);
nor U1617 (N_1617,N_1178,N_1219);
or U1618 (N_1618,N_976,N_839);
nor U1619 (N_1619,N_1381,N_1304);
or U1620 (N_1620,N_1293,N_867);
xor U1621 (N_1621,N_1409,N_959);
or U1622 (N_1622,N_1166,N_1203);
nor U1623 (N_1623,N_1020,N_1235);
nand U1624 (N_1624,N_1039,N_956);
nand U1625 (N_1625,N_1401,N_1014);
xor U1626 (N_1626,N_1099,N_1002);
xor U1627 (N_1627,N_958,N_978);
nand U1628 (N_1628,N_1270,N_1080);
or U1629 (N_1629,N_1061,N_1358);
or U1630 (N_1630,N_847,N_940);
nor U1631 (N_1631,N_1222,N_1199);
or U1632 (N_1632,N_1032,N_1427);
or U1633 (N_1633,N_1153,N_1079);
and U1634 (N_1634,N_1462,N_1459);
and U1635 (N_1635,N_900,N_1285);
nor U1636 (N_1636,N_984,N_1387);
xor U1637 (N_1637,N_765,N_1479);
xor U1638 (N_1638,N_894,N_948);
nand U1639 (N_1639,N_760,N_1133);
nand U1640 (N_1640,N_1107,N_1230);
nor U1641 (N_1641,N_1368,N_1201);
nor U1642 (N_1642,N_1338,N_1388);
xnor U1643 (N_1643,N_1111,N_1044);
nand U1644 (N_1644,N_846,N_999);
xor U1645 (N_1645,N_1029,N_1117);
and U1646 (N_1646,N_849,N_1339);
nand U1647 (N_1647,N_1384,N_1441);
nor U1648 (N_1648,N_1485,N_1223);
and U1649 (N_1649,N_1081,N_1043);
xor U1650 (N_1650,N_1298,N_992);
nand U1651 (N_1651,N_790,N_1151);
nand U1652 (N_1652,N_1128,N_1426);
nand U1653 (N_1653,N_1121,N_969);
and U1654 (N_1654,N_1094,N_962);
or U1655 (N_1655,N_1112,N_1138);
xnor U1656 (N_1656,N_954,N_1278);
or U1657 (N_1657,N_1149,N_1077);
nor U1658 (N_1658,N_1154,N_1326);
nor U1659 (N_1659,N_1498,N_1259);
and U1660 (N_1660,N_1167,N_1448);
or U1661 (N_1661,N_1308,N_1422);
and U1662 (N_1662,N_942,N_799);
nand U1663 (N_1663,N_913,N_1279);
or U1664 (N_1664,N_1256,N_1247);
and U1665 (N_1665,N_1157,N_794);
xor U1666 (N_1666,N_1122,N_1273);
or U1667 (N_1667,N_1468,N_1109);
xor U1668 (N_1668,N_929,N_1225);
nand U1669 (N_1669,N_1103,N_759);
and U1670 (N_1670,N_828,N_872);
xnor U1671 (N_1671,N_922,N_1476);
nand U1672 (N_1672,N_937,N_1251);
and U1673 (N_1673,N_1450,N_933);
and U1674 (N_1674,N_834,N_1470);
or U1675 (N_1675,N_835,N_844);
and U1676 (N_1676,N_782,N_1475);
and U1677 (N_1677,N_1265,N_863);
nor U1678 (N_1678,N_1228,N_893);
xor U1679 (N_1679,N_1209,N_1182);
or U1680 (N_1680,N_1249,N_1428);
nand U1681 (N_1681,N_1134,N_1063);
nand U1682 (N_1682,N_1454,N_1300);
nand U1683 (N_1683,N_994,N_1137);
nor U1684 (N_1684,N_1116,N_1393);
xnor U1685 (N_1685,N_1309,N_853);
or U1686 (N_1686,N_1161,N_1481);
or U1687 (N_1687,N_907,N_1421);
nor U1688 (N_1688,N_869,N_1102);
nand U1689 (N_1689,N_1062,N_1386);
or U1690 (N_1690,N_1016,N_1361);
or U1691 (N_1691,N_1410,N_788);
nor U1692 (N_1692,N_757,N_1131);
xnor U1693 (N_1693,N_1181,N_957);
nand U1694 (N_1694,N_1425,N_1082);
or U1695 (N_1695,N_1204,N_924);
and U1696 (N_1696,N_883,N_1363);
and U1697 (N_1697,N_979,N_1415);
or U1698 (N_1698,N_1068,N_927);
or U1699 (N_1699,N_833,N_1311);
or U1700 (N_1700,N_751,N_1408);
nand U1701 (N_1701,N_783,N_789);
nor U1702 (N_1702,N_1420,N_1083);
xnor U1703 (N_1703,N_877,N_918);
and U1704 (N_1704,N_1086,N_1389);
or U1705 (N_1705,N_1331,N_915);
nand U1706 (N_1706,N_1218,N_1146);
xnor U1707 (N_1707,N_771,N_1022);
nand U1708 (N_1708,N_882,N_1319);
nor U1709 (N_1709,N_1035,N_826);
or U1710 (N_1710,N_1164,N_1139);
nand U1711 (N_1711,N_1034,N_1493);
or U1712 (N_1712,N_871,N_801);
nand U1713 (N_1713,N_1208,N_935);
nor U1714 (N_1714,N_777,N_1049);
nand U1715 (N_1715,N_1396,N_1158);
nand U1716 (N_1716,N_806,N_857);
nor U1717 (N_1717,N_1385,N_1297);
or U1718 (N_1718,N_1174,N_752);
and U1719 (N_1719,N_1327,N_906);
and U1720 (N_1720,N_812,N_1089);
xnor U1721 (N_1721,N_1092,N_1497);
or U1722 (N_1722,N_1156,N_1372);
nor U1723 (N_1723,N_1371,N_1085);
nor U1724 (N_1724,N_896,N_1290);
nand U1725 (N_1725,N_1144,N_920);
xnor U1726 (N_1726,N_879,N_1010);
xnor U1727 (N_1727,N_1008,N_1012);
nor U1728 (N_1728,N_885,N_919);
xor U1729 (N_1729,N_995,N_1373);
xor U1730 (N_1730,N_778,N_890);
xor U1731 (N_1731,N_1224,N_1135);
and U1732 (N_1732,N_1072,N_1351);
nor U1733 (N_1733,N_910,N_1471);
xnor U1734 (N_1734,N_1271,N_1018);
xor U1735 (N_1735,N_1433,N_891);
or U1736 (N_1736,N_1214,N_815);
xor U1737 (N_1737,N_1472,N_1163);
nand U1738 (N_1738,N_1250,N_1337);
xnor U1739 (N_1739,N_797,N_1490);
or U1740 (N_1740,N_949,N_1244);
nor U1741 (N_1741,N_850,N_971);
xor U1742 (N_1742,N_1302,N_1266);
or U1743 (N_1743,N_780,N_1009);
and U1744 (N_1744,N_1243,N_1318);
or U1745 (N_1745,N_1095,N_1330);
nor U1746 (N_1746,N_1088,N_932);
or U1747 (N_1747,N_972,N_993);
nor U1748 (N_1748,N_901,N_989);
xnor U1749 (N_1749,N_1119,N_1312);
nor U1750 (N_1750,N_1324,N_997);
nor U1751 (N_1751,N_1041,N_755);
or U1752 (N_1752,N_1096,N_1398);
and U1753 (N_1753,N_1093,N_851);
xnor U1754 (N_1754,N_1057,N_1074);
and U1755 (N_1755,N_1261,N_1206);
nand U1756 (N_1756,N_1411,N_986);
or U1757 (N_1757,N_1257,N_1101);
xnor U1758 (N_1758,N_1180,N_862);
and U1759 (N_1759,N_1211,N_1024);
or U1760 (N_1760,N_1026,N_758);
nor U1761 (N_1761,N_1474,N_981);
nand U1762 (N_1762,N_1050,N_1442);
nor U1763 (N_1763,N_1045,N_1011);
nand U1764 (N_1764,N_1403,N_944);
nand U1765 (N_1765,N_1467,N_843);
or U1766 (N_1766,N_1352,N_931);
or U1767 (N_1767,N_1127,N_852);
or U1768 (N_1768,N_860,N_1323);
nand U1769 (N_1769,N_1003,N_1118);
nand U1770 (N_1770,N_1280,N_772);
nand U1771 (N_1771,N_1447,N_975);
and U1772 (N_1772,N_982,N_985);
xor U1773 (N_1773,N_813,N_855);
xor U1774 (N_1774,N_1380,N_966);
and U1775 (N_1775,N_1007,N_1494);
nor U1776 (N_1776,N_1491,N_899);
and U1777 (N_1777,N_1065,N_951);
or U1778 (N_1778,N_1186,N_1391);
and U1779 (N_1779,N_773,N_873);
and U1780 (N_1780,N_1382,N_1364);
nand U1781 (N_1781,N_1185,N_1192);
nand U1782 (N_1782,N_1168,N_822);
xor U1783 (N_1783,N_1060,N_1440);
and U1784 (N_1784,N_1120,N_947);
xor U1785 (N_1785,N_842,N_1438);
nand U1786 (N_1786,N_1066,N_1492);
and U1787 (N_1787,N_1281,N_805);
nand U1788 (N_1788,N_889,N_1321);
and U1789 (N_1789,N_1305,N_1314);
xnor U1790 (N_1790,N_1460,N_829);
xnor U1791 (N_1791,N_1176,N_930);
or U1792 (N_1792,N_898,N_1289);
or U1793 (N_1793,N_1332,N_1071);
and U1794 (N_1794,N_1275,N_1416);
and U1795 (N_1795,N_1152,N_1030);
xor U1796 (N_1796,N_1341,N_1374);
nor U1797 (N_1797,N_803,N_1268);
xnor U1798 (N_1798,N_912,N_1412);
or U1799 (N_1799,N_814,N_1269);
nand U1800 (N_1800,N_1058,N_1202);
nand U1801 (N_1801,N_1400,N_1025);
and U1802 (N_1802,N_1375,N_1263);
xor U1803 (N_1803,N_868,N_1419);
or U1804 (N_1804,N_1418,N_1473);
and U1805 (N_1805,N_1328,N_1310);
or U1806 (N_1806,N_1150,N_897);
and U1807 (N_1807,N_1288,N_825);
nand U1808 (N_1808,N_1126,N_1136);
nor U1809 (N_1809,N_1344,N_836);
nor U1810 (N_1810,N_1264,N_1287);
nand U1811 (N_1811,N_786,N_1019);
nand U1812 (N_1812,N_1437,N_946);
nand U1813 (N_1813,N_1098,N_1140);
xnor U1814 (N_1814,N_1461,N_1366);
or U1815 (N_1815,N_904,N_1360);
nand U1816 (N_1816,N_1260,N_831);
xor U1817 (N_1817,N_1169,N_1108);
nor U1818 (N_1818,N_1315,N_1252);
xor U1819 (N_1819,N_1350,N_1489);
nand U1820 (N_1820,N_810,N_1413);
nand U1821 (N_1821,N_1238,N_1336);
and U1822 (N_1822,N_1097,N_1277);
nor U1823 (N_1823,N_1055,N_770);
or U1824 (N_1824,N_1110,N_1392);
nor U1825 (N_1825,N_1463,N_1429);
and U1826 (N_1826,N_925,N_874);
xnor U1827 (N_1827,N_856,N_1254);
nor U1828 (N_1828,N_1197,N_1477);
and U1829 (N_1829,N_905,N_1006);
nor U1830 (N_1830,N_1444,N_967);
or U1831 (N_1831,N_950,N_1284);
or U1832 (N_1832,N_1234,N_902);
or U1833 (N_1833,N_774,N_1191);
xor U1834 (N_1834,N_1084,N_807);
or U1835 (N_1835,N_766,N_1233);
xnor U1836 (N_1836,N_1443,N_1215);
xnor U1837 (N_1837,N_1466,N_1258);
xor U1838 (N_1838,N_1125,N_1272);
and U1839 (N_1839,N_1414,N_1221);
nand U1840 (N_1840,N_1495,N_1456);
nor U1841 (N_1841,N_1130,N_1424);
and U1842 (N_1842,N_955,N_1307);
or U1843 (N_1843,N_1237,N_973);
nand U1844 (N_1844,N_819,N_1405);
or U1845 (N_1845,N_796,N_1160);
nand U1846 (N_1846,N_1195,N_1216);
and U1847 (N_1847,N_1115,N_787);
nand U1848 (N_1848,N_1046,N_784);
nor U1849 (N_1849,N_775,N_837);
xnor U1850 (N_1850,N_1075,N_767);
xor U1851 (N_1851,N_1000,N_795);
nand U1852 (N_1852,N_960,N_1064);
nor U1853 (N_1853,N_1015,N_938);
nand U1854 (N_1854,N_1033,N_750);
or U1855 (N_1855,N_1001,N_1439);
or U1856 (N_1856,N_1340,N_1038);
xnor U1857 (N_1857,N_1299,N_1170);
xnor U1858 (N_1858,N_1343,N_1196);
or U1859 (N_1859,N_1317,N_1037);
xor U1860 (N_1860,N_845,N_840);
nor U1861 (N_1861,N_1017,N_1232);
nor U1862 (N_1862,N_1184,N_1175);
and U1863 (N_1863,N_1435,N_1407);
xor U1864 (N_1864,N_1306,N_838);
and U1865 (N_1865,N_934,N_1142);
or U1866 (N_1866,N_1316,N_1322);
xnor U1867 (N_1867,N_1404,N_1070);
and U1868 (N_1868,N_1399,N_1446);
and U1869 (N_1869,N_914,N_785);
or U1870 (N_1870,N_1113,N_1334);
nor U1871 (N_1871,N_802,N_875);
nand U1872 (N_1872,N_817,N_1488);
xor U1873 (N_1873,N_1129,N_1004);
nor U1874 (N_1874,N_1027,N_1213);
or U1875 (N_1875,N_1339,N_936);
nand U1876 (N_1876,N_1121,N_1430);
or U1877 (N_1877,N_894,N_953);
or U1878 (N_1878,N_1113,N_1205);
xnor U1879 (N_1879,N_1438,N_1112);
nor U1880 (N_1880,N_1462,N_1048);
xor U1881 (N_1881,N_818,N_1012);
or U1882 (N_1882,N_1409,N_876);
and U1883 (N_1883,N_1094,N_1365);
and U1884 (N_1884,N_756,N_918);
and U1885 (N_1885,N_1021,N_921);
xor U1886 (N_1886,N_1289,N_919);
nand U1887 (N_1887,N_857,N_771);
or U1888 (N_1888,N_1268,N_998);
nand U1889 (N_1889,N_1156,N_1149);
nand U1890 (N_1890,N_1396,N_786);
or U1891 (N_1891,N_1111,N_782);
or U1892 (N_1892,N_1279,N_822);
xnor U1893 (N_1893,N_1261,N_854);
nor U1894 (N_1894,N_1078,N_770);
and U1895 (N_1895,N_963,N_812);
nor U1896 (N_1896,N_1078,N_957);
or U1897 (N_1897,N_1063,N_1049);
nand U1898 (N_1898,N_1402,N_1007);
nor U1899 (N_1899,N_990,N_773);
nor U1900 (N_1900,N_1052,N_1347);
nor U1901 (N_1901,N_828,N_1382);
or U1902 (N_1902,N_1053,N_973);
nor U1903 (N_1903,N_989,N_1358);
and U1904 (N_1904,N_766,N_973);
or U1905 (N_1905,N_973,N_1318);
nor U1906 (N_1906,N_1446,N_1209);
nor U1907 (N_1907,N_1319,N_1002);
xnor U1908 (N_1908,N_1394,N_876);
nand U1909 (N_1909,N_1064,N_1024);
xnor U1910 (N_1910,N_1404,N_1107);
nand U1911 (N_1911,N_760,N_1115);
nor U1912 (N_1912,N_1476,N_912);
or U1913 (N_1913,N_967,N_942);
nand U1914 (N_1914,N_1081,N_1030);
and U1915 (N_1915,N_1379,N_1453);
xor U1916 (N_1916,N_865,N_1445);
or U1917 (N_1917,N_1227,N_986);
nand U1918 (N_1918,N_1031,N_1191);
and U1919 (N_1919,N_877,N_820);
nor U1920 (N_1920,N_1370,N_1128);
or U1921 (N_1921,N_1283,N_1339);
nor U1922 (N_1922,N_1432,N_993);
nor U1923 (N_1923,N_879,N_1357);
nor U1924 (N_1924,N_1476,N_1252);
or U1925 (N_1925,N_966,N_1288);
or U1926 (N_1926,N_1266,N_995);
nor U1927 (N_1927,N_957,N_873);
and U1928 (N_1928,N_797,N_819);
nand U1929 (N_1929,N_964,N_1431);
nor U1930 (N_1930,N_1328,N_1316);
or U1931 (N_1931,N_1154,N_1242);
nor U1932 (N_1932,N_957,N_1021);
xor U1933 (N_1933,N_1172,N_787);
xor U1934 (N_1934,N_944,N_1107);
nand U1935 (N_1935,N_1192,N_1087);
nor U1936 (N_1936,N_958,N_1389);
xor U1937 (N_1937,N_1449,N_1459);
nand U1938 (N_1938,N_1148,N_1023);
nor U1939 (N_1939,N_760,N_781);
nor U1940 (N_1940,N_774,N_870);
nor U1941 (N_1941,N_1334,N_782);
and U1942 (N_1942,N_855,N_874);
nand U1943 (N_1943,N_944,N_1351);
or U1944 (N_1944,N_993,N_827);
nor U1945 (N_1945,N_1030,N_1315);
xnor U1946 (N_1946,N_942,N_1225);
nand U1947 (N_1947,N_944,N_1321);
nor U1948 (N_1948,N_787,N_756);
and U1949 (N_1949,N_1358,N_1457);
and U1950 (N_1950,N_1203,N_864);
and U1951 (N_1951,N_1119,N_1077);
nand U1952 (N_1952,N_1135,N_895);
nand U1953 (N_1953,N_824,N_1149);
nor U1954 (N_1954,N_1368,N_1123);
nor U1955 (N_1955,N_1005,N_1314);
nand U1956 (N_1956,N_763,N_1156);
or U1957 (N_1957,N_924,N_1253);
nor U1958 (N_1958,N_1164,N_1419);
or U1959 (N_1959,N_1124,N_768);
and U1960 (N_1960,N_1345,N_1083);
nor U1961 (N_1961,N_1372,N_947);
nand U1962 (N_1962,N_1006,N_1261);
or U1963 (N_1963,N_756,N_1495);
xor U1964 (N_1964,N_1323,N_841);
nand U1965 (N_1965,N_923,N_1125);
nand U1966 (N_1966,N_1198,N_1176);
xor U1967 (N_1967,N_900,N_1149);
nor U1968 (N_1968,N_1338,N_1377);
nand U1969 (N_1969,N_1488,N_1077);
nor U1970 (N_1970,N_1194,N_1456);
xnor U1971 (N_1971,N_1364,N_1189);
nand U1972 (N_1972,N_885,N_1037);
nor U1973 (N_1973,N_966,N_1123);
nor U1974 (N_1974,N_1203,N_1202);
and U1975 (N_1975,N_818,N_811);
xor U1976 (N_1976,N_1225,N_1293);
xnor U1977 (N_1977,N_950,N_891);
and U1978 (N_1978,N_1336,N_1064);
and U1979 (N_1979,N_1246,N_988);
and U1980 (N_1980,N_1262,N_922);
xnor U1981 (N_1981,N_1179,N_1181);
and U1982 (N_1982,N_1419,N_1323);
nor U1983 (N_1983,N_1124,N_823);
nor U1984 (N_1984,N_784,N_1111);
and U1985 (N_1985,N_821,N_1428);
or U1986 (N_1986,N_1036,N_892);
or U1987 (N_1987,N_1288,N_880);
nor U1988 (N_1988,N_1184,N_1013);
nand U1989 (N_1989,N_986,N_1238);
or U1990 (N_1990,N_806,N_1061);
nand U1991 (N_1991,N_946,N_1402);
nor U1992 (N_1992,N_873,N_1040);
or U1993 (N_1993,N_845,N_1339);
nor U1994 (N_1994,N_765,N_1194);
and U1995 (N_1995,N_876,N_1343);
nand U1996 (N_1996,N_942,N_1247);
xor U1997 (N_1997,N_1105,N_1449);
nor U1998 (N_1998,N_894,N_885);
and U1999 (N_1999,N_850,N_1423);
nand U2000 (N_2000,N_1210,N_1149);
xnor U2001 (N_2001,N_952,N_1241);
or U2002 (N_2002,N_799,N_1119);
or U2003 (N_2003,N_990,N_851);
and U2004 (N_2004,N_1462,N_1025);
xor U2005 (N_2005,N_930,N_852);
nand U2006 (N_2006,N_821,N_1377);
xnor U2007 (N_2007,N_811,N_1189);
xor U2008 (N_2008,N_928,N_977);
and U2009 (N_2009,N_1345,N_785);
or U2010 (N_2010,N_944,N_836);
and U2011 (N_2011,N_1044,N_1191);
xor U2012 (N_2012,N_949,N_880);
and U2013 (N_2013,N_1384,N_918);
and U2014 (N_2014,N_1391,N_879);
xnor U2015 (N_2015,N_767,N_931);
nor U2016 (N_2016,N_1324,N_977);
or U2017 (N_2017,N_1169,N_1031);
nand U2018 (N_2018,N_865,N_1118);
or U2019 (N_2019,N_1496,N_1370);
and U2020 (N_2020,N_1135,N_973);
xnor U2021 (N_2021,N_1398,N_1130);
xor U2022 (N_2022,N_1409,N_1464);
or U2023 (N_2023,N_1096,N_1277);
or U2024 (N_2024,N_1498,N_1184);
or U2025 (N_2025,N_1019,N_1302);
and U2026 (N_2026,N_1467,N_750);
and U2027 (N_2027,N_1301,N_1005);
nand U2028 (N_2028,N_842,N_890);
xnor U2029 (N_2029,N_1073,N_1070);
nand U2030 (N_2030,N_946,N_992);
and U2031 (N_2031,N_871,N_1120);
xnor U2032 (N_2032,N_1152,N_972);
xnor U2033 (N_2033,N_1462,N_1302);
and U2034 (N_2034,N_807,N_1082);
or U2035 (N_2035,N_797,N_1469);
and U2036 (N_2036,N_1149,N_1207);
or U2037 (N_2037,N_929,N_792);
and U2038 (N_2038,N_791,N_1325);
and U2039 (N_2039,N_1159,N_1499);
nand U2040 (N_2040,N_1159,N_1200);
xor U2041 (N_2041,N_947,N_1137);
and U2042 (N_2042,N_849,N_1313);
or U2043 (N_2043,N_986,N_1299);
nor U2044 (N_2044,N_826,N_1031);
nor U2045 (N_2045,N_1146,N_1195);
xnor U2046 (N_2046,N_809,N_872);
nor U2047 (N_2047,N_792,N_1029);
xor U2048 (N_2048,N_942,N_1384);
xnor U2049 (N_2049,N_1476,N_1350);
and U2050 (N_2050,N_1384,N_1432);
or U2051 (N_2051,N_813,N_1270);
and U2052 (N_2052,N_1437,N_1083);
xnor U2053 (N_2053,N_999,N_1385);
nor U2054 (N_2054,N_920,N_1355);
xor U2055 (N_2055,N_1234,N_945);
nand U2056 (N_2056,N_1362,N_1352);
or U2057 (N_2057,N_780,N_1015);
nor U2058 (N_2058,N_1410,N_795);
nor U2059 (N_2059,N_1302,N_1441);
nand U2060 (N_2060,N_1131,N_1485);
or U2061 (N_2061,N_1109,N_1349);
xnor U2062 (N_2062,N_1290,N_991);
nor U2063 (N_2063,N_965,N_929);
xor U2064 (N_2064,N_1091,N_879);
nand U2065 (N_2065,N_871,N_1118);
xnor U2066 (N_2066,N_905,N_878);
and U2067 (N_2067,N_1154,N_1257);
nor U2068 (N_2068,N_930,N_1398);
xnor U2069 (N_2069,N_979,N_1141);
nor U2070 (N_2070,N_1425,N_924);
nor U2071 (N_2071,N_1397,N_1305);
and U2072 (N_2072,N_1247,N_1131);
or U2073 (N_2073,N_1003,N_1232);
nor U2074 (N_2074,N_908,N_1049);
and U2075 (N_2075,N_1343,N_1314);
or U2076 (N_2076,N_1456,N_800);
and U2077 (N_2077,N_1003,N_1458);
or U2078 (N_2078,N_907,N_836);
nor U2079 (N_2079,N_1205,N_1254);
or U2080 (N_2080,N_1113,N_1290);
nand U2081 (N_2081,N_1239,N_1421);
xnor U2082 (N_2082,N_1250,N_1130);
nor U2083 (N_2083,N_1205,N_1497);
or U2084 (N_2084,N_1178,N_1171);
and U2085 (N_2085,N_1081,N_1366);
nand U2086 (N_2086,N_881,N_837);
nand U2087 (N_2087,N_1258,N_888);
or U2088 (N_2088,N_804,N_937);
or U2089 (N_2089,N_890,N_1320);
nor U2090 (N_2090,N_1483,N_995);
nand U2091 (N_2091,N_1114,N_896);
and U2092 (N_2092,N_1278,N_963);
and U2093 (N_2093,N_1372,N_762);
xnor U2094 (N_2094,N_1402,N_1417);
nand U2095 (N_2095,N_1384,N_1466);
and U2096 (N_2096,N_1273,N_1380);
nor U2097 (N_2097,N_1323,N_968);
nand U2098 (N_2098,N_1317,N_1212);
xor U2099 (N_2099,N_790,N_1482);
or U2100 (N_2100,N_916,N_935);
and U2101 (N_2101,N_1451,N_1318);
or U2102 (N_2102,N_1248,N_967);
xnor U2103 (N_2103,N_863,N_1244);
xor U2104 (N_2104,N_1138,N_763);
nand U2105 (N_2105,N_1362,N_1348);
and U2106 (N_2106,N_1347,N_1065);
nor U2107 (N_2107,N_1279,N_1146);
nand U2108 (N_2108,N_1013,N_1024);
xnor U2109 (N_2109,N_1217,N_938);
and U2110 (N_2110,N_1064,N_776);
nand U2111 (N_2111,N_1220,N_876);
and U2112 (N_2112,N_1342,N_844);
nand U2113 (N_2113,N_785,N_1182);
or U2114 (N_2114,N_1320,N_1072);
nor U2115 (N_2115,N_1236,N_1045);
and U2116 (N_2116,N_1018,N_993);
xor U2117 (N_2117,N_1253,N_1043);
and U2118 (N_2118,N_1104,N_960);
or U2119 (N_2119,N_1375,N_1233);
nand U2120 (N_2120,N_1489,N_1088);
and U2121 (N_2121,N_1308,N_1459);
xor U2122 (N_2122,N_1406,N_874);
and U2123 (N_2123,N_762,N_824);
nand U2124 (N_2124,N_1275,N_1000);
nor U2125 (N_2125,N_929,N_1417);
nand U2126 (N_2126,N_1244,N_1002);
xnor U2127 (N_2127,N_1193,N_1051);
xnor U2128 (N_2128,N_945,N_939);
xnor U2129 (N_2129,N_1263,N_853);
and U2130 (N_2130,N_1072,N_966);
xor U2131 (N_2131,N_1159,N_1267);
or U2132 (N_2132,N_1215,N_1400);
and U2133 (N_2133,N_893,N_1420);
or U2134 (N_2134,N_1451,N_1300);
and U2135 (N_2135,N_1045,N_1195);
nor U2136 (N_2136,N_1459,N_1375);
nor U2137 (N_2137,N_1360,N_891);
or U2138 (N_2138,N_1139,N_1417);
and U2139 (N_2139,N_1127,N_1497);
and U2140 (N_2140,N_1077,N_1155);
nand U2141 (N_2141,N_951,N_1200);
and U2142 (N_2142,N_1328,N_826);
xnor U2143 (N_2143,N_926,N_1237);
or U2144 (N_2144,N_1013,N_1272);
xnor U2145 (N_2145,N_1221,N_1316);
or U2146 (N_2146,N_822,N_1012);
xnor U2147 (N_2147,N_1025,N_942);
or U2148 (N_2148,N_949,N_1153);
nor U2149 (N_2149,N_1168,N_857);
nand U2150 (N_2150,N_914,N_1018);
nand U2151 (N_2151,N_906,N_812);
xor U2152 (N_2152,N_930,N_1016);
nor U2153 (N_2153,N_1307,N_1013);
xnor U2154 (N_2154,N_824,N_1145);
and U2155 (N_2155,N_1311,N_1414);
xor U2156 (N_2156,N_1290,N_1224);
nor U2157 (N_2157,N_1158,N_1029);
and U2158 (N_2158,N_1478,N_1023);
nand U2159 (N_2159,N_1060,N_853);
xnor U2160 (N_2160,N_1079,N_1367);
or U2161 (N_2161,N_1227,N_1048);
nor U2162 (N_2162,N_754,N_1496);
xnor U2163 (N_2163,N_794,N_942);
and U2164 (N_2164,N_1453,N_1203);
or U2165 (N_2165,N_1453,N_1194);
nor U2166 (N_2166,N_1066,N_941);
or U2167 (N_2167,N_1083,N_1070);
nand U2168 (N_2168,N_953,N_1375);
or U2169 (N_2169,N_865,N_1337);
xnor U2170 (N_2170,N_1327,N_774);
or U2171 (N_2171,N_885,N_1295);
xnor U2172 (N_2172,N_1007,N_1485);
or U2173 (N_2173,N_1357,N_852);
or U2174 (N_2174,N_1279,N_969);
nand U2175 (N_2175,N_751,N_791);
nor U2176 (N_2176,N_916,N_1311);
nand U2177 (N_2177,N_867,N_1092);
and U2178 (N_2178,N_1251,N_1488);
xor U2179 (N_2179,N_861,N_1367);
nor U2180 (N_2180,N_1141,N_1453);
or U2181 (N_2181,N_780,N_1448);
xor U2182 (N_2182,N_805,N_1416);
or U2183 (N_2183,N_1489,N_1065);
xor U2184 (N_2184,N_1454,N_1296);
xor U2185 (N_2185,N_1052,N_1119);
or U2186 (N_2186,N_1097,N_1342);
or U2187 (N_2187,N_1227,N_796);
or U2188 (N_2188,N_954,N_1208);
xnor U2189 (N_2189,N_1142,N_795);
nor U2190 (N_2190,N_793,N_1403);
or U2191 (N_2191,N_1242,N_1408);
and U2192 (N_2192,N_844,N_947);
xor U2193 (N_2193,N_1038,N_1170);
or U2194 (N_2194,N_1412,N_869);
nor U2195 (N_2195,N_847,N_1325);
and U2196 (N_2196,N_1078,N_1076);
or U2197 (N_2197,N_1078,N_1446);
nand U2198 (N_2198,N_1327,N_1346);
and U2199 (N_2199,N_1128,N_1394);
and U2200 (N_2200,N_851,N_854);
nand U2201 (N_2201,N_1470,N_1122);
nor U2202 (N_2202,N_776,N_824);
and U2203 (N_2203,N_1017,N_1331);
nand U2204 (N_2204,N_794,N_1176);
nor U2205 (N_2205,N_1024,N_989);
nand U2206 (N_2206,N_916,N_1383);
and U2207 (N_2207,N_753,N_1162);
and U2208 (N_2208,N_1477,N_1360);
xor U2209 (N_2209,N_1352,N_1471);
or U2210 (N_2210,N_1406,N_1309);
xor U2211 (N_2211,N_1060,N_1413);
xor U2212 (N_2212,N_1163,N_1428);
or U2213 (N_2213,N_1089,N_1226);
or U2214 (N_2214,N_1017,N_1276);
nor U2215 (N_2215,N_893,N_1213);
xnor U2216 (N_2216,N_899,N_1449);
xor U2217 (N_2217,N_1097,N_765);
nor U2218 (N_2218,N_1368,N_1418);
and U2219 (N_2219,N_833,N_1193);
or U2220 (N_2220,N_1477,N_841);
nor U2221 (N_2221,N_1418,N_1057);
or U2222 (N_2222,N_1060,N_1235);
nor U2223 (N_2223,N_886,N_850);
xnor U2224 (N_2224,N_816,N_948);
and U2225 (N_2225,N_1484,N_791);
nor U2226 (N_2226,N_1145,N_958);
or U2227 (N_2227,N_808,N_1442);
or U2228 (N_2228,N_1402,N_982);
nand U2229 (N_2229,N_786,N_775);
nor U2230 (N_2230,N_941,N_1241);
or U2231 (N_2231,N_866,N_831);
nor U2232 (N_2232,N_1055,N_1115);
nand U2233 (N_2233,N_1076,N_1182);
nand U2234 (N_2234,N_943,N_1245);
nand U2235 (N_2235,N_774,N_811);
nor U2236 (N_2236,N_1133,N_1387);
xor U2237 (N_2237,N_1199,N_917);
xnor U2238 (N_2238,N_961,N_1451);
nand U2239 (N_2239,N_1425,N_892);
nand U2240 (N_2240,N_1130,N_768);
or U2241 (N_2241,N_885,N_1300);
xnor U2242 (N_2242,N_1151,N_956);
xor U2243 (N_2243,N_1443,N_1356);
and U2244 (N_2244,N_1177,N_1335);
nor U2245 (N_2245,N_937,N_1267);
nor U2246 (N_2246,N_1148,N_1156);
and U2247 (N_2247,N_1236,N_1097);
xor U2248 (N_2248,N_1087,N_920);
or U2249 (N_2249,N_1072,N_1084);
or U2250 (N_2250,N_1521,N_1987);
or U2251 (N_2251,N_1792,N_2011);
and U2252 (N_2252,N_1804,N_2096);
or U2253 (N_2253,N_2065,N_1964);
and U2254 (N_2254,N_2063,N_2099);
xor U2255 (N_2255,N_1678,N_2037);
nand U2256 (N_2256,N_2050,N_2212);
xor U2257 (N_2257,N_1886,N_1864);
nand U2258 (N_2258,N_1865,N_2126);
or U2259 (N_2259,N_1984,N_2129);
nor U2260 (N_2260,N_2230,N_1978);
and U2261 (N_2261,N_1879,N_2058);
nor U2262 (N_2262,N_1797,N_2167);
nor U2263 (N_2263,N_1663,N_1604);
and U2264 (N_2264,N_2205,N_2130);
or U2265 (N_2265,N_1893,N_1715);
nor U2266 (N_2266,N_1720,N_1581);
or U2267 (N_2267,N_1747,N_1700);
and U2268 (N_2268,N_2054,N_1749);
nor U2269 (N_2269,N_2172,N_1901);
xor U2270 (N_2270,N_1612,N_1946);
and U2271 (N_2271,N_2202,N_2238);
and U2272 (N_2272,N_2155,N_1807);
and U2273 (N_2273,N_2068,N_1756);
nor U2274 (N_2274,N_1955,N_2215);
nor U2275 (N_2275,N_1515,N_1600);
nor U2276 (N_2276,N_1814,N_1971);
nor U2277 (N_2277,N_1793,N_1989);
nor U2278 (N_2278,N_1525,N_1970);
or U2279 (N_2279,N_1800,N_2176);
xnor U2280 (N_2280,N_1717,N_1507);
nor U2281 (N_2281,N_2119,N_1991);
nor U2282 (N_2282,N_2049,N_1550);
nor U2283 (N_2283,N_1707,N_1504);
and U2284 (N_2284,N_2061,N_1687);
and U2285 (N_2285,N_2160,N_1783);
nand U2286 (N_2286,N_2208,N_1745);
and U2287 (N_2287,N_1968,N_1874);
nor U2288 (N_2288,N_2234,N_1895);
xnor U2289 (N_2289,N_2093,N_1727);
nand U2290 (N_2290,N_2200,N_2169);
nand U2291 (N_2291,N_1817,N_2152);
nand U2292 (N_2292,N_1579,N_1966);
nand U2293 (N_2293,N_1734,N_2243);
and U2294 (N_2294,N_1796,N_1698);
nor U2295 (N_2295,N_1903,N_1902);
nand U2296 (N_2296,N_1860,N_1910);
nor U2297 (N_2297,N_1670,N_1780);
xnor U2298 (N_2298,N_1943,N_1643);
nand U2299 (N_2299,N_1812,N_1679);
and U2300 (N_2300,N_1650,N_1706);
or U2301 (N_2301,N_1543,N_1832);
and U2302 (N_2302,N_1609,N_1854);
nand U2303 (N_2303,N_1847,N_2166);
nand U2304 (N_2304,N_2240,N_1782);
nand U2305 (N_2305,N_1763,N_1922);
xor U2306 (N_2306,N_2123,N_1787);
xor U2307 (N_2307,N_1620,N_1969);
xor U2308 (N_2308,N_1956,N_2084);
nand U2309 (N_2309,N_2022,N_2016);
nor U2310 (N_2310,N_2007,N_1547);
nor U2311 (N_2311,N_1658,N_2105);
xor U2312 (N_2312,N_1960,N_1795);
and U2313 (N_2313,N_2122,N_1798);
and U2314 (N_2314,N_1733,N_1644);
xnor U2315 (N_2315,N_1574,N_1711);
nand U2316 (N_2316,N_1685,N_1501);
xnor U2317 (N_2317,N_1815,N_1738);
nor U2318 (N_2318,N_1597,N_2070);
or U2319 (N_2319,N_1988,N_1545);
nand U2320 (N_2320,N_2199,N_2170);
xor U2321 (N_2321,N_1889,N_1518);
nand U2322 (N_2322,N_1646,N_1615);
and U2323 (N_2323,N_1535,N_2127);
nor U2324 (N_2324,N_1972,N_2108);
or U2325 (N_2325,N_1843,N_1746);
nor U2326 (N_2326,N_1858,N_1775);
or U2327 (N_2327,N_2125,N_1630);
xnor U2328 (N_2328,N_1911,N_1701);
or U2329 (N_2329,N_1973,N_1994);
nor U2330 (N_2330,N_1769,N_1674);
nand U2331 (N_2331,N_2110,N_1666);
or U2332 (N_2332,N_1710,N_1827);
xor U2333 (N_2333,N_1506,N_2048);
or U2334 (N_2334,N_1870,N_1526);
nor U2335 (N_2335,N_1880,N_1849);
xnor U2336 (N_2336,N_1686,N_1897);
nand U2337 (N_2337,N_1824,N_1592);
nor U2338 (N_2338,N_1873,N_2220);
and U2339 (N_2339,N_1781,N_1764);
xnor U2340 (N_2340,N_1513,N_1801);
nor U2341 (N_2341,N_1836,N_2174);
nor U2342 (N_2342,N_1754,N_2005);
and U2343 (N_2343,N_2087,N_1599);
nand U2344 (N_2344,N_1912,N_1657);
nor U2345 (N_2345,N_2203,N_1534);
nor U2346 (N_2346,N_1840,N_2244);
xnor U2347 (N_2347,N_2227,N_2221);
nand U2348 (N_2348,N_1790,N_1692);
xnor U2349 (N_2349,N_1726,N_2144);
nand U2350 (N_2350,N_1661,N_1928);
and U2351 (N_2351,N_2242,N_1786);
xor U2352 (N_2352,N_2235,N_1848);
xnor U2353 (N_2353,N_1983,N_1605);
nor U2354 (N_2354,N_2150,N_2164);
nor U2355 (N_2355,N_2131,N_1736);
and U2356 (N_2356,N_1993,N_1582);
or U2357 (N_2357,N_1565,N_1938);
or U2358 (N_2358,N_1958,N_1841);
xor U2359 (N_2359,N_1751,N_1779);
or U2360 (N_2360,N_1619,N_1869);
nor U2361 (N_2361,N_1926,N_2113);
or U2362 (N_2362,N_2028,N_1583);
nor U2363 (N_2363,N_2025,N_2153);
or U2364 (N_2364,N_1693,N_1768);
and U2365 (N_2365,N_1682,N_2151);
or U2366 (N_2366,N_2219,N_1681);
and U2367 (N_2367,N_1549,N_1668);
nor U2368 (N_2368,N_1859,N_1766);
or U2369 (N_2369,N_2083,N_2239);
nor U2370 (N_2370,N_1940,N_1566);
nand U2371 (N_2371,N_1555,N_2159);
nor U2372 (N_2372,N_2165,N_2080);
or U2373 (N_2373,N_1514,N_1662);
and U2374 (N_2374,N_1923,N_2141);
xnor U2375 (N_2375,N_1502,N_1517);
and U2376 (N_2376,N_2228,N_2034);
nor U2377 (N_2377,N_2038,N_2211);
nor U2378 (N_2378,N_1632,N_1559);
or U2379 (N_2379,N_2163,N_1997);
or U2380 (N_2380,N_2232,N_1572);
nor U2381 (N_2381,N_2222,N_1721);
nor U2382 (N_2382,N_1810,N_1825);
and U2383 (N_2383,N_1838,N_2161);
nand U2384 (N_2384,N_1982,N_1683);
nand U2385 (N_2385,N_1741,N_1739);
or U2386 (N_2386,N_2157,N_2006);
and U2387 (N_2387,N_1755,N_1742);
or U2388 (N_2388,N_2008,N_1845);
or U2389 (N_2389,N_1837,N_2075);
or U2390 (N_2390,N_2020,N_1919);
and U2391 (N_2391,N_1607,N_2158);
nor U2392 (N_2392,N_1640,N_2001);
xnor U2393 (N_2393,N_1877,N_1918);
or U2394 (N_2394,N_2247,N_1974);
nand U2395 (N_2395,N_1732,N_2079);
xnor U2396 (N_2396,N_2014,N_1820);
and U2397 (N_2397,N_1855,N_1842);
or U2398 (N_2398,N_2194,N_1653);
xnor U2399 (N_2399,N_2109,N_1618);
or U2400 (N_2400,N_1949,N_1907);
xnor U2401 (N_2401,N_2004,N_2045);
and U2402 (N_2402,N_1505,N_2002);
or U2403 (N_2403,N_2095,N_1729);
or U2404 (N_2404,N_2135,N_2017);
nand U2405 (N_2405,N_1558,N_1771);
and U2406 (N_2406,N_1649,N_1999);
and U2407 (N_2407,N_2100,N_1676);
nand U2408 (N_2408,N_2101,N_1688);
nor U2409 (N_2409,N_1977,N_1882);
xor U2410 (N_2410,N_1906,N_2213);
or U2411 (N_2411,N_1713,N_1696);
nor U2412 (N_2412,N_1799,N_1898);
and U2413 (N_2413,N_1675,N_1896);
nor U2414 (N_2414,N_2206,N_2249);
xnor U2415 (N_2415,N_1709,N_1917);
and U2416 (N_2416,N_1740,N_1654);
nand U2417 (N_2417,N_1806,N_1638);
and U2418 (N_2418,N_1627,N_1611);
xnor U2419 (N_2419,N_1703,N_2140);
nor U2420 (N_2420,N_2223,N_2031);
xnor U2421 (N_2421,N_1932,N_1635);
nor U2422 (N_2422,N_1822,N_1636);
nor U2423 (N_2423,N_2055,N_1894);
xor U2424 (N_2424,N_2074,N_1631);
or U2425 (N_2425,N_2188,N_1878);
nand U2426 (N_2426,N_1762,N_1951);
or U2427 (N_2427,N_1996,N_2143);
or U2428 (N_2428,N_1594,N_1965);
xnor U2429 (N_2429,N_1660,N_2136);
nand U2430 (N_2430,N_1705,N_1899);
or U2431 (N_2431,N_1595,N_1770);
or U2432 (N_2432,N_1778,N_1908);
or U2433 (N_2433,N_1765,N_1818);
or U2434 (N_2434,N_2069,N_1823);
xnor U2435 (N_2435,N_2046,N_2175);
xnor U2436 (N_2436,N_1867,N_1881);
xor U2437 (N_2437,N_1642,N_1924);
nand U2438 (N_2438,N_2116,N_1725);
nand U2439 (N_2439,N_1816,N_2104);
xnor U2440 (N_2440,N_2179,N_1904);
xnor U2441 (N_2441,N_1890,N_2012);
or U2442 (N_2442,N_1563,N_1761);
nand U2443 (N_2443,N_2111,N_1861);
xnor U2444 (N_2444,N_2177,N_2027);
xnor U2445 (N_2445,N_1645,N_1937);
nor U2446 (N_2446,N_1655,N_1634);
or U2447 (N_2447,N_1524,N_1647);
xnor U2448 (N_2448,N_1708,N_1578);
nor U2449 (N_2449,N_2142,N_1830);
xor U2450 (N_2450,N_2071,N_2224);
xor U2451 (N_2451,N_1617,N_1641);
nor U2452 (N_2452,N_1509,N_2032);
or U2453 (N_2453,N_1735,N_1500);
xnor U2454 (N_2454,N_2021,N_2145);
xor U2455 (N_2455,N_2193,N_1802);
nand U2456 (N_2456,N_2197,N_2088);
nor U2457 (N_2457,N_2191,N_2236);
xor U2458 (N_2458,N_1794,N_1856);
nor U2459 (N_2459,N_1748,N_1819);
or U2460 (N_2460,N_1834,N_2216);
and U2461 (N_2461,N_1892,N_2039);
xor U2462 (N_2462,N_1690,N_1835);
nor U2463 (N_2463,N_1979,N_1998);
xnor U2464 (N_2464,N_1909,N_2214);
xor U2465 (N_2465,N_1571,N_1995);
and U2466 (N_2466,N_1954,N_1750);
and U2467 (N_2467,N_2178,N_1947);
and U2468 (N_2468,N_1875,N_1633);
xnor U2469 (N_2469,N_2225,N_2098);
and U2470 (N_2470,N_1531,N_1961);
nor U2471 (N_2471,N_1624,N_1863);
and U2472 (N_2472,N_1557,N_1689);
and U2473 (N_2473,N_1637,N_1844);
nand U2474 (N_2474,N_1546,N_2052);
and U2475 (N_2475,N_1811,N_1813);
nand U2476 (N_2476,N_2231,N_2066);
or U2477 (N_2477,N_2171,N_1850);
nor U2478 (N_2478,N_1744,N_1948);
xnor U2479 (N_2479,N_2138,N_2137);
xnor U2480 (N_2480,N_1933,N_2128);
or U2481 (N_2481,N_2024,N_1503);
xnor U2482 (N_2482,N_1610,N_1785);
nand U2483 (N_2483,N_2040,N_1665);
and U2484 (N_2484,N_1914,N_2204);
nand U2485 (N_2485,N_2187,N_2154);
or U2486 (N_2486,N_2033,N_1602);
xor U2487 (N_2487,N_2036,N_1936);
xor U2488 (N_2488,N_1639,N_1872);
or U2489 (N_2489,N_1986,N_2076);
xor U2490 (N_2490,N_2091,N_1772);
and U2491 (N_2491,N_1731,N_1934);
nor U2492 (N_2492,N_1885,N_2009);
nor U2493 (N_2493,N_1510,N_1608);
nand U2494 (N_2494,N_2156,N_1803);
and U2495 (N_2495,N_1833,N_1808);
nand U2496 (N_2496,N_1539,N_2015);
xnor U2497 (N_2497,N_1930,N_2062);
xnor U2498 (N_2498,N_2134,N_1536);
nor U2499 (N_2499,N_1829,N_1699);
xor U2500 (N_2500,N_2162,N_1629);
nand U2501 (N_2501,N_1588,N_2233);
and U2502 (N_2502,N_1552,N_2000);
and U2503 (N_2503,N_2117,N_2120);
and U2504 (N_2504,N_1883,N_2018);
and U2505 (N_2505,N_1931,N_2090);
and U2506 (N_2506,N_1743,N_1718);
and U2507 (N_2507,N_1656,N_1585);
and U2508 (N_2508,N_2185,N_1777);
xnor U2509 (N_2509,N_2189,N_1564);
xor U2510 (N_2510,N_2064,N_1520);
nor U2511 (N_2511,N_1680,N_1598);
xnor U2512 (N_2512,N_2073,N_2181);
and U2513 (N_2513,N_1773,N_1568);
xnor U2514 (N_2514,N_1508,N_1788);
or U2515 (N_2515,N_1719,N_1659);
and U2516 (N_2516,N_1915,N_1759);
nor U2517 (N_2517,N_1553,N_2057);
and U2518 (N_2518,N_1570,N_2067);
or U2519 (N_2519,N_2229,N_1776);
xnor U2520 (N_2520,N_1580,N_1868);
xor U2521 (N_2521,N_1704,N_2133);
nor U2522 (N_2522,N_2148,N_1567);
xor U2523 (N_2523,N_2051,N_2026);
xor U2524 (N_2524,N_1537,N_1789);
nand U2525 (N_2525,N_1569,N_1851);
nand U2526 (N_2526,N_1957,N_1593);
or U2527 (N_2527,N_2173,N_2226);
or U2528 (N_2528,N_2201,N_1853);
or U2529 (N_2529,N_2180,N_2077);
or U2530 (N_2530,N_1826,N_2146);
or U2531 (N_2531,N_1962,N_1616);
xor U2532 (N_2532,N_1760,N_1723);
xor U2533 (N_2533,N_2198,N_2089);
nor U2534 (N_2534,N_1846,N_2210);
nand U2535 (N_2535,N_1981,N_2245);
nand U2536 (N_2536,N_1876,N_1541);
nand U2537 (N_2537,N_1540,N_1542);
nor U2538 (N_2538,N_2060,N_1603);
or U2539 (N_2539,N_1671,N_1884);
nor U2540 (N_2540,N_2072,N_1625);
or U2541 (N_2541,N_1523,N_2086);
and U2542 (N_2542,N_1621,N_1556);
nand U2543 (N_2543,N_1929,N_1925);
xor U2544 (N_2544,N_2035,N_2121);
and U2545 (N_2545,N_2047,N_1648);
and U2546 (N_2546,N_2168,N_1672);
and U2547 (N_2547,N_1577,N_1590);
or U2548 (N_2548,N_1544,N_1601);
or U2549 (N_2549,N_2023,N_1554);
nor U2550 (N_2550,N_1652,N_1712);
xor U2551 (N_2551,N_1888,N_2114);
or U2552 (N_2552,N_2184,N_2097);
or U2553 (N_2553,N_2209,N_1606);
nand U2554 (N_2554,N_2010,N_1673);
nor U2555 (N_2555,N_1677,N_1664);
xnor U2556 (N_2556,N_1623,N_1560);
or U2557 (N_2557,N_2041,N_1691);
nor U2558 (N_2558,N_2092,N_1767);
nand U2559 (N_2559,N_1774,N_1573);
xnor U2560 (N_2560,N_1697,N_1828);
xnor U2561 (N_2561,N_2081,N_2044);
or U2562 (N_2562,N_2132,N_1791);
or U2563 (N_2563,N_2147,N_1952);
xor U2564 (N_2564,N_1941,N_2078);
nand U2565 (N_2565,N_1651,N_1942);
nand U2566 (N_2566,N_1913,N_1512);
and U2567 (N_2567,N_1730,N_1905);
nand U2568 (N_2568,N_1626,N_1939);
and U2569 (N_2569,N_1562,N_1587);
xor U2570 (N_2570,N_1728,N_1866);
xor U2571 (N_2571,N_1591,N_1667);
nor U2572 (N_2572,N_1530,N_2102);
nand U2573 (N_2573,N_2218,N_1722);
and U2574 (N_2574,N_1809,N_2019);
or U2575 (N_2575,N_1967,N_2237);
xnor U2576 (N_2576,N_1519,N_1529);
and U2577 (N_2577,N_2192,N_1980);
nor U2578 (N_2578,N_2059,N_2182);
and U2579 (N_2579,N_1784,N_1945);
or U2580 (N_2580,N_2118,N_2139);
nor U2581 (N_2581,N_1857,N_2082);
and U2582 (N_2582,N_1992,N_1758);
nand U2583 (N_2583,N_1716,N_2029);
nor U2584 (N_2584,N_1927,N_1935);
nand U2585 (N_2585,N_1737,N_1589);
xnor U2586 (N_2586,N_1596,N_1714);
or U2587 (N_2587,N_1576,N_1622);
xor U2588 (N_2588,N_2103,N_1724);
or U2589 (N_2589,N_1516,N_2124);
xor U2590 (N_2590,N_1527,N_1533);
or U2591 (N_2591,N_1891,N_2094);
xnor U2592 (N_2592,N_1528,N_1669);
or U2593 (N_2593,N_2003,N_1538);
or U2594 (N_2594,N_1551,N_1586);
nand U2595 (N_2595,N_2013,N_1821);
and U2596 (N_2596,N_2115,N_2241);
nand U2597 (N_2597,N_1613,N_2053);
nand U2598 (N_2598,N_1950,N_1921);
nor U2599 (N_2599,N_2183,N_1959);
or U2600 (N_2600,N_1702,N_2085);
xor U2601 (N_2601,N_1920,N_1548);
xor U2602 (N_2602,N_1831,N_1975);
and U2603 (N_2603,N_1985,N_1628);
and U2604 (N_2604,N_1695,N_1805);
nand U2605 (N_2605,N_2190,N_1852);
xor U2606 (N_2606,N_1684,N_2217);
nand U2607 (N_2607,N_1944,N_2207);
nor U2608 (N_2608,N_1953,N_1511);
nand U2609 (N_2609,N_2195,N_2186);
nor U2610 (N_2610,N_1614,N_1916);
or U2611 (N_2611,N_2056,N_2149);
and U2612 (N_2612,N_1887,N_2246);
nor U2613 (N_2613,N_2112,N_2042);
or U2614 (N_2614,N_1839,N_2196);
nor U2615 (N_2615,N_1753,N_2248);
or U2616 (N_2616,N_1584,N_1862);
nand U2617 (N_2617,N_2107,N_1963);
or U2618 (N_2618,N_1522,N_2106);
and U2619 (N_2619,N_1976,N_1575);
and U2620 (N_2620,N_1561,N_1990);
xor U2621 (N_2621,N_1900,N_2030);
nand U2622 (N_2622,N_1694,N_1532);
nor U2623 (N_2623,N_2043,N_1757);
xnor U2624 (N_2624,N_1752,N_1871);
or U2625 (N_2625,N_2029,N_1826);
nor U2626 (N_2626,N_1711,N_2106);
xnor U2627 (N_2627,N_1790,N_1709);
nor U2628 (N_2628,N_1969,N_2212);
xnor U2629 (N_2629,N_1955,N_2048);
and U2630 (N_2630,N_1521,N_1560);
xor U2631 (N_2631,N_1632,N_2244);
xor U2632 (N_2632,N_1744,N_1611);
and U2633 (N_2633,N_1890,N_2017);
nand U2634 (N_2634,N_2117,N_1868);
and U2635 (N_2635,N_1510,N_1873);
and U2636 (N_2636,N_2197,N_2024);
or U2637 (N_2637,N_2211,N_1674);
xor U2638 (N_2638,N_2100,N_2198);
nand U2639 (N_2639,N_2220,N_1879);
xnor U2640 (N_2640,N_2193,N_1780);
nand U2641 (N_2641,N_1808,N_2096);
nor U2642 (N_2642,N_1961,N_2071);
nand U2643 (N_2643,N_1968,N_1921);
nor U2644 (N_2644,N_1682,N_1805);
xor U2645 (N_2645,N_1887,N_2102);
nor U2646 (N_2646,N_1692,N_1878);
or U2647 (N_2647,N_1776,N_1690);
xnor U2648 (N_2648,N_1629,N_1667);
and U2649 (N_2649,N_1767,N_1668);
nor U2650 (N_2650,N_2135,N_2060);
xor U2651 (N_2651,N_2092,N_1717);
or U2652 (N_2652,N_2210,N_2225);
nand U2653 (N_2653,N_2126,N_2141);
nand U2654 (N_2654,N_1795,N_1610);
or U2655 (N_2655,N_2192,N_1762);
and U2656 (N_2656,N_1538,N_1811);
and U2657 (N_2657,N_1715,N_1760);
nor U2658 (N_2658,N_2144,N_1697);
nor U2659 (N_2659,N_1653,N_1890);
nand U2660 (N_2660,N_1849,N_1939);
or U2661 (N_2661,N_1724,N_2096);
xor U2662 (N_2662,N_1769,N_1766);
nor U2663 (N_2663,N_1553,N_1897);
nor U2664 (N_2664,N_1573,N_2099);
or U2665 (N_2665,N_2098,N_1830);
and U2666 (N_2666,N_1947,N_1814);
xor U2667 (N_2667,N_1813,N_1575);
nor U2668 (N_2668,N_1896,N_2194);
or U2669 (N_2669,N_1722,N_1823);
xor U2670 (N_2670,N_1939,N_1764);
and U2671 (N_2671,N_2210,N_1785);
nor U2672 (N_2672,N_1769,N_1970);
or U2673 (N_2673,N_1763,N_1613);
xnor U2674 (N_2674,N_1736,N_1819);
or U2675 (N_2675,N_2117,N_1605);
xnor U2676 (N_2676,N_1997,N_1671);
or U2677 (N_2677,N_1947,N_1696);
or U2678 (N_2678,N_1553,N_1536);
or U2679 (N_2679,N_1586,N_2162);
or U2680 (N_2680,N_2172,N_1532);
nor U2681 (N_2681,N_1873,N_2245);
or U2682 (N_2682,N_1799,N_1917);
or U2683 (N_2683,N_1782,N_1762);
xnor U2684 (N_2684,N_1793,N_1839);
and U2685 (N_2685,N_1764,N_2134);
or U2686 (N_2686,N_2187,N_1556);
or U2687 (N_2687,N_2204,N_1974);
nand U2688 (N_2688,N_1522,N_1792);
and U2689 (N_2689,N_1993,N_2069);
xnor U2690 (N_2690,N_2199,N_1821);
xor U2691 (N_2691,N_2147,N_1652);
or U2692 (N_2692,N_1507,N_1696);
nand U2693 (N_2693,N_2006,N_1609);
xor U2694 (N_2694,N_1745,N_1555);
nor U2695 (N_2695,N_2219,N_1981);
and U2696 (N_2696,N_2090,N_1654);
or U2697 (N_2697,N_1985,N_2228);
nor U2698 (N_2698,N_1771,N_1779);
nand U2699 (N_2699,N_1582,N_1809);
nand U2700 (N_2700,N_2022,N_1686);
or U2701 (N_2701,N_1857,N_1789);
or U2702 (N_2702,N_1605,N_1668);
xor U2703 (N_2703,N_1741,N_1568);
or U2704 (N_2704,N_1822,N_1517);
nand U2705 (N_2705,N_1506,N_2195);
xor U2706 (N_2706,N_2145,N_1956);
or U2707 (N_2707,N_2135,N_2118);
nand U2708 (N_2708,N_1738,N_1880);
or U2709 (N_2709,N_1770,N_2038);
xnor U2710 (N_2710,N_1756,N_2238);
and U2711 (N_2711,N_1666,N_2101);
and U2712 (N_2712,N_1623,N_1501);
or U2713 (N_2713,N_2248,N_1968);
and U2714 (N_2714,N_1849,N_2021);
or U2715 (N_2715,N_1538,N_1531);
xnor U2716 (N_2716,N_1723,N_2196);
nor U2717 (N_2717,N_2061,N_1923);
or U2718 (N_2718,N_2022,N_2074);
xor U2719 (N_2719,N_1964,N_1957);
and U2720 (N_2720,N_1643,N_1832);
xor U2721 (N_2721,N_1747,N_1824);
or U2722 (N_2722,N_1555,N_1744);
xnor U2723 (N_2723,N_2019,N_1742);
xnor U2724 (N_2724,N_1548,N_2108);
nor U2725 (N_2725,N_2176,N_2033);
or U2726 (N_2726,N_1955,N_2160);
or U2727 (N_2727,N_2125,N_2011);
nor U2728 (N_2728,N_1620,N_1710);
or U2729 (N_2729,N_1871,N_1819);
or U2730 (N_2730,N_1768,N_2004);
nor U2731 (N_2731,N_1569,N_1977);
xnor U2732 (N_2732,N_2053,N_2051);
nor U2733 (N_2733,N_1955,N_1858);
nand U2734 (N_2734,N_1511,N_1525);
xor U2735 (N_2735,N_2011,N_1665);
nand U2736 (N_2736,N_2002,N_1680);
nand U2737 (N_2737,N_1502,N_1604);
nor U2738 (N_2738,N_1754,N_2072);
xnor U2739 (N_2739,N_2212,N_1672);
or U2740 (N_2740,N_1852,N_1899);
nand U2741 (N_2741,N_1912,N_1651);
xor U2742 (N_2742,N_1695,N_1852);
nor U2743 (N_2743,N_1575,N_1773);
nor U2744 (N_2744,N_2069,N_1664);
nor U2745 (N_2745,N_2061,N_1770);
xor U2746 (N_2746,N_2055,N_1988);
xor U2747 (N_2747,N_2044,N_1846);
xnor U2748 (N_2748,N_2150,N_1971);
or U2749 (N_2749,N_1945,N_1630);
and U2750 (N_2750,N_1620,N_1784);
and U2751 (N_2751,N_1660,N_2244);
and U2752 (N_2752,N_2226,N_1864);
or U2753 (N_2753,N_2160,N_1873);
xor U2754 (N_2754,N_1546,N_1960);
and U2755 (N_2755,N_1974,N_2052);
nand U2756 (N_2756,N_1763,N_1902);
nand U2757 (N_2757,N_1694,N_1985);
nand U2758 (N_2758,N_1917,N_2059);
xnor U2759 (N_2759,N_1918,N_1746);
nor U2760 (N_2760,N_2172,N_1866);
or U2761 (N_2761,N_1859,N_2141);
nand U2762 (N_2762,N_2204,N_2018);
nand U2763 (N_2763,N_1964,N_1537);
nand U2764 (N_2764,N_2193,N_1941);
nor U2765 (N_2765,N_1602,N_1578);
and U2766 (N_2766,N_2159,N_1852);
and U2767 (N_2767,N_1692,N_1590);
xor U2768 (N_2768,N_1693,N_1626);
xor U2769 (N_2769,N_1660,N_2125);
nor U2770 (N_2770,N_1579,N_1752);
or U2771 (N_2771,N_1574,N_1900);
or U2772 (N_2772,N_2247,N_1552);
nor U2773 (N_2773,N_2223,N_1708);
xnor U2774 (N_2774,N_1791,N_1549);
nand U2775 (N_2775,N_2011,N_2244);
or U2776 (N_2776,N_2151,N_1993);
and U2777 (N_2777,N_1921,N_1652);
nand U2778 (N_2778,N_2148,N_1707);
xnor U2779 (N_2779,N_1557,N_1965);
nand U2780 (N_2780,N_1525,N_1947);
or U2781 (N_2781,N_1738,N_2098);
xnor U2782 (N_2782,N_1620,N_1889);
or U2783 (N_2783,N_1769,N_1551);
xnor U2784 (N_2784,N_1866,N_1643);
xnor U2785 (N_2785,N_1606,N_1560);
nor U2786 (N_2786,N_1903,N_1745);
or U2787 (N_2787,N_1851,N_1617);
or U2788 (N_2788,N_1617,N_1708);
xor U2789 (N_2789,N_1855,N_2147);
and U2790 (N_2790,N_2173,N_1806);
nand U2791 (N_2791,N_2223,N_1654);
or U2792 (N_2792,N_1635,N_2011);
nand U2793 (N_2793,N_2153,N_1934);
nor U2794 (N_2794,N_1896,N_1558);
nand U2795 (N_2795,N_1768,N_1652);
nand U2796 (N_2796,N_1893,N_1644);
nand U2797 (N_2797,N_2167,N_1829);
xnor U2798 (N_2798,N_1940,N_2091);
xnor U2799 (N_2799,N_1753,N_1847);
xnor U2800 (N_2800,N_1897,N_2045);
nand U2801 (N_2801,N_1723,N_1755);
nor U2802 (N_2802,N_2197,N_1752);
and U2803 (N_2803,N_2130,N_2224);
or U2804 (N_2804,N_1737,N_2184);
and U2805 (N_2805,N_2231,N_2164);
or U2806 (N_2806,N_1884,N_1669);
nand U2807 (N_2807,N_1739,N_1735);
nor U2808 (N_2808,N_1998,N_1507);
or U2809 (N_2809,N_1725,N_1779);
nor U2810 (N_2810,N_2084,N_1995);
xor U2811 (N_2811,N_1970,N_1833);
or U2812 (N_2812,N_1897,N_1968);
and U2813 (N_2813,N_1571,N_1633);
xor U2814 (N_2814,N_1978,N_1909);
nand U2815 (N_2815,N_2171,N_1749);
xor U2816 (N_2816,N_1635,N_1898);
nand U2817 (N_2817,N_1699,N_2207);
or U2818 (N_2818,N_2085,N_1687);
xnor U2819 (N_2819,N_2030,N_1865);
and U2820 (N_2820,N_2229,N_1566);
xnor U2821 (N_2821,N_1680,N_1608);
or U2822 (N_2822,N_2191,N_1872);
nand U2823 (N_2823,N_1906,N_1529);
xor U2824 (N_2824,N_2176,N_1818);
nor U2825 (N_2825,N_1914,N_2115);
nor U2826 (N_2826,N_1591,N_1514);
nor U2827 (N_2827,N_1723,N_1591);
nor U2828 (N_2828,N_1515,N_2160);
nor U2829 (N_2829,N_1710,N_2116);
xor U2830 (N_2830,N_1708,N_2043);
and U2831 (N_2831,N_1876,N_1805);
or U2832 (N_2832,N_2001,N_2023);
xnor U2833 (N_2833,N_1581,N_1805);
nand U2834 (N_2834,N_1503,N_1842);
nand U2835 (N_2835,N_2134,N_2228);
and U2836 (N_2836,N_2115,N_1626);
and U2837 (N_2837,N_1726,N_1555);
nand U2838 (N_2838,N_1926,N_1966);
and U2839 (N_2839,N_1515,N_1890);
xnor U2840 (N_2840,N_1633,N_1771);
nor U2841 (N_2841,N_1776,N_2214);
or U2842 (N_2842,N_1538,N_2070);
nor U2843 (N_2843,N_1705,N_2108);
xnor U2844 (N_2844,N_2124,N_1801);
xor U2845 (N_2845,N_1955,N_2142);
and U2846 (N_2846,N_1602,N_1774);
nand U2847 (N_2847,N_1528,N_1797);
nand U2848 (N_2848,N_1603,N_2096);
or U2849 (N_2849,N_1749,N_1745);
nor U2850 (N_2850,N_2042,N_1683);
and U2851 (N_2851,N_1669,N_2158);
xnor U2852 (N_2852,N_1908,N_2142);
and U2853 (N_2853,N_2066,N_1561);
nand U2854 (N_2854,N_2140,N_2225);
and U2855 (N_2855,N_2012,N_2023);
and U2856 (N_2856,N_1898,N_1757);
nand U2857 (N_2857,N_1730,N_1690);
nor U2858 (N_2858,N_2181,N_2010);
or U2859 (N_2859,N_2136,N_2202);
xnor U2860 (N_2860,N_1547,N_1545);
xnor U2861 (N_2861,N_2012,N_1623);
xnor U2862 (N_2862,N_2187,N_1522);
nand U2863 (N_2863,N_1677,N_1560);
nor U2864 (N_2864,N_1982,N_2126);
nor U2865 (N_2865,N_1798,N_1806);
nand U2866 (N_2866,N_1529,N_2232);
or U2867 (N_2867,N_1716,N_1683);
or U2868 (N_2868,N_1558,N_1997);
xor U2869 (N_2869,N_2022,N_1593);
nor U2870 (N_2870,N_1935,N_2181);
nand U2871 (N_2871,N_2162,N_1928);
nand U2872 (N_2872,N_1543,N_1888);
nand U2873 (N_2873,N_2244,N_1743);
nor U2874 (N_2874,N_2128,N_2041);
nand U2875 (N_2875,N_1730,N_1935);
and U2876 (N_2876,N_1939,N_2180);
xnor U2877 (N_2877,N_1940,N_1503);
nor U2878 (N_2878,N_1991,N_1956);
or U2879 (N_2879,N_1909,N_1989);
xor U2880 (N_2880,N_1648,N_2248);
xnor U2881 (N_2881,N_2205,N_2061);
xnor U2882 (N_2882,N_2111,N_1905);
and U2883 (N_2883,N_1595,N_2091);
nand U2884 (N_2884,N_1952,N_2119);
or U2885 (N_2885,N_2074,N_1990);
nand U2886 (N_2886,N_1534,N_2189);
xor U2887 (N_2887,N_2064,N_2218);
or U2888 (N_2888,N_1586,N_1706);
nor U2889 (N_2889,N_1533,N_2208);
nor U2890 (N_2890,N_2085,N_1683);
xnor U2891 (N_2891,N_2094,N_1689);
xor U2892 (N_2892,N_1864,N_1979);
nor U2893 (N_2893,N_2130,N_1646);
xnor U2894 (N_2894,N_2167,N_2084);
nand U2895 (N_2895,N_1695,N_1972);
nor U2896 (N_2896,N_1902,N_1982);
and U2897 (N_2897,N_2223,N_1599);
nor U2898 (N_2898,N_2168,N_1925);
or U2899 (N_2899,N_1556,N_1971);
nand U2900 (N_2900,N_2133,N_2095);
or U2901 (N_2901,N_1565,N_1964);
and U2902 (N_2902,N_1918,N_1558);
xnor U2903 (N_2903,N_2008,N_1873);
and U2904 (N_2904,N_1918,N_1816);
or U2905 (N_2905,N_2215,N_1865);
and U2906 (N_2906,N_1953,N_2044);
nand U2907 (N_2907,N_1541,N_1783);
xor U2908 (N_2908,N_2047,N_1700);
xnor U2909 (N_2909,N_1674,N_2179);
nand U2910 (N_2910,N_2117,N_1993);
and U2911 (N_2911,N_1861,N_2161);
xor U2912 (N_2912,N_2159,N_2075);
or U2913 (N_2913,N_1859,N_1760);
xor U2914 (N_2914,N_2112,N_2211);
and U2915 (N_2915,N_1942,N_1911);
and U2916 (N_2916,N_1741,N_1895);
or U2917 (N_2917,N_1862,N_1741);
or U2918 (N_2918,N_2069,N_2065);
and U2919 (N_2919,N_2102,N_1956);
or U2920 (N_2920,N_1547,N_2109);
xnor U2921 (N_2921,N_2110,N_1532);
xnor U2922 (N_2922,N_1510,N_2084);
or U2923 (N_2923,N_1539,N_1780);
nor U2924 (N_2924,N_1724,N_1949);
or U2925 (N_2925,N_1523,N_1944);
nor U2926 (N_2926,N_1654,N_2217);
or U2927 (N_2927,N_2140,N_2119);
nor U2928 (N_2928,N_1738,N_2070);
xnor U2929 (N_2929,N_1511,N_1637);
or U2930 (N_2930,N_1805,N_1848);
and U2931 (N_2931,N_1780,N_1830);
and U2932 (N_2932,N_2006,N_1698);
and U2933 (N_2933,N_1572,N_2017);
xnor U2934 (N_2934,N_1762,N_1941);
and U2935 (N_2935,N_1742,N_2131);
xor U2936 (N_2936,N_1658,N_1554);
and U2937 (N_2937,N_2077,N_2028);
nor U2938 (N_2938,N_1991,N_2207);
nand U2939 (N_2939,N_2227,N_2124);
nor U2940 (N_2940,N_1832,N_1764);
and U2941 (N_2941,N_2052,N_1895);
nor U2942 (N_2942,N_2218,N_1513);
and U2943 (N_2943,N_1838,N_1611);
nor U2944 (N_2944,N_1941,N_2001);
nor U2945 (N_2945,N_1828,N_2227);
nand U2946 (N_2946,N_2183,N_2083);
or U2947 (N_2947,N_2181,N_2196);
xnor U2948 (N_2948,N_1716,N_2158);
and U2949 (N_2949,N_2064,N_1984);
xor U2950 (N_2950,N_1672,N_2246);
and U2951 (N_2951,N_2009,N_2145);
and U2952 (N_2952,N_2135,N_1581);
or U2953 (N_2953,N_2148,N_2018);
and U2954 (N_2954,N_1700,N_2127);
nand U2955 (N_2955,N_1807,N_1826);
nand U2956 (N_2956,N_1500,N_1727);
xnor U2957 (N_2957,N_1540,N_2126);
nand U2958 (N_2958,N_1911,N_2147);
nand U2959 (N_2959,N_2135,N_2248);
or U2960 (N_2960,N_1961,N_1573);
or U2961 (N_2961,N_1728,N_1908);
nor U2962 (N_2962,N_1697,N_1589);
nand U2963 (N_2963,N_2122,N_1633);
nor U2964 (N_2964,N_1978,N_1851);
or U2965 (N_2965,N_2094,N_2009);
and U2966 (N_2966,N_1958,N_2180);
xor U2967 (N_2967,N_1509,N_1503);
xnor U2968 (N_2968,N_2240,N_1864);
xor U2969 (N_2969,N_2144,N_2202);
nor U2970 (N_2970,N_1892,N_1599);
xor U2971 (N_2971,N_2096,N_1737);
nor U2972 (N_2972,N_1909,N_2156);
and U2973 (N_2973,N_2247,N_1736);
xnor U2974 (N_2974,N_2091,N_1878);
and U2975 (N_2975,N_1773,N_1926);
or U2976 (N_2976,N_1634,N_1607);
nor U2977 (N_2977,N_2240,N_1595);
nand U2978 (N_2978,N_1809,N_1588);
xnor U2979 (N_2979,N_2004,N_1749);
nor U2980 (N_2980,N_1717,N_1695);
nand U2981 (N_2981,N_1927,N_2182);
nor U2982 (N_2982,N_2059,N_2169);
or U2983 (N_2983,N_2124,N_2118);
nor U2984 (N_2984,N_1971,N_1942);
nand U2985 (N_2985,N_1599,N_2157);
nor U2986 (N_2986,N_2197,N_2099);
nand U2987 (N_2987,N_1922,N_1983);
nand U2988 (N_2988,N_1941,N_1962);
or U2989 (N_2989,N_1569,N_2107);
and U2990 (N_2990,N_2235,N_1838);
nand U2991 (N_2991,N_1683,N_2077);
nor U2992 (N_2992,N_1871,N_1698);
and U2993 (N_2993,N_1723,N_1767);
or U2994 (N_2994,N_1926,N_1749);
and U2995 (N_2995,N_1524,N_1880);
xnor U2996 (N_2996,N_1594,N_2240);
or U2997 (N_2997,N_1964,N_1625);
nand U2998 (N_2998,N_1903,N_1766);
and U2999 (N_2999,N_2249,N_2007);
xnor UO_0 (O_0,N_2364,N_2502);
or UO_1 (O_1,N_2856,N_2619);
nor UO_2 (O_2,N_2984,N_2966);
and UO_3 (O_3,N_2718,N_2826);
and UO_4 (O_4,N_2373,N_2506);
xor UO_5 (O_5,N_2857,N_2492);
and UO_6 (O_6,N_2566,N_2746);
nor UO_7 (O_7,N_2845,N_2976);
and UO_8 (O_8,N_2766,N_2251);
xnor UO_9 (O_9,N_2963,N_2776);
nand UO_10 (O_10,N_2353,N_2460);
or UO_11 (O_11,N_2836,N_2275);
xnor UO_12 (O_12,N_2899,N_2866);
xnor UO_13 (O_13,N_2707,N_2729);
nand UO_14 (O_14,N_2303,N_2938);
nand UO_15 (O_15,N_2280,N_2659);
or UO_16 (O_16,N_2795,N_2980);
xnor UO_17 (O_17,N_2444,N_2310);
or UO_18 (O_18,N_2508,N_2287);
xor UO_19 (O_19,N_2309,N_2810);
xnor UO_20 (O_20,N_2332,N_2634);
nor UO_21 (O_21,N_2789,N_2904);
nand UO_22 (O_22,N_2575,N_2784);
and UO_23 (O_23,N_2390,N_2485);
nor UO_24 (O_24,N_2726,N_2289);
or UO_25 (O_25,N_2891,N_2643);
nand UO_26 (O_26,N_2898,N_2903);
and UO_27 (O_27,N_2633,N_2380);
nor UO_28 (O_28,N_2354,N_2305);
xor UO_29 (O_29,N_2312,N_2782);
xor UO_30 (O_30,N_2340,N_2816);
or UO_31 (O_31,N_2739,N_2604);
and UO_32 (O_32,N_2931,N_2421);
nor UO_33 (O_33,N_2438,N_2314);
and UO_34 (O_34,N_2467,N_2759);
nor UO_35 (O_35,N_2946,N_2284);
or UO_36 (O_36,N_2409,N_2468);
nand UO_37 (O_37,N_2547,N_2709);
and UO_38 (O_38,N_2551,N_2525);
and UO_39 (O_39,N_2655,N_2334);
nand UO_40 (O_40,N_2529,N_2840);
nor UO_41 (O_41,N_2626,N_2324);
xnor UO_42 (O_42,N_2939,N_2477);
or UO_43 (O_43,N_2417,N_2660);
xor UO_44 (O_44,N_2806,N_2777);
or UO_45 (O_45,N_2649,N_2620);
nand UO_46 (O_46,N_2997,N_2702);
nor UO_47 (O_47,N_2600,N_2863);
nand UO_48 (O_48,N_2694,N_2374);
nor UO_49 (O_49,N_2539,N_2657);
xnor UO_50 (O_50,N_2775,N_2809);
nor UO_51 (O_51,N_2935,N_2577);
nand UO_52 (O_52,N_2674,N_2763);
nand UO_53 (O_53,N_2791,N_2676);
nand UO_54 (O_54,N_2808,N_2268);
or UO_55 (O_55,N_2905,N_2347);
nor UO_56 (O_56,N_2503,N_2738);
nor UO_57 (O_57,N_2814,N_2326);
nor UO_58 (O_58,N_2977,N_2802);
and UO_59 (O_59,N_2741,N_2871);
xor UO_60 (O_60,N_2507,N_2951);
nor UO_61 (O_61,N_2489,N_2779);
xor UO_62 (O_62,N_2627,N_2682);
xor UO_63 (O_63,N_2786,N_2533);
nand UO_64 (O_64,N_2261,N_2953);
nand UO_65 (O_65,N_2257,N_2757);
nor UO_66 (O_66,N_2341,N_2900);
or UO_67 (O_67,N_2815,N_2865);
and UO_68 (O_68,N_2599,N_2988);
nand UO_69 (O_69,N_2753,N_2979);
nor UO_70 (O_70,N_2915,N_2668);
and UO_71 (O_71,N_2427,N_2523);
or UO_72 (O_72,N_2800,N_2567);
and UO_73 (O_73,N_2999,N_2839);
nor UO_74 (O_74,N_2949,N_2495);
or UO_75 (O_75,N_2990,N_2907);
xnor UO_76 (O_76,N_2527,N_2872);
nand UO_77 (O_77,N_2570,N_2748);
xnor UO_78 (O_78,N_2879,N_2259);
nand UO_79 (O_79,N_2638,N_2996);
or UO_80 (O_80,N_2365,N_2476);
nand UO_81 (O_81,N_2834,N_2440);
and UO_82 (O_82,N_2881,N_2419);
nor UO_83 (O_83,N_2631,N_2392);
xnor UO_84 (O_84,N_2315,N_2986);
xor UO_85 (O_85,N_2511,N_2725);
xor UO_86 (O_86,N_2798,N_2540);
nor UO_87 (O_87,N_2869,N_2370);
nand UO_88 (O_88,N_2496,N_2610);
xnor UO_89 (O_89,N_2947,N_2703);
or UO_90 (O_90,N_2393,N_2859);
nor UO_91 (O_91,N_2351,N_2338);
nor UO_92 (O_92,N_2811,N_2630);
nor UO_93 (O_93,N_2952,N_2394);
or UO_94 (O_94,N_2424,N_2428);
and UO_95 (O_95,N_2388,N_2743);
nand UO_96 (O_96,N_2520,N_2756);
or UO_97 (O_97,N_2618,N_2406);
nand UO_98 (O_98,N_2723,N_2677);
nand UO_99 (O_99,N_2958,N_2528);
and UO_100 (O_100,N_2475,N_2956);
xor UO_101 (O_101,N_2835,N_2851);
xor UO_102 (O_102,N_2458,N_2778);
nor UO_103 (O_103,N_2629,N_2480);
or UO_104 (O_104,N_2501,N_2942);
nor UO_105 (O_105,N_2472,N_2654);
nand UO_106 (O_106,N_2552,N_2342);
and UO_107 (O_107,N_2293,N_2889);
nand UO_108 (O_108,N_2422,N_2514);
nor UO_109 (O_109,N_2328,N_2787);
or UO_110 (O_110,N_2329,N_2945);
and UO_111 (O_111,N_2862,N_2363);
and UO_112 (O_112,N_2758,N_2425);
nor UO_113 (O_113,N_2932,N_2437);
xnor UO_114 (O_114,N_2269,N_2505);
xor UO_115 (O_115,N_2396,N_2369);
nand UO_116 (O_116,N_2955,N_2608);
and UO_117 (O_117,N_2372,N_2561);
nand UO_118 (O_118,N_2436,N_2876);
nor UO_119 (O_119,N_2559,N_2598);
and UO_120 (O_120,N_2727,N_2691);
xor UO_121 (O_121,N_2482,N_2488);
and UO_122 (O_122,N_2543,N_2300);
xnor UO_123 (O_123,N_2715,N_2362);
xnor UO_124 (O_124,N_2637,N_2262);
and UO_125 (O_125,N_2833,N_2724);
and UO_126 (O_126,N_2770,N_2441);
nand UO_127 (O_127,N_2658,N_2882);
nand UO_128 (O_128,N_2473,N_2957);
nand UO_129 (O_129,N_2978,N_2418);
nand UO_130 (O_130,N_2639,N_2398);
xnor UO_131 (O_131,N_2673,N_2717);
xnor UO_132 (O_132,N_2645,N_2337);
nand UO_133 (O_133,N_2500,N_2302);
nand UO_134 (O_134,N_2678,N_2581);
nand UO_135 (O_135,N_2565,N_2360);
and UO_136 (O_136,N_2968,N_2930);
or UO_137 (O_137,N_2410,N_2737);
or UO_138 (O_138,N_2812,N_2260);
xnor UO_139 (O_139,N_2531,N_2716);
nor UO_140 (O_140,N_2982,N_2896);
nand UO_141 (O_141,N_2288,N_2319);
or UO_142 (O_142,N_2925,N_2647);
nor UO_143 (O_143,N_2317,N_2359);
nand UO_144 (O_144,N_2974,N_2278);
nor UO_145 (O_145,N_2803,N_2587);
or UO_146 (O_146,N_2585,N_2959);
or UO_147 (O_147,N_2885,N_2731);
nor UO_148 (O_148,N_2550,N_2254);
or UO_149 (O_149,N_2744,N_2923);
and UO_150 (O_150,N_2431,N_2415);
and UO_151 (O_151,N_2271,N_2653);
and UO_152 (O_152,N_2623,N_2728);
nor UO_153 (O_153,N_2367,N_2940);
or UO_154 (O_154,N_2336,N_2447);
or UO_155 (O_155,N_2936,N_2345);
or UO_156 (O_156,N_2563,N_2250);
nor UO_157 (O_157,N_2265,N_2686);
or UO_158 (O_158,N_2446,N_2343);
and UO_159 (O_159,N_2594,N_2695);
nand UO_160 (O_160,N_2252,N_2771);
nand UO_161 (O_161,N_2868,N_2995);
nor UO_162 (O_162,N_2920,N_2895);
nand UO_163 (O_163,N_2697,N_2435);
xnor UO_164 (O_164,N_2961,N_2267);
or UO_165 (O_165,N_2730,N_2586);
and UO_166 (O_166,N_2632,N_2366);
or UO_167 (O_167,N_2909,N_2858);
or UO_168 (O_168,N_2813,N_2413);
nor UO_169 (O_169,N_2376,N_2384);
and UO_170 (O_170,N_2964,N_2576);
nor UO_171 (O_171,N_2847,N_2555);
nand UO_172 (O_172,N_2368,N_2679);
and UO_173 (O_173,N_2513,N_2442);
nor UO_174 (O_174,N_2675,N_2589);
and UO_175 (O_175,N_2998,N_2687);
xnor UO_176 (O_176,N_2377,N_2464);
or UO_177 (O_177,N_2644,N_2642);
xnor UO_178 (O_178,N_2283,N_2263);
xor UO_179 (O_179,N_2348,N_2453);
xor UO_180 (O_180,N_2621,N_2516);
xor UO_181 (O_181,N_2823,N_2509);
xor UO_182 (O_182,N_2625,N_2320);
xnor UO_183 (O_183,N_2486,N_2892);
xnor UO_184 (O_184,N_2785,N_2297);
or UO_185 (O_185,N_2706,N_2937);
nor UO_186 (O_186,N_2451,N_2841);
nor UO_187 (O_187,N_2306,N_2830);
and UO_188 (O_188,N_2426,N_2828);
and UO_189 (O_189,N_2635,N_2713);
nor UO_190 (O_190,N_2965,N_2433);
nand UO_191 (O_191,N_2596,N_2296);
xnor UO_192 (O_192,N_2805,N_2407);
nor UO_193 (O_193,N_2666,N_2875);
nor UO_194 (O_194,N_2454,N_2801);
or UO_195 (O_195,N_2684,N_2878);
xnor UO_196 (O_196,N_2960,N_2403);
xor UO_197 (O_197,N_2807,N_2975);
and UO_198 (O_198,N_2754,N_2860);
nor UO_199 (O_199,N_2535,N_2579);
and UO_200 (O_200,N_2378,N_2688);
nor UO_201 (O_201,N_2667,N_2591);
xnor UO_202 (O_202,N_2669,N_2499);
nor UO_203 (O_203,N_2944,N_2661);
and UO_204 (O_204,N_2530,N_2652);
or UO_205 (O_205,N_2412,N_2479);
nand UO_206 (O_206,N_2361,N_2641);
xnor UO_207 (O_207,N_2783,N_2358);
nand UO_208 (O_208,N_2294,N_2843);
or UO_209 (O_209,N_2542,N_2408);
and UO_210 (O_210,N_2416,N_2853);
or UO_211 (O_211,N_2818,N_2462);
and UO_212 (O_212,N_2870,N_2640);
or UO_213 (O_213,N_2656,N_2804);
xnor UO_214 (O_214,N_2922,N_2749);
or UO_215 (O_215,N_2449,N_2928);
nand UO_216 (O_216,N_2967,N_2616);
xor UO_217 (O_217,N_2933,N_2512);
or UO_218 (O_218,N_2689,N_2556);
and UO_219 (O_219,N_2609,N_2912);
nand UO_220 (O_220,N_2734,N_2430);
xnor UO_221 (O_221,N_2582,N_2750);
nand UO_222 (O_222,N_2612,N_2402);
nand UO_223 (O_223,N_2295,N_2651);
nor UO_224 (O_224,N_2762,N_2434);
nor UO_225 (O_225,N_2597,N_2711);
or UO_226 (O_226,N_2256,N_2515);
nand UO_227 (O_227,N_2395,N_2973);
xor UO_228 (O_228,N_2852,N_2710);
nor UO_229 (O_229,N_2544,N_2327);
and UO_230 (O_230,N_2821,N_2397);
nand UO_231 (O_231,N_2494,N_2824);
or UO_232 (O_232,N_2751,N_2712);
or UO_233 (O_233,N_2487,N_2483);
or UO_234 (O_234,N_2258,N_2588);
nand UO_235 (O_235,N_2375,N_2767);
and UO_236 (O_236,N_2736,N_2569);
nor UO_237 (O_237,N_2423,N_2827);
xnor UO_238 (O_238,N_2918,N_2672);
xor UO_239 (O_239,N_2574,N_2613);
xor UO_240 (O_240,N_2848,N_2831);
xor UO_241 (O_241,N_2281,N_2429);
xor UO_242 (O_242,N_2481,N_2298);
nor UO_243 (O_243,N_2333,N_2573);
nor UO_244 (O_244,N_2273,N_2985);
and UO_245 (O_245,N_2850,N_2386);
nor UO_246 (O_246,N_2548,N_2465);
and UO_247 (O_247,N_2617,N_2680);
xnor UO_248 (O_248,N_2941,N_2989);
xnor UO_249 (O_249,N_2471,N_2264);
and UO_250 (O_250,N_2253,N_2391);
nand UO_251 (O_251,N_2636,N_2304);
nand UO_252 (O_252,N_2322,N_2714);
xor UO_253 (O_253,N_2571,N_2411);
nand UO_254 (O_254,N_2740,N_2906);
or UO_255 (O_255,N_2755,N_2606);
nand UO_256 (O_256,N_2450,N_2796);
nor UO_257 (O_257,N_2765,N_2330);
and UO_258 (O_258,N_2484,N_2291);
nor UO_259 (O_259,N_2615,N_2286);
nor UO_260 (O_260,N_2292,N_2972);
nor UO_261 (O_261,N_2719,N_2704);
or UO_262 (O_262,N_2399,N_2558);
and UO_263 (O_263,N_2735,N_2352);
and UO_264 (O_264,N_2914,N_2873);
or UO_265 (O_265,N_2646,N_2628);
nand UO_266 (O_266,N_2837,N_2318);
xor UO_267 (O_267,N_2768,N_2401);
nor UO_268 (O_268,N_2562,N_2389);
or UO_269 (O_269,N_2901,N_2781);
xnor UO_270 (O_270,N_2877,N_2720);
xor UO_271 (O_271,N_2276,N_2919);
nand UO_272 (O_272,N_2705,N_2902);
or UO_273 (O_273,N_2607,N_2498);
or UO_274 (O_274,N_2538,N_2557);
nand UO_275 (O_275,N_2560,N_2325);
nand UO_276 (O_276,N_2690,N_2916);
nor UO_277 (O_277,N_2553,N_2510);
and UO_278 (O_278,N_2708,N_2886);
or UO_279 (O_279,N_2722,N_2760);
nor UO_280 (O_280,N_2272,N_2917);
xnor UO_281 (O_281,N_2456,N_2478);
nor UO_282 (O_282,N_2432,N_2908);
nand UO_283 (O_283,N_2316,N_2578);
xnor UO_284 (O_284,N_2534,N_2355);
nor UO_285 (O_285,N_2545,N_2832);
nor UO_286 (O_286,N_2983,N_2371);
nand UO_287 (O_287,N_2842,N_2470);
xnor UO_288 (O_288,N_2405,N_2455);
nand UO_289 (O_289,N_2681,N_2913);
and UO_290 (O_290,N_2971,N_2466);
nor UO_291 (O_291,N_2864,N_2624);
xnor UO_292 (O_292,N_2614,N_2890);
nor UO_293 (O_293,N_2400,N_2954);
nor UO_294 (O_294,N_2910,N_2443);
and UO_295 (O_295,N_2874,N_2993);
and UO_296 (O_296,N_2752,N_2692);
nand UO_297 (O_297,N_2897,N_2474);
nor UO_298 (O_298,N_2339,N_2349);
xnor UO_299 (O_299,N_2817,N_2825);
and UO_300 (O_300,N_2350,N_2323);
xor UO_301 (O_301,N_2445,N_2546);
nor UO_302 (O_302,N_2346,N_2670);
nand UO_303 (O_303,N_2927,N_2279);
xor UO_304 (O_304,N_2622,N_2452);
nor UO_305 (O_305,N_2780,N_2650);
xnor UO_306 (O_306,N_2987,N_2448);
xnor UO_307 (O_307,N_2537,N_2700);
nand UO_308 (O_308,N_2457,N_2950);
and UO_309 (O_309,N_2344,N_2794);
nand UO_310 (O_310,N_2934,N_2601);
nor UO_311 (O_311,N_2526,N_2469);
or UO_312 (O_312,N_2356,N_2603);
xnor UO_313 (O_313,N_2820,N_2266);
nor UO_314 (O_314,N_2962,N_2549);
xnor UO_315 (O_315,N_2911,N_2519);
or UO_316 (O_316,N_2788,N_2335);
or UO_317 (O_317,N_2490,N_2383);
nand UO_318 (O_318,N_2829,N_2924);
nor UO_319 (O_319,N_2887,N_2721);
or UO_320 (O_320,N_2459,N_2255);
nand UO_321 (O_321,N_2307,N_2867);
xnor UO_322 (O_322,N_2844,N_2521);
nand UO_323 (O_323,N_2381,N_2991);
nand UO_324 (O_324,N_2792,N_2693);
nor UO_325 (O_325,N_2308,N_2894);
nand UO_326 (O_326,N_2994,N_2313);
xor UO_327 (O_327,N_2948,N_2772);
or UO_328 (O_328,N_2282,N_2592);
xnor UO_329 (O_329,N_2285,N_2532);
xor UO_330 (O_330,N_2884,N_2854);
nand UO_331 (O_331,N_2970,N_2439);
nand UO_332 (O_332,N_2568,N_2888);
or UO_333 (O_333,N_2517,N_2745);
nor UO_334 (O_334,N_2969,N_2536);
xnor UO_335 (O_335,N_2819,N_2699);
nand UO_336 (O_336,N_2926,N_2733);
xor UO_337 (O_337,N_2270,N_2420);
nor UO_338 (O_338,N_2404,N_2883);
and UO_339 (O_339,N_2611,N_2732);
or UO_340 (O_340,N_2929,N_2921);
or UO_341 (O_341,N_2769,N_2671);
or UO_342 (O_342,N_2493,N_2290);
nor UO_343 (O_343,N_2522,N_2605);
and UO_344 (O_344,N_2855,N_2698);
nor UO_345 (O_345,N_2822,N_2379);
or UO_346 (O_346,N_2665,N_2701);
xnor UO_347 (O_347,N_2880,N_2747);
and UO_348 (O_348,N_2584,N_2663);
nand UO_349 (O_349,N_2463,N_2838);
xor UO_350 (O_350,N_2943,N_2764);
and UO_351 (O_351,N_2662,N_2590);
and UO_352 (O_352,N_2331,N_2277);
and UO_353 (O_353,N_2799,N_2761);
nand UO_354 (O_354,N_2491,N_2861);
nor UO_355 (O_355,N_2648,N_2518);
or UO_356 (O_356,N_2846,N_2564);
or UO_357 (O_357,N_2299,N_2696);
and UO_358 (O_358,N_2773,N_2593);
nand UO_359 (O_359,N_2382,N_2385);
nand UO_360 (O_360,N_2583,N_2414);
nand UO_361 (O_361,N_2595,N_2554);
nor UO_362 (O_362,N_2602,N_2664);
xnor UO_363 (O_363,N_2541,N_2742);
nand UO_364 (O_364,N_2524,N_2387);
or UO_365 (O_365,N_2357,N_2797);
xor UO_366 (O_366,N_2580,N_2992);
nor UO_367 (O_367,N_2461,N_2793);
xor UO_368 (O_368,N_2504,N_2683);
and UO_369 (O_369,N_2301,N_2981);
nor UO_370 (O_370,N_2790,N_2311);
nand UO_371 (O_371,N_2274,N_2849);
and UO_372 (O_372,N_2685,N_2321);
and UO_373 (O_373,N_2893,N_2774);
nor UO_374 (O_374,N_2497,N_2572);
or UO_375 (O_375,N_2391,N_2337);
and UO_376 (O_376,N_2317,N_2438);
nand UO_377 (O_377,N_2297,N_2760);
xor UO_378 (O_378,N_2378,N_2374);
xor UO_379 (O_379,N_2639,N_2292);
xor UO_380 (O_380,N_2646,N_2562);
and UO_381 (O_381,N_2560,N_2938);
or UO_382 (O_382,N_2758,N_2323);
nor UO_383 (O_383,N_2704,N_2429);
nor UO_384 (O_384,N_2320,N_2480);
nor UO_385 (O_385,N_2602,N_2414);
xor UO_386 (O_386,N_2436,N_2552);
or UO_387 (O_387,N_2324,N_2853);
and UO_388 (O_388,N_2604,N_2312);
xor UO_389 (O_389,N_2632,N_2992);
or UO_390 (O_390,N_2374,N_2498);
xor UO_391 (O_391,N_2628,N_2490);
or UO_392 (O_392,N_2734,N_2658);
xnor UO_393 (O_393,N_2330,N_2919);
or UO_394 (O_394,N_2301,N_2282);
nand UO_395 (O_395,N_2877,N_2908);
nor UO_396 (O_396,N_2664,N_2561);
xnor UO_397 (O_397,N_2436,N_2316);
or UO_398 (O_398,N_2862,N_2730);
or UO_399 (O_399,N_2744,N_2410);
nor UO_400 (O_400,N_2575,N_2565);
nor UO_401 (O_401,N_2571,N_2996);
or UO_402 (O_402,N_2412,N_2275);
and UO_403 (O_403,N_2286,N_2552);
nand UO_404 (O_404,N_2615,N_2362);
nor UO_405 (O_405,N_2636,N_2598);
xor UO_406 (O_406,N_2263,N_2676);
nand UO_407 (O_407,N_2754,N_2374);
nand UO_408 (O_408,N_2441,N_2864);
xnor UO_409 (O_409,N_2816,N_2550);
nand UO_410 (O_410,N_2869,N_2734);
or UO_411 (O_411,N_2629,N_2587);
or UO_412 (O_412,N_2321,N_2368);
xnor UO_413 (O_413,N_2627,N_2283);
nor UO_414 (O_414,N_2361,N_2395);
xnor UO_415 (O_415,N_2933,N_2300);
or UO_416 (O_416,N_2476,N_2251);
and UO_417 (O_417,N_2366,N_2840);
xor UO_418 (O_418,N_2797,N_2956);
and UO_419 (O_419,N_2502,N_2555);
or UO_420 (O_420,N_2460,N_2885);
nand UO_421 (O_421,N_2537,N_2448);
or UO_422 (O_422,N_2814,N_2885);
xor UO_423 (O_423,N_2578,N_2370);
or UO_424 (O_424,N_2412,N_2635);
and UO_425 (O_425,N_2348,N_2286);
and UO_426 (O_426,N_2427,N_2876);
and UO_427 (O_427,N_2462,N_2613);
or UO_428 (O_428,N_2399,N_2897);
xnor UO_429 (O_429,N_2500,N_2491);
xor UO_430 (O_430,N_2337,N_2903);
or UO_431 (O_431,N_2361,N_2995);
or UO_432 (O_432,N_2677,N_2534);
and UO_433 (O_433,N_2457,N_2371);
or UO_434 (O_434,N_2983,N_2595);
xnor UO_435 (O_435,N_2641,N_2408);
nor UO_436 (O_436,N_2932,N_2985);
and UO_437 (O_437,N_2657,N_2429);
nand UO_438 (O_438,N_2705,N_2566);
and UO_439 (O_439,N_2496,N_2639);
or UO_440 (O_440,N_2275,N_2905);
or UO_441 (O_441,N_2499,N_2952);
nand UO_442 (O_442,N_2361,N_2801);
xor UO_443 (O_443,N_2650,N_2435);
and UO_444 (O_444,N_2412,N_2391);
nand UO_445 (O_445,N_2535,N_2540);
xor UO_446 (O_446,N_2447,N_2821);
nor UO_447 (O_447,N_2988,N_2252);
nor UO_448 (O_448,N_2831,N_2959);
nand UO_449 (O_449,N_2877,N_2579);
nand UO_450 (O_450,N_2460,N_2769);
nor UO_451 (O_451,N_2883,N_2465);
nor UO_452 (O_452,N_2749,N_2981);
nor UO_453 (O_453,N_2577,N_2417);
nor UO_454 (O_454,N_2994,N_2493);
or UO_455 (O_455,N_2763,N_2250);
nand UO_456 (O_456,N_2291,N_2457);
and UO_457 (O_457,N_2831,N_2513);
xnor UO_458 (O_458,N_2373,N_2362);
or UO_459 (O_459,N_2565,N_2620);
and UO_460 (O_460,N_2579,N_2684);
nand UO_461 (O_461,N_2924,N_2939);
xnor UO_462 (O_462,N_2850,N_2668);
nand UO_463 (O_463,N_2265,N_2737);
or UO_464 (O_464,N_2668,N_2667);
nor UO_465 (O_465,N_2555,N_2643);
or UO_466 (O_466,N_2472,N_2931);
xor UO_467 (O_467,N_2683,N_2456);
xor UO_468 (O_468,N_2874,N_2914);
or UO_469 (O_469,N_2482,N_2476);
and UO_470 (O_470,N_2838,N_2692);
xor UO_471 (O_471,N_2889,N_2671);
nand UO_472 (O_472,N_2891,N_2501);
and UO_473 (O_473,N_2518,N_2905);
and UO_474 (O_474,N_2574,N_2659);
and UO_475 (O_475,N_2311,N_2983);
nor UO_476 (O_476,N_2404,N_2303);
and UO_477 (O_477,N_2699,N_2491);
and UO_478 (O_478,N_2776,N_2901);
nor UO_479 (O_479,N_2423,N_2782);
xor UO_480 (O_480,N_2252,N_2626);
or UO_481 (O_481,N_2645,N_2342);
and UO_482 (O_482,N_2526,N_2854);
or UO_483 (O_483,N_2656,N_2683);
or UO_484 (O_484,N_2958,N_2596);
and UO_485 (O_485,N_2447,N_2719);
and UO_486 (O_486,N_2700,N_2876);
or UO_487 (O_487,N_2769,N_2981);
xnor UO_488 (O_488,N_2886,N_2413);
xnor UO_489 (O_489,N_2832,N_2613);
xnor UO_490 (O_490,N_2343,N_2252);
nand UO_491 (O_491,N_2889,N_2591);
nor UO_492 (O_492,N_2888,N_2485);
xor UO_493 (O_493,N_2289,N_2784);
and UO_494 (O_494,N_2770,N_2899);
or UO_495 (O_495,N_2346,N_2713);
nor UO_496 (O_496,N_2910,N_2590);
xor UO_497 (O_497,N_2789,N_2275);
nand UO_498 (O_498,N_2440,N_2942);
and UO_499 (O_499,N_2922,N_2581);
endmodule