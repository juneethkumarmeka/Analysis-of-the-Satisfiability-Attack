module basic_500_3000_500_6_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_472,In_225);
or U1 (N_1,In_155,In_279);
and U2 (N_2,In_42,In_131);
and U3 (N_3,In_83,In_118);
and U4 (N_4,In_398,In_369);
and U5 (N_5,In_420,In_257);
nand U6 (N_6,In_374,In_50);
nor U7 (N_7,In_482,In_382);
or U8 (N_8,In_18,In_254);
or U9 (N_9,In_97,In_253);
nand U10 (N_10,In_82,In_370);
and U11 (N_11,In_256,In_128);
nor U12 (N_12,In_192,In_477);
nor U13 (N_13,In_443,In_229);
or U14 (N_14,In_232,In_452);
nand U15 (N_15,In_153,In_189);
nor U16 (N_16,In_412,In_204);
or U17 (N_17,In_179,In_22);
and U18 (N_18,In_246,In_379);
nor U19 (N_19,In_133,In_381);
nand U20 (N_20,In_483,In_223);
and U21 (N_21,In_292,In_162);
or U22 (N_22,In_116,In_315);
and U23 (N_23,In_307,In_212);
or U24 (N_24,In_180,In_245);
and U25 (N_25,In_270,In_260);
or U26 (N_26,In_49,In_235);
nand U27 (N_27,In_394,In_144);
nor U28 (N_28,In_213,In_274);
nand U29 (N_29,In_309,In_161);
xor U30 (N_30,In_69,In_15);
or U31 (N_31,In_182,In_322);
or U32 (N_32,In_29,In_347);
nor U33 (N_33,In_132,In_284);
or U34 (N_34,In_291,In_303);
nand U35 (N_35,In_54,In_39);
nor U36 (N_36,In_485,In_259);
and U37 (N_37,In_159,In_311);
or U38 (N_38,In_173,In_198);
nor U39 (N_39,In_368,In_160);
and U40 (N_40,In_334,In_419);
or U41 (N_41,In_226,In_336);
nand U42 (N_42,In_111,In_436);
nand U43 (N_43,In_194,In_267);
or U44 (N_44,In_312,In_397);
and U45 (N_45,In_172,In_393);
nor U46 (N_46,In_202,In_211);
nor U47 (N_47,In_104,In_154);
nand U48 (N_48,In_59,In_114);
or U49 (N_49,In_283,In_359);
nand U50 (N_50,In_31,In_142);
or U51 (N_51,In_310,In_70);
or U52 (N_52,In_422,In_352);
nor U53 (N_53,In_484,In_112);
nand U54 (N_54,In_72,In_2);
and U55 (N_55,In_20,In_134);
or U56 (N_56,In_209,In_439);
and U57 (N_57,In_300,In_187);
or U58 (N_58,In_366,In_158);
nor U59 (N_59,In_288,In_169);
or U60 (N_60,In_333,In_199);
nor U61 (N_61,In_152,In_375);
or U62 (N_62,In_13,In_215);
and U63 (N_63,In_9,In_136);
nand U64 (N_64,In_289,In_120);
or U65 (N_65,In_197,In_34);
and U66 (N_66,In_490,In_98);
xor U67 (N_67,In_335,In_447);
nand U68 (N_68,In_200,In_430);
or U69 (N_69,In_88,In_266);
nand U70 (N_70,In_344,In_105);
or U71 (N_71,In_247,In_65);
and U72 (N_72,In_250,In_305);
nand U73 (N_73,In_489,In_421);
nor U74 (N_74,In_217,In_26);
or U75 (N_75,In_101,In_32);
nor U76 (N_76,In_499,In_295);
nor U77 (N_77,In_3,In_342);
and U78 (N_78,In_220,In_40);
nand U79 (N_79,In_61,In_92);
nor U80 (N_80,In_328,In_361);
or U81 (N_81,In_349,In_383);
or U82 (N_82,In_5,In_73);
or U83 (N_83,In_207,In_411);
and U84 (N_84,In_406,In_285);
or U85 (N_85,In_353,In_167);
nand U86 (N_86,In_45,In_319);
and U87 (N_87,In_302,In_265);
nor U88 (N_88,In_377,In_468);
or U89 (N_89,In_221,In_362);
or U90 (N_90,In_455,In_330);
xor U91 (N_91,In_478,In_273);
or U92 (N_92,In_338,In_389);
and U93 (N_93,In_448,In_86);
nor U94 (N_94,In_316,In_299);
or U95 (N_95,In_364,In_437);
or U96 (N_96,In_214,In_135);
nor U97 (N_97,In_405,In_454);
and U98 (N_98,In_294,In_23);
nand U99 (N_99,In_208,In_297);
nand U100 (N_100,In_296,In_44);
nand U101 (N_101,In_280,In_261);
and U102 (N_102,In_216,In_277);
or U103 (N_103,In_282,In_47);
nand U104 (N_104,In_143,In_323);
nor U105 (N_105,In_473,In_456);
or U106 (N_106,In_355,In_122);
and U107 (N_107,In_409,In_176);
nor U108 (N_108,In_440,In_290);
or U109 (N_109,In_170,In_41);
nor U110 (N_110,In_264,In_96);
nor U111 (N_111,In_298,In_175);
nor U112 (N_112,In_475,In_51);
and U113 (N_113,In_391,In_164);
or U114 (N_114,In_35,In_137);
nand U115 (N_115,In_237,In_228);
nand U116 (N_116,In_460,In_196);
nor U117 (N_117,In_354,In_317);
and U118 (N_118,In_0,In_206);
and U119 (N_119,In_166,In_387);
nand U120 (N_120,In_465,In_56);
and U121 (N_121,In_190,In_320);
or U122 (N_122,In_392,In_76);
and U123 (N_123,In_481,In_8);
nand U124 (N_124,In_373,In_269);
nor U125 (N_125,In_149,In_174);
or U126 (N_126,In_62,In_314);
and U127 (N_127,In_81,In_399);
or U128 (N_128,In_231,In_21);
nand U129 (N_129,In_145,In_24);
and U130 (N_130,In_219,In_242);
nand U131 (N_131,In_445,In_474);
nand U132 (N_132,In_90,In_400);
nand U133 (N_133,In_453,In_402);
or U134 (N_134,In_123,In_146);
nor U135 (N_135,In_60,In_195);
or U136 (N_136,In_433,In_110);
and U137 (N_137,In_331,In_230);
and U138 (N_138,In_345,In_469);
or U139 (N_139,In_441,In_327);
nand U140 (N_140,In_360,In_156);
nor U141 (N_141,In_203,In_129);
nor U142 (N_142,In_11,In_466);
nand U143 (N_143,In_497,In_415);
and U144 (N_144,In_95,In_488);
or U145 (N_145,In_376,In_102);
nor U146 (N_146,In_262,In_446);
nor U147 (N_147,In_495,In_163);
nand U148 (N_148,In_94,In_459);
nor U149 (N_149,In_413,In_240);
or U150 (N_150,In_462,In_363);
or U151 (N_151,In_30,In_125);
nand U152 (N_152,In_340,In_151);
nand U153 (N_153,In_395,In_67);
nor U154 (N_154,In_332,In_470);
nor U155 (N_155,In_358,In_263);
nand U156 (N_156,In_463,In_74);
and U157 (N_157,In_386,In_367);
nand U158 (N_158,In_432,In_341);
nor U159 (N_159,In_286,In_66);
nand U160 (N_160,In_486,In_52);
or U161 (N_161,In_181,In_165);
and U162 (N_162,In_404,In_416);
xnor U163 (N_163,In_390,In_168);
nor U164 (N_164,In_434,In_58);
nor U165 (N_165,In_321,In_25);
nand U166 (N_166,In_14,In_479);
or U167 (N_167,In_318,In_238);
nand U168 (N_168,In_147,In_278);
nor U169 (N_169,In_7,In_449);
nor U170 (N_170,In_185,In_201);
nor U171 (N_171,In_6,In_494);
nor U172 (N_172,In_178,In_304);
nand U173 (N_173,In_244,In_343);
nand U174 (N_174,In_268,In_329);
nand U175 (N_175,In_464,In_275);
or U176 (N_176,In_19,In_27);
and U177 (N_177,In_301,In_138);
and U178 (N_178,In_141,In_458);
or U179 (N_179,In_222,In_414);
nor U180 (N_180,In_372,In_293);
nor U181 (N_181,In_384,In_426);
and U182 (N_182,In_348,In_193);
or U183 (N_183,In_79,In_276);
nand U184 (N_184,In_281,In_80);
nand U185 (N_185,In_385,In_117);
and U186 (N_186,In_55,In_325);
nand U187 (N_187,In_423,In_106);
nand U188 (N_188,In_427,In_43);
or U189 (N_189,In_77,In_17);
or U190 (N_190,In_444,In_467);
or U191 (N_191,In_127,In_417);
or U192 (N_192,In_357,In_487);
or U193 (N_193,In_139,In_157);
or U194 (N_194,In_126,In_255);
or U195 (N_195,In_272,In_403);
and U196 (N_196,In_183,In_150);
or U197 (N_197,In_442,In_46);
and U198 (N_198,In_100,In_356);
or U199 (N_199,In_130,In_140);
and U200 (N_200,In_401,In_480);
and U201 (N_201,In_93,In_287);
nor U202 (N_202,In_224,In_103);
or U203 (N_203,In_99,In_57);
nand U204 (N_204,In_451,In_498);
nand U205 (N_205,In_418,In_84);
nor U206 (N_206,In_53,In_12);
nor U207 (N_207,In_113,In_471);
or U208 (N_208,In_124,In_68);
nor U209 (N_209,In_408,In_431);
or U210 (N_210,In_258,In_236);
or U211 (N_211,In_78,In_4);
and U212 (N_212,In_239,In_271);
or U213 (N_213,In_380,In_324);
and U214 (N_214,In_365,In_191);
and U215 (N_215,In_33,In_493);
or U216 (N_216,In_91,In_85);
and U217 (N_217,In_119,In_308);
nor U218 (N_218,In_410,In_346);
or U219 (N_219,In_28,In_71);
or U220 (N_220,In_371,In_457);
nand U221 (N_221,In_435,In_249);
and U222 (N_222,In_337,In_115);
or U223 (N_223,In_107,In_496);
or U224 (N_224,In_248,In_461);
nand U225 (N_225,In_177,In_227);
nor U226 (N_226,In_407,In_424);
and U227 (N_227,In_252,In_184);
xnor U228 (N_228,In_148,In_251);
nor U229 (N_229,In_63,In_339);
nor U230 (N_230,In_313,In_241);
nand U231 (N_231,In_491,In_428);
and U232 (N_232,In_234,In_476);
or U233 (N_233,In_186,In_10);
nand U234 (N_234,In_87,In_425);
or U235 (N_235,In_109,In_171);
and U236 (N_236,In_48,In_210);
nand U237 (N_237,In_450,In_36);
nand U238 (N_238,In_306,In_388);
nand U239 (N_239,In_218,In_16);
nor U240 (N_240,In_378,In_429);
nor U241 (N_241,In_326,In_188);
and U242 (N_242,In_121,In_108);
or U243 (N_243,In_37,In_75);
nand U244 (N_244,In_350,In_38);
nor U245 (N_245,In_89,In_233);
or U246 (N_246,In_492,In_351);
or U247 (N_247,In_1,In_438);
nor U248 (N_248,In_243,In_205);
nor U249 (N_249,In_64,In_396);
nand U250 (N_250,In_23,In_201);
nand U251 (N_251,In_409,In_256);
nor U252 (N_252,In_396,In_372);
nor U253 (N_253,In_142,In_221);
and U254 (N_254,In_338,In_477);
and U255 (N_255,In_461,In_118);
nor U256 (N_256,In_499,In_164);
or U257 (N_257,In_44,In_347);
or U258 (N_258,In_100,In_184);
or U259 (N_259,In_203,In_294);
nor U260 (N_260,In_179,In_398);
and U261 (N_261,In_164,In_261);
nand U262 (N_262,In_337,In_48);
nor U263 (N_263,In_133,In_376);
and U264 (N_264,In_255,In_47);
and U265 (N_265,In_25,In_48);
and U266 (N_266,In_326,In_97);
nor U267 (N_267,In_185,In_259);
or U268 (N_268,In_165,In_241);
nand U269 (N_269,In_234,In_498);
and U270 (N_270,In_470,In_347);
nand U271 (N_271,In_219,In_353);
nand U272 (N_272,In_430,In_310);
and U273 (N_273,In_47,In_495);
and U274 (N_274,In_353,In_115);
or U275 (N_275,In_261,In_272);
or U276 (N_276,In_217,In_317);
nand U277 (N_277,In_386,In_138);
or U278 (N_278,In_81,In_193);
or U279 (N_279,In_432,In_268);
and U280 (N_280,In_332,In_230);
or U281 (N_281,In_11,In_145);
nand U282 (N_282,In_237,In_409);
and U283 (N_283,In_253,In_70);
nand U284 (N_284,In_174,In_186);
or U285 (N_285,In_240,In_269);
or U286 (N_286,In_164,In_283);
and U287 (N_287,In_216,In_74);
nor U288 (N_288,In_7,In_10);
nand U289 (N_289,In_209,In_66);
or U290 (N_290,In_46,In_26);
and U291 (N_291,In_19,In_421);
and U292 (N_292,In_287,In_331);
or U293 (N_293,In_244,In_408);
nand U294 (N_294,In_13,In_168);
nand U295 (N_295,In_59,In_57);
nor U296 (N_296,In_109,In_151);
and U297 (N_297,In_100,In_448);
or U298 (N_298,In_175,In_12);
nor U299 (N_299,In_344,In_375);
nor U300 (N_300,In_68,In_443);
nor U301 (N_301,In_471,In_445);
nand U302 (N_302,In_217,In_336);
nand U303 (N_303,In_87,In_411);
nor U304 (N_304,In_153,In_141);
nor U305 (N_305,In_198,In_207);
or U306 (N_306,In_381,In_219);
or U307 (N_307,In_219,In_351);
nand U308 (N_308,In_365,In_489);
nor U309 (N_309,In_12,In_259);
xor U310 (N_310,In_249,In_21);
nand U311 (N_311,In_458,In_157);
and U312 (N_312,In_485,In_56);
and U313 (N_313,In_73,In_234);
or U314 (N_314,In_202,In_444);
nor U315 (N_315,In_53,In_144);
nor U316 (N_316,In_406,In_198);
nand U317 (N_317,In_15,In_42);
or U318 (N_318,In_362,In_330);
nand U319 (N_319,In_20,In_230);
nand U320 (N_320,In_462,In_81);
and U321 (N_321,In_34,In_288);
and U322 (N_322,In_278,In_452);
nor U323 (N_323,In_379,In_472);
or U324 (N_324,In_3,In_378);
and U325 (N_325,In_136,In_14);
nor U326 (N_326,In_401,In_348);
nand U327 (N_327,In_129,In_70);
and U328 (N_328,In_144,In_31);
nor U329 (N_329,In_275,In_140);
nor U330 (N_330,In_243,In_169);
nor U331 (N_331,In_298,In_456);
nand U332 (N_332,In_15,In_357);
nand U333 (N_333,In_40,In_10);
nor U334 (N_334,In_274,In_82);
and U335 (N_335,In_33,In_292);
or U336 (N_336,In_391,In_67);
or U337 (N_337,In_141,In_349);
nand U338 (N_338,In_40,In_214);
and U339 (N_339,In_115,In_178);
nor U340 (N_340,In_493,In_63);
and U341 (N_341,In_195,In_177);
and U342 (N_342,In_253,In_322);
or U343 (N_343,In_288,In_199);
or U344 (N_344,In_229,In_471);
nand U345 (N_345,In_165,In_166);
nor U346 (N_346,In_206,In_168);
and U347 (N_347,In_424,In_6);
or U348 (N_348,In_205,In_484);
and U349 (N_349,In_63,In_300);
and U350 (N_350,In_87,In_387);
nor U351 (N_351,In_139,In_345);
and U352 (N_352,In_258,In_345);
and U353 (N_353,In_480,In_324);
nand U354 (N_354,In_277,In_286);
nand U355 (N_355,In_147,In_174);
or U356 (N_356,In_165,In_69);
or U357 (N_357,In_362,In_352);
nand U358 (N_358,In_241,In_432);
and U359 (N_359,In_481,In_464);
nor U360 (N_360,In_63,In_73);
nand U361 (N_361,In_256,In_414);
nand U362 (N_362,In_476,In_46);
nand U363 (N_363,In_379,In_27);
or U364 (N_364,In_80,In_145);
and U365 (N_365,In_147,In_263);
nor U366 (N_366,In_55,In_154);
and U367 (N_367,In_83,In_333);
or U368 (N_368,In_345,In_57);
nand U369 (N_369,In_497,In_499);
and U370 (N_370,In_443,In_457);
and U371 (N_371,In_207,In_172);
nor U372 (N_372,In_477,In_349);
and U373 (N_373,In_429,In_35);
nand U374 (N_374,In_421,In_250);
and U375 (N_375,In_78,In_151);
and U376 (N_376,In_223,In_98);
and U377 (N_377,In_151,In_342);
nor U378 (N_378,In_124,In_206);
or U379 (N_379,In_183,In_355);
xor U380 (N_380,In_295,In_70);
or U381 (N_381,In_233,In_271);
nand U382 (N_382,In_427,In_455);
nand U383 (N_383,In_75,In_6);
or U384 (N_384,In_9,In_477);
or U385 (N_385,In_193,In_283);
or U386 (N_386,In_14,In_191);
and U387 (N_387,In_109,In_404);
nand U388 (N_388,In_27,In_171);
nand U389 (N_389,In_307,In_420);
nand U390 (N_390,In_460,In_83);
nand U391 (N_391,In_1,In_55);
or U392 (N_392,In_208,In_168);
nand U393 (N_393,In_462,In_420);
nand U394 (N_394,In_102,In_35);
nand U395 (N_395,In_33,In_127);
or U396 (N_396,In_133,In_140);
nand U397 (N_397,In_217,In_459);
nor U398 (N_398,In_327,In_433);
nand U399 (N_399,In_190,In_168);
nand U400 (N_400,In_271,In_101);
or U401 (N_401,In_350,In_117);
and U402 (N_402,In_481,In_19);
nor U403 (N_403,In_473,In_301);
and U404 (N_404,In_146,In_83);
and U405 (N_405,In_0,In_191);
or U406 (N_406,In_458,In_80);
nor U407 (N_407,In_298,In_68);
nor U408 (N_408,In_232,In_426);
nor U409 (N_409,In_382,In_148);
nor U410 (N_410,In_309,In_81);
nor U411 (N_411,In_489,In_317);
or U412 (N_412,In_489,In_155);
nor U413 (N_413,In_118,In_478);
nor U414 (N_414,In_392,In_209);
or U415 (N_415,In_28,In_306);
and U416 (N_416,In_308,In_270);
nand U417 (N_417,In_344,In_347);
nand U418 (N_418,In_55,In_136);
and U419 (N_419,In_374,In_301);
xor U420 (N_420,In_203,In_464);
and U421 (N_421,In_330,In_413);
or U422 (N_422,In_99,In_64);
nor U423 (N_423,In_303,In_392);
nor U424 (N_424,In_257,In_82);
or U425 (N_425,In_386,In_451);
nor U426 (N_426,In_442,In_320);
nor U427 (N_427,In_11,In_412);
nor U428 (N_428,In_174,In_0);
or U429 (N_429,In_219,In_121);
nor U430 (N_430,In_257,In_191);
and U431 (N_431,In_289,In_4);
and U432 (N_432,In_439,In_9);
nor U433 (N_433,In_489,In_27);
xnor U434 (N_434,In_89,In_165);
nand U435 (N_435,In_385,In_301);
nand U436 (N_436,In_26,In_429);
and U437 (N_437,In_267,In_97);
and U438 (N_438,In_119,In_256);
and U439 (N_439,In_303,In_337);
and U440 (N_440,In_153,In_88);
nand U441 (N_441,In_165,In_250);
nor U442 (N_442,In_473,In_287);
and U443 (N_443,In_219,In_285);
and U444 (N_444,In_157,In_223);
nor U445 (N_445,In_81,In_302);
nor U446 (N_446,In_491,In_466);
nor U447 (N_447,In_368,In_87);
or U448 (N_448,In_255,In_436);
and U449 (N_449,In_416,In_356);
and U450 (N_450,In_138,In_471);
nand U451 (N_451,In_377,In_230);
nand U452 (N_452,In_264,In_496);
or U453 (N_453,In_101,In_219);
and U454 (N_454,In_447,In_18);
or U455 (N_455,In_450,In_217);
nor U456 (N_456,In_392,In_157);
nor U457 (N_457,In_101,In_233);
or U458 (N_458,In_225,In_51);
nor U459 (N_459,In_113,In_360);
and U460 (N_460,In_145,In_492);
or U461 (N_461,In_137,In_483);
and U462 (N_462,In_174,In_284);
and U463 (N_463,In_124,In_10);
and U464 (N_464,In_142,In_382);
xor U465 (N_465,In_346,In_465);
nand U466 (N_466,In_142,In_270);
and U467 (N_467,In_427,In_465);
and U468 (N_468,In_13,In_275);
and U469 (N_469,In_289,In_292);
and U470 (N_470,In_29,In_457);
or U471 (N_471,In_333,In_217);
or U472 (N_472,In_171,In_456);
or U473 (N_473,In_361,In_13);
nor U474 (N_474,In_389,In_222);
or U475 (N_475,In_226,In_91);
and U476 (N_476,In_192,In_71);
nand U477 (N_477,In_287,In_217);
nand U478 (N_478,In_163,In_76);
and U479 (N_479,In_471,In_378);
nor U480 (N_480,In_328,In_7);
nand U481 (N_481,In_326,In_450);
or U482 (N_482,In_188,In_43);
and U483 (N_483,In_123,In_152);
nor U484 (N_484,In_220,In_185);
or U485 (N_485,In_343,In_166);
nand U486 (N_486,In_329,In_40);
or U487 (N_487,In_196,In_472);
and U488 (N_488,In_386,In_245);
nor U489 (N_489,In_473,In_211);
nor U490 (N_490,In_56,In_98);
nor U491 (N_491,In_197,In_371);
nor U492 (N_492,In_313,In_227);
and U493 (N_493,In_386,In_177);
or U494 (N_494,In_144,In_2);
nor U495 (N_495,In_347,In_77);
nand U496 (N_496,In_487,In_79);
and U497 (N_497,In_290,In_190);
nand U498 (N_498,In_16,In_73);
or U499 (N_499,In_352,In_259);
nand U500 (N_500,N_109,N_360);
nor U501 (N_501,N_395,N_444);
and U502 (N_502,N_384,N_397);
or U503 (N_503,N_299,N_349);
or U504 (N_504,N_436,N_197);
nor U505 (N_505,N_68,N_31);
nand U506 (N_506,N_117,N_99);
nand U507 (N_507,N_276,N_406);
nand U508 (N_508,N_58,N_171);
nor U509 (N_509,N_93,N_187);
or U510 (N_510,N_465,N_253);
nor U511 (N_511,N_326,N_199);
nor U512 (N_512,N_402,N_289);
and U513 (N_513,N_261,N_420);
nand U514 (N_514,N_466,N_7);
and U515 (N_515,N_365,N_305);
nor U516 (N_516,N_39,N_316);
nor U517 (N_517,N_104,N_138);
xor U518 (N_518,N_27,N_449);
or U519 (N_519,N_270,N_181);
nand U520 (N_520,N_461,N_135);
nor U521 (N_521,N_67,N_63);
nand U522 (N_522,N_419,N_306);
or U523 (N_523,N_491,N_370);
nand U524 (N_524,N_48,N_437);
xor U525 (N_525,N_154,N_344);
or U526 (N_526,N_248,N_149);
and U527 (N_527,N_340,N_488);
nor U528 (N_528,N_164,N_36);
and U529 (N_529,N_453,N_490);
nor U530 (N_530,N_390,N_237);
nand U531 (N_531,N_5,N_214);
and U532 (N_532,N_217,N_247);
and U533 (N_533,N_336,N_274);
nand U534 (N_534,N_464,N_317);
nand U535 (N_535,N_80,N_339);
xor U536 (N_536,N_169,N_298);
and U537 (N_537,N_242,N_28);
nor U538 (N_538,N_376,N_119);
nor U539 (N_539,N_50,N_189);
and U540 (N_540,N_489,N_106);
nand U541 (N_541,N_100,N_160);
nor U542 (N_542,N_126,N_405);
or U543 (N_543,N_128,N_16);
nand U544 (N_544,N_13,N_215);
nand U545 (N_545,N_355,N_127);
nor U546 (N_546,N_252,N_179);
and U547 (N_547,N_140,N_312);
nand U548 (N_548,N_266,N_441);
and U549 (N_549,N_57,N_327);
or U550 (N_550,N_224,N_467);
nand U551 (N_551,N_219,N_469);
and U552 (N_552,N_14,N_265);
or U553 (N_553,N_358,N_485);
nor U554 (N_554,N_451,N_329);
and U555 (N_555,N_262,N_51);
or U556 (N_556,N_331,N_124);
nand U557 (N_557,N_22,N_120);
and U558 (N_558,N_474,N_300);
and U559 (N_559,N_385,N_426);
nand U560 (N_560,N_278,N_92);
or U561 (N_561,N_146,N_174);
and U562 (N_562,N_351,N_211);
or U563 (N_563,N_35,N_462);
nand U564 (N_564,N_379,N_123);
nor U565 (N_565,N_62,N_56);
or U566 (N_566,N_408,N_4);
and U567 (N_567,N_378,N_328);
or U568 (N_568,N_495,N_87);
or U569 (N_569,N_368,N_313);
and U570 (N_570,N_221,N_223);
nand U571 (N_571,N_264,N_193);
xor U572 (N_572,N_134,N_170);
or U573 (N_573,N_269,N_161);
or U574 (N_574,N_144,N_256);
nand U575 (N_575,N_244,N_184);
and U576 (N_576,N_400,N_333);
nand U577 (N_577,N_69,N_347);
nand U578 (N_578,N_91,N_319);
nor U579 (N_579,N_2,N_431);
and U580 (N_580,N_111,N_168);
and U581 (N_581,N_345,N_295);
nand U582 (N_582,N_238,N_52);
xor U583 (N_583,N_251,N_387);
nand U584 (N_584,N_70,N_482);
and U585 (N_585,N_407,N_335);
and U586 (N_586,N_225,N_9);
nor U587 (N_587,N_226,N_367);
nor U588 (N_588,N_115,N_83);
nor U589 (N_589,N_157,N_425);
nand U590 (N_590,N_112,N_37);
nand U591 (N_591,N_43,N_103);
xor U592 (N_592,N_353,N_77);
nor U593 (N_593,N_381,N_228);
nor U594 (N_594,N_352,N_84);
or U595 (N_595,N_195,N_210);
nand U596 (N_596,N_396,N_290);
and U597 (N_597,N_363,N_3);
and U598 (N_598,N_372,N_229);
nor U599 (N_599,N_393,N_343);
and U600 (N_600,N_121,N_125);
and U601 (N_601,N_143,N_220);
nand U602 (N_602,N_216,N_325);
nand U603 (N_603,N_45,N_222);
nor U604 (N_604,N_59,N_75);
nor U605 (N_605,N_296,N_452);
or U606 (N_606,N_19,N_8);
and U607 (N_607,N_416,N_279);
or U608 (N_608,N_64,N_356);
or U609 (N_609,N_101,N_424);
or U610 (N_610,N_342,N_472);
and U611 (N_611,N_131,N_475);
nand U612 (N_612,N_173,N_362);
or U613 (N_613,N_292,N_341);
or U614 (N_614,N_139,N_324);
and U615 (N_615,N_71,N_422);
nor U616 (N_616,N_359,N_245);
nor U617 (N_617,N_213,N_205);
nand U618 (N_618,N_130,N_81);
or U619 (N_619,N_209,N_439);
nor U620 (N_620,N_54,N_255);
or U621 (N_621,N_456,N_191);
nand U622 (N_622,N_357,N_203);
nand U623 (N_623,N_95,N_497);
and U624 (N_624,N_309,N_481);
or U625 (N_625,N_41,N_243);
nor U626 (N_626,N_311,N_460);
nor U627 (N_627,N_96,N_320);
or U628 (N_628,N_304,N_133);
nor U629 (N_629,N_230,N_301);
nor U630 (N_630,N_24,N_204);
nand U631 (N_631,N_334,N_55);
nand U632 (N_632,N_231,N_142);
or U633 (N_633,N_116,N_239);
and U634 (N_634,N_90,N_373);
nor U635 (N_635,N_94,N_183);
and U636 (N_636,N_180,N_442);
and U637 (N_637,N_177,N_61);
nor U638 (N_638,N_283,N_182);
and U639 (N_639,N_30,N_136);
or U640 (N_640,N_236,N_188);
or U641 (N_641,N_459,N_207);
nor U642 (N_642,N_40,N_20);
and U643 (N_643,N_132,N_158);
nor U644 (N_644,N_414,N_273);
nor U645 (N_645,N_468,N_318);
and U646 (N_646,N_487,N_33);
nor U647 (N_647,N_389,N_401);
and U648 (N_648,N_354,N_47);
or U649 (N_649,N_473,N_369);
and U650 (N_650,N_293,N_186);
and U651 (N_651,N_302,N_294);
or U652 (N_652,N_44,N_152);
or U653 (N_653,N_26,N_218);
or U654 (N_654,N_268,N_15);
nand U655 (N_655,N_286,N_162);
or U656 (N_656,N_282,N_122);
nor U657 (N_657,N_185,N_12);
nor U658 (N_658,N_235,N_23);
and U659 (N_659,N_201,N_386);
nand U660 (N_660,N_249,N_73);
and U661 (N_661,N_454,N_105);
nand U662 (N_662,N_153,N_438);
and U663 (N_663,N_78,N_263);
and U664 (N_664,N_267,N_178);
and U665 (N_665,N_445,N_34);
and U666 (N_666,N_108,N_435);
nor U667 (N_667,N_165,N_323);
nor U668 (N_668,N_60,N_254);
nor U669 (N_669,N_1,N_163);
or U670 (N_670,N_0,N_42);
or U671 (N_671,N_76,N_257);
nand U672 (N_672,N_196,N_348);
and U673 (N_673,N_374,N_88);
nand U674 (N_674,N_89,N_291);
nand U675 (N_675,N_307,N_428);
nor U676 (N_676,N_110,N_308);
nor U677 (N_677,N_32,N_498);
nor U678 (N_678,N_477,N_403);
nand U679 (N_679,N_478,N_382);
nor U680 (N_680,N_72,N_303);
nor U681 (N_681,N_212,N_148);
or U682 (N_682,N_145,N_29);
nor U683 (N_683,N_337,N_480);
xnor U684 (N_684,N_383,N_11);
nor U685 (N_685,N_330,N_113);
and U686 (N_686,N_53,N_496);
and U687 (N_687,N_150,N_366);
nor U688 (N_688,N_484,N_38);
nor U689 (N_689,N_440,N_198);
or U690 (N_690,N_206,N_6);
nor U691 (N_691,N_391,N_155);
nand U692 (N_692,N_486,N_97);
or U693 (N_693,N_375,N_494);
and U694 (N_694,N_492,N_322);
and U695 (N_695,N_151,N_280);
nor U696 (N_696,N_297,N_246);
and U697 (N_697,N_272,N_102);
xnor U698 (N_698,N_194,N_250);
nand U699 (N_699,N_271,N_338);
nor U700 (N_700,N_404,N_74);
nor U701 (N_701,N_277,N_192);
nand U702 (N_702,N_394,N_166);
or U703 (N_703,N_259,N_281);
or U704 (N_704,N_399,N_432);
nor U705 (N_705,N_200,N_172);
nor U706 (N_706,N_463,N_227);
nand U707 (N_707,N_240,N_380);
nand U708 (N_708,N_447,N_415);
nand U709 (N_709,N_364,N_458);
nand U710 (N_710,N_417,N_287);
and U711 (N_711,N_25,N_470);
nand U712 (N_712,N_65,N_457);
nor U713 (N_713,N_175,N_314);
and U714 (N_714,N_423,N_85);
or U715 (N_715,N_202,N_232);
nor U716 (N_716,N_388,N_476);
or U717 (N_717,N_241,N_377);
nand U718 (N_718,N_421,N_361);
nand U719 (N_719,N_159,N_471);
or U720 (N_720,N_208,N_409);
and U721 (N_721,N_66,N_17);
nor U722 (N_722,N_190,N_114);
or U723 (N_723,N_82,N_147);
or U724 (N_724,N_392,N_350);
nor U725 (N_725,N_371,N_137);
nand U726 (N_726,N_98,N_430);
nand U727 (N_727,N_260,N_499);
nor U728 (N_728,N_411,N_493);
nand U729 (N_729,N_46,N_450);
and U730 (N_730,N_433,N_448);
and U731 (N_731,N_315,N_129);
nand U732 (N_732,N_413,N_176);
nor U733 (N_733,N_49,N_427);
and U734 (N_734,N_455,N_79);
and U735 (N_735,N_332,N_118);
or U736 (N_736,N_86,N_233);
nor U737 (N_737,N_285,N_418);
or U738 (N_738,N_258,N_443);
nor U739 (N_739,N_483,N_410);
and U740 (N_740,N_21,N_412);
nor U741 (N_741,N_288,N_321);
and U742 (N_742,N_275,N_234);
and U743 (N_743,N_10,N_107);
nand U744 (N_744,N_434,N_446);
and U745 (N_745,N_284,N_18);
or U746 (N_746,N_156,N_479);
nor U747 (N_747,N_429,N_167);
or U748 (N_748,N_398,N_141);
xnor U749 (N_749,N_346,N_310);
nand U750 (N_750,N_329,N_132);
or U751 (N_751,N_497,N_440);
and U752 (N_752,N_11,N_297);
nor U753 (N_753,N_367,N_105);
nor U754 (N_754,N_412,N_50);
nand U755 (N_755,N_429,N_218);
nor U756 (N_756,N_44,N_138);
nor U757 (N_757,N_283,N_362);
or U758 (N_758,N_45,N_279);
nand U759 (N_759,N_255,N_78);
and U760 (N_760,N_376,N_11);
nand U761 (N_761,N_430,N_437);
nand U762 (N_762,N_477,N_80);
and U763 (N_763,N_240,N_232);
nor U764 (N_764,N_308,N_283);
or U765 (N_765,N_8,N_11);
nand U766 (N_766,N_103,N_74);
or U767 (N_767,N_1,N_232);
or U768 (N_768,N_117,N_155);
or U769 (N_769,N_402,N_144);
nor U770 (N_770,N_15,N_345);
xnor U771 (N_771,N_316,N_101);
nor U772 (N_772,N_387,N_18);
and U773 (N_773,N_14,N_38);
nand U774 (N_774,N_257,N_391);
and U775 (N_775,N_496,N_176);
nor U776 (N_776,N_110,N_171);
nor U777 (N_777,N_152,N_132);
nand U778 (N_778,N_460,N_253);
or U779 (N_779,N_81,N_80);
and U780 (N_780,N_290,N_160);
or U781 (N_781,N_341,N_83);
nand U782 (N_782,N_391,N_356);
nor U783 (N_783,N_476,N_99);
and U784 (N_784,N_117,N_143);
nand U785 (N_785,N_339,N_52);
nor U786 (N_786,N_164,N_244);
and U787 (N_787,N_486,N_274);
and U788 (N_788,N_469,N_77);
and U789 (N_789,N_249,N_260);
nand U790 (N_790,N_463,N_181);
and U791 (N_791,N_170,N_399);
nor U792 (N_792,N_195,N_300);
nor U793 (N_793,N_215,N_237);
and U794 (N_794,N_401,N_243);
nand U795 (N_795,N_276,N_186);
or U796 (N_796,N_238,N_417);
nor U797 (N_797,N_224,N_21);
nor U798 (N_798,N_42,N_358);
and U799 (N_799,N_124,N_113);
and U800 (N_800,N_56,N_356);
nand U801 (N_801,N_242,N_308);
and U802 (N_802,N_376,N_343);
and U803 (N_803,N_318,N_63);
nor U804 (N_804,N_51,N_23);
and U805 (N_805,N_465,N_147);
or U806 (N_806,N_319,N_10);
nor U807 (N_807,N_18,N_376);
nor U808 (N_808,N_258,N_303);
nand U809 (N_809,N_232,N_360);
and U810 (N_810,N_413,N_319);
nand U811 (N_811,N_346,N_347);
or U812 (N_812,N_191,N_215);
and U813 (N_813,N_46,N_408);
nor U814 (N_814,N_326,N_317);
or U815 (N_815,N_378,N_158);
or U816 (N_816,N_26,N_107);
or U817 (N_817,N_38,N_267);
or U818 (N_818,N_429,N_357);
and U819 (N_819,N_65,N_129);
nand U820 (N_820,N_468,N_238);
nor U821 (N_821,N_192,N_246);
or U822 (N_822,N_375,N_310);
nor U823 (N_823,N_215,N_147);
nand U824 (N_824,N_206,N_300);
nor U825 (N_825,N_419,N_216);
and U826 (N_826,N_408,N_357);
nand U827 (N_827,N_496,N_302);
nor U828 (N_828,N_30,N_67);
and U829 (N_829,N_217,N_348);
nor U830 (N_830,N_428,N_16);
nor U831 (N_831,N_334,N_201);
nor U832 (N_832,N_190,N_284);
and U833 (N_833,N_273,N_191);
nor U834 (N_834,N_0,N_166);
nand U835 (N_835,N_391,N_85);
and U836 (N_836,N_325,N_483);
and U837 (N_837,N_391,N_486);
nor U838 (N_838,N_83,N_385);
nand U839 (N_839,N_218,N_356);
nand U840 (N_840,N_160,N_476);
and U841 (N_841,N_92,N_236);
and U842 (N_842,N_281,N_5);
nor U843 (N_843,N_291,N_42);
or U844 (N_844,N_350,N_89);
or U845 (N_845,N_255,N_168);
nand U846 (N_846,N_170,N_366);
and U847 (N_847,N_188,N_217);
and U848 (N_848,N_78,N_386);
nor U849 (N_849,N_51,N_439);
nand U850 (N_850,N_224,N_331);
and U851 (N_851,N_135,N_145);
nor U852 (N_852,N_34,N_470);
nor U853 (N_853,N_335,N_6);
and U854 (N_854,N_55,N_475);
nor U855 (N_855,N_154,N_421);
or U856 (N_856,N_405,N_164);
or U857 (N_857,N_224,N_273);
nor U858 (N_858,N_383,N_381);
and U859 (N_859,N_119,N_321);
nor U860 (N_860,N_39,N_67);
or U861 (N_861,N_403,N_244);
and U862 (N_862,N_187,N_424);
nand U863 (N_863,N_485,N_215);
nand U864 (N_864,N_424,N_220);
nand U865 (N_865,N_243,N_447);
and U866 (N_866,N_441,N_204);
and U867 (N_867,N_122,N_479);
or U868 (N_868,N_57,N_421);
nor U869 (N_869,N_205,N_299);
nor U870 (N_870,N_266,N_80);
nand U871 (N_871,N_363,N_139);
nor U872 (N_872,N_440,N_179);
and U873 (N_873,N_296,N_138);
or U874 (N_874,N_180,N_438);
nor U875 (N_875,N_462,N_174);
nor U876 (N_876,N_329,N_206);
nand U877 (N_877,N_318,N_68);
and U878 (N_878,N_288,N_141);
nor U879 (N_879,N_269,N_353);
nor U880 (N_880,N_265,N_153);
xnor U881 (N_881,N_95,N_87);
and U882 (N_882,N_430,N_398);
and U883 (N_883,N_193,N_270);
nand U884 (N_884,N_62,N_54);
or U885 (N_885,N_183,N_7);
and U886 (N_886,N_284,N_237);
nor U887 (N_887,N_312,N_419);
nand U888 (N_888,N_44,N_161);
xor U889 (N_889,N_149,N_131);
or U890 (N_890,N_95,N_242);
nor U891 (N_891,N_311,N_15);
and U892 (N_892,N_51,N_0);
nor U893 (N_893,N_37,N_173);
nor U894 (N_894,N_305,N_386);
or U895 (N_895,N_162,N_424);
nand U896 (N_896,N_190,N_24);
and U897 (N_897,N_70,N_448);
and U898 (N_898,N_3,N_386);
nor U899 (N_899,N_249,N_265);
nor U900 (N_900,N_61,N_326);
or U901 (N_901,N_224,N_127);
nand U902 (N_902,N_29,N_51);
nand U903 (N_903,N_225,N_273);
nor U904 (N_904,N_423,N_327);
xnor U905 (N_905,N_326,N_430);
or U906 (N_906,N_149,N_444);
or U907 (N_907,N_1,N_11);
nand U908 (N_908,N_357,N_94);
nand U909 (N_909,N_170,N_68);
or U910 (N_910,N_126,N_193);
nor U911 (N_911,N_18,N_394);
nor U912 (N_912,N_20,N_370);
or U913 (N_913,N_270,N_465);
or U914 (N_914,N_182,N_242);
or U915 (N_915,N_4,N_499);
and U916 (N_916,N_243,N_297);
or U917 (N_917,N_396,N_47);
or U918 (N_918,N_245,N_161);
nand U919 (N_919,N_192,N_363);
or U920 (N_920,N_382,N_310);
or U921 (N_921,N_461,N_78);
nand U922 (N_922,N_478,N_63);
nand U923 (N_923,N_356,N_342);
nor U924 (N_924,N_299,N_409);
nand U925 (N_925,N_135,N_460);
nand U926 (N_926,N_143,N_37);
nor U927 (N_927,N_117,N_98);
nand U928 (N_928,N_377,N_373);
nor U929 (N_929,N_219,N_305);
nor U930 (N_930,N_33,N_405);
and U931 (N_931,N_335,N_23);
nor U932 (N_932,N_209,N_460);
and U933 (N_933,N_449,N_144);
or U934 (N_934,N_104,N_212);
nor U935 (N_935,N_241,N_245);
or U936 (N_936,N_339,N_61);
or U937 (N_937,N_127,N_212);
nand U938 (N_938,N_464,N_69);
nor U939 (N_939,N_29,N_75);
or U940 (N_940,N_277,N_207);
nor U941 (N_941,N_118,N_164);
and U942 (N_942,N_475,N_295);
and U943 (N_943,N_77,N_446);
and U944 (N_944,N_92,N_369);
or U945 (N_945,N_166,N_367);
nand U946 (N_946,N_65,N_142);
nand U947 (N_947,N_18,N_493);
and U948 (N_948,N_188,N_472);
and U949 (N_949,N_366,N_451);
nor U950 (N_950,N_292,N_498);
and U951 (N_951,N_348,N_3);
or U952 (N_952,N_56,N_437);
and U953 (N_953,N_85,N_162);
nor U954 (N_954,N_379,N_397);
and U955 (N_955,N_175,N_171);
nor U956 (N_956,N_408,N_73);
nand U957 (N_957,N_408,N_152);
nor U958 (N_958,N_450,N_9);
nand U959 (N_959,N_443,N_463);
nand U960 (N_960,N_426,N_339);
nand U961 (N_961,N_56,N_231);
nand U962 (N_962,N_435,N_306);
nor U963 (N_963,N_380,N_228);
and U964 (N_964,N_239,N_92);
and U965 (N_965,N_416,N_326);
and U966 (N_966,N_128,N_71);
nand U967 (N_967,N_222,N_23);
nand U968 (N_968,N_141,N_171);
nand U969 (N_969,N_199,N_177);
nand U970 (N_970,N_388,N_444);
and U971 (N_971,N_332,N_382);
and U972 (N_972,N_418,N_469);
or U973 (N_973,N_131,N_8);
or U974 (N_974,N_355,N_475);
and U975 (N_975,N_93,N_455);
nand U976 (N_976,N_326,N_173);
or U977 (N_977,N_304,N_226);
or U978 (N_978,N_146,N_178);
or U979 (N_979,N_272,N_458);
nand U980 (N_980,N_5,N_221);
and U981 (N_981,N_430,N_246);
and U982 (N_982,N_372,N_226);
and U983 (N_983,N_321,N_404);
nand U984 (N_984,N_68,N_131);
nand U985 (N_985,N_485,N_170);
xnor U986 (N_986,N_47,N_52);
or U987 (N_987,N_402,N_14);
and U988 (N_988,N_258,N_155);
or U989 (N_989,N_106,N_419);
and U990 (N_990,N_129,N_276);
nand U991 (N_991,N_307,N_81);
nor U992 (N_992,N_34,N_241);
or U993 (N_993,N_144,N_73);
or U994 (N_994,N_43,N_319);
nand U995 (N_995,N_92,N_271);
nand U996 (N_996,N_445,N_268);
or U997 (N_997,N_402,N_159);
nand U998 (N_998,N_261,N_377);
or U999 (N_999,N_70,N_36);
nor U1000 (N_1000,N_529,N_549);
and U1001 (N_1001,N_883,N_710);
nor U1002 (N_1002,N_881,N_760);
nor U1003 (N_1003,N_745,N_641);
and U1004 (N_1004,N_698,N_598);
nand U1005 (N_1005,N_665,N_919);
and U1006 (N_1006,N_930,N_993);
nand U1007 (N_1007,N_691,N_786);
or U1008 (N_1008,N_530,N_878);
and U1009 (N_1009,N_850,N_650);
nand U1010 (N_1010,N_532,N_709);
and U1011 (N_1011,N_540,N_574);
nor U1012 (N_1012,N_992,N_704);
or U1013 (N_1013,N_946,N_884);
and U1014 (N_1014,N_563,N_829);
and U1015 (N_1015,N_871,N_923);
nand U1016 (N_1016,N_679,N_629);
nand U1017 (N_1017,N_505,N_973);
and U1018 (N_1018,N_990,N_651);
nand U1019 (N_1019,N_949,N_776);
or U1020 (N_1020,N_766,N_795);
and U1021 (N_1021,N_703,N_890);
nand U1022 (N_1022,N_644,N_761);
or U1023 (N_1023,N_824,N_654);
or U1024 (N_1024,N_711,N_769);
xnor U1025 (N_1025,N_569,N_979);
and U1026 (N_1026,N_667,N_578);
nor U1027 (N_1027,N_697,N_562);
nor U1028 (N_1028,N_610,N_921);
nand U1029 (N_1029,N_669,N_891);
nor U1030 (N_1030,N_594,N_660);
or U1031 (N_1031,N_823,N_767);
or U1032 (N_1032,N_974,N_655);
nand U1033 (N_1033,N_879,N_646);
nor U1034 (N_1034,N_758,N_920);
nor U1035 (N_1035,N_794,N_945);
and U1036 (N_1036,N_896,N_603);
or U1037 (N_1037,N_846,N_686);
or U1038 (N_1038,N_936,N_814);
or U1039 (N_1039,N_510,N_753);
nand U1040 (N_1040,N_955,N_750);
nand U1041 (N_1041,N_685,N_674);
nand U1042 (N_1042,N_770,N_803);
nor U1043 (N_1043,N_820,N_601);
xor U1044 (N_1044,N_783,N_564);
nor U1045 (N_1045,N_707,N_922);
nor U1046 (N_1046,N_980,N_589);
nor U1047 (N_1047,N_966,N_619);
nand U1048 (N_1048,N_643,N_793);
and U1049 (N_1049,N_799,N_577);
nand U1050 (N_1050,N_757,N_721);
and U1051 (N_1051,N_501,N_845);
nor U1052 (N_1052,N_587,N_746);
nor U1053 (N_1053,N_908,N_940);
or U1054 (N_1054,N_841,N_672);
or U1055 (N_1055,N_995,N_560);
and U1056 (N_1056,N_642,N_625);
or U1057 (N_1057,N_907,N_666);
or U1058 (N_1058,N_680,N_544);
nor U1059 (N_1059,N_780,N_886);
nor U1060 (N_1060,N_899,N_606);
or U1061 (N_1061,N_618,N_627);
or U1062 (N_1062,N_602,N_938);
nor U1063 (N_1063,N_866,N_503);
and U1064 (N_1064,N_694,N_706);
or U1065 (N_1065,N_843,N_984);
and U1066 (N_1066,N_838,N_559);
xnor U1067 (N_1067,N_839,N_781);
nand U1068 (N_1068,N_914,N_621);
or U1069 (N_1069,N_668,N_673);
nand U1070 (N_1070,N_880,N_634);
or U1071 (N_1071,N_844,N_546);
nor U1072 (N_1072,N_681,N_678);
or U1073 (N_1073,N_897,N_613);
or U1074 (N_1074,N_658,N_515);
and U1075 (N_1075,N_999,N_657);
nor U1076 (N_1076,N_944,N_916);
and U1077 (N_1077,N_591,N_818);
nand U1078 (N_1078,N_608,N_616);
or U1079 (N_1079,N_821,N_759);
nor U1080 (N_1080,N_726,N_526);
and U1081 (N_1081,N_933,N_519);
nor U1082 (N_1082,N_904,N_701);
nand U1083 (N_1083,N_531,N_538);
nand U1084 (N_1084,N_763,N_804);
or U1085 (N_1085,N_715,N_954);
nand U1086 (N_1086,N_988,N_533);
nor U1087 (N_1087,N_645,N_848);
nand U1088 (N_1088,N_663,N_557);
nor U1089 (N_1089,N_552,N_942);
nor U1090 (N_1090,N_637,N_514);
and U1091 (N_1091,N_611,N_732);
nor U1092 (N_1092,N_527,N_893);
nand U1093 (N_1093,N_813,N_702);
nand U1094 (N_1094,N_777,N_649);
nor U1095 (N_1095,N_830,N_885);
nor U1096 (N_1096,N_507,N_797);
nand U1097 (N_1097,N_571,N_545);
or U1098 (N_1098,N_730,N_772);
nand U1099 (N_1099,N_805,N_860);
or U1100 (N_1100,N_985,N_689);
nand U1101 (N_1101,N_963,N_947);
and U1102 (N_1102,N_652,N_909);
nor U1103 (N_1103,N_582,N_934);
nand U1104 (N_1104,N_892,N_956);
or U1105 (N_1105,N_828,N_605);
nor U1106 (N_1106,N_748,N_517);
nand U1107 (N_1107,N_851,N_653);
nand U1108 (N_1108,N_690,N_600);
or U1109 (N_1109,N_957,N_539);
nor U1110 (N_1110,N_599,N_849);
and U1111 (N_1111,N_719,N_688);
or U1112 (N_1112,N_926,N_989);
or U1113 (N_1113,N_811,N_981);
nor U1114 (N_1114,N_521,N_874);
nand U1115 (N_1115,N_536,N_854);
or U1116 (N_1116,N_903,N_792);
or U1117 (N_1117,N_834,N_617);
and U1118 (N_1118,N_717,N_740);
nand U1119 (N_1119,N_856,N_534);
or U1120 (N_1120,N_692,N_831);
and U1121 (N_1121,N_822,N_796);
nor U1122 (N_1122,N_508,N_877);
or U1123 (N_1123,N_743,N_550);
nor U1124 (N_1124,N_768,N_506);
or U1125 (N_1125,N_960,N_982);
nand U1126 (N_1126,N_789,N_581);
or U1127 (N_1127,N_819,N_593);
nor U1128 (N_1128,N_631,N_867);
nor U1129 (N_1129,N_572,N_548);
nand U1130 (N_1130,N_716,N_784);
nand U1131 (N_1131,N_615,N_713);
nor U1132 (N_1132,N_551,N_778);
nor U1133 (N_1133,N_764,N_810);
nand U1134 (N_1134,N_958,N_728);
nor U1135 (N_1135,N_827,N_971);
nand U1136 (N_1136,N_628,N_788);
or U1137 (N_1137,N_976,N_500);
nor U1138 (N_1138,N_928,N_579);
and U1139 (N_1139,N_870,N_873);
nor U1140 (N_1140,N_809,N_755);
nand U1141 (N_1141,N_939,N_970);
or U1142 (N_1142,N_895,N_925);
nor U1143 (N_1143,N_935,N_576);
or U1144 (N_1144,N_638,N_596);
nor U1145 (N_1145,N_585,N_623);
nand U1146 (N_1146,N_962,N_951);
nand U1147 (N_1147,N_901,N_541);
nor U1148 (N_1148,N_953,N_670);
and U1149 (N_1149,N_977,N_659);
and U1150 (N_1150,N_937,N_543);
nor U1151 (N_1151,N_575,N_520);
or U1152 (N_1152,N_699,N_558);
nand U1153 (N_1153,N_913,N_727);
nand U1154 (N_1154,N_910,N_861);
nand U1155 (N_1155,N_556,N_900);
nor U1156 (N_1156,N_733,N_840);
or U1157 (N_1157,N_554,N_537);
nor U1158 (N_1158,N_887,N_798);
nand U1159 (N_1159,N_927,N_588);
nor U1160 (N_1160,N_917,N_852);
nor U1161 (N_1161,N_965,N_725);
nor U1162 (N_1162,N_647,N_662);
or U1163 (N_1163,N_911,N_518);
nor U1164 (N_1164,N_742,N_918);
nor U1165 (N_1165,N_722,N_782);
and U1166 (N_1166,N_693,N_773);
and U1167 (N_1167,N_528,N_718);
and U1168 (N_1168,N_708,N_570);
nor U1169 (N_1169,N_876,N_524);
nor U1170 (N_1170,N_565,N_676);
nand U1171 (N_1171,N_547,N_889);
nand U1172 (N_1172,N_636,N_986);
and U1173 (N_1173,N_705,N_620);
and U1174 (N_1174,N_535,N_696);
nor U1175 (N_1175,N_864,N_592);
nor U1176 (N_1176,N_682,N_941);
or U1177 (N_1177,N_857,N_671);
nor U1178 (N_1178,N_888,N_630);
nor U1179 (N_1179,N_633,N_561);
nor U1180 (N_1180,N_744,N_751);
nand U1181 (N_1181,N_905,N_948);
nor U1182 (N_1182,N_695,N_734);
nor U1183 (N_1183,N_567,N_875);
or U1184 (N_1184,N_800,N_855);
and U1185 (N_1185,N_833,N_997);
nand U1186 (N_1186,N_836,N_952);
or U1187 (N_1187,N_931,N_775);
xnor U1188 (N_1188,N_683,N_724);
and U1189 (N_1189,N_816,N_736);
nor U1190 (N_1190,N_584,N_894);
and U1191 (N_1191,N_677,N_512);
nand U1192 (N_1192,N_622,N_684);
nor U1193 (N_1193,N_714,N_983);
and U1194 (N_1194,N_968,N_648);
nand U1195 (N_1195,N_853,N_604);
or U1196 (N_1196,N_502,N_932);
and U1197 (N_1197,N_614,N_807);
nor U1198 (N_1198,N_590,N_509);
xnor U1199 (N_1199,N_835,N_862);
nor U1200 (N_1200,N_924,N_858);
nor U1201 (N_1201,N_865,N_586);
nand U1202 (N_1202,N_929,N_504);
and U1203 (N_1203,N_675,N_664);
or U1204 (N_1204,N_806,N_523);
nor U1205 (N_1205,N_756,N_752);
and U1206 (N_1206,N_729,N_762);
nor U1207 (N_1207,N_656,N_738);
and U1208 (N_1208,N_516,N_737);
and U1209 (N_1209,N_912,N_640);
nor U1210 (N_1210,N_791,N_712);
or U1211 (N_1211,N_720,N_969);
and U1212 (N_1212,N_967,N_731);
and U1213 (N_1213,N_790,N_972);
nor U1214 (N_1214,N_525,N_661);
nor U1215 (N_1215,N_826,N_700);
nor U1216 (N_1216,N_868,N_542);
and U1217 (N_1217,N_566,N_754);
nand U1218 (N_1218,N_635,N_869);
nor U1219 (N_1219,N_595,N_801);
xor U1220 (N_1220,N_832,N_994);
nor U1221 (N_1221,N_607,N_872);
nor U1222 (N_1222,N_555,N_749);
or U1223 (N_1223,N_609,N_943);
or U1224 (N_1224,N_915,N_902);
nor U1225 (N_1225,N_747,N_975);
nor U1226 (N_1226,N_959,N_808);
and U1227 (N_1227,N_612,N_802);
or U1228 (N_1228,N_687,N_812);
or U1229 (N_1229,N_847,N_739);
nand U1230 (N_1230,N_573,N_991);
and U1231 (N_1231,N_624,N_779);
nand U1232 (N_1232,N_735,N_950);
and U1233 (N_1233,N_580,N_859);
nor U1234 (N_1234,N_996,N_964);
or U1235 (N_1235,N_882,N_639);
or U1236 (N_1236,N_583,N_961);
and U1237 (N_1237,N_817,N_765);
or U1238 (N_1238,N_553,N_978);
nand U1239 (N_1239,N_568,N_513);
nand U1240 (N_1240,N_774,N_511);
nor U1241 (N_1241,N_785,N_863);
and U1242 (N_1242,N_987,N_597);
nand U1243 (N_1243,N_906,N_825);
and U1244 (N_1244,N_815,N_741);
nor U1245 (N_1245,N_842,N_837);
nor U1246 (N_1246,N_632,N_626);
nand U1247 (N_1247,N_522,N_771);
nor U1248 (N_1248,N_998,N_723);
and U1249 (N_1249,N_787,N_898);
nor U1250 (N_1250,N_815,N_738);
nand U1251 (N_1251,N_944,N_935);
or U1252 (N_1252,N_608,N_820);
nor U1253 (N_1253,N_947,N_595);
nand U1254 (N_1254,N_539,N_524);
nand U1255 (N_1255,N_808,N_657);
nand U1256 (N_1256,N_606,N_865);
nand U1257 (N_1257,N_973,N_542);
nor U1258 (N_1258,N_711,N_761);
and U1259 (N_1259,N_972,N_887);
nor U1260 (N_1260,N_807,N_612);
or U1261 (N_1261,N_958,N_646);
nand U1262 (N_1262,N_584,N_557);
or U1263 (N_1263,N_934,N_834);
nor U1264 (N_1264,N_911,N_677);
or U1265 (N_1265,N_868,N_672);
or U1266 (N_1266,N_745,N_800);
or U1267 (N_1267,N_860,N_685);
nand U1268 (N_1268,N_863,N_992);
nor U1269 (N_1269,N_670,N_620);
or U1270 (N_1270,N_521,N_756);
nor U1271 (N_1271,N_727,N_805);
nand U1272 (N_1272,N_957,N_873);
nor U1273 (N_1273,N_840,N_779);
or U1274 (N_1274,N_825,N_845);
nand U1275 (N_1275,N_569,N_883);
and U1276 (N_1276,N_933,N_901);
nand U1277 (N_1277,N_630,N_835);
and U1278 (N_1278,N_912,N_794);
nand U1279 (N_1279,N_874,N_932);
nand U1280 (N_1280,N_760,N_508);
and U1281 (N_1281,N_861,N_953);
or U1282 (N_1282,N_780,N_964);
or U1283 (N_1283,N_970,N_798);
nand U1284 (N_1284,N_747,N_711);
nor U1285 (N_1285,N_696,N_512);
nand U1286 (N_1286,N_772,N_798);
nor U1287 (N_1287,N_903,N_558);
nor U1288 (N_1288,N_558,N_544);
nand U1289 (N_1289,N_852,N_554);
nor U1290 (N_1290,N_682,N_769);
or U1291 (N_1291,N_981,N_657);
nand U1292 (N_1292,N_928,N_860);
and U1293 (N_1293,N_523,N_991);
nor U1294 (N_1294,N_950,N_646);
or U1295 (N_1295,N_693,N_887);
xnor U1296 (N_1296,N_815,N_894);
or U1297 (N_1297,N_914,N_927);
and U1298 (N_1298,N_654,N_825);
nor U1299 (N_1299,N_758,N_699);
and U1300 (N_1300,N_885,N_587);
and U1301 (N_1301,N_542,N_749);
nand U1302 (N_1302,N_918,N_505);
and U1303 (N_1303,N_548,N_663);
nand U1304 (N_1304,N_679,N_823);
xor U1305 (N_1305,N_622,N_692);
or U1306 (N_1306,N_549,N_581);
nor U1307 (N_1307,N_546,N_892);
nand U1308 (N_1308,N_549,N_997);
nand U1309 (N_1309,N_974,N_540);
nand U1310 (N_1310,N_620,N_859);
nand U1311 (N_1311,N_561,N_559);
nor U1312 (N_1312,N_545,N_850);
and U1313 (N_1313,N_986,N_797);
nand U1314 (N_1314,N_757,N_599);
and U1315 (N_1315,N_556,N_972);
nand U1316 (N_1316,N_507,N_982);
or U1317 (N_1317,N_585,N_598);
nand U1318 (N_1318,N_619,N_649);
and U1319 (N_1319,N_867,N_879);
nand U1320 (N_1320,N_540,N_636);
or U1321 (N_1321,N_747,N_870);
nand U1322 (N_1322,N_705,N_638);
or U1323 (N_1323,N_808,N_832);
nor U1324 (N_1324,N_566,N_939);
or U1325 (N_1325,N_725,N_899);
or U1326 (N_1326,N_741,N_689);
or U1327 (N_1327,N_902,N_858);
or U1328 (N_1328,N_735,N_962);
nor U1329 (N_1329,N_691,N_889);
nor U1330 (N_1330,N_970,N_694);
or U1331 (N_1331,N_917,N_542);
nor U1332 (N_1332,N_545,N_768);
or U1333 (N_1333,N_730,N_911);
or U1334 (N_1334,N_979,N_848);
or U1335 (N_1335,N_952,N_780);
nand U1336 (N_1336,N_984,N_897);
nor U1337 (N_1337,N_585,N_648);
or U1338 (N_1338,N_686,N_795);
nor U1339 (N_1339,N_512,N_600);
or U1340 (N_1340,N_944,N_878);
nand U1341 (N_1341,N_663,N_840);
or U1342 (N_1342,N_852,N_535);
nor U1343 (N_1343,N_939,N_978);
or U1344 (N_1344,N_525,N_759);
and U1345 (N_1345,N_569,N_980);
or U1346 (N_1346,N_994,N_742);
or U1347 (N_1347,N_764,N_502);
nor U1348 (N_1348,N_605,N_673);
and U1349 (N_1349,N_817,N_558);
nand U1350 (N_1350,N_570,N_620);
and U1351 (N_1351,N_954,N_809);
or U1352 (N_1352,N_622,N_881);
nor U1353 (N_1353,N_511,N_807);
nor U1354 (N_1354,N_742,N_552);
or U1355 (N_1355,N_926,N_712);
and U1356 (N_1356,N_735,N_560);
nand U1357 (N_1357,N_550,N_615);
nor U1358 (N_1358,N_571,N_718);
nor U1359 (N_1359,N_571,N_900);
or U1360 (N_1360,N_783,N_507);
nor U1361 (N_1361,N_542,N_536);
nor U1362 (N_1362,N_997,N_898);
and U1363 (N_1363,N_541,N_970);
nand U1364 (N_1364,N_877,N_913);
and U1365 (N_1365,N_897,N_801);
and U1366 (N_1366,N_964,N_774);
or U1367 (N_1367,N_644,N_713);
and U1368 (N_1368,N_793,N_535);
nor U1369 (N_1369,N_823,N_872);
nor U1370 (N_1370,N_601,N_503);
nor U1371 (N_1371,N_956,N_550);
nor U1372 (N_1372,N_939,N_832);
and U1373 (N_1373,N_688,N_566);
nand U1374 (N_1374,N_976,N_821);
nand U1375 (N_1375,N_838,N_900);
nand U1376 (N_1376,N_965,N_899);
and U1377 (N_1377,N_778,N_943);
nand U1378 (N_1378,N_799,N_980);
and U1379 (N_1379,N_772,N_762);
nor U1380 (N_1380,N_544,N_710);
nand U1381 (N_1381,N_806,N_905);
nand U1382 (N_1382,N_850,N_732);
or U1383 (N_1383,N_508,N_641);
or U1384 (N_1384,N_721,N_526);
or U1385 (N_1385,N_596,N_540);
nor U1386 (N_1386,N_772,N_953);
nor U1387 (N_1387,N_800,N_645);
nand U1388 (N_1388,N_566,N_515);
nor U1389 (N_1389,N_680,N_650);
nand U1390 (N_1390,N_726,N_611);
nand U1391 (N_1391,N_929,N_597);
nand U1392 (N_1392,N_970,N_521);
nor U1393 (N_1393,N_602,N_570);
nand U1394 (N_1394,N_777,N_591);
nor U1395 (N_1395,N_568,N_875);
or U1396 (N_1396,N_609,N_871);
nor U1397 (N_1397,N_767,N_985);
or U1398 (N_1398,N_855,N_845);
and U1399 (N_1399,N_832,N_838);
or U1400 (N_1400,N_546,N_636);
and U1401 (N_1401,N_953,N_832);
or U1402 (N_1402,N_632,N_542);
nand U1403 (N_1403,N_575,N_930);
nand U1404 (N_1404,N_662,N_599);
nand U1405 (N_1405,N_809,N_609);
and U1406 (N_1406,N_980,N_643);
nor U1407 (N_1407,N_927,N_744);
xor U1408 (N_1408,N_900,N_899);
or U1409 (N_1409,N_764,N_526);
nor U1410 (N_1410,N_679,N_828);
nand U1411 (N_1411,N_662,N_976);
nor U1412 (N_1412,N_567,N_509);
nand U1413 (N_1413,N_986,N_583);
or U1414 (N_1414,N_614,N_831);
nand U1415 (N_1415,N_775,N_552);
or U1416 (N_1416,N_730,N_976);
and U1417 (N_1417,N_549,N_749);
or U1418 (N_1418,N_671,N_914);
nand U1419 (N_1419,N_820,N_999);
or U1420 (N_1420,N_666,N_795);
and U1421 (N_1421,N_584,N_966);
and U1422 (N_1422,N_867,N_572);
and U1423 (N_1423,N_635,N_632);
nor U1424 (N_1424,N_673,N_692);
nor U1425 (N_1425,N_833,N_508);
nand U1426 (N_1426,N_841,N_942);
and U1427 (N_1427,N_961,N_645);
nor U1428 (N_1428,N_560,N_547);
or U1429 (N_1429,N_585,N_532);
nor U1430 (N_1430,N_881,N_819);
nand U1431 (N_1431,N_857,N_513);
and U1432 (N_1432,N_922,N_646);
nand U1433 (N_1433,N_810,N_684);
or U1434 (N_1434,N_733,N_570);
nand U1435 (N_1435,N_594,N_530);
or U1436 (N_1436,N_587,N_524);
or U1437 (N_1437,N_569,N_585);
nand U1438 (N_1438,N_723,N_515);
and U1439 (N_1439,N_565,N_689);
or U1440 (N_1440,N_602,N_668);
nand U1441 (N_1441,N_850,N_897);
nor U1442 (N_1442,N_772,N_889);
or U1443 (N_1443,N_935,N_575);
and U1444 (N_1444,N_866,N_711);
nand U1445 (N_1445,N_950,N_621);
nor U1446 (N_1446,N_898,N_768);
and U1447 (N_1447,N_610,N_706);
or U1448 (N_1448,N_646,N_517);
nand U1449 (N_1449,N_616,N_915);
nor U1450 (N_1450,N_888,N_940);
and U1451 (N_1451,N_699,N_666);
nand U1452 (N_1452,N_821,N_828);
nor U1453 (N_1453,N_503,N_592);
and U1454 (N_1454,N_842,N_510);
and U1455 (N_1455,N_789,N_799);
and U1456 (N_1456,N_757,N_586);
or U1457 (N_1457,N_763,N_585);
nor U1458 (N_1458,N_738,N_530);
or U1459 (N_1459,N_981,N_758);
nor U1460 (N_1460,N_602,N_789);
nor U1461 (N_1461,N_933,N_947);
and U1462 (N_1462,N_521,N_872);
or U1463 (N_1463,N_538,N_988);
nor U1464 (N_1464,N_993,N_531);
and U1465 (N_1465,N_784,N_798);
nand U1466 (N_1466,N_951,N_875);
and U1467 (N_1467,N_896,N_555);
nor U1468 (N_1468,N_703,N_833);
and U1469 (N_1469,N_713,N_564);
and U1470 (N_1470,N_916,N_539);
nand U1471 (N_1471,N_927,N_776);
and U1472 (N_1472,N_797,N_925);
nor U1473 (N_1473,N_652,N_758);
and U1474 (N_1474,N_642,N_691);
nand U1475 (N_1475,N_968,N_574);
or U1476 (N_1476,N_640,N_846);
nor U1477 (N_1477,N_733,N_731);
nor U1478 (N_1478,N_675,N_837);
or U1479 (N_1479,N_515,N_910);
or U1480 (N_1480,N_588,N_784);
nand U1481 (N_1481,N_516,N_974);
nor U1482 (N_1482,N_504,N_937);
nor U1483 (N_1483,N_518,N_585);
nor U1484 (N_1484,N_576,N_683);
nand U1485 (N_1485,N_590,N_925);
and U1486 (N_1486,N_885,N_692);
or U1487 (N_1487,N_768,N_543);
or U1488 (N_1488,N_839,N_811);
nand U1489 (N_1489,N_655,N_956);
nand U1490 (N_1490,N_975,N_606);
and U1491 (N_1491,N_976,N_553);
nand U1492 (N_1492,N_758,N_946);
nand U1493 (N_1493,N_736,N_580);
nand U1494 (N_1494,N_780,N_800);
and U1495 (N_1495,N_655,N_864);
and U1496 (N_1496,N_987,N_897);
nor U1497 (N_1497,N_593,N_841);
or U1498 (N_1498,N_949,N_725);
nor U1499 (N_1499,N_998,N_806);
or U1500 (N_1500,N_1234,N_1405);
nand U1501 (N_1501,N_1394,N_1002);
or U1502 (N_1502,N_1153,N_1077);
nor U1503 (N_1503,N_1458,N_1158);
and U1504 (N_1504,N_1066,N_1028);
or U1505 (N_1505,N_1436,N_1197);
nand U1506 (N_1506,N_1376,N_1316);
nand U1507 (N_1507,N_1265,N_1274);
and U1508 (N_1508,N_1457,N_1352);
and U1509 (N_1509,N_1312,N_1406);
nor U1510 (N_1510,N_1164,N_1085);
nor U1511 (N_1511,N_1160,N_1184);
or U1512 (N_1512,N_1128,N_1208);
nand U1513 (N_1513,N_1313,N_1178);
and U1514 (N_1514,N_1303,N_1020);
and U1515 (N_1515,N_1472,N_1180);
and U1516 (N_1516,N_1110,N_1431);
nor U1517 (N_1517,N_1395,N_1356);
or U1518 (N_1518,N_1209,N_1256);
nor U1519 (N_1519,N_1091,N_1491);
or U1520 (N_1520,N_1157,N_1022);
or U1521 (N_1521,N_1404,N_1133);
nand U1522 (N_1522,N_1040,N_1246);
nand U1523 (N_1523,N_1034,N_1493);
or U1524 (N_1524,N_1042,N_1068);
nand U1525 (N_1525,N_1206,N_1433);
or U1526 (N_1526,N_1357,N_1452);
and U1527 (N_1527,N_1203,N_1414);
and U1528 (N_1528,N_1266,N_1241);
nand U1529 (N_1529,N_1338,N_1318);
nor U1530 (N_1530,N_1393,N_1127);
nand U1531 (N_1531,N_1039,N_1400);
and U1532 (N_1532,N_1396,N_1044);
or U1533 (N_1533,N_1378,N_1314);
nor U1534 (N_1534,N_1479,N_1169);
or U1535 (N_1535,N_1451,N_1262);
nor U1536 (N_1536,N_1407,N_1024);
nor U1537 (N_1537,N_1337,N_1415);
or U1538 (N_1538,N_1089,N_1079);
nor U1539 (N_1539,N_1432,N_1186);
and U1540 (N_1540,N_1008,N_1289);
or U1541 (N_1541,N_1456,N_1345);
and U1542 (N_1542,N_1271,N_1492);
or U1543 (N_1543,N_1360,N_1224);
or U1544 (N_1544,N_1446,N_1001);
and U1545 (N_1545,N_1300,N_1087);
nor U1546 (N_1546,N_1263,N_1238);
and U1547 (N_1547,N_1216,N_1166);
nand U1548 (N_1548,N_1041,N_1468);
and U1549 (N_1549,N_1424,N_1278);
nand U1550 (N_1550,N_1134,N_1410);
nor U1551 (N_1551,N_1305,N_1346);
and U1552 (N_1552,N_1107,N_1189);
and U1553 (N_1553,N_1444,N_1130);
and U1554 (N_1554,N_1227,N_1143);
or U1555 (N_1555,N_1385,N_1140);
nor U1556 (N_1556,N_1488,N_1299);
or U1557 (N_1557,N_1397,N_1429);
nand U1558 (N_1558,N_1200,N_1382);
nand U1559 (N_1559,N_1082,N_1236);
nor U1560 (N_1560,N_1102,N_1188);
nand U1561 (N_1561,N_1269,N_1247);
nand U1562 (N_1562,N_1273,N_1230);
nand U1563 (N_1563,N_1170,N_1076);
nand U1564 (N_1564,N_1416,N_1417);
nand U1565 (N_1565,N_1389,N_1288);
nand U1566 (N_1566,N_1375,N_1471);
and U1567 (N_1567,N_1245,N_1442);
or U1568 (N_1568,N_1137,N_1330);
and U1569 (N_1569,N_1267,N_1162);
or U1570 (N_1570,N_1086,N_1254);
nand U1571 (N_1571,N_1408,N_1398);
and U1572 (N_1572,N_1161,N_1075);
nor U1573 (N_1573,N_1402,N_1467);
nand U1574 (N_1574,N_1048,N_1094);
or U1575 (N_1575,N_1013,N_1210);
nor U1576 (N_1576,N_1469,N_1235);
and U1577 (N_1577,N_1369,N_1276);
nor U1578 (N_1578,N_1486,N_1191);
and U1579 (N_1579,N_1012,N_1005);
or U1580 (N_1580,N_1037,N_1030);
and U1581 (N_1581,N_1117,N_1006);
or U1582 (N_1582,N_1251,N_1481);
nor U1583 (N_1583,N_1201,N_1449);
or U1584 (N_1584,N_1126,N_1152);
or U1585 (N_1585,N_1100,N_1344);
nand U1586 (N_1586,N_1131,N_1232);
nor U1587 (N_1587,N_1093,N_1035);
or U1588 (N_1588,N_1302,N_1307);
nor U1589 (N_1589,N_1466,N_1092);
or U1590 (N_1590,N_1196,N_1242);
nand U1591 (N_1591,N_1215,N_1124);
and U1592 (N_1592,N_1199,N_1147);
and U1593 (N_1593,N_1325,N_1074);
xnor U1594 (N_1594,N_1290,N_1220);
or U1595 (N_1595,N_1212,N_1448);
and U1596 (N_1596,N_1115,N_1195);
nor U1597 (N_1597,N_1401,N_1061);
or U1598 (N_1598,N_1310,N_1261);
nand U1599 (N_1599,N_1171,N_1248);
nor U1600 (N_1600,N_1150,N_1237);
or U1601 (N_1601,N_1440,N_1244);
and U1602 (N_1602,N_1049,N_1328);
and U1603 (N_1603,N_1098,N_1004);
and U1604 (N_1604,N_1309,N_1175);
or U1605 (N_1605,N_1000,N_1460);
or U1606 (N_1606,N_1045,N_1239);
and U1607 (N_1607,N_1252,N_1461);
nor U1608 (N_1608,N_1319,N_1478);
and U1609 (N_1609,N_1023,N_1168);
and U1610 (N_1610,N_1067,N_1327);
nand U1611 (N_1611,N_1340,N_1294);
nand U1612 (N_1612,N_1057,N_1361);
or U1613 (N_1613,N_1109,N_1194);
and U1614 (N_1614,N_1351,N_1202);
nand U1615 (N_1615,N_1050,N_1112);
or U1616 (N_1616,N_1167,N_1282);
and U1617 (N_1617,N_1439,N_1308);
nor U1618 (N_1618,N_1179,N_1285);
nand U1619 (N_1619,N_1193,N_1497);
nor U1620 (N_1620,N_1487,N_1499);
nor U1621 (N_1621,N_1476,N_1443);
or U1622 (N_1622,N_1151,N_1033);
nor U1623 (N_1623,N_1441,N_1253);
and U1624 (N_1624,N_1297,N_1214);
nand U1625 (N_1625,N_1296,N_1025);
nand U1626 (N_1626,N_1059,N_1229);
nand U1627 (N_1627,N_1103,N_1058);
and U1628 (N_1628,N_1428,N_1384);
or U1629 (N_1629,N_1258,N_1324);
or U1630 (N_1630,N_1007,N_1386);
nor U1631 (N_1631,N_1146,N_1380);
and U1632 (N_1632,N_1069,N_1104);
nor U1633 (N_1633,N_1010,N_1226);
or U1634 (N_1634,N_1187,N_1029);
and U1635 (N_1635,N_1217,N_1342);
and U1636 (N_1636,N_1459,N_1081);
or U1637 (N_1637,N_1257,N_1122);
nand U1638 (N_1638,N_1304,N_1490);
nand U1639 (N_1639,N_1264,N_1225);
or U1640 (N_1640,N_1176,N_1015);
nor U1641 (N_1641,N_1207,N_1331);
nand U1642 (N_1642,N_1099,N_1463);
nand U1643 (N_1643,N_1095,N_1329);
and U1644 (N_1644,N_1036,N_1121);
or U1645 (N_1645,N_1326,N_1475);
or U1646 (N_1646,N_1341,N_1155);
nor U1647 (N_1647,N_1047,N_1072);
and U1648 (N_1648,N_1306,N_1280);
nor U1649 (N_1649,N_1465,N_1392);
nand U1650 (N_1650,N_1489,N_1419);
nand U1651 (N_1651,N_1343,N_1359);
nand U1652 (N_1652,N_1371,N_1019);
nor U1653 (N_1653,N_1445,N_1368);
or U1654 (N_1654,N_1473,N_1333);
or U1655 (N_1655,N_1367,N_1347);
nor U1656 (N_1656,N_1470,N_1183);
or U1657 (N_1657,N_1144,N_1383);
or U1658 (N_1658,N_1348,N_1277);
or U1659 (N_1659,N_1477,N_1139);
nand U1660 (N_1660,N_1495,N_1374);
or U1661 (N_1661,N_1064,N_1260);
nor U1662 (N_1662,N_1355,N_1283);
nand U1663 (N_1663,N_1218,N_1287);
and U1664 (N_1664,N_1223,N_1125);
nor U1665 (N_1665,N_1450,N_1435);
or U1666 (N_1666,N_1185,N_1250);
or U1667 (N_1667,N_1113,N_1339);
nor U1668 (N_1668,N_1377,N_1447);
nand U1669 (N_1669,N_1159,N_1420);
nor U1670 (N_1670,N_1181,N_1026);
or U1671 (N_1671,N_1454,N_1101);
or U1672 (N_1672,N_1106,N_1156);
and U1673 (N_1673,N_1221,N_1228);
and U1674 (N_1674,N_1480,N_1320);
or U1675 (N_1675,N_1363,N_1334);
nor U1676 (N_1676,N_1390,N_1434);
or U1677 (N_1677,N_1043,N_1198);
and U1678 (N_1678,N_1027,N_1123);
or U1679 (N_1679,N_1425,N_1118);
and U1680 (N_1680,N_1354,N_1174);
nor U1681 (N_1681,N_1135,N_1083);
nor U1682 (N_1682,N_1409,N_1494);
and U1683 (N_1683,N_1243,N_1272);
nand U1684 (N_1684,N_1323,N_1060);
or U1685 (N_1685,N_1119,N_1009);
and U1686 (N_1686,N_1284,N_1381);
nand U1687 (N_1687,N_1213,N_1054);
and U1688 (N_1688,N_1279,N_1053);
and U1689 (N_1689,N_1423,N_1293);
nand U1690 (N_1690,N_1301,N_1172);
nor U1691 (N_1691,N_1090,N_1496);
and U1692 (N_1692,N_1014,N_1016);
and U1693 (N_1693,N_1182,N_1038);
nand U1694 (N_1694,N_1173,N_1364);
or U1695 (N_1695,N_1281,N_1298);
nor U1696 (N_1696,N_1219,N_1154);
and U1697 (N_1697,N_1056,N_1474);
nand U1698 (N_1698,N_1138,N_1295);
nand U1699 (N_1699,N_1464,N_1192);
and U1700 (N_1700,N_1379,N_1455);
xnor U1701 (N_1701,N_1096,N_1268);
and U1702 (N_1702,N_1055,N_1063);
and U1703 (N_1703,N_1391,N_1165);
nor U1704 (N_1704,N_1366,N_1141);
nor U1705 (N_1705,N_1412,N_1205);
nor U1706 (N_1706,N_1108,N_1011);
nor U1707 (N_1707,N_1421,N_1498);
nand U1708 (N_1708,N_1211,N_1116);
nor U1709 (N_1709,N_1422,N_1003);
and U1710 (N_1710,N_1105,N_1021);
or U1711 (N_1711,N_1438,N_1413);
nand U1712 (N_1712,N_1411,N_1046);
and U1713 (N_1713,N_1372,N_1259);
or U1714 (N_1714,N_1204,N_1084);
and U1715 (N_1715,N_1070,N_1336);
or U1716 (N_1716,N_1163,N_1145);
or U1717 (N_1717,N_1051,N_1142);
nand U1718 (N_1718,N_1317,N_1071);
nor U1719 (N_1719,N_1291,N_1177);
or U1720 (N_1720,N_1233,N_1418);
and U1721 (N_1721,N_1315,N_1031);
or U1722 (N_1722,N_1190,N_1018);
or U1723 (N_1723,N_1335,N_1132);
nor U1724 (N_1724,N_1097,N_1311);
and U1725 (N_1725,N_1275,N_1353);
and U1726 (N_1726,N_1358,N_1365);
or U1727 (N_1727,N_1111,N_1149);
nand U1728 (N_1728,N_1052,N_1332);
or U1729 (N_1729,N_1350,N_1482);
or U1730 (N_1730,N_1120,N_1483);
and U1731 (N_1731,N_1032,N_1255);
nand U1732 (N_1732,N_1129,N_1437);
or U1733 (N_1733,N_1362,N_1322);
or U1734 (N_1734,N_1292,N_1062);
or U1735 (N_1735,N_1484,N_1321);
nand U1736 (N_1736,N_1430,N_1249);
or U1737 (N_1737,N_1017,N_1080);
or U1738 (N_1738,N_1240,N_1427);
and U1739 (N_1739,N_1073,N_1078);
nand U1740 (N_1740,N_1222,N_1370);
nand U1741 (N_1741,N_1373,N_1231);
nand U1742 (N_1742,N_1462,N_1399);
and U1743 (N_1743,N_1114,N_1388);
or U1744 (N_1744,N_1148,N_1349);
nor U1745 (N_1745,N_1387,N_1270);
nand U1746 (N_1746,N_1065,N_1453);
and U1747 (N_1747,N_1426,N_1485);
nor U1748 (N_1748,N_1403,N_1136);
and U1749 (N_1749,N_1286,N_1088);
or U1750 (N_1750,N_1174,N_1477);
and U1751 (N_1751,N_1007,N_1274);
and U1752 (N_1752,N_1341,N_1103);
and U1753 (N_1753,N_1406,N_1126);
xor U1754 (N_1754,N_1072,N_1014);
nand U1755 (N_1755,N_1483,N_1480);
nor U1756 (N_1756,N_1092,N_1064);
or U1757 (N_1757,N_1325,N_1102);
nand U1758 (N_1758,N_1184,N_1429);
nor U1759 (N_1759,N_1152,N_1401);
and U1760 (N_1760,N_1022,N_1061);
nor U1761 (N_1761,N_1121,N_1065);
or U1762 (N_1762,N_1264,N_1305);
or U1763 (N_1763,N_1164,N_1358);
or U1764 (N_1764,N_1060,N_1422);
nand U1765 (N_1765,N_1358,N_1298);
or U1766 (N_1766,N_1449,N_1358);
and U1767 (N_1767,N_1093,N_1393);
nor U1768 (N_1768,N_1409,N_1417);
nand U1769 (N_1769,N_1116,N_1263);
or U1770 (N_1770,N_1138,N_1427);
nand U1771 (N_1771,N_1358,N_1156);
or U1772 (N_1772,N_1408,N_1385);
nand U1773 (N_1773,N_1129,N_1435);
and U1774 (N_1774,N_1428,N_1345);
nand U1775 (N_1775,N_1189,N_1191);
nand U1776 (N_1776,N_1207,N_1082);
nand U1777 (N_1777,N_1068,N_1024);
or U1778 (N_1778,N_1403,N_1228);
and U1779 (N_1779,N_1144,N_1058);
nor U1780 (N_1780,N_1236,N_1320);
or U1781 (N_1781,N_1410,N_1209);
or U1782 (N_1782,N_1184,N_1409);
and U1783 (N_1783,N_1017,N_1058);
nor U1784 (N_1784,N_1074,N_1062);
nand U1785 (N_1785,N_1332,N_1494);
nand U1786 (N_1786,N_1035,N_1410);
nor U1787 (N_1787,N_1030,N_1070);
nand U1788 (N_1788,N_1203,N_1032);
or U1789 (N_1789,N_1424,N_1005);
nor U1790 (N_1790,N_1072,N_1181);
and U1791 (N_1791,N_1468,N_1126);
nand U1792 (N_1792,N_1024,N_1385);
or U1793 (N_1793,N_1468,N_1332);
and U1794 (N_1794,N_1048,N_1434);
and U1795 (N_1795,N_1257,N_1031);
nor U1796 (N_1796,N_1090,N_1139);
or U1797 (N_1797,N_1200,N_1036);
nand U1798 (N_1798,N_1051,N_1031);
and U1799 (N_1799,N_1204,N_1285);
or U1800 (N_1800,N_1094,N_1126);
nand U1801 (N_1801,N_1417,N_1308);
or U1802 (N_1802,N_1278,N_1165);
nand U1803 (N_1803,N_1396,N_1108);
nor U1804 (N_1804,N_1324,N_1189);
or U1805 (N_1805,N_1027,N_1112);
and U1806 (N_1806,N_1076,N_1055);
nor U1807 (N_1807,N_1224,N_1315);
and U1808 (N_1808,N_1212,N_1198);
xnor U1809 (N_1809,N_1332,N_1116);
or U1810 (N_1810,N_1307,N_1346);
and U1811 (N_1811,N_1372,N_1174);
and U1812 (N_1812,N_1409,N_1044);
nor U1813 (N_1813,N_1270,N_1157);
nor U1814 (N_1814,N_1330,N_1356);
and U1815 (N_1815,N_1491,N_1439);
or U1816 (N_1816,N_1113,N_1185);
nor U1817 (N_1817,N_1410,N_1173);
nand U1818 (N_1818,N_1437,N_1197);
nand U1819 (N_1819,N_1191,N_1012);
nor U1820 (N_1820,N_1444,N_1004);
nand U1821 (N_1821,N_1414,N_1273);
and U1822 (N_1822,N_1477,N_1314);
and U1823 (N_1823,N_1263,N_1081);
nand U1824 (N_1824,N_1305,N_1106);
nand U1825 (N_1825,N_1116,N_1342);
nand U1826 (N_1826,N_1266,N_1360);
nand U1827 (N_1827,N_1407,N_1109);
nand U1828 (N_1828,N_1325,N_1208);
or U1829 (N_1829,N_1345,N_1196);
nor U1830 (N_1830,N_1466,N_1341);
nand U1831 (N_1831,N_1250,N_1262);
nand U1832 (N_1832,N_1322,N_1403);
nor U1833 (N_1833,N_1319,N_1477);
nor U1834 (N_1834,N_1489,N_1315);
nor U1835 (N_1835,N_1299,N_1351);
nor U1836 (N_1836,N_1367,N_1440);
xnor U1837 (N_1837,N_1062,N_1042);
nor U1838 (N_1838,N_1372,N_1162);
and U1839 (N_1839,N_1096,N_1250);
and U1840 (N_1840,N_1028,N_1396);
nor U1841 (N_1841,N_1272,N_1332);
or U1842 (N_1842,N_1034,N_1482);
nor U1843 (N_1843,N_1442,N_1432);
or U1844 (N_1844,N_1435,N_1415);
or U1845 (N_1845,N_1153,N_1208);
and U1846 (N_1846,N_1358,N_1217);
nor U1847 (N_1847,N_1350,N_1139);
or U1848 (N_1848,N_1309,N_1167);
nor U1849 (N_1849,N_1421,N_1048);
and U1850 (N_1850,N_1295,N_1003);
nand U1851 (N_1851,N_1180,N_1009);
or U1852 (N_1852,N_1053,N_1366);
and U1853 (N_1853,N_1482,N_1093);
nand U1854 (N_1854,N_1040,N_1471);
nor U1855 (N_1855,N_1142,N_1429);
nor U1856 (N_1856,N_1136,N_1205);
and U1857 (N_1857,N_1333,N_1089);
nand U1858 (N_1858,N_1157,N_1351);
nand U1859 (N_1859,N_1481,N_1495);
nor U1860 (N_1860,N_1449,N_1307);
nor U1861 (N_1861,N_1483,N_1347);
or U1862 (N_1862,N_1357,N_1369);
nand U1863 (N_1863,N_1353,N_1315);
and U1864 (N_1864,N_1346,N_1284);
and U1865 (N_1865,N_1387,N_1182);
nand U1866 (N_1866,N_1232,N_1186);
and U1867 (N_1867,N_1226,N_1472);
and U1868 (N_1868,N_1281,N_1243);
nor U1869 (N_1869,N_1465,N_1399);
or U1870 (N_1870,N_1414,N_1432);
nand U1871 (N_1871,N_1472,N_1432);
nor U1872 (N_1872,N_1348,N_1095);
nor U1873 (N_1873,N_1011,N_1126);
and U1874 (N_1874,N_1048,N_1309);
nor U1875 (N_1875,N_1294,N_1299);
nor U1876 (N_1876,N_1254,N_1089);
nand U1877 (N_1877,N_1062,N_1309);
and U1878 (N_1878,N_1300,N_1349);
or U1879 (N_1879,N_1080,N_1040);
nor U1880 (N_1880,N_1057,N_1282);
nor U1881 (N_1881,N_1282,N_1496);
or U1882 (N_1882,N_1364,N_1019);
nand U1883 (N_1883,N_1084,N_1450);
nand U1884 (N_1884,N_1453,N_1083);
and U1885 (N_1885,N_1251,N_1001);
nand U1886 (N_1886,N_1319,N_1230);
nor U1887 (N_1887,N_1018,N_1061);
nand U1888 (N_1888,N_1351,N_1162);
or U1889 (N_1889,N_1003,N_1093);
and U1890 (N_1890,N_1396,N_1477);
or U1891 (N_1891,N_1151,N_1352);
or U1892 (N_1892,N_1357,N_1370);
or U1893 (N_1893,N_1227,N_1074);
or U1894 (N_1894,N_1208,N_1022);
and U1895 (N_1895,N_1053,N_1392);
nor U1896 (N_1896,N_1350,N_1245);
and U1897 (N_1897,N_1333,N_1160);
nand U1898 (N_1898,N_1317,N_1231);
nand U1899 (N_1899,N_1188,N_1338);
and U1900 (N_1900,N_1328,N_1400);
nand U1901 (N_1901,N_1275,N_1473);
nor U1902 (N_1902,N_1416,N_1117);
or U1903 (N_1903,N_1041,N_1213);
or U1904 (N_1904,N_1160,N_1477);
or U1905 (N_1905,N_1109,N_1477);
and U1906 (N_1906,N_1000,N_1149);
and U1907 (N_1907,N_1174,N_1082);
nor U1908 (N_1908,N_1018,N_1129);
nand U1909 (N_1909,N_1144,N_1387);
nand U1910 (N_1910,N_1369,N_1355);
or U1911 (N_1911,N_1022,N_1265);
or U1912 (N_1912,N_1255,N_1454);
and U1913 (N_1913,N_1336,N_1496);
nor U1914 (N_1914,N_1241,N_1434);
nand U1915 (N_1915,N_1066,N_1057);
and U1916 (N_1916,N_1231,N_1388);
or U1917 (N_1917,N_1488,N_1268);
nor U1918 (N_1918,N_1080,N_1424);
or U1919 (N_1919,N_1335,N_1290);
nand U1920 (N_1920,N_1041,N_1249);
and U1921 (N_1921,N_1002,N_1177);
nand U1922 (N_1922,N_1437,N_1158);
or U1923 (N_1923,N_1476,N_1315);
and U1924 (N_1924,N_1044,N_1113);
nor U1925 (N_1925,N_1097,N_1308);
nor U1926 (N_1926,N_1070,N_1270);
nor U1927 (N_1927,N_1452,N_1490);
and U1928 (N_1928,N_1146,N_1454);
and U1929 (N_1929,N_1417,N_1433);
nor U1930 (N_1930,N_1442,N_1162);
and U1931 (N_1931,N_1355,N_1271);
or U1932 (N_1932,N_1224,N_1120);
nor U1933 (N_1933,N_1249,N_1242);
nor U1934 (N_1934,N_1121,N_1027);
nand U1935 (N_1935,N_1422,N_1491);
nor U1936 (N_1936,N_1037,N_1398);
or U1937 (N_1937,N_1143,N_1315);
and U1938 (N_1938,N_1454,N_1290);
nor U1939 (N_1939,N_1283,N_1322);
and U1940 (N_1940,N_1302,N_1448);
nor U1941 (N_1941,N_1242,N_1080);
and U1942 (N_1942,N_1063,N_1053);
or U1943 (N_1943,N_1496,N_1018);
nor U1944 (N_1944,N_1330,N_1205);
nand U1945 (N_1945,N_1305,N_1061);
and U1946 (N_1946,N_1145,N_1400);
and U1947 (N_1947,N_1323,N_1358);
and U1948 (N_1948,N_1243,N_1169);
or U1949 (N_1949,N_1497,N_1152);
and U1950 (N_1950,N_1034,N_1231);
and U1951 (N_1951,N_1061,N_1089);
nor U1952 (N_1952,N_1234,N_1459);
and U1953 (N_1953,N_1280,N_1344);
nor U1954 (N_1954,N_1027,N_1089);
and U1955 (N_1955,N_1150,N_1059);
or U1956 (N_1956,N_1295,N_1304);
and U1957 (N_1957,N_1373,N_1255);
nor U1958 (N_1958,N_1472,N_1423);
or U1959 (N_1959,N_1322,N_1223);
and U1960 (N_1960,N_1386,N_1288);
and U1961 (N_1961,N_1381,N_1289);
or U1962 (N_1962,N_1160,N_1353);
and U1963 (N_1963,N_1208,N_1264);
nand U1964 (N_1964,N_1453,N_1294);
nand U1965 (N_1965,N_1326,N_1458);
nor U1966 (N_1966,N_1089,N_1038);
nor U1967 (N_1967,N_1323,N_1185);
and U1968 (N_1968,N_1436,N_1455);
or U1969 (N_1969,N_1181,N_1369);
nand U1970 (N_1970,N_1056,N_1164);
nand U1971 (N_1971,N_1171,N_1393);
nor U1972 (N_1972,N_1243,N_1323);
nor U1973 (N_1973,N_1482,N_1238);
nor U1974 (N_1974,N_1048,N_1465);
or U1975 (N_1975,N_1135,N_1428);
nand U1976 (N_1976,N_1388,N_1323);
xor U1977 (N_1977,N_1264,N_1016);
and U1978 (N_1978,N_1445,N_1248);
nor U1979 (N_1979,N_1422,N_1135);
and U1980 (N_1980,N_1426,N_1148);
nor U1981 (N_1981,N_1367,N_1445);
or U1982 (N_1982,N_1433,N_1015);
nor U1983 (N_1983,N_1173,N_1284);
or U1984 (N_1984,N_1107,N_1078);
nor U1985 (N_1985,N_1347,N_1475);
or U1986 (N_1986,N_1216,N_1041);
and U1987 (N_1987,N_1193,N_1205);
nor U1988 (N_1988,N_1333,N_1364);
and U1989 (N_1989,N_1248,N_1176);
or U1990 (N_1990,N_1063,N_1431);
nand U1991 (N_1991,N_1499,N_1338);
nand U1992 (N_1992,N_1210,N_1036);
nand U1993 (N_1993,N_1162,N_1125);
nand U1994 (N_1994,N_1083,N_1464);
nor U1995 (N_1995,N_1460,N_1333);
or U1996 (N_1996,N_1052,N_1044);
nand U1997 (N_1997,N_1110,N_1182);
nand U1998 (N_1998,N_1201,N_1117);
and U1999 (N_1999,N_1433,N_1475);
nor U2000 (N_2000,N_1781,N_1511);
and U2001 (N_2001,N_1973,N_1977);
and U2002 (N_2002,N_1642,N_1840);
nor U2003 (N_2003,N_1917,N_1676);
or U2004 (N_2004,N_1925,N_1600);
or U2005 (N_2005,N_1724,N_1556);
or U2006 (N_2006,N_1660,N_1830);
nand U2007 (N_2007,N_1786,N_1992);
or U2008 (N_2008,N_1738,N_1718);
or U2009 (N_2009,N_1613,N_1650);
and U2010 (N_2010,N_1929,N_1606);
nor U2011 (N_2011,N_1548,N_1599);
nand U2012 (N_2012,N_1741,N_1959);
nand U2013 (N_2013,N_1557,N_1501);
or U2014 (N_2014,N_1554,N_1566);
or U2015 (N_2015,N_1631,N_1920);
nor U2016 (N_2016,N_1957,N_1540);
nor U2017 (N_2017,N_1697,N_1839);
nor U2018 (N_2018,N_1657,N_1536);
nor U2019 (N_2019,N_1698,N_1691);
and U2020 (N_2020,N_1968,N_1755);
and U2021 (N_2021,N_1869,N_1623);
nand U2022 (N_2022,N_1928,N_1774);
and U2023 (N_2023,N_1727,N_1616);
nand U2024 (N_2024,N_1822,N_1763);
nand U2025 (N_2025,N_1687,N_1885);
or U2026 (N_2026,N_1978,N_1633);
nand U2027 (N_2027,N_1500,N_1998);
nor U2028 (N_2028,N_1710,N_1761);
nor U2029 (N_2029,N_1884,N_1926);
or U2030 (N_2030,N_1862,N_1739);
or U2031 (N_2031,N_1700,N_1817);
nand U2032 (N_2032,N_1812,N_1612);
and U2033 (N_2033,N_1652,N_1983);
and U2034 (N_2034,N_1578,N_1630);
and U2035 (N_2035,N_1668,N_1894);
nand U2036 (N_2036,N_1619,N_1605);
or U2037 (N_2037,N_1598,N_1748);
or U2038 (N_2038,N_1561,N_1962);
or U2039 (N_2039,N_1503,N_1914);
nand U2040 (N_2040,N_1510,N_1584);
and U2041 (N_2041,N_1726,N_1728);
xnor U2042 (N_2042,N_1916,N_1678);
or U2043 (N_2043,N_1883,N_1931);
nor U2044 (N_2044,N_1994,N_1997);
nor U2045 (N_2045,N_1861,N_1634);
and U2046 (N_2046,N_1614,N_1843);
xor U2047 (N_2047,N_1942,N_1859);
nand U2048 (N_2048,N_1641,N_1952);
or U2049 (N_2049,N_1541,N_1620);
nor U2050 (N_2050,N_1841,N_1800);
nor U2051 (N_2051,N_1853,N_1525);
and U2052 (N_2052,N_1629,N_1564);
nand U2053 (N_2053,N_1826,N_1856);
or U2054 (N_2054,N_1984,N_1672);
and U2055 (N_2055,N_1995,N_1581);
nand U2056 (N_2056,N_1801,N_1814);
and U2057 (N_2057,N_1508,N_1517);
and U2058 (N_2058,N_1744,N_1935);
and U2059 (N_2059,N_1574,N_1535);
and U2060 (N_2060,N_1610,N_1794);
nand U2061 (N_2061,N_1745,N_1523);
nor U2062 (N_2062,N_1910,N_1505);
nand U2063 (N_2063,N_1834,N_1770);
and U2064 (N_2064,N_1866,N_1733);
nand U2065 (N_2065,N_1778,N_1988);
or U2066 (N_2066,N_1956,N_1887);
and U2067 (N_2067,N_1751,N_1563);
nand U2068 (N_2068,N_1756,N_1646);
and U2069 (N_2069,N_1663,N_1787);
or U2070 (N_2070,N_1680,N_1527);
nor U2071 (N_2071,N_1732,N_1767);
nand U2072 (N_2072,N_1922,N_1526);
nor U2073 (N_2073,N_1793,N_1902);
and U2074 (N_2074,N_1693,N_1873);
nor U2075 (N_2075,N_1520,N_1851);
nor U2076 (N_2076,N_1542,N_1864);
nand U2077 (N_2077,N_1719,N_1655);
and U2078 (N_2078,N_1569,N_1836);
and U2079 (N_2079,N_1624,N_1838);
and U2080 (N_2080,N_1950,N_1980);
and U2081 (N_2081,N_1833,N_1971);
nand U2082 (N_2082,N_1701,N_1626);
and U2083 (N_2083,N_1588,N_1848);
nand U2084 (N_2084,N_1712,N_1986);
nor U2085 (N_2085,N_1709,N_1516);
nand U2086 (N_2086,N_1627,N_1722);
and U2087 (N_2087,N_1919,N_1683);
nand U2088 (N_2088,N_1878,N_1832);
nand U2089 (N_2089,N_1937,N_1562);
and U2090 (N_2090,N_1538,N_1515);
and U2091 (N_2091,N_1820,N_1549);
and U2092 (N_2092,N_1965,N_1954);
nor U2093 (N_2093,N_1559,N_1669);
and U2094 (N_2094,N_1593,N_1675);
nor U2095 (N_2095,N_1874,N_1784);
nand U2096 (N_2096,N_1580,N_1647);
and U2097 (N_2097,N_1775,N_1876);
and U2098 (N_2098,N_1529,N_1713);
or U2099 (N_2099,N_1604,N_1560);
nor U2100 (N_2100,N_1742,N_1509);
nand U2101 (N_2101,N_1813,N_1597);
nand U2102 (N_2102,N_1696,N_1837);
nor U2103 (N_2103,N_1790,N_1880);
nand U2104 (N_2104,N_1805,N_1753);
and U2105 (N_2105,N_1844,N_1939);
or U2106 (N_2106,N_1512,N_1818);
or U2107 (N_2107,N_1684,N_1667);
nand U2108 (N_2108,N_1618,N_1651);
nand U2109 (N_2109,N_1904,N_1632);
or U2110 (N_2110,N_1653,N_1783);
nand U2111 (N_2111,N_1737,N_1635);
nand U2112 (N_2112,N_1544,N_1644);
nor U2113 (N_2113,N_1847,N_1567);
or U2114 (N_2114,N_1649,N_1764);
and U2115 (N_2115,N_1821,N_1846);
nand U2116 (N_2116,N_1682,N_1735);
and U2117 (N_2117,N_1802,N_1565);
and U2118 (N_2118,N_1879,N_1587);
nor U2119 (N_2119,N_1865,N_1731);
and U2120 (N_2120,N_1758,N_1946);
nor U2121 (N_2121,N_1749,N_1762);
nand U2122 (N_2122,N_1850,N_1720);
and U2123 (N_2123,N_1795,N_1534);
nand U2124 (N_2124,N_1779,N_1857);
or U2125 (N_2125,N_1934,N_1570);
nor U2126 (N_2126,N_1611,N_1699);
nand U2127 (N_2127,N_1546,N_1552);
xnor U2128 (N_2128,N_1918,N_1897);
and U2129 (N_2129,N_1637,N_1768);
and U2130 (N_2130,N_1594,N_1903);
or U2131 (N_2131,N_1706,N_1703);
or U2132 (N_2132,N_1785,N_1842);
or U2133 (N_2133,N_1702,N_1961);
or U2134 (N_2134,N_1743,N_1661);
nand U2135 (N_2135,N_1674,N_1777);
and U2136 (N_2136,N_1572,N_1648);
nand U2137 (N_2137,N_1924,N_1579);
or U2138 (N_2138,N_1662,N_1524);
nor U2139 (N_2139,N_1530,N_1927);
and U2140 (N_2140,N_1900,N_1776);
nand U2141 (N_2141,N_1789,N_1940);
and U2142 (N_2142,N_1507,N_1615);
and U2143 (N_2143,N_1949,N_1886);
nor U2144 (N_2144,N_1845,N_1829);
nand U2145 (N_2145,N_1819,N_1982);
nor U2146 (N_2146,N_1602,N_1858);
or U2147 (N_2147,N_1799,N_1608);
and U2148 (N_2148,N_1625,N_1725);
or U2149 (N_2149,N_1547,N_1960);
nor U2150 (N_2150,N_1628,N_1985);
nand U2151 (N_2151,N_1673,N_1506);
and U2152 (N_2152,N_1810,N_1659);
nor U2153 (N_2153,N_1948,N_1930);
nor U2154 (N_2154,N_1870,N_1911);
or U2155 (N_2155,N_1899,N_1955);
nor U2156 (N_2156,N_1736,N_1601);
or U2157 (N_2157,N_1970,N_1622);
or U2158 (N_2158,N_1972,N_1893);
and U2159 (N_2159,N_1979,N_1824);
and U2160 (N_2160,N_1679,N_1502);
and U2161 (N_2161,N_1750,N_1849);
nor U2162 (N_2162,N_1989,N_1825);
or U2163 (N_2163,N_1640,N_1991);
nor U2164 (N_2164,N_1933,N_1558);
nor U2165 (N_2165,N_1976,N_1772);
and U2166 (N_2166,N_1792,N_1730);
or U2167 (N_2167,N_1798,N_1656);
and U2168 (N_2168,N_1589,N_1908);
and U2169 (N_2169,N_1747,N_1882);
or U2170 (N_2170,N_1823,N_1607);
and U2171 (N_2171,N_1717,N_1532);
nor U2172 (N_2172,N_1892,N_1708);
and U2173 (N_2173,N_1695,N_1686);
nor U2174 (N_2174,N_1681,N_1573);
and U2175 (N_2175,N_1513,N_1707);
nand U2176 (N_2176,N_1746,N_1582);
nor U2177 (N_2177,N_1831,N_1636);
nand U2178 (N_2178,N_1592,N_1685);
and U2179 (N_2179,N_1936,N_1704);
and U2180 (N_2180,N_1754,N_1975);
nand U2181 (N_2181,N_1855,N_1877);
nor U2182 (N_2182,N_1796,N_1692);
and U2183 (N_2183,N_1639,N_1944);
nand U2184 (N_2184,N_1591,N_1854);
or U2185 (N_2185,N_1907,N_1782);
nand U2186 (N_2186,N_1543,N_1553);
nand U2187 (N_2187,N_1808,N_1945);
nand U2188 (N_2188,N_1987,N_1689);
nor U2189 (N_2189,N_1938,N_1941);
or U2190 (N_2190,N_1953,N_1958);
nor U2191 (N_2191,N_1913,N_1771);
and U2192 (N_2192,N_1734,N_1645);
nor U2193 (N_2193,N_1690,N_1827);
and U2194 (N_2194,N_1514,N_1550);
nand U2195 (N_2195,N_1664,N_1881);
nor U2196 (N_2196,N_1964,N_1773);
nand U2197 (N_2197,N_1895,N_1555);
nor U2198 (N_2198,N_1568,N_1804);
nor U2199 (N_2199,N_1677,N_1888);
xnor U2200 (N_2200,N_1809,N_1551);
and U2201 (N_2201,N_1576,N_1863);
nor U2202 (N_2202,N_1996,N_1828);
and U2203 (N_2203,N_1522,N_1638);
nor U2204 (N_2204,N_1947,N_1871);
nor U2205 (N_2205,N_1803,N_1835);
or U2206 (N_2206,N_1729,N_1723);
nand U2207 (N_2207,N_1577,N_1806);
nor U2208 (N_2208,N_1889,N_1752);
xnor U2209 (N_2209,N_1575,N_1815);
or U2210 (N_2210,N_1688,N_1585);
and U2211 (N_2211,N_1896,N_1951);
nand U2212 (N_2212,N_1766,N_1872);
or U2213 (N_2213,N_1504,N_1721);
and U2214 (N_2214,N_1898,N_1943);
and U2215 (N_2215,N_1531,N_1969);
and U2216 (N_2216,N_1654,N_1780);
nor U2217 (N_2217,N_1967,N_1963);
nor U2218 (N_2218,N_1537,N_1816);
nor U2219 (N_2219,N_1528,N_1788);
nand U2220 (N_2220,N_1765,N_1521);
or U2221 (N_2221,N_1759,N_1852);
or U2222 (N_2222,N_1905,N_1658);
and U2223 (N_2223,N_1912,N_1583);
or U2224 (N_2224,N_1757,N_1545);
and U2225 (N_2225,N_1666,N_1716);
or U2226 (N_2226,N_1715,N_1999);
nand U2227 (N_2227,N_1595,N_1791);
xor U2228 (N_2228,N_1890,N_1993);
nor U2229 (N_2229,N_1586,N_1974);
or U2230 (N_2230,N_1811,N_1603);
or U2231 (N_2231,N_1671,N_1769);
nand U2232 (N_2232,N_1909,N_1533);
or U2233 (N_2233,N_1807,N_1921);
nand U2234 (N_2234,N_1617,N_1571);
nor U2235 (N_2235,N_1705,N_1868);
or U2236 (N_2236,N_1966,N_1891);
and U2237 (N_2237,N_1860,N_1665);
nand U2238 (N_2238,N_1694,N_1797);
or U2239 (N_2239,N_1643,N_1906);
and U2240 (N_2240,N_1915,N_1990);
and U2241 (N_2241,N_1670,N_1539);
or U2242 (N_2242,N_1981,N_1714);
nand U2243 (N_2243,N_1596,N_1740);
nor U2244 (N_2244,N_1923,N_1590);
nand U2245 (N_2245,N_1867,N_1519);
or U2246 (N_2246,N_1932,N_1609);
nand U2247 (N_2247,N_1621,N_1711);
nor U2248 (N_2248,N_1518,N_1875);
nand U2249 (N_2249,N_1760,N_1901);
nor U2250 (N_2250,N_1763,N_1794);
nor U2251 (N_2251,N_1526,N_1918);
or U2252 (N_2252,N_1895,N_1854);
nor U2253 (N_2253,N_1684,N_1949);
and U2254 (N_2254,N_1736,N_1782);
nand U2255 (N_2255,N_1886,N_1759);
or U2256 (N_2256,N_1649,N_1733);
nor U2257 (N_2257,N_1877,N_1873);
nor U2258 (N_2258,N_1755,N_1979);
nor U2259 (N_2259,N_1768,N_1990);
or U2260 (N_2260,N_1581,N_1952);
and U2261 (N_2261,N_1524,N_1534);
and U2262 (N_2262,N_1929,N_1801);
or U2263 (N_2263,N_1821,N_1859);
and U2264 (N_2264,N_1668,N_1758);
and U2265 (N_2265,N_1783,N_1707);
nor U2266 (N_2266,N_1815,N_1705);
or U2267 (N_2267,N_1547,N_1992);
or U2268 (N_2268,N_1919,N_1984);
and U2269 (N_2269,N_1529,N_1813);
nand U2270 (N_2270,N_1543,N_1994);
and U2271 (N_2271,N_1814,N_1667);
nand U2272 (N_2272,N_1746,N_1539);
nor U2273 (N_2273,N_1816,N_1708);
and U2274 (N_2274,N_1570,N_1697);
nor U2275 (N_2275,N_1592,N_1560);
nor U2276 (N_2276,N_1632,N_1778);
nor U2277 (N_2277,N_1989,N_1949);
nor U2278 (N_2278,N_1970,N_1931);
and U2279 (N_2279,N_1819,N_1791);
nand U2280 (N_2280,N_1979,N_1632);
nand U2281 (N_2281,N_1542,N_1981);
nand U2282 (N_2282,N_1756,N_1817);
and U2283 (N_2283,N_1679,N_1526);
or U2284 (N_2284,N_1728,N_1586);
nand U2285 (N_2285,N_1935,N_1543);
nor U2286 (N_2286,N_1956,N_1659);
nor U2287 (N_2287,N_1699,N_1718);
nand U2288 (N_2288,N_1738,N_1742);
nor U2289 (N_2289,N_1766,N_1598);
and U2290 (N_2290,N_1678,N_1943);
nand U2291 (N_2291,N_1586,N_1637);
nor U2292 (N_2292,N_1600,N_1791);
nor U2293 (N_2293,N_1717,N_1719);
or U2294 (N_2294,N_1614,N_1961);
and U2295 (N_2295,N_1869,N_1825);
and U2296 (N_2296,N_1638,N_1631);
nand U2297 (N_2297,N_1795,N_1505);
nor U2298 (N_2298,N_1555,N_1738);
and U2299 (N_2299,N_1897,N_1651);
nand U2300 (N_2300,N_1882,N_1660);
nor U2301 (N_2301,N_1772,N_1686);
or U2302 (N_2302,N_1712,N_1676);
or U2303 (N_2303,N_1551,N_1783);
nand U2304 (N_2304,N_1652,N_1517);
and U2305 (N_2305,N_1542,N_1963);
nand U2306 (N_2306,N_1541,N_1945);
or U2307 (N_2307,N_1939,N_1679);
nor U2308 (N_2308,N_1676,N_1579);
or U2309 (N_2309,N_1657,N_1660);
nor U2310 (N_2310,N_1573,N_1884);
and U2311 (N_2311,N_1815,N_1613);
nand U2312 (N_2312,N_1889,N_1867);
and U2313 (N_2313,N_1530,N_1520);
nor U2314 (N_2314,N_1593,N_1826);
or U2315 (N_2315,N_1531,N_1686);
nor U2316 (N_2316,N_1814,N_1815);
and U2317 (N_2317,N_1767,N_1892);
nor U2318 (N_2318,N_1516,N_1943);
or U2319 (N_2319,N_1752,N_1855);
nor U2320 (N_2320,N_1694,N_1841);
nor U2321 (N_2321,N_1678,N_1562);
nor U2322 (N_2322,N_1878,N_1518);
nand U2323 (N_2323,N_1949,N_1634);
nand U2324 (N_2324,N_1682,N_1587);
or U2325 (N_2325,N_1948,N_1709);
and U2326 (N_2326,N_1573,N_1682);
and U2327 (N_2327,N_1613,N_1708);
and U2328 (N_2328,N_1814,N_1956);
nor U2329 (N_2329,N_1686,N_1864);
and U2330 (N_2330,N_1903,N_1804);
nand U2331 (N_2331,N_1811,N_1833);
nor U2332 (N_2332,N_1883,N_1968);
nor U2333 (N_2333,N_1711,N_1669);
or U2334 (N_2334,N_1829,N_1733);
nand U2335 (N_2335,N_1689,N_1883);
or U2336 (N_2336,N_1894,N_1760);
or U2337 (N_2337,N_1569,N_1824);
nand U2338 (N_2338,N_1551,N_1592);
nor U2339 (N_2339,N_1555,N_1755);
nor U2340 (N_2340,N_1636,N_1733);
nor U2341 (N_2341,N_1506,N_1679);
and U2342 (N_2342,N_1944,N_1956);
nor U2343 (N_2343,N_1981,N_1624);
nand U2344 (N_2344,N_1557,N_1699);
and U2345 (N_2345,N_1854,N_1533);
and U2346 (N_2346,N_1783,N_1520);
and U2347 (N_2347,N_1587,N_1881);
nand U2348 (N_2348,N_1863,N_1797);
nand U2349 (N_2349,N_1956,N_1837);
and U2350 (N_2350,N_1502,N_1996);
nor U2351 (N_2351,N_1932,N_1805);
and U2352 (N_2352,N_1912,N_1974);
nor U2353 (N_2353,N_1627,N_1868);
and U2354 (N_2354,N_1523,N_1920);
or U2355 (N_2355,N_1864,N_1664);
or U2356 (N_2356,N_1580,N_1797);
or U2357 (N_2357,N_1910,N_1636);
or U2358 (N_2358,N_1638,N_1565);
nor U2359 (N_2359,N_1885,N_1584);
nand U2360 (N_2360,N_1896,N_1919);
nand U2361 (N_2361,N_1531,N_1964);
nand U2362 (N_2362,N_1912,N_1931);
and U2363 (N_2363,N_1593,N_1516);
or U2364 (N_2364,N_1697,N_1611);
and U2365 (N_2365,N_1669,N_1712);
nand U2366 (N_2366,N_1702,N_1940);
or U2367 (N_2367,N_1812,N_1765);
nor U2368 (N_2368,N_1828,N_1612);
xor U2369 (N_2369,N_1970,N_1605);
and U2370 (N_2370,N_1958,N_1540);
nand U2371 (N_2371,N_1619,N_1517);
nor U2372 (N_2372,N_1685,N_1702);
and U2373 (N_2373,N_1773,N_1714);
nor U2374 (N_2374,N_1559,N_1535);
nor U2375 (N_2375,N_1609,N_1878);
or U2376 (N_2376,N_1837,N_1500);
nand U2377 (N_2377,N_1612,N_1931);
nand U2378 (N_2378,N_1644,N_1624);
or U2379 (N_2379,N_1708,N_1711);
nor U2380 (N_2380,N_1887,N_1663);
nor U2381 (N_2381,N_1714,N_1676);
nor U2382 (N_2382,N_1632,N_1945);
or U2383 (N_2383,N_1849,N_1993);
xnor U2384 (N_2384,N_1956,N_1553);
nor U2385 (N_2385,N_1767,N_1935);
and U2386 (N_2386,N_1701,N_1864);
nand U2387 (N_2387,N_1966,N_1504);
or U2388 (N_2388,N_1823,N_1792);
and U2389 (N_2389,N_1625,N_1741);
nor U2390 (N_2390,N_1551,N_1887);
nand U2391 (N_2391,N_1944,N_1870);
and U2392 (N_2392,N_1833,N_1583);
nand U2393 (N_2393,N_1529,N_1709);
and U2394 (N_2394,N_1866,N_1606);
nand U2395 (N_2395,N_1851,N_1607);
and U2396 (N_2396,N_1737,N_1756);
and U2397 (N_2397,N_1582,N_1506);
and U2398 (N_2398,N_1691,N_1919);
or U2399 (N_2399,N_1955,N_1522);
nand U2400 (N_2400,N_1528,N_1983);
nand U2401 (N_2401,N_1834,N_1812);
and U2402 (N_2402,N_1595,N_1785);
nor U2403 (N_2403,N_1810,N_1567);
nand U2404 (N_2404,N_1607,N_1614);
nor U2405 (N_2405,N_1851,N_1519);
nand U2406 (N_2406,N_1925,N_1711);
or U2407 (N_2407,N_1852,N_1574);
nand U2408 (N_2408,N_1695,N_1598);
nand U2409 (N_2409,N_1598,N_1518);
and U2410 (N_2410,N_1582,N_1817);
nand U2411 (N_2411,N_1617,N_1504);
or U2412 (N_2412,N_1725,N_1688);
nor U2413 (N_2413,N_1855,N_1878);
or U2414 (N_2414,N_1611,N_1574);
nor U2415 (N_2415,N_1776,N_1746);
or U2416 (N_2416,N_1719,N_1622);
or U2417 (N_2417,N_1740,N_1667);
or U2418 (N_2418,N_1735,N_1506);
nand U2419 (N_2419,N_1529,N_1945);
nand U2420 (N_2420,N_1834,N_1736);
nor U2421 (N_2421,N_1680,N_1948);
and U2422 (N_2422,N_1925,N_1831);
nand U2423 (N_2423,N_1931,N_1833);
and U2424 (N_2424,N_1509,N_1668);
nand U2425 (N_2425,N_1762,N_1549);
or U2426 (N_2426,N_1809,N_1601);
and U2427 (N_2427,N_1980,N_1691);
and U2428 (N_2428,N_1642,N_1859);
or U2429 (N_2429,N_1995,N_1509);
nand U2430 (N_2430,N_1629,N_1584);
or U2431 (N_2431,N_1704,N_1543);
nor U2432 (N_2432,N_1596,N_1786);
nand U2433 (N_2433,N_1985,N_1561);
and U2434 (N_2434,N_1641,N_1850);
nand U2435 (N_2435,N_1928,N_1897);
or U2436 (N_2436,N_1705,N_1960);
nand U2437 (N_2437,N_1614,N_1503);
and U2438 (N_2438,N_1713,N_1884);
or U2439 (N_2439,N_1804,N_1746);
or U2440 (N_2440,N_1778,N_1896);
and U2441 (N_2441,N_1913,N_1604);
nand U2442 (N_2442,N_1660,N_1922);
or U2443 (N_2443,N_1832,N_1675);
nor U2444 (N_2444,N_1964,N_1863);
and U2445 (N_2445,N_1947,N_1733);
nor U2446 (N_2446,N_1849,N_1681);
or U2447 (N_2447,N_1512,N_1523);
and U2448 (N_2448,N_1827,N_1968);
nand U2449 (N_2449,N_1507,N_1875);
or U2450 (N_2450,N_1987,N_1925);
or U2451 (N_2451,N_1825,N_1719);
nand U2452 (N_2452,N_1800,N_1813);
and U2453 (N_2453,N_1842,N_1748);
and U2454 (N_2454,N_1987,N_1511);
or U2455 (N_2455,N_1705,N_1898);
xnor U2456 (N_2456,N_1606,N_1980);
or U2457 (N_2457,N_1985,N_1720);
and U2458 (N_2458,N_1865,N_1732);
or U2459 (N_2459,N_1925,N_1981);
or U2460 (N_2460,N_1721,N_1914);
nor U2461 (N_2461,N_1929,N_1841);
or U2462 (N_2462,N_1619,N_1708);
xnor U2463 (N_2463,N_1830,N_1560);
nor U2464 (N_2464,N_1803,N_1998);
nand U2465 (N_2465,N_1745,N_1736);
or U2466 (N_2466,N_1626,N_1984);
and U2467 (N_2467,N_1946,N_1859);
or U2468 (N_2468,N_1637,N_1954);
or U2469 (N_2469,N_1892,N_1689);
and U2470 (N_2470,N_1790,N_1884);
nand U2471 (N_2471,N_1573,N_1654);
or U2472 (N_2472,N_1668,N_1745);
nor U2473 (N_2473,N_1964,N_1614);
nor U2474 (N_2474,N_1930,N_1525);
and U2475 (N_2475,N_1702,N_1949);
nand U2476 (N_2476,N_1968,N_1608);
or U2477 (N_2477,N_1935,N_1663);
nor U2478 (N_2478,N_1709,N_1795);
or U2479 (N_2479,N_1755,N_1777);
nand U2480 (N_2480,N_1864,N_1643);
or U2481 (N_2481,N_1753,N_1755);
or U2482 (N_2482,N_1648,N_1830);
and U2483 (N_2483,N_1593,N_1780);
and U2484 (N_2484,N_1786,N_1856);
or U2485 (N_2485,N_1944,N_1638);
and U2486 (N_2486,N_1899,N_1641);
nand U2487 (N_2487,N_1573,N_1658);
and U2488 (N_2488,N_1521,N_1600);
nor U2489 (N_2489,N_1800,N_1972);
nand U2490 (N_2490,N_1910,N_1509);
nor U2491 (N_2491,N_1799,N_1630);
nand U2492 (N_2492,N_1885,N_1644);
nor U2493 (N_2493,N_1562,N_1970);
or U2494 (N_2494,N_1951,N_1957);
nand U2495 (N_2495,N_1595,N_1864);
or U2496 (N_2496,N_1883,N_1515);
nand U2497 (N_2497,N_1673,N_1532);
or U2498 (N_2498,N_1744,N_1972);
nor U2499 (N_2499,N_1765,N_1917);
and U2500 (N_2500,N_2098,N_2131);
nand U2501 (N_2501,N_2050,N_2234);
or U2502 (N_2502,N_2117,N_2102);
nand U2503 (N_2503,N_2378,N_2188);
or U2504 (N_2504,N_2205,N_2403);
or U2505 (N_2505,N_2232,N_2096);
or U2506 (N_2506,N_2200,N_2428);
nand U2507 (N_2507,N_2390,N_2173);
nand U2508 (N_2508,N_2481,N_2391);
nand U2509 (N_2509,N_2105,N_2058);
or U2510 (N_2510,N_2444,N_2048);
nand U2511 (N_2511,N_2268,N_2278);
or U2512 (N_2512,N_2256,N_2328);
nand U2513 (N_2513,N_2263,N_2239);
nand U2514 (N_2514,N_2492,N_2347);
or U2515 (N_2515,N_2147,N_2397);
or U2516 (N_2516,N_2228,N_2178);
nor U2517 (N_2517,N_2143,N_2130);
and U2518 (N_2518,N_2359,N_2419);
nand U2519 (N_2519,N_2482,N_2047);
nand U2520 (N_2520,N_2355,N_2377);
and U2521 (N_2521,N_2259,N_2317);
or U2522 (N_2522,N_2455,N_2211);
nand U2523 (N_2523,N_2091,N_2070);
nor U2524 (N_2524,N_2494,N_2320);
nand U2525 (N_2525,N_2134,N_2158);
or U2526 (N_2526,N_2474,N_2398);
or U2527 (N_2527,N_2285,N_2413);
nor U2528 (N_2528,N_2324,N_2407);
nand U2529 (N_2529,N_2190,N_2249);
or U2530 (N_2530,N_2323,N_2055);
nor U2531 (N_2531,N_2289,N_2282);
or U2532 (N_2532,N_2451,N_2184);
nand U2533 (N_2533,N_2141,N_2418);
nor U2534 (N_2534,N_2318,N_2425);
nor U2535 (N_2535,N_2356,N_2148);
nand U2536 (N_2536,N_2108,N_2459);
nand U2537 (N_2537,N_2156,N_2023);
and U2538 (N_2538,N_2111,N_2422);
or U2539 (N_2539,N_2260,N_2498);
nand U2540 (N_2540,N_2138,N_2110);
or U2541 (N_2541,N_2243,N_2449);
and U2542 (N_2542,N_2273,N_2463);
and U2543 (N_2543,N_2342,N_2199);
and U2544 (N_2544,N_2040,N_2496);
nand U2545 (N_2545,N_2274,N_2415);
nand U2546 (N_2546,N_2401,N_2394);
nand U2547 (N_2547,N_2475,N_2251);
nor U2548 (N_2548,N_2155,N_2170);
nor U2549 (N_2549,N_2406,N_2385);
nor U2550 (N_2550,N_2340,N_2389);
and U2551 (N_2551,N_2265,N_2189);
nor U2552 (N_2552,N_2396,N_2171);
or U2553 (N_2553,N_2333,N_2215);
nand U2554 (N_2554,N_2126,N_2045);
xnor U2555 (N_2555,N_2242,N_2379);
and U2556 (N_2556,N_2016,N_2345);
nand U2557 (N_2557,N_2341,N_2434);
or U2558 (N_2558,N_2497,N_2465);
and U2559 (N_2559,N_2247,N_2272);
or U2560 (N_2560,N_2077,N_2061);
and U2561 (N_2561,N_2002,N_2408);
nor U2562 (N_2562,N_2063,N_2420);
nand U2563 (N_2563,N_2489,N_2034);
and U2564 (N_2564,N_2095,N_2325);
nand U2565 (N_2565,N_2386,N_2322);
nor U2566 (N_2566,N_2024,N_2309);
xor U2567 (N_2567,N_2248,N_2220);
or U2568 (N_2568,N_2001,N_2270);
and U2569 (N_2569,N_2468,N_2014);
nor U2570 (N_2570,N_2209,N_2246);
or U2571 (N_2571,N_2319,N_2290);
nor U2572 (N_2572,N_2043,N_2357);
and U2573 (N_2573,N_2219,N_2182);
and U2574 (N_2574,N_2181,N_2331);
nand U2575 (N_2575,N_2009,N_2367);
and U2576 (N_2576,N_2329,N_2075);
or U2577 (N_2577,N_2227,N_2392);
nand U2578 (N_2578,N_2064,N_2140);
or U2579 (N_2579,N_2099,N_2216);
and U2580 (N_2580,N_2438,N_2166);
and U2581 (N_2581,N_2037,N_2010);
nor U2582 (N_2582,N_2471,N_2454);
or U2583 (N_2583,N_2297,N_2383);
nor U2584 (N_2584,N_2253,N_2381);
nand U2585 (N_2585,N_2443,N_2177);
and U2586 (N_2586,N_2291,N_2193);
nand U2587 (N_2587,N_2281,N_2313);
or U2588 (N_2588,N_2145,N_2476);
nand U2589 (N_2589,N_2083,N_2262);
nand U2590 (N_2590,N_2339,N_2167);
nor U2591 (N_2591,N_2092,N_2087);
and U2592 (N_2592,N_2195,N_2351);
nor U2593 (N_2593,N_2296,N_2467);
nor U2594 (N_2594,N_2312,N_2019);
and U2595 (N_2595,N_2373,N_2128);
nor U2596 (N_2596,N_2186,N_2028);
nand U2597 (N_2597,N_2052,N_2264);
or U2598 (N_2598,N_2433,N_2026);
nand U2599 (N_2599,N_2124,N_2258);
and U2600 (N_2600,N_2240,N_2306);
nor U2601 (N_2601,N_2431,N_2213);
and U2602 (N_2602,N_2121,N_2033);
or U2603 (N_2603,N_2197,N_2196);
nor U2604 (N_2604,N_2107,N_2473);
nor U2605 (N_2605,N_2301,N_2169);
and U2606 (N_2606,N_2218,N_2079);
or U2607 (N_2607,N_2088,N_2041);
or U2608 (N_2608,N_2106,N_2152);
nor U2609 (N_2609,N_2022,N_2090);
or U2610 (N_2610,N_2187,N_2020);
and U2611 (N_2611,N_2000,N_2336);
nor U2612 (N_2612,N_2343,N_2032);
nor U2613 (N_2613,N_2412,N_2206);
nor U2614 (N_2614,N_2038,N_2305);
and U2615 (N_2615,N_2267,N_2157);
and U2616 (N_2616,N_2025,N_2423);
or U2617 (N_2617,N_2376,N_2279);
nand U2618 (N_2618,N_2030,N_2424);
nand U2619 (N_2619,N_2144,N_2299);
nand U2620 (N_2620,N_2487,N_2409);
and U2621 (N_2621,N_2066,N_2185);
or U2622 (N_2622,N_2115,N_2006);
and U2623 (N_2623,N_2484,N_2294);
or U2624 (N_2624,N_2230,N_2007);
nor U2625 (N_2625,N_2175,N_2238);
and U2626 (N_2626,N_2337,N_2136);
or U2627 (N_2627,N_2172,N_2348);
or U2628 (N_2628,N_2370,N_2316);
or U2629 (N_2629,N_2085,N_2114);
or U2630 (N_2630,N_2217,N_2269);
or U2631 (N_2631,N_2466,N_2133);
nor U2632 (N_2632,N_2039,N_2310);
nand U2633 (N_2633,N_2462,N_2123);
or U2634 (N_2634,N_2335,N_2160);
nand U2635 (N_2635,N_2212,N_2224);
nor U2636 (N_2636,N_2076,N_2372);
nand U2637 (N_2637,N_2477,N_2071);
nor U2638 (N_2638,N_2067,N_2132);
and U2639 (N_2639,N_2308,N_2352);
nor U2640 (N_2640,N_2469,N_2456);
or U2641 (N_2641,N_2125,N_2499);
or U2642 (N_2642,N_2003,N_2452);
nand U2643 (N_2643,N_2118,N_2146);
nand U2644 (N_2644,N_2364,N_2480);
nand U2645 (N_2645,N_2153,N_2060);
and U2646 (N_2646,N_2369,N_2168);
or U2647 (N_2647,N_2446,N_2395);
nor U2648 (N_2648,N_2151,N_2084);
and U2649 (N_2649,N_2194,N_2012);
nand U2650 (N_2650,N_2065,N_2271);
nor U2651 (N_2651,N_2387,N_2008);
or U2652 (N_2652,N_2180,N_2137);
or U2653 (N_2653,N_2074,N_2056);
nor U2654 (N_2654,N_2458,N_2283);
nor U2655 (N_2655,N_2235,N_2027);
nand U2656 (N_2656,N_2013,N_2059);
nor U2657 (N_2657,N_2236,N_2275);
nand U2658 (N_2658,N_2049,N_2223);
or U2659 (N_2659,N_2244,N_2210);
nor U2660 (N_2660,N_2104,N_2461);
and U2661 (N_2661,N_2307,N_2101);
nand U2662 (N_2662,N_2165,N_2405);
or U2663 (N_2663,N_2414,N_2159);
nor U2664 (N_2664,N_2161,N_2371);
or U2665 (N_2665,N_2127,N_2327);
and U2666 (N_2666,N_2284,N_2326);
or U2667 (N_2667,N_2162,N_2457);
nand U2668 (N_2668,N_2198,N_2287);
and U2669 (N_2669,N_2349,N_2361);
nand U2670 (N_2670,N_2426,N_2353);
and U2671 (N_2671,N_2005,N_2250);
and U2672 (N_2672,N_2081,N_2366);
nand U2673 (N_2673,N_2429,N_2417);
nor U2674 (N_2674,N_2314,N_2208);
nor U2675 (N_2675,N_2411,N_2150);
or U2676 (N_2676,N_2277,N_2241);
nand U2677 (N_2677,N_2053,N_2113);
nand U2678 (N_2678,N_2338,N_2436);
and U2679 (N_2679,N_2062,N_2464);
xor U2680 (N_2680,N_2495,N_2112);
and U2681 (N_2681,N_2254,N_2447);
nand U2682 (N_2682,N_2441,N_2202);
or U2683 (N_2683,N_2103,N_2226);
or U2684 (N_2684,N_2298,N_2015);
or U2685 (N_2685,N_2344,N_2448);
or U2686 (N_2686,N_2404,N_2094);
or U2687 (N_2687,N_2057,N_2183);
nand U2688 (N_2688,N_2334,N_2430);
nor U2689 (N_2689,N_2288,N_2164);
or U2690 (N_2690,N_2483,N_2393);
or U2691 (N_2691,N_2051,N_2191);
and U2692 (N_2692,N_2054,N_2089);
or U2693 (N_2693,N_2354,N_2490);
nor U2694 (N_2694,N_2029,N_2266);
nor U2695 (N_2695,N_2179,N_2302);
and U2696 (N_2696,N_2321,N_2068);
or U2697 (N_2697,N_2276,N_2491);
nand U2698 (N_2698,N_2031,N_2078);
nand U2699 (N_2699,N_2439,N_2255);
and U2700 (N_2700,N_2375,N_2116);
or U2701 (N_2701,N_2470,N_2214);
nor U2702 (N_2702,N_2437,N_2368);
and U2703 (N_2703,N_2416,N_2350);
nor U2704 (N_2704,N_2432,N_2072);
nor U2705 (N_2705,N_2100,N_2488);
nor U2706 (N_2706,N_2261,N_2035);
nand U2707 (N_2707,N_2201,N_2435);
and U2708 (N_2708,N_2384,N_2086);
nand U2709 (N_2709,N_2080,N_2311);
nor U2710 (N_2710,N_2069,N_2374);
nor U2711 (N_2711,N_2427,N_2093);
and U2712 (N_2712,N_2402,N_2365);
and U2713 (N_2713,N_2460,N_2479);
and U2714 (N_2714,N_2445,N_2149);
nor U2715 (N_2715,N_2221,N_2486);
nand U2716 (N_2716,N_2280,N_2011);
nor U2717 (N_2717,N_2119,N_2135);
or U2718 (N_2718,N_2303,N_2382);
nor U2719 (N_2719,N_2346,N_2493);
and U2720 (N_2720,N_2222,N_2192);
nand U2721 (N_2721,N_2004,N_2225);
and U2722 (N_2722,N_2450,N_2017);
and U2723 (N_2723,N_2400,N_2257);
or U2724 (N_2724,N_2122,N_2330);
nand U2725 (N_2725,N_2442,N_2142);
nand U2726 (N_2726,N_2315,N_2358);
or U2727 (N_2727,N_2440,N_2363);
and U2728 (N_2728,N_2293,N_2021);
and U2729 (N_2729,N_2304,N_2485);
or U2730 (N_2730,N_2472,N_2120);
nor U2731 (N_2731,N_2203,N_2097);
nor U2732 (N_2732,N_2410,N_2036);
nor U2733 (N_2733,N_2042,N_2421);
nor U2734 (N_2734,N_2129,N_2388);
nand U2735 (N_2735,N_2295,N_2286);
nand U2736 (N_2736,N_2478,N_2453);
and U2737 (N_2737,N_2229,N_2292);
or U2738 (N_2738,N_2176,N_2380);
and U2739 (N_2739,N_2174,N_2163);
or U2740 (N_2740,N_2044,N_2237);
and U2741 (N_2741,N_2073,N_2082);
nand U2742 (N_2742,N_2233,N_2332);
or U2743 (N_2743,N_2231,N_2204);
or U2744 (N_2744,N_2109,N_2362);
nand U2745 (N_2745,N_2399,N_2139);
nor U2746 (N_2746,N_2245,N_2300);
nor U2747 (N_2747,N_2018,N_2046);
nand U2748 (N_2748,N_2207,N_2252);
or U2749 (N_2749,N_2360,N_2154);
or U2750 (N_2750,N_2455,N_2119);
or U2751 (N_2751,N_2300,N_2250);
nand U2752 (N_2752,N_2060,N_2481);
and U2753 (N_2753,N_2182,N_2016);
nand U2754 (N_2754,N_2171,N_2409);
nand U2755 (N_2755,N_2101,N_2116);
or U2756 (N_2756,N_2422,N_2415);
nand U2757 (N_2757,N_2220,N_2408);
and U2758 (N_2758,N_2372,N_2077);
or U2759 (N_2759,N_2141,N_2108);
or U2760 (N_2760,N_2408,N_2494);
or U2761 (N_2761,N_2320,N_2192);
and U2762 (N_2762,N_2227,N_2151);
and U2763 (N_2763,N_2415,N_2045);
or U2764 (N_2764,N_2206,N_2124);
nor U2765 (N_2765,N_2055,N_2017);
nor U2766 (N_2766,N_2216,N_2108);
and U2767 (N_2767,N_2485,N_2410);
nor U2768 (N_2768,N_2212,N_2118);
nand U2769 (N_2769,N_2303,N_2370);
nor U2770 (N_2770,N_2460,N_2291);
or U2771 (N_2771,N_2419,N_2150);
nand U2772 (N_2772,N_2484,N_2268);
and U2773 (N_2773,N_2117,N_2139);
nand U2774 (N_2774,N_2046,N_2147);
nor U2775 (N_2775,N_2387,N_2346);
nor U2776 (N_2776,N_2181,N_2150);
and U2777 (N_2777,N_2429,N_2199);
and U2778 (N_2778,N_2066,N_2484);
nand U2779 (N_2779,N_2402,N_2161);
or U2780 (N_2780,N_2391,N_2462);
nor U2781 (N_2781,N_2450,N_2193);
or U2782 (N_2782,N_2011,N_2080);
nand U2783 (N_2783,N_2433,N_2157);
xor U2784 (N_2784,N_2148,N_2414);
and U2785 (N_2785,N_2297,N_2101);
and U2786 (N_2786,N_2032,N_2012);
and U2787 (N_2787,N_2108,N_2319);
nand U2788 (N_2788,N_2060,N_2017);
and U2789 (N_2789,N_2281,N_2377);
nor U2790 (N_2790,N_2248,N_2359);
and U2791 (N_2791,N_2467,N_2316);
nor U2792 (N_2792,N_2151,N_2349);
nand U2793 (N_2793,N_2048,N_2432);
nand U2794 (N_2794,N_2062,N_2140);
nor U2795 (N_2795,N_2276,N_2205);
nor U2796 (N_2796,N_2327,N_2226);
nand U2797 (N_2797,N_2041,N_2037);
nand U2798 (N_2798,N_2130,N_2334);
and U2799 (N_2799,N_2426,N_2181);
or U2800 (N_2800,N_2411,N_2021);
nor U2801 (N_2801,N_2047,N_2488);
nor U2802 (N_2802,N_2015,N_2212);
nand U2803 (N_2803,N_2270,N_2249);
nand U2804 (N_2804,N_2217,N_2478);
or U2805 (N_2805,N_2047,N_2379);
nand U2806 (N_2806,N_2447,N_2001);
nor U2807 (N_2807,N_2057,N_2231);
and U2808 (N_2808,N_2163,N_2320);
nand U2809 (N_2809,N_2435,N_2497);
and U2810 (N_2810,N_2218,N_2469);
nand U2811 (N_2811,N_2219,N_2327);
nand U2812 (N_2812,N_2475,N_2042);
and U2813 (N_2813,N_2156,N_2039);
or U2814 (N_2814,N_2234,N_2103);
or U2815 (N_2815,N_2496,N_2494);
nand U2816 (N_2816,N_2293,N_2009);
and U2817 (N_2817,N_2035,N_2141);
nor U2818 (N_2818,N_2257,N_2166);
nand U2819 (N_2819,N_2485,N_2258);
and U2820 (N_2820,N_2238,N_2131);
nand U2821 (N_2821,N_2027,N_2438);
and U2822 (N_2822,N_2174,N_2232);
nor U2823 (N_2823,N_2367,N_2108);
and U2824 (N_2824,N_2145,N_2047);
nor U2825 (N_2825,N_2231,N_2280);
or U2826 (N_2826,N_2109,N_2250);
and U2827 (N_2827,N_2059,N_2397);
or U2828 (N_2828,N_2485,N_2094);
and U2829 (N_2829,N_2444,N_2436);
and U2830 (N_2830,N_2366,N_2227);
and U2831 (N_2831,N_2073,N_2276);
nand U2832 (N_2832,N_2197,N_2036);
and U2833 (N_2833,N_2244,N_2169);
nor U2834 (N_2834,N_2113,N_2451);
and U2835 (N_2835,N_2123,N_2124);
nand U2836 (N_2836,N_2069,N_2100);
nor U2837 (N_2837,N_2498,N_2292);
nand U2838 (N_2838,N_2470,N_2372);
xor U2839 (N_2839,N_2117,N_2026);
or U2840 (N_2840,N_2041,N_2443);
or U2841 (N_2841,N_2370,N_2053);
or U2842 (N_2842,N_2429,N_2288);
and U2843 (N_2843,N_2031,N_2448);
and U2844 (N_2844,N_2155,N_2380);
nand U2845 (N_2845,N_2218,N_2049);
nand U2846 (N_2846,N_2343,N_2094);
nor U2847 (N_2847,N_2343,N_2496);
nor U2848 (N_2848,N_2319,N_2004);
nand U2849 (N_2849,N_2302,N_2476);
or U2850 (N_2850,N_2104,N_2452);
nand U2851 (N_2851,N_2406,N_2104);
and U2852 (N_2852,N_2068,N_2011);
and U2853 (N_2853,N_2133,N_2417);
or U2854 (N_2854,N_2438,N_2117);
and U2855 (N_2855,N_2343,N_2452);
or U2856 (N_2856,N_2206,N_2315);
and U2857 (N_2857,N_2154,N_2412);
nand U2858 (N_2858,N_2377,N_2041);
or U2859 (N_2859,N_2024,N_2174);
and U2860 (N_2860,N_2376,N_2374);
nor U2861 (N_2861,N_2360,N_2355);
nor U2862 (N_2862,N_2307,N_2477);
nand U2863 (N_2863,N_2028,N_2209);
or U2864 (N_2864,N_2173,N_2034);
nor U2865 (N_2865,N_2351,N_2146);
and U2866 (N_2866,N_2398,N_2461);
and U2867 (N_2867,N_2230,N_2154);
or U2868 (N_2868,N_2372,N_2408);
and U2869 (N_2869,N_2301,N_2499);
and U2870 (N_2870,N_2216,N_2113);
nand U2871 (N_2871,N_2398,N_2409);
nand U2872 (N_2872,N_2136,N_2452);
nor U2873 (N_2873,N_2107,N_2159);
nor U2874 (N_2874,N_2090,N_2406);
or U2875 (N_2875,N_2144,N_2325);
nand U2876 (N_2876,N_2107,N_2332);
and U2877 (N_2877,N_2195,N_2224);
nor U2878 (N_2878,N_2132,N_2487);
nand U2879 (N_2879,N_2446,N_2295);
and U2880 (N_2880,N_2025,N_2451);
or U2881 (N_2881,N_2308,N_2375);
and U2882 (N_2882,N_2240,N_2431);
nor U2883 (N_2883,N_2043,N_2250);
or U2884 (N_2884,N_2155,N_2395);
nor U2885 (N_2885,N_2196,N_2442);
and U2886 (N_2886,N_2200,N_2100);
nor U2887 (N_2887,N_2024,N_2476);
and U2888 (N_2888,N_2485,N_2434);
nand U2889 (N_2889,N_2306,N_2262);
or U2890 (N_2890,N_2469,N_2369);
or U2891 (N_2891,N_2453,N_2055);
nor U2892 (N_2892,N_2388,N_2031);
or U2893 (N_2893,N_2258,N_2287);
nor U2894 (N_2894,N_2068,N_2476);
or U2895 (N_2895,N_2051,N_2388);
nor U2896 (N_2896,N_2426,N_2445);
and U2897 (N_2897,N_2310,N_2111);
or U2898 (N_2898,N_2331,N_2366);
nor U2899 (N_2899,N_2221,N_2304);
nor U2900 (N_2900,N_2171,N_2407);
or U2901 (N_2901,N_2357,N_2151);
nor U2902 (N_2902,N_2334,N_2053);
nand U2903 (N_2903,N_2432,N_2262);
or U2904 (N_2904,N_2215,N_2498);
nor U2905 (N_2905,N_2421,N_2452);
and U2906 (N_2906,N_2431,N_2340);
nand U2907 (N_2907,N_2239,N_2343);
and U2908 (N_2908,N_2416,N_2302);
nor U2909 (N_2909,N_2401,N_2377);
and U2910 (N_2910,N_2233,N_2255);
and U2911 (N_2911,N_2322,N_2443);
nor U2912 (N_2912,N_2226,N_2479);
nor U2913 (N_2913,N_2116,N_2455);
and U2914 (N_2914,N_2165,N_2390);
or U2915 (N_2915,N_2085,N_2358);
and U2916 (N_2916,N_2292,N_2163);
and U2917 (N_2917,N_2476,N_2455);
nand U2918 (N_2918,N_2038,N_2149);
or U2919 (N_2919,N_2315,N_2258);
or U2920 (N_2920,N_2207,N_2043);
xor U2921 (N_2921,N_2482,N_2003);
and U2922 (N_2922,N_2295,N_2440);
nor U2923 (N_2923,N_2083,N_2191);
or U2924 (N_2924,N_2036,N_2134);
nor U2925 (N_2925,N_2014,N_2395);
nand U2926 (N_2926,N_2049,N_2056);
and U2927 (N_2927,N_2394,N_2132);
or U2928 (N_2928,N_2255,N_2403);
nor U2929 (N_2929,N_2013,N_2051);
and U2930 (N_2930,N_2202,N_2068);
and U2931 (N_2931,N_2375,N_2118);
nand U2932 (N_2932,N_2207,N_2137);
nand U2933 (N_2933,N_2043,N_2243);
nand U2934 (N_2934,N_2439,N_2134);
or U2935 (N_2935,N_2340,N_2376);
nor U2936 (N_2936,N_2081,N_2299);
nand U2937 (N_2937,N_2277,N_2320);
or U2938 (N_2938,N_2459,N_2389);
nor U2939 (N_2939,N_2135,N_2024);
and U2940 (N_2940,N_2336,N_2367);
nor U2941 (N_2941,N_2487,N_2178);
or U2942 (N_2942,N_2121,N_2132);
or U2943 (N_2943,N_2451,N_2264);
or U2944 (N_2944,N_2436,N_2334);
or U2945 (N_2945,N_2380,N_2036);
nor U2946 (N_2946,N_2162,N_2355);
nor U2947 (N_2947,N_2300,N_2289);
and U2948 (N_2948,N_2058,N_2145);
or U2949 (N_2949,N_2101,N_2076);
xor U2950 (N_2950,N_2493,N_2344);
nand U2951 (N_2951,N_2125,N_2237);
and U2952 (N_2952,N_2328,N_2169);
or U2953 (N_2953,N_2022,N_2193);
xnor U2954 (N_2954,N_2213,N_2080);
nand U2955 (N_2955,N_2160,N_2009);
and U2956 (N_2956,N_2475,N_2082);
nor U2957 (N_2957,N_2324,N_2181);
nand U2958 (N_2958,N_2392,N_2090);
xor U2959 (N_2959,N_2464,N_2300);
nand U2960 (N_2960,N_2165,N_2489);
nand U2961 (N_2961,N_2134,N_2087);
nand U2962 (N_2962,N_2287,N_2166);
nand U2963 (N_2963,N_2299,N_2393);
and U2964 (N_2964,N_2201,N_2238);
nor U2965 (N_2965,N_2271,N_2317);
nor U2966 (N_2966,N_2163,N_2000);
nand U2967 (N_2967,N_2306,N_2422);
nand U2968 (N_2968,N_2344,N_2342);
nor U2969 (N_2969,N_2311,N_2451);
nand U2970 (N_2970,N_2265,N_2266);
or U2971 (N_2971,N_2204,N_2005);
or U2972 (N_2972,N_2311,N_2099);
nor U2973 (N_2973,N_2118,N_2013);
and U2974 (N_2974,N_2305,N_2125);
and U2975 (N_2975,N_2429,N_2095);
nor U2976 (N_2976,N_2453,N_2036);
or U2977 (N_2977,N_2227,N_2448);
nor U2978 (N_2978,N_2266,N_2392);
and U2979 (N_2979,N_2099,N_2052);
nor U2980 (N_2980,N_2423,N_2469);
nor U2981 (N_2981,N_2283,N_2461);
or U2982 (N_2982,N_2436,N_2026);
nor U2983 (N_2983,N_2428,N_2201);
nor U2984 (N_2984,N_2165,N_2366);
or U2985 (N_2985,N_2057,N_2170);
or U2986 (N_2986,N_2243,N_2197);
or U2987 (N_2987,N_2186,N_2112);
nor U2988 (N_2988,N_2493,N_2327);
nand U2989 (N_2989,N_2213,N_2243);
and U2990 (N_2990,N_2339,N_2264);
or U2991 (N_2991,N_2197,N_2139);
nor U2992 (N_2992,N_2268,N_2028);
nand U2993 (N_2993,N_2348,N_2375);
nand U2994 (N_2994,N_2123,N_2311);
or U2995 (N_2995,N_2141,N_2383);
nand U2996 (N_2996,N_2401,N_2117);
nor U2997 (N_2997,N_2093,N_2254);
and U2998 (N_2998,N_2147,N_2032);
nor U2999 (N_2999,N_2482,N_2133);
nand UO_0 (O_0,N_2900,N_2715);
or UO_1 (O_1,N_2571,N_2887);
or UO_2 (O_2,N_2832,N_2575);
and UO_3 (O_3,N_2682,N_2968);
or UO_4 (O_4,N_2954,N_2933);
nand UO_5 (O_5,N_2927,N_2716);
nor UO_6 (O_6,N_2607,N_2854);
nor UO_7 (O_7,N_2622,N_2949);
and UO_8 (O_8,N_2969,N_2879);
and UO_9 (O_9,N_2655,N_2899);
and UO_10 (O_10,N_2602,N_2986);
and UO_11 (O_11,N_2877,N_2881);
nor UO_12 (O_12,N_2936,N_2620);
or UO_13 (O_13,N_2651,N_2611);
and UO_14 (O_14,N_2627,N_2805);
and UO_15 (O_15,N_2993,N_2835);
nor UO_16 (O_16,N_2865,N_2791);
and UO_17 (O_17,N_2649,N_2723);
or UO_18 (O_18,N_2593,N_2907);
and UO_19 (O_19,N_2758,N_2856);
or UO_20 (O_20,N_2921,N_2924);
nand UO_21 (O_21,N_2834,N_2995);
and UO_22 (O_22,N_2663,N_2944);
and UO_23 (O_23,N_2714,N_2688);
or UO_24 (O_24,N_2870,N_2871);
nor UO_25 (O_25,N_2517,N_2823);
and UO_26 (O_26,N_2772,N_2676);
nand UO_27 (O_27,N_2669,N_2516);
and UO_28 (O_28,N_2630,N_2761);
nor UO_29 (O_29,N_2822,N_2556);
and UO_30 (O_30,N_2629,N_2690);
nand UO_31 (O_31,N_2643,N_2652);
and UO_32 (O_32,N_2803,N_2868);
or UO_33 (O_33,N_2527,N_2519);
nor UO_34 (O_34,N_2759,N_2780);
or UO_35 (O_35,N_2732,N_2963);
nand UO_36 (O_36,N_2683,N_2660);
or UO_37 (O_37,N_2743,N_2635);
or UO_38 (O_38,N_2557,N_2522);
nor UO_39 (O_39,N_2808,N_2932);
and UO_40 (O_40,N_2699,N_2838);
or UO_41 (O_41,N_2955,N_2615);
and UO_42 (O_42,N_2529,N_2976);
nand UO_43 (O_43,N_2513,N_2566);
and UO_44 (O_44,N_2794,N_2554);
and UO_45 (O_45,N_2935,N_2801);
nand UO_46 (O_46,N_2540,N_2819);
nand UO_47 (O_47,N_2594,N_2746);
nor UO_48 (O_48,N_2654,N_2750);
and UO_49 (O_49,N_2563,N_2719);
or UO_50 (O_50,N_2918,N_2781);
and UO_51 (O_51,N_2608,N_2561);
and UO_52 (O_52,N_2942,N_2987);
xnor UO_53 (O_53,N_2694,N_2795);
or UO_54 (O_54,N_2667,N_2790);
nor UO_55 (O_55,N_2768,N_2988);
nor UO_56 (O_56,N_2731,N_2916);
nand UO_57 (O_57,N_2775,N_2587);
and UO_58 (O_58,N_2866,N_2526);
nor UO_59 (O_59,N_2757,N_2592);
or UO_60 (O_60,N_2770,N_2626);
nor UO_61 (O_61,N_2679,N_2510);
nor UO_62 (O_62,N_2911,N_2931);
nand UO_63 (O_63,N_2930,N_2539);
or UO_64 (O_64,N_2825,N_2502);
or UO_65 (O_65,N_2804,N_2906);
or UO_66 (O_66,N_2733,N_2984);
nand UO_67 (O_67,N_2765,N_2600);
and UO_68 (O_68,N_2953,N_2747);
and UO_69 (O_69,N_2618,N_2829);
or UO_70 (O_70,N_2598,N_2590);
nor UO_71 (O_71,N_2541,N_2863);
or UO_72 (O_72,N_2905,N_2712);
or UO_73 (O_73,N_2724,N_2555);
nor UO_74 (O_74,N_2709,N_2549);
nor UO_75 (O_75,N_2606,N_2585);
xnor UO_76 (O_76,N_2559,N_2753);
or UO_77 (O_77,N_2547,N_2928);
nand UO_78 (O_78,N_2671,N_2754);
nand UO_79 (O_79,N_2853,N_2939);
and UO_80 (O_80,N_2505,N_2730);
nor UO_81 (O_81,N_2558,N_2810);
nand UO_82 (O_82,N_2596,N_2901);
and UO_83 (O_83,N_2903,N_2703);
or UO_84 (O_84,N_2837,N_2678);
nor UO_85 (O_85,N_2811,N_2893);
or UO_86 (O_86,N_2873,N_2574);
nand UO_87 (O_87,N_2553,N_2511);
nor UO_88 (O_88,N_2970,N_2710);
nand UO_89 (O_89,N_2830,N_2704);
and UO_90 (O_90,N_2929,N_2894);
or UO_91 (O_91,N_2507,N_2612);
nand UO_92 (O_92,N_2512,N_2827);
and UO_93 (O_93,N_2779,N_2833);
nand UO_94 (O_94,N_2677,N_2670);
nand UO_95 (O_95,N_2745,N_2910);
and UO_96 (O_96,N_2764,N_2562);
nand UO_97 (O_97,N_2782,N_2914);
nor UO_98 (O_98,N_2544,N_2767);
nand UO_99 (O_99,N_2972,N_2581);
and UO_100 (O_100,N_2545,N_2521);
or UO_101 (O_101,N_2964,N_2614);
or UO_102 (O_102,N_2740,N_2628);
nand UO_103 (O_103,N_2909,N_2951);
nor UO_104 (O_104,N_2705,N_2623);
nand UO_105 (O_105,N_2657,N_2604);
nor UO_106 (O_106,N_2826,N_2736);
or UO_107 (O_107,N_2849,N_2691);
or UO_108 (O_108,N_2619,N_2824);
nand UO_109 (O_109,N_2855,N_2996);
nor UO_110 (O_110,N_2713,N_2722);
nand UO_111 (O_111,N_2839,N_2673);
and UO_112 (O_112,N_2828,N_2845);
nor UO_113 (O_113,N_2568,N_2599);
and UO_114 (O_114,N_2636,N_2800);
nor UO_115 (O_115,N_2610,N_2728);
nor UO_116 (O_116,N_2565,N_2888);
nand UO_117 (O_117,N_2852,N_2898);
nor UO_118 (O_118,N_2613,N_2597);
and UO_119 (O_119,N_2576,N_2880);
nor UO_120 (O_120,N_2978,N_2895);
nor UO_121 (O_121,N_2625,N_2889);
nand UO_122 (O_122,N_2981,N_2798);
nand UO_123 (O_123,N_2760,N_2664);
and UO_124 (O_124,N_2861,N_2892);
nor UO_125 (O_125,N_2950,N_2520);
and UO_126 (O_126,N_2872,N_2749);
or UO_127 (O_127,N_2624,N_2518);
or UO_128 (O_128,N_2737,N_2595);
nand UO_129 (O_129,N_2701,N_2786);
nor UO_130 (O_130,N_2662,N_2904);
nor UO_131 (O_131,N_2584,N_2666);
nand UO_132 (O_132,N_2774,N_2846);
or UO_133 (O_133,N_2843,N_2778);
nand UO_134 (O_134,N_2840,N_2501);
nor UO_135 (O_135,N_2958,N_2902);
nor UO_136 (O_136,N_2831,N_2857);
nor UO_137 (O_137,N_2658,N_2659);
and UO_138 (O_138,N_2616,N_2862);
nor UO_139 (O_139,N_2725,N_2640);
nor UO_140 (O_140,N_2965,N_2572);
nand UO_141 (O_141,N_2579,N_2792);
nand UO_142 (O_142,N_2789,N_2818);
nor UO_143 (O_143,N_2807,N_2860);
nor UO_144 (O_144,N_2686,N_2528);
and UO_145 (O_145,N_2708,N_2882);
and UO_146 (O_146,N_2923,N_2680);
nor UO_147 (O_147,N_2564,N_2546);
nor UO_148 (O_148,N_2684,N_2943);
nand UO_149 (O_149,N_2509,N_2656);
or UO_150 (O_150,N_2920,N_2836);
nor UO_151 (O_151,N_2925,N_2848);
nand UO_152 (O_152,N_2992,N_2739);
or UO_153 (O_153,N_2644,N_2864);
or UO_154 (O_154,N_2681,N_2582);
or UO_155 (O_155,N_2959,N_2583);
nor UO_156 (O_156,N_2858,N_2915);
and UO_157 (O_157,N_2700,N_2886);
nand UO_158 (O_158,N_2755,N_2784);
or UO_159 (O_159,N_2696,N_2821);
and UO_160 (O_160,N_2633,N_2702);
and UO_161 (O_161,N_2934,N_2941);
or UO_162 (O_162,N_2638,N_2983);
and UO_163 (O_163,N_2515,N_2639);
or UO_164 (O_164,N_2551,N_2717);
nand UO_165 (O_165,N_2601,N_2738);
and UO_166 (O_166,N_2776,N_2752);
nand UO_167 (O_167,N_2817,N_2711);
nor UO_168 (O_168,N_2744,N_2734);
xor UO_169 (O_169,N_2875,N_2591);
and UO_170 (O_170,N_2689,N_2799);
nor UO_171 (O_171,N_2844,N_2977);
nor UO_172 (O_172,N_2530,N_2506);
nor UO_173 (O_173,N_2634,N_2535);
or UO_174 (O_174,N_2637,N_2525);
nand UO_175 (O_175,N_2937,N_2569);
or UO_176 (O_176,N_2726,N_2707);
nor UO_177 (O_177,N_2979,N_2815);
xnor UO_178 (O_178,N_2756,N_2645);
and UO_179 (O_179,N_2922,N_2721);
nand UO_180 (O_180,N_2806,N_2550);
nand UO_181 (O_181,N_2531,N_2945);
nand UO_182 (O_182,N_2814,N_2588);
or UO_183 (O_183,N_2891,N_2997);
or UO_184 (O_184,N_2998,N_2956);
nor UO_185 (O_185,N_2991,N_2990);
nor UO_186 (O_186,N_2809,N_2890);
or UO_187 (O_187,N_2542,N_2741);
nor UO_188 (O_188,N_2971,N_2567);
nor UO_189 (O_189,N_2771,N_2793);
nor UO_190 (O_190,N_2999,N_2777);
or UO_191 (O_191,N_2693,N_2876);
and UO_192 (O_192,N_2533,N_2573);
and UO_193 (O_193,N_2797,N_2646);
and UO_194 (O_194,N_2742,N_2578);
nor UO_195 (O_195,N_2867,N_2503);
and UO_196 (O_196,N_2665,N_2695);
nor UO_197 (O_197,N_2570,N_2982);
or UO_198 (O_198,N_2967,N_2692);
nand UO_199 (O_199,N_2919,N_2548);
and UO_200 (O_200,N_2947,N_2698);
nor UO_201 (O_201,N_2674,N_2642);
and UO_202 (O_202,N_2994,N_2813);
nor UO_203 (O_203,N_2908,N_2632);
nor UO_204 (O_204,N_2985,N_2847);
nand UO_205 (O_205,N_2560,N_2787);
or UO_206 (O_206,N_2885,N_2966);
or UO_207 (O_207,N_2538,N_2974);
nor UO_208 (O_208,N_2523,N_2841);
and UO_209 (O_209,N_2729,N_2812);
nor UO_210 (O_210,N_2524,N_2536);
or UO_211 (O_211,N_2883,N_2647);
nand UO_212 (O_212,N_2975,N_2842);
or UO_213 (O_213,N_2816,N_2661);
and UO_214 (O_214,N_2897,N_2605);
xor UO_215 (O_215,N_2884,N_2617);
nand UO_216 (O_216,N_2957,N_2718);
or UO_217 (O_217,N_2859,N_2577);
nor UO_218 (O_218,N_2766,N_2668);
and UO_219 (O_219,N_2727,N_2514);
nor UO_220 (O_220,N_2980,N_2926);
nand UO_221 (O_221,N_2961,N_2504);
nand UO_222 (O_222,N_2783,N_2973);
nor UO_223 (O_223,N_2762,N_2672);
nand UO_224 (O_224,N_2653,N_2706);
nor UO_225 (O_225,N_2748,N_2940);
xnor UO_226 (O_226,N_2621,N_2500);
nand UO_227 (O_227,N_2802,N_2720);
nand UO_228 (O_228,N_2648,N_2552);
xnor UO_229 (O_229,N_2687,N_2869);
and UO_230 (O_230,N_2769,N_2773);
nor UO_231 (O_231,N_2960,N_2675);
nand UO_232 (O_232,N_2917,N_2962);
nor UO_233 (O_233,N_2603,N_2631);
nor UO_234 (O_234,N_2851,N_2796);
or UO_235 (O_235,N_2641,N_2735);
nor UO_236 (O_236,N_2586,N_2609);
nor UO_237 (O_237,N_2537,N_2874);
nand UO_238 (O_238,N_2788,N_2850);
and UO_239 (O_239,N_2763,N_2878);
or UO_240 (O_240,N_2508,N_2913);
nor UO_241 (O_241,N_2534,N_2896);
nor UO_242 (O_242,N_2785,N_2751);
nor UO_243 (O_243,N_2532,N_2952);
nand UO_244 (O_244,N_2948,N_2685);
nand UO_245 (O_245,N_2580,N_2946);
and UO_246 (O_246,N_2912,N_2650);
nand UO_247 (O_247,N_2589,N_2820);
nand UO_248 (O_248,N_2697,N_2938);
or UO_249 (O_249,N_2989,N_2543);
or UO_250 (O_250,N_2523,N_2766);
or UO_251 (O_251,N_2648,N_2556);
and UO_252 (O_252,N_2752,N_2771);
and UO_253 (O_253,N_2541,N_2800);
nand UO_254 (O_254,N_2590,N_2592);
xnor UO_255 (O_255,N_2564,N_2838);
nor UO_256 (O_256,N_2841,N_2814);
and UO_257 (O_257,N_2932,N_2804);
nand UO_258 (O_258,N_2983,N_2770);
or UO_259 (O_259,N_2851,N_2852);
and UO_260 (O_260,N_2537,N_2619);
nand UO_261 (O_261,N_2929,N_2986);
and UO_262 (O_262,N_2608,N_2968);
and UO_263 (O_263,N_2760,N_2819);
nand UO_264 (O_264,N_2619,N_2939);
nor UO_265 (O_265,N_2727,N_2865);
nand UO_266 (O_266,N_2885,N_2916);
nor UO_267 (O_267,N_2760,N_2519);
or UO_268 (O_268,N_2739,N_2910);
xor UO_269 (O_269,N_2577,N_2583);
and UO_270 (O_270,N_2803,N_2538);
and UO_271 (O_271,N_2845,N_2825);
nand UO_272 (O_272,N_2667,N_2602);
xor UO_273 (O_273,N_2921,N_2582);
and UO_274 (O_274,N_2898,N_2521);
nand UO_275 (O_275,N_2804,N_2852);
nor UO_276 (O_276,N_2842,N_2844);
or UO_277 (O_277,N_2954,N_2918);
or UO_278 (O_278,N_2901,N_2913);
or UO_279 (O_279,N_2962,N_2615);
nand UO_280 (O_280,N_2872,N_2728);
or UO_281 (O_281,N_2885,N_2929);
nand UO_282 (O_282,N_2784,N_2620);
nand UO_283 (O_283,N_2822,N_2765);
and UO_284 (O_284,N_2882,N_2679);
and UO_285 (O_285,N_2810,N_2513);
and UO_286 (O_286,N_2757,N_2602);
and UO_287 (O_287,N_2740,N_2680);
and UO_288 (O_288,N_2675,N_2887);
or UO_289 (O_289,N_2923,N_2990);
nand UO_290 (O_290,N_2775,N_2510);
nand UO_291 (O_291,N_2756,N_2972);
and UO_292 (O_292,N_2978,N_2711);
nor UO_293 (O_293,N_2634,N_2658);
nand UO_294 (O_294,N_2932,N_2677);
and UO_295 (O_295,N_2685,N_2738);
nand UO_296 (O_296,N_2603,N_2909);
or UO_297 (O_297,N_2557,N_2539);
nand UO_298 (O_298,N_2503,N_2724);
nor UO_299 (O_299,N_2563,N_2887);
nand UO_300 (O_300,N_2617,N_2930);
nand UO_301 (O_301,N_2506,N_2514);
nand UO_302 (O_302,N_2501,N_2678);
or UO_303 (O_303,N_2658,N_2696);
and UO_304 (O_304,N_2588,N_2512);
nor UO_305 (O_305,N_2664,N_2854);
or UO_306 (O_306,N_2913,N_2581);
or UO_307 (O_307,N_2698,N_2823);
and UO_308 (O_308,N_2692,N_2619);
nor UO_309 (O_309,N_2502,N_2924);
or UO_310 (O_310,N_2588,N_2615);
or UO_311 (O_311,N_2933,N_2561);
nand UO_312 (O_312,N_2939,N_2995);
xor UO_313 (O_313,N_2561,N_2567);
or UO_314 (O_314,N_2733,N_2567);
or UO_315 (O_315,N_2718,N_2662);
nand UO_316 (O_316,N_2631,N_2529);
or UO_317 (O_317,N_2806,N_2876);
or UO_318 (O_318,N_2950,N_2954);
nor UO_319 (O_319,N_2698,N_2728);
nand UO_320 (O_320,N_2599,N_2851);
nand UO_321 (O_321,N_2992,N_2590);
nand UO_322 (O_322,N_2553,N_2791);
and UO_323 (O_323,N_2814,N_2834);
and UO_324 (O_324,N_2503,N_2553);
nor UO_325 (O_325,N_2515,N_2923);
nand UO_326 (O_326,N_2815,N_2612);
nor UO_327 (O_327,N_2646,N_2562);
or UO_328 (O_328,N_2754,N_2524);
nand UO_329 (O_329,N_2954,N_2632);
or UO_330 (O_330,N_2810,N_2912);
nand UO_331 (O_331,N_2677,N_2526);
or UO_332 (O_332,N_2843,N_2997);
and UO_333 (O_333,N_2794,N_2884);
nand UO_334 (O_334,N_2644,N_2749);
nand UO_335 (O_335,N_2785,N_2921);
or UO_336 (O_336,N_2968,N_2847);
and UO_337 (O_337,N_2804,N_2888);
or UO_338 (O_338,N_2848,N_2542);
or UO_339 (O_339,N_2539,N_2998);
or UO_340 (O_340,N_2890,N_2783);
nand UO_341 (O_341,N_2639,N_2571);
nand UO_342 (O_342,N_2929,N_2703);
and UO_343 (O_343,N_2690,N_2876);
nand UO_344 (O_344,N_2989,N_2606);
or UO_345 (O_345,N_2661,N_2875);
and UO_346 (O_346,N_2747,N_2620);
nor UO_347 (O_347,N_2560,N_2661);
nor UO_348 (O_348,N_2670,N_2530);
and UO_349 (O_349,N_2603,N_2809);
nand UO_350 (O_350,N_2771,N_2505);
nand UO_351 (O_351,N_2892,N_2560);
nor UO_352 (O_352,N_2610,N_2520);
and UO_353 (O_353,N_2789,N_2914);
nand UO_354 (O_354,N_2528,N_2918);
and UO_355 (O_355,N_2869,N_2737);
and UO_356 (O_356,N_2839,N_2898);
nand UO_357 (O_357,N_2714,N_2695);
nand UO_358 (O_358,N_2912,N_2855);
nand UO_359 (O_359,N_2679,N_2823);
nor UO_360 (O_360,N_2864,N_2988);
or UO_361 (O_361,N_2864,N_2623);
or UO_362 (O_362,N_2914,N_2575);
nor UO_363 (O_363,N_2913,N_2796);
nor UO_364 (O_364,N_2515,N_2698);
and UO_365 (O_365,N_2863,N_2942);
nand UO_366 (O_366,N_2992,N_2697);
nor UO_367 (O_367,N_2603,N_2967);
nor UO_368 (O_368,N_2720,N_2773);
nor UO_369 (O_369,N_2949,N_2951);
and UO_370 (O_370,N_2967,N_2789);
nand UO_371 (O_371,N_2618,N_2867);
and UO_372 (O_372,N_2597,N_2932);
and UO_373 (O_373,N_2987,N_2717);
nor UO_374 (O_374,N_2654,N_2503);
nor UO_375 (O_375,N_2969,N_2917);
nand UO_376 (O_376,N_2678,N_2520);
xor UO_377 (O_377,N_2794,N_2915);
nor UO_378 (O_378,N_2613,N_2788);
and UO_379 (O_379,N_2509,N_2729);
or UO_380 (O_380,N_2771,N_2632);
nand UO_381 (O_381,N_2938,N_2742);
or UO_382 (O_382,N_2959,N_2856);
and UO_383 (O_383,N_2989,N_2662);
xor UO_384 (O_384,N_2640,N_2751);
or UO_385 (O_385,N_2925,N_2852);
and UO_386 (O_386,N_2567,N_2860);
nor UO_387 (O_387,N_2701,N_2875);
or UO_388 (O_388,N_2968,N_2928);
or UO_389 (O_389,N_2910,N_2967);
or UO_390 (O_390,N_2757,N_2737);
and UO_391 (O_391,N_2938,N_2894);
nand UO_392 (O_392,N_2897,N_2703);
nand UO_393 (O_393,N_2940,N_2636);
or UO_394 (O_394,N_2821,N_2568);
or UO_395 (O_395,N_2908,N_2739);
and UO_396 (O_396,N_2973,N_2846);
or UO_397 (O_397,N_2979,N_2517);
xnor UO_398 (O_398,N_2789,N_2740);
and UO_399 (O_399,N_2636,N_2515);
and UO_400 (O_400,N_2792,N_2620);
or UO_401 (O_401,N_2544,N_2762);
nor UO_402 (O_402,N_2826,N_2767);
and UO_403 (O_403,N_2844,N_2558);
or UO_404 (O_404,N_2932,N_2889);
or UO_405 (O_405,N_2763,N_2501);
nand UO_406 (O_406,N_2574,N_2992);
or UO_407 (O_407,N_2659,N_2913);
nor UO_408 (O_408,N_2915,N_2923);
nand UO_409 (O_409,N_2594,N_2831);
or UO_410 (O_410,N_2792,N_2768);
or UO_411 (O_411,N_2617,N_2742);
nand UO_412 (O_412,N_2914,N_2790);
or UO_413 (O_413,N_2831,N_2922);
or UO_414 (O_414,N_2870,N_2897);
or UO_415 (O_415,N_2551,N_2661);
xnor UO_416 (O_416,N_2988,N_2503);
or UO_417 (O_417,N_2799,N_2511);
and UO_418 (O_418,N_2643,N_2859);
and UO_419 (O_419,N_2784,N_2552);
nor UO_420 (O_420,N_2821,N_2640);
and UO_421 (O_421,N_2852,N_2662);
and UO_422 (O_422,N_2553,N_2715);
nand UO_423 (O_423,N_2910,N_2876);
or UO_424 (O_424,N_2859,N_2951);
nor UO_425 (O_425,N_2881,N_2824);
or UO_426 (O_426,N_2540,N_2574);
and UO_427 (O_427,N_2760,N_2940);
nand UO_428 (O_428,N_2973,N_2591);
and UO_429 (O_429,N_2998,N_2988);
nand UO_430 (O_430,N_2924,N_2856);
nor UO_431 (O_431,N_2803,N_2738);
or UO_432 (O_432,N_2582,N_2801);
or UO_433 (O_433,N_2756,N_2803);
nor UO_434 (O_434,N_2750,N_2718);
nor UO_435 (O_435,N_2754,N_2963);
nor UO_436 (O_436,N_2673,N_2555);
and UO_437 (O_437,N_2828,N_2961);
nor UO_438 (O_438,N_2978,N_2669);
and UO_439 (O_439,N_2699,N_2575);
nand UO_440 (O_440,N_2623,N_2704);
nand UO_441 (O_441,N_2943,N_2961);
nand UO_442 (O_442,N_2674,N_2703);
or UO_443 (O_443,N_2670,N_2958);
or UO_444 (O_444,N_2770,N_2551);
nor UO_445 (O_445,N_2805,N_2585);
or UO_446 (O_446,N_2930,N_2661);
nand UO_447 (O_447,N_2684,N_2979);
and UO_448 (O_448,N_2891,N_2591);
and UO_449 (O_449,N_2736,N_2783);
or UO_450 (O_450,N_2852,N_2641);
and UO_451 (O_451,N_2820,N_2887);
nand UO_452 (O_452,N_2833,N_2759);
nor UO_453 (O_453,N_2836,N_2812);
nand UO_454 (O_454,N_2641,N_2690);
nand UO_455 (O_455,N_2690,N_2786);
nand UO_456 (O_456,N_2694,N_2961);
nor UO_457 (O_457,N_2928,N_2898);
and UO_458 (O_458,N_2893,N_2623);
xor UO_459 (O_459,N_2675,N_2601);
or UO_460 (O_460,N_2906,N_2553);
nand UO_461 (O_461,N_2555,N_2513);
nand UO_462 (O_462,N_2912,N_2982);
nand UO_463 (O_463,N_2665,N_2874);
or UO_464 (O_464,N_2503,N_2969);
and UO_465 (O_465,N_2795,N_2668);
or UO_466 (O_466,N_2791,N_2742);
nand UO_467 (O_467,N_2837,N_2719);
nor UO_468 (O_468,N_2651,N_2783);
and UO_469 (O_469,N_2960,N_2626);
or UO_470 (O_470,N_2679,N_2853);
nand UO_471 (O_471,N_2669,N_2624);
nor UO_472 (O_472,N_2847,N_2825);
or UO_473 (O_473,N_2791,N_2623);
or UO_474 (O_474,N_2582,N_2637);
and UO_475 (O_475,N_2550,N_2874);
and UO_476 (O_476,N_2704,N_2592);
nor UO_477 (O_477,N_2861,N_2902);
nand UO_478 (O_478,N_2873,N_2730);
nor UO_479 (O_479,N_2865,N_2590);
or UO_480 (O_480,N_2752,N_2573);
or UO_481 (O_481,N_2786,N_2916);
nor UO_482 (O_482,N_2887,N_2985);
nand UO_483 (O_483,N_2782,N_2938);
nor UO_484 (O_484,N_2889,N_2892);
nand UO_485 (O_485,N_2737,N_2759);
and UO_486 (O_486,N_2511,N_2670);
nand UO_487 (O_487,N_2968,N_2988);
and UO_488 (O_488,N_2545,N_2919);
and UO_489 (O_489,N_2922,N_2503);
nor UO_490 (O_490,N_2912,N_2835);
and UO_491 (O_491,N_2891,N_2903);
and UO_492 (O_492,N_2893,N_2618);
or UO_493 (O_493,N_2625,N_2665);
or UO_494 (O_494,N_2501,N_2734);
nor UO_495 (O_495,N_2933,N_2844);
nor UO_496 (O_496,N_2554,N_2564);
nor UO_497 (O_497,N_2837,N_2741);
or UO_498 (O_498,N_2789,N_2718);
nand UO_499 (O_499,N_2883,N_2692);
endmodule