module basic_1000_10000_1500_20_levels_2xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_392,In_459);
nor U1 (N_1,In_268,In_573);
or U2 (N_2,In_235,In_52);
nand U3 (N_3,In_804,In_753);
or U4 (N_4,In_817,In_360);
and U5 (N_5,In_670,In_289);
and U6 (N_6,In_358,In_13);
nand U7 (N_7,In_529,In_744);
xnor U8 (N_8,In_852,In_485);
xor U9 (N_9,In_497,In_935);
nor U10 (N_10,In_836,In_291);
and U11 (N_11,In_283,In_953);
or U12 (N_12,In_583,In_287);
and U13 (N_13,In_226,In_212);
or U14 (N_14,In_930,In_613);
nand U15 (N_15,In_559,In_684);
xnor U16 (N_16,In_404,In_565);
nor U17 (N_17,In_669,In_709);
nor U18 (N_18,In_203,In_356);
nor U19 (N_19,In_822,In_255);
and U20 (N_20,In_393,In_674);
nand U21 (N_21,In_812,In_476);
and U22 (N_22,In_138,In_985);
or U23 (N_23,In_845,In_607);
nor U24 (N_24,In_734,In_856);
and U25 (N_25,In_948,In_411);
and U26 (N_26,In_696,In_929);
nor U27 (N_27,In_387,In_251);
and U28 (N_28,In_994,In_717);
nand U29 (N_29,In_75,In_584);
nor U30 (N_30,In_708,In_762);
and U31 (N_31,In_471,In_232);
and U32 (N_32,In_130,In_964);
or U33 (N_33,In_659,In_545);
nor U34 (N_34,In_945,In_707);
and U35 (N_35,In_963,In_389);
nand U36 (N_36,In_769,In_40);
nor U37 (N_37,In_265,In_344);
nand U38 (N_38,In_305,In_464);
nor U39 (N_39,In_221,In_763);
nand U40 (N_40,In_775,In_57);
nor U41 (N_41,In_423,In_540);
or U42 (N_42,In_338,In_436);
xnor U43 (N_43,In_323,In_598);
nand U44 (N_44,In_957,In_81);
nand U45 (N_45,In_714,In_51);
and U46 (N_46,In_427,In_304);
nand U47 (N_47,In_509,In_313);
and U48 (N_48,In_80,In_60);
xor U49 (N_49,In_388,In_473);
and U50 (N_50,In_122,In_862);
nor U51 (N_51,In_194,In_172);
or U52 (N_52,In_248,In_556);
nor U53 (N_53,In_240,In_376);
or U54 (N_54,In_332,In_553);
nand U55 (N_55,In_335,In_858);
or U56 (N_56,In_887,In_815);
nor U57 (N_57,In_415,In_230);
and U58 (N_58,In_46,In_403);
and U59 (N_59,In_113,In_803);
or U60 (N_60,In_550,In_72);
or U61 (N_61,In_683,In_166);
or U62 (N_62,In_294,In_6);
and U63 (N_63,In_791,In_569);
nand U64 (N_64,In_89,In_516);
nor U65 (N_65,In_183,In_266);
or U66 (N_66,In_174,In_41);
nor U67 (N_67,In_570,In_560);
nand U68 (N_68,In_342,In_44);
or U69 (N_69,In_641,In_377);
nor U70 (N_70,In_206,In_209);
or U71 (N_71,In_431,In_698);
nor U72 (N_72,In_872,In_712);
or U73 (N_73,In_292,In_827);
or U74 (N_74,In_874,In_549);
and U75 (N_75,In_768,In_347);
xnor U76 (N_76,In_502,In_594);
and U77 (N_77,In_159,In_622);
and U78 (N_78,In_618,In_894);
and U79 (N_79,In_56,In_102);
and U80 (N_80,In_54,In_794);
nand U81 (N_81,In_917,In_207);
xor U82 (N_82,In_229,In_178);
nor U83 (N_83,In_308,In_574);
nor U84 (N_84,In_451,In_654);
or U85 (N_85,In_861,In_976);
and U86 (N_86,In_329,In_345);
nor U87 (N_87,In_910,In_48);
nor U88 (N_88,In_297,In_301);
and U89 (N_89,In_114,In_515);
and U90 (N_90,In_397,In_49);
nand U91 (N_91,In_430,In_83);
and U92 (N_92,In_939,In_807);
nand U93 (N_93,In_878,In_399);
nor U94 (N_94,In_264,In_364);
xnor U95 (N_95,In_156,In_608);
or U96 (N_96,In_315,In_866);
nor U97 (N_97,In_562,In_832);
and U98 (N_98,In_468,In_907);
or U99 (N_99,In_577,In_928);
nand U100 (N_100,In_390,In_742);
nand U101 (N_101,In_489,In_153);
xor U102 (N_102,In_441,In_919);
and U103 (N_103,In_331,In_93);
or U104 (N_104,In_733,In_774);
or U105 (N_105,In_630,In_117);
nand U106 (N_106,In_579,In_681);
nand U107 (N_107,In_262,In_300);
and U108 (N_108,In_539,In_228);
nand U109 (N_109,In_310,In_846);
and U110 (N_110,In_980,In_472);
nor U111 (N_111,In_373,In_567);
nor U112 (N_112,In_968,In_299);
or U113 (N_113,In_648,In_655);
or U114 (N_114,In_317,In_326);
nor U115 (N_115,In_946,In_367);
or U116 (N_116,In_951,In_754);
or U117 (N_117,In_790,In_84);
nand U118 (N_118,In_28,In_62);
and U119 (N_119,In_278,In_564);
nand U120 (N_120,In_470,In_220);
nor U121 (N_121,In_600,In_391);
or U122 (N_122,In_844,In_327);
nand U123 (N_123,In_616,In_810);
and U124 (N_124,In_64,In_692);
nor U125 (N_125,In_841,In_958);
nor U126 (N_126,In_523,In_309);
xor U127 (N_127,In_177,In_334);
and U128 (N_128,In_371,In_546);
nand U129 (N_129,In_311,In_18);
and U130 (N_130,In_284,In_30);
and U131 (N_131,In_971,In_39);
nor U132 (N_132,In_133,In_109);
and U133 (N_133,In_168,In_580);
nor U134 (N_134,In_795,In_433);
nand U135 (N_135,In_414,In_261);
and U136 (N_136,In_179,In_250);
and U137 (N_137,In_704,In_873);
and U138 (N_138,In_947,In_913);
or U139 (N_139,In_596,In_282);
and U140 (N_140,In_79,In_325);
or U141 (N_141,In_854,In_418);
nor U142 (N_142,In_591,In_626);
nand U143 (N_143,In_285,In_426);
nand U144 (N_144,In_814,In_219);
or U145 (N_145,In_990,In_806);
and U146 (N_146,In_2,In_944);
and U147 (N_147,In_756,In_86);
and U148 (N_148,In_989,In_189);
nor U149 (N_149,In_745,In_611);
or U150 (N_150,In_69,In_429);
nand U151 (N_151,In_888,In_105);
nand U152 (N_152,In_355,In_528);
or U153 (N_153,In_760,In_526);
nor U154 (N_154,In_719,In_952);
nor U155 (N_155,In_413,In_838);
nand U156 (N_156,In_767,In_123);
or U157 (N_157,In_307,In_274);
nor U158 (N_158,In_771,In_672);
and U159 (N_159,In_91,In_800);
and U160 (N_160,In_9,In_524);
and U161 (N_161,In_269,In_370);
nand U162 (N_162,In_749,In_766);
and U163 (N_163,In_8,In_22);
xnor U164 (N_164,In_972,In_855);
nor U165 (N_165,In_909,In_925);
nand U166 (N_166,In_503,In_384);
or U167 (N_167,In_0,In_78);
and U168 (N_168,In_34,In_184);
nand U169 (N_169,In_821,In_737);
nand U170 (N_170,In_517,In_893);
or U171 (N_171,In_296,In_330);
and U172 (N_172,In_870,In_181);
nand U173 (N_173,In_490,In_755);
and U174 (N_174,In_372,In_597);
or U175 (N_175,In_632,In_288);
and U176 (N_176,In_341,In_617);
and U177 (N_177,In_563,In_465);
or U178 (N_178,In_537,In_736);
xor U179 (N_179,In_357,In_970);
and U180 (N_180,In_339,In_969);
and U181 (N_181,In_934,In_190);
and U182 (N_182,In_351,In_780);
nand U183 (N_183,In_170,In_25);
or U184 (N_184,In_215,In_131);
and U185 (N_185,In_223,In_992);
nor U186 (N_186,In_53,In_561);
or U187 (N_187,In_381,In_757);
and U188 (N_188,In_35,In_880);
and U189 (N_189,In_112,In_881);
nand U190 (N_190,In_536,In_162);
nor U191 (N_191,In_513,In_995);
or U192 (N_192,In_378,In_735);
nor U193 (N_193,In_442,In_157);
nor U194 (N_194,In_628,In_204);
nand U195 (N_195,In_127,In_374);
nor U196 (N_196,In_555,In_967);
or U197 (N_197,In_965,In_635);
nand U198 (N_198,In_314,In_143);
or U199 (N_199,In_306,In_743);
nand U200 (N_200,In_31,In_77);
nor U201 (N_201,In_759,In_336);
nor U202 (N_202,In_3,In_900);
nor U203 (N_203,In_276,In_789);
and U204 (N_204,In_514,In_100);
and U205 (N_205,In_446,In_605);
and U206 (N_206,In_407,In_802);
and U207 (N_207,In_652,In_751);
or U208 (N_208,In_346,In_581);
or U209 (N_209,In_676,In_544);
nand U210 (N_210,In_463,In_152);
and U211 (N_211,In_303,In_784);
or U212 (N_212,In_864,In_90);
and U213 (N_213,In_740,In_587);
and U214 (N_214,In_542,In_481);
or U215 (N_215,In_424,In_987);
or U216 (N_216,In_918,In_891);
and U217 (N_217,In_222,In_482);
nand U218 (N_218,In_343,In_531);
nand U219 (N_219,In_128,In_601);
nand U220 (N_220,In_125,In_216);
nand U221 (N_221,In_61,In_4);
xor U222 (N_222,In_825,In_911);
or U223 (N_223,In_716,In_405);
nand U224 (N_224,In_631,In_396);
nor U225 (N_225,In_729,In_408);
nand U226 (N_226,In_551,In_36);
or U227 (N_227,In_460,In_615);
and U228 (N_228,In_614,In_350);
or U229 (N_229,In_328,In_7);
and U230 (N_230,In_857,In_12);
or U231 (N_231,In_779,In_21);
or U232 (N_232,In_653,In_43);
nand U233 (N_233,In_422,In_663);
or U234 (N_234,In_538,In_499);
nor U235 (N_235,In_772,In_643);
and U236 (N_236,In_55,In_828);
nor U237 (N_237,In_649,In_849);
nand U238 (N_238,In_210,In_275);
nand U239 (N_239,In_318,In_662);
xnor U240 (N_240,In_993,In_548);
or U241 (N_241,In_205,In_139);
and U242 (N_242,In_859,In_955);
nor U243 (N_243,In_227,In_988);
nor U244 (N_244,In_466,In_245);
nor U245 (N_245,In_478,In_715);
nor U246 (N_246,In_983,In_107);
or U247 (N_247,In_58,In_369);
or U248 (N_248,In_694,In_723);
and U249 (N_249,In_142,In_850);
and U250 (N_250,In_434,In_211);
xor U251 (N_251,In_406,In_706);
nor U252 (N_252,In_185,In_214);
or U253 (N_253,In_820,In_787);
or U254 (N_254,In_400,In_690);
and U255 (N_255,In_624,In_354);
and U256 (N_256,In_23,In_96);
nand U257 (N_257,In_14,In_146);
nor U258 (N_258,In_260,In_977);
or U259 (N_259,In_510,In_5);
or U260 (N_260,In_272,In_87);
xor U261 (N_261,In_101,In_905);
nor U262 (N_262,In_457,In_239);
nor U263 (N_263,In_758,In_45);
and U264 (N_264,In_428,In_382);
or U265 (N_265,In_785,In_650);
nor U266 (N_266,In_187,In_410);
xnor U267 (N_267,In_448,In_511);
and U268 (N_268,In_94,In_671);
and U269 (N_269,In_445,In_202);
or U270 (N_270,In_518,In_504);
nor U271 (N_271,In_664,In_960);
and U272 (N_272,In_454,In_645);
nand U273 (N_273,In_116,In_586);
nor U274 (N_274,In_621,In_991);
or U275 (N_275,In_137,In_847);
and U276 (N_276,In_799,In_498);
nor U277 (N_277,In_477,In_678);
nand U278 (N_278,In_686,In_543);
and U279 (N_279,In_950,In_180);
and U280 (N_280,In_770,In_629);
nand U281 (N_281,In_164,In_135);
xor U282 (N_282,In_134,In_363);
nand U283 (N_283,In_927,In_398);
nand U284 (N_284,In_765,In_277);
nand U285 (N_285,In_394,In_961);
xor U286 (N_286,In_158,In_612);
nand U287 (N_287,In_996,In_242);
and U288 (N_288,In_782,In_417);
nand U289 (N_289,In_981,In_924);
nand U290 (N_290,In_163,In_193);
and U291 (N_291,In_270,In_777);
and U292 (N_292,In_20,In_824);
and U293 (N_293,In_85,In_440);
nand U294 (N_294,In_682,In_456);
nor U295 (N_295,In_340,In_816);
or U296 (N_296,In_324,In_484);
nor U297 (N_297,In_699,In_585);
nor U298 (N_298,In_711,In_271);
nor U299 (N_299,In_798,In_902);
nand U300 (N_300,In_667,In_47);
and U301 (N_301,In_797,In_68);
nor U302 (N_302,In_71,In_811);
and U303 (N_303,In_450,In_444);
or U304 (N_304,In_604,In_488);
and U305 (N_305,In_160,In_17);
nand U306 (N_306,In_851,In_906);
and U307 (N_307,In_727,In_196);
and U308 (N_308,In_732,In_148);
nor U309 (N_309,In_722,In_786);
and U310 (N_310,In_973,In_241);
or U311 (N_311,In_111,In_582);
nor U312 (N_312,In_439,In_962);
nand U313 (N_313,In_38,In_954);
nand U314 (N_314,In_140,In_890);
and U315 (N_315,In_959,In_898);
nor U316 (N_316,In_530,In_932);
or U317 (N_317,In_199,In_161);
or U318 (N_318,In_984,In_480);
nor U319 (N_319,In_233,In_256);
nor U320 (N_320,In_487,In_558);
or U321 (N_321,In_644,In_750);
nand U322 (N_322,In_595,In_82);
and U323 (N_323,In_519,In_730);
nand U324 (N_324,In_169,In_108);
and U325 (N_325,In_966,In_147);
and U326 (N_326,In_512,In_703);
nor U327 (N_327,In_247,In_244);
or U328 (N_328,In_668,In_462);
nor U329 (N_329,In_124,In_88);
and U330 (N_330,In_267,In_119);
and U331 (N_331,In_349,In_295);
and U332 (N_332,In_547,In_368);
nor U333 (N_333,In_829,In_914);
nand U334 (N_334,In_486,In_923);
and U335 (N_335,In_610,In_366);
or U336 (N_336,In_126,In_637);
and U337 (N_337,In_541,In_104);
nand U338 (N_338,In_361,In_435);
nor U339 (N_339,In_720,In_141);
nand U340 (N_340,In_830,In_748);
nand U341 (N_341,In_575,In_493);
nand U342 (N_342,In_491,In_997);
nor U343 (N_343,In_195,In_273);
nor U344 (N_344,In_685,In_680);
and U345 (N_345,In_359,In_884);
and U346 (N_346,In_29,In_677);
nand U347 (N_347,In_420,In_432);
nand U348 (N_348,In_636,In_805);
xnor U349 (N_349,In_974,In_19);
nor U350 (N_350,In_693,In_32);
and U351 (N_351,In_298,In_495);
nand U352 (N_352,In_533,In_571);
and U353 (N_353,In_103,In_73);
and U354 (N_354,In_479,In_938);
or U355 (N_355,In_721,In_171);
or U356 (N_356,In_129,In_98);
nor U357 (N_357,In_876,In_728);
or U358 (N_358,In_741,In_293);
nor U359 (N_359,In_280,In_640);
nor U360 (N_360,In_634,In_165);
and U361 (N_361,In_725,In_895);
nor U362 (N_362,In_937,In_975);
and U363 (N_363,In_263,In_982);
nor U364 (N_364,In_590,In_657);
nor U365 (N_365,In_192,In_506);
or U366 (N_366,In_236,In_24);
nand U367 (N_367,In_593,In_421);
nand U368 (N_368,In_15,In_679);
nand U369 (N_369,In_362,In_176);
or U370 (N_370,In_120,In_348);
and U371 (N_371,In_182,In_74);
nor U372 (N_372,In_792,In_688);
or U373 (N_373,In_258,In_826);
nand U374 (N_374,In_201,In_606);
nor U375 (N_375,In_752,In_835);
xor U376 (N_376,In_395,In_375);
and U377 (N_377,In_818,In_449);
nor U378 (N_378,In_702,In_173);
nand U379 (N_379,In_554,In_312);
or U380 (N_380,In_149,In_380);
and U381 (N_381,In_59,In_188);
or U382 (N_382,In_281,In_522);
nand U383 (N_383,In_505,In_474);
xor U384 (N_384,In_877,In_10);
nand U385 (N_385,In_118,In_986);
or U386 (N_386,In_197,In_875);
nand U387 (N_387,In_231,In_402);
or U388 (N_388,In_458,In_921);
nor U389 (N_389,In_447,In_998);
nor U390 (N_390,In_11,In_132);
and U391 (N_391,In_319,In_724);
nand U392 (N_392,In_213,In_922);
and U393 (N_393,In_666,In_286);
and U394 (N_394,In_746,In_437);
or U395 (N_395,In_687,In_892);
or U396 (N_396,In_661,In_623);
and U397 (N_397,In_796,In_903);
nand U398 (N_398,In_191,In_700);
nor U399 (N_399,In_520,In_246);
and U400 (N_400,In_257,In_452);
or U401 (N_401,In_778,In_453);
and U402 (N_402,In_602,In_483);
nor U403 (N_403,In_882,In_869);
or U404 (N_404,In_200,In_808);
and U405 (N_405,In_842,In_92);
and U406 (N_406,In_302,In_475);
xnor U407 (N_407,In_237,In_942);
and U408 (N_408,In_110,In_889);
or U409 (N_409,In_834,In_186);
nand U410 (N_410,In_253,In_713);
nand U411 (N_411,In_238,In_175);
nand U412 (N_412,In_321,In_710);
and U413 (N_413,In_943,In_115);
and U414 (N_414,In_940,In_492);
nand U415 (N_415,In_383,In_572);
nand U416 (N_416,In_508,In_106);
nand U417 (N_417,In_224,In_689);
and U418 (N_418,In_867,In_651);
nor U419 (N_419,In_705,In_697);
xnor U420 (N_420,In_904,In_63);
and U421 (N_421,In_576,In_501);
nand U422 (N_422,In_290,In_999);
nor U423 (N_423,In_883,In_409);
nand U424 (N_424,In_809,In_978);
nand U425 (N_425,In_33,In_65);
or U426 (N_426,In_535,In_379);
nor U427 (N_427,In_879,In_568);
or U428 (N_428,In_525,In_656);
nor U429 (N_429,In_863,In_527);
nor U430 (N_430,In_781,In_701);
and U431 (N_431,In_788,In_658);
and U432 (N_432,In_899,In_783);
nor U433 (N_433,In_916,In_837);
nand U434 (N_434,In_401,In_675);
nor U435 (N_435,In_620,In_726);
or U436 (N_436,In_912,In_599);
and U437 (N_437,In_337,In_896);
xor U438 (N_438,In_813,In_908);
nor U439 (N_439,In_521,In_425);
xnor U440 (N_440,In_642,In_494);
nand U441 (N_441,In_901,In_588);
and U442 (N_442,In_121,In_933);
nand U443 (N_443,In_469,In_461);
nand U444 (N_444,In_76,In_831);
nand U445 (N_445,In_67,In_167);
and U446 (N_446,In_145,In_467);
and U447 (N_447,In_217,In_316);
nand U448 (N_448,In_865,In_915);
nand U449 (N_449,In_144,In_695);
or U450 (N_450,In_151,In_853);
or U451 (N_451,In_225,In_95);
xor U452 (N_452,In_665,In_234);
and U453 (N_453,In_731,In_333);
xor U454 (N_454,In_773,In_936);
or U455 (N_455,In_739,In_500);
and U456 (N_456,In_412,In_557);
nor U457 (N_457,In_897,In_249);
nor U458 (N_458,In_419,In_931);
nor U459 (N_459,In_496,In_871);
or U460 (N_460,In_691,In_26);
and U461 (N_461,In_150,In_603);
and U462 (N_462,In_208,In_99);
and U463 (N_463,In_926,In_252);
nor U464 (N_464,In_136,In_761);
and U465 (N_465,In_979,In_385);
nand U466 (N_466,In_353,In_552);
xnor U467 (N_467,In_1,In_619);
nor U468 (N_468,In_352,In_534);
or U469 (N_469,In_848,In_70);
or U470 (N_470,In_97,In_860);
nand U471 (N_471,In_386,In_801);
nor U472 (N_472,In_840,In_823);
or U473 (N_473,In_443,In_455);
nor U474 (N_474,In_633,In_322);
and U475 (N_475,In_638,In_279);
and U476 (N_476,In_776,In_647);
and U477 (N_477,In_566,In_155);
or U478 (N_478,In_609,In_42);
nor U479 (N_479,In_747,In_320);
or U480 (N_480,In_886,In_941);
nand U481 (N_481,In_66,In_885);
nor U482 (N_482,In_673,In_16);
nor U483 (N_483,In_254,In_218);
nand U484 (N_484,In_956,In_833);
nor U485 (N_485,In_764,In_843);
nand U486 (N_486,In_243,In_639);
xor U487 (N_487,In_949,In_589);
or U488 (N_488,In_819,In_50);
nor U489 (N_489,In_507,In_718);
nor U490 (N_490,In_868,In_793);
and U491 (N_491,In_920,In_660);
or U492 (N_492,In_154,In_532);
nand U493 (N_493,In_198,In_578);
nor U494 (N_494,In_27,In_259);
or U495 (N_495,In_646,In_625);
nand U496 (N_496,In_37,In_839);
nor U497 (N_497,In_365,In_627);
nand U498 (N_498,In_592,In_738);
or U499 (N_499,In_438,In_416);
nor U500 (N_500,N_439,N_64);
nor U501 (N_501,N_261,N_119);
nand U502 (N_502,N_272,N_363);
nand U503 (N_503,N_71,N_114);
nor U504 (N_504,N_332,N_72);
nor U505 (N_505,N_69,N_446);
nor U506 (N_506,N_312,N_136);
nor U507 (N_507,N_374,N_11);
nor U508 (N_508,N_269,N_264);
nor U509 (N_509,N_390,N_422);
nand U510 (N_510,N_495,N_150);
nor U511 (N_511,N_486,N_224);
or U512 (N_512,N_279,N_465);
or U513 (N_513,N_395,N_113);
or U514 (N_514,N_499,N_493);
xnor U515 (N_515,N_194,N_437);
nor U516 (N_516,N_449,N_87);
nand U517 (N_517,N_387,N_302);
nor U518 (N_518,N_67,N_230);
and U519 (N_519,N_303,N_248);
nor U520 (N_520,N_421,N_348);
and U521 (N_521,N_30,N_386);
and U522 (N_522,N_433,N_219);
nand U523 (N_523,N_100,N_480);
nor U524 (N_524,N_94,N_398);
and U525 (N_525,N_44,N_369);
nor U526 (N_526,N_223,N_444);
nand U527 (N_527,N_249,N_301);
nand U528 (N_528,N_297,N_56);
nor U529 (N_529,N_12,N_405);
or U530 (N_530,N_227,N_165);
and U531 (N_531,N_181,N_209);
xnor U532 (N_532,N_406,N_5);
nand U533 (N_533,N_442,N_484);
nor U534 (N_534,N_372,N_307);
nor U535 (N_535,N_61,N_323);
nand U536 (N_536,N_337,N_419);
nand U537 (N_537,N_21,N_392);
or U538 (N_538,N_3,N_490);
nand U539 (N_539,N_304,N_10);
nor U540 (N_540,N_184,N_466);
nor U541 (N_541,N_339,N_393);
xor U542 (N_542,N_360,N_259);
or U543 (N_543,N_149,N_389);
or U544 (N_544,N_212,N_48);
nor U545 (N_545,N_144,N_89);
or U546 (N_546,N_330,N_497);
nor U547 (N_547,N_345,N_265);
or U548 (N_548,N_143,N_6);
or U549 (N_549,N_161,N_475);
nor U550 (N_550,N_138,N_185);
nor U551 (N_551,N_318,N_53);
and U552 (N_552,N_322,N_229);
nand U553 (N_553,N_376,N_256);
nand U554 (N_554,N_49,N_358);
nor U555 (N_555,N_244,N_134);
or U556 (N_556,N_166,N_431);
and U557 (N_557,N_274,N_472);
nor U558 (N_558,N_139,N_57);
and U559 (N_559,N_409,N_489);
or U560 (N_560,N_84,N_154);
nor U561 (N_561,N_483,N_397);
nand U562 (N_562,N_383,N_305);
nor U563 (N_563,N_354,N_146);
and U564 (N_564,N_208,N_120);
xnor U565 (N_565,N_445,N_147);
and U566 (N_566,N_81,N_316);
and U567 (N_567,N_321,N_356);
nand U568 (N_568,N_105,N_474);
and U569 (N_569,N_122,N_325);
nand U570 (N_570,N_171,N_40);
and U571 (N_571,N_467,N_359);
nor U572 (N_572,N_461,N_291);
and U573 (N_573,N_310,N_476);
or U574 (N_574,N_388,N_257);
xnor U575 (N_575,N_167,N_39);
nor U576 (N_576,N_189,N_317);
and U577 (N_577,N_306,N_286);
and U578 (N_578,N_468,N_121);
or U579 (N_579,N_328,N_457);
and U580 (N_580,N_59,N_186);
and U581 (N_581,N_233,N_13);
or U582 (N_582,N_17,N_463);
nand U583 (N_583,N_108,N_164);
and U584 (N_584,N_454,N_29);
nor U585 (N_585,N_311,N_34);
or U586 (N_586,N_206,N_326);
and U587 (N_587,N_80,N_438);
and U588 (N_588,N_399,N_96);
nand U589 (N_589,N_443,N_62);
nor U590 (N_590,N_288,N_382);
nor U591 (N_591,N_263,N_412);
nor U592 (N_592,N_293,N_308);
nand U593 (N_593,N_349,N_357);
or U594 (N_594,N_287,N_137);
or U595 (N_595,N_205,N_459);
nand U596 (N_596,N_76,N_416);
nand U597 (N_597,N_384,N_37);
and U598 (N_598,N_267,N_469);
and U599 (N_599,N_447,N_148);
or U600 (N_600,N_116,N_155);
or U601 (N_601,N_403,N_411);
and U602 (N_602,N_225,N_236);
or U603 (N_603,N_340,N_51);
nor U604 (N_604,N_319,N_131);
nor U605 (N_605,N_343,N_109);
or U606 (N_606,N_292,N_456);
or U607 (N_607,N_430,N_156);
or U608 (N_608,N_367,N_283);
nor U609 (N_609,N_462,N_218);
nor U610 (N_610,N_141,N_213);
and U611 (N_611,N_169,N_140);
nand U612 (N_612,N_425,N_429);
nor U613 (N_613,N_498,N_246);
nand U614 (N_614,N_452,N_262);
and U615 (N_615,N_440,N_377);
nor U616 (N_616,N_414,N_385);
nand U617 (N_617,N_361,N_176);
nand U618 (N_618,N_241,N_70);
and U619 (N_619,N_333,N_232);
xnor U620 (N_620,N_38,N_35);
nand U621 (N_621,N_8,N_295);
nand U622 (N_622,N_99,N_74);
nor U623 (N_623,N_247,N_355);
and U624 (N_624,N_404,N_273);
or U625 (N_625,N_86,N_487);
nor U626 (N_626,N_401,N_88);
nor U627 (N_627,N_423,N_396);
and U628 (N_628,N_102,N_371);
nor U629 (N_629,N_210,N_496);
xor U630 (N_630,N_441,N_19);
nand U631 (N_631,N_177,N_2);
nor U632 (N_632,N_216,N_54);
nand U633 (N_633,N_128,N_296);
and U634 (N_634,N_129,N_193);
nor U635 (N_635,N_217,N_127);
or U636 (N_636,N_103,N_42);
nor U637 (N_637,N_255,N_182);
and U638 (N_638,N_254,N_36);
and U639 (N_639,N_178,N_124);
and U640 (N_640,N_491,N_91);
nor U641 (N_641,N_488,N_118);
and U642 (N_642,N_471,N_130);
nor U643 (N_643,N_207,N_329);
nand U644 (N_644,N_168,N_192);
and U645 (N_645,N_183,N_33);
nand U646 (N_646,N_180,N_107);
nand U647 (N_647,N_198,N_417);
nor U648 (N_648,N_26,N_25);
nor U649 (N_649,N_174,N_320);
or U650 (N_650,N_60,N_215);
nand U651 (N_651,N_142,N_90);
nor U652 (N_652,N_222,N_126);
nand U653 (N_653,N_9,N_407);
and U654 (N_654,N_197,N_1);
nor U655 (N_655,N_300,N_199);
nor U656 (N_656,N_350,N_27);
nor U657 (N_657,N_115,N_47);
or U658 (N_658,N_314,N_16);
and U659 (N_659,N_334,N_450);
or U660 (N_660,N_191,N_344);
or U661 (N_661,N_201,N_7);
nand U662 (N_662,N_77,N_453);
and U663 (N_663,N_46,N_458);
xor U664 (N_664,N_50,N_352);
nand U665 (N_665,N_117,N_110);
nor U666 (N_666,N_24,N_242);
nor U667 (N_667,N_170,N_370);
or U668 (N_668,N_200,N_313);
nand U669 (N_669,N_160,N_0);
nor U670 (N_670,N_111,N_335);
nand U671 (N_671,N_83,N_132);
nor U672 (N_672,N_31,N_14);
or U673 (N_673,N_494,N_270);
nor U674 (N_674,N_282,N_123);
and U675 (N_675,N_175,N_250);
nor U676 (N_676,N_55,N_20);
and U677 (N_677,N_492,N_362);
nand U678 (N_678,N_92,N_226);
and U679 (N_679,N_478,N_485);
nand U680 (N_680,N_464,N_451);
and U681 (N_681,N_4,N_93);
or U682 (N_682,N_435,N_294);
and U683 (N_683,N_101,N_432);
or U684 (N_684,N_157,N_187);
or U685 (N_685,N_290,N_342);
nor U686 (N_686,N_373,N_43);
nand U687 (N_687,N_15,N_158);
nand U688 (N_688,N_145,N_73);
nor U689 (N_689,N_221,N_234);
nand U690 (N_690,N_97,N_366);
or U691 (N_691,N_173,N_428);
nand U692 (N_692,N_298,N_473);
or U693 (N_693,N_280,N_394);
and U694 (N_694,N_275,N_82);
and U695 (N_695,N_195,N_331);
nor U696 (N_696,N_240,N_434);
or U697 (N_697,N_239,N_28);
nand U698 (N_698,N_336,N_112);
or U699 (N_699,N_231,N_79);
nand U700 (N_700,N_277,N_271);
nand U701 (N_701,N_228,N_418);
or U702 (N_702,N_188,N_202);
nand U703 (N_703,N_276,N_284);
and U704 (N_704,N_18,N_235);
nor U705 (N_705,N_163,N_85);
nor U706 (N_706,N_402,N_266);
and U707 (N_707,N_41,N_32);
and U708 (N_708,N_368,N_448);
or U709 (N_709,N_162,N_365);
and U710 (N_710,N_253,N_203);
and U711 (N_711,N_309,N_125);
nand U712 (N_712,N_341,N_415);
and U713 (N_713,N_214,N_104);
and U714 (N_714,N_391,N_460);
and U715 (N_715,N_455,N_346);
or U716 (N_716,N_375,N_299);
nand U717 (N_717,N_420,N_98);
nand U718 (N_718,N_324,N_400);
nand U719 (N_719,N_364,N_172);
and U720 (N_720,N_381,N_289);
or U721 (N_721,N_426,N_436);
or U722 (N_722,N_135,N_281);
and U723 (N_723,N_45,N_424);
nor U724 (N_724,N_327,N_22);
nand U725 (N_725,N_252,N_477);
nand U726 (N_726,N_315,N_285);
and U727 (N_727,N_238,N_220);
and U728 (N_728,N_204,N_278);
or U729 (N_729,N_153,N_23);
nor U730 (N_730,N_413,N_133);
and U731 (N_731,N_427,N_152);
and U732 (N_732,N_251,N_211);
nand U733 (N_733,N_75,N_68);
and U734 (N_734,N_353,N_260);
and U735 (N_735,N_65,N_379);
and U736 (N_736,N_63,N_151);
and U737 (N_737,N_258,N_479);
nor U738 (N_738,N_482,N_58);
and U739 (N_739,N_470,N_408);
or U740 (N_740,N_78,N_66);
and U741 (N_741,N_380,N_338);
nor U742 (N_742,N_237,N_245);
and U743 (N_743,N_243,N_410);
nand U744 (N_744,N_347,N_179);
nor U745 (N_745,N_268,N_481);
nand U746 (N_746,N_95,N_106);
or U747 (N_747,N_378,N_196);
or U748 (N_748,N_351,N_190);
nor U749 (N_749,N_52,N_159);
and U750 (N_750,N_83,N_187);
or U751 (N_751,N_46,N_329);
and U752 (N_752,N_287,N_486);
and U753 (N_753,N_163,N_69);
nor U754 (N_754,N_29,N_485);
nand U755 (N_755,N_52,N_368);
and U756 (N_756,N_129,N_215);
or U757 (N_757,N_8,N_215);
nand U758 (N_758,N_326,N_105);
or U759 (N_759,N_354,N_455);
or U760 (N_760,N_291,N_82);
nand U761 (N_761,N_120,N_431);
nand U762 (N_762,N_145,N_24);
nand U763 (N_763,N_311,N_272);
and U764 (N_764,N_400,N_86);
nand U765 (N_765,N_393,N_364);
nand U766 (N_766,N_445,N_433);
and U767 (N_767,N_169,N_81);
nand U768 (N_768,N_60,N_91);
nand U769 (N_769,N_110,N_285);
nand U770 (N_770,N_13,N_34);
or U771 (N_771,N_164,N_249);
nand U772 (N_772,N_108,N_426);
nor U773 (N_773,N_38,N_79);
or U774 (N_774,N_350,N_66);
nor U775 (N_775,N_314,N_359);
nor U776 (N_776,N_25,N_266);
or U777 (N_777,N_61,N_256);
nand U778 (N_778,N_227,N_411);
nor U779 (N_779,N_28,N_349);
xor U780 (N_780,N_9,N_491);
nand U781 (N_781,N_334,N_41);
nor U782 (N_782,N_86,N_15);
xor U783 (N_783,N_67,N_199);
nand U784 (N_784,N_402,N_88);
or U785 (N_785,N_405,N_148);
or U786 (N_786,N_371,N_366);
or U787 (N_787,N_90,N_370);
nor U788 (N_788,N_191,N_476);
nand U789 (N_789,N_345,N_90);
xnor U790 (N_790,N_58,N_279);
and U791 (N_791,N_169,N_274);
and U792 (N_792,N_112,N_420);
nand U793 (N_793,N_483,N_151);
and U794 (N_794,N_479,N_54);
and U795 (N_795,N_199,N_136);
nand U796 (N_796,N_39,N_448);
nand U797 (N_797,N_407,N_304);
and U798 (N_798,N_44,N_206);
nand U799 (N_799,N_163,N_488);
nor U800 (N_800,N_495,N_246);
nor U801 (N_801,N_147,N_461);
nand U802 (N_802,N_80,N_327);
nand U803 (N_803,N_436,N_109);
nor U804 (N_804,N_77,N_475);
nand U805 (N_805,N_10,N_483);
nand U806 (N_806,N_37,N_440);
nand U807 (N_807,N_346,N_257);
nor U808 (N_808,N_444,N_100);
nand U809 (N_809,N_459,N_293);
and U810 (N_810,N_224,N_148);
nor U811 (N_811,N_491,N_253);
or U812 (N_812,N_144,N_73);
nor U813 (N_813,N_167,N_27);
nand U814 (N_814,N_278,N_453);
nor U815 (N_815,N_225,N_151);
nor U816 (N_816,N_151,N_96);
nand U817 (N_817,N_267,N_482);
nor U818 (N_818,N_322,N_201);
and U819 (N_819,N_155,N_291);
nor U820 (N_820,N_446,N_150);
or U821 (N_821,N_26,N_179);
nand U822 (N_822,N_8,N_474);
and U823 (N_823,N_126,N_34);
nor U824 (N_824,N_130,N_457);
nor U825 (N_825,N_470,N_304);
and U826 (N_826,N_46,N_409);
xnor U827 (N_827,N_369,N_490);
nand U828 (N_828,N_191,N_49);
nor U829 (N_829,N_496,N_67);
nor U830 (N_830,N_387,N_309);
nor U831 (N_831,N_389,N_370);
nor U832 (N_832,N_164,N_180);
and U833 (N_833,N_38,N_313);
and U834 (N_834,N_67,N_167);
or U835 (N_835,N_209,N_475);
nor U836 (N_836,N_353,N_399);
nor U837 (N_837,N_107,N_206);
nor U838 (N_838,N_158,N_487);
or U839 (N_839,N_313,N_456);
nor U840 (N_840,N_398,N_7);
nand U841 (N_841,N_389,N_456);
nand U842 (N_842,N_449,N_276);
and U843 (N_843,N_267,N_485);
or U844 (N_844,N_240,N_450);
nand U845 (N_845,N_157,N_90);
and U846 (N_846,N_231,N_153);
or U847 (N_847,N_456,N_429);
or U848 (N_848,N_32,N_181);
or U849 (N_849,N_361,N_435);
or U850 (N_850,N_150,N_241);
nand U851 (N_851,N_468,N_51);
xnor U852 (N_852,N_114,N_408);
nand U853 (N_853,N_339,N_162);
nor U854 (N_854,N_481,N_167);
or U855 (N_855,N_48,N_147);
and U856 (N_856,N_229,N_320);
nor U857 (N_857,N_15,N_281);
and U858 (N_858,N_61,N_369);
nand U859 (N_859,N_176,N_168);
nand U860 (N_860,N_137,N_409);
or U861 (N_861,N_490,N_10);
nor U862 (N_862,N_141,N_387);
or U863 (N_863,N_431,N_123);
xor U864 (N_864,N_344,N_25);
nor U865 (N_865,N_141,N_337);
and U866 (N_866,N_420,N_440);
and U867 (N_867,N_24,N_385);
and U868 (N_868,N_334,N_207);
and U869 (N_869,N_309,N_369);
nor U870 (N_870,N_465,N_119);
nand U871 (N_871,N_240,N_116);
and U872 (N_872,N_493,N_487);
nand U873 (N_873,N_256,N_66);
nor U874 (N_874,N_440,N_211);
nor U875 (N_875,N_279,N_482);
nor U876 (N_876,N_460,N_224);
and U877 (N_877,N_157,N_365);
and U878 (N_878,N_357,N_260);
nand U879 (N_879,N_223,N_343);
nor U880 (N_880,N_315,N_132);
or U881 (N_881,N_204,N_82);
nand U882 (N_882,N_74,N_183);
and U883 (N_883,N_362,N_250);
or U884 (N_884,N_247,N_185);
nand U885 (N_885,N_44,N_323);
nor U886 (N_886,N_335,N_317);
nand U887 (N_887,N_34,N_160);
nand U888 (N_888,N_54,N_263);
nor U889 (N_889,N_30,N_8);
nor U890 (N_890,N_376,N_421);
and U891 (N_891,N_430,N_345);
and U892 (N_892,N_11,N_269);
and U893 (N_893,N_56,N_405);
or U894 (N_894,N_349,N_66);
nand U895 (N_895,N_271,N_20);
and U896 (N_896,N_430,N_95);
and U897 (N_897,N_21,N_220);
nor U898 (N_898,N_208,N_303);
and U899 (N_899,N_464,N_405);
nand U900 (N_900,N_475,N_41);
nor U901 (N_901,N_149,N_200);
nand U902 (N_902,N_20,N_497);
and U903 (N_903,N_395,N_180);
and U904 (N_904,N_136,N_111);
and U905 (N_905,N_287,N_458);
nand U906 (N_906,N_390,N_420);
or U907 (N_907,N_147,N_185);
or U908 (N_908,N_119,N_350);
nand U909 (N_909,N_363,N_289);
nand U910 (N_910,N_224,N_228);
xor U911 (N_911,N_210,N_69);
nor U912 (N_912,N_359,N_257);
nand U913 (N_913,N_271,N_283);
nor U914 (N_914,N_108,N_354);
nor U915 (N_915,N_71,N_435);
or U916 (N_916,N_182,N_415);
nand U917 (N_917,N_410,N_68);
nand U918 (N_918,N_73,N_88);
or U919 (N_919,N_166,N_439);
and U920 (N_920,N_443,N_193);
nor U921 (N_921,N_450,N_78);
or U922 (N_922,N_110,N_246);
or U923 (N_923,N_444,N_155);
xnor U924 (N_924,N_339,N_175);
or U925 (N_925,N_471,N_451);
nor U926 (N_926,N_413,N_378);
and U927 (N_927,N_466,N_204);
nor U928 (N_928,N_325,N_261);
nor U929 (N_929,N_29,N_187);
and U930 (N_930,N_493,N_489);
or U931 (N_931,N_239,N_295);
or U932 (N_932,N_428,N_196);
and U933 (N_933,N_112,N_127);
and U934 (N_934,N_350,N_222);
and U935 (N_935,N_301,N_254);
and U936 (N_936,N_209,N_174);
or U937 (N_937,N_441,N_331);
nor U938 (N_938,N_162,N_13);
and U939 (N_939,N_303,N_302);
or U940 (N_940,N_207,N_105);
or U941 (N_941,N_72,N_235);
nor U942 (N_942,N_170,N_418);
or U943 (N_943,N_343,N_131);
and U944 (N_944,N_310,N_404);
nand U945 (N_945,N_293,N_15);
nor U946 (N_946,N_4,N_102);
nor U947 (N_947,N_122,N_272);
or U948 (N_948,N_324,N_268);
nand U949 (N_949,N_357,N_467);
or U950 (N_950,N_241,N_312);
nand U951 (N_951,N_413,N_328);
and U952 (N_952,N_214,N_175);
nor U953 (N_953,N_268,N_492);
nor U954 (N_954,N_121,N_206);
or U955 (N_955,N_271,N_55);
and U956 (N_956,N_311,N_324);
and U957 (N_957,N_105,N_254);
or U958 (N_958,N_52,N_335);
or U959 (N_959,N_64,N_122);
or U960 (N_960,N_324,N_23);
and U961 (N_961,N_204,N_83);
nor U962 (N_962,N_252,N_66);
or U963 (N_963,N_229,N_197);
and U964 (N_964,N_442,N_407);
or U965 (N_965,N_179,N_104);
nand U966 (N_966,N_420,N_469);
nor U967 (N_967,N_121,N_140);
nand U968 (N_968,N_79,N_98);
and U969 (N_969,N_496,N_348);
nor U970 (N_970,N_61,N_297);
or U971 (N_971,N_240,N_465);
and U972 (N_972,N_249,N_170);
nor U973 (N_973,N_447,N_425);
xor U974 (N_974,N_266,N_479);
or U975 (N_975,N_95,N_189);
or U976 (N_976,N_26,N_133);
nor U977 (N_977,N_36,N_15);
nor U978 (N_978,N_379,N_307);
nand U979 (N_979,N_224,N_213);
nand U980 (N_980,N_440,N_256);
or U981 (N_981,N_379,N_316);
xnor U982 (N_982,N_288,N_166);
nand U983 (N_983,N_13,N_86);
nor U984 (N_984,N_348,N_252);
or U985 (N_985,N_349,N_284);
and U986 (N_986,N_400,N_274);
nor U987 (N_987,N_119,N_299);
and U988 (N_988,N_253,N_159);
nand U989 (N_989,N_80,N_128);
and U990 (N_990,N_345,N_407);
or U991 (N_991,N_414,N_291);
nor U992 (N_992,N_399,N_469);
and U993 (N_993,N_108,N_32);
and U994 (N_994,N_258,N_0);
or U995 (N_995,N_250,N_347);
nor U996 (N_996,N_145,N_327);
or U997 (N_997,N_123,N_447);
nor U998 (N_998,N_98,N_365);
nor U999 (N_999,N_347,N_231);
nor U1000 (N_1000,N_579,N_584);
nor U1001 (N_1001,N_553,N_538);
and U1002 (N_1002,N_652,N_655);
nor U1003 (N_1003,N_621,N_635);
nor U1004 (N_1004,N_509,N_608);
nand U1005 (N_1005,N_850,N_702);
nor U1006 (N_1006,N_982,N_744);
nor U1007 (N_1007,N_925,N_851);
or U1008 (N_1008,N_611,N_686);
xor U1009 (N_1009,N_764,N_727);
and U1010 (N_1010,N_984,N_836);
or U1011 (N_1011,N_663,N_950);
nor U1012 (N_1012,N_999,N_591);
nor U1013 (N_1013,N_594,N_846);
xor U1014 (N_1014,N_586,N_954);
nand U1015 (N_1015,N_771,N_810);
nor U1016 (N_1016,N_529,N_865);
nor U1017 (N_1017,N_902,N_794);
nor U1018 (N_1018,N_958,N_772);
or U1019 (N_1019,N_914,N_882);
nand U1020 (N_1020,N_543,N_770);
nor U1021 (N_1021,N_828,N_881);
nand U1022 (N_1022,N_540,N_880);
nor U1023 (N_1023,N_749,N_811);
nor U1024 (N_1024,N_820,N_546);
nor U1025 (N_1025,N_903,N_863);
nor U1026 (N_1026,N_994,N_573);
nor U1027 (N_1027,N_570,N_607);
nand U1028 (N_1028,N_626,N_517);
or U1029 (N_1029,N_756,N_629);
nand U1030 (N_1030,N_760,N_980);
and U1031 (N_1031,N_766,N_979);
nand U1032 (N_1032,N_932,N_685);
or U1033 (N_1033,N_666,N_716);
or U1034 (N_1034,N_730,N_550);
nand U1035 (N_1035,N_651,N_912);
nor U1036 (N_1036,N_557,N_796);
nand U1037 (N_1037,N_735,N_575);
nand U1038 (N_1038,N_693,N_637);
nor U1039 (N_1039,N_696,N_753);
nand U1040 (N_1040,N_514,N_977);
nor U1041 (N_1041,N_717,N_737);
nand U1042 (N_1042,N_878,N_734);
or U1043 (N_1043,N_551,N_567);
or U1044 (N_1044,N_838,N_501);
or U1045 (N_1045,N_833,N_713);
nand U1046 (N_1046,N_832,N_996);
nor U1047 (N_1047,N_556,N_634);
nor U1048 (N_1048,N_962,N_720);
and U1049 (N_1049,N_620,N_502);
and U1050 (N_1050,N_513,N_624);
or U1051 (N_1051,N_969,N_587);
nor U1052 (N_1052,N_719,N_671);
nand U1053 (N_1053,N_905,N_712);
and U1054 (N_1054,N_944,N_532);
or U1055 (N_1055,N_929,N_909);
and U1056 (N_1056,N_915,N_622);
nor U1057 (N_1057,N_898,N_845);
nor U1058 (N_1058,N_707,N_877);
nand U1059 (N_1059,N_806,N_653);
and U1060 (N_1060,N_780,N_741);
and U1061 (N_1061,N_554,N_662);
nand U1062 (N_1062,N_606,N_699);
nand U1063 (N_1063,N_528,N_933);
nor U1064 (N_1064,N_839,N_612);
nand U1065 (N_1065,N_987,N_904);
nor U1066 (N_1066,N_849,N_911);
nand U1067 (N_1067,N_640,N_534);
or U1068 (N_1068,N_757,N_595);
and U1069 (N_1069,N_787,N_510);
nand U1070 (N_1070,N_761,N_886);
and U1071 (N_1071,N_822,N_598);
nor U1072 (N_1072,N_544,N_873);
and U1073 (N_1073,N_507,N_889);
and U1074 (N_1074,N_648,N_660);
nor U1075 (N_1075,N_868,N_805);
nand U1076 (N_1076,N_938,N_945);
nor U1077 (N_1077,N_879,N_870);
and U1078 (N_1078,N_649,N_636);
nand U1079 (N_1079,N_542,N_650);
or U1080 (N_1080,N_960,N_688);
or U1081 (N_1081,N_853,N_799);
nand U1082 (N_1082,N_885,N_616);
xor U1083 (N_1083,N_539,N_890);
or U1084 (N_1084,N_992,N_827);
nor U1085 (N_1085,N_858,N_826);
and U1086 (N_1086,N_891,N_565);
or U1087 (N_1087,N_559,N_661);
nor U1088 (N_1088,N_767,N_816);
nor U1089 (N_1089,N_808,N_812);
and U1090 (N_1090,N_601,N_842);
or U1091 (N_1091,N_789,N_931);
nor U1092 (N_1092,N_856,N_710);
nand U1093 (N_1093,N_678,N_899);
and U1094 (N_1094,N_792,N_680);
or U1095 (N_1095,N_644,N_630);
nor U1096 (N_1096,N_817,N_500);
and U1097 (N_1097,N_829,N_701);
and U1098 (N_1098,N_689,N_562);
or U1099 (N_1099,N_961,N_888);
and U1100 (N_1100,N_941,N_927);
or U1101 (N_1101,N_729,N_536);
and U1102 (N_1102,N_940,N_871);
and U1103 (N_1103,N_779,N_837);
nand U1104 (N_1104,N_921,N_642);
nor U1105 (N_1105,N_520,N_964);
and U1106 (N_1106,N_643,N_831);
or U1107 (N_1107,N_568,N_993);
nor U1108 (N_1108,N_647,N_677);
or U1109 (N_1109,N_801,N_956);
or U1110 (N_1110,N_599,N_522);
and U1111 (N_1111,N_907,N_617);
and U1112 (N_1112,N_535,N_580);
or U1113 (N_1113,N_582,N_900);
nand U1114 (N_1114,N_596,N_955);
or U1115 (N_1115,N_659,N_623);
and U1116 (N_1116,N_813,N_997);
and U1117 (N_1117,N_600,N_602);
nand U1118 (N_1118,N_862,N_807);
nor U1119 (N_1119,N_775,N_963);
nor U1120 (N_1120,N_913,N_683);
nor U1121 (N_1121,N_852,N_848);
and U1122 (N_1122,N_555,N_706);
and U1123 (N_1123,N_672,N_967);
or U1124 (N_1124,N_973,N_521);
nor U1125 (N_1125,N_625,N_786);
or U1126 (N_1126,N_687,N_527);
and U1127 (N_1127,N_769,N_721);
nor U1128 (N_1128,N_571,N_561);
or U1129 (N_1129,N_782,N_566);
or U1130 (N_1130,N_924,N_943);
and U1131 (N_1131,N_860,N_609);
or U1132 (N_1132,N_815,N_814);
and U1133 (N_1133,N_694,N_926);
nor U1134 (N_1134,N_645,N_773);
nor U1135 (N_1135,N_558,N_819);
or U1136 (N_1136,N_919,N_667);
nand U1137 (N_1137,N_872,N_972);
or U1138 (N_1138,N_783,N_793);
or U1139 (N_1139,N_681,N_949);
nor U1140 (N_1140,N_768,N_930);
nor U1141 (N_1141,N_968,N_947);
or U1142 (N_1142,N_697,N_581);
and U1143 (N_1143,N_746,N_966);
and U1144 (N_1144,N_970,N_923);
nor U1145 (N_1145,N_859,N_525);
or U1146 (N_1146,N_658,N_603);
or U1147 (N_1147,N_818,N_533);
and U1148 (N_1148,N_804,N_883);
or U1149 (N_1149,N_765,N_763);
nor U1150 (N_1150,N_952,N_627);
and U1151 (N_1151,N_511,N_530);
nand U1152 (N_1152,N_965,N_563);
and U1153 (N_1153,N_847,N_908);
nand U1154 (N_1154,N_781,N_593);
and U1155 (N_1155,N_917,N_638);
and U1156 (N_1156,N_995,N_725);
and U1157 (N_1157,N_714,N_590);
or U1158 (N_1158,N_572,N_726);
nor U1159 (N_1159,N_942,N_646);
or U1160 (N_1160,N_974,N_703);
xor U1161 (N_1161,N_830,N_758);
nand U1162 (N_1162,N_928,N_615);
nand U1163 (N_1163,N_610,N_524);
nand U1164 (N_1164,N_824,N_560);
nand U1165 (N_1165,N_739,N_738);
and U1166 (N_1166,N_935,N_742);
and U1167 (N_1167,N_916,N_875);
nor U1168 (N_1168,N_988,N_975);
and U1169 (N_1169,N_631,N_785);
or U1170 (N_1170,N_657,N_946);
or U1171 (N_1171,N_633,N_777);
or U1172 (N_1172,N_548,N_841);
and U1173 (N_1173,N_867,N_605);
or U1174 (N_1174,N_669,N_844);
xnor U1175 (N_1175,N_989,N_731);
and U1176 (N_1176,N_894,N_800);
or U1177 (N_1177,N_887,N_733);
or U1178 (N_1178,N_704,N_691);
or U1179 (N_1179,N_695,N_545);
nand U1180 (N_1180,N_537,N_795);
nor U1181 (N_1181,N_797,N_675);
or U1182 (N_1182,N_547,N_531);
nor U1183 (N_1183,N_759,N_990);
nand U1184 (N_1184,N_656,N_654);
xnor U1185 (N_1185,N_670,N_512);
nor U1186 (N_1186,N_778,N_585);
xnor U1187 (N_1187,N_700,N_523);
nand U1188 (N_1188,N_515,N_589);
nor U1189 (N_1189,N_665,N_978);
nor U1190 (N_1190,N_869,N_985);
nor U1191 (N_1191,N_751,N_576);
and U1192 (N_1192,N_857,N_708);
nand U1193 (N_1193,N_791,N_673);
or U1194 (N_1194,N_505,N_809);
or U1195 (N_1195,N_574,N_526);
and U1196 (N_1196,N_840,N_866);
nand U1197 (N_1197,N_564,N_948);
and U1198 (N_1198,N_798,N_516);
nor U1199 (N_1199,N_549,N_821);
or U1200 (N_1200,N_748,N_506);
and U1201 (N_1201,N_628,N_577);
or U1202 (N_1202,N_711,N_698);
and U1203 (N_1203,N_774,N_802);
nand U1204 (N_1204,N_951,N_690);
or U1205 (N_1205,N_752,N_676);
xor U1206 (N_1206,N_981,N_892);
and U1207 (N_1207,N_745,N_854);
and U1208 (N_1208,N_939,N_718);
xnor U1209 (N_1209,N_583,N_834);
nor U1210 (N_1210,N_998,N_541);
and U1211 (N_1211,N_934,N_604);
nor U1212 (N_1212,N_991,N_619);
and U1213 (N_1213,N_728,N_552);
or U1214 (N_1214,N_971,N_895);
and U1215 (N_1215,N_674,N_641);
nand U1216 (N_1216,N_922,N_709);
or U1217 (N_1217,N_918,N_743);
or U1218 (N_1218,N_901,N_664);
or U1219 (N_1219,N_503,N_884);
or U1220 (N_1220,N_679,N_784);
nand U1221 (N_1221,N_790,N_618);
or U1222 (N_1222,N_723,N_724);
or U1223 (N_1223,N_588,N_861);
or U1224 (N_1224,N_614,N_803);
and U1225 (N_1225,N_632,N_613);
or U1226 (N_1226,N_747,N_639);
or U1227 (N_1227,N_976,N_508);
or U1228 (N_1228,N_519,N_855);
nor U1229 (N_1229,N_504,N_910);
nor U1230 (N_1230,N_762,N_740);
nor U1231 (N_1231,N_843,N_893);
nand U1232 (N_1232,N_668,N_736);
and U1233 (N_1233,N_682,N_825);
nand U1234 (N_1234,N_569,N_986);
nor U1235 (N_1235,N_835,N_983);
or U1236 (N_1236,N_876,N_597);
or U1237 (N_1237,N_684,N_959);
and U1238 (N_1238,N_776,N_906);
nand U1239 (N_1239,N_578,N_754);
and U1240 (N_1240,N_750,N_896);
and U1241 (N_1241,N_823,N_692);
nor U1242 (N_1242,N_957,N_755);
and U1243 (N_1243,N_788,N_705);
nand U1244 (N_1244,N_874,N_722);
and U1245 (N_1245,N_864,N_732);
or U1246 (N_1246,N_715,N_518);
nand U1247 (N_1247,N_897,N_920);
and U1248 (N_1248,N_592,N_936);
or U1249 (N_1249,N_953,N_937);
and U1250 (N_1250,N_676,N_689);
or U1251 (N_1251,N_721,N_669);
nor U1252 (N_1252,N_674,N_508);
and U1253 (N_1253,N_888,N_600);
and U1254 (N_1254,N_575,N_880);
nand U1255 (N_1255,N_814,N_856);
nand U1256 (N_1256,N_929,N_756);
or U1257 (N_1257,N_796,N_892);
nor U1258 (N_1258,N_946,N_888);
or U1259 (N_1259,N_905,N_708);
and U1260 (N_1260,N_931,N_553);
or U1261 (N_1261,N_978,N_831);
and U1262 (N_1262,N_534,N_656);
or U1263 (N_1263,N_528,N_721);
nand U1264 (N_1264,N_677,N_917);
and U1265 (N_1265,N_537,N_636);
nand U1266 (N_1266,N_504,N_579);
or U1267 (N_1267,N_536,N_597);
nor U1268 (N_1268,N_522,N_529);
nor U1269 (N_1269,N_769,N_506);
and U1270 (N_1270,N_896,N_957);
nand U1271 (N_1271,N_733,N_868);
nor U1272 (N_1272,N_575,N_669);
nand U1273 (N_1273,N_842,N_923);
or U1274 (N_1274,N_736,N_717);
and U1275 (N_1275,N_711,N_658);
nand U1276 (N_1276,N_830,N_670);
nand U1277 (N_1277,N_883,N_932);
nor U1278 (N_1278,N_945,N_514);
nand U1279 (N_1279,N_570,N_773);
and U1280 (N_1280,N_821,N_733);
nand U1281 (N_1281,N_703,N_898);
or U1282 (N_1282,N_574,N_901);
or U1283 (N_1283,N_659,N_893);
or U1284 (N_1284,N_726,N_731);
nand U1285 (N_1285,N_739,N_978);
nand U1286 (N_1286,N_947,N_604);
or U1287 (N_1287,N_822,N_627);
or U1288 (N_1288,N_822,N_523);
nand U1289 (N_1289,N_791,N_947);
or U1290 (N_1290,N_937,N_852);
xor U1291 (N_1291,N_862,N_511);
and U1292 (N_1292,N_845,N_506);
or U1293 (N_1293,N_676,N_637);
nand U1294 (N_1294,N_686,N_823);
nand U1295 (N_1295,N_567,N_970);
nor U1296 (N_1296,N_697,N_708);
or U1297 (N_1297,N_781,N_709);
and U1298 (N_1298,N_757,N_650);
and U1299 (N_1299,N_611,N_504);
or U1300 (N_1300,N_799,N_889);
nor U1301 (N_1301,N_603,N_880);
nor U1302 (N_1302,N_528,N_752);
nor U1303 (N_1303,N_762,N_746);
nand U1304 (N_1304,N_656,N_894);
nor U1305 (N_1305,N_553,N_694);
nand U1306 (N_1306,N_734,N_733);
nor U1307 (N_1307,N_560,N_935);
and U1308 (N_1308,N_662,N_865);
nand U1309 (N_1309,N_678,N_676);
nand U1310 (N_1310,N_851,N_949);
or U1311 (N_1311,N_710,N_919);
or U1312 (N_1312,N_990,N_848);
and U1313 (N_1313,N_507,N_832);
nand U1314 (N_1314,N_847,N_522);
nand U1315 (N_1315,N_598,N_612);
nand U1316 (N_1316,N_940,N_886);
and U1317 (N_1317,N_611,N_625);
and U1318 (N_1318,N_715,N_778);
or U1319 (N_1319,N_704,N_639);
nand U1320 (N_1320,N_740,N_654);
or U1321 (N_1321,N_735,N_974);
nand U1322 (N_1322,N_761,N_995);
nor U1323 (N_1323,N_984,N_532);
nor U1324 (N_1324,N_935,N_558);
or U1325 (N_1325,N_804,N_669);
nor U1326 (N_1326,N_576,N_795);
and U1327 (N_1327,N_730,N_679);
and U1328 (N_1328,N_980,N_978);
nand U1329 (N_1329,N_686,N_996);
nand U1330 (N_1330,N_655,N_791);
nor U1331 (N_1331,N_905,N_569);
nand U1332 (N_1332,N_570,N_525);
nand U1333 (N_1333,N_978,N_878);
nor U1334 (N_1334,N_801,N_971);
nand U1335 (N_1335,N_629,N_643);
nand U1336 (N_1336,N_848,N_821);
nand U1337 (N_1337,N_546,N_845);
nor U1338 (N_1338,N_690,N_696);
and U1339 (N_1339,N_542,N_920);
or U1340 (N_1340,N_829,N_681);
nand U1341 (N_1341,N_672,N_558);
or U1342 (N_1342,N_554,N_503);
or U1343 (N_1343,N_897,N_533);
or U1344 (N_1344,N_708,N_532);
nand U1345 (N_1345,N_684,N_767);
xor U1346 (N_1346,N_909,N_766);
nand U1347 (N_1347,N_808,N_720);
and U1348 (N_1348,N_744,N_600);
nor U1349 (N_1349,N_883,N_924);
nor U1350 (N_1350,N_505,N_596);
and U1351 (N_1351,N_985,N_507);
or U1352 (N_1352,N_533,N_507);
nor U1353 (N_1353,N_514,N_691);
nor U1354 (N_1354,N_949,N_890);
nand U1355 (N_1355,N_998,N_749);
and U1356 (N_1356,N_553,N_701);
nor U1357 (N_1357,N_620,N_563);
nor U1358 (N_1358,N_518,N_709);
and U1359 (N_1359,N_515,N_799);
and U1360 (N_1360,N_648,N_512);
or U1361 (N_1361,N_550,N_859);
nand U1362 (N_1362,N_625,N_822);
nor U1363 (N_1363,N_626,N_631);
nand U1364 (N_1364,N_899,N_938);
or U1365 (N_1365,N_754,N_572);
nor U1366 (N_1366,N_651,N_529);
or U1367 (N_1367,N_679,N_895);
nor U1368 (N_1368,N_811,N_882);
nand U1369 (N_1369,N_902,N_777);
or U1370 (N_1370,N_611,N_728);
nor U1371 (N_1371,N_603,N_914);
or U1372 (N_1372,N_500,N_637);
or U1373 (N_1373,N_780,N_883);
and U1374 (N_1374,N_706,N_630);
or U1375 (N_1375,N_788,N_838);
and U1376 (N_1376,N_806,N_782);
or U1377 (N_1377,N_948,N_957);
or U1378 (N_1378,N_714,N_660);
and U1379 (N_1379,N_706,N_525);
nor U1380 (N_1380,N_679,N_929);
nor U1381 (N_1381,N_777,N_603);
or U1382 (N_1382,N_692,N_779);
nor U1383 (N_1383,N_522,N_840);
nor U1384 (N_1384,N_897,N_605);
nand U1385 (N_1385,N_586,N_511);
xor U1386 (N_1386,N_776,N_540);
and U1387 (N_1387,N_801,N_947);
nand U1388 (N_1388,N_624,N_554);
nor U1389 (N_1389,N_914,N_647);
xnor U1390 (N_1390,N_543,N_821);
and U1391 (N_1391,N_674,N_950);
nor U1392 (N_1392,N_642,N_534);
and U1393 (N_1393,N_599,N_742);
or U1394 (N_1394,N_958,N_753);
nor U1395 (N_1395,N_878,N_515);
nor U1396 (N_1396,N_503,N_771);
and U1397 (N_1397,N_803,N_606);
and U1398 (N_1398,N_811,N_677);
or U1399 (N_1399,N_927,N_729);
or U1400 (N_1400,N_577,N_557);
nor U1401 (N_1401,N_812,N_682);
and U1402 (N_1402,N_940,N_789);
or U1403 (N_1403,N_722,N_841);
and U1404 (N_1404,N_743,N_714);
and U1405 (N_1405,N_612,N_852);
xor U1406 (N_1406,N_745,N_701);
or U1407 (N_1407,N_583,N_858);
nand U1408 (N_1408,N_868,N_784);
xor U1409 (N_1409,N_876,N_772);
nor U1410 (N_1410,N_911,N_780);
or U1411 (N_1411,N_690,N_816);
and U1412 (N_1412,N_552,N_508);
and U1413 (N_1413,N_656,N_558);
and U1414 (N_1414,N_547,N_997);
nand U1415 (N_1415,N_522,N_937);
or U1416 (N_1416,N_793,N_971);
or U1417 (N_1417,N_649,N_525);
or U1418 (N_1418,N_914,N_621);
nand U1419 (N_1419,N_833,N_993);
nand U1420 (N_1420,N_678,N_904);
and U1421 (N_1421,N_819,N_932);
nand U1422 (N_1422,N_613,N_639);
and U1423 (N_1423,N_805,N_640);
and U1424 (N_1424,N_622,N_599);
or U1425 (N_1425,N_965,N_741);
nand U1426 (N_1426,N_921,N_977);
and U1427 (N_1427,N_737,N_929);
nand U1428 (N_1428,N_617,N_515);
and U1429 (N_1429,N_663,N_509);
nand U1430 (N_1430,N_731,N_767);
and U1431 (N_1431,N_654,N_833);
or U1432 (N_1432,N_905,N_737);
nor U1433 (N_1433,N_697,N_746);
nor U1434 (N_1434,N_648,N_566);
or U1435 (N_1435,N_632,N_935);
or U1436 (N_1436,N_995,N_553);
nand U1437 (N_1437,N_757,N_618);
nand U1438 (N_1438,N_900,N_505);
and U1439 (N_1439,N_796,N_974);
or U1440 (N_1440,N_893,N_627);
nor U1441 (N_1441,N_714,N_984);
nor U1442 (N_1442,N_973,N_723);
xor U1443 (N_1443,N_549,N_675);
or U1444 (N_1444,N_936,N_639);
nor U1445 (N_1445,N_775,N_675);
nor U1446 (N_1446,N_638,N_822);
or U1447 (N_1447,N_568,N_706);
or U1448 (N_1448,N_858,N_827);
and U1449 (N_1449,N_986,N_761);
or U1450 (N_1450,N_592,N_727);
or U1451 (N_1451,N_550,N_757);
nor U1452 (N_1452,N_889,N_692);
nor U1453 (N_1453,N_868,N_928);
nand U1454 (N_1454,N_997,N_873);
nand U1455 (N_1455,N_621,N_848);
nand U1456 (N_1456,N_706,N_836);
or U1457 (N_1457,N_901,N_708);
and U1458 (N_1458,N_905,N_654);
or U1459 (N_1459,N_615,N_820);
nor U1460 (N_1460,N_969,N_542);
nand U1461 (N_1461,N_636,N_604);
or U1462 (N_1462,N_813,N_720);
and U1463 (N_1463,N_806,N_558);
or U1464 (N_1464,N_662,N_921);
and U1465 (N_1465,N_815,N_632);
nand U1466 (N_1466,N_800,N_954);
nand U1467 (N_1467,N_600,N_766);
or U1468 (N_1468,N_907,N_990);
nand U1469 (N_1469,N_849,N_795);
nor U1470 (N_1470,N_962,N_893);
and U1471 (N_1471,N_585,N_838);
and U1472 (N_1472,N_522,N_615);
nand U1473 (N_1473,N_944,N_965);
or U1474 (N_1474,N_766,N_676);
nor U1475 (N_1475,N_628,N_890);
nand U1476 (N_1476,N_917,N_974);
nand U1477 (N_1477,N_592,N_994);
and U1478 (N_1478,N_748,N_685);
and U1479 (N_1479,N_731,N_772);
or U1480 (N_1480,N_671,N_776);
xnor U1481 (N_1481,N_930,N_873);
and U1482 (N_1482,N_924,N_860);
xnor U1483 (N_1483,N_680,N_985);
and U1484 (N_1484,N_611,N_743);
nor U1485 (N_1485,N_594,N_644);
or U1486 (N_1486,N_635,N_663);
nand U1487 (N_1487,N_801,N_610);
xnor U1488 (N_1488,N_930,N_805);
and U1489 (N_1489,N_918,N_725);
nor U1490 (N_1490,N_803,N_865);
or U1491 (N_1491,N_844,N_801);
nand U1492 (N_1492,N_519,N_677);
or U1493 (N_1493,N_910,N_841);
nand U1494 (N_1494,N_763,N_740);
or U1495 (N_1495,N_655,N_711);
nor U1496 (N_1496,N_704,N_852);
nand U1497 (N_1497,N_680,N_502);
nor U1498 (N_1498,N_705,N_896);
nand U1499 (N_1499,N_780,N_510);
or U1500 (N_1500,N_1153,N_1381);
nor U1501 (N_1501,N_1185,N_1321);
or U1502 (N_1502,N_1215,N_1335);
nor U1503 (N_1503,N_1428,N_1259);
nand U1504 (N_1504,N_1328,N_1161);
and U1505 (N_1505,N_1006,N_1405);
nor U1506 (N_1506,N_1273,N_1093);
or U1507 (N_1507,N_1134,N_1418);
and U1508 (N_1508,N_1026,N_1411);
or U1509 (N_1509,N_1069,N_1071);
nor U1510 (N_1510,N_1446,N_1010);
or U1511 (N_1511,N_1477,N_1124);
and U1512 (N_1512,N_1081,N_1156);
and U1513 (N_1513,N_1334,N_1080);
or U1514 (N_1514,N_1284,N_1186);
nand U1515 (N_1515,N_1396,N_1345);
nand U1516 (N_1516,N_1159,N_1406);
nor U1517 (N_1517,N_1272,N_1278);
nand U1518 (N_1518,N_1052,N_1075);
nand U1519 (N_1519,N_1481,N_1299);
and U1520 (N_1520,N_1262,N_1129);
nor U1521 (N_1521,N_1043,N_1166);
or U1522 (N_1522,N_1363,N_1077);
and U1523 (N_1523,N_1230,N_1297);
nand U1524 (N_1524,N_1160,N_1233);
nor U1525 (N_1525,N_1167,N_1184);
nand U1526 (N_1526,N_1423,N_1304);
or U1527 (N_1527,N_1490,N_1264);
or U1528 (N_1528,N_1285,N_1174);
nor U1529 (N_1529,N_1229,N_1462);
and U1530 (N_1530,N_1361,N_1349);
or U1531 (N_1531,N_1275,N_1420);
nor U1532 (N_1532,N_1128,N_1137);
and U1533 (N_1533,N_1019,N_1385);
or U1534 (N_1534,N_1394,N_1136);
nand U1535 (N_1535,N_1003,N_1115);
nor U1536 (N_1536,N_1450,N_1182);
nand U1537 (N_1537,N_1101,N_1469);
and U1538 (N_1538,N_1047,N_1203);
nand U1539 (N_1539,N_1370,N_1117);
nor U1540 (N_1540,N_1293,N_1051);
nor U1541 (N_1541,N_1024,N_1076);
or U1542 (N_1542,N_1060,N_1120);
nand U1543 (N_1543,N_1465,N_1483);
nor U1544 (N_1544,N_1130,N_1053);
nand U1545 (N_1545,N_1073,N_1302);
nor U1546 (N_1546,N_1365,N_1493);
nand U1547 (N_1547,N_1257,N_1286);
xor U1548 (N_1548,N_1427,N_1360);
nand U1549 (N_1549,N_1072,N_1131);
or U1550 (N_1550,N_1187,N_1241);
and U1551 (N_1551,N_1225,N_1288);
nand U1552 (N_1552,N_1373,N_1031);
nand U1553 (N_1553,N_1213,N_1484);
nand U1554 (N_1554,N_1212,N_1029);
nand U1555 (N_1555,N_1154,N_1313);
nand U1556 (N_1556,N_1012,N_1305);
or U1557 (N_1557,N_1315,N_1416);
nor U1558 (N_1558,N_1020,N_1219);
nor U1559 (N_1559,N_1092,N_1104);
or U1560 (N_1560,N_1338,N_1352);
nor U1561 (N_1561,N_1004,N_1150);
or U1562 (N_1562,N_1414,N_1118);
or U1563 (N_1563,N_1391,N_1256);
nand U1564 (N_1564,N_1417,N_1169);
and U1565 (N_1565,N_1408,N_1290);
nand U1566 (N_1566,N_1249,N_1119);
or U1567 (N_1567,N_1366,N_1384);
nand U1568 (N_1568,N_1441,N_1298);
nand U1569 (N_1569,N_1114,N_1362);
and U1570 (N_1570,N_1274,N_1001);
nand U1571 (N_1571,N_1308,N_1250);
or U1572 (N_1572,N_1211,N_1070);
nand U1573 (N_1573,N_1466,N_1439);
nand U1574 (N_1574,N_1377,N_1289);
nor U1575 (N_1575,N_1096,N_1436);
nand U1576 (N_1576,N_1191,N_1261);
or U1577 (N_1577,N_1336,N_1422);
or U1578 (N_1578,N_1132,N_1198);
or U1579 (N_1579,N_1082,N_1235);
nand U1580 (N_1580,N_1374,N_1309);
nor U1581 (N_1581,N_1492,N_1044);
xnor U1582 (N_1582,N_1463,N_1183);
nand U1583 (N_1583,N_1399,N_1068);
or U1584 (N_1584,N_1434,N_1364);
nor U1585 (N_1585,N_1403,N_1193);
nand U1586 (N_1586,N_1295,N_1133);
nand U1587 (N_1587,N_1479,N_1437);
nand U1588 (N_1588,N_1448,N_1276);
or U1589 (N_1589,N_1277,N_1158);
nor U1590 (N_1590,N_1351,N_1379);
nor U1591 (N_1591,N_1471,N_1218);
nand U1592 (N_1592,N_1111,N_1039);
and U1593 (N_1593,N_1267,N_1472);
and U1594 (N_1594,N_1413,N_1192);
nor U1595 (N_1595,N_1487,N_1449);
and U1596 (N_1596,N_1234,N_1337);
nand U1597 (N_1597,N_1210,N_1240);
or U1598 (N_1598,N_1435,N_1320);
nand U1599 (N_1599,N_1332,N_1461);
nor U1600 (N_1600,N_1054,N_1066);
nand U1601 (N_1601,N_1110,N_1214);
nor U1602 (N_1602,N_1045,N_1036);
xor U1603 (N_1603,N_1369,N_1453);
or U1604 (N_1604,N_1410,N_1447);
nand U1605 (N_1605,N_1057,N_1400);
nand U1606 (N_1606,N_1344,N_1190);
nand U1607 (N_1607,N_1444,N_1002);
nor U1608 (N_1608,N_1202,N_1244);
nand U1609 (N_1609,N_1025,N_1094);
and U1610 (N_1610,N_1401,N_1179);
or U1611 (N_1611,N_1312,N_1063);
or U1612 (N_1612,N_1311,N_1226);
nor U1613 (N_1613,N_1474,N_1173);
or U1614 (N_1614,N_1314,N_1074);
nor U1615 (N_1615,N_1497,N_1245);
or U1616 (N_1616,N_1037,N_1280);
nand U1617 (N_1617,N_1392,N_1078);
nand U1618 (N_1618,N_1357,N_1189);
and U1619 (N_1619,N_1412,N_1170);
xor U1620 (N_1620,N_1064,N_1419);
or U1621 (N_1621,N_1407,N_1017);
nor U1622 (N_1622,N_1271,N_1103);
and U1623 (N_1623,N_1079,N_1318);
nand U1624 (N_1624,N_1227,N_1177);
or U1625 (N_1625,N_1347,N_1316);
and U1626 (N_1626,N_1329,N_1108);
xnor U1627 (N_1627,N_1388,N_1116);
nor U1628 (N_1628,N_1383,N_1459);
nor U1629 (N_1629,N_1088,N_1232);
xor U1630 (N_1630,N_1102,N_1488);
or U1631 (N_1631,N_1404,N_1018);
and U1632 (N_1632,N_1440,N_1062);
nor U1633 (N_1633,N_1270,N_1209);
nor U1634 (N_1634,N_1485,N_1112);
nor U1635 (N_1635,N_1042,N_1331);
nor U1636 (N_1636,N_1443,N_1430);
and U1637 (N_1637,N_1236,N_1098);
nand U1638 (N_1638,N_1172,N_1475);
nand U1639 (N_1639,N_1030,N_1005);
or U1640 (N_1640,N_1171,N_1491);
nand U1641 (N_1641,N_1028,N_1000);
and U1642 (N_1642,N_1220,N_1178);
nor U1643 (N_1643,N_1323,N_1216);
or U1644 (N_1644,N_1055,N_1395);
and U1645 (N_1645,N_1127,N_1105);
nand U1646 (N_1646,N_1432,N_1205);
nor U1647 (N_1647,N_1135,N_1498);
or U1648 (N_1648,N_1372,N_1109);
and U1649 (N_1649,N_1100,N_1222);
nor U1650 (N_1650,N_1126,N_1067);
nor U1651 (N_1651,N_1356,N_1035);
nand U1652 (N_1652,N_1470,N_1468);
and U1653 (N_1653,N_1367,N_1342);
nand U1654 (N_1654,N_1023,N_1138);
and U1655 (N_1655,N_1355,N_1393);
nor U1656 (N_1656,N_1168,N_1188);
nand U1657 (N_1657,N_1121,N_1324);
nor U1658 (N_1658,N_1496,N_1228);
and U1659 (N_1659,N_1007,N_1354);
nand U1660 (N_1660,N_1322,N_1348);
and U1661 (N_1661,N_1339,N_1433);
and U1662 (N_1662,N_1317,N_1265);
nor U1663 (N_1663,N_1353,N_1162);
or U1664 (N_1664,N_1397,N_1330);
and U1665 (N_1665,N_1201,N_1251);
nand U1666 (N_1666,N_1438,N_1486);
and U1667 (N_1667,N_1380,N_1223);
or U1668 (N_1668,N_1248,N_1180);
nand U1669 (N_1669,N_1139,N_1011);
or U1670 (N_1670,N_1008,N_1382);
and U1671 (N_1671,N_1346,N_1199);
nand U1672 (N_1672,N_1152,N_1303);
and U1673 (N_1673,N_1032,N_1058);
nor U1674 (N_1674,N_1239,N_1455);
nor U1675 (N_1675,N_1141,N_1084);
or U1676 (N_1676,N_1164,N_1155);
or U1677 (N_1677,N_1489,N_1340);
nor U1678 (N_1678,N_1375,N_1125);
nand U1679 (N_1679,N_1386,N_1341);
nor U1680 (N_1680,N_1425,N_1061);
and U1681 (N_1681,N_1143,N_1269);
nor U1682 (N_1682,N_1095,N_1059);
nand U1683 (N_1683,N_1421,N_1123);
and U1684 (N_1684,N_1294,N_1194);
and U1685 (N_1685,N_1247,N_1196);
nor U1686 (N_1686,N_1473,N_1107);
and U1687 (N_1687,N_1144,N_1258);
nand U1688 (N_1688,N_1282,N_1056);
nor U1689 (N_1689,N_1378,N_1181);
nand U1690 (N_1690,N_1113,N_1283);
nor U1691 (N_1691,N_1106,N_1260);
and U1692 (N_1692,N_1325,N_1246);
nand U1693 (N_1693,N_1480,N_1390);
and U1694 (N_1694,N_1279,N_1207);
nor U1695 (N_1695,N_1221,N_1224);
nand U1696 (N_1696,N_1009,N_1457);
and U1697 (N_1697,N_1310,N_1090);
and U1698 (N_1698,N_1494,N_1281);
nor U1699 (N_1699,N_1217,N_1319);
nand U1700 (N_1700,N_1175,N_1254);
and U1701 (N_1701,N_1049,N_1099);
nand U1702 (N_1702,N_1034,N_1402);
and U1703 (N_1703,N_1027,N_1476);
and U1704 (N_1704,N_1454,N_1176);
nor U1705 (N_1705,N_1033,N_1022);
nand U1706 (N_1706,N_1263,N_1040);
or U1707 (N_1707,N_1266,N_1291);
nand U1708 (N_1708,N_1343,N_1255);
nor U1709 (N_1709,N_1038,N_1376);
nor U1710 (N_1710,N_1296,N_1086);
or U1711 (N_1711,N_1165,N_1452);
nor U1712 (N_1712,N_1333,N_1206);
nor U1713 (N_1713,N_1021,N_1142);
nor U1714 (N_1714,N_1458,N_1197);
or U1715 (N_1715,N_1268,N_1445);
or U1716 (N_1716,N_1147,N_1013);
and U1717 (N_1717,N_1495,N_1148);
or U1718 (N_1718,N_1253,N_1327);
nor U1719 (N_1719,N_1358,N_1467);
nor U1720 (N_1720,N_1387,N_1243);
and U1721 (N_1721,N_1163,N_1252);
nor U1722 (N_1722,N_1242,N_1200);
xor U1723 (N_1723,N_1237,N_1389);
nor U1724 (N_1724,N_1122,N_1359);
or U1725 (N_1725,N_1300,N_1145);
and U1726 (N_1726,N_1231,N_1482);
nand U1727 (N_1727,N_1442,N_1204);
and U1728 (N_1728,N_1464,N_1499);
and U1729 (N_1729,N_1016,N_1048);
and U1730 (N_1730,N_1050,N_1091);
nor U1731 (N_1731,N_1429,N_1083);
nand U1732 (N_1732,N_1151,N_1015);
and U1733 (N_1733,N_1149,N_1087);
nor U1734 (N_1734,N_1307,N_1195);
and U1735 (N_1735,N_1089,N_1157);
and U1736 (N_1736,N_1097,N_1460);
nand U1737 (N_1737,N_1208,N_1292);
or U1738 (N_1738,N_1415,N_1426);
nand U1739 (N_1739,N_1431,N_1398);
nand U1740 (N_1740,N_1478,N_1085);
nor U1741 (N_1741,N_1014,N_1301);
or U1742 (N_1742,N_1146,N_1326);
or U1743 (N_1743,N_1140,N_1456);
nand U1744 (N_1744,N_1287,N_1238);
and U1745 (N_1745,N_1424,N_1409);
nor U1746 (N_1746,N_1046,N_1065);
or U1747 (N_1747,N_1350,N_1306);
and U1748 (N_1748,N_1368,N_1451);
or U1749 (N_1749,N_1371,N_1041);
or U1750 (N_1750,N_1484,N_1236);
and U1751 (N_1751,N_1255,N_1326);
nand U1752 (N_1752,N_1383,N_1093);
or U1753 (N_1753,N_1328,N_1014);
nand U1754 (N_1754,N_1307,N_1035);
and U1755 (N_1755,N_1338,N_1470);
or U1756 (N_1756,N_1133,N_1153);
nor U1757 (N_1757,N_1293,N_1038);
nor U1758 (N_1758,N_1005,N_1442);
and U1759 (N_1759,N_1478,N_1030);
nor U1760 (N_1760,N_1175,N_1385);
and U1761 (N_1761,N_1001,N_1096);
nand U1762 (N_1762,N_1089,N_1111);
and U1763 (N_1763,N_1244,N_1112);
nor U1764 (N_1764,N_1242,N_1493);
nor U1765 (N_1765,N_1368,N_1058);
and U1766 (N_1766,N_1082,N_1469);
or U1767 (N_1767,N_1248,N_1473);
or U1768 (N_1768,N_1291,N_1382);
or U1769 (N_1769,N_1334,N_1277);
nor U1770 (N_1770,N_1493,N_1485);
and U1771 (N_1771,N_1267,N_1253);
or U1772 (N_1772,N_1354,N_1200);
nor U1773 (N_1773,N_1176,N_1324);
or U1774 (N_1774,N_1331,N_1230);
and U1775 (N_1775,N_1045,N_1429);
nand U1776 (N_1776,N_1044,N_1323);
and U1777 (N_1777,N_1139,N_1366);
nor U1778 (N_1778,N_1185,N_1211);
and U1779 (N_1779,N_1388,N_1254);
nor U1780 (N_1780,N_1394,N_1405);
and U1781 (N_1781,N_1075,N_1245);
nand U1782 (N_1782,N_1336,N_1230);
and U1783 (N_1783,N_1408,N_1234);
and U1784 (N_1784,N_1173,N_1067);
or U1785 (N_1785,N_1162,N_1349);
or U1786 (N_1786,N_1208,N_1128);
and U1787 (N_1787,N_1155,N_1447);
and U1788 (N_1788,N_1196,N_1121);
nor U1789 (N_1789,N_1113,N_1107);
and U1790 (N_1790,N_1351,N_1214);
and U1791 (N_1791,N_1337,N_1324);
nor U1792 (N_1792,N_1030,N_1369);
nor U1793 (N_1793,N_1062,N_1379);
and U1794 (N_1794,N_1321,N_1132);
and U1795 (N_1795,N_1198,N_1379);
nand U1796 (N_1796,N_1017,N_1375);
or U1797 (N_1797,N_1160,N_1052);
and U1798 (N_1798,N_1101,N_1090);
nand U1799 (N_1799,N_1131,N_1379);
nand U1800 (N_1800,N_1422,N_1366);
nand U1801 (N_1801,N_1264,N_1000);
or U1802 (N_1802,N_1460,N_1330);
nor U1803 (N_1803,N_1367,N_1487);
nor U1804 (N_1804,N_1138,N_1216);
nand U1805 (N_1805,N_1439,N_1407);
nor U1806 (N_1806,N_1014,N_1460);
nor U1807 (N_1807,N_1492,N_1077);
and U1808 (N_1808,N_1296,N_1225);
nor U1809 (N_1809,N_1023,N_1343);
and U1810 (N_1810,N_1185,N_1035);
and U1811 (N_1811,N_1075,N_1495);
and U1812 (N_1812,N_1033,N_1405);
nor U1813 (N_1813,N_1080,N_1081);
and U1814 (N_1814,N_1000,N_1142);
or U1815 (N_1815,N_1428,N_1373);
nand U1816 (N_1816,N_1476,N_1241);
nor U1817 (N_1817,N_1403,N_1021);
nand U1818 (N_1818,N_1115,N_1283);
or U1819 (N_1819,N_1242,N_1256);
or U1820 (N_1820,N_1338,N_1111);
xor U1821 (N_1821,N_1263,N_1339);
nor U1822 (N_1822,N_1390,N_1473);
nor U1823 (N_1823,N_1333,N_1230);
nor U1824 (N_1824,N_1140,N_1413);
and U1825 (N_1825,N_1250,N_1418);
and U1826 (N_1826,N_1048,N_1256);
nand U1827 (N_1827,N_1216,N_1090);
nor U1828 (N_1828,N_1481,N_1478);
and U1829 (N_1829,N_1006,N_1494);
or U1830 (N_1830,N_1162,N_1252);
nor U1831 (N_1831,N_1174,N_1065);
nand U1832 (N_1832,N_1492,N_1457);
or U1833 (N_1833,N_1027,N_1451);
and U1834 (N_1834,N_1205,N_1409);
or U1835 (N_1835,N_1439,N_1199);
and U1836 (N_1836,N_1403,N_1414);
nand U1837 (N_1837,N_1445,N_1393);
nand U1838 (N_1838,N_1477,N_1419);
and U1839 (N_1839,N_1385,N_1214);
nor U1840 (N_1840,N_1094,N_1331);
nor U1841 (N_1841,N_1113,N_1057);
nand U1842 (N_1842,N_1280,N_1098);
nor U1843 (N_1843,N_1465,N_1002);
or U1844 (N_1844,N_1022,N_1382);
nand U1845 (N_1845,N_1156,N_1296);
nand U1846 (N_1846,N_1034,N_1176);
or U1847 (N_1847,N_1451,N_1144);
or U1848 (N_1848,N_1351,N_1489);
and U1849 (N_1849,N_1158,N_1392);
nor U1850 (N_1850,N_1283,N_1035);
or U1851 (N_1851,N_1227,N_1386);
or U1852 (N_1852,N_1169,N_1228);
nand U1853 (N_1853,N_1268,N_1020);
nand U1854 (N_1854,N_1085,N_1440);
nor U1855 (N_1855,N_1404,N_1231);
nor U1856 (N_1856,N_1085,N_1130);
nand U1857 (N_1857,N_1178,N_1419);
nand U1858 (N_1858,N_1082,N_1465);
and U1859 (N_1859,N_1469,N_1001);
nor U1860 (N_1860,N_1280,N_1335);
nor U1861 (N_1861,N_1002,N_1445);
nand U1862 (N_1862,N_1293,N_1427);
nor U1863 (N_1863,N_1007,N_1429);
or U1864 (N_1864,N_1430,N_1123);
nor U1865 (N_1865,N_1024,N_1186);
nor U1866 (N_1866,N_1275,N_1353);
nor U1867 (N_1867,N_1030,N_1015);
or U1868 (N_1868,N_1308,N_1059);
nand U1869 (N_1869,N_1230,N_1400);
and U1870 (N_1870,N_1444,N_1459);
and U1871 (N_1871,N_1150,N_1274);
and U1872 (N_1872,N_1099,N_1268);
and U1873 (N_1873,N_1170,N_1262);
nor U1874 (N_1874,N_1423,N_1231);
and U1875 (N_1875,N_1278,N_1062);
nor U1876 (N_1876,N_1347,N_1445);
and U1877 (N_1877,N_1140,N_1214);
and U1878 (N_1878,N_1253,N_1474);
nand U1879 (N_1879,N_1303,N_1012);
or U1880 (N_1880,N_1042,N_1477);
nor U1881 (N_1881,N_1345,N_1045);
and U1882 (N_1882,N_1206,N_1087);
nand U1883 (N_1883,N_1487,N_1475);
or U1884 (N_1884,N_1211,N_1178);
nor U1885 (N_1885,N_1007,N_1001);
or U1886 (N_1886,N_1406,N_1069);
nor U1887 (N_1887,N_1273,N_1328);
nand U1888 (N_1888,N_1361,N_1330);
and U1889 (N_1889,N_1105,N_1365);
nor U1890 (N_1890,N_1414,N_1490);
and U1891 (N_1891,N_1235,N_1296);
nand U1892 (N_1892,N_1208,N_1286);
and U1893 (N_1893,N_1412,N_1090);
or U1894 (N_1894,N_1332,N_1050);
nor U1895 (N_1895,N_1370,N_1124);
and U1896 (N_1896,N_1434,N_1482);
or U1897 (N_1897,N_1347,N_1115);
and U1898 (N_1898,N_1231,N_1318);
or U1899 (N_1899,N_1332,N_1436);
nor U1900 (N_1900,N_1364,N_1137);
and U1901 (N_1901,N_1045,N_1432);
or U1902 (N_1902,N_1053,N_1453);
or U1903 (N_1903,N_1246,N_1138);
and U1904 (N_1904,N_1197,N_1199);
or U1905 (N_1905,N_1193,N_1498);
nor U1906 (N_1906,N_1318,N_1013);
or U1907 (N_1907,N_1448,N_1218);
nand U1908 (N_1908,N_1156,N_1168);
nor U1909 (N_1909,N_1255,N_1177);
nor U1910 (N_1910,N_1473,N_1089);
nand U1911 (N_1911,N_1006,N_1032);
and U1912 (N_1912,N_1060,N_1007);
nor U1913 (N_1913,N_1121,N_1429);
nor U1914 (N_1914,N_1223,N_1193);
nor U1915 (N_1915,N_1050,N_1037);
or U1916 (N_1916,N_1154,N_1480);
or U1917 (N_1917,N_1423,N_1418);
and U1918 (N_1918,N_1487,N_1086);
nand U1919 (N_1919,N_1072,N_1313);
or U1920 (N_1920,N_1422,N_1159);
nor U1921 (N_1921,N_1259,N_1452);
or U1922 (N_1922,N_1452,N_1290);
or U1923 (N_1923,N_1286,N_1130);
or U1924 (N_1924,N_1236,N_1353);
or U1925 (N_1925,N_1346,N_1434);
or U1926 (N_1926,N_1239,N_1208);
nand U1927 (N_1927,N_1240,N_1151);
or U1928 (N_1928,N_1149,N_1386);
or U1929 (N_1929,N_1243,N_1487);
or U1930 (N_1930,N_1389,N_1455);
nor U1931 (N_1931,N_1048,N_1233);
or U1932 (N_1932,N_1374,N_1422);
nor U1933 (N_1933,N_1223,N_1095);
or U1934 (N_1934,N_1294,N_1001);
nand U1935 (N_1935,N_1465,N_1152);
and U1936 (N_1936,N_1498,N_1086);
nor U1937 (N_1937,N_1013,N_1374);
nor U1938 (N_1938,N_1028,N_1298);
or U1939 (N_1939,N_1158,N_1115);
or U1940 (N_1940,N_1368,N_1012);
nor U1941 (N_1941,N_1358,N_1464);
nand U1942 (N_1942,N_1477,N_1016);
nand U1943 (N_1943,N_1080,N_1078);
or U1944 (N_1944,N_1219,N_1491);
xor U1945 (N_1945,N_1362,N_1255);
nand U1946 (N_1946,N_1147,N_1252);
nor U1947 (N_1947,N_1411,N_1168);
or U1948 (N_1948,N_1066,N_1333);
or U1949 (N_1949,N_1009,N_1296);
and U1950 (N_1950,N_1114,N_1205);
or U1951 (N_1951,N_1138,N_1462);
or U1952 (N_1952,N_1093,N_1204);
nor U1953 (N_1953,N_1178,N_1354);
nor U1954 (N_1954,N_1166,N_1143);
xor U1955 (N_1955,N_1484,N_1114);
and U1956 (N_1956,N_1412,N_1301);
nor U1957 (N_1957,N_1289,N_1242);
nor U1958 (N_1958,N_1224,N_1460);
nor U1959 (N_1959,N_1343,N_1198);
or U1960 (N_1960,N_1271,N_1116);
nand U1961 (N_1961,N_1442,N_1339);
and U1962 (N_1962,N_1053,N_1131);
nand U1963 (N_1963,N_1149,N_1291);
nor U1964 (N_1964,N_1460,N_1253);
nor U1965 (N_1965,N_1031,N_1015);
nand U1966 (N_1966,N_1366,N_1356);
and U1967 (N_1967,N_1160,N_1239);
nor U1968 (N_1968,N_1314,N_1015);
nand U1969 (N_1969,N_1258,N_1193);
and U1970 (N_1970,N_1346,N_1324);
nor U1971 (N_1971,N_1131,N_1246);
and U1972 (N_1972,N_1153,N_1376);
and U1973 (N_1973,N_1050,N_1262);
or U1974 (N_1974,N_1337,N_1401);
and U1975 (N_1975,N_1439,N_1321);
nor U1976 (N_1976,N_1012,N_1083);
nand U1977 (N_1977,N_1427,N_1157);
nor U1978 (N_1978,N_1294,N_1329);
nand U1979 (N_1979,N_1407,N_1384);
and U1980 (N_1980,N_1055,N_1386);
and U1981 (N_1981,N_1341,N_1065);
nand U1982 (N_1982,N_1169,N_1133);
and U1983 (N_1983,N_1233,N_1484);
nor U1984 (N_1984,N_1400,N_1391);
nor U1985 (N_1985,N_1264,N_1402);
and U1986 (N_1986,N_1378,N_1002);
nand U1987 (N_1987,N_1455,N_1354);
or U1988 (N_1988,N_1474,N_1021);
nand U1989 (N_1989,N_1250,N_1422);
nand U1990 (N_1990,N_1148,N_1210);
and U1991 (N_1991,N_1465,N_1243);
and U1992 (N_1992,N_1471,N_1000);
nor U1993 (N_1993,N_1276,N_1494);
nor U1994 (N_1994,N_1377,N_1265);
or U1995 (N_1995,N_1066,N_1151);
nor U1996 (N_1996,N_1447,N_1199);
and U1997 (N_1997,N_1311,N_1302);
nor U1998 (N_1998,N_1450,N_1038);
nor U1999 (N_1999,N_1017,N_1309);
nor U2000 (N_2000,N_1900,N_1645);
and U2001 (N_2001,N_1802,N_1831);
nand U2002 (N_2002,N_1731,N_1924);
nor U2003 (N_2003,N_1657,N_1874);
and U2004 (N_2004,N_1991,N_1581);
or U2005 (N_2005,N_1713,N_1681);
nor U2006 (N_2006,N_1971,N_1979);
nand U2007 (N_2007,N_1764,N_1895);
or U2008 (N_2008,N_1605,N_1674);
nand U2009 (N_2009,N_1826,N_1894);
nor U2010 (N_2010,N_1663,N_1532);
xnor U2011 (N_2011,N_1509,N_1824);
nor U2012 (N_2012,N_1662,N_1568);
nand U2013 (N_2013,N_1743,N_1806);
nor U2014 (N_2014,N_1504,N_1821);
nor U2015 (N_2015,N_1520,N_1539);
and U2016 (N_2016,N_1813,N_1890);
nand U2017 (N_2017,N_1703,N_1603);
or U2018 (N_2018,N_1975,N_1592);
or U2019 (N_2019,N_1968,N_1849);
or U2020 (N_2020,N_1801,N_1667);
and U2021 (N_2021,N_1962,N_1919);
nand U2022 (N_2022,N_1763,N_1685);
nand U2023 (N_2023,N_1661,N_1948);
nand U2024 (N_2024,N_1896,N_1565);
and U2025 (N_2025,N_1954,N_1625);
nor U2026 (N_2026,N_1993,N_1814);
nand U2027 (N_2027,N_1519,N_1771);
and U2028 (N_2028,N_1629,N_1669);
nand U2029 (N_2029,N_1654,N_1745);
or U2030 (N_2030,N_1728,N_1545);
nor U2031 (N_2031,N_1570,N_1827);
or U2032 (N_2032,N_1778,N_1647);
and U2033 (N_2033,N_1637,N_1877);
nor U2034 (N_2034,N_1698,N_1952);
and U2035 (N_2035,N_1977,N_1988);
or U2036 (N_2036,N_1942,N_1632);
and U2037 (N_2037,N_1766,N_1705);
nor U2038 (N_2038,N_1733,N_1571);
and U2039 (N_2039,N_1558,N_1535);
nand U2040 (N_2040,N_1641,N_1950);
nor U2041 (N_2041,N_1867,N_1583);
nand U2042 (N_2042,N_1501,N_1747);
and U2043 (N_2043,N_1578,N_1823);
xnor U2044 (N_2044,N_1837,N_1816);
and U2045 (N_2045,N_1608,N_1903);
or U2046 (N_2046,N_1609,N_1527);
nor U2047 (N_2047,N_1542,N_1686);
or U2048 (N_2048,N_1836,N_1744);
nand U2049 (N_2049,N_1712,N_1742);
nor U2050 (N_2050,N_1631,N_1636);
nor U2051 (N_2051,N_1708,N_1951);
nand U2052 (N_2052,N_1739,N_1551);
nand U2053 (N_2053,N_1999,N_1798);
or U2054 (N_2054,N_1815,N_1678);
and U2055 (N_2055,N_1844,N_1723);
nand U2056 (N_2056,N_1648,N_1664);
or U2057 (N_2057,N_1875,N_1704);
nand U2058 (N_2058,N_1537,N_1619);
nor U2059 (N_2059,N_1659,N_1893);
nand U2060 (N_2060,N_1671,N_1762);
or U2061 (N_2061,N_1920,N_1553);
or U2062 (N_2062,N_1853,N_1697);
or U2063 (N_2063,N_1575,N_1561);
and U2064 (N_2064,N_1595,N_1524);
and U2065 (N_2065,N_1732,N_1953);
and U2066 (N_2066,N_1923,N_1774);
and U2067 (N_2067,N_1635,N_1935);
nor U2068 (N_2068,N_1508,N_1984);
nand U2069 (N_2069,N_1755,N_1886);
and U2070 (N_2070,N_1630,N_1850);
and U2071 (N_2071,N_1871,N_1576);
nor U2072 (N_2072,N_1819,N_1973);
and U2073 (N_2073,N_1714,N_1624);
xor U2074 (N_2074,N_1696,N_1792);
nand U2075 (N_2075,N_1758,N_1695);
and U2076 (N_2076,N_1925,N_1776);
nor U2077 (N_2077,N_1722,N_1868);
and U2078 (N_2078,N_1775,N_1756);
or U2079 (N_2079,N_1773,N_1549);
nand U2080 (N_2080,N_1721,N_1869);
nand U2081 (N_2081,N_1932,N_1986);
nor U2082 (N_2082,N_1585,N_1794);
nand U2083 (N_2083,N_1516,N_1943);
and U2084 (N_2084,N_1599,N_1502);
or U2085 (N_2085,N_1807,N_1596);
nand U2086 (N_2086,N_1682,N_1781);
or U2087 (N_2087,N_1547,N_1769);
nor U2088 (N_2088,N_1691,N_1512);
and U2089 (N_2089,N_1729,N_1891);
and U2090 (N_2090,N_1618,N_1761);
nand U2091 (N_2091,N_1934,N_1963);
or U2092 (N_2092,N_1767,N_1646);
or U2093 (N_2093,N_1848,N_1960);
nand U2094 (N_2094,N_1898,N_1670);
xor U2095 (N_2095,N_1878,N_1857);
nor U2096 (N_2096,N_1944,N_1974);
nor U2097 (N_2097,N_1789,N_1799);
nand U2098 (N_2098,N_1525,N_1530);
nor U2099 (N_2099,N_1846,N_1909);
nor U2100 (N_2100,N_1959,N_1796);
nand U2101 (N_2101,N_1779,N_1843);
and U2102 (N_2102,N_1594,N_1786);
and U2103 (N_2103,N_1899,N_1741);
nand U2104 (N_2104,N_1562,N_1882);
or U2105 (N_2105,N_1638,N_1734);
or U2106 (N_2106,N_1680,N_1990);
nor U2107 (N_2107,N_1817,N_1690);
nor U2108 (N_2108,N_1727,N_1737);
nand U2109 (N_2109,N_1969,N_1892);
xnor U2110 (N_2110,N_1926,N_1677);
nand U2111 (N_2111,N_1910,N_1863);
nand U2112 (N_2112,N_1541,N_1679);
and U2113 (N_2113,N_1811,N_1835);
or U2114 (N_2114,N_1995,N_1621);
or U2115 (N_2115,N_1666,N_1534);
or U2116 (N_2116,N_1901,N_1675);
nor U2117 (N_2117,N_1724,N_1538);
nand U2118 (N_2118,N_1511,N_1945);
and U2119 (N_2119,N_1665,N_1845);
or U2120 (N_2120,N_1966,N_1555);
xor U2121 (N_2121,N_1589,N_1876);
and U2122 (N_2122,N_1569,N_1611);
or U2123 (N_2123,N_1860,N_1548);
and U2124 (N_2124,N_1588,N_1804);
nand U2125 (N_2125,N_1726,N_1812);
nand U2126 (N_2126,N_1644,N_1964);
and U2127 (N_2127,N_1917,N_1828);
nor U2128 (N_2128,N_1760,N_1870);
xor U2129 (N_2129,N_1556,N_1614);
nor U2130 (N_2130,N_1607,N_1597);
and U2131 (N_2131,N_1840,N_1694);
nor U2132 (N_2132,N_1572,N_1692);
nand U2133 (N_2133,N_1579,N_1683);
or U2134 (N_2134,N_1655,N_1980);
nor U2135 (N_2135,N_1858,N_1718);
and U2136 (N_2136,N_1559,N_1883);
and U2137 (N_2137,N_1866,N_1930);
or U2138 (N_2138,N_1981,N_1931);
nor U2139 (N_2139,N_1855,N_1546);
or U2140 (N_2140,N_1830,N_1985);
or U2141 (N_2141,N_1591,N_1955);
and U2142 (N_2142,N_1780,N_1639);
nand U2143 (N_2143,N_1693,N_1617);
or U2144 (N_2144,N_1808,N_1822);
and U2145 (N_2145,N_1939,N_1790);
nand U2146 (N_2146,N_1753,N_1913);
nand U2147 (N_2147,N_1847,N_1649);
or U2148 (N_2148,N_1716,N_1918);
or U2149 (N_2149,N_1751,N_1584);
nor U2150 (N_2150,N_1526,N_1515);
or U2151 (N_2151,N_1795,N_1933);
nand U2152 (N_2152,N_1938,N_1998);
nor U2153 (N_2153,N_1916,N_1908);
or U2154 (N_2154,N_1543,N_1772);
and U2155 (N_2155,N_1905,N_1967);
nor U2156 (N_2156,N_1702,N_1533);
and U2157 (N_2157,N_1521,N_1622);
and U2158 (N_2158,N_1859,N_1841);
or U2159 (N_2159,N_1805,N_1862);
and U2160 (N_2160,N_1921,N_1904);
nand U2161 (N_2161,N_1593,N_1915);
nor U2162 (N_2162,N_1707,N_1554);
nand U2163 (N_2163,N_1610,N_1616);
or U2164 (N_2164,N_1660,N_1518);
and U2165 (N_2165,N_1884,N_1937);
or U2166 (N_2166,N_1522,N_1582);
or U2167 (N_2167,N_1577,N_1650);
and U2168 (N_2168,N_1927,N_1791);
nor U2169 (N_2169,N_1627,N_1961);
nand U2170 (N_2170,N_1709,N_1580);
and U2171 (N_2171,N_1958,N_1688);
or U2172 (N_2172,N_1834,N_1528);
nor U2173 (N_2173,N_1606,N_1989);
nand U2174 (N_2174,N_1689,N_1566);
or U2175 (N_2175,N_1613,N_1851);
nor U2176 (N_2176,N_1861,N_1784);
or U2177 (N_2177,N_1803,N_1972);
nand U2178 (N_2178,N_1914,N_1782);
or U2179 (N_2179,N_1601,N_1873);
nor U2180 (N_2180,N_1949,N_1941);
nor U2181 (N_2181,N_1736,N_1902);
and U2182 (N_2182,N_1982,N_1651);
nand U2183 (N_2183,N_1626,N_1500);
nand U2184 (N_2184,N_1672,N_1765);
and U2185 (N_2185,N_1946,N_1656);
nor U2186 (N_2186,N_1852,N_1623);
nor U2187 (N_2187,N_1720,N_1740);
or U2188 (N_2188,N_1947,N_1643);
or U2189 (N_2189,N_1864,N_1965);
nor U2190 (N_2190,N_1604,N_1996);
nor U2191 (N_2191,N_1881,N_1560);
nor U2192 (N_2192,N_1505,N_1701);
and U2193 (N_2193,N_1800,N_1983);
and U2194 (N_2194,N_1897,N_1587);
nor U2195 (N_2195,N_1785,N_1970);
nand U2196 (N_2196,N_1563,N_1880);
nand U2197 (N_2197,N_1829,N_1717);
or U2198 (N_2198,N_1749,N_1768);
or U2199 (N_2199,N_1906,N_1658);
nor U2200 (N_2200,N_1872,N_1992);
and U2201 (N_2201,N_1940,N_1503);
or U2202 (N_2202,N_1820,N_1818);
nor U2203 (N_2203,N_1653,N_1600);
nand U2204 (N_2204,N_1706,N_1976);
or U2205 (N_2205,N_1633,N_1652);
nand U2206 (N_2206,N_1809,N_1833);
or U2207 (N_2207,N_1907,N_1531);
nand U2208 (N_2208,N_1770,N_1810);
nand U2209 (N_2209,N_1911,N_1725);
nor U2210 (N_2210,N_1738,N_1987);
nor U2211 (N_2211,N_1719,N_1517);
and U2212 (N_2212,N_1620,N_1787);
or U2213 (N_2213,N_1676,N_1540);
nand U2214 (N_2214,N_1825,N_1957);
nor U2215 (N_2215,N_1842,N_1839);
or U2216 (N_2216,N_1832,N_1564);
nor U2217 (N_2217,N_1634,N_1668);
and U2218 (N_2218,N_1752,N_1759);
or U2219 (N_2219,N_1615,N_1567);
or U2220 (N_2220,N_1889,N_1888);
and U2221 (N_2221,N_1673,N_1838);
nor U2222 (N_2222,N_1710,N_1590);
nor U2223 (N_2223,N_1865,N_1557);
nand U2224 (N_2224,N_1552,N_1523);
xor U2225 (N_2225,N_1687,N_1628);
or U2226 (N_2226,N_1856,N_1550);
nor U2227 (N_2227,N_1797,N_1885);
and U2228 (N_2228,N_1956,N_1715);
nand U2229 (N_2229,N_1912,N_1929);
nor U2230 (N_2230,N_1684,N_1586);
and U2231 (N_2231,N_1750,N_1612);
or U2232 (N_2232,N_1536,N_1978);
nor U2233 (N_2233,N_1854,N_1699);
or U2234 (N_2234,N_1514,N_1783);
xor U2235 (N_2235,N_1793,N_1602);
and U2236 (N_2236,N_1598,N_1513);
nand U2237 (N_2237,N_1994,N_1640);
nor U2238 (N_2238,N_1700,N_1997);
or U2239 (N_2239,N_1748,N_1510);
nor U2240 (N_2240,N_1544,N_1928);
and U2241 (N_2241,N_1507,N_1573);
nor U2242 (N_2242,N_1746,N_1711);
and U2243 (N_2243,N_1574,N_1754);
nor U2244 (N_2244,N_1879,N_1757);
or U2245 (N_2245,N_1642,N_1777);
nand U2246 (N_2246,N_1887,N_1788);
nand U2247 (N_2247,N_1529,N_1936);
nand U2248 (N_2248,N_1922,N_1735);
and U2249 (N_2249,N_1730,N_1506);
and U2250 (N_2250,N_1960,N_1610);
and U2251 (N_2251,N_1667,N_1739);
or U2252 (N_2252,N_1537,N_1633);
and U2253 (N_2253,N_1801,N_1852);
nor U2254 (N_2254,N_1757,N_1705);
or U2255 (N_2255,N_1998,N_1951);
nand U2256 (N_2256,N_1589,N_1553);
or U2257 (N_2257,N_1988,N_1696);
nor U2258 (N_2258,N_1524,N_1630);
or U2259 (N_2259,N_1606,N_1634);
or U2260 (N_2260,N_1939,N_1596);
or U2261 (N_2261,N_1728,N_1667);
nand U2262 (N_2262,N_1776,N_1504);
nor U2263 (N_2263,N_1618,N_1516);
nor U2264 (N_2264,N_1999,N_1738);
and U2265 (N_2265,N_1998,N_1746);
or U2266 (N_2266,N_1572,N_1844);
and U2267 (N_2267,N_1989,N_1708);
and U2268 (N_2268,N_1522,N_1514);
nand U2269 (N_2269,N_1970,N_1703);
nor U2270 (N_2270,N_1817,N_1751);
nor U2271 (N_2271,N_1610,N_1889);
nand U2272 (N_2272,N_1748,N_1840);
and U2273 (N_2273,N_1981,N_1973);
nor U2274 (N_2274,N_1812,N_1999);
and U2275 (N_2275,N_1528,N_1786);
nand U2276 (N_2276,N_1642,N_1906);
or U2277 (N_2277,N_1726,N_1983);
nand U2278 (N_2278,N_1848,N_1687);
and U2279 (N_2279,N_1528,N_1572);
or U2280 (N_2280,N_1557,N_1773);
xnor U2281 (N_2281,N_1502,N_1907);
and U2282 (N_2282,N_1906,N_1767);
nand U2283 (N_2283,N_1725,N_1715);
and U2284 (N_2284,N_1787,N_1903);
and U2285 (N_2285,N_1972,N_1926);
and U2286 (N_2286,N_1983,N_1783);
nand U2287 (N_2287,N_1952,N_1632);
and U2288 (N_2288,N_1932,N_1818);
or U2289 (N_2289,N_1514,N_1517);
nand U2290 (N_2290,N_1861,N_1853);
or U2291 (N_2291,N_1501,N_1771);
nand U2292 (N_2292,N_1833,N_1547);
nor U2293 (N_2293,N_1723,N_1679);
nor U2294 (N_2294,N_1576,N_1932);
nand U2295 (N_2295,N_1795,N_1734);
nand U2296 (N_2296,N_1820,N_1827);
and U2297 (N_2297,N_1956,N_1695);
or U2298 (N_2298,N_1962,N_1807);
or U2299 (N_2299,N_1713,N_1726);
or U2300 (N_2300,N_1812,N_1550);
nor U2301 (N_2301,N_1695,N_1986);
and U2302 (N_2302,N_1547,N_1831);
nor U2303 (N_2303,N_1553,N_1947);
nand U2304 (N_2304,N_1607,N_1684);
nand U2305 (N_2305,N_1705,N_1880);
xnor U2306 (N_2306,N_1929,N_1566);
nor U2307 (N_2307,N_1737,N_1575);
nor U2308 (N_2308,N_1683,N_1737);
or U2309 (N_2309,N_1881,N_1688);
and U2310 (N_2310,N_1922,N_1794);
nor U2311 (N_2311,N_1582,N_1844);
nor U2312 (N_2312,N_1768,N_1697);
or U2313 (N_2313,N_1599,N_1854);
xnor U2314 (N_2314,N_1605,N_1675);
and U2315 (N_2315,N_1951,N_1939);
or U2316 (N_2316,N_1966,N_1855);
and U2317 (N_2317,N_1550,N_1626);
nand U2318 (N_2318,N_1851,N_1644);
and U2319 (N_2319,N_1874,N_1669);
and U2320 (N_2320,N_1534,N_1711);
and U2321 (N_2321,N_1742,N_1719);
nor U2322 (N_2322,N_1775,N_1766);
nor U2323 (N_2323,N_1799,N_1635);
or U2324 (N_2324,N_1516,N_1736);
and U2325 (N_2325,N_1821,N_1974);
or U2326 (N_2326,N_1516,N_1740);
nor U2327 (N_2327,N_1748,N_1920);
or U2328 (N_2328,N_1516,N_1771);
nand U2329 (N_2329,N_1748,N_1821);
nand U2330 (N_2330,N_1929,N_1953);
and U2331 (N_2331,N_1964,N_1724);
and U2332 (N_2332,N_1759,N_1901);
and U2333 (N_2333,N_1859,N_1519);
or U2334 (N_2334,N_1601,N_1683);
nor U2335 (N_2335,N_1514,N_1558);
xnor U2336 (N_2336,N_1845,N_1676);
and U2337 (N_2337,N_1797,N_1783);
and U2338 (N_2338,N_1923,N_1714);
xor U2339 (N_2339,N_1550,N_1822);
nand U2340 (N_2340,N_1892,N_1661);
nand U2341 (N_2341,N_1728,N_1677);
nand U2342 (N_2342,N_1856,N_1953);
and U2343 (N_2343,N_1982,N_1609);
or U2344 (N_2344,N_1775,N_1740);
nand U2345 (N_2345,N_1821,N_1718);
and U2346 (N_2346,N_1892,N_1960);
nand U2347 (N_2347,N_1924,N_1635);
nand U2348 (N_2348,N_1608,N_1981);
nand U2349 (N_2349,N_1868,N_1933);
and U2350 (N_2350,N_1513,N_1961);
and U2351 (N_2351,N_1947,N_1816);
nand U2352 (N_2352,N_1529,N_1743);
nand U2353 (N_2353,N_1553,N_1654);
and U2354 (N_2354,N_1856,N_1738);
and U2355 (N_2355,N_1697,N_1842);
nand U2356 (N_2356,N_1866,N_1902);
nand U2357 (N_2357,N_1508,N_1712);
xor U2358 (N_2358,N_1976,N_1595);
and U2359 (N_2359,N_1692,N_1752);
or U2360 (N_2360,N_1728,N_1689);
nand U2361 (N_2361,N_1924,N_1907);
and U2362 (N_2362,N_1944,N_1628);
nand U2363 (N_2363,N_1745,N_1882);
xor U2364 (N_2364,N_1728,N_1619);
or U2365 (N_2365,N_1851,N_1833);
nand U2366 (N_2366,N_1811,N_1568);
nand U2367 (N_2367,N_1652,N_1615);
nor U2368 (N_2368,N_1736,N_1570);
nor U2369 (N_2369,N_1669,N_1628);
nor U2370 (N_2370,N_1985,N_1839);
nand U2371 (N_2371,N_1887,N_1761);
or U2372 (N_2372,N_1527,N_1752);
nor U2373 (N_2373,N_1960,N_1713);
and U2374 (N_2374,N_1988,N_1727);
or U2375 (N_2375,N_1616,N_1544);
nor U2376 (N_2376,N_1662,N_1957);
nor U2377 (N_2377,N_1952,N_1979);
nand U2378 (N_2378,N_1704,N_1991);
and U2379 (N_2379,N_1731,N_1980);
nand U2380 (N_2380,N_1995,N_1925);
nor U2381 (N_2381,N_1645,N_1774);
or U2382 (N_2382,N_1724,N_1638);
and U2383 (N_2383,N_1617,N_1599);
nor U2384 (N_2384,N_1933,N_1908);
and U2385 (N_2385,N_1925,N_1881);
nand U2386 (N_2386,N_1506,N_1549);
and U2387 (N_2387,N_1992,N_1863);
and U2388 (N_2388,N_1504,N_1680);
or U2389 (N_2389,N_1831,N_1647);
and U2390 (N_2390,N_1686,N_1844);
nor U2391 (N_2391,N_1552,N_1706);
and U2392 (N_2392,N_1885,N_1892);
or U2393 (N_2393,N_1891,N_1937);
nand U2394 (N_2394,N_1986,N_1691);
nand U2395 (N_2395,N_1549,N_1584);
or U2396 (N_2396,N_1974,N_1878);
nor U2397 (N_2397,N_1642,N_1952);
or U2398 (N_2398,N_1579,N_1926);
or U2399 (N_2399,N_1920,N_1974);
nor U2400 (N_2400,N_1864,N_1891);
and U2401 (N_2401,N_1900,N_1893);
or U2402 (N_2402,N_1906,N_1511);
nand U2403 (N_2403,N_1925,N_1950);
nor U2404 (N_2404,N_1884,N_1613);
nor U2405 (N_2405,N_1967,N_1977);
and U2406 (N_2406,N_1706,N_1513);
or U2407 (N_2407,N_1832,N_1954);
and U2408 (N_2408,N_1596,N_1877);
and U2409 (N_2409,N_1899,N_1567);
nand U2410 (N_2410,N_1693,N_1820);
nor U2411 (N_2411,N_1519,N_1728);
nand U2412 (N_2412,N_1717,N_1567);
or U2413 (N_2413,N_1668,N_1956);
nand U2414 (N_2414,N_1994,N_1762);
nor U2415 (N_2415,N_1573,N_1872);
and U2416 (N_2416,N_1735,N_1639);
nor U2417 (N_2417,N_1633,N_1700);
nand U2418 (N_2418,N_1544,N_1531);
nor U2419 (N_2419,N_1632,N_1924);
xnor U2420 (N_2420,N_1773,N_1709);
or U2421 (N_2421,N_1890,N_1584);
nor U2422 (N_2422,N_1627,N_1917);
or U2423 (N_2423,N_1818,N_1624);
nor U2424 (N_2424,N_1715,N_1519);
and U2425 (N_2425,N_1610,N_1679);
nand U2426 (N_2426,N_1813,N_1937);
xnor U2427 (N_2427,N_1637,N_1973);
or U2428 (N_2428,N_1945,N_1923);
nor U2429 (N_2429,N_1837,N_1850);
and U2430 (N_2430,N_1536,N_1648);
or U2431 (N_2431,N_1871,N_1983);
and U2432 (N_2432,N_1568,N_1608);
and U2433 (N_2433,N_1686,N_1572);
and U2434 (N_2434,N_1934,N_1601);
nand U2435 (N_2435,N_1822,N_1976);
and U2436 (N_2436,N_1585,N_1936);
nor U2437 (N_2437,N_1598,N_1762);
and U2438 (N_2438,N_1878,N_1855);
nand U2439 (N_2439,N_1982,N_1537);
or U2440 (N_2440,N_1772,N_1753);
xnor U2441 (N_2441,N_1901,N_1946);
and U2442 (N_2442,N_1962,N_1544);
and U2443 (N_2443,N_1663,N_1764);
or U2444 (N_2444,N_1980,N_1896);
and U2445 (N_2445,N_1641,N_1657);
or U2446 (N_2446,N_1592,N_1721);
xnor U2447 (N_2447,N_1825,N_1992);
nor U2448 (N_2448,N_1833,N_1556);
and U2449 (N_2449,N_1805,N_1717);
nor U2450 (N_2450,N_1665,N_1812);
xnor U2451 (N_2451,N_1819,N_1723);
or U2452 (N_2452,N_1899,N_1687);
and U2453 (N_2453,N_1753,N_1834);
or U2454 (N_2454,N_1949,N_1789);
and U2455 (N_2455,N_1966,N_1795);
or U2456 (N_2456,N_1989,N_1665);
and U2457 (N_2457,N_1678,N_1756);
and U2458 (N_2458,N_1798,N_1751);
nor U2459 (N_2459,N_1577,N_1884);
and U2460 (N_2460,N_1854,N_1752);
and U2461 (N_2461,N_1733,N_1823);
nand U2462 (N_2462,N_1974,N_1586);
and U2463 (N_2463,N_1687,N_1958);
xor U2464 (N_2464,N_1870,N_1762);
or U2465 (N_2465,N_1713,N_1901);
or U2466 (N_2466,N_1500,N_1710);
or U2467 (N_2467,N_1544,N_1693);
or U2468 (N_2468,N_1618,N_1631);
nor U2469 (N_2469,N_1507,N_1946);
nor U2470 (N_2470,N_1560,N_1704);
and U2471 (N_2471,N_1640,N_1542);
and U2472 (N_2472,N_1706,N_1841);
or U2473 (N_2473,N_1852,N_1948);
or U2474 (N_2474,N_1774,N_1998);
nand U2475 (N_2475,N_1904,N_1708);
nor U2476 (N_2476,N_1569,N_1934);
nand U2477 (N_2477,N_1986,N_1543);
xnor U2478 (N_2478,N_1642,N_1844);
nand U2479 (N_2479,N_1690,N_1700);
or U2480 (N_2480,N_1502,N_1812);
nand U2481 (N_2481,N_1529,N_1701);
or U2482 (N_2482,N_1839,N_1502);
and U2483 (N_2483,N_1608,N_1864);
and U2484 (N_2484,N_1943,N_1606);
nor U2485 (N_2485,N_1928,N_1851);
or U2486 (N_2486,N_1622,N_1730);
and U2487 (N_2487,N_1537,N_1734);
nor U2488 (N_2488,N_1958,N_1599);
or U2489 (N_2489,N_1687,N_1885);
or U2490 (N_2490,N_1612,N_1596);
and U2491 (N_2491,N_1520,N_1703);
and U2492 (N_2492,N_1539,N_1572);
nor U2493 (N_2493,N_1612,N_1886);
nor U2494 (N_2494,N_1543,N_1729);
nand U2495 (N_2495,N_1721,N_1635);
and U2496 (N_2496,N_1640,N_1578);
nor U2497 (N_2497,N_1993,N_1651);
nor U2498 (N_2498,N_1548,N_1552);
or U2499 (N_2499,N_1522,N_1989);
or U2500 (N_2500,N_2212,N_2455);
xor U2501 (N_2501,N_2311,N_2190);
nor U2502 (N_2502,N_2316,N_2430);
nand U2503 (N_2503,N_2437,N_2009);
or U2504 (N_2504,N_2420,N_2302);
xnor U2505 (N_2505,N_2000,N_2098);
nor U2506 (N_2506,N_2491,N_2135);
or U2507 (N_2507,N_2165,N_2072);
nor U2508 (N_2508,N_2277,N_2206);
nand U2509 (N_2509,N_2419,N_2363);
nor U2510 (N_2510,N_2450,N_2287);
or U2511 (N_2511,N_2228,N_2324);
nand U2512 (N_2512,N_2063,N_2344);
and U2513 (N_2513,N_2458,N_2162);
and U2514 (N_2514,N_2319,N_2096);
or U2515 (N_2515,N_2275,N_2456);
or U2516 (N_2516,N_2118,N_2390);
nand U2517 (N_2517,N_2409,N_2156);
or U2518 (N_2518,N_2066,N_2236);
nor U2519 (N_2519,N_2052,N_2478);
nand U2520 (N_2520,N_2237,N_2352);
nor U2521 (N_2521,N_2106,N_2073);
or U2522 (N_2522,N_2358,N_2086);
and U2523 (N_2523,N_2123,N_2383);
nand U2524 (N_2524,N_2153,N_2188);
nand U2525 (N_2525,N_2137,N_2305);
nor U2526 (N_2526,N_2029,N_2253);
or U2527 (N_2527,N_2464,N_2360);
nand U2528 (N_2528,N_2496,N_2145);
nor U2529 (N_2529,N_2293,N_2020);
or U2530 (N_2530,N_2144,N_2048);
nor U2531 (N_2531,N_2278,N_2315);
nand U2532 (N_2532,N_2076,N_2421);
nand U2533 (N_2533,N_2095,N_2012);
nand U2534 (N_2534,N_2022,N_2025);
nor U2535 (N_2535,N_2428,N_2151);
or U2536 (N_2536,N_2157,N_2424);
nand U2537 (N_2537,N_2308,N_2047);
or U2538 (N_2538,N_2323,N_2097);
or U2539 (N_2539,N_2267,N_2355);
nor U2540 (N_2540,N_2062,N_2480);
and U2541 (N_2541,N_2032,N_2349);
nand U2542 (N_2542,N_2172,N_2265);
nor U2543 (N_2543,N_2446,N_2069);
or U2544 (N_2544,N_2109,N_2329);
nor U2545 (N_2545,N_2138,N_2250);
nor U2546 (N_2546,N_2413,N_2005);
nand U2547 (N_2547,N_2330,N_2297);
and U2548 (N_2548,N_2334,N_2122);
or U2549 (N_2549,N_2040,N_2343);
nor U2550 (N_2550,N_2241,N_2093);
nand U2551 (N_2551,N_2353,N_2373);
nor U2552 (N_2552,N_2403,N_2264);
or U2553 (N_2553,N_2199,N_2222);
nand U2554 (N_2554,N_2204,N_2402);
nand U2555 (N_2555,N_2408,N_2395);
or U2556 (N_2556,N_2028,N_2415);
nor U2557 (N_2557,N_2434,N_2339);
nor U2558 (N_2558,N_2386,N_2271);
or U2559 (N_2559,N_2024,N_2036);
and U2560 (N_2560,N_2218,N_2488);
or U2561 (N_2561,N_2479,N_2059);
or U2562 (N_2562,N_2201,N_2083);
nand U2563 (N_2563,N_2061,N_2307);
and U2564 (N_2564,N_2008,N_2259);
nand U2565 (N_2565,N_2019,N_2078);
or U2566 (N_2566,N_2459,N_2198);
or U2567 (N_2567,N_2382,N_2171);
and U2568 (N_2568,N_2336,N_2080);
or U2569 (N_2569,N_2341,N_2276);
nor U2570 (N_2570,N_2077,N_2202);
and U2571 (N_2571,N_2010,N_2346);
or U2572 (N_2572,N_2347,N_2159);
nor U2573 (N_2573,N_2294,N_2401);
and U2574 (N_2574,N_2033,N_2404);
nand U2575 (N_2575,N_2070,N_2013);
nor U2576 (N_2576,N_2089,N_2388);
or U2577 (N_2577,N_2107,N_2291);
nand U2578 (N_2578,N_2467,N_2397);
or U2579 (N_2579,N_2499,N_2181);
nand U2580 (N_2580,N_2104,N_2440);
and U2581 (N_2581,N_2435,N_2414);
or U2582 (N_2582,N_2379,N_2282);
nand U2583 (N_2583,N_2231,N_2444);
nand U2584 (N_2584,N_2189,N_2152);
or U2585 (N_2585,N_2274,N_2090);
nand U2586 (N_2586,N_2211,N_2389);
and U2587 (N_2587,N_2163,N_2304);
or U2588 (N_2588,N_2303,N_2494);
nor U2589 (N_2589,N_2338,N_2006);
or U2590 (N_2590,N_2067,N_2313);
and U2591 (N_2591,N_2015,N_2247);
or U2592 (N_2592,N_2233,N_2016);
nor U2593 (N_2593,N_2234,N_2454);
nor U2594 (N_2594,N_2057,N_2217);
nand U2595 (N_2595,N_2261,N_2405);
nand U2596 (N_2596,N_2179,N_2001);
nor U2597 (N_2597,N_2257,N_2037);
and U2598 (N_2598,N_2492,N_2101);
and U2599 (N_2599,N_2485,N_2200);
and U2600 (N_2600,N_2372,N_2134);
or U2601 (N_2601,N_2442,N_2045);
nor U2602 (N_2602,N_2387,N_2108);
nand U2603 (N_2603,N_2481,N_2018);
nand U2604 (N_2604,N_2381,N_2238);
nand U2605 (N_2605,N_2273,N_2486);
nand U2606 (N_2606,N_2342,N_2164);
or U2607 (N_2607,N_2411,N_2457);
or U2608 (N_2608,N_2088,N_2490);
or U2609 (N_2609,N_2392,N_2380);
and U2610 (N_2610,N_2367,N_2141);
nand U2611 (N_2611,N_2416,N_2384);
nand U2612 (N_2612,N_2180,N_2474);
or U2613 (N_2613,N_2429,N_2143);
and U2614 (N_2614,N_2394,N_2406);
xnor U2615 (N_2615,N_2223,N_2055);
nor U2616 (N_2616,N_2116,N_2262);
nand U2617 (N_2617,N_2128,N_2468);
nor U2618 (N_2618,N_2209,N_2205);
or U2619 (N_2619,N_2482,N_2364);
or U2620 (N_2620,N_2325,N_2023);
nor U2621 (N_2621,N_2493,N_2301);
xnor U2622 (N_2622,N_2445,N_2105);
nand U2623 (N_2623,N_2284,N_2350);
nand U2624 (N_2624,N_2431,N_2131);
nor U2625 (N_2625,N_2487,N_2299);
and U2626 (N_2626,N_2232,N_2017);
or U2627 (N_2627,N_2438,N_2044);
and U2628 (N_2628,N_2327,N_2071);
or U2629 (N_2629,N_2176,N_2099);
nor U2630 (N_2630,N_2082,N_2225);
or U2631 (N_2631,N_2377,N_2398);
or U2632 (N_2632,N_2322,N_2150);
nand U2633 (N_2633,N_2192,N_2340);
nor U2634 (N_2634,N_2331,N_2207);
or U2635 (N_2635,N_2208,N_2195);
nor U2636 (N_2636,N_2014,N_2193);
or U2637 (N_2637,N_2348,N_2079);
and U2638 (N_2638,N_2436,N_2332);
nor U2639 (N_2639,N_2391,N_2053);
and U2640 (N_2640,N_2248,N_2425);
and U2641 (N_2641,N_2357,N_2443);
or U2642 (N_2642,N_2058,N_2177);
and U2643 (N_2643,N_2452,N_2281);
and U2644 (N_2644,N_2043,N_2385);
nor U2645 (N_2645,N_2127,N_2147);
nor U2646 (N_2646,N_2423,N_2256);
nor U2647 (N_2647,N_2448,N_2003);
and U2648 (N_2648,N_2412,N_2031);
or U2649 (N_2649,N_2114,N_2251);
and U2650 (N_2650,N_2060,N_2451);
and U2651 (N_2651,N_2466,N_2170);
xnor U2652 (N_2652,N_2258,N_2132);
nand U2653 (N_2653,N_2174,N_2469);
or U2654 (N_2654,N_2167,N_2084);
nor U2655 (N_2655,N_2146,N_2102);
or U2656 (N_2656,N_2300,N_2449);
and U2657 (N_2657,N_2161,N_2136);
nor U2658 (N_2658,N_2441,N_2187);
nand U2659 (N_2659,N_2244,N_2113);
and U2660 (N_2660,N_2354,N_2166);
nor U2661 (N_2661,N_2268,N_2473);
nor U2662 (N_2662,N_2475,N_2290);
nand U2663 (N_2663,N_2288,N_2042);
nand U2664 (N_2664,N_2068,N_2011);
and U2665 (N_2665,N_2214,N_2002);
and U2666 (N_2666,N_2056,N_2393);
nand U2667 (N_2667,N_2286,N_2169);
nor U2668 (N_2668,N_2314,N_2034);
nand U2669 (N_2669,N_2368,N_2220);
or U2670 (N_2670,N_2280,N_2260);
and U2671 (N_2671,N_2312,N_2221);
or U2672 (N_2672,N_2476,N_2194);
and U2673 (N_2673,N_2410,N_2463);
nand U2674 (N_2674,N_2175,N_2465);
or U2675 (N_2675,N_2270,N_2335);
and U2676 (N_2676,N_2337,N_2119);
nand U2677 (N_2677,N_2054,N_2252);
nand U2678 (N_2678,N_2115,N_2117);
nand U2679 (N_2679,N_2407,N_2296);
nand U2680 (N_2680,N_2472,N_2110);
and U2681 (N_2681,N_2453,N_2439);
nand U2682 (N_2682,N_2320,N_2112);
and U2683 (N_2683,N_2263,N_2046);
nor U2684 (N_2684,N_2471,N_2085);
and U2685 (N_2685,N_2378,N_2210);
nand U2686 (N_2686,N_2292,N_2168);
xnor U2687 (N_2687,N_2255,N_2038);
or U2688 (N_2688,N_2216,N_2422);
nor U2689 (N_2689,N_2362,N_2140);
nand U2690 (N_2690,N_2139,N_2470);
and U2691 (N_2691,N_2155,N_2371);
or U2692 (N_2692,N_2120,N_2447);
nand U2693 (N_2693,N_2495,N_2149);
and U2694 (N_2694,N_2142,N_2121);
nand U2695 (N_2695,N_2091,N_2460);
nor U2696 (N_2696,N_2326,N_2186);
or U2697 (N_2697,N_2087,N_2432);
nand U2698 (N_2698,N_2483,N_2160);
or U2699 (N_2699,N_2396,N_2092);
or U2700 (N_2700,N_2100,N_2285);
nand U2701 (N_2701,N_2184,N_2370);
nor U2702 (N_2702,N_2185,N_2249);
nand U2703 (N_2703,N_2345,N_2213);
or U2704 (N_2704,N_2321,N_2369);
and U2705 (N_2705,N_2427,N_2298);
nor U2706 (N_2706,N_2178,N_2283);
or U2707 (N_2707,N_2081,N_2375);
nand U2708 (N_2708,N_2418,N_2242);
and U2709 (N_2709,N_2361,N_2351);
nand U2710 (N_2710,N_2498,N_2399);
nor U2711 (N_2711,N_2049,N_2289);
nand U2712 (N_2712,N_2039,N_2374);
nor U2713 (N_2713,N_2318,N_2103);
nor U2714 (N_2714,N_2461,N_2215);
xnor U2715 (N_2715,N_2365,N_2021);
nor U2716 (N_2716,N_2004,N_2245);
and U2717 (N_2717,N_2130,N_2239);
nor U2718 (N_2718,N_2462,N_2191);
nor U2719 (N_2719,N_2227,N_2328);
nor U2720 (N_2720,N_2196,N_2050);
nand U2721 (N_2721,N_2148,N_2173);
or U2722 (N_2722,N_2417,N_2197);
and U2723 (N_2723,N_2433,N_2306);
or U2724 (N_2724,N_2426,N_2266);
nor U2725 (N_2725,N_2158,N_2124);
and U2726 (N_2726,N_2246,N_2254);
and U2727 (N_2727,N_2041,N_2133);
nor U2728 (N_2728,N_2333,N_2243);
xnor U2729 (N_2729,N_2094,N_2269);
nor U2730 (N_2730,N_2489,N_2356);
nand U2731 (N_2731,N_2230,N_2051);
nor U2732 (N_2732,N_2235,N_2126);
nor U2733 (N_2733,N_2030,N_2366);
or U2734 (N_2734,N_2310,N_2154);
and U2735 (N_2735,N_2272,N_2065);
nand U2736 (N_2736,N_2219,N_2240);
nand U2737 (N_2737,N_2203,N_2027);
nand U2738 (N_2738,N_2359,N_2182);
nor U2739 (N_2739,N_2229,N_2026);
and U2740 (N_2740,N_2075,N_2497);
or U2741 (N_2741,N_2183,N_2309);
and U2742 (N_2742,N_2111,N_2400);
nor U2743 (N_2743,N_2477,N_2064);
and U2744 (N_2744,N_2224,N_2007);
nor U2745 (N_2745,N_2295,N_2226);
nand U2746 (N_2746,N_2279,N_2125);
nor U2747 (N_2747,N_2074,N_2035);
or U2748 (N_2748,N_2317,N_2129);
and U2749 (N_2749,N_2376,N_2484);
nor U2750 (N_2750,N_2052,N_2403);
and U2751 (N_2751,N_2401,N_2012);
and U2752 (N_2752,N_2386,N_2343);
or U2753 (N_2753,N_2306,N_2481);
and U2754 (N_2754,N_2279,N_2094);
nor U2755 (N_2755,N_2097,N_2039);
and U2756 (N_2756,N_2042,N_2178);
nand U2757 (N_2757,N_2480,N_2343);
or U2758 (N_2758,N_2097,N_2428);
xor U2759 (N_2759,N_2221,N_2082);
and U2760 (N_2760,N_2149,N_2446);
nor U2761 (N_2761,N_2135,N_2164);
nand U2762 (N_2762,N_2041,N_2141);
and U2763 (N_2763,N_2071,N_2469);
nor U2764 (N_2764,N_2441,N_2407);
nand U2765 (N_2765,N_2419,N_2287);
nand U2766 (N_2766,N_2160,N_2277);
nor U2767 (N_2767,N_2481,N_2496);
or U2768 (N_2768,N_2400,N_2489);
nand U2769 (N_2769,N_2179,N_2217);
and U2770 (N_2770,N_2039,N_2321);
or U2771 (N_2771,N_2028,N_2060);
or U2772 (N_2772,N_2382,N_2220);
nand U2773 (N_2773,N_2074,N_2107);
nand U2774 (N_2774,N_2030,N_2181);
nand U2775 (N_2775,N_2322,N_2014);
nand U2776 (N_2776,N_2280,N_2304);
or U2777 (N_2777,N_2458,N_2489);
nand U2778 (N_2778,N_2074,N_2304);
and U2779 (N_2779,N_2293,N_2381);
nand U2780 (N_2780,N_2412,N_2117);
or U2781 (N_2781,N_2102,N_2479);
and U2782 (N_2782,N_2446,N_2078);
nand U2783 (N_2783,N_2403,N_2431);
nor U2784 (N_2784,N_2354,N_2489);
and U2785 (N_2785,N_2340,N_2204);
nand U2786 (N_2786,N_2441,N_2290);
nor U2787 (N_2787,N_2262,N_2309);
or U2788 (N_2788,N_2309,N_2450);
xnor U2789 (N_2789,N_2042,N_2291);
or U2790 (N_2790,N_2168,N_2313);
and U2791 (N_2791,N_2185,N_2457);
or U2792 (N_2792,N_2049,N_2026);
and U2793 (N_2793,N_2026,N_2286);
and U2794 (N_2794,N_2038,N_2160);
and U2795 (N_2795,N_2060,N_2027);
and U2796 (N_2796,N_2323,N_2363);
or U2797 (N_2797,N_2422,N_2035);
and U2798 (N_2798,N_2014,N_2240);
and U2799 (N_2799,N_2468,N_2476);
and U2800 (N_2800,N_2173,N_2188);
or U2801 (N_2801,N_2394,N_2216);
and U2802 (N_2802,N_2037,N_2006);
and U2803 (N_2803,N_2429,N_2202);
and U2804 (N_2804,N_2123,N_2214);
nand U2805 (N_2805,N_2107,N_2196);
nor U2806 (N_2806,N_2087,N_2398);
or U2807 (N_2807,N_2494,N_2369);
nand U2808 (N_2808,N_2498,N_2343);
or U2809 (N_2809,N_2001,N_2249);
nor U2810 (N_2810,N_2033,N_2076);
nand U2811 (N_2811,N_2401,N_2056);
and U2812 (N_2812,N_2450,N_2364);
or U2813 (N_2813,N_2328,N_2437);
nand U2814 (N_2814,N_2345,N_2026);
and U2815 (N_2815,N_2399,N_2187);
nand U2816 (N_2816,N_2275,N_2413);
and U2817 (N_2817,N_2335,N_2481);
nand U2818 (N_2818,N_2452,N_2193);
nand U2819 (N_2819,N_2114,N_2496);
nand U2820 (N_2820,N_2367,N_2399);
nor U2821 (N_2821,N_2328,N_2082);
nor U2822 (N_2822,N_2479,N_2204);
nand U2823 (N_2823,N_2377,N_2044);
nor U2824 (N_2824,N_2370,N_2463);
and U2825 (N_2825,N_2360,N_2461);
nand U2826 (N_2826,N_2206,N_2485);
and U2827 (N_2827,N_2398,N_2077);
nor U2828 (N_2828,N_2076,N_2287);
or U2829 (N_2829,N_2303,N_2110);
or U2830 (N_2830,N_2122,N_2026);
and U2831 (N_2831,N_2493,N_2384);
nand U2832 (N_2832,N_2290,N_2025);
nor U2833 (N_2833,N_2060,N_2321);
nand U2834 (N_2834,N_2292,N_2223);
nand U2835 (N_2835,N_2472,N_2156);
nor U2836 (N_2836,N_2451,N_2266);
and U2837 (N_2837,N_2423,N_2241);
or U2838 (N_2838,N_2012,N_2094);
nand U2839 (N_2839,N_2298,N_2476);
and U2840 (N_2840,N_2229,N_2188);
nand U2841 (N_2841,N_2118,N_2034);
nor U2842 (N_2842,N_2052,N_2488);
nor U2843 (N_2843,N_2077,N_2440);
nand U2844 (N_2844,N_2235,N_2445);
nor U2845 (N_2845,N_2420,N_2445);
nand U2846 (N_2846,N_2187,N_2492);
nand U2847 (N_2847,N_2314,N_2135);
or U2848 (N_2848,N_2217,N_2168);
nor U2849 (N_2849,N_2110,N_2300);
nor U2850 (N_2850,N_2244,N_2432);
and U2851 (N_2851,N_2450,N_2384);
nor U2852 (N_2852,N_2292,N_2231);
nand U2853 (N_2853,N_2130,N_2006);
nor U2854 (N_2854,N_2334,N_2428);
nor U2855 (N_2855,N_2218,N_2443);
and U2856 (N_2856,N_2494,N_2021);
and U2857 (N_2857,N_2119,N_2125);
nand U2858 (N_2858,N_2094,N_2181);
xnor U2859 (N_2859,N_2465,N_2316);
or U2860 (N_2860,N_2441,N_2220);
or U2861 (N_2861,N_2252,N_2499);
nor U2862 (N_2862,N_2025,N_2029);
and U2863 (N_2863,N_2416,N_2348);
nor U2864 (N_2864,N_2448,N_2407);
or U2865 (N_2865,N_2039,N_2208);
and U2866 (N_2866,N_2330,N_2176);
xnor U2867 (N_2867,N_2259,N_2247);
nor U2868 (N_2868,N_2356,N_2272);
and U2869 (N_2869,N_2451,N_2173);
nor U2870 (N_2870,N_2375,N_2440);
nand U2871 (N_2871,N_2197,N_2201);
nor U2872 (N_2872,N_2255,N_2494);
or U2873 (N_2873,N_2112,N_2079);
xnor U2874 (N_2874,N_2264,N_2427);
nor U2875 (N_2875,N_2124,N_2252);
or U2876 (N_2876,N_2243,N_2108);
nor U2877 (N_2877,N_2348,N_2264);
nand U2878 (N_2878,N_2068,N_2434);
or U2879 (N_2879,N_2474,N_2148);
nand U2880 (N_2880,N_2498,N_2006);
nor U2881 (N_2881,N_2140,N_2405);
nor U2882 (N_2882,N_2196,N_2416);
nor U2883 (N_2883,N_2217,N_2285);
nand U2884 (N_2884,N_2482,N_2243);
or U2885 (N_2885,N_2335,N_2364);
or U2886 (N_2886,N_2464,N_2241);
nand U2887 (N_2887,N_2419,N_2264);
xor U2888 (N_2888,N_2290,N_2376);
nor U2889 (N_2889,N_2092,N_2346);
nor U2890 (N_2890,N_2421,N_2006);
nand U2891 (N_2891,N_2358,N_2130);
and U2892 (N_2892,N_2273,N_2272);
or U2893 (N_2893,N_2324,N_2171);
and U2894 (N_2894,N_2220,N_2476);
or U2895 (N_2895,N_2278,N_2331);
xnor U2896 (N_2896,N_2009,N_2311);
nand U2897 (N_2897,N_2071,N_2058);
xor U2898 (N_2898,N_2213,N_2305);
nor U2899 (N_2899,N_2153,N_2164);
or U2900 (N_2900,N_2037,N_2066);
nor U2901 (N_2901,N_2276,N_2161);
nand U2902 (N_2902,N_2405,N_2257);
nor U2903 (N_2903,N_2028,N_2131);
nor U2904 (N_2904,N_2434,N_2162);
or U2905 (N_2905,N_2071,N_2214);
nand U2906 (N_2906,N_2332,N_2334);
nand U2907 (N_2907,N_2105,N_2469);
and U2908 (N_2908,N_2029,N_2322);
and U2909 (N_2909,N_2313,N_2488);
or U2910 (N_2910,N_2315,N_2260);
nand U2911 (N_2911,N_2359,N_2303);
nor U2912 (N_2912,N_2285,N_2311);
nand U2913 (N_2913,N_2116,N_2413);
or U2914 (N_2914,N_2259,N_2173);
or U2915 (N_2915,N_2252,N_2185);
and U2916 (N_2916,N_2179,N_2195);
nand U2917 (N_2917,N_2134,N_2327);
nand U2918 (N_2918,N_2351,N_2476);
nand U2919 (N_2919,N_2118,N_2361);
nor U2920 (N_2920,N_2328,N_2135);
or U2921 (N_2921,N_2349,N_2399);
nand U2922 (N_2922,N_2431,N_2051);
nand U2923 (N_2923,N_2346,N_2452);
nand U2924 (N_2924,N_2234,N_2177);
nor U2925 (N_2925,N_2137,N_2175);
and U2926 (N_2926,N_2093,N_2362);
or U2927 (N_2927,N_2320,N_2081);
nand U2928 (N_2928,N_2169,N_2442);
or U2929 (N_2929,N_2266,N_2411);
and U2930 (N_2930,N_2106,N_2004);
xnor U2931 (N_2931,N_2210,N_2398);
nor U2932 (N_2932,N_2336,N_2483);
or U2933 (N_2933,N_2460,N_2030);
or U2934 (N_2934,N_2195,N_2218);
nor U2935 (N_2935,N_2225,N_2036);
nor U2936 (N_2936,N_2480,N_2180);
nor U2937 (N_2937,N_2272,N_2484);
nand U2938 (N_2938,N_2483,N_2062);
or U2939 (N_2939,N_2206,N_2024);
nor U2940 (N_2940,N_2158,N_2349);
nor U2941 (N_2941,N_2011,N_2380);
or U2942 (N_2942,N_2224,N_2262);
nand U2943 (N_2943,N_2061,N_2187);
or U2944 (N_2944,N_2333,N_2198);
nor U2945 (N_2945,N_2260,N_2365);
and U2946 (N_2946,N_2303,N_2466);
and U2947 (N_2947,N_2308,N_2031);
and U2948 (N_2948,N_2444,N_2180);
xnor U2949 (N_2949,N_2443,N_2003);
nor U2950 (N_2950,N_2153,N_2357);
nand U2951 (N_2951,N_2285,N_2492);
nand U2952 (N_2952,N_2323,N_2391);
nand U2953 (N_2953,N_2114,N_2273);
and U2954 (N_2954,N_2445,N_2215);
nor U2955 (N_2955,N_2187,N_2302);
nand U2956 (N_2956,N_2247,N_2253);
nor U2957 (N_2957,N_2436,N_2429);
xnor U2958 (N_2958,N_2480,N_2329);
and U2959 (N_2959,N_2355,N_2176);
or U2960 (N_2960,N_2133,N_2030);
nand U2961 (N_2961,N_2310,N_2372);
nand U2962 (N_2962,N_2131,N_2219);
or U2963 (N_2963,N_2161,N_2152);
xor U2964 (N_2964,N_2031,N_2483);
and U2965 (N_2965,N_2335,N_2198);
nand U2966 (N_2966,N_2426,N_2290);
and U2967 (N_2967,N_2332,N_2292);
or U2968 (N_2968,N_2376,N_2466);
nand U2969 (N_2969,N_2139,N_2418);
nor U2970 (N_2970,N_2480,N_2133);
or U2971 (N_2971,N_2041,N_2323);
and U2972 (N_2972,N_2121,N_2048);
and U2973 (N_2973,N_2367,N_2065);
xnor U2974 (N_2974,N_2014,N_2201);
and U2975 (N_2975,N_2116,N_2429);
nand U2976 (N_2976,N_2337,N_2335);
and U2977 (N_2977,N_2323,N_2249);
or U2978 (N_2978,N_2400,N_2241);
and U2979 (N_2979,N_2155,N_2153);
nor U2980 (N_2980,N_2291,N_2153);
nand U2981 (N_2981,N_2459,N_2275);
or U2982 (N_2982,N_2238,N_2173);
or U2983 (N_2983,N_2494,N_2009);
nor U2984 (N_2984,N_2481,N_2145);
and U2985 (N_2985,N_2355,N_2008);
or U2986 (N_2986,N_2079,N_2084);
or U2987 (N_2987,N_2199,N_2458);
nand U2988 (N_2988,N_2061,N_2001);
nor U2989 (N_2989,N_2026,N_2401);
or U2990 (N_2990,N_2098,N_2497);
nand U2991 (N_2991,N_2397,N_2330);
nand U2992 (N_2992,N_2293,N_2323);
or U2993 (N_2993,N_2306,N_2000);
nand U2994 (N_2994,N_2223,N_2204);
nand U2995 (N_2995,N_2451,N_2319);
or U2996 (N_2996,N_2190,N_2016);
nor U2997 (N_2997,N_2279,N_2259);
and U2998 (N_2998,N_2401,N_2429);
nor U2999 (N_2999,N_2404,N_2311);
or U3000 (N_3000,N_2864,N_2934);
xnor U3001 (N_3001,N_2641,N_2959);
or U3002 (N_3002,N_2653,N_2504);
and U3003 (N_3003,N_2648,N_2767);
nor U3004 (N_3004,N_2503,N_2736);
nor U3005 (N_3005,N_2585,N_2887);
nor U3006 (N_3006,N_2670,N_2536);
nor U3007 (N_3007,N_2576,N_2924);
nor U3008 (N_3008,N_2973,N_2785);
and U3009 (N_3009,N_2899,N_2601);
nand U3010 (N_3010,N_2805,N_2710);
and U3011 (N_3011,N_2730,N_2573);
nand U3012 (N_3012,N_2796,N_2662);
or U3013 (N_3013,N_2669,N_2609);
or U3014 (N_3014,N_2949,N_2633);
nand U3015 (N_3015,N_2786,N_2904);
nand U3016 (N_3016,N_2510,N_2920);
nor U3017 (N_3017,N_2562,N_2844);
nand U3018 (N_3018,N_2945,N_2881);
nor U3019 (N_3019,N_2741,N_2671);
nor U3020 (N_3020,N_2718,N_2518);
and U3021 (N_3021,N_2908,N_2657);
nor U3022 (N_3022,N_2880,N_2624);
or U3023 (N_3023,N_2995,N_2651);
nand U3024 (N_3024,N_2631,N_2513);
and U3025 (N_3025,N_2758,N_2909);
nand U3026 (N_3026,N_2658,N_2993);
and U3027 (N_3027,N_2647,N_2808);
or U3028 (N_3028,N_2673,N_2519);
and U3029 (N_3029,N_2614,N_2849);
nor U3030 (N_3030,N_2680,N_2531);
nor U3031 (N_3031,N_2582,N_2878);
nand U3032 (N_3032,N_2528,N_2763);
nand U3033 (N_3033,N_2687,N_2543);
or U3034 (N_3034,N_2867,N_2622);
nor U3035 (N_3035,N_2912,N_2726);
nand U3036 (N_3036,N_2996,N_2630);
nand U3037 (N_3037,N_2723,N_2728);
or U3038 (N_3038,N_2558,N_2884);
and U3039 (N_3039,N_2509,N_2744);
or U3040 (N_3040,N_2516,N_2906);
nand U3041 (N_3041,N_2532,N_2937);
nand U3042 (N_3042,N_2674,N_2533);
and U3043 (N_3043,N_2889,N_2848);
or U3044 (N_3044,N_2646,N_2733);
nor U3045 (N_3045,N_2713,N_2637);
or U3046 (N_3046,N_2656,N_2965);
nand U3047 (N_3047,N_2623,N_2618);
nand U3048 (N_3048,N_2501,N_2709);
and U3049 (N_3049,N_2832,N_2526);
and U3050 (N_3050,N_2850,N_2695);
or U3051 (N_3051,N_2791,N_2911);
and U3052 (N_3052,N_2705,N_2659);
nor U3053 (N_3053,N_2749,N_2682);
and U3054 (N_3054,N_2634,N_2777);
nor U3055 (N_3055,N_2795,N_2968);
nand U3056 (N_3056,N_2925,N_2552);
nand U3057 (N_3057,N_2701,N_2628);
or U3058 (N_3058,N_2661,N_2708);
or U3059 (N_3059,N_2928,N_2553);
or U3060 (N_3060,N_2690,N_2769);
nor U3061 (N_3061,N_2551,N_2566);
nor U3062 (N_3062,N_2824,N_2907);
or U3063 (N_3063,N_2716,N_2650);
or U3064 (N_3064,N_2955,N_2745);
nand U3065 (N_3065,N_2780,N_2626);
or U3066 (N_3066,N_2982,N_2948);
and U3067 (N_3067,N_2714,N_2883);
and U3068 (N_3068,N_2966,N_2765);
nor U3069 (N_3069,N_2704,N_2766);
or U3070 (N_3070,N_2933,N_2644);
and U3071 (N_3071,N_2679,N_2688);
and U3072 (N_3072,N_2967,N_2860);
and U3073 (N_3073,N_2514,N_2592);
nor U3074 (N_3074,N_2869,N_2865);
and U3075 (N_3075,N_2971,N_2613);
and U3076 (N_3076,N_2581,N_2580);
nor U3077 (N_3077,N_2876,N_2746);
nand U3078 (N_3078,N_2610,N_2579);
and U3079 (N_3079,N_2508,N_2843);
or U3080 (N_3080,N_2840,N_2607);
and U3081 (N_3081,N_2681,N_2892);
or U3082 (N_3082,N_2923,N_2793);
nor U3083 (N_3083,N_2890,N_2706);
or U3084 (N_3084,N_2675,N_2962);
or U3085 (N_3085,N_2771,N_2655);
or U3086 (N_3086,N_2814,N_2806);
or U3087 (N_3087,N_2594,N_2555);
nand U3088 (N_3088,N_2753,N_2632);
or U3089 (N_3089,N_2699,N_2783);
xor U3090 (N_3090,N_2983,N_2807);
or U3091 (N_3091,N_2667,N_2590);
or U3092 (N_3092,N_2755,N_2523);
and U3093 (N_3093,N_2963,N_2550);
nor U3094 (N_3094,N_2625,N_2642);
or U3095 (N_3095,N_2980,N_2604);
nand U3096 (N_3096,N_2936,N_2639);
nor U3097 (N_3097,N_2717,N_2740);
and U3098 (N_3098,N_2927,N_2542);
and U3099 (N_3099,N_2943,N_2559);
nor U3100 (N_3100,N_2729,N_2764);
or U3101 (N_3101,N_2839,N_2831);
and U3102 (N_3102,N_2629,N_2683);
or U3103 (N_3103,N_2539,N_2752);
nand U3104 (N_3104,N_2697,N_2739);
and U3105 (N_3105,N_2847,N_2627);
nor U3106 (N_3106,N_2931,N_2851);
nand U3107 (N_3107,N_2801,N_2544);
and U3108 (N_3108,N_2569,N_2506);
or U3109 (N_3109,N_2578,N_2762);
or U3110 (N_3110,N_2507,N_2898);
or U3111 (N_3111,N_2868,N_2685);
and U3112 (N_3112,N_2882,N_2602);
and U3113 (N_3113,N_2571,N_2872);
and U3114 (N_3114,N_2502,N_2692);
xnor U3115 (N_3115,N_2998,N_2874);
xnor U3116 (N_3116,N_2854,N_2938);
nor U3117 (N_3117,N_2829,N_2951);
or U3118 (N_3118,N_2790,N_2921);
nand U3119 (N_3119,N_2960,N_2702);
nor U3120 (N_3120,N_2525,N_2902);
nor U3121 (N_3121,N_2852,N_2735);
or U3122 (N_3122,N_2577,N_2810);
nand U3123 (N_3123,N_2556,N_2813);
nand U3124 (N_3124,N_2608,N_2800);
and U3125 (N_3125,N_2879,N_2694);
nand U3126 (N_3126,N_2922,N_2989);
or U3127 (N_3127,N_2640,N_2893);
and U3128 (N_3128,N_2593,N_2835);
nand U3129 (N_3129,N_2522,N_2530);
and U3130 (N_3130,N_2597,N_2564);
or U3131 (N_3131,N_2886,N_2970);
nand U3132 (N_3132,N_2822,N_2885);
nor U3133 (N_3133,N_2621,N_2969);
or U3134 (N_3134,N_2759,N_2595);
nand U3135 (N_3135,N_2720,N_2816);
nor U3136 (N_3136,N_2798,N_2981);
nor U3137 (N_3137,N_2956,N_2787);
nand U3138 (N_3138,N_2821,N_2802);
nor U3139 (N_3139,N_2722,N_2616);
and U3140 (N_3140,N_2599,N_2684);
nor U3141 (N_3141,N_2914,N_2567);
nor U3142 (N_3142,N_2678,N_2823);
nand U3143 (N_3143,N_2529,N_2845);
and U3144 (N_3144,N_2779,N_2561);
or U3145 (N_3145,N_2775,N_2589);
and U3146 (N_3146,N_2985,N_2547);
nand U3147 (N_3147,N_2660,N_2797);
nand U3148 (N_3148,N_2570,N_2990);
or U3149 (N_3149,N_2819,N_2903);
and U3150 (N_3150,N_2603,N_2900);
nor U3151 (N_3151,N_2774,N_2841);
or U3152 (N_3152,N_2871,N_2859);
or U3153 (N_3153,N_2804,N_2707);
nand U3154 (N_3154,N_2789,N_2500);
nand U3155 (N_3155,N_2999,N_2505);
nand U3156 (N_3156,N_2545,N_2615);
and U3157 (N_3157,N_2930,N_2935);
or U3158 (N_3158,N_2842,N_2803);
nor U3159 (N_3159,N_2792,N_2815);
and U3160 (N_3160,N_2870,N_2919);
nor U3161 (N_3161,N_2711,N_2664);
or U3162 (N_3162,N_2611,N_2916);
or U3163 (N_3163,N_2944,N_2760);
nor U3164 (N_3164,N_2747,N_2668);
nand U3165 (N_3165,N_2897,N_2932);
and U3166 (N_3166,N_2591,N_2712);
and U3167 (N_3167,N_2541,N_2940);
nand U3168 (N_3168,N_2612,N_2548);
nor U3169 (N_3169,N_2988,N_2677);
nand U3170 (N_3170,N_2979,N_2583);
nor U3171 (N_3171,N_2619,N_2950);
or U3172 (N_3172,N_2992,N_2748);
nand U3173 (N_3173,N_2858,N_2877);
and U3174 (N_3174,N_2820,N_2875);
or U3175 (N_3175,N_2857,N_2895);
nor U3176 (N_3176,N_2987,N_2794);
nor U3177 (N_3177,N_2836,N_2588);
or U3178 (N_3178,N_2978,N_2521);
and U3179 (N_3179,N_2957,N_2584);
nor U3180 (N_3180,N_2773,N_2863);
nor U3181 (N_3181,N_2649,N_2698);
or U3182 (N_3182,N_2511,N_2838);
or U3183 (N_3183,N_2861,N_2654);
nand U3184 (N_3184,N_2587,N_2663);
nor U3185 (N_3185,N_2535,N_2941);
nand U3186 (N_3186,N_2974,N_2913);
and U3187 (N_3187,N_2942,N_2905);
or U3188 (N_3188,N_2926,N_2703);
or U3189 (N_3189,N_2776,N_2693);
xnor U3190 (N_3190,N_2984,N_2738);
nand U3191 (N_3191,N_2947,N_2575);
or U3192 (N_3192,N_2751,N_2818);
or U3193 (N_3193,N_2652,N_2524);
nor U3194 (N_3194,N_2617,N_2954);
and U3195 (N_3195,N_2598,N_2826);
or U3196 (N_3196,N_2828,N_2896);
and U3197 (N_3197,N_2565,N_2606);
nor U3198 (N_3198,N_2901,N_2772);
nand U3199 (N_3199,N_2554,N_2605);
and U3200 (N_3200,N_2915,N_2645);
nand U3201 (N_3201,N_2853,N_2817);
or U3202 (N_3202,N_2515,N_2986);
nor U3203 (N_3203,N_2991,N_2727);
and U3204 (N_3204,N_2620,N_2834);
nor U3205 (N_3205,N_2563,N_2856);
or U3206 (N_3206,N_2972,N_2691);
nand U3207 (N_3207,N_2696,N_2918);
or U3208 (N_3208,N_2600,N_2574);
or U3209 (N_3209,N_2976,N_2846);
and U3210 (N_3210,N_2686,N_2952);
and U3211 (N_3211,N_2743,N_2731);
nor U3212 (N_3212,N_2724,N_2862);
nor U3213 (N_3213,N_2873,N_2737);
nand U3214 (N_3214,N_2666,N_2557);
nand U3215 (N_3215,N_2977,N_2754);
nor U3216 (N_3216,N_2888,N_2596);
nor U3217 (N_3217,N_2781,N_2586);
nand U3218 (N_3218,N_2961,N_2917);
and U3219 (N_3219,N_2742,N_2546);
nand U3220 (N_3220,N_2891,N_2830);
and U3221 (N_3221,N_2512,N_2721);
or U3222 (N_3222,N_2534,N_2549);
and U3223 (N_3223,N_2540,N_2750);
nand U3224 (N_3224,N_2827,N_2572);
nand U3225 (N_3225,N_2756,N_2538);
or U3226 (N_3226,N_2812,N_2719);
and U3227 (N_3227,N_2958,N_2568);
nand U3228 (N_3228,N_2809,N_2725);
and U3229 (N_3229,N_2689,N_2527);
nand U3230 (N_3230,N_2964,N_2757);
or U3231 (N_3231,N_2975,N_2939);
or U3232 (N_3232,N_2784,N_2782);
xor U3233 (N_3233,N_2946,N_2833);
or U3234 (N_3234,N_2811,N_2894);
or U3235 (N_3235,N_2732,N_2761);
nand U3236 (N_3236,N_2537,N_2929);
nand U3237 (N_3237,N_2700,N_2676);
xor U3238 (N_3238,N_2643,N_2768);
xnor U3239 (N_3239,N_2825,N_2778);
nand U3240 (N_3240,N_2638,N_2517);
or U3241 (N_3241,N_2560,N_2734);
nand U3242 (N_3242,N_2953,N_2770);
and U3243 (N_3243,N_2635,N_2866);
xor U3244 (N_3244,N_2665,N_2636);
and U3245 (N_3245,N_2837,N_2715);
nor U3246 (N_3246,N_2520,N_2910);
nand U3247 (N_3247,N_2855,N_2997);
nand U3248 (N_3248,N_2799,N_2788);
xnor U3249 (N_3249,N_2672,N_2994);
nor U3250 (N_3250,N_2782,N_2968);
or U3251 (N_3251,N_2964,N_2642);
nor U3252 (N_3252,N_2654,N_2721);
nor U3253 (N_3253,N_2853,N_2653);
and U3254 (N_3254,N_2604,N_2795);
nand U3255 (N_3255,N_2511,N_2900);
nand U3256 (N_3256,N_2706,N_2545);
and U3257 (N_3257,N_2685,N_2899);
nor U3258 (N_3258,N_2971,N_2727);
or U3259 (N_3259,N_2675,N_2669);
or U3260 (N_3260,N_2652,N_2948);
or U3261 (N_3261,N_2580,N_2958);
or U3262 (N_3262,N_2577,N_2731);
or U3263 (N_3263,N_2826,N_2653);
xnor U3264 (N_3264,N_2583,N_2713);
or U3265 (N_3265,N_2892,N_2856);
nor U3266 (N_3266,N_2655,N_2739);
and U3267 (N_3267,N_2663,N_2577);
and U3268 (N_3268,N_2566,N_2897);
and U3269 (N_3269,N_2741,N_2912);
nand U3270 (N_3270,N_2725,N_2585);
nand U3271 (N_3271,N_2564,N_2873);
xnor U3272 (N_3272,N_2775,N_2933);
nand U3273 (N_3273,N_2537,N_2945);
or U3274 (N_3274,N_2905,N_2772);
nor U3275 (N_3275,N_2857,N_2901);
nor U3276 (N_3276,N_2973,N_2609);
or U3277 (N_3277,N_2719,N_2950);
xor U3278 (N_3278,N_2720,N_2941);
nor U3279 (N_3279,N_2775,N_2683);
nand U3280 (N_3280,N_2840,N_2900);
or U3281 (N_3281,N_2915,N_2912);
or U3282 (N_3282,N_2597,N_2957);
or U3283 (N_3283,N_2505,N_2767);
nand U3284 (N_3284,N_2598,N_2715);
or U3285 (N_3285,N_2603,N_2651);
nand U3286 (N_3286,N_2747,N_2768);
or U3287 (N_3287,N_2863,N_2874);
or U3288 (N_3288,N_2509,N_2736);
nand U3289 (N_3289,N_2670,N_2596);
and U3290 (N_3290,N_2602,N_2741);
or U3291 (N_3291,N_2676,N_2770);
and U3292 (N_3292,N_2964,N_2649);
or U3293 (N_3293,N_2779,N_2786);
and U3294 (N_3294,N_2762,N_2902);
nand U3295 (N_3295,N_2813,N_2830);
or U3296 (N_3296,N_2905,N_2906);
and U3297 (N_3297,N_2626,N_2832);
nand U3298 (N_3298,N_2869,N_2947);
and U3299 (N_3299,N_2750,N_2559);
nor U3300 (N_3300,N_2763,N_2523);
nand U3301 (N_3301,N_2626,N_2731);
and U3302 (N_3302,N_2752,N_2895);
xor U3303 (N_3303,N_2698,N_2877);
nor U3304 (N_3304,N_2688,N_2743);
nor U3305 (N_3305,N_2621,N_2882);
nor U3306 (N_3306,N_2940,N_2578);
and U3307 (N_3307,N_2879,N_2507);
xnor U3308 (N_3308,N_2885,N_2922);
and U3309 (N_3309,N_2512,N_2985);
and U3310 (N_3310,N_2897,N_2780);
nand U3311 (N_3311,N_2786,N_2575);
or U3312 (N_3312,N_2643,N_2739);
nand U3313 (N_3313,N_2979,N_2996);
nand U3314 (N_3314,N_2552,N_2701);
nand U3315 (N_3315,N_2707,N_2732);
nand U3316 (N_3316,N_2575,N_2814);
and U3317 (N_3317,N_2973,N_2682);
or U3318 (N_3318,N_2733,N_2589);
or U3319 (N_3319,N_2797,N_2778);
nand U3320 (N_3320,N_2604,N_2780);
or U3321 (N_3321,N_2575,N_2861);
or U3322 (N_3322,N_2570,N_2739);
or U3323 (N_3323,N_2675,N_2926);
and U3324 (N_3324,N_2891,N_2671);
or U3325 (N_3325,N_2596,N_2727);
nor U3326 (N_3326,N_2929,N_2868);
nor U3327 (N_3327,N_2672,N_2870);
nand U3328 (N_3328,N_2807,N_2948);
or U3329 (N_3329,N_2746,N_2883);
nor U3330 (N_3330,N_2580,N_2833);
or U3331 (N_3331,N_2859,N_2704);
or U3332 (N_3332,N_2977,N_2747);
or U3333 (N_3333,N_2854,N_2972);
or U3334 (N_3334,N_2885,N_2817);
and U3335 (N_3335,N_2597,N_2817);
or U3336 (N_3336,N_2851,N_2793);
nand U3337 (N_3337,N_2989,N_2589);
nor U3338 (N_3338,N_2772,N_2532);
nand U3339 (N_3339,N_2555,N_2900);
and U3340 (N_3340,N_2820,N_2631);
nand U3341 (N_3341,N_2597,N_2890);
nor U3342 (N_3342,N_2963,N_2744);
and U3343 (N_3343,N_2708,N_2954);
nand U3344 (N_3344,N_2719,N_2620);
and U3345 (N_3345,N_2785,N_2682);
or U3346 (N_3346,N_2677,N_2747);
or U3347 (N_3347,N_2581,N_2706);
nand U3348 (N_3348,N_2503,N_2942);
nor U3349 (N_3349,N_2582,N_2817);
or U3350 (N_3350,N_2890,N_2609);
or U3351 (N_3351,N_2541,N_2725);
or U3352 (N_3352,N_2938,N_2572);
nor U3353 (N_3353,N_2881,N_2645);
xnor U3354 (N_3354,N_2585,N_2519);
and U3355 (N_3355,N_2596,N_2634);
nand U3356 (N_3356,N_2807,N_2785);
nand U3357 (N_3357,N_2662,N_2574);
nand U3358 (N_3358,N_2794,N_2951);
or U3359 (N_3359,N_2663,N_2817);
or U3360 (N_3360,N_2629,N_2778);
or U3361 (N_3361,N_2698,N_2662);
or U3362 (N_3362,N_2659,N_2986);
nand U3363 (N_3363,N_2906,N_2607);
nand U3364 (N_3364,N_2959,N_2820);
and U3365 (N_3365,N_2609,N_2521);
and U3366 (N_3366,N_2789,N_2823);
nor U3367 (N_3367,N_2997,N_2610);
nand U3368 (N_3368,N_2578,N_2693);
and U3369 (N_3369,N_2934,N_2818);
nor U3370 (N_3370,N_2626,N_2985);
and U3371 (N_3371,N_2702,N_2577);
and U3372 (N_3372,N_2959,N_2586);
and U3373 (N_3373,N_2664,N_2972);
nor U3374 (N_3374,N_2968,N_2984);
xnor U3375 (N_3375,N_2973,N_2663);
nand U3376 (N_3376,N_2649,N_2501);
nor U3377 (N_3377,N_2713,N_2963);
nand U3378 (N_3378,N_2744,N_2969);
nand U3379 (N_3379,N_2756,N_2517);
nand U3380 (N_3380,N_2900,N_2934);
nand U3381 (N_3381,N_2558,N_2556);
nor U3382 (N_3382,N_2621,N_2805);
or U3383 (N_3383,N_2816,N_2652);
or U3384 (N_3384,N_2648,N_2932);
or U3385 (N_3385,N_2513,N_2596);
nand U3386 (N_3386,N_2505,N_2690);
nor U3387 (N_3387,N_2548,N_2918);
nand U3388 (N_3388,N_2827,N_2634);
nor U3389 (N_3389,N_2620,N_2614);
nand U3390 (N_3390,N_2759,N_2827);
and U3391 (N_3391,N_2811,N_2985);
xnor U3392 (N_3392,N_2903,N_2667);
xnor U3393 (N_3393,N_2589,N_2962);
nand U3394 (N_3394,N_2862,N_2546);
nor U3395 (N_3395,N_2991,N_2678);
nor U3396 (N_3396,N_2870,N_2770);
nor U3397 (N_3397,N_2981,N_2622);
nand U3398 (N_3398,N_2839,N_2827);
nand U3399 (N_3399,N_2961,N_2614);
nand U3400 (N_3400,N_2542,N_2723);
and U3401 (N_3401,N_2680,N_2822);
nand U3402 (N_3402,N_2694,N_2691);
and U3403 (N_3403,N_2628,N_2960);
nand U3404 (N_3404,N_2798,N_2754);
nor U3405 (N_3405,N_2864,N_2900);
nand U3406 (N_3406,N_2657,N_2910);
nor U3407 (N_3407,N_2847,N_2791);
nor U3408 (N_3408,N_2965,N_2874);
and U3409 (N_3409,N_2508,N_2624);
nand U3410 (N_3410,N_2885,N_2567);
nor U3411 (N_3411,N_2598,N_2845);
nand U3412 (N_3412,N_2601,N_2998);
nand U3413 (N_3413,N_2991,N_2721);
or U3414 (N_3414,N_2835,N_2540);
nor U3415 (N_3415,N_2613,N_2962);
nor U3416 (N_3416,N_2613,N_2632);
nor U3417 (N_3417,N_2731,N_2859);
nand U3418 (N_3418,N_2515,N_2517);
and U3419 (N_3419,N_2755,N_2719);
and U3420 (N_3420,N_2869,N_2797);
nor U3421 (N_3421,N_2925,N_2673);
nand U3422 (N_3422,N_2790,N_2869);
nor U3423 (N_3423,N_2595,N_2709);
or U3424 (N_3424,N_2909,N_2713);
and U3425 (N_3425,N_2621,N_2586);
or U3426 (N_3426,N_2671,N_2629);
or U3427 (N_3427,N_2574,N_2809);
nor U3428 (N_3428,N_2660,N_2698);
and U3429 (N_3429,N_2550,N_2789);
nand U3430 (N_3430,N_2784,N_2660);
nand U3431 (N_3431,N_2526,N_2922);
nand U3432 (N_3432,N_2928,N_2946);
nor U3433 (N_3433,N_2521,N_2679);
nor U3434 (N_3434,N_2529,N_2796);
and U3435 (N_3435,N_2561,N_2523);
nand U3436 (N_3436,N_2687,N_2571);
or U3437 (N_3437,N_2669,N_2685);
or U3438 (N_3438,N_2984,N_2504);
xor U3439 (N_3439,N_2991,N_2549);
and U3440 (N_3440,N_2966,N_2820);
nor U3441 (N_3441,N_2601,N_2973);
or U3442 (N_3442,N_2872,N_2568);
nand U3443 (N_3443,N_2803,N_2920);
nor U3444 (N_3444,N_2639,N_2623);
or U3445 (N_3445,N_2934,N_2836);
and U3446 (N_3446,N_2874,N_2818);
nand U3447 (N_3447,N_2957,N_2937);
nor U3448 (N_3448,N_2568,N_2829);
nand U3449 (N_3449,N_2982,N_2840);
nor U3450 (N_3450,N_2762,N_2981);
xnor U3451 (N_3451,N_2596,N_2752);
or U3452 (N_3452,N_2666,N_2892);
and U3453 (N_3453,N_2517,N_2966);
or U3454 (N_3454,N_2685,N_2699);
and U3455 (N_3455,N_2876,N_2712);
and U3456 (N_3456,N_2818,N_2510);
nor U3457 (N_3457,N_2703,N_2564);
or U3458 (N_3458,N_2682,N_2792);
nand U3459 (N_3459,N_2559,N_2882);
nor U3460 (N_3460,N_2785,N_2877);
nand U3461 (N_3461,N_2671,N_2682);
nor U3462 (N_3462,N_2797,N_2816);
or U3463 (N_3463,N_2873,N_2660);
nor U3464 (N_3464,N_2535,N_2765);
and U3465 (N_3465,N_2760,N_2557);
nor U3466 (N_3466,N_2580,N_2776);
or U3467 (N_3467,N_2947,N_2505);
and U3468 (N_3468,N_2953,N_2861);
nor U3469 (N_3469,N_2864,N_2994);
nor U3470 (N_3470,N_2505,N_2937);
and U3471 (N_3471,N_2927,N_2852);
and U3472 (N_3472,N_2871,N_2985);
and U3473 (N_3473,N_2758,N_2951);
and U3474 (N_3474,N_2570,N_2539);
and U3475 (N_3475,N_2669,N_2904);
and U3476 (N_3476,N_2762,N_2779);
or U3477 (N_3477,N_2583,N_2971);
nor U3478 (N_3478,N_2827,N_2735);
nor U3479 (N_3479,N_2593,N_2975);
or U3480 (N_3480,N_2625,N_2654);
or U3481 (N_3481,N_2816,N_2937);
nand U3482 (N_3482,N_2544,N_2686);
nor U3483 (N_3483,N_2947,N_2717);
nand U3484 (N_3484,N_2846,N_2528);
and U3485 (N_3485,N_2507,N_2740);
or U3486 (N_3486,N_2528,N_2748);
nor U3487 (N_3487,N_2683,N_2519);
xor U3488 (N_3488,N_2748,N_2979);
nor U3489 (N_3489,N_2987,N_2952);
nand U3490 (N_3490,N_2714,N_2873);
or U3491 (N_3491,N_2738,N_2501);
nand U3492 (N_3492,N_2515,N_2688);
and U3493 (N_3493,N_2725,N_2591);
nand U3494 (N_3494,N_2575,N_2935);
nor U3495 (N_3495,N_2568,N_2723);
and U3496 (N_3496,N_2789,N_2644);
nand U3497 (N_3497,N_2632,N_2715);
nor U3498 (N_3498,N_2779,N_2661);
or U3499 (N_3499,N_2729,N_2728);
and U3500 (N_3500,N_3324,N_3002);
or U3501 (N_3501,N_3359,N_3055);
nor U3502 (N_3502,N_3229,N_3201);
nand U3503 (N_3503,N_3266,N_3335);
nor U3504 (N_3504,N_3188,N_3400);
nor U3505 (N_3505,N_3309,N_3197);
and U3506 (N_3506,N_3088,N_3447);
nor U3507 (N_3507,N_3288,N_3427);
nand U3508 (N_3508,N_3111,N_3429);
and U3509 (N_3509,N_3273,N_3126);
or U3510 (N_3510,N_3062,N_3118);
nand U3511 (N_3511,N_3185,N_3217);
nor U3512 (N_3512,N_3078,N_3005);
or U3513 (N_3513,N_3124,N_3457);
nor U3514 (N_3514,N_3173,N_3020);
or U3515 (N_3515,N_3121,N_3384);
and U3516 (N_3516,N_3054,N_3450);
nand U3517 (N_3517,N_3113,N_3103);
nand U3518 (N_3518,N_3112,N_3455);
and U3519 (N_3519,N_3144,N_3393);
or U3520 (N_3520,N_3477,N_3049);
nand U3521 (N_3521,N_3465,N_3230);
nand U3522 (N_3522,N_3134,N_3255);
nor U3523 (N_3523,N_3192,N_3349);
nand U3524 (N_3524,N_3275,N_3278);
and U3525 (N_3525,N_3093,N_3323);
nor U3526 (N_3526,N_3357,N_3166);
nand U3527 (N_3527,N_3026,N_3004);
or U3528 (N_3528,N_3364,N_3321);
xnor U3529 (N_3529,N_3253,N_3237);
or U3530 (N_3530,N_3058,N_3448);
or U3531 (N_3531,N_3141,N_3155);
or U3532 (N_3532,N_3090,N_3046);
or U3533 (N_3533,N_3437,N_3325);
or U3534 (N_3534,N_3122,N_3047);
nor U3535 (N_3535,N_3070,N_3310);
nand U3536 (N_3536,N_3249,N_3159);
or U3537 (N_3537,N_3360,N_3085);
or U3538 (N_3538,N_3394,N_3351);
nor U3539 (N_3539,N_3081,N_3101);
nor U3540 (N_3540,N_3180,N_3304);
nor U3541 (N_3541,N_3276,N_3379);
and U3542 (N_3542,N_3277,N_3095);
nor U3543 (N_3543,N_3153,N_3072);
and U3544 (N_3544,N_3075,N_3080);
and U3545 (N_3545,N_3162,N_3445);
and U3546 (N_3546,N_3387,N_3116);
and U3547 (N_3547,N_3438,N_3066);
nand U3548 (N_3548,N_3428,N_3163);
nand U3549 (N_3549,N_3301,N_3326);
nor U3550 (N_3550,N_3274,N_3038);
nor U3551 (N_3551,N_3355,N_3411);
xnor U3552 (N_3552,N_3403,N_3099);
or U3553 (N_3553,N_3143,N_3263);
or U3554 (N_3554,N_3297,N_3286);
nor U3555 (N_3555,N_3036,N_3202);
nand U3556 (N_3556,N_3439,N_3287);
or U3557 (N_3557,N_3133,N_3389);
or U3558 (N_3558,N_3493,N_3446);
or U3559 (N_3559,N_3014,N_3233);
and U3560 (N_3560,N_3084,N_3092);
nor U3561 (N_3561,N_3495,N_3187);
or U3562 (N_3562,N_3258,N_3397);
or U3563 (N_3563,N_3425,N_3454);
nor U3564 (N_3564,N_3262,N_3399);
nor U3565 (N_3565,N_3151,N_3214);
or U3566 (N_3566,N_3369,N_3198);
nand U3567 (N_3567,N_3030,N_3234);
nor U3568 (N_3568,N_3145,N_3097);
nand U3569 (N_3569,N_3183,N_3486);
nor U3570 (N_3570,N_3045,N_3102);
or U3571 (N_3571,N_3096,N_3021);
and U3572 (N_3572,N_3068,N_3009);
or U3573 (N_3573,N_3337,N_3373);
and U3574 (N_3574,N_3247,N_3320);
and U3575 (N_3575,N_3347,N_3430);
nor U3576 (N_3576,N_3472,N_3057);
or U3577 (N_3577,N_3031,N_3125);
and U3578 (N_3578,N_3327,N_3231);
and U3579 (N_3579,N_3462,N_3223);
or U3580 (N_3580,N_3254,N_3205);
nand U3581 (N_3581,N_3395,N_3140);
or U3582 (N_3582,N_3060,N_3458);
nor U3583 (N_3583,N_3160,N_3339);
nand U3584 (N_3584,N_3407,N_3041);
nor U3585 (N_3585,N_3268,N_3479);
nor U3586 (N_3586,N_3176,N_3476);
or U3587 (N_3587,N_3181,N_3494);
and U3588 (N_3588,N_3006,N_3353);
or U3589 (N_3589,N_3216,N_3418);
and U3590 (N_3590,N_3414,N_3423);
nand U3591 (N_3591,N_3182,N_3239);
or U3592 (N_3592,N_3289,N_3451);
nand U3593 (N_3593,N_3256,N_3361);
nand U3594 (N_3594,N_3138,N_3385);
or U3595 (N_3595,N_3149,N_3232);
or U3596 (N_3596,N_3100,N_3257);
nand U3597 (N_3597,N_3416,N_3105);
xor U3598 (N_3598,N_3039,N_3492);
and U3599 (N_3599,N_3366,N_3293);
and U3600 (N_3600,N_3392,N_3073);
nor U3601 (N_3601,N_3468,N_3435);
nand U3602 (N_3602,N_3108,N_3044);
or U3603 (N_3603,N_3146,N_3065);
nor U3604 (N_3604,N_3388,N_3147);
nand U3605 (N_3605,N_3128,N_3033);
or U3606 (N_3606,N_3077,N_3299);
nand U3607 (N_3607,N_3220,N_3442);
or U3608 (N_3608,N_3136,N_3441);
nand U3609 (N_3609,N_3246,N_3312);
or U3610 (N_3610,N_3298,N_3331);
or U3611 (N_3611,N_3482,N_3485);
nor U3612 (N_3612,N_3235,N_3212);
and U3613 (N_3613,N_3292,N_3022);
or U3614 (N_3614,N_3264,N_3076);
or U3615 (N_3615,N_3089,N_3025);
or U3616 (N_3616,N_3110,N_3417);
xor U3617 (N_3617,N_3332,N_3383);
or U3618 (N_3618,N_3377,N_3431);
nor U3619 (N_3619,N_3483,N_3484);
nand U3620 (N_3620,N_3224,N_3087);
and U3621 (N_3621,N_3291,N_3378);
nand U3622 (N_3622,N_3380,N_3426);
and U3623 (N_3623,N_3043,N_3440);
nor U3624 (N_3624,N_3114,N_3382);
xnor U3625 (N_3625,N_3210,N_3157);
and U3626 (N_3626,N_3470,N_3251);
or U3627 (N_3627,N_3244,N_3107);
and U3628 (N_3628,N_3011,N_3053);
and U3629 (N_3629,N_3333,N_3071);
or U3630 (N_3630,N_3218,N_3329);
or U3631 (N_3631,N_3091,N_3199);
and U3632 (N_3632,N_3409,N_3203);
nor U3633 (N_3633,N_3074,N_3415);
nor U3634 (N_3634,N_3139,N_3015);
and U3635 (N_3635,N_3158,N_3156);
and U3636 (N_3636,N_3282,N_3245);
and U3637 (N_3637,N_3420,N_3348);
or U3638 (N_3638,N_3432,N_3316);
nor U3639 (N_3639,N_3196,N_3318);
or U3640 (N_3640,N_3226,N_3132);
and U3641 (N_3641,N_3069,N_3017);
nor U3642 (N_3642,N_3040,N_3236);
nor U3643 (N_3643,N_3109,N_3261);
nand U3644 (N_3644,N_3152,N_3059);
xnor U3645 (N_3645,N_3123,N_3010);
nor U3646 (N_3646,N_3413,N_3478);
and U3647 (N_3647,N_3209,N_3161);
or U3648 (N_3648,N_3148,N_3365);
nor U3649 (N_3649,N_3131,N_3311);
nand U3650 (N_3650,N_3082,N_3048);
or U3651 (N_3651,N_3167,N_3368);
nor U3652 (N_3652,N_3260,N_3241);
or U3653 (N_3653,N_3221,N_3165);
or U3654 (N_3654,N_3338,N_3305);
or U3655 (N_3655,N_3193,N_3308);
or U3656 (N_3656,N_3227,N_3408);
nor U3657 (N_3657,N_3200,N_3172);
nor U3658 (N_3658,N_3027,N_3453);
nand U3659 (N_3659,N_3028,N_3404);
or U3660 (N_3660,N_3307,N_3345);
nor U3661 (N_3661,N_3341,N_3350);
nor U3662 (N_3662,N_3490,N_3272);
nand U3663 (N_3663,N_3184,N_3313);
or U3664 (N_3664,N_3186,N_3238);
nand U3665 (N_3665,N_3050,N_3051);
and U3666 (N_3666,N_3488,N_3007);
and U3667 (N_3667,N_3381,N_3164);
nor U3668 (N_3668,N_3179,N_3248);
or U3669 (N_3669,N_3390,N_3376);
and U3670 (N_3670,N_3279,N_3037);
nand U3671 (N_3671,N_3497,N_3315);
nand U3672 (N_3672,N_3356,N_3314);
and U3673 (N_3673,N_3271,N_3016);
and U3674 (N_3674,N_3391,N_3104);
and U3675 (N_3675,N_3029,N_3240);
nand U3676 (N_3676,N_3269,N_3370);
or U3677 (N_3677,N_3024,N_3285);
nor U3678 (N_3678,N_3023,N_3137);
nor U3679 (N_3679,N_3334,N_3410);
or U3680 (N_3680,N_3150,N_3018);
nand U3681 (N_3681,N_3032,N_3222);
nor U3682 (N_3682,N_3375,N_3094);
and U3683 (N_3683,N_3499,N_3191);
or U3684 (N_3684,N_3443,N_3317);
or U3685 (N_3685,N_3467,N_3405);
nand U3686 (N_3686,N_3322,N_3215);
and U3687 (N_3687,N_3174,N_3436);
nor U3688 (N_3688,N_3295,N_3463);
nor U3689 (N_3689,N_3265,N_3280);
or U3690 (N_3690,N_3098,N_3211);
and U3691 (N_3691,N_3178,N_3464);
or U3692 (N_3692,N_3401,N_3396);
nor U3693 (N_3693,N_3406,N_3194);
nor U3694 (N_3694,N_3019,N_3303);
nand U3695 (N_3695,N_3300,N_3296);
or U3696 (N_3696,N_3056,N_3067);
or U3697 (N_3697,N_3419,N_3129);
or U3698 (N_3698,N_3213,N_3371);
nand U3699 (N_3699,N_3469,N_3270);
nor U3700 (N_3700,N_3252,N_3460);
nand U3701 (N_3701,N_3306,N_3421);
nor U3702 (N_3702,N_3475,N_3452);
or U3703 (N_3703,N_3473,N_3374);
nand U3704 (N_3704,N_3363,N_3346);
or U3705 (N_3705,N_3079,N_3000);
nor U3706 (N_3706,N_3424,N_3003);
and U3707 (N_3707,N_3120,N_3228);
nand U3708 (N_3708,N_3250,N_3219);
or U3709 (N_3709,N_3127,N_3175);
nand U3710 (N_3710,N_3281,N_3117);
and U3711 (N_3711,N_3034,N_3344);
or U3712 (N_3712,N_3106,N_3284);
or U3713 (N_3713,N_3154,N_3177);
or U3714 (N_3714,N_3474,N_3362);
and U3715 (N_3715,N_3189,N_3480);
nand U3716 (N_3716,N_3456,N_3358);
and U3717 (N_3717,N_3498,N_3471);
or U3718 (N_3718,N_3061,N_3459);
nand U3719 (N_3719,N_3496,N_3243);
nor U3720 (N_3720,N_3168,N_3242);
nand U3721 (N_3721,N_3386,N_3290);
nand U3722 (N_3722,N_3086,N_3422);
nor U3723 (N_3723,N_3135,N_3013);
nand U3724 (N_3724,N_3328,N_3012);
and U3725 (N_3725,N_3319,N_3064);
xnor U3726 (N_3726,N_3170,N_3402);
nor U3727 (N_3727,N_3208,N_3206);
nand U3728 (N_3728,N_3491,N_3195);
or U3729 (N_3729,N_3142,N_3481);
nor U3730 (N_3730,N_3412,N_3302);
and U3731 (N_3731,N_3204,N_3169);
and U3732 (N_3732,N_3372,N_3267);
nand U3733 (N_3733,N_3001,N_3352);
xnor U3734 (N_3734,N_3035,N_3283);
and U3735 (N_3735,N_3354,N_3466);
nand U3736 (N_3736,N_3119,N_3444);
nor U3737 (N_3737,N_3207,N_3434);
and U3738 (N_3738,N_3433,N_3330);
nor U3739 (N_3739,N_3449,N_3343);
nand U3740 (N_3740,N_3342,N_3052);
and U3741 (N_3741,N_3294,N_3259);
and U3742 (N_3742,N_3115,N_3171);
or U3743 (N_3743,N_3487,N_3063);
nor U3744 (N_3744,N_3367,N_3398);
nand U3745 (N_3745,N_3336,N_3190);
nand U3746 (N_3746,N_3489,N_3008);
nor U3747 (N_3747,N_3083,N_3340);
and U3748 (N_3748,N_3130,N_3225);
nor U3749 (N_3749,N_3042,N_3461);
nor U3750 (N_3750,N_3288,N_3027);
or U3751 (N_3751,N_3394,N_3332);
and U3752 (N_3752,N_3373,N_3202);
and U3753 (N_3753,N_3185,N_3408);
nor U3754 (N_3754,N_3032,N_3329);
or U3755 (N_3755,N_3308,N_3337);
nor U3756 (N_3756,N_3190,N_3209);
and U3757 (N_3757,N_3113,N_3161);
or U3758 (N_3758,N_3031,N_3172);
and U3759 (N_3759,N_3200,N_3376);
nor U3760 (N_3760,N_3099,N_3122);
nor U3761 (N_3761,N_3093,N_3000);
nor U3762 (N_3762,N_3444,N_3252);
and U3763 (N_3763,N_3166,N_3265);
nor U3764 (N_3764,N_3061,N_3242);
nor U3765 (N_3765,N_3063,N_3462);
nor U3766 (N_3766,N_3496,N_3163);
and U3767 (N_3767,N_3491,N_3191);
nor U3768 (N_3768,N_3309,N_3387);
or U3769 (N_3769,N_3220,N_3396);
nor U3770 (N_3770,N_3059,N_3425);
or U3771 (N_3771,N_3349,N_3024);
or U3772 (N_3772,N_3293,N_3282);
and U3773 (N_3773,N_3063,N_3261);
nand U3774 (N_3774,N_3182,N_3058);
or U3775 (N_3775,N_3030,N_3077);
nor U3776 (N_3776,N_3400,N_3488);
nor U3777 (N_3777,N_3097,N_3478);
nand U3778 (N_3778,N_3227,N_3169);
and U3779 (N_3779,N_3273,N_3191);
nand U3780 (N_3780,N_3306,N_3428);
or U3781 (N_3781,N_3323,N_3054);
nor U3782 (N_3782,N_3257,N_3316);
and U3783 (N_3783,N_3485,N_3309);
nand U3784 (N_3784,N_3029,N_3050);
nand U3785 (N_3785,N_3260,N_3290);
and U3786 (N_3786,N_3034,N_3463);
nand U3787 (N_3787,N_3448,N_3280);
nand U3788 (N_3788,N_3279,N_3246);
and U3789 (N_3789,N_3461,N_3097);
nand U3790 (N_3790,N_3048,N_3458);
nor U3791 (N_3791,N_3158,N_3299);
or U3792 (N_3792,N_3365,N_3085);
or U3793 (N_3793,N_3138,N_3273);
and U3794 (N_3794,N_3126,N_3374);
nand U3795 (N_3795,N_3406,N_3293);
nand U3796 (N_3796,N_3115,N_3292);
nor U3797 (N_3797,N_3162,N_3211);
and U3798 (N_3798,N_3050,N_3163);
and U3799 (N_3799,N_3288,N_3042);
or U3800 (N_3800,N_3300,N_3133);
or U3801 (N_3801,N_3401,N_3024);
and U3802 (N_3802,N_3165,N_3060);
and U3803 (N_3803,N_3080,N_3295);
nand U3804 (N_3804,N_3390,N_3031);
nand U3805 (N_3805,N_3127,N_3154);
nor U3806 (N_3806,N_3305,N_3331);
nand U3807 (N_3807,N_3379,N_3439);
or U3808 (N_3808,N_3145,N_3408);
nand U3809 (N_3809,N_3072,N_3052);
and U3810 (N_3810,N_3141,N_3125);
nand U3811 (N_3811,N_3470,N_3431);
xnor U3812 (N_3812,N_3411,N_3002);
and U3813 (N_3813,N_3360,N_3186);
xor U3814 (N_3814,N_3290,N_3253);
nor U3815 (N_3815,N_3452,N_3227);
or U3816 (N_3816,N_3365,N_3035);
and U3817 (N_3817,N_3037,N_3346);
and U3818 (N_3818,N_3222,N_3120);
nor U3819 (N_3819,N_3037,N_3143);
and U3820 (N_3820,N_3354,N_3279);
or U3821 (N_3821,N_3470,N_3186);
nand U3822 (N_3822,N_3281,N_3336);
nand U3823 (N_3823,N_3102,N_3167);
nand U3824 (N_3824,N_3095,N_3134);
or U3825 (N_3825,N_3491,N_3249);
nand U3826 (N_3826,N_3407,N_3142);
and U3827 (N_3827,N_3408,N_3495);
nor U3828 (N_3828,N_3182,N_3334);
or U3829 (N_3829,N_3267,N_3139);
nor U3830 (N_3830,N_3006,N_3476);
nor U3831 (N_3831,N_3268,N_3414);
and U3832 (N_3832,N_3075,N_3459);
and U3833 (N_3833,N_3398,N_3473);
and U3834 (N_3834,N_3208,N_3268);
nor U3835 (N_3835,N_3197,N_3130);
or U3836 (N_3836,N_3332,N_3491);
or U3837 (N_3837,N_3493,N_3235);
nand U3838 (N_3838,N_3337,N_3253);
or U3839 (N_3839,N_3455,N_3010);
and U3840 (N_3840,N_3201,N_3392);
nor U3841 (N_3841,N_3188,N_3229);
nor U3842 (N_3842,N_3271,N_3278);
and U3843 (N_3843,N_3338,N_3125);
or U3844 (N_3844,N_3005,N_3309);
and U3845 (N_3845,N_3219,N_3188);
or U3846 (N_3846,N_3297,N_3068);
nand U3847 (N_3847,N_3007,N_3333);
or U3848 (N_3848,N_3399,N_3276);
nor U3849 (N_3849,N_3192,N_3169);
nor U3850 (N_3850,N_3260,N_3448);
nand U3851 (N_3851,N_3486,N_3260);
or U3852 (N_3852,N_3495,N_3342);
and U3853 (N_3853,N_3270,N_3397);
nor U3854 (N_3854,N_3016,N_3289);
or U3855 (N_3855,N_3233,N_3299);
nor U3856 (N_3856,N_3437,N_3267);
nand U3857 (N_3857,N_3274,N_3081);
and U3858 (N_3858,N_3461,N_3267);
xor U3859 (N_3859,N_3183,N_3018);
nand U3860 (N_3860,N_3386,N_3256);
nor U3861 (N_3861,N_3013,N_3008);
nor U3862 (N_3862,N_3236,N_3466);
nor U3863 (N_3863,N_3251,N_3122);
nand U3864 (N_3864,N_3077,N_3476);
nor U3865 (N_3865,N_3443,N_3396);
nand U3866 (N_3866,N_3030,N_3025);
and U3867 (N_3867,N_3213,N_3464);
nand U3868 (N_3868,N_3471,N_3122);
nor U3869 (N_3869,N_3305,N_3276);
or U3870 (N_3870,N_3195,N_3255);
nor U3871 (N_3871,N_3188,N_3221);
or U3872 (N_3872,N_3131,N_3278);
and U3873 (N_3873,N_3333,N_3155);
nor U3874 (N_3874,N_3335,N_3390);
nor U3875 (N_3875,N_3206,N_3369);
nor U3876 (N_3876,N_3218,N_3443);
or U3877 (N_3877,N_3457,N_3430);
and U3878 (N_3878,N_3024,N_3039);
or U3879 (N_3879,N_3152,N_3005);
nand U3880 (N_3880,N_3032,N_3003);
xnor U3881 (N_3881,N_3263,N_3369);
and U3882 (N_3882,N_3456,N_3202);
and U3883 (N_3883,N_3253,N_3010);
or U3884 (N_3884,N_3199,N_3341);
and U3885 (N_3885,N_3453,N_3055);
or U3886 (N_3886,N_3201,N_3185);
or U3887 (N_3887,N_3185,N_3172);
or U3888 (N_3888,N_3218,N_3113);
nand U3889 (N_3889,N_3250,N_3205);
and U3890 (N_3890,N_3396,N_3481);
and U3891 (N_3891,N_3135,N_3208);
and U3892 (N_3892,N_3465,N_3378);
or U3893 (N_3893,N_3424,N_3404);
nor U3894 (N_3894,N_3065,N_3223);
and U3895 (N_3895,N_3473,N_3381);
nor U3896 (N_3896,N_3342,N_3436);
nand U3897 (N_3897,N_3351,N_3278);
nand U3898 (N_3898,N_3166,N_3471);
xor U3899 (N_3899,N_3454,N_3333);
or U3900 (N_3900,N_3424,N_3120);
nand U3901 (N_3901,N_3400,N_3358);
nor U3902 (N_3902,N_3386,N_3163);
xnor U3903 (N_3903,N_3345,N_3098);
xor U3904 (N_3904,N_3443,N_3430);
nor U3905 (N_3905,N_3430,N_3314);
nor U3906 (N_3906,N_3496,N_3467);
and U3907 (N_3907,N_3023,N_3178);
nor U3908 (N_3908,N_3271,N_3407);
nand U3909 (N_3909,N_3384,N_3234);
nand U3910 (N_3910,N_3079,N_3011);
nor U3911 (N_3911,N_3447,N_3426);
or U3912 (N_3912,N_3182,N_3106);
nor U3913 (N_3913,N_3387,N_3093);
nand U3914 (N_3914,N_3005,N_3301);
nor U3915 (N_3915,N_3209,N_3204);
nor U3916 (N_3916,N_3345,N_3015);
nor U3917 (N_3917,N_3438,N_3014);
nor U3918 (N_3918,N_3428,N_3019);
nand U3919 (N_3919,N_3110,N_3085);
nor U3920 (N_3920,N_3479,N_3216);
or U3921 (N_3921,N_3106,N_3103);
or U3922 (N_3922,N_3467,N_3011);
nor U3923 (N_3923,N_3191,N_3150);
or U3924 (N_3924,N_3463,N_3257);
nor U3925 (N_3925,N_3101,N_3242);
nand U3926 (N_3926,N_3489,N_3062);
or U3927 (N_3927,N_3164,N_3482);
xnor U3928 (N_3928,N_3259,N_3423);
nor U3929 (N_3929,N_3247,N_3160);
and U3930 (N_3930,N_3332,N_3481);
or U3931 (N_3931,N_3251,N_3080);
nand U3932 (N_3932,N_3309,N_3091);
nor U3933 (N_3933,N_3021,N_3111);
and U3934 (N_3934,N_3140,N_3319);
and U3935 (N_3935,N_3265,N_3003);
nand U3936 (N_3936,N_3296,N_3428);
and U3937 (N_3937,N_3161,N_3406);
nand U3938 (N_3938,N_3137,N_3493);
and U3939 (N_3939,N_3469,N_3473);
and U3940 (N_3940,N_3333,N_3386);
nor U3941 (N_3941,N_3398,N_3147);
or U3942 (N_3942,N_3284,N_3262);
nand U3943 (N_3943,N_3469,N_3156);
nand U3944 (N_3944,N_3451,N_3013);
or U3945 (N_3945,N_3296,N_3317);
xnor U3946 (N_3946,N_3027,N_3351);
nor U3947 (N_3947,N_3149,N_3438);
and U3948 (N_3948,N_3241,N_3124);
nand U3949 (N_3949,N_3288,N_3425);
or U3950 (N_3950,N_3026,N_3494);
or U3951 (N_3951,N_3279,N_3323);
nand U3952 (N_3952,N_3178,N_3342);
xor U3953 (N_3953,N_3373,N_3402);
or U3954 (N_3954,N_3106,N_3285);
and U3955 (N_3955,N_3130,N_3412);
nor U3956 (N_3956,N_3425,N_3003);
or U3957 (N_3957,N_3370,N_3015);
and U3958 (N_3958,N_3218,N_3322);
nor U3959 (N_3959,N_3351,N_3172);
nand U3960 (N_3960,N_3117,N_3186);
nand U3961 (N_3961,N_3277,N_3473);
or U3962 (N_3962,N_3130,N_3325);
and U3963 (N_3963,N_3297,N_3352);
or U3964 (N_3964,N_3075,N_3423);
or U3965 (N_3965,N_3190,N_3366);
or U3966 (N_3966,N_3129,N_3055);
nor U3967 (N_3967,N_3018,N_3314);
nor U3968 (N_3968,N_3358,N_3424);
nor U3969 (N_3969,N_3164,N_3498);
or U3970 (N_3970,N_3177,N_3014);
and U3971 (N_3971,N_3187,N_3123);
nor U3972 (N_3972,N_3328,N_3006);
or U3973 (N_3973,N_3226,N_3367);
nor U3974 (N_3974,N_3456,N_3105);
or U3975 (N_3975,N_3200,N_3092);
and U3976 (N_3976,N_3146,N_3016);
or U3977 (N_3977,N_3252,N_3313);
nand U3978 (N_3978,N_3283,N_3034);
and U3979 (N_3979,N_3100,N_3113);
nand U3980 (N_3980,N_3397,N_3421);
and U3981 (N_3981,N_3052,N_3210);
and U3982 (N_3982,N_3015,N_3172);
nor U3983 (N_3983,N_3046,N_3417);
nor U3984 (N_3984,N_3276,N_3189);
nor U3985 (N_3985,N_3068,N_3045);
nand U3986 (N_3986,N_3162,N_3104);
nand U3987 (N_3987,N_3248,N_3021);
or U3988 (N_3988,N_3177,N_3193);
nor U3989 (N_3989,N_3345,N_3072);
and U3990 (N_3990,N_3075,N_3237);
nor U3991 (N_3991,N_3469,N_3035);
xor U3992 (N_3992,N_3166,N_3074);
nand U3993 (N_3993,N_3022,N_3375);
and U3994 (N_3994,N_3153,N_3113);
and U3995 (N_3995,N_3383,N_3273);
nor U3996 (N_3996,N_3149,N_3406);
nand U3997 (N_3997,N_3160,N_3299);
or U3998 (N_3998,N_3307,N_3285);
nor U3999 (N_3999,N_3424,N_3433);
xnor U4000 (N_4000,N_3951,N_3669);
nor U4001 (N_4001,N_3687,N_3608);
nor U4002 (N_4002,N_3915,N_3550);
nor U4003 (N_4003,N_3805,N_3662);
and U4004 (N_4004,N_3749,N_3965);
nor U4005 (N_4005,N_3971,N_3892);
nand U4006 (N_4006,N_3712,N_3584);
nand U4007 (N_4007,N_3543,N_3997);
nand U4008 (N_4008,N_3974,N_3876);
nand U4009 (N_4009,N_3606,N_3764);
nor U4010 (N_4010,N_3586,N_3504);
nand U4011 (N_4011,N_3638,N_3848);
or U4012 (N_4012,N_3804,N_3928);
and U4013 (N_4013,N_3635,N_3897);
or U4014 (N_4014,N_3990,N_3941);
nand U4015 (N_4015,N_3976,N_3904);
nand U4016 (N_4016,N_3614,N_3818);
nor U4017 (N_4017,N_3806,N_3851);
or U4018 (N_4018,N_3936,N_3514);
and U4019 (N_4019,N_3700,N_3587);
nor U4020 (N_4020,N_3722,N_3561);
nand U4021 (N_4021,N_3744,N_3678);
or U4022 (N_4022,N_3991,N_3726);
and U4023 (N_4023,N_3684,N_3782);
nor U4024 (N_4024,N_3945,N_3665);
nor U4025 (N_4025,N_3560,N_3742);
and U4026 (N_4026,N_3835,N_3544);
nand U4027 (N_4027,N_3900,N_3772);
nor U4028 (N_4028,N_3747,N_3503);
or U4029 (N_4029,N_3612,N_3884);
or U4030 (N_4030,N_3737,N_3640);
and U4031 (N_4031,N_3953,N_3570);
or U4032 (N_4032,N_3911,N_3754);
or U4033 (N_4033,N_3758,N_3661);
and U4034 (N_4034,N_3527,N_3889);
or U4035 (N_4035,N_3960,N_3532);
or U4036 (N_4036,N_3610,N_3625);
and U4037 (N_4037,N_3617,N_3807);
nor U4038 (N_4038,N_3856,N_3718);
or U4039 (N_4039,N_3675,N_3773);
nor U4040 (N_4040,N_3930,N_3699);
and U4041 (N_4041,N_3698,N_3731);
or U4042 (N_4042,N_3756,N_3899);
nand U4043 (N_4043,N_3812,N_3701);
or U4044 (N_4044,N_3557,N_3748);
nor U4045 (N_4045,N_3888,N_3826);
nand U4046 (N_4046,N_3735,N_3705);
nor U4047 (N_4047,N_3575,N_3738);
and U4048 (N_4048,N_3829,N_3693);
nand U4049 (N_4049,N_3592,N_3548);
or U4050 (N_4050,N_3688,N_3502);
or U4051 (N_4051,N_3916,N_3950);
nand U4052 (N_4052,N_3552,N_3602);
nor U4053 (N_4053,N_3598,N_3942);
nand U4054 (N_4054,N_3949,N_3647);
nor U4055 (N_4055,N_3834,N_3792);
and U4056 (N_4056,N_3717,N_3978);
and U4057 (N_4057,N_3719,N_3946);
and U4058 (N_4058,N_3566,N_3538);
nand U4059 (N_4059,N_3879,N_3524);
and U4060 (N_4060,N_3767,N_3788);
and U4061 (N_4061,N_3968,N_3702);
nand U4062 (N_4062,N_3667,N_3676);
or U4063 (N_4063,N_3952,N_3556);
nand U4064 (N_4064,N_3793,N_3808);
nor U4065 (N_4065,N_3810,N_3873);
or U4066 (N_4066,N_3721,N_3816);
nor U4067 (N_4067,N_3781,N_3506);
nor U4068 (N_4068,N_3644,N_3565);
nand U4069 (N_4069,N_3992,N_3551);
and U4070 (N_4070,N_3609,N_3740);
nand U4071 (N_4071,N_3890,N_3594);
or U4072 (N_4072,N_3853,N_3878);
and U4073 (N_4073,N_3755,N_3935);
or U4074 (N_4074,N_3639,N_3857);
or U4075 (N_4075,N_3983,N_3901);
or U4076 (N_4076,N_3515,N_3814);
xor U4077 (N_4077,N_3875,N_3648);
nand U4078 (N_4078,N_3802,N_3618);
nor U4079 (N_4079,N_3547,N_3613);
xnor U4080 (N_4080,N_3832,N_3530);
nand U4081 (N_4081,N_3521,N_3574);
and U4082 (N_4082,N_3939,N_3633);
or U4083 (N_4083,N_3862,N_3553);
nor U4084 (N_4084,N_3562,N_3512);
nand U4085 (N_4085,N_3604,N_3616);
or U4086 (N_4086,N_3933,N_3671);
nor U4087 (N_4087,N_3603,N_3760);
or U4088 (N_4088,N_3985,N_3670);
nor U4089 (N_4089,N_3860,N_3572);
or U4090 (N_4090,N_3993,N_3607);
nand U4091 (N_4091,N_3868,N_3745);
or U4092 (N_4092,N_3882,N_3843);
or U4093 (N_4093,N_3771,N_3822);
and U4094 (N_4094,N_3659,N_3836);
and U4095 (N_4095,N_3679,N_3922);
nand U4096 (N_4096,N_3967,N_3864);
nand U4097 (N_4097,N_3918,N_3513);
or U4098 (N_4098,N_3927,N_3919);
nand U4099 (N_4099,N_3519,N_3711);
and U4100 (N_4100,N_3716,N_3925);
and U4101 (N_4101,N_3668,N_3894);
and U4102 (N_4102,N_3697,N_3599);
and U4103 (N_4103,N_3528,N_3710);
nor U4104 (N_4104,N_3923,N_3652);
nand U4105 (N_4105,N_3902,N_3752);
or U4106 (N_4106,N_3563,N_3629);
and U4107 (N_4107,N_3650,N_3893);
and U4108 (N_4108,N_3943,N_3877);
or U4109 (N_4109,N_3507,N_3725);
nand U4110 (N_4110,N_3837,N_3695);
or U4111 (N_4111,N_3982,N_3932);
nand U4112 (N_4112,N_3645,N_3770);
nand U4113 (N_4113,N_3987,N_3981);
and U4114 (N_4114,N_3641,N_3526);
and U4115 (N_4115,N_3558,N_3820);
nor U4116 (N_4116,N_3909,N_3580);
or U4117 (N_4117,N_3801,N_3654);
nor U4118 (N_4118,N_3605,N_3830);
or U4119 (N_4119,N_3871,N_3611);
nor U4120 (N_4120,N_3912,N_3582);
nand U4121 (N_4121,N_3954,N_3692);
and U4122 (N_4122,N_3914,N_3757);
or U4123 (N_4123,N_3841,N_3510);
or U4124 (N_4124,N_3948,N_3903);
and U4125 (N_4125,N_3833,N_3555);
nand U4126 (N_4126,N_3730,N_3531);
and U4127 (N_4127,N_3989,N_3784);
and U4128 (N_4128,N_3739,N_3913);
nand U4129 (N_4129,N_3880,N_3601);
nand U4130 (N_4130,N_3621,N_3959);
nand U4131 (N_4131,N_3958,N_3777);
nand U4132 (N_4132,N_3940,N_3628);
and U4133 (N_4133,N_3746,N_3803);
nand U4134 (N_4134,N_3597,N_3724);
nand U4135 (N_4135,N_3714,N_3651);
or U4136 (N_4136,N_3559,N_3674);
nand U4137 (N_4137,N_3720,N_3783);
nand U4138 (N_4138,N_3799,N_3984);
or U4139 (N_4139,N_3655,N_3680);
nor U4140 (N_4140,N_3986,N_3677);
nand U4141 (N_4141,N_3500,N_3774);
and U4142 (N_4142,N_3931,N_3998);
and U4143 (N_4143,N_3649,N_3637);
nor U4144 (N_4144,N_3588,N_3850);
or U4145 (N_4145,N_3765,N_3769);
and U4146 (N_4146,N_3620,N_3685);
nor U4147 (N_4147,N_3536,N_3794);
and U4148 (N_4148,N_3861,N_3529);
and U4149 (N_4149,N_3980,N_3977);
and U4150 (N_4150,N_3780,N_3908);
or U4151 (N_4151,N_3589,N_3751);
and U4152 (N_4152,N_3694,N_3569);
nand U4153 (N_4153,N_3966,N_3706);
nand U4154 (N_4154,N_3576,N_3713);
nand U4155 (N_4155,N_3775,N_3673);
nor U4156 (N_4156,N_3535,N_3944);
and U4157 (N_4157,N_3627,N_3790);
or U4158 (N_4158,N_3631,N_3579);
nand U4159 (N_4159,N_3623,N_3663);
or U4160 (N_4160,N_3938,N_3591);
or U4161 (N_4161,N_3866,N_3929);
nand U4162 (N_4162,N_3859,N_3682);
nand U4163 (N_4163,N_3509,N_3729);
and U4164 (N_4164,N_3956,N_3615);
nand U4165 (N_4165,N_3750,N_3549);
or U4166 (N_4166,N_3955,N_3917);
nor U4167 (N_4167,N_3683,N_3821);
or U4168 (N_4168,N_3568,N_3518);
and U4169 (N_4169,N_3858,N_3786);
or U4170 (N_4170,N_3844,N_3508);
or U4171 (N_4171,N_3846,N_3653);
nand U4172 (N_4172,N_3728,N_3578);
nand U4173 (N_4173,N_3595,N_3619);
nor U4174 (N_4174,N_3957,N_3567);
nor U4175 (N_4175,N_3534,N_3874);
nand U4176 (N_4176,N_3734,N_3704);
or U4177 (N_4177,N_3691,N_3854);
nor U4178 (N_4178,N_3828,N_3554);
or U4179 (N_4179,N_3525,N_3642);
nor U4180 (N_4180,N_3824,N_3907);
nand U4181 (N_4181,N_3845,N_3753);
nor U4182 (N_4182,N_3847,N_3800);
and U4183 (N_4183,N_3947,N_3827);
or U4184 (N_4184,N_3863,N_3995);
nand U4185 (N_4185,N_3522,N_3672);
and U4186 (N_4186,N_3811,N_3779);
or U4187 (N_4187,N_3516,N_3732);
nand U4188 (N_4188,N_3798,N_3520);
or U4189 (N_4189,N_3924,N_3964);
and U4190 (N_4190,N_3823,N_3994);
nand U4191 (N_4191,N_3763,N_3539);
xnor U4192 (N_4192,N_3795,N_3869);
and U4193 (N_4193,N_3590,N_3660);
nor U4194 (N_4194,N_3926,N_3778);
nand U4195 (N_4195,N_3896,N_3715);
and U4196 (N_4196,N_3624,N_3839);
and U4197 (N_4197,N_3962,N_3961);
and U4198 (N_4198,N_3761,N_3690);
and U4199 (N_4199,N_3921,N_3577);
or U4200 (N_4200,N_3870,N_3583);
and U4201 (N_4201,N_3523,N_3809);
and U4202 (N_4202,N_3643,N_3842);
and U4203 (N_4203,N_3813,N_3664);
or U4204 (N_4204,N_3666,N_3979);
or U4205 (N_4205,N_3585,N_3886);
nand U4206 (N_4206,N_3825,N_3972);
nor U4207 (N_4207,N_3840,N_3564);
or U4208 (N_4208,N_3630,N_3727);
and U4209 (N_4209,N_3872,N_3831);
or U4210 (N_4210,N_3849,N_3838);
nor U4211 (N_4211,N_3681,N_3634);
or U4212 (N_4212,N_3571,N_3545);
nand U4213 (N_4213,N_3656,N_3895);
nor U4214 (N_4214,N_3626,N_3776);
and U4215 (N_4215,N_3581,N_3787);
and U4216 (N_4216,N_3791,N_3885);
nor U4217 (N_4217,N_3759,N_3906);
nor U4218 (N_4218,N_3540,N_3658);
nor U4219 (N_4219,N_3970,N_3593);
or U4220 (N_4220,N_3815,N_3689);
nand U4221 (N_4221,N_3785,N_3546);
or U4222 (N_4222,N_3797,N_3969);
or U4223 (N_4223,N_3517,N_3696);
nand U4224 (N_4224,N_3999,N_3867);
nand U4225 (N_4225,N_3622,N_3511);
nor U4226 (N_4226,N_3686,N_3646);
nand U4227 (N_4227,N_3819,N_3852);
and U4228 (N_4228,N_3736,N_3723);
or U4229 (N_4229,N_3766,N_3501);
nor U4230 (N_4230,N_3898,N_3636);
or U4231 (N_4231,N_3505,N_3533);
nor U4232 (N_4232,N_3703,N_3817);
nor U4233 (N_4233,N_3600,N_3865);
or U4234 (N_4234,N_3743,N_3937);
nand U4235 (N_4235,N_3789,N_3596);
nor U4236 (N_4236,N_3988,N_3762);
and U4237 (N_4237,N_3920,N_3573);
and U4238 (N_4238,N_3768,N_3881);
and U4239 (N_4239,N_3709,N_3934);
nand U4240 (N_4240,N_3973,N_3632);
nor U4241 (N_4241,N_3708,N_3796);
and U4242 (N_4242,N_3707,N_3542);
nor U4243 (N_4243,N_3996,N_3537);
and U4244 (N_4244,N_3883,N_3741);
nor U4245 (N_4245,N_3855,N_3891);
and U4246 (N_4246,N_3657,N_3975);
nand U4247 (N_4247,N_3910,N_3541);
nor U4248 (N_4248,N_3887,N_3905);
nor U4249 (N_4249,N_3733,N_3963);
nor U4250 (N_4250,N_3695,N_3725);
and U4251 (N_4251,N_3689,N_3970);
or U4252 (N_4252,N_3811,N_3951);
nor U4253 (N_4253,N_3527,N_3946);
and U4254 (N_4254,N_3565,N_3991);
nand U4255 (N_4255,N_3608,N_3916);
and U4256 (N_4256,N_3574,N_3994);
nor U4257 (N_4257,N_3843,N_3759);
nand U4258 (N_4258,N_3593,N_3764);
xor U4259 (N_4259,N_3691,N_3898);
and U4260 (N_4260,N_3661,N_3865);
nand U4261 (N_4261,N_3895,N_3690);
nand U4262 (N_4262,N_3923,N_3562);
nor U4263 (N_4263,N_3548,N_3614);
nor U4264 (N_4264,N_3705,N_3547);
or U4265 (N_4265,N_3781,N_3792);
nand U4266 (N_4266,N_3912,N_3659);
nand U4267 (N_4267,N_3556,N_3754);
nor U4268 (N_4268,N_3825,N_3697);
nand U4269 (N_4269,N_3755,N_3977);
nor U4270 (N_4270,N_3524,N_3817);
or U4271 (N_4271,N_3777,N_3872);
nand U4272 (N_4272,N_3530,N_3527);
or U4273 (N_4273,N_3944,N_3862);
and U4274 (N_4274,N_3925,N_3625);
nand U4275 (N_4275,N_3604,N_3820);
and U4276 (N_4276,N_3535,N_3719);
and U4277 (N_4277,N_3523,N_3975);
or U4278 (N_4278,N_3888,N_3898);
nor U4279 (N_4279,N_3983,N_3602);
and U4280 (N_4280,N_3602,N_3860);
and U4281 (N_4281,N_3794,N_3611);
nor U4282 (N_4282,N_3858,N_3890);
nor U4283 (N_4283,N_3814,N_3891);
and U4284 (N_4284,N_3893,N_3568);
nand U4285 (N_4285,N_3886,N_3815);
nor U4286 (N_4286,N_3941,N_3980);
nor U4287 (N_4287,N_3715,N_3725);
or U4288 (N_4288,N_3590,N_3521);
and U4289 (N_4289,N_3730,N_3897);
or U4290 (N_4290,N_3715,N_3548);
nand U4291 (N_4291,N_3645,N_3831);
nor U4292 (N_4292,N_3602,N_3578);
or U4293 (N_4293,N_3528,N_3627);
nand U4294 (N_4294,N_3959,N_3726);
nand U4295 (N_4295,N_3554,N_3718);
nor U4296 (N_4296,N_3915,N_3971);
or U4297 (N_4297,N_3801,N_3800);
nor U4298 (N_4298,N_3744,N_3886);
xnor U4299 (N_4299,N_3893,N_3840);
and U4300 (N_4300,N_3899,N_3832);
nor U4301 (N_4301,N_3780,N_3748);
or U4302 (N_4302,N_3632,N_3993);
and U4303 (N_4303,N_3634,N_3650);
nor U4304 (N_4304,N_3606,N_3600);
or U4305 (N_4305,N_3838,N_3654);
and U4306 (N_4306,N_3639,N_3955);
nand U4307 (N_4307,N_3931,N_3886);
or U4308 (N_4308,N_3861,N_3949);
or U4309 (N_4309,N_3658,N_3661);
nor U4310 (N_4310,N_3664,N_3750);
or U4311 (N_4311,N_3648,N_3596);
nor U4312 (N_4312,N_3743,N_3776);
or U4313 (N_4313,N_3749,N_3993);
nor U4314 (N_4314,N_3606,N_3598);
xnor U4315 (N_4315,N_3755,N_3539);
or U4316 (N_4316,N_3745,N_3681);
nand U4317 (N_4317,N_3590,N_3618);
nor U4318 (N_4318,N_3765,N_3732);
nand U4319 (N_4319,N_3649,N_3911);
nand U4320 (N_4320,N_3652,N_3577);
nor U4321 (N_4321,N_3658,N_3951);
and U4322 (N_4322,N_3851,N_3625);
or U4323 (N_4323,N_3808,N_3897);
nand U4324 (N_4324,N_3701,N_3972);
and U4325 (N_4325,N_3668,N_3910);
nand U4326 (N_4326,N_3988,N_3707);
nor U4327 (N_4327,N_3913,N_3546);
nor U4328 (N_4328,N_3937,N_3822);
nand U4329 (N_4329,N_3981,N_3614);
nand U4330 (N_4330,N_3862,N_3735);
or U4331 (N_4331,N_3734,N_3669);
or U4332 (N_4332,N_3537,N_3917);
and U4333 (N_4333,N_3902,N_3882);
nand U4334 (N_4334,N_3845,N_3543);
or U4335 (N_4335,N_3807,N_3620);
and U4336 (N_4336,N_3640,N_3825);
nor U4337 (N_4337,N_3688,N_3956);
and U4338 (N_4338,N_3830,N_3894);
or U4339 (N_4339,N_3555,N_3980);
nand U4340 (N_4340,N_3555,N_3923);
nand U4341 (N_4341,N_3755,N_3747);
xor U4342 (N_4342,N_3782,N_3707);
or U4343 (N_4343,N_3564,N_3720);
nand U4344 (N_4344,N_3903,N_3947);
or U4345 (N_4345,N_3703,N_3780);
or U4346 (N_4346,N_3844,N_3538);
xnor U4347 (N_4347,N_3878,N_3896);
and U4348 (N_4348,N_3636,N_3913);
or U4349 (N_4349,N_3983,N_3506);
and U4350 (N_4350,N_3591,N_3751);
nand U4351 (N_4351,N_3531,N_3803);
nor U4352 (N_4352,N_3552,N_3826);
nand U4353 (N_4353,N_3925,N_3527);
nor U4354 (N_4354,N_3850,N_3600);
nand U4355 (N_4355,N_3682,N_3890);
nand U4356 (N_4356,N_3515,N_3917);
nand U4357 (N_4357,N_3689,N_3938);
nand U4358 (N_4358,N_3615,N_3761);
and U4359 (N_4359,N_3578,N_3708);
or U4360 (N_4360,N_3938,N_3565);
and U4361 (N_4361,N_3581,N_3669);
nor U4362 (N_4362,N_3654,N_3699);
nor U4363 (N_4363,N_3992,N_3609);
nor U4364 (N_4364,N_3759,N_3772);
or U4365 (N_4365,N_3768,N_3512);
nand U4366 (N_4366,N_3685,N_3944);
nor U4367 (N_4367,N_3991,N_3608);
nor U4368 (N_4368,N_3715,N_3975);
nor U4369 (N_4369,N_3860,N_3892);
or U4370 (N_4370,N_3916,N_3809);
and U4371 (N_4371,N_3535,N_3800);
nor U4372 (N_4372,N_3779,N_3565);
nand U4373 (N_4373,N_3743,N_3708);
or U4374 (N_4374,N_3792,N_3593);
nand U4375 (N_4375,N_3647,N_3753);
or U4376 (N_4376,N_3822,N_3750);
or U4377 (N_4377,N_3833,N_3797);
and U4378 (N_4378,N_3837,N_3712);
nand U4379 (N_4379,N_3722,N_3693);
nor U4380 (N_4380,N_3523,N_3531);
nor U4381 (N_4381,N_3551,N_3682);
nand U4382 (N_4382,N_3665,N_3705);
or U4383 (N_4383,N_3879,N_3548);
nor U4384 (N_4384,N_3591,N_3611);
nor U4385 (N_4385,N_3983,N_3657);
or U4386 (N_4386,N_3992,N_3850);
and U4387 (N_4387,N_3624,N_3722);
nor U4388 (N_4388,N_3559,N_3681);
and U4389 (N_4389,N_3949,N_3702);
and U4390 (N_4390,N_3733,N_3965);
and U4391 (N_4391,N_3746,N_3885);
nor U4392 (N_4392,N_3632,N_3701);
or U4393 (N_4393,N_3642,N_3702);
and U4394 (N_4394,N_3980,N_3707);
xnor U4395 (N_4395,N_3877,N_3784);
and U4396 (N_4396,N_3943,N_3566);
and U4397 (N_4397,N_3664,N_3858);
and U4398 (N_4398,N_3531,N_3505);
nor U4399 (N_4399,N_3863,N_3914);
or U4400 (N_4400,N_3760,N_3630);
or U4401 (N_4401,N_3649,N_3739);
nor U4402 (N_4402,N_3635,N_3679);
nand U4403 (N_4403,N_3955,N_3644);
xor U4404 (N_4404,N_3798,N_3933);
and U4405 (N_4405,N_3744,N_3962);
or U4406 (N_4406,N_3859,N_3754);
or U4407 (N_4407,N_3572,N_3897);
or U4408 (N_4408,N_3533,N_3996);
and U4409 (N_4409,N_3943,N_3700);
nand U4410 (N_4410,N_3632,N_3512);
or U4411 (N_4411,N_3731,N_3948);
nor U4412 (N_4412,N_3627,N_3566);
xor U4413 (N_4413,N_3855,N_3569);
nor U4414 (N_4414,N_3969,N_3528);
nor U4415 (N_4415,N_3654,N_3641);
and U4416 (N_4416,N_3697,N_3549);
nand U4417 (N_4417,N_3533,N_3564);
nor U4418 (N_4418,N_3850,N_3572);
and U4419 (N_4419,N_3872,N_3507);
and U4420 (N_4420,N_3651,N_3652);
and U4421 (N_4421,N_3659,N_3763);
nand U4422 (N_4422,N_3660,N_3947);
and U4423 (N_4423,N_3995,N_3853);
nand U4424 (N_4424,N_3881,N_3505);
or U4425 (N_4425,N_3874,N_3681);
or U4426 (N_4426,N_3874,N_3883);
or U4427 (N_4427,N_3937,N_3568);
and U4428 (N_4428,N_3614,N_3846);
nor U4429 (N_4429,N_3925,N_3850);
or U4430 (N_4430,N_3898,N_3669);
nand U4431 (N_4431,N_3673,N_3831);
and U4432 (N_4432,N_3932,N_3525);
nor U4433 (N_4433,N_3778,N_3665);
and U4434 (N_4434,N_3551,N_3710);
or U4435 (N_4435,N_3921,N_3630);
nand U4436 (N_4436,N_3717,N_3614);
and U4437 (N_4437,N_3772,N_3523);
and U4438 (N_4438,N_3756,N_3981);
nand U4439 (N_4439,N_3720,N_3776);
nand U4440 (N_4440,N_3845,N_3629);
nor U4441 (N_4441,N_3561,N_3535);
nor U4442 (N_4442,N_3512,N_3544);
nor U4443 (N_4443,N_3682,N_3978);
nor U4444 (N_4444,N_3638,N_3532);
or U4445 (N_4445,N_3957,N_3836);
and U4446 (N_4446,N_3522,N_3721);
and U4447 (N_4447,N_3563,N_3798);
xor U4448 (N_4448,N_3801,N_3603);
nand U4449 (N_4449,N_3882,N_3697);
and U4450 (N_4450,N_3844,N_3824);
nand U4451 (N_4451,N_3820,N_3779);
nand U4452 (N_4452,N_3763,N_3536);
and U4453 (N_4453,N_3546,N_3967);
or U4454 (N_4454,N_3608,N_3837);
nor U4455 (N_4455,N_3562,N_3841);
and U4456 (N_4456,N_3890,N_3789);
nand U4457 (N_4457,N_3681,N_3582);
or U4458 (N_4458,N_3709,N_3861);
nor U4459 (N_4459,N_3964,N_3749);
or U4460 (N_4460,N_3596,N_3948);
nand U4461 (N_4461,N_3885,N_3931);
or U4462 (N_4462,N_3896,N_3854);
or U4463 (N_4463,N_3706,N_3586);
nand U4464 (N_4464,N_3706,N_3890);
or U4465 (N_4465,N_3793,N_3755);
nor U4466 (N_4466,N_3597,N_3905);
and U4467 (N_4467,N_3736,N_3814);
and U4468 (N_4468,N_3629,N_3905);
and U4469 (N_4469,N_3809,N_3878);
and U4470 (N_4470,N_3508,N_3824);
nor U4471 (N_4471,N_3746,N_3726);
and U4472 (N_4472,N_3646,N_3898);
and U4473 (N_4473,N_3800,N_3511);
or U4474 (N_4474,N_3644,N_3946);
nor U4475 (N_4475,N_3619,N_3766);
or U4476 (N_4476,N_3788,N_3702);
nor U4477 (N_4477,N_3835,N_3964);
nand U4478 (N_4478,N_3688,N_3850);
nor U4479 (N_4479,N_3803,N_3668);
and U4480 (N_4480,N_3572,N_3782);
nand U4481 (N_4481,N_3951,N_3924);
or U4482 (N_4482,N_3535,N_3976);
and U4483 (N_4483,N_3903,N_3673);
nand U4484 (N_4484,N_3945,N_3656);
nand U4485 (N_4485,N_3924,N_3709);
nor U4486 (N_4486,N_3687,N_3521);
or U4487 (N_4487,N_3569,N_3803);
and U4488 (N_4488,N_3758,N_3703);
nand U4489 (N_4489,N_3725,N_3965);
nor U4490 (N_4490,N_3585,N_3744);
nand U4491 (N_4491,N_3791,N_3514);
and U4492 (N_4492,N_3884,N_3659);
and U4493 (N_4493,N_3995,N_3575);
nand U4494 (N_4494,N_3569,N_3732);
nor U4495 (N_4495,N_3705,N_3579);
nand U4496 (N_4496,N_3788,N_3947);
nor U4497 (N_4497,N_3630,N_3970);
nor U4498 (N_4498,N_3637,N_3931);
nor U4499 (N_4499,N_3960,N_3610);
nand U4500 (N_4500,N_4152,N_4349);
nand U4501 (N_4501,N_4385,N_4125);
nor U4502 (N_4502,N_4045,N_4437);
and U4503 (N_4503,N_4314,N_4000);
nor U4504 (N_4504,N_4137,N_4283);
nand U4505 (N_4505,N_4475,N_4172);
nand U4506 (N_4506,N_4061,N_4033);
or U4507 (N_4507,N_4438,N_4022);
nand U4508 (N_4508,N_4354,N_4259);
or U4509 (N_4509,N_4043,N_4367);
nor U4510 (N_4510,N_4315,N_4491);
or U4511 (N_4511,N_4405,N_4142);
nand U4512 (N_4512,N_4424,N_4490);
nand U4513 (N_4513,N_4285,N_4143);
or U4514 (N_4514,N_4038,N_4151);
nand U4515 (N_4515,N_4436,N_4433);
or U4516 (N_4516,N_4295,N_4399);
or U4517 (N_4517,N_4124,N_4128);
nand U4518 (N_4518,N_4266,N_4458);
and U4519 (N_4519,N_4431,N_4463);
or U4520 (N_4520,N_4177,N_4341);
or U4521 (N_4521,N_4225,N_4374);
nand U4522 (N_4522,N_4292,N_4461);
and U4523 (N_4523,N_4272,N_4174);
nand U4524 (N_4524,N_4443,N_4345);
or U4525 (N_4525,N_4060,N_4157);
nand U4526 (N_4526,N_4440,N_4231);
or U4527 (N_4527,N_4370,N_4120);
nor U4528 (N_4528,N_4027,N_4485);
nor U4529 (N_4529,N_4401,N_4300);
and U4530 (N_4530,N_4081,N_4209);
or U4531 (N_4531,N_4105,N_4403);
or U4532 (N_4532,N_4323,N_4183);
nand U4533 (N_4533,N_4141,N_4132);
and U4534 (N_4534,N_4025,N_4145);
or U4535 (N_4535,N_4013,N_4052);
and U4536 (N_4536,N_4050,N_4393);
and U4537 (N_4537,N_4104,N_4406);
or U4538 (N_4538,N_4037,N_4087);
nor U4539 (N_4539,N_4469,N_4054);
nor U4540 (N_4540,N_4304,N_4211);
xor U4541 (N_4541,N_4257,N_4428);
nor U4542 (N_4542,N_4254,N_4416);
nor U4543 (N_4543,N_4115,N_4144);
or U4544 (N_4544,N_4189,N_4070);
or U4545 (N_4545,N_4414,N_4150);
or U4546 (N_4546,N_4237,N_4378);
nand U4547 (N_4547,N_4123,N_4277);
nand U4548 (N_4548,N_4200,N_4146);
nor U4549 (N_4549,N_4351,N_4094);
or U4550 (N_4550,N_4460,N_4446);
nor U4551 (N_4551,N_4488,N_4334);
nand U4552 (N_4552,N_4243,N_4324);
and U4553 (N_4553,N_4455,N_4441);
and U4554 (N_4554,N_4319,N_4357);
nor U4555 (N_4555,N_4239,N_4148);
nand U4556 (N_4556,N_4079,N_4307);
nand U4557 (N_4557,N_4364,N_4264);
nor U4558 (N_4558,N_4008,N_4019);
nor U4559 (N_4559,N_4076,N_4289);
nor U4560 (N_4560,N_4130,N_4365);
and U4561 (N_4561,N_4193,N_4109);
nor U4562 (N_4562,N_4486,N_4082);
nor U4563 (N_4563,N_4179,N_4470);
or U4564 (N_4564,N_4096,N_4339);
nor U4565 (N_4565,N_4227,N_4030);
nand U4566 (N_4566,N_4474,N_4260);
or U4567 (N_4567,N_4497,N_4242);
nand U4568 (N_4568,N_4164,N_4078);
or U4569 (N_4569,N_4086,N_4282);
xnor U4570 (N_4570,N_4232,N_4217);
nor U4571 (N_4571,N_4298,N_4447);
and U4572 (N_4572,N_4454,N_4473);
nor U4573 (N_4573,N_4095,N_4340);
nand U4574 (N_4574,N_4024,N_4212);
and U4575 (N_4575,N_4034,N_4176);
or U4576 (N_4576,N_4249,N_4267);
and U4577 (N_4577,N_4149,N_4090);
nand U4578 (N_4578,N_4333,N_4253);
or U4579 (N_4579,N_4065,N_4114);
nor U4580 (N_4580,N_4317,N_4201);
nand U4581 (N_4581,N_4041,N_4384);
nor U4582 (N_4582,N_4325,N_4139);
and U4583 (N_4583,N_4064,N_4493);
or U4584 (N_4584,N_4245,N_4388);
nor U4585 (N_4585,N_4080,N_4326);
or U4586 (N_4586,N_4091,N_4156);
and U4587 (N_4587,N_4417,N_4450);
nand U4588 (N_4588,N_4359,N_4067);
nand U4589 (N_4589,N_4336,N_4097);
nand U4590 (N_4590,N_4166,N_4444);
or U4591 (N_4591,N_4484,N_4412);
or U4592 (N_4592,N_4422,N_4400);
nand U4593 (N_4593,N_4425,N_4346);
nor U4594 (N_4594,N_4330,N_4467);
and U4595 (N_4595,N_4495,N_4187);
or U4596 (N_4596,N_4386,N_4396);
and U4597 (N_4597,N_4499,N_4026);
and U4598 (N_4598,N_4219,N_4310);
nor U4599 (N_4599,N_4280,N_4498);
or U4600 (N_4600,N_4459,N_4236);
and U4601 (N_4601,N_4246,N_4186);
and U4602 (N_4602,N_4274,N_4286);
nand U4603 (N_4603,N_4464,N_4153);
nor U4604 (N_4604,N_4299,N_4119);
nand U4605 (N_4605,N_4205,N_4049);
and U4606 (N_4606,N_4244,N_4126);
or U4607 (N_4607,N_4099,N_4462);
nor U4608 (N_4608,N_4077,N_4398);
and U4609 (N_4609,N_4407,N_4453);
and U4610 (N_4610,N_4221,N_4110);
nand U4611 (N_4611,N_4291,N_4048);
nor U4612 (N_4612,N_4430,N_4442);
nor U4613 (N_4613,N_4207,N_4308);
nor U4614 (N_4614,N_4039,N_4083);
and U4615 (N_4615,N_4181,N_4046);
or U4616 (N_4616,N_4210,N_4262);
nand U4617 (N_4617,N_4465,N_4409);
or U4618 (N_4618,N_4103,N_4411);
nor U4619 (N_4619,N_4456,N_4418);
or U4620 (N_4620,N_4057,N_4016);
nand U4621 (N_4621,N_4047,N_4483);
nor U4622 (N_4622,N_4014,N_4387);
and U4623 (N_4623,N_4352,N_4101);
and U4624 (N_4624,N_4371,N_4092);
nand U4625 (N_4625,N_4098,N_4466);
nand U4626 (N_4626,N_4328,N_4084);
and U4627 (N_4627,N_4382,N_4158);
and U4628 (N_4628,N_4363,N_4389);
nor U4629 (N_4629,N_4452,N_4439);
nand U4630 (N_4630,N_4215,N_4127);
or U4631 (N_4631,N_4372,N_4163);
or U4632 (N_4632,N_4147,N_4068);
nor U4633 (N_4633,N_4226,N_4492);
or U4634 (N_4634,N_4111,N_4121);
and U4635 (N_4635,N_4036,N_4481);
nand U4636 (N_4636,N_4251,N_4250);
and U4637 (N_4637,N_4290,N_4348);
nand U4638 (N_4638,N_4356,N_4162);
nand U4639 (N_4639,N_4294,N_4408);
or U4640 (N_4640,N_4020,N_4276);
or U4641 (N_4641,N_4305,N_4224);
nor U4642 (N_4642,N_4032,N_4358);
or U4643 (N_4643,N_4381,N_4191);
nor U4644 (N_4644,N_4368,N_4471);
nand U4645 (N_4645,N_4380,N_4252);
nor U4646 (N_4646,N_4180,N_4154);
nand U4647 (N_4647,N_4185,N_4268);
nor U4648 (N_4648,N_4161,N_4190);
nor U4649 (N_4649,N_4035,N_4001);
and U4650 (N_4650,N_4197,N_4220);
nand U4651 (N_4651,N_4093,N_4017);
nor U4652 (N_4652,N_4496,N_4122);
and U4653 (N_4653,N_4106,N_4168);
nor U4654 (N_4654,N_4420,N_4131);
nor U4655 (N_4655,N_4331,N_4353);
or U4656 (N_4656,N_4136,N_4021);
and U4657 (N_4657,N_4195,N_4373);
nand U4658 (N_4658,N_4015,N_4165);
and U4659 (N_4659,N_4265,N_4029);
and U4660 (N_4660,N_4023,N_4002);
or U4661 (N_4661,N_4214,N_4432);
nand U4662 (N_4662,N_4012,N_4392);
nand U4663 (N_4663,N_4489,N_4275);
or U4664 (N_4664,N_4167,N_4322);
nand U4665 (N_4665,N_4263,N_4301);
and U4666 (N_4666,N_4062,N_4413);
xor U4667 (N_4667,N_4184,N_4306);
or U4668 (N_4668,N_4391,N_4297);
and U4669 (N_4669,N_4222,N_4028);
and U4670 (N_4670,N_4332,N_4476);
or U4671 (N_4671,N_4108,N_4366);
or U4672 (N_4672,N_4051,N_4451);
nand U4673 (N_4673,N_4230,N_4318);
or U4674 (N_4674,N_4006,N_4479);
nand U4675 (N_4675,N_4112,N_4009);
nand U4676 (N_4676,N_4063,N_4194);
or U4677 (N_4677,N_4040,N_4261);
and U4678 (N_4678,N_4390,N_4445);
nand U4679 (N_4679,N_4247,N_4404);
nor U4680 (N_4680,N_4281,N_4102);
or U4681 (N_4681,N_4178,N_4415);
or U4682 (N_4682,N_4160,N_4256);
nor U4683 (N_4683,N_4419,N_4196);
or U4684 (N_4684,N_4229,N_4004);
or U4685 (N_4685,N_4271,N_4360);
nor U4686 (N_4686,N_4296,N_4171);
nor U4687 (N_4687,N_4206,N_4423);
and U4688 (N_4688,N_4233,N_4394);
or U4689 (N_4689,N_4369,N_4182);
or U4690 (N_4690,N_4118,N_4003);
nand U4691 (N_4691,N_4449,N_4329);
or U4692 (N_4692,N_4059,N_4042);
nor U4693 (N_4693,N_4175,N_4117);
nand U4694 (N_4694,N_4395,N_4288);
nand U4695 (N_4695,N_4347,N_4427);
or U4696 (N_4696,N_4069,N_4056);
nand U4697 (N_4697,N_4216,N_4173);
or U4698 (N_4698,N_4159,N_4134);
nor U4699 (N_4699,N_4335,N_4170);
or U4700 (N_4700,N_4255,N_4478);
nand U4701 (N_4701,N_4066,N_4075);
and U4702 (N_4702,N_4313,N_4107);
or U4703 (N_4703,N_4343,N_4434);
or U4704 (N_4704,N_4203,N_4435);
nand U4705 (N_4705,N_4248,N_4129);
nand U4706 (N_4706,N_4113,N_4031);
and U4707 (N_4707,N_4278,N_4477);
nand U4708 (N_4708,N_4344,N_4426);
nor U4709 (N_4709,N_4338,N_4018);
nand U4710 (N_4710,N_4058,N_4169);
nand U4711 (N_4711,N_4055,N_4073);
nand U4712 (N_4712,N_4379,N_4342);
nor U4713 (N_4713,N_4355,N_4457);
nand U4714 (N_4714,N_4402,N_4472);
nand U4715 (N_4715,N_4258,N_4273);
and U4716 (N_4716,N_4053,N_4234);
nand U4717 (N_4717,N_4240,N_4135);
or U4718 (N_4718,N_4072,N_4074);
or U4719 (N_4719,N_4133,N_4487);
or U4720 (N_4720,N_4238,N_4312);
nor U4721 (N_4721,N_4044,N_4376);
nor U4722 (N_4722,N_4089,N_4213);
nand U4723 (N_4723,N_4480,N_4208);
and U4724 (N_4724,N_4429,N_4303);
and U4725 (N_4725,N_4007,N_4361);
or U4726 (N_4726,N_4010,N_4088);
nand U4727 (N_4727,N_4350,N_4320);
or U4728 (N_4728,N_4377,N_4302);
or U4729 (N_4729,N_4155,N_4005);
or U4730 (N_4730,N_4223,N_4116);
or U4731 (N_4731,N_4309,N_4362);
nor U4732 (N_4732,N_4011,N_4284);
nor U4733 (N_4733,N_4100,N_4494);
nand U4734 (N_4734,N_4279,N_4337);
nor U4735 (N_4735,N_4375,N_4241);
nand U4736 (N_4736,N_4269,N_4293);
nor U4737 (N_4737,N_4287,N_4383);
nand U4738 (N_4738,N_4218,N_4235);
xor U4739 (N_4739,N_4198,N_4410);
nor U4740 (N_4740,N_4204,N_4316);
nor U4741 (N_4741,N_4327,N_4199);
nor U4742 (N_4742,N_4140,N_4448);
nand U4743 (N_4743,N_4071,N_4421);
or U4744 (N_4744,N_4188,N_4202);
nor U4745 (N_4745,N_4468,N_4138);
and U4746 (N_4746,N_4482,N_4397);
nand U4747 (N_4747,N_4321,N_4192);
nand U4748 (N_4748,N_4311,N_4085);
and U4749 (N_4749,N_4228,N_4270);
and U4750 (N_4750,N_4328,N_4290);
and U4751 (N_4751,N_4441,N_4244);
nor U4752 (N_4752,N_4084,N_4157);
and U4753 (N_4753,N_4112,N_4479);
or U4754 (N_4754,N_4295,N_4314);
nor U4755 (N_4755,N_4021,N_4425);
nand U4756 (N_4756,N_4264,N_4302);
nor U4757 (N_4757,N_4445,N_4163);
and U4758 (N_4758,N_4040,N_4415);
or U4759 (N_4759,N_4497,N_4126);
nand U4760 (N_4760,N_4458,N_4293);
nand U4761 (N_4761,N_4115,N_4032);
nand U4762 (N_4762,N_4483,N_4065);
nand U4763 (N_4763,N_4120,N_4236);
nor U4764 (N_4764,N_4439,N_4384);
nand U4765 (N_4765,N_4420,N_4476);
or U4766 (N_4766,N_4072,N_4254);
nand U4767 (N_4767,N_4248,N_4342);
and U4768 (N_4768,N_4065,N_4098);
xor U4769 (N_4769,N_4429,N_4445);
or U4770 (N_4770,N_4202,N_4360);
nor U4771 (N_4771,N_4298,N_4370);
nand U4772 (N_4772,N_4053,N_4039);
xor U4773 (N_4773,N_4277,N_4146);
nor U4774 (N_4774,N_4195,N_4425);
and U4775 (N_4775,N_4289,N_4385);
and U4776 (N_4776,N_4348,N_4044);
xnor U4777 (N_4777,N_4464,N_4466);
or U4778 (N_4778,N_4486,N_4079);
nand U4779 (N_4779,N_4145,N_4379);
and U4780 (N_4780,N_4497,N_4100);
nand U4781 (N_4781,N_4375,N_4430);
and U4782 (N_4782,N_4499,N_4001);
nand U4783 (N_4783,N_4415,N_4481);
nor U4784 (N_4784,N_4272,N_4379);
and U4785 (N_4785,N_4295,N_4470);
and U4786 (N_4786,N_4116,N_4137);
nor U4787 (N_4787,N_4311,N_4349);
or U4788 (N_4788,N_4314,N_4173);
or U4789 (N_4789,N_4227,N_4278);
xor U4790 (N_4790,N_4360,N_4273);
and U4791 (N_4791,N_4316,N_4215);
nand U4792 (N_4792,N_4484,N_4243);
nor U4793 (N_4793,N_4452,N_4322);
nor U4794 (N_4794,N_4410,N_4107);
nor U4795 (N_4795,N_4462,N_4084);
or U4796 (N_4796,N_4264,N_4281);
nor U4797 (N_4797,N_4396,N_4499);
nand U4798 (N_4798,N_4412,N_4233);
nand U4799 (N_4799,N_4377,N_4055);
and U4800 (N_4800,N_4450,N_4370);
and U4801 (N_4801,N_4006,N_4331);
nor U4802 (N_4802,N_4011,N_4414);
nand U4803 (N_4803,N_4330,N_4432);
nand U4804 (N_4804,N_4144,N_4361);
or U4805 (N_4805,N_4368,N_4146);
or U4806 (N_4806,N_4062,N_4303);
or U4807 (N_4807,N_4335,N_4348);
and U4808 (N_4808,N_4304,N_4264);
and U4809 (N_4809,N_4320,N_4396);
and U4810 (N_4810,N_4165,N_4043);
and U4811 (N_4811,N_4086,N_4215);
or U4812 (N_4812,N_4314,N_4326);
and U4813 (N_4813,N_4429,N_4423);
nor U4814 (N_4814,N_4474,N_4083);
or U4815 (N_4815,N_4132,N_4443);
nor U4816 (N_4816,N_4418,N_4370);
nor U4817 (N_4817,N_4174,N_4342);
nor U4818 (N_4818,N_4396,N_4344);
and U4819 (N_4819,N_4231,N_4126);
and U4820 (N_4820,N_4232,N_4011);
or U4821 (N_4821,N_4404,N_4420);
nand U4822 (N_4822,N_4123,N_4223);
and U4823 (N_4823,N_4217,N_4146);
nor U4824 (N_4824,N_4301,N_4112);
and U4825 (N_4825,N_4111,N_4099);
and U4826 (N_4826,N_4264,N_4405);
and U4827 (N_4827,N_4182,N_4051);
nor U4828 (N_4828,N_4277,N_4066);
and U4829 (N_4829,N_4173,N_4192);
and U4830 (N_4830,N_4287,N_4014);
and U4831 (N_4831,N_4388,N_4336);
nand U4832 (N_4832,N_4296,N_4093);
nor U4833 (N_4833,N_4419,N_4116);
nand U4834 (N_4834,N_4001,N_4243);
nand U4835 (N_4835,N_4134,N_4274);
or U4836 (N_4836,N_4185,N_4460);
or U4837 (N_4837,N_4155,N_4360);
and U4838 (N_4838,N_4417,N_4174);
or U4839 (N_4839,N_4358,N_4008);
and U4840 (N_4840,N_4041,N_4093);
or U4841 (N_4841,N_4063,N_4306);
and U4842 (N_4842,N_4176,N_4116);
and U4843 (N_4843,N_4119,N_4173);
and U4844 (N_4844,N_4482,N_4140);
nand U4845 (N_4845,N_4187,N_4330);
nand U4846 (N_4846,N_4208,N_4273);
or U4847 (N_4847,N_4257,N_4302);
nand U4848 (N_4848,N_4169,N_4046);
nand U4849 (N_4849,N_4436,N_4205);
or U4850 (N_4850,N_4187,N_4180);
or U4851 (N_4851,N_4178,N_4266);
nand U4852 (N_4852,N_4408,N_4220);
nor U4853 (N_4853,N_4495,N_4440);
or U4854 (N_4854,N_4273,N_4148);
and U4855 (N_4855,N_4056,N_4046);
and U4856 (N_4856,N_4156,N_4011);
nor U4857 (N_4857,N_4467,N_4342);
or U4858 (N_4858,N_4283,N_4236);
nand U4859 (N_4859,N_4334,N_4428);
and U4860 (N_4860,N_4402,N_4053);
and U4861 (N_4861,N_4408,N_4134);
or U4862 (N_4862,N_4297,N_4069);
nand U4863 (N_4863,N_4466,N_4256);
or U4864 (N_4864,N_4409,N_4195);
or U4865 (N_4865,N_4288,N_4094);
or U4866 (N_4866,N_4457,N_4013);
nand U4867 (N_4867,N_4060,N_4459);
or U4868 (N_4868,N_4009,N_4375);
and U4869 (N_4869,N_4470,N_4392);
and U4870 (N_4870,N_4256,N_4431);
or U4871 (N_4871,N_4097,N_4396);
or U4872 (N_4872,N_4231,N_4317);
and U4873 (N_4873,N_4423,N_4239);
or U4874 (N_4874,N_4316,N_4387);
nand U4875 (N_4875,N_4079,N_4065);
xor U4876 (N_4876,N_4371,N_4188);
nand U4877 (N_4877,N_4224,N_4183);
or U4878 (N_4878,N_4115,N_4367);
nand U4879 (N_4879,N_4405,N_4216);
nand U4880 (N_4880,N_4480,N_4162);
or U4881 (N_4881,N_4146,N_4358);
nor U4882 (N_4882,N_4128,N_4159);
nand U4883 (N_4883,N_4288,N_4356);
xnor U4884 (N_4884,N_4434,N_4385);
nand U4885 (N_4885,N_4315,N_4049);
and U4886 (N_4886,N_4400,N_4314);
and U4887 (N_4887,N_4440,N_4119);
nor U4888 (N_4888,N_4131,N_4121);
xor U4889 (N_4889,N_4260,N_4388);
and U4890 (N_4890,N_4092,N_4311);
xnor U4891 (N_4891,N_4000,N_4465);
nand U4892 (N_4892,N_4165,N_4480);
nand U4893 (N_4893,N_4088,N_4266);
nor U4894 (N_4894,N_4494,N_4475);
and U4895 (N_4895,N_4471,N_4026);
nand U4896 (N_4896,N_4118,N_4300);
nand U4897 (N_4897,N_4260,N_4076);
nor U4898 (N_4898,N_4308,N_4335);
nor U4899 (N_4899,N_4299,N_4473);
and U4900 (N_4900,N_4167,N_4199);
and U4901 (N_4901,N_4478,N_4197);
and U4902 (N_4902,N_4068,N_4497);
and U4903 (N_4903,N_4273,N_4249);
and U4904 (N_4904,N_4285,N_4369);
nand U4905 (N_4905,N_4418,N_4115);
nor U4906 (N_4906,N_4408,N_4474);
nand U4907 (N_4907,N_4317,N_4185);
and U4908 (N_4908,N_4206,N_4443);
nor U4909 (N_4909,N_4257,N_4389);
nor U4910 (N_4910,N_4117,N_4260);
nor U4911 (N_4911,N_4363,N_4071);
or U4912 (N_4912,N_4441,N_4352);
and U4913 (N_4913,N_4110,N_4169);
nor U4914 (N_4914,N_4372,N_4345);
nand U4915 (N_4915,N_4175,N_4078);
nor U4916 (N_4916,N_4005,N_4141);
xnor U4917 (N_4917,N_4326,N_4139);
nand U4918 (N_4918,N_4205,N_4433);
and U4919 (N_4919,N_4010,N_4265);
or U4920 (N_4920,N_4242,N_4317);
nor U4921 (N_4921,N_4336,N_4127);
or U4922 (N_4922,N_4334,N_4462);
nand U4923 (N_4923,N_4104,N_4091);
and U4924 (N_4924,N_4221,N_4285);
nor U4925 (N_4925,N_4365,N_4073);
or U4926 (N_4926,N_4206,N_4117);
or U4927 (N_4927,N_4132,N_4190);
or U4928 (N_4928,N_4309,N_4094);
or U4929 (N_4929,N_4070,N_4157);
nor U4930 (N_4930,N_4032,N_4336);
nand U4931 (N_4931,N_4455,N_4401);
xnor U4932 (N_4932,N_4161,N_4421);
nand U4933 (N_4933,N_4110,N_4172);
nor U4934 (N_4934,N_4409,N_4291);
and U4935 (N_4935,N_4080,N_4153);
nor U4936 (N_4936,N_4130,N_4217);
nor U4937 (N_4937,N_4389,N_4157);
nand U4938 (N_4938,N_4263,N_4341);
and U4939 (N_4939,N_4400,N_4388);
nor U4940 (N_4940,N_4298,N_4201);
nor U4941 (N_4941,N_4251,N_4150);
nor U4942 (N_4942,N_4175,N_4090);
or U4943 (N_4943,N_4282,N_4307);
or U4944 (N_4944,N_4461,N_4007);
nor U4945 (N_4945,N_4481,N_4190);
or U4946 (N_4946,N_4152,N_4085);
or U4947 (N_4947,N_4419,N_4428);
or U4948 (N_4948,N_4359,N_4321);
nand U4949 (N_4949,N_4343,N_4177);
nand U4950 (N_4950,N_4481,N_4273);
nand U4951 (N_4951,N_4143,N_4004);
nor U4952 (N_4952,N_4070,N_4093);
or U4953 (N_4953,N_4390,N_4163);
nand U4954 (N_4954,N_4194,N_4219);
nand U4955 (N_4955,N_4128,N_4409);
nor U4956 (N_4956,N_4407,N_4399);
nor U4957 (N_4957,N_4017,N_4327);
nand U4958 (N_4958,N_4316,N_4354);
and U4959 (N_4959,N_4424,N_4275);
or U4960 (N_4960,N_4036,N_4187);
or U4961 (N_4961,N_4471,N_4294);
nand U4962 (N_4962,N_4352,N_4080);
nor U4963 (N_4963,N_4151,N_4321);
nor U4964 (N_4964,N_4120,N_4441);
and U4965 (N_4965,N_4436,N_4471);
nand U4966 (N_4966,N_4273,N_4151);
and U4967 (N_4967,N_4338,N_4323);
or U4968 (N_4968,N_4338,N_4249);
or U4969 (N_4969,N_4496,N_4047);
and U4970 (N_4970,N_4329,N_4139);
or U4971 (N_4971,N_4094,N_4484);
nand U4972 (N_4972,N_4320,N_4028);
or U4973 (N_4973,N_4447,N_4169);
nand U4974 (N_4974,N_4259,N_4442);
nand U4975 (N_4975,N_4132,N_4268);
or U4976 (N_4976,N_4089,N_4498);
nor U4977 (N_4977,N_4270,N_4249);
xnor U4978 (N_4978,N_4164,N_4431);
nor U4979 (N_4979,N_4171,N_4240);
nand U4980 (N_4980,N_4400,N_4390);
nor U4981 (N_4981,N_4362,N_4445);
nor U4982 (N_4982,N_4484,N_4213);
or U4983 (N_4983,N_4093,N_4293);
and U4984 (N_4984,N_4049,N_4099);
nand U4985 (N_4985,N_4294,N_4137);
and U4986 (N_4986,N_4044,N_4041);
or U4987 (N_4987,N_4312,N_4440);
nor U4988 (N_4988,N_4451,N_4025);
and U4989 (N_4989,N_4107,N_4361);
or U4990 (N_4990,N_4294,N_4330);
nor U4991 (N_4991,N_4364,N_4162);
or U4992 (N_4992,N_4168,N_4377);
or U4993 (N_4993,N_4221,N_4230);
or U4994 (N_4994,N_4198,N_4190);
nor U4995 (N_4995,N_4352,N_4411);
nand U4996 (N_4996,N_4310,N_4196);
and U4997 (N_4997,N_4126,N_4227);
nand U4998 (N_4998,N_4226,N_4116);
nor U4999 (N_4999,N_4497,N_4026);
nor U5000 (N_5000,N_4884,N_4978);
or U5001 (N_5001,N_4612,N_4907);
nor U5002 (N_5002,N_4925,N_4609);
and U5003 (N_5003,N_4622,N_4506);
nand U5004 (N_5004,N_4672,N_4995);
and U5005 (N_5005,N_4673,N_4762);
and U5006 (N_5006,N_4620,N_4811);
or U5007 (N_5007,N_4727,N_4851);
nand U5008 (N_5008,N_4555,N_4946);
xnor U5009 (N_5009,N_4537,N_4550);
and U5010 (N_5010,N_4823,N_4618);
nor U5011 (N_5011,N_4879,N_4531);
nor U5012 (N_5012,N_4610,N_4633);
or U5013 (N_5013,N_4717,N_4522);
nor U5014 (N_5014,N_4999,N_4720);
and U5015 (N_5015,N_4819,N_4895);
nor U5016 (N_5016,N_4665,N_4986);
or U5017 (N_5017,N_4931,N_4745);
nand U5018 (N_5018,N_4586,N_4913);
nor U5019 (N_5019,N_4554,N_4509);
nor U5020 (N_5020,N_4645,N_4687);
nand U5021 (N_5021,N_4847,N_4683);
and U5022 (N_5022,N_4625,N_4602);
nor U5023 (N_5023,N_4575,N_4750);
nand U5024 (N_5024,N_4505,N_4979);
nor U5025 (N_5025,N_4841,N_4923);
nor U5026 (N_5026,N_4772,N_4974);
and U5027 (N_5027,N_4890,N_4523);
nor U5028 (N_5028,N_4903,N_4840);
nand U5029 (N_5029,N_4992,N_4648);
and U5030 (N_5030,N_4632,N_4716);
or U5031 (N_5031,N_4686,N_4810);
and U5032 (N_5032,N_4794,N_4713);
nand U5033 (N_5033,N_4773,N_4566);
or U5034 (N_5034,N_4545,N_4561);
nor U5035 (N_5035,N_4829,N_4926);
nor U5036 (N_5036,N_4538,N_4594);
nand U5037 (N_5037,N_4709,N_4831);
or U5038 (N_5038,N_4571,N_4953);
nor U5039 (N_5039,N_4621,N_4661);
xor U5040 (N_5040,N_4824,N_4919);
nor U5041 (N_5041,N_4732,N_4805);
nand U5042 (N_5042,N_4611,N_4998);
or U5043 (N_5043,N_4603,N_4968);
nor U5044 (N_5044,N_4941,N_4821);
nand U5045 (N_5045,N_4776,N_4500);
nor U5046 (N_5046,N_4548,N_4598);
or U5047 (N_5047,N_4796,N_4797);
or U5048 (N_5048,N_4886,N_4552);
nor U5049 (N_5049,N_4912,N_4910);
or U5050 (N_5050,N_4614,N_4589);
xnor U5051 (N_5051,N_4744,N_4534);
and U5052 (N_5052,N_4742,N_4736);
and U5053 (N_5053,N_4634,N_4551);
and U5054 (N_5054,N_4660,N_4905);
xnor U5055 (N_5055,N_4863,N_4993);
nor U5056 (N_5056,N_4607,N_4958);
nor U5057 (N_5057,N_4857,N_4578);
or U5058 (N_5058,N_4868,N_4597);
nor U5059 (N_5059,N_4615,N_4984);
or U5060 (N_5060,N_4936,N_4567);
or U5061 (N_5061,N_4767,N_4674);
nor U5062 (N_5062,N_4526,N_4825);
and U5063 (N_5063,N_4569,N_4681);
nand U5064 (N_5064,N_4543,N_4802);
nor U5065 (N_5065,N_4771,N_4558);
or U5066 (N_5066,N_4641,N_4664);
or U5067 (N_5067,N_4937,N_4954);
and U5068 (N_5068,N_4836,N_4737);
nor U5069 (N_5069,N_4966,N_4734);
nand U5070 (N_5070,N_4536,N_4549);
or U5071 (N_5071,N_4553,N_4828);
or U5072 (N_5072,N_4924,N_4718);
and U5073 (N_5073,N_4662,N_4693);
nand U5074 (N_5074,N_4647,N_4964);
or U5075 (N_5075,N_4535,N_4588);
or U5076 (N_5076,N_4761,N_4540);
or U5077 (N_5077,N_4635,N_4948);
or U5078 (N_5078,N_4712,N_4972);
nor U5079 (N_5079,N_4763,N_4636);
and U5080 (N_5080,N_4657,N_4581);
nor U5081 (N_5081,N_4908,N_4666);
or U5082 (N_5082,N_4568,N_4617);
nand U5083 (N_5083,N_4752,N_4976);
or U5084 (N_5084,N_4503,N_4897);
and U5085 (N_5085,N_4738,N_4596);
nand U5086 (N_5086,N_4853,N_4932);
xor U5087 (N_5087,N_4658,N_4803);
or U5088 (N_5088,N_4837,N_4669);
nand U5089 (N_5089,N_4985,N_4699);
nand U5090 (N_5090,N_4580,N_4870);
nand U5091 (N_5091,N_4730,N_4832);
nor U5092 (N_5092,N_4671,N_4963);
nor U5093 (N_5093,N_4756,N_4640);
nand U5094 (N_5094,N_4957,N_4677);
nor U5095 (N_5095,N_4875,N_4921);
nor U5096 (N_5096,N_4808,N_4547);
or U5097 (N_5097,N_4842,N_4934);
nor U5098 (N_5098,N_4511,N_4818);
and U5099 (N_5099,N_4945,N_4869);
nor U5100 (N_5100,N_4512,N_4876);
nor U5101 (N_5101,N_4758,N_4630);
nand U5102 (N_5102,N_4891,N_4601);
or U5103 (N_5103,N_4955,N_4753);
or U5104 (N_5104,N_4676,N_4795);
and U5105 (N_5105,N_4881,N_4711);
nand U5106 (N_5106,N_4817,N_4746);
nor U5107 (N_5107,N_4760,N_4639);
and U5108 (N_5108,N_4565,N_4965);
and U5109 (N_5109,N_4988,N_4827);
and U5110 (N_5110,N_4577,N_4951);
and U5111 (N_5111,N_4695,N_4502);
nand U5112 (N_5112,N_4694,N_4714);
nor U5113 (N_5113,N_4994,N_4651);
nor U5114 (N_5114,N_4864,N_4678);
and U5115 (N_5115,N_4990,N_4690);
nor U5116 (N_5116,N_4606,N_4781);
or U5117 (N_5117,N_4587,N_4906);
or U5118 (N_5118,N_4613,N_4754);
and U5119 (N_5119,N_4679,N_4521);
and U5120 (N_5120,N_4806,N_4708);
or U5121 (N_5121,N_4574,N_4838);
or U5122 (N_5122,N_4939,N_4515);
nor U5123 (N_5123,N_4680,N_4685);
or U5124 (N_5124,N_4975,N_4860);
nor U5125 (N_5125,N_4980,N_4922);
and U5126 (N_5126,N_4759,N_4780);
nand U5127 (N_5127,N_4570,N_4766);
nor U5128 (N_5128,N_4592,N_4843);
and U5129 (N_5129,N_4942,N_4705);
nand U5130 (N_5130,N_4917,N_4916);
xnor U5131 (N_5131,N_4777,N_4544);
and U5132 (N_5132,N_4816,N_4944);
or U5133 (N_5133,N_4724,N_4804);
and U5134 (N_5134,N_4629,N_4563);
and U5135 (N_5135,N_4790,N_4682);
nand U5136 (N_5136,N_4519,N_4774);
and U5137 (N_5137,N_4595,N_4967);
xor U5138 (N_5138,N_4987,N_4539);
nor U5139 (N_5139,N_4969,N_4542);
nor U5140 (N_5140,N_4728,N_4909);
or U5141 (N_5141,N_4848,N_4740);
and U5142 (N_5142,N_4960,N_4541);
nor U5143 (N_5143,N_4893,N_4862);
xor U5144 (N_5144,N_4751,N_4513);
nor U5145 (N_5145,N_4530,N_4726);
nor U5146 (N_5146,N_4582,N_4904);
nor U5147 (N_5147,N_4920,N_4982);
nor U5148 (N_5148,N_4562,N_4631);
nor U5149 (N_5149,N_4572,N_4835);
nor U5150 (N_5150,N_4775,N_4918);
nand U5151 (N_5151,N_4815,N_4623);
nand U5152 (N_5152,N_4779,N_4525);
nor U5153 (N_5153,N_4915,N_4956);
nor U5154 (N_5154,N_4989,N_4970);
or U5155 (N_5155,N_4556,N_4789);
nor U5156 (N_5156,N_4722,N_4559);
and U5157 (N_5157,N_4959,N_4719);
nor U5158 (N_5158,N_4793,N_4649);
or U5159 (N_5159,N_4809,N_4688);
or U5160 (N_5160,N_4943,N_4770);
xnor U5161 (N_5161,N_4834,N_4877);
nand U5162 (N_5162,N_4813,N_4782);
and U5163 (N_5163,N_4599,N_4533);
nand U5164 (N_5164,N_4739,N_4644);
or U5165 (N_5165,N_4675,N_4872);
nor U5166 (N_5166,N_4873,N_4799);
nand U5167 (N_5167,N_4757,N_4659);
or U5168 (N_5168,N_4784,N_4667);
nand U5169 (N_5169,N_4723,N_4604);
nand U5170 (N_5170,N_4684,N_4930);
xor U5171 (N_5171,N_4697,N_4791);
or U5172 (N_5172,N_4501,N_4590);
nand U5173 (N_5173,N_4997,N_4654);
nor U5174 (N_5174,N_4991,N_4643);
or U5175 (N_5175,N_4801,N_4689);
nor U5176 (N_5176,N_4899,N_4514);
nor U5177 (N_5177,N_4977,N_4844);
nor U5178 (N_5178,N_4755,N_4888);
and U5179 (N_5179,N_4783,N_4652);
nor U5180 (N_5180,N_4528,N_4961);
nand U5181 (N_5181,N_4894,N_4725);
and U5182 (N_5182,N_4619,N_4778);
or U5183 (N_5183,N_4769,N_4593);
nor U5184 (N_5184,N_4950,N_4787);
nor U5185 (N_5185,N_4764,N_4765);
or U5186 (N_5186,N_4933,N_4878);
nor U5187 (N_5187,N_4785,N_4792);
nor U5188 (N_5188,N_4655,N_4733);
or U5189 (N_5189,N_4715,N_4898);
nand U5190 (N_5190,N_4576,N_4929);
and U5191 (N_5191,N_4628,N_4928);
nor U5192 (N_5192,N_4646,N_4616);
nor U5193 (N_5193,N_4889,N_4874);
nor U5194 (N_5194,N_4650,N_4703);
nand U5195 (N_5195,N_4518,N_4527);
or U5196 (N_5196,N_4573,N_4627);
and U5197 (N_5197,N_4983,N_4871);
and U5198 (N_5198,N_4887,N_4900);
or U5199 (N_5199,N_4902,N_4663);
and U5200 (N_5200,N_4600,N_4626);
and U5201 (N_5201,N_4882,N_4704);
and U5202 (N_5202,N_4935,N_4798);
or U5203 (N_5203,N_4524,N_4911);
nand U5204 (N_5204,N_4865,N_4668);
nand U5205 (N_5205,N_4546,N_4856);
or U5206 (N_5206,N_4814,N_4845);
or U5207 (N_5207,N_4748,N_4642);
or U5208 (N_5208,N_4656,N_4585);
nand U5209 (N_5209,N_4880,N_4698);
nand U5210 (N_5210,N_4508,N_4885);
or U5211 (N_5211,N_4850,N_4517);
and U5212 (N_5212,N_4826,N_4892);
nor U5213 (N_5213,N_4608,N_4812);
nor U5214 (N_5214,N_4691,N_4854);
and U5215 (N_5215,N_4952,N_4516);
nand U5216 (N_5216,N_4624,N_4866);
and U5217 (N_5217,N_4706,N_4529);
or U5218 (N_5218,N_4996,N_4883);
and U5219 (N_5219,N_4507,N_4532);
and U5220 (N_5220,N_4949,N_4579);
or U5221 (N_5221,N_4867,N_4855);
and U5222 (N_5222,N_4820,N_4710);
nor U5223 (N_5223,N_4701,N_4981);
nor U5224 (N_5224,N_4735,N_4653);
nor U5225 (N_5225,N_4973,N_4788);
nor U5226 (N_5226,N_4914,N_4731);
or U5227 (N_5227,N_4510,N_4927);
nor U5228 (N_5228,N_4807,N_4938);
and U5229 (N_5229,N_4557,N_4741);
and U5230 (N_5230,N_4696,N_4591);
or U5231 (N_5231,N_4729,N_4833);
or U5232 (N_5232,N_4504,N_4822);
nand U5233 (N_5233,N_4859,N_4940);
and U5234 (N_5234,N_4849,N_4584);
or U5235 (N_5235,N_4670,N_4743);
or U5236 (N_5236,N_4721,N_4896);
nor U5237 (N_5237,N_4692,N_4638);
nand U5238 (N_5238,N_4861,N_4947);
nor U5239 (N_5239,N_4768,N_4962);
xor U5240 (N_5240,N_4707,N_4858);
and U5241 (N_5241,N_4800,N_4846);
nor U5242 (N_5242,N_4702,N_4971);
nor U5243 (N_5243,N_4852,N_4749);
nor U5244 (N_5244,N_4520,N_4901);
nand U5245 (N_5245,N_4605,N_4839);
or U5246 (N_5246,N_4564,N_4637);
nor U5247 (N_5247,N_4747,N_4700);
or U5248 (N_5248,N_4786,N_4560);
nor U5249 (N_5249,N_4583,N_4830);
or U5250 (N_5250,N_4927,N_4756);
nor U5251 (N_5251,N_4579,N_4644);
nand U5252 (N_5252,N_4775,N_4769);
or U5253 (N_5253,N_4684,N_4908);
nor U5254 (N_5254,N_4775,N_4637);
nand U5255 (N_5255,N_4912,N_4998);
and U5256 (N_5256,N_4603,N_4756);
or U5257 (N_5257,N_4940,N_4737);
or U5258 (N_5258,N_4824,N_4578);
or U5259 (N_5259,N_4878,N_4603);
nand U5260 (N_5260,N_4506,N_4891);
nand U5261 (N_5261,N_4969,N_4709);
xnor U5262 (N_5262,N_4668,N_4947);
nand U5263 (N_5263,N_4806,N_4807);
and U5264 (N_5264,N_4757,N_4640);
nor U5265 (N_5265,N_4628,N_4643);
and U5266 (N_5266,N_4505,N_4819);
or U5267 (N_5267,N_4767,N_4694);
nor U5268 (N_5268,N_4827,N_4726);
and U5269 (N_5269,N_4550,N_4528);
and U5270 (N_5270,N_4941,N_4900);
or U5271 (N_5271,N_4552,N_4969);
and U5272 (N_5272,N_4521,N_4590);
or U5273 (N_5273,N_4902,N_4559);
or U5274 (N_5274,N_4948,N_4693);
xnor U5275 (N_5275,N_4654,N_4855);
nor U5276 (N_5276,N_4628,N_4792);
or U5277 (N_5277,N_4791,N_4524);
nor U5278 (N_5278,N_4571,N_4585);
nor U5279 (N_5279,N_4872,N_4638);
or U5280 (N_5280,N_4666,N_4821);
and U5281 (N_5281,N_4968,N_4722);
or U5282 (N_5282,N_4759,N_4702);
nor U5283 (N_5283,N_4616,N_4887);
or U5284 (N_5284,N_4529,N_4992);
nor U5285 (N_5285,N_4729,N_4582);
and U5286 (N_5286,N_4883,N_4832);
nor U5287 (N_5287,N_4881,N_4972);
nand U5288 (N_5288,N_4714,N_4817);
nand U5289 (N_5289,N_4901,N_4922);
and U5290 (N_5290,N_4997,N_4826);
nand U5291 (N_5291,N_4670,N_4785);
nor U5292 (N_5292,N_4519,N_4920);
and U5293 (N_5293,N_4943,N_4896);
xor U5294 (N_5294,N_4816,N_4569);
or U5295 (N_5295,N_4859,N_4501);
nand U5296 (N_5296,N_4532,N_4803);
nand U5297 (N_5297,N_4921,N_4926);
and U5298 (N_5298,N_4916,N_4801);
or U5299 (N_5299,N_4990,N_4810);
nor U5300 (N_5300,N_4911,N_4518);
or U5301 (N_5301,N_4952,N_4858);
nor U5302 (N_5302,N_4527,N_4574);
or U5303 (N_5303,N_4672,N_4934);
and U5304 (N_5304,N_4709,N_4899);
nand U5305 (N_5305,N_4539,N_4841);
or U5306 (N_5306,N_4713,N_4961);
or U5307 (N_5307,N_4961,N_4856);
and U5308 (N_5308,N_4789,N_4719);
nor U5309 (N_5309,N_4948,N_4826);
nand U5310 (N_5310,N_4740,N_4701);
and U5311 (N_5311,N_4714,N_4930);
and U5312 (N_5312,N_4532,N_4920);
or U5313 (N_5313,N_4873,N_4679);
nand U5314 (N_5314,N_4787,N_4750);
nor U5315 (N_5315,N_4978,N_4826);
and U5316 (N_5316,N_4857,N_4635);
and U5317 (N_5317,N_4939,N_4938);
xnor U5318 (N_5318,N_4719,N_4685);
or U5319 (N_5319,N_4521,N_4953);
or U5320 (N_5320,N_4589,N_4504);
nor U5321 (N_5321,N_4973,N_4982);
nor U5322 (N_5322,N_4662,N_4801);
or U5323 (N_5323,N_4694,N_4814);
or U5324 (N_5324,N_4637,N_4576);
and U5325 (N_5325,N_4864,N_4943);
or U5326 (N_5326,N_4987,N_4686);
and U5327 (N_5327,N_4615,N_4953);
or U5328 (N_5328,N_4934,N_4965);
nand U5329 (N_5329,N_4568,N_4862);
nor U5330 (N_5330,N_4962,N_4798);
or U5331 (N_5331,N_4510,N_4991);
nor U5332 (N_5332,N_4547,N_4870);
xor U5333 (N_5333,N_4546,N_4592);
nand U5334 (N_5334,N_4580,N_4529);
nand U5335 (N_5335,N_4608,N_4671);
and U5336 (N_5336,N_4708,N_4610);
nand U5337 (N_5337,N_4683,N_4729);
and U5338 (N_5338,N_4796,N_4768);
xor U5339 (N_5339,N_4592,N_4616);
xor U5340 (N_5340,N_4915,N_4674);
and U5341 (N_5341,N_4508,N_4568);
xnor U5342 (N_5342,N_4985,N_4859);
nand U5343 (N_5343,N_4963,N_4827);
nor U5344 (N_5344,N_4658,N_4757);
nor U5345 (N_5345,N_4509,N_4815);
nand U5346 (N_5346,N_4693,N_4667);
and U5347 (N_5347,N_4709,N_4936);
nand U5348 (N_5348,N_4751,N_4974);
nand U5349 (N_5349,N_4731,N_4840);
nor U5350 (N_5350,N_4825,N_4634);
or U5351 (N_5351,N_4849,N_4506);
and U5352 (N_5352,N_4919,N_4964);
and U5353 (N_5353,N_4736,N_4549);
or U5354 (N_5354,N_4677,N_4627);
or U5355 (N_5355,N_4620,N_4861);
nor U5356 (N_5356,N_4505,N_4511);
nor U5357 (N_5357,N_4808,N_4527);
and U5358 (N_5358,N_4694,N_4873);
or U5359 (N_5359,N_4834,N_4538);
nor U5360 (N_5360,N_4779,N_4947);
and U5361 (N_5361,N_4910,N_4762);
nor U5362 (N_5362,N_4590,N_4586);
nand U5363 (N_5363,N_4829,N_4943);
or U5364 (N_5364,N_4622,N_4868);
nand U5365 (N_5365,N_4684,N_4816);
nor U5366 (N_5366,N_4606,N_4845);
nor U5367 (N_5367,N_4540,N_4644);
nand U5368 (N_5368,N_4698,N_4888);
and U5369 (N_5369,N_4949,N_4616);
nand U5370 (N_5370,N_4850,N_4838);
nand U5371 (N_5371,N_4793,N_4736);
and U5372 (N_5372,N_4825,N_4730);
nand U5373 (N_5373,N_4574,N_4795);
and U5374 (N_5374,N_4861,N_4740);
or U5375 (N_5375,N_4847,N_4909);
or U5376 (N_5376,N_4685,N_4614);
nor U5377 (N_5377,N_4840,N_4868);
and U5378 (N_5378,N_4686,N_4825);
nor U5379 (N_5379,N_4733,N_4626);
or U5380 (N_5380,N_4540,N_4993);
and U5381 (N_5381,N_4851,N_4983);
nor U5382 (N_5382,N_4577,N_4967);
and U5383 (N_5383,N_4925,N_4559);
nand U5384 (N_5384,N_4915,N_4823);
and U5385 (N_5385,N_4653,N_4828);
nand U5386 (N_5386,N_4882,N_4936);
and U5387 (N_5387,N_4747,N_4682);
nand U5388 (N_5388,N_4612,N_4717);
nor U5389 (N_5389,N_4725,N_4937);
and U5390 (N_5390,N_4894,N_4748);
nand U5391 (N_5391,N_4617,N_4779);
nor U5392 (N_5392,N_4734,N_4534);
and U5393 (N_5393,N_4864,N_4727);
and U5394 (N_5394,N_4604,N_4880);
and U5395 (N_5395,N_4589,N_4586);
or U5396 (N_5396,N_4681,N_4676);
nand U5397 (N_5397,N_4927,N_4798);
or U5398 (N_5398,N_4730,N_4713);
and U5399 (N_5399,N_4943,N_4752);
nand U5400 (N_5400,N_4931,N_4922);
nor U5401 (N_5401,N_4896,N_4668);
and U5402 (N_5402,N_4574,N_4531);
nand U5403 (N_5403,N_4522,N_4610);
and U5404 (N_5404,N_4921,N_4646);
or U5405 (N_5405,N_4634,N_4860);
xor U5406 (N_5406,N_4958,N_4904);
nand U5407 (N_5407,N_4850,N_4786);
nor U5408 (N_5408,N_4945,N_4516);
nor U5409 (N_5409,N_4722,N_4771);
and U5410 (N_5410,N_4768,N_4638);
nand U5411 (N_5411,N_4954,N_4628);
nand U5412 (N_5412,N_4783,N_4974);
nor U5413 (N_5413,N_4696,N_4649);
and U5414 (N_5414,N_4822,N_4850);
nand U5415 (N_5415,N_4692,N_4574);
nand U5416 (N_5416,N_4925,N_4753);
nand U5417 (N_5417,N_4935,N_4881);
nand U5418 (N_5418,N_4910,N_4649);
nand U5419 (N_5419,N_4506,N_4862);
and U5420 (N_5420,N_4523,N_4849);
nor U5421 (N_5421,N_4515,N_4788);
nor U5422 (N_5422,N_4686,N_4719);
or U5423 (N_5423,N_4900,N_4621);
and U5424 (N_5424,N_4977,N_4950);
or U5425 (N_5425,N_4598,N_4793);
or U5426 (N_5426,N_4619,N_4639);
nor U5427 (N_5427,N_4567,N_4796);
and U5428 (N_5428,N_4944,N_4858);
or U5429 (N_5429,N_4546,N_4707);
nand U5430 (N_5430,N_4638,N_4511);
and U5431 (N_5431,N_4504,N_4979);
nor U5432 (N_5432,N_4534,N_4759);
nor U5433 (N_5433,N_4866,N_4570);
and U5434 (N_5434,N_4860,N_4759);
and U5435 (N_5435,N_4708,N_4583);
nor U5436 (N_5436,N_4864,N_4926);
or U5437 (N_5437,N_4863,N_4529);
and U5438 (N_5438,N_4507,N_4862);
and U5439 (N_5439,N_4645,N_4621);
or U5440 (N_5440,N_4974,N_4679);
nand U5441 (N_5441,N_4802,N_4997);
and U5442 (N_5442,N_4688,N_4516);
and U5443 (N_5443,N_4749,N_4667);
or U5444 (N_5444,N_4514,N_4675);
and U5445 (N_5445,N_4763,N_4539);
nor U5446 (N_5446,N_4868,N_4586);
nor U5447 (N_5447,N_4777,N_4690);
nor U5448 (N_5448,N_4547,N_4566);
and U5449 (N_5449,N_4626,N_4916);
and U5450 (N_5450,N_4804,N_4684);
and U5451 (N_5451,N_4753,N_4841);
or U5452 (N_5452,N_4654,N_4830);
nor U5453 (N_5453,N_4742,N_4579);
and U5454 (N_5454,N_4880,N_4941);
nor U5455 (N_5455,N_4618,N_4541);
nor U5456 (N_5456,N_4616,N_4510);
nor U5457 (N_5457,N_4594,N_4845);
or U5458 (N_5458,N_4531,N_4655);
or U5459 (N_5459,N_4640,N_4625);
nand U5460 (N_5460,N_4965,N_4513);
nor U5461 (N_5461,N_4895,N_4748);
nand U5462 (N_5462,N_4603,N_4895);
xnor U5463 (N_5463,N_4964,N_4888);
and U5464 (N_5464,N_4904,N_4673);
or U5465 (N_5465,N_4516,N_4909);
nor U5466 (N_5466,N_4563,N_4929);
or U5467 (N_5467,N_4980,N_4628);
nand U5468 (N_5468,N_4682,N_4608);
and U5469 (N_5469,N_4662,N_4672);
nor U5470 (N_5470,N_4919,N_4565);
and U5471 (N_5471,N_4617,N_4923);
or U5472 (N_5472,N_4941,N_4849);
xnor U5473 (N_5473,N_4984,N_4838);
and U5474 (N_5474,N_4546,N_4502);
and U5475 (N_5475,N_4864,N_4692);
nor U5476 (N_5476,N_4540,N_4739);
nand U5477 (N_5477,N_4663,N_4696);
nor U5478 (N_5478,N_4654,N_4517);
nor U5479 (N_5479,N_4597,N_4885);
nand U5480 (N_5480,N_4634,N_4609);
or U5481 (N_5481,N_4891,N_4761);
xor U5482 (N_5482,N_4945,N_4865);
or U5483 (N_5483,N_4647,N_4636);
or U5484 (N_5484,N_4535,N_4953);
and U5485 (N_5485,N_4512,N_4786);
nor U5486 (N_5486,N_4988,N_4595);
nand U5487 (N_5487,N_4792,N_4903);
nand U5488 (N_5488,N_4866,N_4595);
nor U5489 (N_5489,N_4752,N_4817);
or U5490 (N_5490,N_4562,N_4768);
nand U5491 (N_5491,N_4546,N_4684);
or U5492 (N_5492,N_4709,N_4663);
and U5493 (N_5493,N_4932,N_4858);
or U5494 (N_5494,N_4938,N_4532);
nor U5495 (N_5495,N_4934,N_4684);
and U5496 (N_5496,N_4969,N_4730);
nand U5497 (N_5497,N_4889,N_4558);
nor U5498 (N_5498,N_4785,N_4860);
or U5499 (N_5499,N_4733,N_4729);
or U5500 (N_5500,N_5023,N_5164);
xor U5501 (N_5501,N_5087,N_5357);
and U5502 (N_5502,N_5011,N_5340);
nand U5503 (N_5503,N_5461,N_5373);
or U5504 (N_5504,N_5449,N_5344);
and U5505 (N_5505,N_5096,N_5367);
nor U5506 (N_5506,N_5138,N_5429);
or U5507 (N_5507,N_5418,N_5471);
or U5508 (N_5508,N_5388,N_5292);
and U5509 (N_5509,N_5168,N_5133);
or U5510 (N_5510,N_5310,N_5350);
or U5511 (N_5511,N_5103,N_5285);
nand U5512 (N_5512,N_5099,N_5142);
nand U5513 (N_5513,N_5490,N_5060);
or U5514 (N_5514,N_5097,N_5448);
nor U5515 (N_5515,N_5355,N_5360);
or U5516 (N_5516,N_5474,N_5270);
and U5517 (N_5517,N_5054,N_5433);
or U5518 (N_5518,N_5372,N_5196);
nor U5519 (N_5519,N_5309,N_5296);
nand U5520 (N_5520,N_5002,N_5352);
and U5521 (N_5521,N_5324,N_5409);
or U5522 (N_5522,N_5226,N_5191);
nand U5523 (N_5523,N_5294,N_5293);
nor U5524 (N_5524,N_5404,N_5442);
and U5525 (N_5525,N_5361,N_5231);
nor U5526 (N_5526,N_5493,N_5106);
xor U5527 (N_5527,N_5094,N_5325);
nand U5528 (N_5528,N_5035,N_5271);
or U5529 (N_5529,N_5261,N_5411);
and U5530 (N_5530,N_5434,N_5304);
nor U5531 (N_5531,N_5439,N_5064);
nor U5532 (N_5532,N_5412,N_5414);
nor U5533 (N_5533,N_5489,N_5326);
or U5534 (N_5534,N_5472,N_5484);
nor U5535 (N_5535,N_5247,N_5118);
nand U5536 (N_5536,N_5494,N_5179);
nand U5537 (N_5537,N_5151,N_5263);
or U5538 (N_5538,N_5214,N_5051);
or U5539 (N_5539,N_5464,N_5177);
or U5540 (N_5540,N_5420,N_5199);
xor U5541 (N_5541,N_5216,N_5445);
nand U5542 (N_5542,N_5217,N_5430);
nor U5543 (N_5543,N_5190,N_5431);
nor U5544 (N_5544,N_5030,N_5497);
or U5545 (N_5545,N_5347,N_5380);
xnor U5546 (N_5546,N_5395,N_5295);
nand U5547 (N_5547,N_5148,N_5056);
nand U5548 (N_5548,N_5165,N_5137);
or U5549 (N_5549,N_5026,N_5045);
and U5550 (N_5550,N_5432,N_5245);
nand U5551 (N_5551,N_5072,N_5341);
and U5552 (N_5552,N_5470,N_5486);
nand U5553 (N_5553,N_5088,N_5032);
nand U5554 (N_5554,N_5206,N_5419);
nand U5555 (N_5555,N_5331,N_5275);
nand U5556 (N_5556,N_5237,N_5076);
nor U5557 (N_5557,N_5382,N_5255);
and U5558 (N_5558,N_5368,N_5406);
and U5559 (N_5559,N_5371,N_5264);
or U5560 (N_5560,N_5182,N_5273);
and U5561 (N_5561,N_5068,N_5391);
and U5562 (N_5562,N_5480,N_5028);
nand U5563 (N_5563,N_5147,N_5450);
or U5564 (N_5564,N_5102,N_5329);
nand U5565 (N_5565,N_5353,N_5443);
nor U5566 (N_5566,N_5456,N_5074);
or U5567 (N_5567,N_5128,N_5356);
nor U5568 (N_5568,N_5283,N_5145);
nand U5569 (N_5569,N_5407,N_5254);
nor U5570 (N_5570,N_5093,N_5223);
or U5571 (N_5571,N_5375,N_5234);
nor U5572 (N_5572,N_5277,N_5062);
nor U5573 (N_5573,N_5159,N_5415);
nand U5574 (N_5574,N_5278,N_5120);
nand U5575 (N_5575,N_5017,N_5410);
and U5576 (N_5576,N_5211,N_5012);
nand U5577 (N_5577,N_5210,N_5390);
nand U5578 (N_5578,N_5114,N_5004);
or U5579 (N_5579,N_5057,N_5466);
nor U5580 (N_5580,N_5303,N_5117);
nand U5581 (N_5581,N_5243,N_5020);
nor U5582 (N_5582,N_5171,N_5042);
nand U5583 (N_5583,N_5343,N_5333);
nand U5584 (N_5584,N_5156,N_5022);
nor U5585 (N_5585,N_5167,N_5485);
nand U5586 (N_5586,N_5358,N_5116);
nor U5587 (N_5587,N_5280,N_5473);
or U5588 (N_5588,N_5065,N_5379);
and U5589 (N_5589,N_5043,N_5351);
and U5590 (N_5590,N_5413,N_5027);
nor U5591 (N_5591,N_5173,N_5198);
and U5592 (N_5592,N_5104,N_5157);
nand U5593 (N_5593,N_5069,N_5495);
or U5594 (N_5594,N_5149,N_5183);
and U5595 (N_5595,N_5327,N_5359);
or U5596 (N_5596,N_5208,N_5115);
nor U5597 (N_5597,N_5284,N_5058);
nor U5598 (N_5598,N_5084,N_5427);
and U5599 (N_5599,N_5140,N_5090);
nor U5600 (N_5600,N_5291,N_5031);
and U5601 (N_5601,N_5338,N_5385);
nand U5602 (N_5602,N_5161,N_5394);
nand U5603 (N_5603,N_5186,N_5135);
xor U5604 (N_5604,N_5328,N_5007);
nor U5605 (N_5605,N_5101,N_5483);
or U5606 (N_5606,N_5317,N_5405);
nand U5607 (N_5607,N_5377,N_5459);
nand U5608 (N_5608,N_5453,N_5279);
or U5609 (N_5609,N_5203,N_5089);
nor U5610 (N_5610,N_5207,N_5320);
and U5611 (N_5611,N_5256,N_5123);
nand U5612 (N_5612,N_5276,N_5300);
and U5613 (N_5613,N_5050,N_5111);
or U5614 (N_5614,N_5193,N_5386);
xnor U5615 (N_5615,N_5000,N_5136);
nand U5616 (N_5616,N_5224,N_5083);
and U5617 (N_5617,N_5323,N_5348);
nand U5618 (N_5618,N_5187,N_5313);
and U5619 (N_5619,N_5399,N_5169);
and U5620 (N_5620,N_5428,N_5205);
nor U5621 (N_5621,N_5318,N_5469);
nand U5622 (N_5622,N_5113,N_5397);
nand U5623 (N_5623,N_5143,N_5176);
nand U5624 (N_5624,N_5152,N_5122);
and U5625 (N_5625,N_5478,N_5053);
and U5626 (N_5626,N_5481,N_5003);
nand U5627 (N_5627,N_5458,N_5455);
nor U5628 (N_5628,N_5095,N_5364);
nor U5629 (N_5629,N_5334,N_5086);
nor U5630 (N_5630,N_5110,N_5370);
and U5631 (N_5631,N_5457,N_5381);
nor U5632 (N_5632,N_5289,N_5259);
nor U5633 (N_5633,N_5024,N_5238);
and U5634 (N_5634,N_5437,N_5048);
nand U5635 (N_5635,N_5257,N_5034);
and U5636 (N_5636,N_5127,N_5105);
or U5637 (N_5637,N_5307,N_5218);
or U5638 (N_5638,N_5366,N_5121);
nor U5639 (N_5639,N_5041,N_5475);
nand U5640 (N_5640,N_5479,N_5321);
or U5641 (N_5641,N_5188,N_5498);
and U5642 (N_5642,N_5487,N_5209);
or U5643 (N_5643,N_5384,N_5311);
xnor U5644 (N_5644,N_5269,N_5134);
nor U5645 (N_5645,N_5287,N_5194);
nor U5646 (N_5646,N_5244,N_5383);
nor U5647 (N_5647,N_5055,N_5202);
nand U5648 (N_5648,N_5335,N_5175);
and U5649 (N_5649,N_5204,N_5248);
nand U5650 (N_5650,N_5233,N_5345);
and U5651 (N_5651,N_5158,N_5192);
nor U5652 (N_5652,N_5378,N_5346);
and U5653 (N_5653,N_5339,N_5132);
nand U5654 (N_5654,N_5236,N_5258);
and U5655 (N_5655,N_5402,N_5421);
nor U5656 (N_5656,N_5129,N_5316);
or U5657 (N_5657,N_5005,N_5290);
or U5658 (N_5658,N_5221,N_5220);
nor U5659 (N_5659,N_5178,N_5301);
or U5660 (N_5660,N_5477,N_5195);
nand U5661 (N_5661,N_5049,N_5067);
and U5662 (N_5662,N_5080,N_5229);
or U5663 (N_5663,N_5125,N_5160);
and U5664 (N_5664,N_5297,N_5426);
nand U5665 (N_5665,N_5365,N_5451);
nand U5666 (N_5666,N_5249,N_5213);
nor U5667 (N_5667,N_5354,N_5150);
and U5668 (N_5668,N_5073,N_5337);
nor U5669 (N_5669,N_5107,N_5197);
nor U5670 (N_5670,N_5059,N_5006);
or U5671 (N_5671,N_5319,N_5025);
nor U5672 (N_5672,N_5462,N_5201);
nand U5673 (N_5673,N_5302,N_5298);
nand U5674 (N_5674,N_5219,N_5342);
nor U5675 (N_5675,N_5392,N_5139);
or U5676 (N_5676,N_5369,N_5100);
nand U5677 (N_5677,N_5240,N_5322);
nand U5678 (N_5678,N_5438,N_5314);
and U5679 (N_5679,N_5460,N_5166);
and U5680 (N_5680,N_5305,N_5425);
and U5681 (N_5681,N_5423,N_5330);
nor U5682 (N_5682,N_5288,N_5155);
and U5683 (N_5683,N_5075,N_5008);
nand U5684 (N_5684,N_5315,N_5131);
nand U5685 (N_5685,N_5267,N_5436);
and U5686 (N_5686,N_5447,N_5010);
or U5687 (N_5687,N_5435,N_5282);
or U5688 (N_5688,N_5441,N_5476);
nand U5689 (N_5689,N_5146,N_5189);
and U5690 (N_5690,N_5374,N_5061);
or U5691 (N_5691,N_5252,N_5130);
or U5692 (N_5692,N_5225,N_5266);
xor U5693 (N_5693,N_5047,N_5037);
nor U5694 (N_5694,N_5440,N_5184);
or U5695 (N_5695,N_5424,N_5235);
nand U5696 (N_5696,N_5021,N_5492);
nand U5697 (N_5697,N_5014,N_5185);
or U5698 (N_5698,N_5268,N_5013);
and U5699 (N_5699,N_5401,N_5299);
nand U5700 (N_5700,N_5082,N_5417);
xor U5701 (N_5701,N_5400,N_5044);
and U5702 (N_5702,N_5009,N_5126);
xor U5703 (N_5703,N_5239,N_5215);
and U5704 (N_5704,N_5071,N_5227);
xnor U5705 (N_5705,N_5468,N_5141);
nor U5706 (N_5706,N_5467,N_5077);
and U5707 (N_5707,N_5001,N_5163);
nand U5708 (N_5708,N_5029,N_5272);
nand U5709 (N_5709,N_5260,N_5228);
nor U5710 (N_5710,N_5066,N_5091);
or U5711 (N_5711,N_5422,N_5242);
and U5712 (N_5712,N_5144,N_5124);
nor U5713 (N_5713,N_5444,N_5262);
and U5714 (N_5714,N_5416,N_5482);
nand U5715 (N_5715,N_5019,N_5396);
and U5716 (N_5716,N_5172,N_5222);
nand U5717 (N_5717,N_5200,N_5253);
nand U5718 (N_5718,N_5387,N_5408);
and U5719 (N_5719,N_5376,N_5403);
and U5720 (N_5720,N_5119,N_5286);
or U5721 (N_5721,N_5241,N_5363);
and U5722 (N_5722,N_5308,N_5362);
or U5723 (N_5723,N_5306,N_5463);
and U5724 (N_5724,N_5108,N_5349);
or U5725 (N_5725,N_5081,N_5499);
or U5726 (N_5726,N_5251,N_5070);
or U5727 (N_5727,N_5465,N_5312);
nor U5728 (N_5728,N_5246,N_5446);
and U5729 (N_5729,N_5018,N_5109);
nor U5730 (N_5730,N_5038,N_5265);
and U5731 (N_5731,N_5332,N_5230);
nor U5732 (N_5732,N_5232,N_5063);
and U5733 (N_5733,N_5488,N_5274);
nand U5734 (N_5734,N_5212,N_5078);
and U5735 (N_5735,N_5154,N_5281);
nand U5736 (N_5736,N_5336,N_5181);
nand U5737 (N_5737,N_5085,N_5098);
nand U5738 (N_5738,N_5393,N_5454);
and U5739 (N_5739,N_5162,N_5036);
nand U5740 (N_5740,N_5180,N_5039);
and U5741 (N_5741,N_5452,N_5079);
and U5742 (N_5742,N_5491,N_5496);
nand U5743 (N_5743,N_5398,N_5016);
or U5744 (N_5744,N_5092,N_5040);
and U5745 (N_5745,N_5052,N_5112);
or U5746 (N_5746,N_5174,N_5250);
or U5747 (N_5747,N_5389,N_5033);
and U5748 (N_5748,N_5170,N_5015);
and U5749 (N_5749,N_5153,N_5046);
nor U5750 (N_5750,N_5427,N_5015);
or U5751 (N_5751,N_5071,N_5356);
nor U5752 (N_5752,N_5298,N_5177);
nor U5753 (N_5753,N_5434,N_5324);
or U5754 (N_5754,N_5003,N_5075);
nor U5755 (N_5755,N_5046,N_5461);
or U5756 (N_5756,N_5398,N_5437);
nand U5757 (N_5757,N_5302,N_5067);
or U5758 (N_5758,N_5058,N_5154);
or U5759 (N_5759,N_5119,N_5479);
or U5760 (N_5760,N_5153,N_5165);
or U5761 (N_5761,N_5010,N_5036);
and U5762 (N_5762,N_5118,N_5234);
nor U5763 (N_5763,N_5299,N_5082);
nor U5764 (N_5764,N_5254,N_5466);
or U5765 (N_5765,N_5397,N_5450);
or U5766 (N_5766,N_5085,N_5031);
and U5767 (N_5767,N_5403,N_5056);
and U5768 (N_5768,N_5382,N_5247);
nand U5769 (N_5769,N_5215,N_5086);
and U5770 (N_5770,N_5006,N_5002);
and U5771 (N_5771,N_5337,N_5305);
or U5772 (N_5772,N_5430,N_5426);
and U5773 (N_5773,N_5348,N_5445);
or U5774 (N_5774,N_5173,N_5133);
nand U5775 (N_5775,N_5345,N_5450);
and U5776 (N_5776,N_5073,N_5022);
nand U5777 (N_5777,N_5088,N_5427);
nor U5778 (N_5778,N_5015,N_5047);
nor U5779 (N_5779,N_5084,N_5244);
xnor U5780 (N_5780,N_5320,N_5165);
nand U5781 (N_5781,N_5324,N_5018);
or U5782 (N_5782,N_5371,N_5405);
nor U5783 (N_5783,N_5080,N_5072);
or U5784 (N_5784,N_5237,N_5100);
nand U5785 (N_5785,N_5033,N_5199);
nor U5786 (N_5786,N_5436,N_5035);
and U5787 (N_5787,N_5063,N_5387);
and U5788 (N_5788,N_5148,N_5114);
nor U5789 (N_5789,N_5329,N_5397);
nor U5790 (N_5790,N_5286,N_5199);
or U5791 (N_5791,N_5488,N_5027);
nand U5792 (N_5792,N_5017,N_5349);
nand U5793 (N_5793,N_5295,N_5028);
and U5794 (N_5794,N_5259,N_5231);
or U5795 (N_5795,N_5200,N_5360);
and U5796 (N_5796,N_5204,N_5294);
and U5797 (N_5797,N_5380,N_5092);
nand U5798 (N_5798,N_5399,N_5167);
nand U5799 (N_5799,N_5354,N_5021);
nor U5800 (N_5800,N_5399,N_5490);
xor U5801 (N_5801,N_5189,N_5293);
nor U5802 (N_5802,N_5427,N_5356);
nand U5803 (N_5803,N_5037,N_5288);
nor U5804 (N_5804,N_5216,N_5386);
and U5805 (N_5805,N_5430,N_5369);
nand U5806 (N_5806,N_5254,N_5474);
or U5807 (N_5807,N_5224,N_5013);
or U5808 (N_5808,N_5035,N_5126);
nor U5809 (N_5809,N_5490,N_5104);
nand U5810 (N_5810,N_5239,N_5218);
and U5811 (N_5811,N_5062,N_5217);
nand U5812 (N_5812,N_5456,N_5421);
xor U5813 (N_5813,N_5395,N_5001);
nand U5814 (N_5814,N_5404,N_5224);
nand U5815 (N_5815,N_5121,N_5081);
nand U5816 (N_5816,N_5121,N_5184);
nand U5817 (N_5817,N_5273,N_5069);
nor U5818 (N_5818,N_5207,N_5424);
or U5819 (N_5819,N_5367,N_5181);
nand U5820 (N_5820,N_5357,N_5319);
or U5821 (N_5821,N_5105,N_5057);
or U5822 (N_5822,N_5369,N_5424);
nor U5823 (N_5823,N_5044,N_5017);
and U5824 (N_5824,N_5494,N_5068);
nand U5825 (N_5825,N_5297,N_5348);
nor U5826 (N_5826,N_5413,N_5016);
nand U5827 (N_5827,N_5113,N_5481);
nor U5828 (N_5828,N_5357,N_5025);
and U5829 (N_5829,N_5011,N_5188);
and U5830 (N_5830,N_5234,N_5185);
and U5831 (N_5831,N_5348,N_5061);
nand U5832 (N_5832,N_5045,N_5030);
or U5833 (N_5833,N_5377,N_5123);
nor U5834 (N_5834,N_5128,N_5049);
nand U5835 (N_5835,N_5017,N_5446);
nor U5836 (N_5836,N_5128,N_5423);
or U5837 (N_5837,N_5225,N_5150);
and U5838 (N_5838,N_5308,N_5327);
nor U5839 (N_5839,N_5301,N_5188);
and U5840 (N_5840,N_5022,N_5368);
or U5841 (N_5841,N_5216,N_5181);
nor U5842 (N_5842,N_5370,N_5430);
nor U5843 (N_5843,N_5475,N_5130);
nand U5844 (N_5844,N_5421,N_5330);
and U5845 (N_5845,N_5106,N_5367);
nand U5846 (N_5846,N_5274,N_5399);
and U5847 (N_5847,N_5171,N_5453);
nor U5848 (N_5848,N_5493,N_5224);
nor U5849 (N_5849,N_5488,N_5071);
and U5850 (N_5850,N_5467,N_5333);
xnor U5851 (N_5851,N_5057,N_5346);
nor U5852 (N_5852,N_5498,N_5108);
or U5853 (N_5853,N_5073,N_5279);
nor U5854 (N_5854,N_5077,N_5021);
and U5855 (N_5855,N_5038,N_5169);
nand U5856 (N_5856,N_5354,N_5096);
xor U5857 (N_5857,N_5255,N_5337);
nand U5858 (N_5858,N_5351,N_5445);
and U5859 (N_5859,N_5115,N_5307);
and U5860 (N_5860,N_5496,N_5492);
nor U5861 (N_5861,N_5136,N_5070);
nor U5862 (N_5862,N_5182,N_5257);
and U5863 (N_5863,N_5039,N_5085);
or U5864 (N_5864,N_5151,N_5413);
nand U5865 (N_5865,N_5052,N_5072);
and U5866 (N_5866,N_5224,N_5069);
nor U5867 (N_5867,N_5216,N_5074);
and U5868 (N_5868,N_5402,N_5429);
or U5869 (N_5869,N_5121,N_5229);
xnor U5870 (N_5870,N_5094,N_5413);
or U5871 (N_5871,N_5441,N_5310);
nor U5872 (N_5872,N_5015,N_5155);
and U5873 (N_5873,N_5364,N_5326);
and U5874 (N_5874,N_5156,N_5241);
nor U5875 (N_5875,N_5393,N_5320);
nor U5876 (N_5876,N_5429,N_5411);
or U5877 (N_5877,N_5457,N_5068);
nand U5878 (N_5878,N_5095,N_5497);
and U5879 (N_5879,N_5233,N_5203);
or U5880 (N_5880,N_5214,N_5477);
and U5881 (N_5881,N_5444,N_5195);
nand U5882 (N_5882,N_5292,N_5027);
or U5883 (N_5883,N_5448,N_5304);
and U5884 (N_5884,N_5496,N_5371);
and U5885 (N_5885,N_5399,N_5057);
or U5886 (N_5886,N_5487,N_5403);
nor U5887 (N_5887,N_5264,N_5328);
or U5888 (N_5888,N_5165,N_5389);
nor U5889 (N_5889,N_5423,N_5296);
or U5890 (N_5890,N_5283,N_5471);
and U5891 (N_5891,N_5281,N_5460);
or U5892 (N_5892,N_5440,N_5289);
nor U5893 (N_5893,N_5428,N_5254);
and U5894 (N_5894,N_5253,N_5172);
nand U5895 (N_5895,N_5008,N_5382);
nand U5896 (N_5896,N_5192,N_5313);
or U5897 (N_5897,N_5157,N_5298);
or U5898 (N_5898,N_5135,N_5499);
nor U5899 (N_5899,N_5026,N_5450);
nor U5900 (N_5900,N_5308,N_5054);
nand U5901 (N_5901,N_5238,N_5284);
nor U5902 (N_5902,N_5214,N_5441);
nand U5903 (N_5903,N_5300,N_5466);
nor U5904 (N_5904,N_5494,N_5357);
and U5905 (N_5905,N_5015,N_5368);
nor U5906 (N_5906,N_5442,N_5366);
or U5907 (N_5907,N_5266,N_5343);
nor U5908 (N_5908,N_5318,N_5286);
nand U5909 (N_5909,N_5047,N_5390);
nand U5910 (N_5910,N_5308,N_5067);
and U5911 (N_5911,N_5263,N_5071);
or U5912 (N_5912,N_5220,N_5093);
and U5913 (N_5913,N_5208,N_5149);
nand U5914 (N_5914,N_5231,N_5098);
nor U5915 (N_5915,N_5470,N_5218);
xor U5916 (N_5916,N_5161,N_5254);
nor U5917 (N_5917,N_5364,N_5139);
nor U5918 (N_5918,N_5401,N_5415);
or U5919 (N_5919,N_5418,N_5395);
or U5920 (N_5920,N_5318,N_5197);
nor U5921 (N_5921,N_5376,N_5395);
or U5922 (N_5922,N_5197,N_5037);
nor U5923 (N_5923,N_5136,N_5175);
nand U5924 (N_5924,N_5341,N_5248);
nor U5925 (N_5925,N_5411,N_5435);
nor U5926 (N_5926,N_5048,N_5391);
or U5927 (N_5927,N_5008,N_5307);
and U5928 (N_5928,N_5197,N_5206);
nor U5929 (N_5929,N_5413,N_5120);
or U5930 (N_5930,N_5028,N_5018);
nand U5931 (N_5931,N_5338,N_5256);
nand U5932 (N_5932,N_5389,N_5370);
nor U5933 (N_5933,N_5049,N_5437);
and U5934 (N_5934,N_5204,N_5038);
or U5935 (N_5935,N_5392,N_5218);
and U5936 (N_5936,N_5018,N_5368);
or U5937 (N_5937,N_5032,N_5492);
and U5938 (N_5938,N_5240,N_5022);
or U5939 (N_5939,N_5290,N_5131);
nor U5940 (N_5940,N_5235,N_5213);
or U5941 (N_5941,N_5397,N_5194);
nor U5942 (N_5942,N_5152,N_5446);
or U5943 (N_5943,N_5247,N_5047);
nand U5944 (N_5944,N_5238,N_5360);
and U5945 (N_5945,N_5449,N_5351);
or U5946 (N_5946,N_5465,N_5068);
nand U5947 (N_5947,N_5212,N_5477);
or U5948 (N_5948,N_5087,N_5323);
nor U5949 (N_5949,N_5087,N_5416);
nor U5950 (N_5950,N_5247,N_5136);
nand U5951 (N_5951,N_5189,N_5367);
nand U5952 (N_5952,N_5162,N_5014);
and U5953 (N_5953,N_5022,N_5206);
nand U5954 (N_5954,N_5156,N_5151);
nor U5955 (N_5955,N_5012,N_5160);
and U5956 (N_5956,N_5327,N_5416);
and U5957 (N_5957,N_5414,N_5284);
nand U5958 (N_5958,N_5147,N_5051);
and U5959 (N_5959,N_5069,N_5151);
and U5960 (N_5960,N_5043,N_5187);
or U5961 (N_5961,N_5496,N_5479);
nand U5962 (N_5962,N_5332,N_5153);
nor U5963 (N_5963,N_5423,N_5121);
nor U5964 (N_5964,N_5315,N_5418);
nor U5965 (N_5965,N_5480,N_5316);
nand U5966 (N_5966,N_5199,N_5279);
and U5967 (N_5967,N_5200,N_5155);
and U5968 (N_5968,N_5272,N_5430);
nand U5969 (N_5969,N_5490,N_5059);
or U5970 (N_5970,N_5417,N_5132);
nor U5971 (N_5971,N_5443,N_5266);
nand U5972 (N_5972,N_5378,N_5169);
nor U5973 (N_5973,N_5305,N_5146);
or U5974 (N_5974,N_5066,N_5448);
and U5975 (N_5975,N_5043,N_5029);
or U5976 (N_5976,N_5407,N_5421);
or U5977 (N_5977,N_5253,N_5322);
nand U5978 (N_5978,N_5378,N_5048);
or U5979 (N_5979,N_5018,N_5301);
and U5980 (N_5980,N_5485,N_5334);
nand U5981 (N_5981,N_5439,N_5124);
nand U5982 (N_5982,N_5095,N_5002);
or U5983 (N_5983,N_5013,N_5437);
and U5984 (N_5984,N_5068,N_5277);
or U5985 (N_5985,N_5042,N_5177);
nor U5986 (N_5986,N_5123,N_5081);
and U5987 (N_5987,N_5324,N_5448);
nor U5988 (N_5988,N_5069,N_5265);
nor U5989 (N_5989,N_5309,N_5038);
nor U5990 (N_5990,N_5231,N_5202);
nor U5991 (N_5991,N_5021,N_5303);
and U5992 (N_5992,N_5442,N_5129);
nor U5993 (N_5993,N_5348,N_5046);
or U5994 (N_5994,N_5111,N_5291);
or U5995 (N_5995,N_5189,N_5167);
or U5996 (N_5996,N_5342,N_5495);
nor U5997 (N_5997,N_5423,N_5046);
and U5998 (N_5998,N_5198,N_5323);
and U5999 (N_5999,N_5393,N_5038);
and U6000 (N_6000,N_5842,N_5816);
and U6001 (N_6001,N_5650,N_5770);
nor U6002 (N_6002,N_5546,N_5672);
nand U6003 (N_6003,N_5877,N_5890);
or U6004 (N_6004,N_5805,N_5804);
or U6005 (N_6005,N_5862,N_5675);
xor U6006 (N_6006,N_5826,N_5752);
and U6007 (N_6007,N_5560,N_5942);
or U6008 (N_6008,N_5745,N_5591);
and U6009 (N_6009,N_5637,N_5943);
nor U6010 (N_6010,N_5663,N_5714);
or U6011 (N_6011,N_5757,N_5506);
nand U6012 (N_6012,N_5711,N_5516);
and U6013 (N_6013,N_5790,N_5548);
nor U6014 (N_6014,N_5630,N_5631);
or U6015 (N_6015,N_5938,N_5901);
xor U6016 (N_6016,N_5824,N_5531);
nor U6017 (N_6017,N_5692,N_5744);
and U6018 (N_6018,N_5551,N_5583);
and U6019 (N_6019,N_5514,N_5620);
and U6020 (N_6020,N_5996,N_5573);
nor U6021 (N_6021,N_5882,N_5553);
and U6022 (N_6022,N_5905,N_5602);
or U6023 (N_6023,N_5661,N_5676);
and U6024 (N_6024,N_5852,N_5798);
or U6025 (N_6025,N_5712,N_5985);
nand U6026 (N_6026,N_5910,N_5728);
and U6027 (N_6027,N_5592,N_5521);
nor U6028 (N_6028,N_5850,N_5892);
or U6029 (N_6029,N_5847,N_5786);
or U6030 (N_6030,N_5549,N_5555);
nand U6031 (N_6031,N_5987,N_5965);
and U6032 (N_6032,N_5912,N_5530);
nand U6033 (N_6033,N_5715,N_5710);
nor U6034 (N_6034,N_5646,N_5505);
nor U6035 (N_6035,N_5833,N_5638);
or U6036 (N_6036,N_5709,N_5541);
xor U6037 (N_6037,N_5590,N_5927);
nand U6038 (N_6038,N_5542,N_5758);
nor U6039 (N_6039,N_5722,N_5754);
nand U6040 (N_6040,N_5688,N_5674);
and U6041 (N_6041,N_5843,N_5642);
or U6042 (N_6042,N_5670,N_5918);
and U6043 (N_6043,N_5500,N_5750);
or U6044 (N_6044,N_5601,N_5569);
and U6045 (N_6045,N_5789,N_5593);
nand U6046 (N_6046,N_5701,N_5515);
or U6047 (N_6047,N_5869,N_5700);
and U6048 (N_6048,N_5976,N_5787);
or U6049 (N_6049,N_5922,N_5823);
and U6050 (N_6050,N_5613,N_5561);
nor U6051 (N_6051,N_5831,N_5993);
or U6052 (N_6052,N_5643,N_5933);
nand U6053 (N_6053,N_5520,N_5753);
and U6054 (N_6054,N_5662,N_5510);
nand U6055 (N_6055,N_5582,N_5828);
or U6056 (N_6056,N_5960,N_5835);
nor U6057 (N_6057,N_5939,N_5717);
and U6058 (N_6058,N_5623,N_5950);
nor U6059 (N_6059,N_5628,N_5654);
nand U6060 (N_6060,N_5866,N_5565);
nand U6061 (N_6061,N_5800,N_5820);
nor U6062 (N_6062,N_5699,N_5647);
or U6063 (N_6063,N_5732,N_5718);
nand U6064 (N_6064,N_5879,N_5810);
and U6065 (N_6065,N_5603,N_5706);
or U6066 (N_6066,N_5973,N_5791);
or U6067 (N_6067,N_5867,N_5773);
or U6068 (N_6068,N_5746,N_5734);
and U6069 (N_6069,N_5951,N_5666);
nor U6070 (N_6070,N_5563,N_5512);
nand U6071 (N_6071,N_5969,N_5598);
and U6072 (N_6072,N_5599,N_5581);
nand U6073 (N_6073,N_5907,N_5839);
nor U6074 (N_6074,N_5802,N_5544);
nand U6075 (N_6075,N_5762,N_5731);
nor U6076 (N_6076,N_5977,N_5739);
nand U6077 (N_6077,N_5838,N_5696);
or U6078 (N_6078,N_5519,N_5697);
or U6079 (N_6079,N_5911,N_5920);
nand U6080 (N_6080,N_5606,N_5702);
or U6081 (N_6081,N_5749,N_5761);
nand U6082 (N_6082,N_5600,N_5868);
or U6083 (N_6083,N_5580,N_5508);
or U6084 (N_6084,N_5668,N_5503);
and U6085 (N_6085,N_5522,N_5854);
nor U6086 (N_6086,N_5884,N_5975);
nand U6087 (N_6087,N_5539,N_5664);
nor U6088 (N_6088,N_5849,N_5625);
nand U6089 (N_6089,N_5629,N_5693);
or U6090 (N_6090,N_5844,N_5764);
xnor U6091 (N_6091,N_5981,N_5878);
nor U6092 (N_6092,N_5946,N_5609);
and U6093 (N_6093,N_5558,N_5747);
nand U6094 (N_6094,N_5622,N_5538);
or U6095 (N_6095,N_5813,N_5963);
nand U6096 (N_6096,N_5990,N_5864);
nand U6097 (N_6097,N_5562,N_5799);
or U6098 (N_6098,N_5574,N_5897);
or U6099 (N_6099,N_5916,N_5829);
and U6100 (N_6100,N_5618,N_5783);
and U6101 (N_6101,N_5924,N_5934);
or U6102 (N_6102,N_5778,N_5932);
or U6103 (N_6103,N_5730,N_5874);
nand U6104 (N_6104,N_5611,N_5614);
or U6105 (N_6105,N_5641,N_5980);
nand U6106 (N_6106,N_5729,N_5794);
or U6107 (N_6107,N_5906,N_5954);
or U6108 (N_6108,N_5713,N_5639);
nand U6109 (N_6109,N_5653,N_5763);
or U6110 (N_6110,N_5527,N_5836);
and U6111 (N_6111,N_5535,N_5891);
nand U6112 (N_6112,N_5979,N_5735);
or U6113 (N_6113,N_5543,N_5955);
nor U6114 (N_6114,N_5814,N_5705);
nand U6115 (N_6115,N_5552,N_5776);
xnor U6116 (N_6116,N_5571,N_5765);
nor U6117 (N_6117,N_5694,N_5504);
or U6118 (N_6118,N_5957,N_5991);
and U6119 (N_6119,N_5930,N_5936);
and U6120 (N_6120,N_5658,N_5743);
nand U6121 (N_6121,N_5526,N_5665);
nand U6122 (N_6122,N_5785,N_5657);
and U6123 (N_6123,N_5883,N_5615);
and U6124 (N_6124,N_5940,N_5656);
or U6125 (N_6125,N_5880,N_5806);
or U6126 (N_6126,N_5627,N_5550);
or U6127 (N_6127,N_5781,N_5587);
nor U6128 (N_6128,N_5994,N_5989);
nor U6129 (N_6129,N_5748,N_5937);
or U6130 (N_6130,N_5695,N_5808);
nand U6131 (N_6131,N_5636,N_5511);
nor U6132 (N_6132,N_5534,N_5788);
nand U6133 (N_6133,N_5997,N_5673);
or U6134 (N_6134,N_5649,N_5859);
nand U6135 (N_6135,N_5983,N_5612);
nand U6136 (N_6136,N_5682,N_5952);
nand U6137 (N_6137,N_5853,N_5691);
or U6138 (N_6138,N_5872,N_5502);
nor U6139 (N_6139,N_5545,N_5733);
or U6140 (N_6140,N_5567,N_5570);
or U6141 (N_6141,N_5958,N_5875);
nand U6142 (N_6142,N_5660,N_5633);
and U6143 (N_6143,N_5564,N_5873);
nor U6144 (N_6144,N_5984,N_5517);
and U6145 (N_6145,N_5988,N_5585);
nand U6146 (N_6146,N_5677,N_5634);
nor U6147 (N_6147,N_5719,N_5982);
and U6148 (N_6148,N_5803,N_5832);
or U6149 (N_6149,N_5681,N_5685);
or U6150 (N_6150,N_5669,N_5815);
or U6151 (N_6151,N_5953,N_5528);
nand U6152 (N_6152,N_5857,N_5617);
nor U6153 (N_6153,N_5848,N_5796);
or U6154 (N_6154,N_5640,N_5568);
nor U6155 (N_6155,N_5588,N_5978);
nor U6156 (N_6156,N_5970,N_5784);
nor U6157 (N_6157,N_5774,N_5959);
nor U6158 (N_6158,N_5554,N_5533);
nand U6159 (N_6159,N_5819,N_5956);
nand U6160 (N_6160,N_5679,N_5888);
and U6161 (N_6161,N_5556,N_5557);
nand U6162 (N_6162,N_5525,N_5851);
and U6163 (N_6163,N_5738,N_5948);
nand U6164 (N_6164,N_5865,N_5651);
or U6165 (N_6165,N_5513,N_5935);
nor U6166 (N_6166,N_5822,N_5886);
and U6167 (N_6167,N_5834,N_5904);
or U6168 (N_6168,N_5579,N_5768);
or U6169 (N_6169,N_5876,N_5547);
or U6170 (N_6170,N_5889,N_5894);
nor U6171 (N_6171,N_5998,N_5610);
or U6172 (N_6172,N_5690,N_5724);
or U6173 (N_6173,N_5689,N_5921);
nor U6174 (N_6174,N_5902,N_5974);
nand U6175 (N_6175,N_5723,N_5594);
nand U6176 (N_6176,N_5777,N_5795);
and U6177 (N_6177,N_5687,N_5652);
and U6178 (N_6178,N_5575,N_5887);
nor U6179 (N_6179,N_5817,N_5586);
nor U6180 (N_6180,N_5725,N_5619);
xor U6181 (N_6181,N_5780,N_5755);
nor U6182 (N_6182,N_5949,N_5779);
and U6183 (N_6183,N_5896,N_5972);
nor U6184 (N_6184,N_5967,N_5596);
nand U6185 (N_6185,N_5576,N_5809);
or U6186 (N_6186,N_5947,N_5999);
nor U6187 (N_6187,N_5968,N_5861);
and U6188 (N_6188,N_5684,N_5792);
or U6189 (N_6189,N_5811,N_5756);
nand U6190 (N_6190,N_5917,N_5584);
or U6191 (N_6191,N_5616,N_5945);
and U6192 (N_6192,N_5807,N_5698);
nor U6193 (N_6193,N_5566,N_5863);
or U6194 (N_6194,N_5966,N_5645);
nor U6195 (N_6195,N_5925,N_5962);
nor U6196 (N_6196,N_5507,N_5821);
nor U6197 (N_6197,N_5532,N_5903);
or U6198 (N_6198,N_5680,N_5772);
nor U6199 (N_6199,N_5915,N_5767);
or U6200 (N_6200,N_5726,N_5881);
nor U6201 (N_6201,N_5621,N_5683);
xnor U6202 (N_6202,N_5841,N_5885);
or U6203 (N_6203,N_5742,N_5572);
nor U6204 (N_6204,N_5736,N_5860);
and U6205 (N_6205,N_5899,N_5626);
and U6206 (N_6206,N_5536,N_5919);
nand U6207 (N_6207,N_5518,N_5928);
nor U6208 (N_6208,N_5825,N_5678);
nor U6209 (N_6209,N_5971,N_5944);
or U6210 (N_6210,N_5659,N_5909);
and U6211 (N_6211,N_5608,N_5737);
nor U6212 (N_6212,N_5992,N_5686);
xor U6213 (N_6213,N_5741,N_5648);
nor U6214 (N_6214,N_5893,N_5870);
and U6215 (N_6215,N_5797,N_5529);
or U6216 (N_6216,N_5707,N_5635);
or U6217 (N_6217,N_5961,N_5855);
xnor U6218 (N_6218,N_5837,N_5858);
or U6219 (N_6219,N_5703,N_5793);
nand U6220 (N_6220,N_5523,N_5856);
and U6221 (N_6221,N_5827,N_5923);
nor U6222 (N_6222,N_5578,N_5605);
nand U6223 (N_6223,N_5607,N_5589);
or U6224 (N_6224,N_5509,N_5577);
nand U6225 (N_6225,N_5644,N_5771);
or U6226 (N_6226,N_5721,N_5830);
nor U6227 (N_6227,N_5812,N_5840);
or U6228 (N_6228,N_5929,N_5624);
and U6229 (N_6229,N_5760,N_5926);
nand U6230 (N_6230,N_5775,N_5524);
and U6231 (N_6231,N_5931,N_5845);
nor U6232 (N_6232,N_5986,N_5740);
nand U6233 (N_6233,N_5964,N_5871);
and U6234 (N_6234,N_5704,N_5537);
nand U6235 (N_6235,N_5941,N_5766);
xnor U6236 (N_6236,N_5727,N_5655);
and U6237 (N_6237,N_5782,N_5540);
and U6238 (N_6238,N_5895,N_5671);
nor U6239 (N_6239,N_5846,N_5759);
nand U6240 (N_6240,N_5913,N_5604);
xor U6241 (N_6241,N_5632,N_5751);
nor U6242 (N_6242,N_5716,N_5995);
nor U6243 (N_6243,N_5720,N_5914);
nand U6244 (N_6244,N_5898,N_5501);
or U6245 (N_6245,N_5908,N_5597);
and U6246 (N_6246,N_5818,N_5595);
and U6247 (N_6247,N_5559,N_5801);
nand U6248 (N_6248,N_5769,N_5708);
nor U6249 (N_6249,N_5667,N_5900);
nand U6250 (N_6250,N_5550,N_5882);
nand U6251 (N_6251,N_5844,N_5805);
nand U6252 (N_6252,N_5575,N_5900);
or U6253 (N_6253,N_5804,N_5612);
or U6254 (N_6254,N_5726,N_5887);
and U6255 (N_6255,N_5827,N_5864);
xor U6256 (N_6256,N_5673,N_5694);
nand U6257 (N_6257,N_5589,N_5936);
and U6258 (N_6258,N_5588,N_5716);
nand U6259 (N_6259,N_5737,N_5930);
nand U6260 (N_6260,N_5730,N_5803);
nand U6261 (N_6261,N_5590,N_5722);
and U6262 (N_6262,N_5928,N_5634);
or U6263 (N_6263,N_5841,N_5884);
and U6264 (N_6264,N_5722,N_5606);
nor U6265 (N_6265,N_5754,N_5858);
nor U6266 (N_6266,N_5594,N_5623);
nor U6267 (N_6267,N_5631,N_5812);
nor U6268 (N_6268,N_5990,N_5608);
and U6269 (N_6269,N_5580,N_5747);
or U6270 (N_6270,N_5598,N_5666);
and U6271 (N_6271,N_5749,N_5897);
or U6272 (N_6272,N_5689,N_5584);
nor U6273 (N_6273,N_5520,N_5727);
or U6274 (N_6274,N_5593,N_5882);
and U6275 (N_6275,N_5514,N_5934);
nand U6276 (N_6276,N_5898,N_5972);
nand U6277 (N_6277,N_5643,N_5732);
nor U6278 (N_6278,N_5551,N_5963);
nand U6279 (N_6279,N_5674,N_5919);
and U6280 (N_6280,N_5919,N_5687);
and U6281 (N_6281,N_5800,N_5847);
and U6282 (N_6282,N_5733,N_5825);
and U6283 (N_6283,N_5626,N_5959);
nor U6284 (N_6284,N_5839,N_5984);
or U6285 (N_6285,N_5677,N_5633);
nand U6286 (N_6286,N_5929,N_5575);
and U6287 (N_6287,N_5848,N_5537);
and U6288 (N_6288,N_5997,N_5512);
or U6289 (N_6289,N_5875,N_5836);
nand U6290 (N_6290,N_5675,N_5512);
or U6291 (N_6291,N_5711,N_5627);
or U6292 (N_6292,N_5745,N_5556);
and U6293 (N_6293,N_5918,N_5684);
or U6294 (N_6294,N_5656,N_5655);
nor U6295 (N_6295,N_5964,N_5749);
nor U6296 (N_6296,N_5627,N_5953);
nand U6297 (N_6297,N_5883,N_5539);
and U6298 (N_6298,N_5874,N_5908);
or U6299 (N_6299,N_5854,N_5925);
nor U6300 (N_6300,N_5633,N_5951);
and U6301 (N_6301,N_5528,N_5862);
and U6302 (N_6302,N_5956,N_5758);
or U6303 (N_6303,N_5866,N_5529);
and U6304 (N_6304,N_5677,N_5790);
nor U6305 (N_6305,N_5515,N_5925);
nand U6306 (N_6306,N_5823,N_5894);
xor U6307 (N_6307,N_5700,N_5917);
nand U6308 (N_6308,N_5884,N_5964);
nor U6309 (N_6309,N_5671,N_5599);
and U6310 (N_6310,N_5698,N_5952);
and U6311 (N_6311,N_5882,N_5595);
and U6312 (N_6312,N_5654,N_5745);
nand U6313 (N_6313,N_5997,N_5565);
nor U6314 (N_6314,N_5830,N_5973);
and U6315 (N_6315,N_5632,N_5604);
nand U6316 (N_6316,N_5604,N_5994);
nor U6317 (N_6317,N_5638,N_5811);
nor U6318 (N_6318,N_5886,N_5817);
nand U6319 (N_6319,N_5818,N_5529);
xnor U6320 (N_6320,N_5840,N_5563);
nand U6321 (N_6321,N_5988,N_5994);
and U6322 (N_6322,N_5644,N_5607);
and U6323 (N_6323,N_5803,N_5693);
nand U6324 (N_6324,N_5938,N_5555);
nor U6325 (N_6325,N_5903,N_5575);
and U6326 (N_6326,N_5744,N_5558);
nand U6327 (N_6327,N_5753,N_5870);
nor U6328 (N_6328,N_5546,N_5641);
nand U6329 (N_6329,N_5848,N_5776);
or U6330 (N_6330,N_5619,N_5700);
and U6331 (N_6331,N_5809,N_5557);
nand U6332 (N_6332,N_5960,N_5646);
nand U6333 (N_6333,N_5908,N_5648);
xor U6334 (N_6334,N_5501,N_5854);
or U6335 (N_6335,N_5650,N_5832);
nand U6336 (N_6336,N_5851,N_5673);
or U6337 (N_6337,N_5973,N_5690);
and U6338 (N_6338,N_5571,N_5502);
nor U6339 (N_6339,N_5553,N_5623);
or U6340 (N_6340,N_5580,N_5802);
and U6341 (N_6341,N_5830,N_5626);
nand U6342 (N_6342,N_5769,N_5765);
nor U6343 (N_6343,N_5993,N_5679);
nand U6344 (N_6344,N_5893,N_5979);
or U6345 (N_6345,N_5752,N_5512);
and U6346 (N_6346,N_5655,N_5523);
nand U6347 (N_6347,N_5990,N_5641);
nand U6348 (N_6348,N_5862,N_5648);
and U6349 (N_6349,N_5570,N_5787);
or U6350 (N_6350,N_5840,N_5805);
and U6351 (N_6351,N_5995,N_5548);
or U6352 (N_6352,N_5826,N_5898);
nor U6353 (N_6353,N_5640,N_5815);
or U6354 (N_6354,N_5672,N_5938);
and U6355 (N_6355,N_5725,N_5958);
or U6356 (N_6356,N_5973,N_5844);
nand U6357 (N_6357,N_5515,N_5804);
or U6358 (N_6358,N_5926,N_5790);
nand U6359 (N_6359,N_5595,N_5931);
or U6360 (N_6360,N_5573,N_5777);
or U6361 (N_6361,N_5855,N_5552);
nand U6362 (N_6362,N_5897,N_5540);
and U6363 (N_6363,N_5877,N_5604);
and U6364 (N_6364,N_5964,N_5536);
nand U6365 (N_6365,N_5721,N_5747);
and U6366 (N_6366,N_5749,N_5821);
nand U6367 (N_6367,N_5863,N_5777);
or U6368 (N_6368,N_5634,N_5740);
nor U6369 (N_6369,N_5733,N_5879);
or U6370 (N_6370,N_5656,N_5688);
and U6371 (N_6371,N_5503,N_5873);
or U6372 (N_6372,N_5963,N_5504);
nor U6373 (N_6373,N_5971,N_5586);
xor U6374 (N_6374,N_5622,N_5667);
or U6375 (N_6375,N_5524,N_5749);
or U6376 (N_6376,N_5540,N_5742);
nor U6377 (N_6377,N_5978,N_5665);
nor U6378 (N_6378,N_5859,N_5664);
and U6379 (N_6379,N_5957,N_5589);
and U6380 (N_6380,N_5515,N_5861);
or U6381 (N_6381,N_5723,N_5930);
or U6382 (N_6382,N_5754,N_5790);
xor U6383 (N_6383,N_5904,N_5792);
or U6384 (N_6384,N_5721,N_5990);
nand U6385 (N_6385,N_5815,N_5864);
or U6386 (N_6386,N_5599,N_5765);
and U6387 (N_6387,N_5603,N_5793);
nor U6388 (N_6388,N_5688,N_5984);
or U6389 (N_6389,N_5515,N_5647);
nor U6390 (N_6390,N_5688,N_5803);
nor U6391 (N_6391,N_5923,N_5916);
nand U6392 (N_6392,N_5586,N_5555);
nand U6393 (N_6393,N_5548,N_5613);
or U6394 (N_6394,N_5937,N_5509);
xnor U6395 (N_6395,N_5952,N_5633);
and U6396 (N_6396,N_5907,N_5510);
nor U6397 (N_6397,N_5749,N_5594);
or U6398 (N_6398,N_5629,N_5589);
nand U6399 (N_6399,N_5782,N_5885);
nor U6400 (N_6400,N_5500,N_5572);
nand U6401 (N_6401,N_5934,N_5611);
nand U6402 (N_6402,N_5966,N_5767);
nor U6403 (N_6403,N_5753,N_5947);
and U6404 (N_6404,N_5618,N_5714);
nand U6405 (N_6405,N_5916,N_5596);
nor U6406 (N_6406,N_5913,N_5666);
nand U6407 (N_6407,N_5520,N_5530);
and U6408 (N_6408,N_5614,N_5835);
nand U6409 (N_6409,N_5687,N_5603);
nor U6410 (N_6410,N_5818,N_5571);
and U6411 (N_6411,N_5616,N_5506);
and U6412 (N_6412,N_5600,N_5807);
and U6413 (N_6413,N_5544,N_5692);
or U6414 (N_6414,N_5891,N_5741);
xor U6415 (N_6415,N_5567,N_5822);
nand U6416 (N_6416,N_5640,N_5890);
nor U6417 (N_6417,N_5722,N_5579);
nand U6418 (N_6418,N_5879,N_5929);
or U6419 (N_6419,N_5744,N_5671);
or U6420 (N_6420,N_5565,N_5782);
and U6421 (N_6421,N_5701,N_5702);
and U6422 (N_6422,N_5757,N_5942);
and U6423 (N_6423,N_5769,N_5576);
nand U6424 (N_6424,N_5872,N_5792);
nand U6425 (N_6425,N_5591,N_5970);
and U6426 (N_6426,N_5797,N_5576);
or U6427 (N_6427,N_5734,N_5666);
and U6428 (N_6428,N_5977,N_5521);
nand U6429 (N_6429,N_5614,N_5992);
and U6430 (N_6430,N_5723,N_5868);
nand U6431 (N_6431,N_5766,N_5709);
nor U6432 (N_6432,N_5842,N_5703);
nor U6433 (N_6433,N_5882,N_5836);
and U6434 (N_6434,N_5922,N_5872);
nor U6435 (N_6435,N_5953,N_5952);
or U6436 (N_6436,N_5844,N_5606);
or U6437 (N_6437,N_5826,N_5717);
or U6438 (N_6438,N_5811,N_5673);
nand U6439 (N_6439,N_5628,N_5672);
and U6440 (N_6440,N_5758,N_5967);
xor U6441 (N_6441,N_5747,N_5641);
or U6442 (N_6442,N_5968,N_5956);
nor U6443 (N_6443,N_5871,N_5850);
and U6444 (N_6444,N_5669,N_5945);
or U6445 (N_6445,N_5878,N_5500);
nor U6446 (N_6446,N_5703,N_5666);
or U6447 (N_6447,N_5522,N_5967);
nor U6448 (N_6448,N_5950,N_5983);
nor U6449 (N_6449,N_5797,N_5670);
nor U6450 (N_6450,N_5677,N_5775);
and U6451 (N_6451,N_5717,N_5536);
or U6452 (N_6452,N_5901,N_5861);
and U6453 (N_6453,N_5726,N_5541);
or U6454 (N_6454,N_5850,N_5649);
nand U6455 (N_6455,N_5921,N_5842);
nor U6456 (N_6456,N_5682,N_5513);
and U6457 (N_6457,N_5880,N_5924);
or U6458 (N_6458,N_5569,N_5968);
nor U6459 (N_6459,N_5685,N_5506);
or U6460 (N_6460,N_5988,N_5942);
and U6461 (N_6461,N_5568,N_5637);
nand U6462 (N_6462,N_5721,N_5641);
nand U6463 (N_6463,N_5745,N_5526);
nor U6464 (N_6464,N_5501,N_5592);
nor U6465 (N_6465,N_5953,N_5509);
nand U6466 (N_6466,N_5708,N_5859);
nor U6467 (N_6467,N_5959,N_5563);
nor U6468 (N_6468,N_5771,N_5572);
nand U6469 (N_6469,N_5559,N_5546);
and U6470 (N_6470,N_5537,N_5751);
and U6471 (N_6471,N_5881,N_5776);
or U6472 (N_6472,N_5880,N_5581);
nand U6473 (N_6473,N_5854,N_5929);
nand U6474 (N_6474,N_5948,N_5778);
and U6475 (N_6475,N_5783,N_5581);
nor U6476 (N_6476,N_5628,N_5949);
xor U6477 (N_6477,N_5796,N_5815);
or U6478 (N_6478,N_5582,N_5937);
nor U6479 (N_6479,N_5695,N_5940);
nand U6480 (N_6480,N_5995,N_5513);
and U6481 (N_6481,N_5949,N_5687);
and U6482 (N_6482,N_5543,N_5949);
nor U6483 (N_6483,N_5604,N_5831);
xor U6484 (N_6484,N_5760,N_5953);
and U6485 (N_6485,N_5632,N_5621);
nor U6486 (N_6486,N_5576,N_5605);
or U6487 (N_6487,N_5687,N_5731);
nand U6488 (N_6488,N_5538,N_5747);
or U6489 (N_6489,N_5969,N_5520);
nor U6490 (N_6490,N_5847,N_5701);
or U6491 (N_6491,N_5516,N_5594);
nand U6492 (N_6492,N_5706,N_5950);
or U6493 (N_6493,N_5731,N_5608);
or U6494 (N_6494,N_5687,N_5825);
or U6495 (N_6495,N_5627,N_5917);
nor U6496 (N_6496,N_5796,N_5635);
nand U6497 (N_6497,N_5514,N_5626);
and U6498 (N_6498,N_5877,N_5533);
nand U6499 (N_6499,N_5524,N_5578);
and U6500 (N_6500,N_6295,N_6467);
or U6501 (N_6501,N_6032,N_6041);
or U6502 (N_6502,N_6352,N_6068);
nand U6503 (N_6503,N_6103,N_6289);
and U6504 (N_6504,N_6403,N_6280);
nor U6505 (N_6505,N_6065,N_6208);
nor U6506 (N_6506,N_6104,N_6482);
xnor U6507 (N_6507,N_6091,N_6227);
nand U6508 (N_6508,N_6464,N_6363);
nand U6509 (N_6509,N_6097,N_6051);
nand U6510 (N_6510,N_6402,N_6343);
or U6511 (N_6511,N_6284,N_6447);
or U6512 (N_6512,N_6146,N_6301);
nor U6513 (N_6513,N_6026,N_6052);
or U6514 (N_6514,N_6364,N_6048);
and U6515 (N_6515,N_6079,N_6281);
and U6516 (N_6516,N_6424,N_6331);
nor U6517 (N_6517,N_6012,N_6130);
nor U6518 (N_6518,N_6255,N_6073);
nor U6519 (N_6519,N_6421,N_6181);
nor U6520 (N_6520,N_6173,N_6209);
or U6521 (N_6521,N_6184,N_6000);
nand U6522 (N_6522,N_6192,N_6047);
nand U6523 (N_6523,N_6201,N_6194);
and U6524 (N_6524,N_6265,N_6136);
xnor U6525 (N_6525,N_6229,N_6231);
and U6526 (N_6526,N_6463,N_6419);
nor U6527 (N_6527,N_6334,N_6472);
nand U6528 (N_6528,N_6101,N_6355);
and U6529 (N_6529,N_6057,N_6242);
nor U6530 (N_6530,N_6155,N_6074);
or U6531 (N_6531,N_6043,N_6034);
or U6532 (N_6532,N_6491,N_6062);
nor U6533 (N_6533,N_6413,N_6011);
nand U6534 (N_6534,N_6028,N_6354);
and U6535 (N_6535,N_6185,N_6374);
nand U6536 (N_6536,N_6398,N_6444);
xnor U6537 (N_6537,N_6238,N_6342);
nor U6538 (N_6538,N_6456,N_6287);
nor U6539 (N_6539,N_6267,N_6159);
or U6540 (N_6540,N_6477,N_6039);
and U6541 (N_6541,N_6106,N_6326);
nand U6542 (N_6542,N_6025,N_6183);
nand U6543 (N_6543,N_6276,N_6266);
nand U6544 (N_6544,N_6246,N_6150);
nor U6545 (N_6545,N_6046,N_6001);
nand U6546 (N_6546,N_6323,N_6022);
or U6547 (N_6547,N_6067,N_6089);
nand U6548 (N_6548,N_6335,N_6061);
and U6549 (N_6549,N_6006,N_6239);
xor U6550 (N_6550,N_6263,N_6158);
nor U6551 (N_6551,N_6215,N_6451);
and U6552 (N_6552,N_6307,N_6291);
nor U6553 (N_6553,N_6296,N_6222);
and U6554 (N_6554,N_6008,N_6056);
or U6555 (N_6555,N_6015,N_6115);
and U6556 (N_6556,N_6492,N_6351);
or U6557 (N_6557,N_6282,N_6260);
nand U6558 (N_6558,N_6216,N_6270);
or U6559 (N_6559,N_6399,N_6198);
nand U6560 (N_6560,N_6415,N_6253);
nor U6561 (N_6561,N_6484,N_6496);
nor U6562 (N_6562,N_6225,N_6371);
and U6563 (N_6563,N_6273,N_6210);
or U6564 (N_6564,N_6095,N_6113);
or U6565 (N_6565,N_6096,N_6373);
or U6566 (N_6566,N_6489,N_6100);
nor U6567 (N_6567,N_6495,N_6176);
and U6568 (N_6568,N_6475,N_6059);
and U6569 (N_6569,N_6426,N_6064);
and U6570 (N_6570,N_6223,N_6336);
nand U6571 (N_6571,N_6414,N_6228);
nand U6572 (N_6572,N_6189,N_6483);
nor U6573 (N_6573,N_6377,N_6237);
and U6574 (N_6574,N_6082,N_6434);
and U6575 (N_6575,N_6197,N_6358);
and U6576 (N_6576,N_6160,N_6429);
and U6577 (N_6577,N_6007,N_6036);
and U6578 (N_6578,N_6166,N_6431);
nor U6579 (N_6579,N_6108,N_6473);
or U6580 (N_6580,N_6353,N_6257);
nor U6581 (N_6581,N_6448,N_6325);
or U6582 (N_6582,N_6345,N_6070);
or U6583 (N_6583,N_6169,N_6163);
nand U6584 (N_6584,N_6376,N_6172);
and U6585 (N_6585,N_6134,N_6144);
nor U6586 (N_6586,N_6387,N_6127);
nor U6587 (N_6587,N_6433,N_6412);
and U6588 (N_6588,N_6439,N_6220);
and U6589 (N_6589,N_6381,N_6436);
nand U6590 (N_6590,N_6205,N_6299);
nand U6591 (N_6591,N_6324,N_6234);
xnor U6592 (N_6592,N_6050,N_6114);
nand U6593 (N_6593,N_6244,N_6102);
nor U6594 (N_6594,N_6303,N_6411);
nor U6595 (N_6595,N_6131,N_6135);
nand U6596 (N_6596,N_6021,N_6151);
nor U6597 (N_6597,N_6124,N_6214);
nand U6598 (N_6598,N_6430,N_6404);
nor U6599 (N_6599,N_6165,N_6143);
or U6600 (N_6600,N_6002,N_6117);
or U6601 (N_6601,N_6081,N_6133);
nor U6602 (N_6602,N_6427,N_6190);
nand U6603 (N_6603,N_6129,N_6119);
or U6604 (N_6604,N_6357,N_6126);
or U6605 (N_6605,N_6031,N_6480);
nor U6606 (N_6606,N_6240,N_6443);
nand U6607 (N_6607,N_6243,N_6112);
nand U6608 (N_6608,N_6494,N_6359);
nand U6609 (N_6609,N_6196,N_6084);
and U6610 (N_6610,N_6379,N_6123);
and U6611 (N_6611,N_6422,N_6288);
nand U6612 (N_6612,N_6320,N_6232);
nor U6613 (N_6613,N_6476,N_6063);
nor U6614 (N_6614,N_6370,N_6395);
nor U6615 (N_6615,N_6252,N_6275);
or U6616 (N_6616,N_6453,N_6177);
nor U6617 (N_6617,N_6272,N_6054);
nor U6618 (N_6618,N_6157,N_6362);
nand U6619 (N_6619,N_6024,N_6072);
or U6620 (N_6620,N_6153,N_6250);
nor U6621 (N_6621,N_6066,N_6003);
nor U6622 (N_6622,N_6093,N_6087);
and U6623 (N_6623,N_6468,N_6236);
or U6624 (N_6624,N_6098,N_6298);
nor U6625 (N_6625,N_6269,N_6300);
or U6626 (N_6626,N_6116,N_6145);
nand U6627 (N_6627,N_6388,N_6302);
nand U6628 (N_6628,N_6040,N_6486);
nor U6629 (N_6629,N_6092,N_6014);
and U6630 (N_6630,N_6204,N_6086);
and U6631 (N_6631,N_6020,N_6442);
or U6632 (N_6632,N_6139,N_6122);
nand U6633 (N_6633,N_6230,N_6372);
nor U6634 (N_6634,N_6361,N_6211);
nand U6635 (N_6635,N_6271,N_6297);
and U6636 (N_6636,N_6200,N_6333);
and U6637 (N_6637,N_6397,N_6401);
or U6638 (N_6638,N_6341,N_6409);
nand U6639 (N_6639,N_6156,N_6154);
nand U6640 (N_6640,N_6389,N_6400);
nor U6641 (N_6641,N_6470,N_6278);
nor U6642 (N_6642,N_6487,N_6187);
nand U6643 (N_6643,N_6105,N_6152);
nor U6644 (N_6644,N_6206,N_6221);
and U6645 (N_6645,N_6202,N_6191);
or U6646 (N_6646,N_6418,N_6274);
and U6647 (N_6647,N_6010,N_6071);
or U6648 (N_6648,N_6249,N_6120);
nand U6649 (N_6649,N_6168,N_6233);
or U6650 (N_6650,N_6340,N_6140);
and U6651 (N_6651,N_6386,N_6245);
nor U6652 (N_6652,N_6290,N_6138);
nand U6653 (N_6653,N_6042,N_6217);
or U6654 (N_6654,N_6369,N_6179);
nor U6655 (N_6655,N_6450,N_6396);
and U6656 (N_6656,N_6294,N_6218);
nor U6657 (N_6657,N_6460,N_6425);
nand U6658 (N_6658,N_6279,N_6083);
nor U6659 (N_6659,N_6368,N_6485);
nor U6660 (N_6660,N_6408,N_6382);
nand U6661 (N_6661,N_6383,N_6348);
and U6662 (N_6662,N_6469,N_6224);
and U6663 (N_6663,N_6167,N_6349);
nand U6664 (N_6664,N_6393,N_6457);
nand U6665 (N_6665,N_6027,N_6023);
or U6666 (N_6666,N_6111,N_6474);
and U6667 (N_6667,N_6164,N_6235);
nand U6668 (N_6668,N_6058,N_6076);
nor U6669 (N_6669,N_6045,N_6219);
or U6670 (N_6670,N_6060,N_6432);
or U6671 (N_6671,N_6019,N_6292);
nand U6672 (N_6672,N_6384,N_6488);
nor U6673 (N_6673,N_6356,N_6213);
or U6674 (N_6674,N_6195,N_6329);
nand U6675 (N_6675,N_6304,N_6033);
or U6676 (N_6676,N_6365,N_6410);
and U6677 (N_6677,N_6435,N_6319);
nand U6678 (N_6678,N_6128,N_6327);
xor U6679 (N_6679,N_6286,N_6277);
or U6680 (N_6680,N_6479,N_6385);
nor U6681 (N_6681,N_6285,N_6121);
and U6682 (N_6682,N_6094,N_6132);
nor U6683 (N_6683,N_6142,N_6254);
or U6684 (N_6684,N_6391,N_6178);
nor U6685 (N_6685,N_6499,N_6446);
nand U6686 (N_6686,N_6258,N_6110);
nor U6687 (N_6687,N_6078,N_6321);
or U6688 (N_6688,N_6174,N_6458);
nand U6689 (N_6689,N_6423,N_6378);
nor U6690 (N_6690,N_6315,N_6309);
nor U6691 (N_6691,N_6080,N_6318);
and U6692 (N_6692,N_6462,N_6420);
nand U6693 (N_6693,N_6264,N_6149);
nor U6694 (N_6694,N_6037,N_6090);
nand U6695 (N_6695,N_6256,N_6322);
and U6696 (N_6696,N_6203,N_6030);
and U6697 (N_6697,N_6199,N_6044);
nand U6698 (N_6698,N_6344,N_6009);
or U6699 (N_6699,N_6171,N_6455);
nor U6700 (N_6700,N_6261,N_6490);
and U6701 (N_6701,N_6449,N_6170);
nor U6702 (N_6702,N_6310,N_6380);
or U6703 (N_6703,N_6350,N_6193);
and U6704 (N_6704,N_6162,N_6259);
or U6705 (N_6705,N_6212,N_6416);
and U6706 (N_6706,N_6375,N_6366);
nand U6707 (N_6707,N_6438,N_6498);
nand U6708 (N_6708,N_6226,N_6445);
or U6709 (N_6709,N_6038,N_6313);
and U6710 (N_6710,N_6088,N_6437);
nand U6711 (N_6711,N_6497,N_6004);
and U6712 (N_6712,N_6182,N_6029);
nand U6713 (N_6713,N_6312,N_6493);
or U6714 (N_6714,N_6268,N_6293);
and U6715 (N_6715,N_6186,N_6016);
nor U6716 (N_6716,N_6316,N_6077);
nor U6717 (N_6717,N_6099,N_6417);
and U6718 (N_6718,N_6018,N_6148);
nand U6719 (N_6719,N_6175,N_6330);
nand U6720 (N_6720,N_6459,N_6390);
and U6721 (N_6721,N_6314,N_6180);
or U6722 (N_6722,N_6405,N_6338);
nand U6723 (N_6723,N_6471,N_6406);
nor U6724 (N_6724,N_6465,N_6055);
or U6725 (N_6725,N_6317,N_6107);
nand U6726 (N_6726,N_6262,N_6251);
and U6727 (N_6727,N_6392,N_6118);
nor U6728 (N_6728,N_6109,N_6481);
and U6729 (N_6729,N_6085,N_6367);
and U6730 (N_6730,N_6035,N_6147);
nor U6731 (N_6731,N_6478,N_6049);
and U6732 (N_6732,N_6075,N_6360);
nor U6733 (N_6733,N_6141,N_6305);
or U6734 (N_6734,N_6053,N_6346);
or U6735 (N_6735,N_6339,N_6428);
or U6736 (N_6736,N_6247,N_6069);
or U6737 (N_6737,N_6241,N_6311);
or U6738 (N_6738,N_6407,N_6137);
and U6739 (N_6739,N_6394,N_6005);
nor U6740 (N_6740,N_6013,N_6248);
or U6741 (N_6741,N_6283,N_6466);
or U6742 (N_6742,N_6337,N_6332);
and U6743 (N_6743,N_6125,N_6347);
or U6744 (N_6744,N_6454,N_6452);
or U6745 (N_6745,N_6188,N_6306);
and U6746 (N_6746,N_6441,N_6440);
or U6747 (N_6747,N_6328,N_6461);
and U6748 (N_6748,N_6017,N_6207);
nor U6749 (N_6749,N_6161,N_6308);
xor U6750 (N_6750,N_6202,N_6131);
or U6751 (N_6751,N_6300,N_6178);
nor U6752 (N_6752,N_6429,N_6482);
and U6753 (N_6753,N_6074,N_6381);
or U6754 (N_6754,N_6485,N_6192);
or U6755 (N_6755,N_6314,N_6391);
nand U6756 (N_6756,N_6146,N_6132);
or U6757 (N_6757,N_6395,N_6204);
nand U6758 (N_6758,N_6350,N_6013);
or U6759 (N_6759,N_6105,N_6039);
or U6760 (N_6760,N_6009,N_6236);
nand U6761 (N_6761,N_6296,N_6267);
and U6762 (N_6762,N_6343,N_6301);
nor U6763 (N_6763,N_6041,N_6099);
nor U6764 (N_6764,N_6303,N_6243);
and U6765 (N_6765,N_6205,N_6383);
and U6766 (N_6766,N_6444,N_6493);
nor U6767 (N_6767,N_6271,N_6484);
nor U6768 (N_6768,N_6404,N_6187);
nor U6769 (N_6769,N_6064,N_6217);
or U6770 (N_6770,N_6091,N_6184);
nor U6771 (N_6771,N_6152,N_6110);
nand U6772 (N_6772,N_6018,N_6443);
nand U6773 (N_6773,N_6448,N_6449);
nor U6774 (N_6774,N_6350,N_6499);
and U6775 (N_6775,N_6249,N_6103);
or U6776 (N_6776,N_6403,N_6392);
nor U6777 (N_6777,N_6165,N_6266);
nand U6778 (N_6778,N_6262,N_6285);
nand U6779 (N_6779,N_6064,N_6041);
nor U6780 (N_6780,N_6350,N_6277);
and U6781 (N_6781,N_6169,N_6303);
and U6782 (N_6782,N_6053,N_6430);
nand U6783 (N_6783,N_6122,N_6166);
or U6784 (N_6784,N_6264,N_6349);
and U6785 (N_6785,N_6375,N_6094);
or U6786 (N_6786,N_6038,N_6105);
or U6787 (N_6787,N_6249,N_6015);
or U6788 (N_6788,N_6438,N_6422);
nand U6789 (N_6789,N_6096,N_6479);
or U6790 (N_6790,N_6176,N_6169);
or U6791 (N_6791,N_6010,N_6234);
nand U6792 (N_6792,N_6041,N_6074);
and U6793 (N_6793,N_6205,N_6332);
and U6794 (N_6794,N_6149,N_6112);
or U6795 (N_6795,N_6436,N_6432);
nand U6796 (N_6796,N_6419,N_6401);
nand U6797 (N_6797,N_6482,N_6189);
nand U6798 (N_6798,N_6100,N_6060);
or U6799 (N_6799,N_6293,N_6025);
nor U6800 (N_6800,N_6425,N_6123);
or U6801 (N_6801,N_6440,N_6113);
and U6802 (N_6802,N_6157,N_6371);
or U6803 (N_6803,N_6205,N_6142);
and U6804 (N_6804,N_6253,N_6385);
or U6805 (N_6805,N_6111,N_6330);
nor U6806 (N_6806,N_6306,N_6365);
nor U6807 (N_6807,N_6316,N_6171);
nor U6808 (N_6808,N_6370,N_6475);
or U6809 (N_6809,N_6158,N_6488);
nor U6810 (N_6810,N_6236,N_6183);
xnor U6811 (N_6811,N_6120,N_6022);
nand U6812 (N_6812,N_6087,N_6345);
and U6813 (N_6813,N_6295,N_6276);
nand U6814 (N_6814,N_6389,N_6130);
or U6815 (N_6815,N_6493,N_6253);
nand U6816 (N_6816,N_6417,N_6326);
nor U6817 (N_6817,N_6116,N_6480);
nand U6818 (N_6818,N_6357,N_6434);
xnor U6819 (N_6819,N_6357,N_6077);
or U6820 (N_6820,N_6271,N_6411);
nor U6821 (N_6821,N_6150,N_6000);
and U6822 (N_6822,N_6201,N_6276);
nand U6823 (N_6823,N_6071,N_6321);
or U6824 (N_6824,N_6212,N_6248);
nand U6825 (N_6825,N_6384,N_6426);
nor U6826 (N_6826,N_6147,N_6379);
nand U6827 (N_6827,N_6459,N_6475);
nor U6828 (N_6828,N_6377,N_6163);
and U6829 (N_6829,N_6284,N_6271);
or U6830 (N_6830,N_6155,N_6436);
and U6831 (N_6831,N_6056,N_6208);
and U6832 (N_6832,N_6071,N_6354);
nand U6833 (N_6833,N_6132,N_6364);
and U6834 (N_6834,N_6110,N_6146);
and U6835 (N_6835,N_6079,N_6494);
and U6836 (N_6836,N_6382,N_6425);
nor U6837 (N_6837,N_6348,N_6258);
or U6838 (N_6838,N_6124,N_6331);
and U6839 (N_6839,N_6495,N_6166);
nor U6840 (N_6840,N_6353,N_6120);
or U6841 (N_6841,N_6417,N_6010);
and U6842 (N_6842,N_6474,N_6497);
nand U6843 (N_6843,N_6035,N_6037);
nor U6844 (N_6844,N_6290,N_6404);
nor U6845 (N_6845,N_6144,N_6463);
and U6846 (N_6846,N_6499,N_6254);
or U6847 (N_6847,N_6159,N_6050);
and U6848 (N_6848,N_6440,N_6177);
nand U6849 (N_6849,N_6358,N_6234);
nor U6850 (N_6850,N_6397,N_6087);
nor U6851 (N_6851,N_6433,N_6479);
xor U6852 (N_6852,N_6421,N_6064);
nor U6853 (N_6853,N_6156,N_6314);
nand U6854 (N_6854,N_6089,N_6434);
and U6855 (N_6855,N_6420,N_6002);
or U6856 (N_6856,N_6127,N_6251);
or U6857 (N_6857,N_6213,N_6276);
nand U6858 (N_6858,N_6205,N_6415);
nand U6859 (N_6859,N_6106,N_6400);
or U6860 (N_6860,N_6489,N_6446);
nor U6861 (N_6861,N_6150,N_6139);
nor U6862 (N_6862,N_6377,N_6430);
nand U6863 (N_6863,N_6484,N_6090);
nand U6864 (N_6864,N_6147,N_6225);
nor U6865 (N_6865,N_6378,N_6415);
or U6866 (N_6866,N_6472,N_6100);
nor U6867 (N_6867,N_6308,N_6409);
and U6868 (N_6868,N_6262,N_6472);
nand U6869 (N_6869,N_6077,N_6258);
nor U6870 (N_6870,N_6185,N_6123);
nand U6871 (N_6871,N_6343,N_6454);
or U6872 (N_6872,N_6089,N_6467);
nand U6873 (N_6873,N_6450,N_6155);
nor U6874 (N_6874,N_6322,N_6469);
nor U6875 (N_6875,N_6020,N_6326);
nand U6876 (N_6876,N_6003,N_6373);
or U6877 (N_6877,N_6356,N_6070);
nand U6878 (N_6878,N_6449,N_6162);
nand U6879 (N_6879,N_6322,N_6299);
nor U6880 (N_6880,N_6389,N_6364);
and U6881 (N_6881,N_6388,N_6246);
nor U6882 (N_6882,N_6154,N_6439);
and U6883 (N_6883,N_6182,N_6082);
nand U6884 (N_6884,N_6126,N_6449);
or U6885 (N_6885,N_6103,N_6162);
and U6886 (N_6886,N_6496,N_6070);
and U6887 (N_6887,N_6015,N_6058);
xnor U6888 (N_6888,N_6064,N_6283);
and U6889 (N_6889,N_6486,N_6072);
nand U6890 (N_6890,N_6203,N_6003);
and U6891 (N_6891,N_6144,N_6167);
nand U6892 (N_6892,N_6003,N_6492);
nor U6893 (N_6893,N_6350,N_6240);
or U6894 (N_6894,N_6496,N_6054);
nor U6895 (N_6895,N_6335,N_6259);
or U6896 (N_6896,N_6075,N_6340);
nand U6897 (N_6897,N_6110,N_6193);
and U6898 (N_6898,N_6326,N_6117);
nor U6899 (N_6899,N_6455,N_6308);
nor U6900 (N_6900,N_6391,N_6277);
xnor U6901 (N_6901,N_6372,N_6366);
and U6902 (N_6902,N_6281,N_6033);
and U6903 (N_6903,N_6219,N_6252);
nor U6904 (N_6904,N_6012,N_6222);
and U6905 (N_6905,N_6227,N_6067);
or U6906 (N_6906,N_6011,N_6179);
nor U6907 (N_6907,N_6339,N_6348);
nand U6908 (N_6908,N_6075,N_6289);
nand U6909 (N_6909,N_6059,N_6028);
nand U6910 (N_6910,N_6109,N_6005);
or U6911 (N_6911,N_6028,N_6361);
nor U6912 (N_6912,N_6454,N_6190);
nor U6913 (N_6913,N_6005,N_6302);
and U6914 (N_6914,N_6219,N_6387);
nor U6915 (N_6915,N_6216,N_6293);
nor U6916 (N_6916,N_6486,N_6051);
nand U6917 (N_6917,N_6474,N_6454);
and U6918 (N_6918,N_6437,N_6369);
or U6919 (N_6919,N_6492,N_6032);
nand U6920 (N_6920,N_6134,N_6257);
nand U6921 (N_6921,N_6254,N_6299);
and U6922 (N_6922,N_6084,N_6223);
nand U6923 (N_6923,N_6435,N_6404);
or U6924 (N_6924,N_6094,N_6325);
or U6925 (N_6925,N_6452,N_6313);
nor U6926 (N_6926,N_6039,N_6247);
nor U6927 (N_6927,N_6342,N_6267);
nand U6928 (N_6928,N_6031,N_6003);
nand U6929 (N_6929,N_6072,N_6129);
or U6930 (N_6930,N_6424,N_6379);
or U6931 (N_6931,N_6470,N_6141);
and U6932 (N_6932,N_6101,N_6175);
nand U6933 (N_6933,N_6319,N_6349);
or U6934 (N_6934,N_6244,N_6423);
nor U6935 (N_6935,N_6307,N_6286);
and U6936 (N_6936,N_6076,N_6132);
or U6937 (N_6937,N_6074,N_6228);
or U6938 (N_6938,N_6330,N_6430);
nand U6939 (N_6939,N_6443,N_6488);
and U6940 (N_6940,N_6262,N_6032);
or U6941 (N_6941,N_6114,N_6317);
nor U6942 (N_6942,N_6358,N_6283);
and U6943 (N_6943,N_6285,N_6066);
or U6944 (N_6944,N_6482,N_6272);
nand U6945 (N_6945,N_6212,N_6007);
nor U6946 (N_6946,N_6318,N_6153);
nor U6947 (N_6947,N_6387,N_6193);
nor U6948 (N_6948,N_6170,N_6257);
nand U6949 (N_6949,N_6351,N_6341);
or U6950 (N_6950,N_6425,N_6048);
nand U6951 (N_6951,N_6112,N_6057);
nor U6952 (N_6952,N_6161,N_6264);
nor U6953 (N_6953,N_6386,N_6358);
nor U6954 (N_6954,N_6445,N_6170);
or U6955 (N_6955,N_6094,N_6355);
nand U6956 (N_6956,N_6457,N_6027);
and U6957 (N_6957,N_6088,N_6167);
or U6958 (N_6958,N_6438,N_6377);
or U6959 (N_6959,N_6012,N_6234);
nand U6960 (N_6960,N_6067,N_6152);
and U6961 (N_6961,N_6421,N_6066);
or U6962 (N_6962,N_6022,N_6012);
nor U6963 (N_6963,N_6240,N_6170);
nand U6964 (N_6964,N_6279,N_6148);
nor U6965 (N_6965,N_6273,N_6090);
nor U6966 (N_6966,N_6223,N_6033);
nor U6967 (N_6967,N_6121,N_6153);
nor U6968 (N_6968,N_6430,N_6190);
or U6969 (N_6969,N_6036,N_6268);
and U6970 (N_6970,N_6480,N_6344);
nor U6971 (N_6971,N_6280,N_6246);
or U6972 (N_6972,N_6067,N_6308);
and U6973 (N_6973,N_6260,N_6353);
nand U6974 (N_6974,N_6336,N_6117);
nor U6975 (N_6975,N_6027,N_6173);
or U6976 (N_6976,N_6136,N_6489);
nand U6977 (N_6977,N_6415,N_6289);
nand U6978 (N_6978,N_6332,N_6214);
and U6979 (N_6979,N_6211,N_6050);
nor U6980 (N_6980,N_6225,N_6276);
and U6981 (N_6981,N_6159,N_6358);
and U6982 (N_6982,N_6417,N_6055);
nand U6983 (N_6983,N_6387,N_6211);
or U6984 (N_6984,N_6002,N_6453);
nand U6985 (N_6985,N_6011,N_6455);
or U6986 (N_6986,N_6259,N_6407);
or U6987 (N_6987,N_6065,N_6220);
or U6988 (N_6988,N_6052,N_6267);
or U6989 (N_6989,N_6367,N_6399);
nor U6990 (N_6990,N_6142,N_6482);
nor U6991 (N_6991,N_6242,N_6470);
nand U6992 (N_6992,N_6282,N_6168);
nand U6993 (N_6993,N_6089,N_6352);
or U6994 (N_6994,N_6420,N_6394);
nand U6995 (N_6995,N_6214,N_6241);
and U6996 (N_6996,N_6303,N_6259);
nand U6997 (N_6997,N_6339,N_6487);
or U6998 (N_6998,N_6401,N_6420);
and U6999 (N_6999,N_6330,N_6392);
or U7000 (N_7000,N_6545,N_6541);
or U7001 (N_7001,N_6750,N_6946);
and U7002 (N_7002,N_6552,N_6897);
and U7003 (N_7003,N_6902,N_6717);
or U7004 (N_7004,N_6779,N_6691);
or U7005 (N_7005,N_6941,N_6736);
xnor U7006 (N_7006,N_6586,N_6727);
nand U7007 (N_7007,N_6653,N_6632);
or U7008 (N_7008,N_6561,N_6607);
or U7009 (N_7009,N_6602,N_6876);
and U7010 (N_7010,N_6765,N_6734);
or U7011 (N_7011,N_6683,N_6543);
or U7012 (N_7012,N_6973,N_6926);
nand U7013 (N_7013,N_6714,N_6771);
nor U7014 (N_7014,N_6540,N_6724);
and U7015 (N_7015,N_6842,N_6977);
nor U7016 (N_7016,N_6752,N_6594);
or U7017 (N_7017,N_6615,N_6888);
nand U7018 (N_7018,N_6682,N_6858);
nor U7019 (N_7019,N_6614,N_6609);
nor U7020 (N_7020,N_6922,N_6535);
nor U7021 (N_7021,N_6699,N_6638);
and U7022 (N_7022,N_6566,N_6984);
or U7023 (N_7023,N_6937,N_6532);
or U7024 (N_7024,N_6511,N_6515);
or U7025 (N_7025,N_6527,N_6673);
nor U7026 (N_7026,N_6994,N_6731);
and U7027 (N_7027,N_6675,N_6898);
nor U7028 (N_7028,N_6934,N_6684);
xnor U7029 (N_7029,N_6957,N_6563);
nor U7030 (N_7030,N_6667,N_6899);
and U7031 (N_7031,N_6835,N_6725);
and U7032 (N_7032,N_6849,N_6965);
nor U7033 (N_7033,N_6960,N_6801);
and U7034 (N_7034,N_6841,N_6840);
or U7035 (N_7035,N_6911,N_6534);
nor U7036 (N_7036,N_6892,N_6914);
nor U7037 (N_7037,N_6533,N_6523);
nand U7038 (N_7038,N_6593,N_6701);
nor U7039 (N_7039,N_6554,N_6744);
nand U7040 (N_7040,N_6516,N_6703);
nand U7041 (N_7041,N_6745,N_6716);
or U7042 (N_7042,N_6610,N_6780);
and U7043 (N_7043,N_6927,N_6695);
or U7044 (N_7044,N_6548,N_6950);
or U7045 (N_7045,N_6650,N_6549);
or U7046 (N_7046,N_6808,N_6597);
and U7047 (N_7047,N_6932,N_6880);
nor U7048 (N_7048,N_6512,N_6847);
or U7049 (N_7049,N_6816,N_6788);
and U7050 (N_7050,N_6974,N_6688);
nor U7051 (N_7051,N_6612,N_6613);
nor U7052 (N_7052,N_6671,N_6786);
xor U7053 (N_7053,N_6666,N_6753);
and U7054 (N_7054,N_6733,N_6850);
nand U7055 (N_7055,N_6944,N_6558);
nand U7056 (N_7056,N_6575,N_6958);
nor U7057 (N_7057,N_6580,N_6544);
or U7058 (N_7058,N_6542,N_6864);
or U7059 (N_7059,N_6879,N_6803);
or U7060 (N_7060,N_6576,N_6508);
and U7061 (N_7061,N_6955,N_6660);
or U7062 (N_7062,N_6737,N_6704);
and U7063 (N_7063,N_6741,N_6935);
and U7064 (N_7064,N_6500,N_6603);
and U7065 (N_7065,N_6793,N_6592);
nor U7066 (N_7066,N_6606,N_6975);
nand U7067 (N_7067,N_6848,N_6949);
or U7068 (N_7068,N_6598,N_6601);
or U7069 (N_7069,N_6505,N_6513);
or U7070 (N_7070,N_6645,N_6806);
nand U7071 (N_7071,N_6551,N_6782);
nor U7072 (N_7072,N_6800,N_6860);
or U7073 (N_7073,N_6812,N_6821);
nand U7074 (N_7074,N_6853,N_6913);
and U7075 (N_7075,N_6528,N_6730);
nand U7076 (N_7076,N_6875,N_6526);
or U7077 (N_7077,N_6751,N_6560);
nor U7078 (N_7078,N_6656,N_6985);
nor U7079 (N_7079,N_6851,N_6986);
or U7080 (N_7080,N_6915,N_6998);
xnor U7081 (N_7081,N_6758,N_6966);
nand U7082 (N_7082,N_6784,N_6546);
or U7083 (N_7083,N_6676,N_6686);
or U7084 (N_7084,N_6828,N_6895);
or U7085 (N_7085,N_6818,N_6877);
or U7086 (N_7086,N_6909,N_6789);
nand U7087 (N_7087,N_6547,N_6951);
nor U7088 (N_7088,N_6905,N_6729);
and U7089 (N_7089,N_6775,N_6945);
nor U7090 (N_7090,N_6881,N_6510);
or U7091 (N_7091,N_6893,N_6796);
nand U7092 (N_7092,N_6923,N_6577);
nor U7093 (N_7093,N_6567,N_6582);
nand U7094 (N_7094,N_6938,N_6988);
and U7095 (N_7095,N_6869,N_6524);
or U7096 (N_7096,N_6755,N_6930);
nor U7097 (N_7097,N_6556,N_6721);
nor U7098 (N_7098,N_6810,N_6962);
nor U7099 (N_7099,N_6630,N_6989);
or U7100 (N_7100,N_6891,N_6872);
and U7101 (N_7101,N_6885,N_6600);
nor U7102 (N_7102,N_6769,N_6863);
nand U7103 (N_7103,N_6936,N_6845);
and U7104 (N_7104,N_6790,N_6919);
or U7105 (N_7105,N_6861,N_6647);
nor U7106 (N_7106,N_6623,N_6629);
nand U7107 (N_7107,N_6642,N_6971);
or U7108 (N_7108,N_6662,N_6611);
nand U7109 (N_7109,N_6992,N_6823);
or U7110 (N_7110,N_6639,N_6735);
xnor U7111 (N_7111,N_6993,N_6762);
nor U7112 (N_7112,N_6652,N_6633);
or U7113 (N_7113,N_6907,N_6759);
or U7114 (N_7114,N_6956,N_6713);
and U7115 (N_7115,N_6857,N_6920);
nor U7116 (N_7116,N_6807,N_6723);
and U7117 (N_7117,N_6748,N_6596);
or U7118 (N_7118,N_6677,N_6952);
and U7119 (N_7119,N_6754,N_6933);
or U7120 (N_7120,N_6627,N_6967);
nand U7121 (N_7121,N_6996,N_6519);
nand U7122 (N_7122,N_6635,N_6792);
nor U7123 (N_7123,N_6870,N_6826);
or U7124 (N_7124,N_6641,N_6979);
or U7125 (N_7125,N_6648,N_6643);
nor U7126 (N_7126,N_6963,N_6504);
or U7127 (N_7127,N_6706,N_6619);
or U7128 (N_7128,N_6862,N_6839);
nor U7129 (N_7129,N_6772,N_6867);
or U7130 (N_7130,N_6700,N_6569);
xnor U7131 (N_7131,N_6530,N_6776);
nand U7132 (N_7132,N_6538,N_6931);
nor U7133 (N_7133,N_6692,N_6702);
or U7134 (N_7134,N_6657,N_6868);
and U7135 (N_7135,N_6697,N_6838);
nor U7136 (N_7136,N_6678,N_6763);
nor U7137 (N_7137,N_6943,N_6708);
xnor U7138 (N_7138,N_6608,N_6707);
and U7139 (N_7139,N_6777,N_6690);
and U7140 (N_7140,N_6559,N_6997);
or U7141 (N_7141,N_6681,N_6659);
and U7142 (N_7142,N_6517,N_6722);
nand U7143 (N_7143,N_6693,N_6756);
or U7144 (N_7144,N_6827,N_6910);
nand U7145 (N_7145,N_6621,N_6795);
or U7146 (N_7146,N_6908,N_6822);
and U7147 (N_7147,N_6987,N_6587);
nor U7148 (N_7148,N_6830,N_6571);
and U7149 (N_7149,N_6694,N_6947);
nand U7150 (N_7150,N_6886,N_6728);
nand U7151 (N_7151,N_6663,N_6742);
or U7152 (N_7152,N_6928,N_6636);
nor U7153 (N_7153,N_6900,N_6770);
xor U7154 (N_7154,N_6904,N_6605);
or U7155 (N_7155,N_6550,N_6815);
or U7156 (N_7156,N_6518,N_6537);
nor U7157 (N_7157,N_6964,N_6761);
and U7158 (N_7158,N_6814,N_6874);
nand U7159 (N_7159,N_6634,N_6674);
xor U7160 (N_7160,N_6732,N_6889);
nand U7161 (N_7161,N_6588,N_6799);
nor U7162 (N_7162,N_6720,N_6573);
xnor U7163 (N_7163,N_6918,N_6809);
or U7164 (N_7164,N_6712,N_6644);
nor U7165 (N_7165,N_6805,N_6747);
and U7166 (N_7166,N_6859,N_6521);
or U7167 (N_7167,N_6832,N_6531);
nand U7168 (N_7168,N_6649,N_6719);
nand U7169 (N_7169,N_6591,N_6766);
nor U7170 (N_7170,N_6651,N_6846);
nor U7171 (N_7171,N_6631,N_6884);
nor U7172 (N_7172,N_6718,N_6628);
and U7173 (N_7173,N_6583,N_6794);
nor U7174 (N_7174,N_6572,N_6968);
or U7175 (N_7175,N_6855,N_6953);
or U7176 (N_7176,N_6764,N_6698);
and U7177 (N_7177,N_6503,N_6620);
or U7178 (N_7178,N_6599,N_6959);
or U7179 (N_7179,N_6749,N_6873);
and U7180 (N_7180,N_6661,N_6804);
and U7181 (N_7181,N_6866,N_6564);
nand U7182 (N_7182,N_6990,N_6646);
and U7183 (N_7183,N_6680,N_6768);
nor U7184 (N_7184,N_6787,N_6579);
and U7185 (N_7185,N_6565,N_6813);
and U7186 (N_7186,N_6921,N_6501);
nor U7187 (N_7187,N_6970,N_6948);
or U7188 (N_7188,N_6562,N_6624);
and U7189 (N_7189,N_6983,N_6520);
nor U7190 (N_7190,N_6882,N_6595);
nand U7191 (N_7191,N_6901,N_6670);
nand U7192 (N_7192,N_6509,N_6865);
or U7193 (N_7193,N_6854,N_6689);
nor U7194 (N_7194,N_6995,N_6555);
nand U7195 (N_7195,N_6916,N_6536);
nor U7196 (N_7196,N_6658,N_6715);
and U7197 (N_7197,N_6890,N_6852);
or U7198 (N_7198,N_6553,N_6883);
nand U7199 (N_7199,N_6981,N_6817);
or U7200 (N_7200,N_6668,N_6570);
nor U7201 (N_7201,N_6696,N_6739);
or U7202 (N_7202,N_6672,N_6726);
or U7203 (N_7203,N_6585,N_6654);
or U7204 (N_7204,N_6925,N_6637);
nand U7205 (N_7205,N_6820,N_6616);
and U7206 (N_7206,N_6640,N_6685);
and U7207 (N_7207,N_6604,N_6502);
and U7208 (N_7208,N_6940,N_6797);
nor U7209 (N_7209,N_6584,N_6767);
nand U7210 (N_7210,N_6655,N_6557);
and U7211 (N_7211,N_6711,N_6906);
and U7212 (N_7212,N_6625,N_6878);
nand U7213 (N_7213,N_6578,N_6924);
and U7214 (N_7214,N_6679,N_6954);
or U7215 (N_7215,N_6590,N_6738);
nand U7216 (N_7216,N_6783,N_6746);
nand U7217 (N_7217,N_6819,N_6514);
or U7218 (N_7218,N_6999,N_6798);
or U7219 (N_7219,N_6781,N_6833);
nor U7220 (N_7220,N_6568,N_6991);
nor U7221 (N_7221,N_6773,N_6980);
nand U7222 (N_7222,N_6969,N_6778);
and U7223 (N_7223,N_6802,N_6837);
xnor U7224 (N_7224,N_6917,N_6836);
nor U7225 (N_7225,N_6939,N_6831);
nor U7226 (N_7226,N_6834,N_6581);
or U7227 (N_7227,N_6912,N_6929);
and U7228 (N_7228,N_6618,N_6825);
or U7229 (N_7229,N_6507,N_6844);
nand U7230 (N_7230,N_6589,N_6785);
nand U7231 (N_7231,N_6829,N_6539);
nand U7232 (N_7232,N_6871,N_6856);
or U7233 (N_7233,N_6811,N_6665);
nand U7234 (N_7234,N_6791,N_6978);
or U7235 (N_7235,N_6617,N_6743);
nand U7236 (N_7236,N_6709,N_6972);
nand U7237 (N_7237,N_6896,N_6622);
and U7238 (N_7238,N_6961,N_6976);
nor U7239 (N_7239,N_6705,N_6824);
nand U7240 (N_7240,N_6903,N_6894);
and U7241 (N_7241,N_6687,N_6982);
nor U7242 (N_7242,N_6774,N_6522);
and U7243 (N_7243,N_6669,N_6887);
and U7244 (N_7244,N_6574,N_6942);
and U7245 (N_7245,N_6710,N_6525);
nand U7246 (N_7246,N_6760,N_6843);
and U7247 (N_7247,N_6626,N_6664);
or U7248 (N_7248,N_6506,N_6740);
or U7249 (N_7249,N_6757,N_6529);
nand U7250 (N_7250,N_6756,N_6761);
and U7251 (N_7251,N_6766,N_6573);
nor U7252 (N_7252,N_6737,N_6870);
or U7253 (N_7253,N_6769,N_6740);
nand U7254 (N_7254,N_6604,N_6995);
nand U7255 (N_7255,N_6645,N_6709);
and U7256 (N_7256,N_6958,N_6692);
xor U7257 (N_7257,N_6621,N_6526);
nor U7258 (N_7258,N_6863,N_6823);
and U7259 (N_7259,N_6934,N_6968);
nor U7260 (N_7260,N_6751,N_6588);
nor U7261 (N_7261,N_6759,N_6972);
and U7262 (N_7262,N_6580,N_6738);
nand U7263 (N_7263,N_6791,N_6572);
xnor U7264 (N_7264,N_6920,N_6816);
or U7265 (N_7265,N_6649,N_6559);
or U7266 (N_7266,N_6661,N_6587);
and U7267 (N_7267,N_6583,N_6844);
or U7268 (N_7268,N_6596,N_6882);
and U7269 (N_7269,N_6902,N_6812);
nand U7270 (N_7270,N_6688,N_6912);
nor U7271 (N_7271,N_6646,N_6820);
and U7272 (N_7272,N_6883,N_6945);
or U7273 (N_7273,N_6559,N_6852);
and U7274 (N_7274,N_6734,N_6950);
and U7275 (N_7275,N_6824,N_6601);
or U7276 (N_7276,N_6949,N_6679);
or U7277 (N_7277,N_6688,N_6714);
and U7278 (N_7278,N_6661,N_6980);
xnor U7279 (N_7279,N_6538,N_6793);
or U7280 (N_7280,N_6695,N_6532);
nor U7281 (N_7281,N_6849,N_6681);
and U7282 (N_7282,N_6634,N_6824);
nand U7283 (N_7283,N_6978,N_6532);
nand U7284 (N_7284,N_6716,N_6648);
and U7285 (N_7285,N_6563,N_6946);
and U7286 (N_7286,N_6813,N_6716);
nor U7287 (N_7287,N_6673,N_6910);
or U7288 (N_7288,N_6639,N_6931);
nor U7289 (N_7289,N_6920,N_6910);
nand U7290 (N_7290,N_6500,N_6581);
nand U7291 (N_7291,N_6739,N_6852);
and U7292 (N_7292,N_6538,N_6731);
nor U7293 (N_7293,N_6884,N_6961);
or U7294 (N_7294,N_6983,N_6928);
or U7295 (N_7295,N_6527,N_6535);
and U7296 (N_7296,N_6987,N_6537);
nor U7297 (N_7297,N_6587,N_6867);
and U7298 (N_7298,N_6840,N_6945);
and U7299 (N_7299,N_6853,N_6944);
or U7300 (N_7300,N_6871,N_6732);
nand U7301 (N_7301,N_6629,N_6587);
and U7302 (N_7302,N_6711,N_6999);
xnor U7303 (N_7303,N_6801,N_6669);
nand U7304 (N_7304,N_6570,N_6951);
nand U7305 (N_7305,N_6707,N_6619);
nor U7306 (N_7306,N_6672,N_6543);
nor U7307 (N_7307,N_6623,N_6985);
nand U7308 (N_7308,N_6620,N_6939);
or U7309 (N_7309,N_6963,N_6703);
nand U7310 (N_7310,N_6847,N_6782);
and U7311 (N_7311,N_6615,N_6898);
nor U7312 (N_7312,N_6734,N_6782);
nor U7313 (N_7313,N_6717,N_6534);
xor U7314 (N_7314,N_6598,N_6696);
nor U7315 (N_7315,N_6956,N_6608);
nand U7316 (N_7316,N_6764,N_6908);
nor U7317 (N_7317,N_6617,N_6523);
or U7318 (N_7318,N_6898,N_6815);
or U7319 (N_7319,N_6733,N_6973);
and U7320 (N_7320,N_6912,N_6655);
nor U7321 (N_7321,N_6874,N_6923);
nand U7322 (N_7322,N_6995,N_6582);
nor U7323 (N_7323,N_6613,N_6911);
or U7324 (N_7324,N_6813,N_6965);
and U7325 (N_7325,N_6661,N_6999);
and U7326 (N_7326,N_6507,N_6798);
nor U7327 (N_7327,N_6824,N_6569);
and U7328 (N_7328,N_6617,N_6656);
and U7329 (N_7329,N_6603,N_6629);
or U7330 (N_7330,N_6605,N_6851);
nand U7331 (N_7331,N_6906,N_6777);
xnor U7332 (N_7332,N_6759,N_6677);
nor U7333 (N_7333,N_6820,N_6841);
nor U7334 (N_7334,N_6541,N_6623);
nor U7335 (N_7335,N_6745,N_6984);
and U7336 (N_7336,N_6971,N_6505);
and U7337 (N_7337,N_6795,N_6700);
nor U7338 (N_7338,N_6529,N_6661);
and U7339 (N_7339,N_6754,N_6526);
nor U7340 (N_7340,N_6992,N_6916);
nand U7341 (N_7341,N_6660,N_6583);
or U7342 (N_7342,N_6658,N_6962);
nand U7343 (N_7343,N_6624,N_6880);
or U7344 (N_7344,N_6691,N_6734);
and U7345 (N_7345,N_6722,N_6901);
nor U7346 (N_7346,N_6971,N_6768);
nand U7347 (N_7347,N_6978,N_6613);
nand U7348 (N_7348,N_6520,N_6660);
nor U7349 (N_7349,N_6742,N_6879);
nand U7350 (N_7350,N_6855,N_6736);
nand U7351 (N_7351,N_6993,N_6688);
and U7352 (N_7352,N_6874,N_6756);
nor U7353 (N_7353,N_6535,N_6814);
and U7354 (N_7354,N_6522,N_6842);
or U7355 (N_7355,N_6537,N_6793);
and U7356 (N_7356,N_6931,N_6807);
nand U7357 (N_7357,N_6815,N_6803);
nor U7358 (N_7358,N_6675,N_6922);
or U7359 (N_7359,N_6759,N_6990);
and U7360 (N_7360,N_6619,N_6953);
nor U7361 (N_7361,N_6695,N_6821);
or U7362 (N_7362,N_6851,N_6754);
and U7363 (N_7363,N_6592,N_6582);
nand U7364 (N_7364,N_6911,N_6813);
nand U7365 (N_7365,N_6792,N_6897);
nor U7366 (N_7366,N_6690,N_6969);
and U7367 (N_7367,N_6524,N_6930);
nand U7368 (N_7368,N_6523,N_6810);
and U7369 (N_7369,N_6698,N_6966);
nand U7370 (N_7370,N_6618,N_6591);
nand U7371 (N_7371,N_6582,N_6512);
or U7372 (N_7372,N_6812,N_6971);
nand U7373 (N_7373,N_6629,N_6579);
xor U7374 (N_7374,N_6818,N_6693);
nor U7375 (N_7375,N_6509,N_6982);
nor U7376 (N_7376,N_6953,N_6916);
and U7377 (N_7377,N_6835,N_6802);
nand U7378 (N_7378,N_6889,N_6702);
nand U7379 (N_7379,N_6886,N_6969);
nor U7380 (N_7380,N_6882,N_6599);
nand U7381 (N_7381,N_6538,N_6987);
or U7382 (N_7382,N_6623,N_6816);
and U7383 (N_7383,N_6709,N_6619);
or U7384 (N_7384,N_6651,N_6764);
or U7385 (N_7385,N_6787,N_6508);
or U7386 (N_7386,N_6851,N_6736);
nand U7387 (N_7387,N_6824,N_6756);
and U7388 (N_7388,N_6835,N_6862);
and U7389 (N_7389,N_6683,N_6818);
and U7390 (N_7390,N_6614,N_6862);
or U7391 (N_7391,N_6711,N_6705);
nand U7392 (N_7392,N_6513,N_6722);
and U7393 (N_7393,N_6885,N_6747);
nand U7394 (N_7394,N_6787,N_6993);
and U7395 (N_7395,N_6804,N_6701);
or U7396 (N_7396,N_6683,N_6822);
nand U7397 (N_7397,N_6821,N_6938);
or U7398 (N_7398,N_6824,N_6654);
or U7399 (N_7399,N_6996,N_6728);
and U7400 (N_7400,N_6906,N_6824);
nor U7401 (N_7401,N_6556,N_6884);
and U7402 (N_7402,N_6558,N_6703);
nor U7403 (N_7403,N_6823,N_6804);
nand U7404 (N_7404,N_6711,N_6959);
and U7405 (N_7405,N_6548,N_6757);
and U7406 (N_7406,N_6676,N_6576);
nand U7407 (N_7407,N_6969,N_6684);
or U7408 (N_7408,N_6805,N_6620);
nor U7409 (N_7409,N_6970,N_6510);
nor U7410 (N_7410,N_6825,N_6576);
or U7411 (N_7411,N_6791,N_6566);
or U7412 (N_7412,N_6817,N_6945);
xnor U7413 (N_7413,N_6652,N_6754);
or U7414 (N_7414,N_6584,N_6973);
or U7415 (N_7415,N_6514,N_6552);
or U7416 (N_7416,N_6840,N_6510);
and U7417 (N_7417,N_6527,N_6989);
and U7418 (N_7418,N_6564,N_6983);
or U7419 (N_7419,N_6710,N_6916);
nor U7420 (N_7420,N_6723,N_6840);
and U7421 (N_7421,N_6706,N_6654);
nand U7422 (N_7422,N_6725,N_6746);
nor U7423 (N_7423,N_6884,N_6511);
and U7424 (N_7424,N_6823,N_6903);
xnor U7425 (N_7425,N_6664,N_6818);
xnor U7426 (N_7426,N_6740,N_6688);
nand U7427 (N_7427,N_6874,N_6937);
or U7428 (N_7428,N_6893,N_6620);
or U7429 (N_7429,N_6585,N_6564);
nand U7430 (N_7430,N_6755,N_6693);
nand U7431 (N_7431,N_6762,N_6657);
nor U7432 (N_7432,N_6701,N_6824);
and U7433 (N_7433,N_6701,N_6722);
and U7434 (N_7434,N_6824,N_6541);
nand U7435 (N_7435,N_6631,N_6933);
or U7436 (N_7436,N_6558,N_6828);
and U7437 (N_7437,N_6659,N_6713);
and U7438 (N_7438,N_6957,N_6674);
or U7439 (N_7439,N_6501,N_6518);
nand U7440 (N_7440,N_6756,N_6896);
nor U7441 (N_7441,N_6824,N_6765);
and U7442 (N_7442,N_6589,N_6928);
and U7443 (N_7443,N_6873,N_6658);
nor U7444 (N_7444,N_6840,N_6738);
and U7445 (N_7445,N_6764,N_6506);
nor U7446 (N_7446,N_6981,N_6538);
nand U7447 (N_7447,N_6822,N_6700);
and U7448 (N_7448,N_6992,N_6808);
or U7449 (N_7449,N_6699,N_6687);
nor U7450 (N_7450,N_6589,N_6891);
and U7451 (N_7451,N_6601,N_6680);
or U7452 (N_7452,N_6929,N_6547);
or U7453 (N_7453,N_6971,N_6895);
and U7454 (N_7454,N_6689,N_6683);
nor U7455 (N_7455,N_6505,N_6556);
or U7456 (N_7456,N_6851,N_6962);
nand U7457 (N_7457,N_6816,N_6905);
nor U7458 (N_7458,N_6629,N_6673);
or U7459 (N_7459,N_6635,N_6542);
or U7460 (N_7460,N_6908,N_6760);
or U7461 (N_7461,N_6730,N_6701);
or U7462 (N_7462,N_6611,N_6844);
nand U7463 (N_7463,N_6869,N_6567);
nand U7464 (N_7464,N_6775,N_6980);
nand U7465 (N_7465,N_6979,N_6546);
and U7466 (N_7466,N_6658,N_6884);
or U7467 (N_7467,N_6639,N_6777);
nor U7468 (N_7468,N_6761,N_6910);
and U7469 (N_7469,N_6556,N_6996);
nor U7470 (N_7470,N_6816,N_6898);
xnor U7471 (N_7471,N_6785,N_6670);
xnor U7472 (N_7472,N_6894,N_6568);
nor U7473 (N_7473,N_6788,N_6810);
nor U7474 (N_7474,N_6827,N_6801);
nand U7475 (N_7475,N_6753,N_6627);
or U7476 (N_7476,N_6881,N_6772);
or U7477 (N_7477,N_6568,N_6839);
nand U7478 (N_7478,N_6588,N_6527);
or U7479 (N_7479,N_6537,N_6686);
nand U7480 (N_7480,N_6771,N_6987);
or U7481 (N_7481,N_6614,N_6933);
nor U7482 (N_7482,N_6520,N_6995);
or U7483 (N_7483,N_6676,N_6840);
or U7484 (N_7484,N_6764,N_6768);
nor U7485 (N_7485,N_6505,N_6783);
or U7486 (N_7486,N_6617,N_6601);
nand U7487 (N_7487,N_6611,N_6696);
nor U7488 (N_7488,N_6986,N_6648);
and U7489 (N_7489,N_6545,N_6865);
and U7490 (N_7490,N_6528,N_6837);
nor U7491 (N_7491,N_6667,N_6924);
or U7492 (N_7492,N_6716,N_6528);
and U7493 (N_7493,N_6595,N_6598);
nand U7494 (N_7494,N_6608,N_6859);
nand U7495 (N_7495,N_6662,N_6926);
nand U7496 (N_7496,N_6923,N_6884);
nor U7497 (N_7497,N_6654,N_6614);
or U7498 (N_7498,N_6744,N_6604);
nand U7499 (N_7499,N_6509,N_6689);
nand U7500 (N_7500,N_7256,N_7004);
nand U7501 (N_7501,N_7212,N_7450);
or U7502 (N_7502,N_7190,N_7264);
nand U7503 (N_7503,N_7204,N_7012);
or U7504 (N_7504,N_7369,N_7001);
and U7505 (N_7505,N_7437,N_7243);
nand U7506 (N_7506,N_7289,N_7439);
nand U7507 (N_7507,N_7087,N_7188);
nor U7508 (N_7508,N_7038,N_7265);
nand U7509 (N_7509,N_7385,N_7206);
nand U7510 (N_7510,N_7388,N_7468);
and U7511 (N_7511,N_7297,N_7014);
nand U7512 (N_7512,N_7063,N_7220);
or U7513 (N_7513,N_7294,N_7183);
nor U7514 (N_7514,N_7241,N_7093);
nor U7515 (N_7515,N_7086,N_7238);
nor U7516 (N_7516,N_7246,N_7406);
and U7517 (N_7517,N_7098,N_7455);
xor U7518 (N_7518,N_7454,N_7025);
or U7519 (N_7519,N_7445,N_7497);
nor U7520 (N_7520,N_7069,N_7193);
or U7521 (N_7521,N_7469,N_7167);
and U7522 (N_7522,N_7210,N_7415);
xor U7523 (N_7523,N_7307,N_7099);
and U7524 (N_7524,N_7104,N_7082);
and U7525 (N_7525,N_7333,N_7114);
or U7526 (N_7526,N_7016,N_7399);
nor U7527 (N_7527,N_7126,N_7225);
nand U7528 (N_7528,N_7000,N_7254);
nor U7529 (N_7529,N_7263,N_7118);
or U7530 (N_7530,N_7235,N_7164);
nand U7531 (N_7531,N_7361,N_7350);
and U7532 (N_7532,N_7481,N_7031);
and U7533 (N_7533,N_7041,N_7440);
nor U7534 (N_7534,N_7182,N_7330);
nor U7535 (N_7535,N_7144,N_7057);
nand U7536 (N_7536,N_7153,N_7302);
nor U7537 (N_7537,N_7127,N_7162);
nand U7538 (N_7538,N_7008,N_7325);
nor U7539 (N_7539,N_7271,N_7366);
nor U7540 (N_7540,N_7131,N_7424);
nor U7541 (N_7541,N_7298,N_7139);
and U7542 (N_7542,N_7384,N_7017);
nand U7543 (N_7543,N_7486,N_7493);
or U7544 (N_7544,N_7213,N_7052);
or U7545 (N_7545,N_7310,N_7077);
nor U7546 (N_7546,N_7261,N_7227);
nor U7547 (N_7547,N_7049,N_7018);
xor U7548 (N_7548,N_7354,N_7102);
nand U7549 (N_7549,N_7426,N_7343);
and U7550 (N_7550,N_7442,N_7059);
or U7551 (N_7551,N_7109,N_7039);
nor U7552 (N_7552,N_7129,N_7386);
and U7553 (N_7553,N_7140,N_7342);
or U7554 (N_7554,N_7376,N_7145);
or U7555 (N_7555,N_7165,N_7085);
or U7556 (N_7556,N_7390,N_7346);
and U7557 (N_7557,N_7159,N_7340);
nand U7558 (N_7558,N_7456,N_7134);
or U7559 (N_7559,N_7048,N_7335);
or U7560 (N_7560,N_7438,N_7436);
and U7561 (N_7561,N_7105,N_7427);
nand U7562 (N_7562,N_7146,N_7095);
xnor U7563 (N_7563,N_7355,N_7176);
or U7564 (N_7564,N_7321,N_7295);
nand U7565 (N_7565,N_7103,N_7215);
or U7566 (N_7566,N_7487,N_7009);
and U7567 (N_7567,N_7470,N_7222);
nor U7568 (N_7568,N_7040,N_7221);
nor U7569 (N_7569,N_7045,N_7150);
nand U7570 (N_7570,N_7071,N_7116);
nand U7571 (N_7571,N_7084,N_7304);
nand U7572 (N_7572,N_7396,N_7021);
nor U7573 (N_7573,N_7351,N_7453);
or U7574 (N_7574,N_7316,N_7180);
nor U7575 (N_7575,N_7312,N_7196);
nand U7576 (N_7576,N_7463,N_7160);
or U7577 (N_7577,N_7423,N_7257);
nor U7578 (N_7578,N_7466,N_7205);
or U7579 (N_7579,N_7447,N_7253);
nor U7580 (N_7580,N_7083,N_7410);
xnor U7581 (N_7581,N_7056,N_7244);
and U7582 (N_7582,N_7135,N_7154);
nor U7583 (N_7583,N_7022,N_7467);
nand U7584 (N_7584,N_7122,N_7349);
xnor U7585 (N_7585,N_7373,N_7251);
nor U7586 (N_7586,N_7090,N_7249);
nor U7587 (N_7587,N_7414,N_7152);
xnor U7588 (N_7588,N_7068,N_7494);
or U7589 (N_7589,N_7359,N_7132);
nand U7590 (N_7590,N_7327,N_7168);
nor U7591 (N_7591,N_7318,N_7451);
xnor U7592 (N_7592,N_7189,N_7051);
or U7593 (N_7593,N_7448,N_7058);
nor U7594 (N_7594,N_7383,N_7428);
nor U7595 (N_7595,N_7460,N_7268);
or U7596 (N_7596,N_7293,N_7080);
nand U7597 (N_7597,N_7203,N_7416);
or U7598 (N_7598,N_7314,N_7231);
or U7599 (N_7599,N_7282,N_7344);
and U7600 (N_7600,N_7322,N_7035);
or U7601 (N_7601,N_7108,N_7496);
nand U7602 (N_7602,N_7337,N_7036);
nand U7603 (N_7603,N_7461,N_7377);
nor U7604 (N_7604,N_7473,N_7197);
and U7605 (N_7605,N_7096,N_7192);
or U7606 (N_7606,N_7280,N_7315);
or U7607 (N_7607,N_7296,N_7136);
and U7608 (N_7608,N_7417,N_7174);
nor U7609 (N_7609,N_7171,N_7360);
nand U7610 (N_7610,N_7237,N_7113);
nor U7611 (N_7611,N_7299,N_7259);
and U7612 (N_7612,N_7065,N_7030);
or U7613 (N_7613,N_7229,N_7395);
and U7614 (N_7614,N_7290,N_7002);
and U7615 (N_7615,N_7248,N_7498);
nand U7616 (N_7616,N_7250,N_7010);
and U7617 (N_7617,N_7007,N_7362);
nand U7618 (N_7618,N_7397,N_7492);
and U7619 (N_7619,N_7483,N_7471);
and U7620 (N_7620,N_7430,N_7358);
and U7621 (N_7621,N_7042,N_7334);
and U7622 (N_7622,N_7005,N_7320);
and U7623 (N_7623,N_7425,N_7209);
and U7624 (N_7624,N_7200,N_7458);
nor U7625 (N_7625,N_7348,N_7207);
nand U7626 (N_7626,N_7173,N_7400);
or U7627 (N_7627,N_7123,N_7392);
nand U7628 (N_7628,N_7138,N_7043);
nand U7629 (N_7629,N_7462,N_7452);
nor U7630 (N_7630,N_7394,N_7181);
and U7631 (N_7631,N_7301,N_7491);
and U7632 (N_7632,N_7247,N_7091);
and U7633 (N_7633,N_7020,N_7378);
nand U7634 (N_7634,N_7357,N_7270);
or U7635 (N_7635,N_7232,N_7158);
xor U7636 (N_7636,N_7233,N_7094);
and U7637 (N_7637,N_7037,N_7236);
or U7638 (N_7638,N_7479,N_7034);
nand U7639 (N_7639,N_7194,N_7124);
nand U7640 (N_7640,N_7186,N_7311);
nand U7641 (N_7641,N_7029,N_7345);
or U7642 (N_7642,N_7081,N_7120);
nand U7643 (N_7643,N_7338,N_7285);
nor U7644 (N_7644,N_7305,N_7465);
or U7645 (N_7645,N_7121,N_7306);
and U7646 (N_7646,N_7089,N_7441);
or U7647 (N_7647,N_7101,N_7157);
and U7648 (N_7648,N_7476,N_7262);
and U7649 (N_7649,N_7364,N_7061);
and U7650 (N_7650,N_7119,N_7475);
nand U7651 (N_7651,N_7053,N_7402);
and U7652 (N_7652,N_7026,N_7365);
or U7653 (N_7653,N_7341,N_7485);
or U7654 (N_7654,N_7488,N_7329);
or U7655 (N_7655,N_7252,N_7279);
nand U7656 (N_7656,N_7177,N_7011);
and U7657 (N_7657,N_7495,N_7013);
or U7658 (N_7658,N_7412,N_7266);
or U7659 (N_7659,N_7179,N_7332);
or U7660 (N_7660,N_7272,N_7273);
and U7661 (N_7661,N_7143,N_7128);
or U7662 (N_7662,N_7133,N_7474);
nand U7663 (N_7663,N_7172,N_7142);
nor U7664 (N_7664,N_7184,N_7387);
and U7665 (N_7665,N_7393,N_7275);
nor U7666 (N_7666,N_7317,N_7352);
nand U7667 (N_7667,N_7398,N_7319);
or U7668 (N_7668,N_7381,N_7431);
and U7669 (N_7669,N_7175,N_7217);
or U7670 (N_7670,N_7218,N_7198);
xor U7671 (N_7671,N_7070,N_7224);
or U7672 (N_7672,N_7240,N_7353);
nand U7673 (N_7673,N_7405,N_7046);
nand U7674 (N_7674,N_7147,N_7490);
and U7675 (N_7675,N_7201,N_7499);
nand U7676 (N_7676,N_7404,N_7409);
nor U7677 (N_7677,N_7006,N_7389);
and U7678 (N_7678,N_7408,N_7478);
nor U7679 (N_7679,N_7418,N_7309);
nand U7680 (N_7680,N_7286,N_7422);
nor U7681 (N_7681,N_7234,N_7472);
and U7682 (N_7682,N_7278,N_7401);
nor U7683 (N_7683,N_7208,N_7434);
nand U7684 (N_7684,N_7161,N_7274);
and U7685 (N_7685,N_7245,N_7166);
nor U7686 (N_7686,N_7075,N_7281);
nor U7687 (N_7687,N_7115,N_7339);
and U7688 (N_7688,N_7382,N_7170);
nor U7689 (N_7689,N_7380,N_7072);
nand U7690 (N_7690,N_7024,N_7284);
and U7691 (N_7691,N_7187,N_7097);
xor U7692 (N_7692,N_7368,N_7420);
nor U7693 (N_7693,N_7027,N_7411);
nor U7694 (N_7694,N_7336,N_7100);
and U7695 (N_7695,N_7211,N_7269);
nand U7696 (N_7696,N_7323,N_7230);
nor U7697 (N_7697,N_7076,N_7375);
and U7698 (N_7698,N_7331,N_7260);
xor U7699 (N_7699,N_7363,N_7156);
or U7700 (N_7700,N_7219,N_7033);
or U7701 (N_7701,N_7356,N_7433);
nor U7702 (N_7702,N_7178,N_7028);
nor U7703 (N_7703,N_7374,N_7258);
or U7704 (N_7704,N_7223,N_7078);
nor U7705 (N_7705,N_7074,N_7226);
nor U7706 (N_7706,N_7313,N_7107);
or U7707 (N_7707,N_7019,N_7066);
and U7708 (N_7708,N_7328,N_7191);
and U7709 (N_7709,N_7276,N_7185);
or U7710 (N_7710,N_7370,N_7047);
nand U7711 (N_7711,N_7459,N_7443);
nor U7712 (N_7712,N_7435,N_7449);
and U7713 (N_7713,N_7239,N_7092);
and U7714 (N_7714,N_7482,N_7287);
nand U7715 (N_7715,N_7148,N_7106);
or U7716 (N_7716,N_7015,N_7073);
nor U7717 (N_7717,N_7267,N_7067);
nand U7718 (N_7718,N_7489,N_7088);
or U7719 (N_7719,N_7308,N_7419);
nand U7720 (N_7720,N_7292,N_7242);
nand U7721 (N_7721,N_7464,N_7117);
nand U7722 (N_7722,N_7023,N_7277);
nor U7723 (N_7723,N_7421,N_7137);
nand U7724 (N_7724,N_7060,N_7169);
and U7725 (N_7725,N_7480,N_7079);
or U7726 (N_7726,N_7155,N_7367);
nor U7727 (N_7727,N_7050,N_7413);
nand U7728 (N_7728,N_7202,N_7032);
and U7729 (N_7729,N_7003,N_7228);
or U7730 (N_7730,N_7444,N_7457);
nand U7731 (N_7731,N_7446,N_7347);
or U7732 (N_7732,N_7141,N_7149);
and U7733 (N_7733,N_7255,N_7195);
and U7734 (N_7734,N_7125,N_7055);
nor U7735 (N_7735,N_7062,N_7300);
nor U7736 (N_7736,N_7477,N_7151);
nand U7737 (N_7737,N_7429,N_7110);
nand U7738 (N_7738,N_7112,N_7054);
nand U7739 (N_7739,N_7379,N_7291);
nor U7740 (N_7740,N_7432,N_7044);
or U7741 (N_7741,N_7372,N_7324);
nand U7742 (N_7742,N_7403,N_7283);
nand U7743 (N_7743,N_7111,N_7216);
nor U7744 (N_7744,N_7199,N_7064);
or U7745 (N_7745,N_7303,N_7288);
and U7746 (N_7746,N_7326,N_7391);
nand U7747 (N_7747,N_7214,N_7130);
and U7748 (N_7748,N_7371,N_7407);
and U7749 (N_7749,N_7484,N_7163);
and U7750 (N_7750,N_7003,N_7145);
or U7751 (N_7751,N_7266,N_7363);
and U7752 (N_7752,N_7234,N_7367);
nor U7753 (N_7753,N_7204,N_7487);
nand U7754 (N_7754,N_7258,N_7098);
or U7755 (N_7755,N_7334,N_7210);
nor U7756 (N_7756,N_7072,N_7254);
and U7757 (N_7757,N_7443,N_7404);
and U7758 (N_7758,N_7415,N_7115);
nor U7759 (N_7759,N_7348,N_7341);
nand U7760 (N_7760,N_7006,N_7310);
nand U7761 (N_7761,N_7247,N_7476);
nand U7762 (N_7762,N_7420,N_7001);
or U7763 (N_7763,N_7288,N_7141);
nor U7764 (N_7764,N_7003,N_7120);
or U7765 (N_7765,N_7072,N_7308);
or U7766 (N_7766,N_7045,N_7176);
and U7767 (N_7767,N_7490,N_7122);
and U7768 (N_7768,N_7476,N_7029);
nand U7769 (N_7769,N_7219,N_7182);
nor U7770 (N_7770,N_7049,N_7052);
nor U7771 (N_7771,N_7274,N_7309);
or U7772 (N_7772,N_7463,N_7330);
and U7773 (N_7773,N_7015,N_7172);
nor U7774 (N_7774,N_7483,N_7170);
nand U7775 (N_7775,N_7386,N_7282);
and U7776 (N_7776,N_7228,N_7399);
and U7777 (N_7777,N_7334,N_7222);
nor U7778 (N_7778,N_7244,N_7005);
nand U7779 (N_7779,N_7360,N_7439);
and U7780 (N_7780,N_7016,N_7141);
nor U7781 (N_7781,N_7250,N_7489);
or U7782 (N_7782,N_7432,N_7363);
nand U7783 (N_7783,N_7437,N_7156);
and U7784 (N_7784,N_7266,N_7253);
or U7785 (N_7785,N_7470,N_7021);
xor U7786 (N_7786,N_7126,N_7459);
nor U7787 (N_7787,N_7117,N_7301);
or U7788 (N_7788,N_7110,N_7176);
and U7789 (N_7789,N_7011,N_7180);
nand U7790 (N_7790,N_7498,N_7278);
nand U7791 (N_7791,N_7323,N_7138);
nor U7792 (N_7792,N_7456,N_7150);
and U7793 (N_7793,N_7000,N_7238);
nand U7794 (N_7794,N_7077,N_7443);
and U7795 (N_7795,N_7062,N_7033);
and U7796 (N_7796,N_7053,N_7091);
xnor U7797 (N_7797,N_7165,N_7468);
and U7798 (N_7798,N_7441,N_7454);
or U7799 (N_7799,N_7176,N_7351);
nand U7800 (N_7800,N_7321,N_7275);
nand U7801 (N_7801,N_7296,N_7376);
nor U7802 (N_7802,N_7000,N_7259);
nand U7803 (N_7803,N_7327,N_7345);
nand U7804 (N_7804,N_7134,N_7168);
and U7805 (N_7805,N_7149,N_7271);
and U7806 (N_7806,N_7175,N_7464);
and U7807 (N_7807,N_7162,N_7130);
nand U7808 (N_7808,N_7120,N_7440);
nor U7809 (N_7809,N_7286,N_7074);
nor U7810 (N_7810,N_7113,N_7427);
nand U7811 (N_7811,N_7424,N_7201);
nand U7812 (N_7812,N_7162,N_7183);
nor U7813 (N_7813,N_7233,N_7302);
nand U7814 (N_7814,N_7072,N_7355);
or U7815 (N_7815,N_7236,N_7166);
nand U7816 (N_7816,N_7398,N_7253);
nor U7817 (N_7817,N_7266,N_7340);
nor U7818 (N_7818,N_7318,N_7270);
or U7819 (N_7819,N_7304,N_7468);
nand U7820 (N_7820,N_7358,N_7295);
or U7821 (N_7821,N_7248,N_7177);
nor U7822 (N_7822,N_7202,N_7383);
nor U7823 (N_7823,N_7154,N_7188);
nand U7824 (N_7824,N_7453,N_7331);
and U7825 (N_7825,N_7394,N_7304);
nor U7826 (N_7826,N_7128,N_7474);
or U7827 (N_7827,N_7089,N_7041);
and U7828 (N_7828,N_7051,N_7459);
nor U7829 (N_7829,N_7459,N_7097);
nor U7830 (N_7830,N_7480,N_7399);
xnor U7831 (N_7831,N_7300,N_7258);
nor U7832 (N_7832,N_7009,N_7235);
and U7833 (N_7833,N_7375,N_7389);
and U7834 (N_7834,N_7444,N_7035);
or U7835 (N_7835,N_7178,N_7299);
nand U7836 (N_7836,N_7412,N_7383);
and U7837 (N_7837,N_7244,N_7181);
xor U7838 (N_7838,N_7438,N_7368);
nand U7839 (N_7839,N_7151,N_7145);
or U7840 (N_7840,N_7137,N_7344);
or U7841 (N_7841,N_7223,N_7351);
nand U7842 (N_7842,N_7181,N_7350);
or U7843 (N_7843,N_7433,N_7005);
and U7844 (N_7844,N_7074,N_7380);
nand U7845 (N_7845,N_7402,N_7405);
nand U7846 (N_7846,N_7452,N_7310);
xnor U7847 (N_7847,N_7424,N_7050);
nand U7848 (N_7848,N_7277,N_7025);
or U7849 (N_7849,N_7369,N_7304);
nor U7850 (N_7850,N_7300,N_7198);
nor U7851 (N_7851,N_7026,N_7392);
or U7852 (N_7852,N_7398,N_7251);
and U7853 (N_7853,N_7396,N_7210);
or U7854 (N_7854,N_7372,N_7221);
nor U7855 (N_7855,N_7157,N_7424);
nor U7856 (N_7856,N_7089,N_7339);
or U7857 (N_7857,N_7124,N_7103);
nor U7858 (N_7858,N_7060,N_7367);
or U7859 (N_7859,N_7253,N_7194);
and U7860 (N_7860,N_7006,N_7499);
nor U7861 (N_7861,N_7037,N_7030);
and U7862 (N_7862,N_7402,N_7303);
or U7863 (N_7863,N_7122,N_7009);
nor U7864 (N_7864,N_7454,N_7006);
nand U7865 (N_7865,N_7339,N_7170);
nand U7866 (N_7866,N_7327,N_7199);
and U7867 (N_7867,N_7069,N_7300);
and U7868 (N_7868,N_7089,N_7302);
and U7869 (N_7869,N_7254,N_7194);
nor U7870 (N_7870,N_7032,N_7189);
nor U7871 (N_7871,N_7082,N_7089);
nor U7872 (N_7872,N_7002,N_7372);
and U7873 (N_7873,N_7388,N_7244);
nand U7874 (N_7874,N_7201,N_7046);
or U7875 (N_7875,N_7432,N_7372);
and U7876 (N_7876,N_7125,N_7071);
nor U7877 (N_7877,N_7456,N_7056);
or U7878 (N_7878,N_7195,N_7092);
nor U7879 (N_7879,N_7064,N_7319);
and U7880 (N_7880,N_7226,N_7173);
nand U7881 (N_7881,N_7342,N_7290);
and U7882 (N_7882,N_7276,N_7329);
nor U7883 (N_7883,N_7039,N_7318);
nand U7884 (N_7884,N_7255,N_7108);
nand U7885 (N_7885,N_7211,N_7368);
or U7886 (N_7886,N_7024,N_7292);
or U7887 (N_7887,N_7394,N_7194);
and U7888 (N_7888,N_7373,N_7360);
and U7889 (N_7889,N_7175,N_7372);
and U7890 (N_7890,N_7111,N_7299);
nor U7891 (N_7891,N_7124,N_7224);
nand U7892 (N_7892,N_7039,N_7151);
xnor U7893 (N_7893,N_7301,N_7327);
or U7894 (N_7894,N_7491,N_7017);
or U7895 (N_7895,N_7065,N_7332);
nand U7896 (N_7896,N_7026,N_7282);
and U7897 (N_7897,N_7129,N_7216);
xnor U7898 (N_7898,N_7276,N_7124);
and U7899 (N_7899,N_7127,N_7256);
nand U7900 (N_7900,N_7010,N_7030);
nor U7901 (N_7901,N_7005,N_7091);
nor U7902 (N_7902,N_7075,N_7068);
and U7903 (N_7903,N_7271,N_7221);
nor U7904 (N_7904,N_7051,N_7260);
nor U7905 (N_7905,N_7137,N_7261);
and U7906 (N_7906,N_7394,N_7171);
nand U7907 (N_7907,N_7147,N_7345);
or U7908 (N_7908,N_7377,N_7170);
nand U7909 (N_7909,N_7169,N_7417);
nand U7910 (N_7910,N_7431,N_7387);
nand U7911 (N_7911,N_7486,N_7123);
and U7912 (N_7912,N_7199,N_7376);
nand U7913 (N_7913,N_7331,N_7391);
and U7914 (N_7914,N_7363,N_7286);
and U7915 (N_7915,N_7063,N_7010);
and U7916 (N_7916,N_7466,N_7331);
or U7917 (N_7917,N_7371,N_7459);
nor U7918 (N_7918,N_7491,N_7449);
nand U7919 (N_7919,N_7114,N_7492);
and U7920 (N_7920,N_7265,N_7046);
nor U7921 (N_7921,N_7245,N_7280);
and U7922 (N_7922,N_7208,N_7203);
nand U7923 (N_7923,N_7062,N_7238);
nand U7924 (N_7924,N_7183,N_7199);
nand U7925 (N_7925,N_7129,N_7230);
and U7926 (N_7926,N_7407,N_7428);
nand U7927 (N_7927,N_7434,N_7310);
nand U7928 (N_7928,N_7317,N_7170);
nor U7929 (N_7929,N_7465,N_7075);
nand U7930 (N_7930,N_7118,N_7132);
or U7931 (N_7931,N_7243,N_7321);
nor U7932 (N_7932,N_7455,N_7259);
and U7933 (N_7933,N_7465,N_7072);
and U7934 (N_7934,N_7403,N_7125);
nand U7935 (N_7935,N_7376,N_7141);
and U7936 (N_7936,N_7452,N_7034);
nor U7937 (N_7937,N_7292,N_7499);
nand U7938 (N_7938,N_7255,N_7407);
or U7939 (N_7939,N_7063,N_7495);
nor U7940 (N_7940,N_7497,N_7249);
nor U7941 (N_7941,N_7040,N_7094);
nor U7942 (N_7942,N_7153,N_7021);
nor U7943 (N_7943,N_7446,N_7401);
nand U7944 (N_7944,N_7047,N_7432);
nand U7945 (N_7945,N_7070,N_7084);
or U7946 (N_7946,N_7061,N_7306);
nand U7947 (N_7947,N_7130,N_7038);
nor U7948 (N_7948,N_7404,N_7425);
nor U7949 (N_7949,N_7477,N_7450);
nor U7950 (N_7950,N_7233,N_7286);
or U7951 (N_7951,N_7005,N_7466);
or U7952 (N_7952,N_7124,N_7049);
nor U7953 (N_7953,N_7471,N_7351);
and U7954 (N_7954,N_7459,N_7017);
or U7955 (N_7955,N_7327,N_7243);
nand U7956 (N_7956,N_7143,N_7318);
nand U7957 (N_7957,N_7324,N_7026);
nor U7958 (N_7958,N_7485,N_7269);
or U7959 (N_7959,N_7156,N_7461);
or U7960 (N_7960,N_7049,N_7109);
nor U7961 (N_7961,N_7382,N_7412);
or U7962 (N_7962,N_7135,N_7339);
nor U7963 (N_7963,N_7039,N_7095);
nor U7964 (N_7964,N_7098,N_7062);
and U7965 (N_7965,N_7255,N_7353);
nor U7966 (N_7966,N_7311,N_7214);
or U7967 (N_7967,N_7301,N_7165);
and U7968 (N_7968,N_7130,N_7043);
and U7969 (N_7969,N_7134,N_7383);
nand U7970 (N_7970,N_7027,N_7021);
or U7971 (N_7971,N_7392,N_7269);
nand U7972 (N_7972,N_7242,N_7485);
nor U7973 (N_7973,N_7389,N_7323);
nor U7974 (N_7974,N_7411,N_7058);
or U7975 (N_7975,N_7049,N_7472);
and U7976 (N_7976,N_7344,N_7258);
and U7977 (N_7977,N_7421,N_7486);
xor U7978 (N_7978,N_7250,N_7289);
nand U7979 (N_7979,N_7174,N_7301);
nand U7980 (N_7980,N_7257,N_7179);
xnor U7981 (N_7981,N_7474,N_7248);
or U7982 (N_7982,N_7354,N_7000);
nor U7983 (N_7983,N_7407,N_7166);
or U7984 (N_7984,N_7481,N_7313);
and U7985 (N_7985,N_7204,N_7417);
or U7986 (N_7986,N_7355,N_7329);
or U7987 (N_7987,N_7420,N_7170);
or U7988 (N_7988,N_7380,N_7342);
and U7989 (N_7989,N_7381,N_7318);
and U7990 (N_7990,N_7148,N_7192);
nor U7991 (N_7991,N_7162,N_7288);
and U7992 (N_7992,N_7133,N_7320);
nand U7993 (N_7993,N_7444,N_7353);
and U7994 (N_7994,N_7138,N_7415);
nand U7995 (N_7995,N_7299,N_7143);
or U7996 (N_7996,N_7333,N_7346);
nor U7997 (N_7997,N_7347,N_7156);
or U7998 (N_7998,N_7224,N_7029);
xnor U7999 (N_7999,N_7152,N_7037);
and U8000 (N_8000,N_7894,N_7857);
or U8001 (N_8001,N_7807,N_7506);
or U8002 (N_8002,N_7595,N_7699);
and U8003 (N_8003,N_7989,N_7937);
or U8004 (N_8004,N_7603,N_7835);
nand U8005 (N_8005,N_7515,N_7765);
and U8006 (N_8006,N_7655,N_7793);
and U8007 (N_8007,N_7553,N_7853);
nand U8008 (N_8008,N_7896,N_7710);
or U8009 (N_8009,N_7675,N_7778);
nor U8010 (N_8010,N_7891,N_7683);
or U8011 (N_8011,N_7505,N_7747);
nor U8012 (N_8012,N_7795,N_7775);
or U8013 (N_8013,N_7789,N_7957);
and U8014 (N_8014,N_7801,N_7913);
or U8015 (N_8015,N_7950,N_7525);
or U8016 (N_8016,N_7735,N_7927);
nor U8017 (N_8017,N_7792,N_7830);
nor U8018 (N_8018,N_7696,N_7674);
or U8019 (N_8019,N_7728,N_7523);
nand U8020 (N_8020,N_7733,N_7871);
and U8021 (N_8021,N_7694,N_7978);
or U8022 (N_8022,N_7885,N_7941);
and U8023 (N_8023,N_7949,N_7856);
or U8024 (N_8024,N_7892,N_7817);
or U8025 (N_8025,N_7685,N_7668);
nor U8026 (N_8026,N_7709,N_7563);
or U8027 (N_8027,N_7863,N_7995);
and U8028 (N_8028,N_7667,N_7832);
nand U8029 (N_8029,N_7681,N_7712);
nand U8030 (N_8030,N_7592,N_7653);
and U8031 (N_8031,N_7504,N_7849);
nor U8032 (N_8032,N_7738,N_7952);
and U8033 (N_8033,N_7970,N_7847);
nor U8034 (N_8034,N_7658,N_7909);
xor U8035 (N_8035,N_7762,N_7917);
and U8036 (N_8036,N_7962,N_7533);
nand U8037 (N_8037,N_7895,N_7814);
nand U8038 (N_8038,N_7774,N_7583);
nand U8039 (N_8039,N_7586,N_7605);
nand U8040 (N_8040,N_7648,N_7898);
and U8041 (N_8041,N_7839,N_7890);
and U8042 (N_8042,N_7868,N_7878);
nand U8043 (N_8043,N_7576,N_7876);
nor U8044 (N_8044,N_7936,N_7600);
and U8045 (N_8045,N_7704,N_7611);
nand U8046 (N_8046,N_7804,N_7959);
and U8047 (N_8047,N_7919,N_7725);
and U8048 (N_8048,N_7811,N_7846);
nor U8049 (N_8049,N_7616,N_7698);
nand U8050 (N_8050,N_7692,N_7633);
nor U8051 (N_8051,N_7921,N_7569);
nor U8052 (N_8052,N_7671,N_7664);
nor U8053 (N_8053,N_7872,N_7755);
nor U8054 (N_8054,N_7954,N_7521);
xnor U8055 (N_8055,N_7622,N_7972);
nor U8056 (N_8056,N_7736,N_7718);
nor U8057 (N_8057,N_7720,N_7968);
nor U8058 (N_8058,N_7751,N_7707);
nor U8059 (N_8059,N_7708,N_7714);
nand U8060 (N_8060,N_7530,N_7851);
or U8061 (N_8061,N_7865,N_7679);
nand U8062 (N_8062,N_7688,N_7503);
and U8063 (N_8063,N_7606,N_7866);
or U8064 (N_8064,N_7854,N_7869);
and U8065 (N_8065,N_7572,N_7527);
nor U8066 (N_8066,N_7887,N_7838);
and U8067 (N_8067,N_7610,N_7982);
nor U8068 (N_8068,N_7634,N_7537);
or U8069 (N_8069,N_7691,N_7790);
nand U8070 (N_8070,N_7643,N_7624);
and U8071 (N_8071,N_7809,N_7686);
or U8072 (N_8072,N_7677,N_7639);
and U8073 (N_8073,N_7629,N_7619);
or U8074 (N_8074,N_7944,N_7621);
nand U8075 (N_8075,N_7964,N_7907);
nand U8076 (N_8076,N_7988,N_7693);
nor U8077 (N_8077,N_7877,N_7780);
nor U8078 (N_8078,N_7557,N_7717);
or U8079 (N_8079,N_7750,N_7594);
nor U8080 (N_8080,N_7934,N_7649);
and U8081 (N_8081,N_7609,N_7697);
or U8082 (N_8082,N_7742,N_7882);
nand U8083 (N_8083,N_7744,N_7690);
or U8084 (N_8084,N_7745,N_7993);
nor U8085 (N_8085,N_7822,N_7620);
or U8086 (N_8086,N_7935,N_7545);
nor U8087 (N_8087,N_7992,N_7925);
and U8088 (N_8088,N_7997,N_7584);
and U8089 (N_8089,N_7975,N_7991);
nand U8090 (N_8090,N_7770,N_7987);
or U8091 (N_8091,N_7884,N_7539);
or U8092 (N_8092,N_7948,N_7731);
nor U8093 (N_8093,N_7874,N_7676);
and U8094 (N_8094,N_7945,N_7973);
nand U8095 (N_8095,N_7580,N_7910);
xor U8096 (N_8096,N_7906,N_7980);
nand U8097 (N_8097,N_7916,N_7821);
nor U8098 (N_8098,N_7590,N_7858);
xor U8099 (N_8099,N_7705,N_7900);
xor U8100 (N_8100,N_7604,N_7538);
and U8101 (N_8101,N_7632,N_7746);
and U8102 (N_8102,N_7815,N_7743);
or U8103 (N_8103,N_7715,N_7631);
or U8104 (N_8104,N_7820,N_7623);
nor U8105 (N_8105,N_7568,N_7591);
nand U8106 (N_8106,N_7519,N_7625);
or U8107 (N_8107,N_7810,N_7646);
or U8108 (N_8108,N_7607,N_7889);
or U8109 (N_8109,N_7544,N_7627);
nor U8110 (N_8110,N_7642,N_7551);
nor U8111 (N_8111,N_7737,N_7641);
nor U8112 (N_8112,N_7756,N_7998);
nand U8113 (N_8113,N_7654,N_7831);
nand U8114 (N_8114,N_7500,N_7776);
nand U8115 (N_8115,N_7645,N_7661);
or U8116 (N_8116,N_7732,N_7946);
nor U8117 (N_8117,N_7902,N_7543);
xnor U8118 (N_8118,N_7908,N_7870);
or U8119 (N_8119,N_7665,N_7930);
and U8120 (N_8120,N_7759,N_7589);
nor U8121 (N_8121,N_7752,N_7764);
or U8122 (N_8122,N_7953,N_7999);
or U8123 (N_8123,N_7501,N_7638);
xnor U8124 (N_8124,N_7888,N_7926);
or U8125 (N_8125,N_7833,N_7798);
nor U8126 (N_8126,N_7836,N_7711);
nor U8127 (N_8127,N_7861,N_7758);
nand U8128 (N_8128,N_7626,N_7662);
or U8129 (N_8129,N_7981,N_7520);
and U8130 (N_8130,N_7787,N_7582);
nand U8131 (N_8131,N_7786,N_7848);
or U8132 (N_8132,N_7531,N_7785);
nand U8133 (N_8133,N_7796,N_7635);
nand U8134 (N_8134,N_7911,N_7976);
nor U8135 (N_8135,N_7922,N_7940);
nand U8136 (N_8136,N_7816,N_7554);
nand U8137 (N_8137,N_7771,N_7779);
nor U8138 (N_8138,N_7651,N_7966);
or U8139 (N_8139,N_7788,N_7640);
nor U8140 (N_8140,N_7573,N_7588);
nand U8141 (N_8141,N_7673,N_7886);
or U8142 (N_8142,N_7719,N_7579);
nand U8143 (N_8143,N_7904,N_7897);
nand U8144 (N_8144,N_7777,N_7529);
and U8145 (N_8145,N_7524,N_7805);
xnor U8146 (N_8146,N_7960,N_7985);
nor U8147 (N_8147,N_7703,N_7542);
and U8148 (N_8148,N_7819,N_7767);
nor U8149 (N_8149,N_7931,N_7628);
nand U8150 (N_8150,N_7799,N_7516);
or U8151 (N_8151,N_7791,N_7602);
and U8152 (N_8152,N_7552,N_7983);
nand U8153 (N_8153,N_7977,N_7630);
or U8154 (N_8154,N_7932,N_7522);
nor U8155 (N_8155,N_7956,N_7502);
or U8156 (N_8156,N_7802,N_7578);
or U8157 (N_8157,N_7867,N_7843);
or U8158 (N_8158,N_7899,N_7761);
or U8159 (N_8159,N_7650,N_7680);
and U8160 (N_8160,N_7612,N_7724);
nand U8161 (N_8161,N_7901,N_7608);
and U8162 (N_8162,N_7560,N_7528);
nor U8163 (N_8163,N_7617,N_7782);
or U8164 (N_8164,N_7647,N_7672);
nand U8165 (N_8165,N_7739,N_7965);
nand U8166 (N_8166,N_7684,N_7749);
nor U8167 (N_8167,N_7581,N_7905);
and U8168 (N_8168,N_7559,N_7864);
nand U8169 (N_8169,N_7852,N_7855);
nand U8170 (N_8170,N_7546,N_7549);
and U8171 (N_8171,N_7535,N_7880);
nor U8172 (N_8172,N_7585,N_7828);
nand U8173 (N_8173,N_7768,N_7912);
nand U8174 (N_8174,N_7984,N_7813);
or U8175 (N_8175,N_7687,N_7618);
nand U8176 (N_8176,N_7825,N_7967);
nor U8177 (N_8177,N_7883,N_7826);
nand U8178 (N_8178,N_7740,N_7824);
or U8179 (N_8179,N_7511,N_7656);
nand U8180 (N_8180,N_7596,N_7689);
nand U8181 (N_8181,N_7526,N_7682);
or U8182 (N_8182,N_7555,N_7772);
or U8183 (N_8183,N_7971,N_7808);
or U8184 (N_8184,N_7850,N_7574);
nor U8185 (N_8185,N_7829,N_7507);
or U8186 (N_8186,N_7567,N_7695);
nor U8187 (N_8187,N_7994,N_7875);
xor U8188 (N_8188,N_7548,N_7760);
nor U8189 (N_8189,N_7512,N_7969);
nor U8190 (N_8190,N_7918,N_7644);
nand U8191 (N_8191,N_7613,N_7769);
or U8192 (N_8192,N_7784,N_7781);
nand U8193 (N_8193,N_7513,N_7514);
nand U8194 (N_8194,N_7859,N_7701);
and U8195 (N_8195,N_7587,N_7963);
nor U8196 (N_8196,N_7734,N_7540);
or U8197 (N_8197,N_7547,N_7844);
or U8198 (N_8198,N_7598,N_7986);
nor U8199 (N_8199,N_7958,N_7722);
nor U8200 (N_8200,N_7669,N_7615);
and U8201 (N_8201,N_7575,N_7827);
nand U8202 (N_8202,N_7893,N_7637);
nand U8203 (N_8203,N_7562,N_7700);
nor U8204 (N_8204,N_7914,N_7881);
nor U8205 (N_8205,N_7534,N_7879);
nor U8206 (N_8206,N_7924,N_7800);
and U8207 (N_8207,N_7794,N_7721);
nand U8208 (N_8208,N_7943,N_7726);
and U8209 (N_8209,N_7518,N_7599);
nand U8210 (N_8210,N_7727,N_7571);
nand U8211 (N_8211,N_7840,N_7577);
or U8212 (N_8212,N_7845,N_7716);
or U8213 (N_8213,N_7510,N_7757);
nor U8214 (N_8214,N_7947,N_7837);
and U8215 (N_8215,N_7601,N_7860);
nand U8216 (N_8216,N_7558,N_7730);
or U8217 (N_8217,N_7713,N_7741);
nor U8218 (N_8218,N_7806,N_7990);
or U8219 (N_8219,N_7823,N_7841);
nor U8220 (N_8220,N_7938,N_7659);
and U8221 (N_8221,N_7564,N_7517);
nand U8222 (N_8222,N_7766,N_7797);
and U8223 (N_8223,N_7753,N_7536);
or U8224 (N_8224,N_7614,N_7812);
xor U8225 (N_8225,N_7652,N_7666);
nor U8226 (N_8226,N_7818,N_7928);
nor U8227 (N_8227,N_7803,N_7834);
nor U8228 (N_8228,N_7748,N_7566);
nand U8229 (N_8229,N_7570,N_7974);
and U8230 (N_8230,N_7783,N_7920);
or U8231 (N_8231,N_7657,N_7597);
or U8232 (N_8232,N_7862,N_7842);
nand U8233 (N_8233,N_7723,N_7763);
nand U8234 (N_8234,N_7903,N_7706);
or U8235 (N_8235,N_7929,N_7678);
or U8236 (N_8236,N_7541,N_7636);
nand U8237 (N_8237,N_7660,N_7561);
or U8238 (N_8238,N_7754,N_7873);
nor U8239 (N_8239,N_7979,N_7961);
nand U8240 (N_8240,N_7702,N_7942);
xor U8241 (N_8241,N_7951,N_7508);
nor U8242 (N_8242,N_7773,N_7996);
and U8243 (N_8243,N_7663,N_7556);
and U8244 (N_8244,N_7565,N_7593);
and U8245 (N_8245,N_7550,N_7670);
nand U8246 (N_8246,N_7532,N_7939);
nor U8247 (N_8247,N_7923,N_7729);
nand U8248 (N_8248,N_7955,N_7933);
nor U8249 (N_8249,N_7509,N_7915);
nor U8250 (N_8250,N_7552,N_7978);
xnor U8251 (N_8251,N_7538,N_7700);
nand U8252 (N_8252,N_7738,N_7961);
and U8253 (N_8253,N_7772,N_7581);
and U8254 (N_8254,N_7939,N_7873);
nor U8255 (N_8255,N_7737,N_7795);
nand U8256 (N_8256,N_7688,N_7546);
or U8257 (N_8257,N_7718,N_7609);
or U8258 (N_8258,N_7599,N_7631);
and U8259 (N_8259,N_7916,N_7698);
nor U8260 (N_8260,N_7733,N_7802);
nand U8261 (N_8261,N_7653,N_7561);
or U8262 (N_8262,N_7993,N_7778);
and U8263 (N_8263,N_7612,N_7899);
nor U8264 (N_8264,N_7808,N_7593);
and U8265 (N_8265,N_7879,N_7669);
nand U8266 (N_8266,N_7913,N_7725);
nand U8267 (N_8267,N_7814,N_7965);
nor U8268 (N_8268,N_7614,N_7766);
and U8269 (N_8269,N_7758,N_7787);
nor U8270 (N_8270,N_7658,N_7768);
and U8271 (N_8271,N_7721,N_7859);
nand U8272 (N_8272,N_7688,N_7718);
nand U8273 (N_8273,N_7822,N_7816);
or U8274 (N_8274,N_7854,N_7887);
and U8275 (N_8275,N_7622,N_7916);
and U8276 (N_8276,N_7566,N_7958);
and U8277 (N_8277,N_7756,N_7824);
or U8278 (N_8278,N_7677,N_7838);
nand U8279 (N_8279,N_7794,N_7955);
and U8280 (N_8280,N_7548,N_7946);
nand U8281 (N_8281,N_7938,N_7515);
and U8282 (N_8282,N_7923,N_7556);
or U8283 (N_8283,N_7876,N_7964);
and U8284 (N_8284,N_7681,N_7668);
nand U8285 (N_8285,N_7616,N_7822);
or U8286 (N_8286,N_7705,N_7512);
nand U8287 (N_8287,N_7706,N_7589);
or U8288 (N_8288,N_7909,N_7643);
nor U8289 (N_8289,N_7746,N_7567);
or U8290 (N_8290,N_7603,N_7794);
nand U8291 (N_8291,N_7681,N_7849);
nor U8292 (N_8292,N_7763,N_7699);
nor U8293 (N_8293,N_7522,N_7844);
nor U8294 (N_8294,N_7520,N_7590);
and U8295 (N_8295,N_7583,N_7695);
nor U8296 (N_8296,N_7552,N_7661);
or U8297 (N_8297,N_7626,N_7560);
and U8298 (N_8298,N_7920,N_7660);
nor U8299 (N_8299,N_7664,N_7503);
nor U8300 (N_8300,N_7779,N_7616);
nor U8301 (N_8301,N_7750,N_7589);
xnor U8302 (N_8302,N_7888,N_7759);
or U8303 (N_8303,N_7773,N_7853);
nand U8304 (N_8304,N_7772,N_7870);
nor U8305 (N_8305,N_7512,N_7758);
nand U8306 (N_8306,N_7519,N_7875);
and U8307 (N_8307,N_7730,N_7837);
nand U8308 (N_8308,N_7646,N_7856);
or U8309 (N_8309,N_7740,N_7869);
nor U8310 (N_8310,N_7693,N_7911);
or U8311 (N_8311,N_7974,N_7908);
or U8312 (N_8312,N_7969,N_7608);
nand U8313 (N_8313,N_7858,N_7652);
nor U8314 (N_8314,N_7889,N_7998);
xnor U8315 (N_8315,N_7757,N_7592);
or U8316 (N_8316,N_7724,N_7787);
or U8317 (N_8317,N_7606,N_7872);
or U8318 (N_8318,N_7577,N_7735);
xor U8319 (N_8319,N_7785,N_7836);
nand U8320 (N_8320,N_7798,N_7930);
nor U8321 (N_8321,N_7906,N_7541);
and U8322 (N_8322,N_7680,N_7624);
and U8323 (N_8323,N_7679,N_7783);
and U8324 (N_8324,N_7813,N_7691);
or U8325 (N_8325,N_7736,N_7559);
or U8326 (N_8326,N_7757,N_7740);
nand U8327 (N_8327,N_7773,N_7708);
or U8328 (N_8328,N_7764,N_7999);
nand U8329 (N_8329,N_7545,N_7980);
nor U8330 (N_8330,N_7568,N_7739);
nor U8331 (N_8331,N_7891,N_7642);
or U8332 (N_8332,N_7551,N_7601);
or U8333 (N_8333,N_7755,N_7912);
nand U8334 (N_8334,N_7534,N_7767);
or U8335 (N_8335,N_7545,N_7589);
nor U8336 (N_8336,N_7922,N_7670);
nor U8337 (N_8337,N_7788,N_7763);
and U8338 (N_8338,N_7545,N_7864);
and U8339 (N_8339,N_7969,N_7940);
nor U8340 (N_8340,N_7751,N_7661);
nor U8341 (N_8341,N_7568,N_7789);
nand U8342 (N_8342,N_7736,N_7892);
nor U8343 (N_8343,N_7710,N_7839);
nor U8344 (N_8344,N_7596,N_7933);
and U8345 (N_8345,N_7898,N_7658);
nand U8346 (N_8346,N_7976,N_7723);
and U8347 (N_8347,N_7614,N_7818);
and U8348 (N_8348,N_7511,N_7874);
and U8349 (N_8349,N_7837,N_7519);
or U8350 (N_8350,N_7790,N_7848);
or U8351 (N_8351,N_7995,N_7691);
and U8352 (N_8352,N_7645,N_7565);
nand U8353 (N_8353,N_7835,N_7976);
nand U8354 (N_8354,N_7681,N_7680);
nand U8355 (N_8355,N_7824,N_7764);
and U8356 (N_8356,N_7678,N_7753);
and U8357 (N_8357,N_7515,N_7907);
nor U8358 (N_8358,N_7965,N_7819);
nor U8359 (N_8359,N_7749,N_7555);
or U8360 (N_8360,N_7609,N_7612);
and U8361 (N_8361,N_7507,N_7506);
and U8362 (N_8362,N_7834,N_7838);
and U8363 (N_8363,N_7774,N_7676);
or U8364 (N_8364,N_7854,N_7755);
nor U8365 (N_8365,N_7951,N_7966);
nand U8366 (N_8366,N_7600,N_7656);
and U8367 (N_8367,N_7823,N_7976);
nor U8368 (N_8368,N_7597,N_7601);
or U8369 (N_8369,N_7898,N_7569);
and U8370 (N_8370,N_7723,N_7658);
or U8371 (N_8371,N_7692,N_7906);
and U8372 (N_8372,N_7863,N_7554);
or U8373 (N_8373,N_7864,N_7892);
nor U8374 (N_8374,N_7913,N_7713);
or U8375 (N_8375,N_7964,N_7510);
and U8376 (N_8376,N_7843,N_7931);
and U8377 (N_8377,N_7784,N_7840);
nor U8378 (N_8378,N_7991,N_7616);
or U8379 (N_8379,N_7628,N_7872);
and U8380 (N_8380,N_7800,N_7694);
nor U8381 (N_8381,N_7526,N_7599);
or U8382 (N_8382,N_7744,N_7736);
or U8383 (N_8383,N_7828,N_7806);
nor U8384 (N_8384,N_7577,N_7896);
or U8385 (N_8385,N_7880,N_7788);
nor U8386 (N_8386,N_7838,N_7616);
or U8387 (N_8387,N_7941,N_7775);
and U8388 (N_8388,N_7795,N_7730);
nand U8389 (N_8389,N_7608,N_7948);
nor U8390 (N_8390,N_7536,N_7738);
nand U8391 (N_8391,N_7528,N_7680);
or U8392 (N_8392,N_7629,N_7891);
nor U8393 (N_8393,N_7985,N_7833);
or U8394 (N_8394,N_7518,N_7661);
nor U8395 (N_8395,N_7992,N_7533);
nor U8396 (N_8396,N_7580,N_7619);
and U8397 (N_8397,N_7823,N_7505);
nor U8398 (N_8398,N_7856,N_7807);
and U8399 (N_8399,N_7926,N_7971);
or U8400 (N_8400,N_7988,N_7824);
and U8401 (N_8401,N_7512,N_7511);
nand U8402 (N_8402,N_7762,N_7633);
or U8403 (N_8403,N_7715,N_7520);
or U8404 (N_8404,N_7934,N_7611);
and U8405 (N_8405,N_7856,N_7969);
nand U8406 (N_8406,N_7604,N_7663);
and U8407 (N_8407,N_7613,N_7793);
and U8408 (N_8408,N_7707,N_7699);
nand U8409 (N_8409,N_7653,N_7956);
nand U8410 (N_8410,N_7575,N_7931);
nor U8411 (N_8411,N_7603,N_7954);
and U8412 (N_8412,N_7636,N_7927);
nor U8413 (N_8413,N_7533,N_7516);
or U8414 (N_8414,N_7771,N_7577);
or U8415 (N_8415,N_7640,N_7965);
or U8416 (N_8416,N_7967,N_7701);
nand U8417 (N_8417,N_7558,N_7536);
and U8418 (N_8418,N_7836,N_7504);
nor U8419 (N_8419,N_7954,N_7505);
xnor U8420 (N_8420,N_7837,N_7676);
and U8421 (N_8421,N_7905,N_7678);
nand U8422 (N_8422,N_7773,N_7859);
nand U8423 (N_8423,N_7643,N_7523);
nand U8424 (N_8424,N_7925,N_7571);
or U8425 (N_8425,N_7971,N_7631);
or U8426 (N_8426,N_7973,N_7700);
or U8427 (N_8427,N_7899,N_7715);
nand U8428 (N_8428,N_7733,N_7714);
and U8429 (N_8429,N_7787,N_7756);
and U8430 (N_8430,N_7990,N_7808);
or U8431 (N_8431,N_7574,N_7599);
xnor U8432 (N_8432,N_7537,N_7548);
xnor U8433 (N_8433,N_7668,N_7634);
and U8434 (N_8434,N_7624,N_7826);
or U8435 (N_8435,N_7871,N_7820);
or U8436 (N_8436,N_7984,N_7601);
nand U8437 (N_8437,N_7947,N_7910);
nor U8438 (N_8438,N_7837,N_7890);
nand U8439 (N_8439,N_7801,N_7795);
nand U8440 (N_8440,N_7648,N_7540);
nand U8441 (N_8441,N_7816,N_7564);
and U8442 (N_8442,N_7670,N_7666);
or U8443 (N_8443,N_7867,N_7728);
and U8444 (N_8444,N_7598,N_7690);
or U8445 (N_8445,N_7700,N_7832);
or U8446 (N_8446,N_7644,N_7566);
and U8447 (N_8447,N_7990,N_7984);
and U8448 (N_8448,N_7755,N_7884);
and U8449 (N_8449,N_7537,N_7855);
and U8450 (N_8450,N_7655,N_7912);
nor U8451 (N_8451,N_7720,N_7754);
or U8452 (N_8452,N_7796,N_7900);
nand U8453 (N_8453,N_7911,N_7719);
nand U8454 (N_8454,N_7931,N_7560);
nor U8455 (N_8455,N_7709,N_7890);
nand U8456 (N_8456,N_7643,N_7749);
or U8457 (N_8457,N_7690,N_7735);
and U8458 (N_8458,N_7681,N_7983);
nor U8459 (N_8459,N_7657,N_7726);
nand U8460 (N_8460,N_7646,N_7723);
nand U8461 (N_8461,N_7530,N_7953);
or U8462 (N_8462,N_7569,N_7627);
nor U8463 (N_8463,N_7976,N_7918);
or U8464 (N_8464,N_7944,N_7720);
or U8465 (N_8465,N_7818,N_7697);
or U8466 (N_8466,N_7910,N_7604);
nand U8467 (N_8467,N_7842,N_7961);
nor U8468 (N_8468,N_7588,N_7897);
and U8469 (N_8469,N_7814,N_7682);
or U8470 (N_8470,N_7612,N_7624);
nand U8471 (N_8471,N_7679,N_7922);
nor U8472 (N_8472,N_7813,N_7968);
and U8473 (N_8473,N_7864,N_7976);
or U8474 (N_8474,N_7996,N_7555);
nand U8475 (N_8475,N_7708,N_7899);
and U8476 (N_8476,N_7723,N_7719);
and U8477 (N_8477,N_7505,N_7576);
nand U8478 (N_8478,N_7537,N_7899);
and U8479 (N_8479,N_7902,N_7594);
and U8480 (N_8480,N_7765,N_7960);
nand U8481 (N_8481,N_7818,N_7645);
nand U8482 (N_8482,N_7966,N_7681);
and U8483 (N_8483,N_7973,N_7876);
and U8484 (N_8484,N_7946,N_7500);
nand U8485 (N_8485,N_7548,N_7921);
nor U8486 (N_8486,N_7658,N_7968);
and U8487 (N_8487,N_7779,N_7862);
or U8488 (N_8488,N_7852,N_7769);
nand U8489 (N_8489,N_7679,N_7937);
or U8490 (N_8490,N_7977,N_7995);
nand U8491 (N_8491,N_7821,N_7694);
and U8492 (N_8492,N_7895,N_7788);
or U8493 (N_8493,N_7958,N_7654);
xnor U8494 (N_8494,N_7615,N_7750);
xnor U8495 (N_8495,N_7509,N_7772);
nand U8496 (N_8496,N_7910,N_7908);
nand U8497 (N_8497,N_7952,N_7935);
nor U8498 (N_8498,N_7581,N_7913);
and U8499 (N_8499,N_7963,N_7865);
and U8500 (N_8500,N_8366,N_8185);
and U8501 (N_8501,N_8465,N_8142);
xnor U8502 (N_8502,N_8126,N_8494);
and U8503 (N_8503,N_8359,N_8081);
nor U8504 (N_8504,N_8368,N_8098);
and U8505 (N_8505,N_8171,N_8316);
nor U8506 (N_8506,N_8281,N_8196);
and U8507 (N_8507,N_8271,N_8493);
and U8508 (N_8508,N_8254,N_8434);
nor U8509 (N_8509,N_8320,N_8016);
or U8510 (N_8510,N_8438,N_8147);
nor U8511 (N_8511,N_8108,N_8045);
or U8512 (N_8512,N_8051,N_8343);
or U8513 (N_8513,N_8236,N_8223);
nand U8514 (N_8514,N_8232,N_8482);
nor U8515 (N_8515,N_8305,N_8445);
or U8516 (N_8516,N_8360,N_8161);
nor U8517 (N_8517,N_8273,N_8308);
and U8518 (N_8518,N_8246,N_8119);
nand U8519 (N_8519,N_8240,N_8158);
nand U8520 (N_8520,N_8398,N_8485);
nor U8521 (N_8521,N_8186,N_8115);
nor U8522 (N_8522,N_8114,N_8310);
and U8523 (N_8523,N_8205,N_8373);
nor U8524 (N_8524,N_8038,N_8128);
nand U8525 (N_8525,N_8064,N_8212);
or U8526 (N_8526,N_8157,N_8391);
and U8527 (N_8527,N_8371,N_8294);
xnor U8528 (N_8528,N_8345,N_8125);
nor U8529 (N_8529,N_8340,N_8027);
and U8530 (N_8530,N_8007,N_8136);
or U8531 (N_8531,N_8089,N_8491);
or U8532 (N_8532,N_8208,N_8261);
nor U8533 (N_8533,N_8000,N_8321);
and U8534 (N_8534,N_8394,N_8036);
and U8535 (N_8535,N_8399,N_8168);
and U8536 (N_8536,N_8484,N_8381);
or U8537 (N_8537,N_8194,N_8293);
nor U8538 (N_8538,N_8182,N_8101);
nand U8539 (N_8539,N_8302,N_8035);
nand U8540 (N_8540,N_8275,N_8059);
or U8541 (N_8541,N_8436,N_8231);
or U8542 (N_8542,N_8370,N_8328);
or U8543 (N_8543,N_8057,N_8303);
nand U8544 (N_8544,N_8113,N_8392);
nor U8545 (N_8545,N_8017,N_8311);
or U8546 (N_8546,N_8228,N_8452);
nor U8547 (N_8547,N_8160,N_8276);
or U8548 (N_8548,N_8496,N_8141);
or U8549 (N_8549,N_8419,N_8230);
nand U8550 (N_8550,N_8033,N_8469);
xnor U8551 (N_8551,N_8030,N_8226);
nor U8552 (N_8552,N_8428,N_8433);
nand U8553 (N_8553,N_8164,N_8331);
nor U8554 (N_8554,N_8424,N_8435);
xnor U8555 (N_8555,N_8074,N_8439);
or U8556 (N_8556,N_8178,N_8325);
and U8557 (N_8557,N_8430,N_8122);
and U8558 (N_8558,N_8449,N_8010);
nor U8559 (N_8559,N_8172,N_8404);
nand U8560 (N_8560,N_8471,N_8129);
nand U8561 (N_8561,N_8247,N_8137);
and U8562 (N_8562,N_8009,N_8354);
nand U8563 (N_8563,N_8227,N_8350);
nor U8564 (N_8564,N_8197,N_8080);
nor U8565 (N_8565,N_8118,N_8183);
or U8566 (N_8566,N_8062,N_8042);
nand U8567 (N_8567,N_8420,N_8324);
or U8568 (N_8568,N_8286,N_8397);
nor U8569 (N_8569,N_8191,N_8029);
or U8570 (N_8570,N_8117,N_8234);
nor U8571 (N_8571,N_8130,N_8289);
and U8572 (N_8572,N_8265,N_8237);
or U8573 (N_8573,N_8049,N_8317);
nand U8574 (N_8574,N_8020,N_8065);
nor U8575 (N_8575,N_8123,N_8039);
and U8576 (N_8576,N_8329,N_8225);
and U8577 (N_8577,N_8002,N_8463);
xnor U8578 (N_8578,N_8330,N_8425);
nand U8579 (N_8579,N_8268,N_8140);
nand U8580 (N_8580,N_8292,N_8283);
nand U8581 (N_8581,N_8159,N_8367);
nand U8582 (N_8582,N_8187,N_8429);
nand U8583 (N_8583,N_8104,N_8335);
or U8584 (N_8584,N_8377,N_8024);
nand U8585 (N_8585,N_8405,N_8127);
xnor U8586 (N_8586,N_8110,N_8264);
nand U8587 (N_8587,N_8400,N_8412);
nand U8588 (N_8588,N_8440,N_8266);
or U8589 (N_8589,N_8387,N_8073);
and U8590 (N_8590,N_8190,N_8426);
or U8591 (N_8591,N_8072,N_8103);
nor U8592 (N_8592,N_8043,N_8132);
or U8593 (N_8593,N_8019,N_8041);
nor U8594 (N_8594,N_8344,N_8006);
or U8595 (N_8595,N_8384,N_8455);
and U8596 (N_8596,N_8409,N_8095);
xor U8597 (N_8597,N_8309,N_8219);
nand U8598 (N_8598,N_8492,N_8477);
nor U8599 (N_8599,N_8166,N_8063);
and U8600 (N_8600,N_8213,N_8393);
nor U8601 (N_8601,N_8150,N_8075);
nand U8602 (N_8602,N_8218,N_8195);
or U8603 (N_8603,N_8388,N_8209);
nand U8604 (N_8604,N_8083,N_8094);
nor U8605 (N_8605,N_8280,N_8107);
or U8606 (N_8606,N_8386,N_8061);
and U8607 (N_8607,N_8028,N_8383);
and U8608 (N_8608,N_8413,N_8044);
and U8609 (N_8609,N_8034,N_8327);
or U8610 (N_8610,N_8479,N_8277);
nand U8611 (N_8611,N_8380,N_8215);
and U8612 (N_8612,N_8198,N_8416);
nand U8613 (N_8613,N_8336,N_8221);
nand U8614 (N_8614,N_8259,N_8018);
nor U8615 (N_8615,N_8406,N_8224);
or U8616 (N_8616,N_8076,N_8222);
nand U8617 (N_8617,N_8288,N_8304);
and U8618 (N_8618,N_8233,N_8053);
xor U8619 (N_8619,N_8274,N_8106);
or U8620 (N_8620,N_8116,N_8427);
and U8621 (N_8621,N_8047,N_8483);
nor U8622 (N_8622,N_8284,N_8023);
or U8623 (N_8623,N_8348,N_8148);
nor U8624 (N_8624,N_8097,N_8055);
nor U8625 (N_8625,N_8100,N_8423);
or U8626 (N_8626,N_8188,N_8249);
and U8627 (N_8627,N_8179,N_8408);
nand U8628 (N_8628,N_8177,N_8184);
and U8629 (N_8629,N_8378,N_8003);
nor U8630 (N_8630,N_8295,N_8472);
or U8631 (N_8631,N_8056,N_8180);
nand U8632 (N_8632,N_8480,N_8453);
nor U8633 (N_8633,N_8096,N_8138);
xnor U8634 (N_8634,N_8014,N_8086);
nand U8635 (N_8635,N_8352,N_8488);
nand U8636 (N_8636,N_8372,N_8454);
or U8637 (N_8637,N_8156,N_8088);
and U8638 (N_8638,N_8342,N_8238);
nor U8639 (N_8639,N_8490,N_8422);
and U8640 (N_8640,N_8257,N_8279);
nand U8641 (N_8641,N_8374,N_8263);
nor U8642 (N_8642,N_8456,N_8058);
and U8643 (N_8643,N_8353,N_8313);
xnor U8644 (N_8644,N_8470,N_8478);
or U8645 (N_8645,N_8270,N_8390);
nand U8646 (N_8646,N_8175,N_8099);
nand U8647 (N_8647,N_8181,N_8012);
and U8648 (N_8648,N_8048,N_8216);
nand U8649 (N_8649,N_8307,N_8458);
nor U8650 (N_8650,N_8193,N_8121);
or U8651 (N_8651,N_8031,N_8133);
nand U8652 (N_8652,N_8446,N_8487);
or U8653 (N_8653,N_8332,N_8369);
nor U8654 (N_8654,N_8206,N_8026);
or U8655 (N_8655,N_8272,N_8203);
xor U8656 (N_8656,N_8414,N_8447);
or U8657 (N_8657,N_8253,N_8199);
nand U8658 (N_8658,N_8068,N_8364);
nor U8659 (N_8659,N_8252,N_8153);
nor U8660 (N_8660,N_8403,N_8432);
and U8661 (N_8661,N_8437,N_8155);
or U8662 (N_8662,N_8069,N_8498);
nor U8663 (N_8663,N_8442,N_8251);
or U8664 (N_8664,N_8319,N_8382);
or U8665 (N_8665,N_8109,N_8001);
nor U8666 (N_8666,N_8267,N_8296);
nand U8667 (N_8667,N_8451,N_8356);
nor U8668 (N_8668,N_8462,N_8385);
or U8669 (N_8669,N_8337,N_8468);
and U8670 (N_8670,N_8476,N_8154);
or U8671 (N_8671,N_8131,N_8375);
nor U8672 (N_8672,N_8464,N_8473);
nand U8673 (N_8673,N_8152,N_8102);
nand U8674 (N_8674,N_8201,N_8050);
and U8675 (N_8675,N_8474,N_8347);
or U8676 (N_8676,N_8376,N_8448);
and U8677 (N_8677,N_8441,N_8411);
xnor U8678 (N_8678,N_8396,N_8489);
and U8679 (N_8679,N_8163,N_8300);
nor U8680 (N_8680,N_8333,N_8084);
nand U8681 (N_8681,N_8202,N_8323);
or U8682 (N_8682,N_8025,N_8457);
and U8683 (N_8683,N_8278,N_8410);
nor U8684 (N_8684,N_8021,N_8461);
or U8685 (N_8685,N_8167,N_8431);
nor U8686 (N_8686,N_8322,N_8389);
and U8687 (N_8687,N_8256,N_8149);
and U8688 (N_8688,N_8314,N_8459);
and U8689 (N_8689,N_8407,N_8402);
and U8690 (N_8690,N_8040,N_8070);
nand U8691 (N_8691,N_8365,N_8105);
nand U8692 (N_8692,N_8143,N_8189);
nand U8693 (N_8693,N_8466,N_8450);
nor U8694 (N_8694,N_8475,N_8015);
or U8695 (N_8695,N_8052,N_8067);
or U8696 (N_8696,N_8214,N_8291);
or U8697 (N_8697,N_8361,N_8022);
nand U8698 (N_8698,N_8290,N_8287);
nand U8699 (N_8699,N_8262,N_8091);
and U8700 (N_8700,N_8162,N_8418);
nand U8701 (N_8701,N_8417,N_8229);
nor U8702 (N_8702,N_8134,N_8349);
nor U8703 (N_8703,N_8243,N_8443);
nand U8704 (N_8704,N_8481,N_8235);
and U8705 (N_8705,N_8093,N_8046);
nand U8706 (N_8706,N_8355,N_8200);
or U8707 (N_8707,N_8255,N_8499);
nor U8708 (N_8708,N_8242,N_8269);
nand U8709 (N_8709,N_8220,N_8165);
nor U8710 (N_8710,N_8297,N_8120);
or U8711 (N_8711,N_8245,N_8357);
nor U8712 (N_8712,N_8079,N_8011);
and U8713 (N_8713,N_8169,N_8082);
or U8714 (N_8714,N_8495,N_8077);
nor U8715 (N_8715,N_8338,N_8486);
nand U8716 (N_8716,N_8146,N_8421);
and U8717 (N_8717,N_8013,N_8087);
nor U8718 (N_8718,N_8111,N_8173);
and U8719 (N_8719,N_8004,N_8444);
xnor U8720 (N_8720,N_8078,N_8250);
or U8721 (N_8721,N_8298,N_8363);
or U8722 (N_8722,N_8318,N_8395);
nor U8723 (N_8723,N_8054,N_8037);
and U8724 (N_8724,N_8326,N_8301);
nor U8725 (N_8725,N_8112,N_8204);
and U8726 (N_8726,N_8341,N_8032);
nor U8727 (N_8727,N_8497,N_8415);
or U8728 (N_8728,N_8285,N_8092);
nor U8729 (N_8729,N_8306,N_8248);
nand U8730 (N_8730,N_8351,N_8174);
nand U8731 (N_8731,N_8460,N_8346);
or U8732 (N_8732,N_8192,N_8085);
nor U8733 (N_8733,N_8170,N_8362);
or U8734 (N_8734,N_8207,N_8312);
and U8735 (N_8735,N_8339,N_8260);
nand U8736 (N_8736,N_8467,N_8258);
and U8737 (N_8737,N_8005,N_8210);
nor U8738 (N_8738,N_8060,N_8139);
and U8739 (N_8739,N_8217,N_8379);
or U8740 (N_8740,N_8008,N_8401);
xor U8741 (N_8741,N_8334,N_8211);
and U8742 (N_8742,N_8239,N_8090);
or U8743 (N_8743,N_8282,N_8241);
nor U8744 (N_8744,N_8176,N_8358);
nor U8745 (N_8745,N_8244,N_8071);
and U8746 (N_8746,N_8145,N_8151);
or U8747 (N_8747,N_8124,N_8144);
nand U8748 (N_8748,N_8299,N_8135);
nand U8749 (N_8749,N_8315,N_8066);
and U8750 (N_8750,N_8216,N_8347);
or U8751 (N_8751,N_8045,N_8472);
nand U8752 (N_8752,N_8389,N_8339);
xnor U8753 (N_8753,N_8110,N_8449);
and U8754 (N_8754,N_8217,N_8110);
or U8755 (N_8755,N_8370,N_8307);
xnor U8756 (N_8756,N_8263,N_8282);
nand U8757 (N_8757,N_8307,N_8095);
and U8758 (N_8758,N_8053,N_8129);
nand U8759 (N_8759,N_8307,N_8302);
nor U8760 (N_8760,N_8433,N_8368);
xnor U8761 (N_8761,N_8147,N_8247);
or U8762 (N_8762,N_8218,N_8499);
nor U8763 (N_8763,N_8060,N_8101);
nor U8764 (N_8764,N_8329,N_8137);
nor U8765 (N_8765,N_8392,N_8443);
nor U8766 (N_8766,N_8056,N_8297);
nand U8767 (N_8767,N_8081,N_8394);
or U8768 (N_8768,N_8285,N_8131);
nand U8769 (N_8769,N_8297,N_8007);
or U8770 (N_8770,N_8162,N_8060);
and U8771 (N_8771,N_8352,N_8379);
nand U8772 (N_8772,N_8096,N_8060);
nand U8773 (N_8773,N_8029,N_8489);
nor U8774 (N_8774,N_8102,N_8352);
or U8775 (N_8775,N_8209,N_8177);
nor U8776 (N_8776,N_8473,N_8033);
and U8777 (N_8777,N_8207,N_8467);
or U8778 (N_8778,N_8061,N_8325);
nand U8779 (N_8779,N_8281,N_8424);
or U8780 (N_8780,N_8276,N_8482);
nor U8781 (N_8781,N_8334,N_8126);
or U8782 (N_8782,N_8267,N_8472);
and U8783 (N_8783,N_8459,N_8222);
nor U8784 (N_8784,N_8126,N_8262);
or U8785 (N_8785,N_8429,N_8448);
nor U8786 (N_8786,N_8185,N_8079);
and U8787 (N_8787,N_8084,N_8469);
nand U8788 (N_8788,N_8361,N_8135);
and U8789 (N_8789,N_8127,N_8052);
nand U8790 (N_8790,N_8357,N_8460);
or U8791 (N_8791,N_8248,N_8054);
or U8792 (N_8792,N_8439,N_8151);
nand U8793 (N_8793,N_8001,N_8459);
nor U8794 (N_8794,N_8414,N_8390);
nor U8795 (N_8795,N_8193,N_8116);
and U8796 (N_8796,N_8428,N_8282);
nor U8797 (N_8797,N_8262,N_8185);
and U8798 (N_8798,N_8298,N_8187);
and U8799 (N_8799,N_8012,N_8007);
and U8800 (N_8800,N_8011,N_8331);
and U8801 (N_8801,N_8013,N_8200);
xnor U8802 (N_8802,N_8470,N_8372);
nor U8803 (N_8803,N_8244,N_8004);
and U8804 (N_8804,N_8025,N_8266);
and U8805 (N_8805,N_8007,N_8406);
and U8806 (N_8806,N_8013,N_8125);
or U8807 (N_8807,N_8127,N_8237);
nor U8808 (N_8808,N_8058,N_8474);
nor U8809 (N_8809,N_8359,N_8324);
or U8810 (N_8810,N_8484,N_8428);
nor U8811 (N_8811,N_8067,N_8161);
and U8812 (N_8812,N_8488,N_8319);
nand U8813 (N_8813,N_8258,N_8030);
nor U8814 (N_8814,N_8077,N_8157);
nand U8815 (N_8815,N_8237,N_8104);
and U8816 (N_8816,N_8463,N_8363);
or U8817 (N_8817,N_8337,N_8206);
or U8818 (N_8818,N_8072,N_8353);
and U8819 (N_8819,N_8230,N_8453);
nor U8820 (N_8820,N_8470,N_8084);
or U8821 (N_8821,N_8274,N_8440);
nand U8822 (N_8822,N_8319,N_8225);
or U8823 (N_8823,N_8383,N_8363);
nand U8824 (N_8824,N_8030,N_8175);
nor U8825 (N_8825,N_8344,N_8127);
or U8826 (N_8826,N_8096,N_8169);
nor U8827 (N_8827,N_8239,N_8017);
nand U8828 (N_8828,N_8420,N_8149);
nor U8829 (N_8829,N_8341,N_8069);
and U8830 (N_8830,N_8220,N_8483);
and U8831 (N_8831,N_8097,N_8290);
and U8832 (N_8832,N_8484,N_8447);
nand U8833 (N_8833,N_8350,N_8308);
and U8834 (N_8834,N_8210,N_8371);
or U8835 (N_8835,N_8277,N_8211);
and U8836 (N_8836,N_8430,N_8240);
or U8837 (N_8837,N_8268,N_8232);
nand U8838 (N_8838,N_8366,N_8166);
and U8839 (N_8839,N_8374,N_8245);
nor U8840 (N_8840,N_8260,N_8193);
and U8841 (N_8841,N_8010,N_8398);
nand U8842 (N_8842,N_8029,N_8497);
or U8843 (N_8843,N_8000,N_8423);
and U8844 (N_8844,N_8103,N_8309);
nand U8845 (N_8845,N_8239,N_8068);
and U8846 (N_8846,N_8475,N_8133);
and U8847 (N_8847,N_8326,N_8113);
or U8848 (N_8848,N_8298,N_8045);
nand U8849 (N_8849,N_8055,N_8284);
nor U8850 (N_8850,N_8002,N_8312);
or U8851 (N_8851,N_8232,N_8489);
or U8852 (N_8852,N_8275,N_8318);
and U8853 (N_8853,N_8342,N_8166);
and U8854 (N_8854,N_8383,N_8324);
nand U8855 (N_8855,N_8046,N_8003);
and U8856 (N_8856,N_8408,N_8157);
nor U8857 (N_8857,N_8222,N_8310);
or U8858 (N_8858,N_8116,N_8391);
and U8859 (N_8859,N_8388,N_8159);
or U8860 (N_8860,N_8198,N_8441);
or U8861 (N_8861,N_8376,N_8154);
and U8862 (N_8862,N_8366,N_8480);
and U8863 (N_8863,N_8497,N_8393);
or U8864 (N_8864,N_8186,N_8187);
and U8865 (N_8865,N_8435,N_8194);
nor U8866 (N_8866,N_8238,N_8130);
or U8867 (N_8867,N_8273,N_8051);
or U8868 (N_8868,N_8352,N_8460);
or U8869 (N_8869,N_8467,N_8400);
or U8870 (N_8870,N_8400,N_8092);
nand U8871 (N_8871,N_8261,N_8292);
or U8872 (N_8872,N_8371,N_8288);
and U8873 (N_8873,N_8218,N_8224);
or U8874 (N_8874,N_8101,N_8271);
or U8875 (N_8875,N_8001,N_8479);
or U8876 (N_8876,N_8445,N_8120);
nand U8877 (N_8877,N_8398,N_8202);
nand U8878 (N_8878,N_8012,N_8308);
or U8879 (N_8879,N_8174,N_8255);
and U8880 (N_8880,N_8223,N_8247);
nor U8881 (N_8881,N_8369,N_8471);
nor U8882 (N_8882,N_8352,N_8191);
xor U8883 (N_8883,N_8355,N_8344);
nor U8884 (N_8884,N_8163,N_8271);
or U8885 (N_8885,N_8302,N_8029);
nor U8886 (N_8886,N_8412,N_8293);
and U8887 (N_8887,N_8025,N_8247);
xor U8888 (N_8888,N_8489,N_8095);
or U8889 (N_8889,N_8099,N_8410);
or U8890 (N_8890,N_8271,N_8228);
nor U8891 (N_8891,N_8223,N_8420);
and U8892 (N_8892,N_8153,N_8386);
or U8893 (N_8893,N_8468,N_8214);
or U8894 (N_8894,N_8066,N_8441);
or U8895 (N_8895,N_8142,N_8460);
or U8896 (N_8896,N_8385,N_8041);
nor U8897 (N_8897,N_8156,N_8397);
and U8898 (N_8898,N_8234,N_8454);
nor U8899 (N_8899,N_8407,N_8364);
nor U8900 (N_8900,N_8095,N_8191);
nor U8901 (N_8901,N_8082,N_8305);
or U8902 (N_8902,N_8373,N_8097);
and U8903 (N_8903,N_8262,N_8379);
and U8904 (N_8904,N_8214,N_8426);
or U8905 (N_8905,N_8189,N_8117);
and U8906 (N_8906,N_8210,N_8410);
and U8907 (N_8907,N_8203,N_8228);
or U8908 (N_8908,N_8404,N_8379);
xnor U8909 (N_8909,N_8158,N_8316);
and U8910 (N_8910,N_8030,N_8373);
nor U8911 (N_8911,N_8423,N_8175);
nand U8912 (N_8912,N_8329,N_8209);
nand U8913 (N_8913,N_8042,N_8193);
nand U8914 (N_8914,N_8299,N_8406);
or U8915 (N_8915,N_8190,N_8237);
nor U8916 (N_8916,N_8278,N_8357);
nor U8917 (N_8917,N_8460,N_8009);
and U8918 (N_8918,N_8483,N_8315);
nor U8919 (N_8919,N_8013,N_8177);
nor U8920 (N_8920,N_8477,N_8097);
and U8921 (N_8921,N_8287,N_8193);
and U8922 (N_8922,N_8310,N_8363);
nor U8923 (N_8923,N_8390,N_8394);
nor U8924 (N_8924,N_8472,N_8377);
or U8925 (N_8925,N_8228,N_8277);
nor U8926 (N_8926,N_8087,N_8340);
or U8927 (N_8927,N_8456,N_8084);
or U8928 (N_8928,N_8120,N_8220);
and U8929 (N_8929,N_8382,N_8448);
or U8930 (N_8930,N_8359,N_8446);
and U8931 (N_8931,N_8497,N_8025);
or U8932 (N_8932,N_8254,N_8221);
xor U8933 (N_8933,N_8447,N_8145);
or U8934 (N_8934,N_8022,N_8348);
nand U8935 (N_8935,N_8367,N_8390);
and U8936 (N_8936,N_8137,N_8313);
and U8937 (N_8937,N_8147,N_8180);
and U8938 (N_8938,N_8357,N_8356);
nand U8939 (N_8939,N_8447,N_8277);
nor U8940 (N_8940,N_8286,N_8304);
and U8941 (N_8941,N_8387,N_8313);
and U8942 (N_8942,N_8030,N_8349);
and U8943 (N_8943,N_8313,N_8029);
nand U8944 (N_8944,N_8068,N_8019);
nor U8945 (N_8945,N_8297,N_8410);
and U8946 (N_8946,N_8499,N_8059);
and U8947 (N_8947,N_8117,N_8467);
nand U8948 (N_8948,N_8223,N_8028);
and U8949 (N_8949,N_8095,N_8368);
or U8950 (N_8950,N_8052,N_8013);
and U8951 (N_8951,N_8322,N_8258);
nand U8952 (N_8952,N_8005,N_8336);
or U8953 (N_8953,N_8439,N_8104);
and U8954 (N_8954,N_8002,N_8374);
or U8955 (N_8955,N_8129,N_8351);
or U8956 (N_8956,N_8112,N_8044);
nor U8957 (N_8957,N_8407,N_8317);
nand U8958 (N_8958,N_8415,N_8029);
nand U8959 (N_8959,N_8151,N_8064);
nor U8960 (N_8960,N_8422,N_8480);
nor U8961 (N_8961,N_8305,N_8440);
nand U8962 (N_8962,N_8234,N_8161);
nor U8963 (N_8963,N_8472,N_8302);
or U8964 (N_8964,N_8200,N_8049);
or U8965 (N_8965,N_8083,N_8222);
nand U8966 (N_8966,N_8425,N_8015);
and U8967 (N_8967,N_8359,N_8109);
nand U8968 (N_8968,N_8080,N_8044);
or U8969 (N_8969,N_8489,N_8187);
nor U8970 (N_8970,N_8074,N_8206);
nor U8971 (N_8971,N_8451,N_8010);
nor U8972 (N_8972,N_8174,N_8298);
nor U8973 (N_8973,N_8348,N_8172);
nand U8974 (N_8974,N_8219,N_8125);
and U8975 (N_8975,N_8026,N_8198);
and U8976 (N_8976,N_8447,N_8453);
nor U8977 (N_8977,N_8222,N_8253);
and U8978 (N_8978,N_8344,N_8484);
and U8979 (N_8979,N_8044,N_8464);
or U8980 (N_8980,N_8027,N_8402);
and U8981 (N_8981,N_8009,N_8262);
and U8982 (N_8982,N_8076,N_8008);
and U8983 (N_8983,N_8405,N_8228);
nand U8984 (N_8984,N_8042,N_8421);
nand U8985 (N_8985,N_8267,N_8000);
and U8986 (N_8986,N_8019,N_8118);
nor U8987 (N_8987,N_8258,N_8407);
and U8988 (N_8988,N_8414,N_8215);
or U8989 (N_8989,N_8283,N_8062);
nand U8990 (N_8990,N_8217,N_8022);
nor U8991 (N_8991,N_8376,N_8201);
nand U8992 (N_8992,N_8299,N_8478);
nand U8993 (N_8993,N_8239,N_8392);
or U8994 (N_8994,N_8268,N_8426);
nor U8995 (N_8995,N_8259,N_8427);
nor U8996 (N_8996,N_8115,N_8207);
and U8997 (N_8997,N_8033,N_8349);
nor U8998 (N_8998,N_8308,N_8400);
nand U8999 (N_8999,N_8494,N_8076);
or U9000 (N_9000,N_8999,N_8509);
or U9001 (N_9001,N_8615,N_8876);
nor U9002 (N_9002,N_8961,N_8755);
and U9003 (N_9003,N_8545,N_8942);
or U9004 (N_9004,N_8874,N_8846);
or U9005 (N_9005,N_8949,N_8866);
or U9006 (N_9006,N_8782,N_8665);
nor U9007 (N_9007,N_8929,N_8784);
and U9008 (N_9008,N_8761,N_8579);
xnor U9009 (N_9009,N_8620,N_8713);
nand U9010 (N_9010,N_8558,N_8610);
or U9011 (N_9011,N_8669,N_8679);
xor U9012 (N_9012,N_8760,N_8756);
or U9013 (N_9013,N_8724,N_8625);
nor U9014 (N_9014,N_8847,N_8611);
and U9015 (N_9015,N_8834,N_8879);
nor U9016 (N_9016,N_8712,N_8648);
xnor U9017 (N_9017,N_8729,N_8740);
nor U9018 (N_9018,N_8593,N_8616);
nand U9019 (N_9019,N_8897,N_8886);
or U9020 (N_9020,N_8766,N_8551);
and U9021 (N_9021,N_8563,N_8829);
or U9022 (N_9022,N_8797,N_8550);
or U9023 (N_9023,N_8697,N_8916);
nand U9024 (N_9024,N_8749,N_8681);
or U9025 (N_9025,N_8612,N_8747);
and U9026 (N_9026,N_8895,N_8944);
nand U9027 (N_9027,N_8753,N_8867);
nor U9028 (N_9028,N_8900,N_8642);
nor U9029 (N_9029,N_8991,N_8792);
nand U9030 (N_9030,N_8614,N_8621);
and U9031 (N_9031,N_8704,N_8532);
or U9032 (N_9032,N_8793,N_8746);
or U9033 (N_9033,N_8561,N_8696);
and U9034 (N_9034,N_8631,N_8959);
or U9035 (N_9035,N_8833,N_8733);
nor U9036 (N_9036,N_8820,N_8940);
or U9037 (N_9037,N_8607,N_8739);
and U9038 (N_9038,N_8645,N_8664);
nand U9039 (N_9039,N_8513,N_8599);
nor U9040 (N_9040,N_8741,N_8884);
or U9041 (N_9041,N_8933,N_8653);
nor U9042 (N_9042,N_8960,N_8915);
and U9043 (N_9043,N_8514,N_8587);
or U9044 (N_9044,N_8821,N_8913);
and U9045 (N_9045,N_8971,N_8844);
and U9046 (N_9046,N_8718,N_8768);
or U9047 (N_9047,N_8671,N_8955);
xnor U9048 (N_9048,N_8994,N_8535);
or U9049 (N_9049,N_8723,N_8938);
and U9050 (N_9050,N_8810,N_8591);
nor U9051 (N_9051,N_8525,N_8826);
nor U9052 (N_9052,N_8928,N_8606);
or U9053 (N_9053,N_8996,N_8619);
nor U9054 (N_9054,N_8809,N_8727);
nand U9055 (N_9055,N_8717,N_8564);
and U9056 (N_9056,N_8780,N_8685);
or U9057 (N_9057,N_8978,N_8658);
or U9058 (N_9058,N_8629,N_8689);
or U9059 (N_9059,N_8701,N_8974);
nand U9060 (N_9060,N_8919,N_8817);
or U9061 (N_9061,N_8730,N_8888);
nor U9062 (N_9062,N_8835,N_8993);
and U9063 (N_9063,N_8666,N_8524);
or U9064 (N_9064,N_8641,N_8774);
or U9065 (N_9065,N_8802,N_8646);
and U9066 (N_9066,N_8904,N_8995);
nand U9067 (N_9067,N_8649,N_8601);
or U9068 (N_9068,N_8586,N_8630);
nor U9069 (N_9069,N_8813,N_8636);
or U9070 (N_9070,N_8687,N_8815);
nand U9071 (N_9071,N_8530,N_8818);
and U9072 (N_9072,N_8538,N_8863);
or U9073 (N_9073,N_8673,N_8592);
and U9074 (N_9074,N_8853,N_8602);
nor U9075 (N_9075,N_8757,N_8656);
nor U9076 (N_9076,N_8751,N_8667);
nor U9077 (N_9077,N_8855,N_8603);
nand U9078 (N_9078,N_8703,N_8738);
nor U9079 (N_9079,N_8506,N_8907);
and U9080 (N_9080,N_8767,N_8519);
nand U9081 (N_9081,N_8883,N_8778);
or U9082 (N_9082,N_8931,N_8790);
or U9083 (N_9083,N_8504,N_8546);
or U9084 (N_9084,N_8568,N_8644);
and U9085 (N_9085,N_8585,N_8939);
and U9086 (N_9086,N_8662,N_8507);
nand U9087 (N_9087,N_8981,N_8694);
nand U9088 (N_9088,N_8677,N_8577);
nand U9089 (N_9089,N_8565,N_8922);
or U9090 (N_9090,N_8805,N_8698);
nand U9091 (N_9091,N_8952,N_8908);
nor U9092 (N_9092,N_8663,N_8567);
and U9093 (N_9093,N_8700,N_8901);
xnor U9094 (N_9094,N_8789,N_8594);
nand U9095 (N_9095,N_8762,N_8882);
or U9096 (N_9096,N_8770,N_8911);
or U9097 (N_9097,N_8896,N_8754);
nand U9098 (N_9098,N_8923,N_8927);
nor U9099 (N_9099,N_8804,N_8779);
and U9100 (N_9100,N_8984,N_8880);
nand U9101 (N_9101,N_8559,N_8693);
or U9102 (N_9102,N_8634,N_8893);
nand U9103 (N_9103,N_8652,N_8842);
and U9104 (N_9104,N_8576,N_8950);
nor U9105 (N_9105,N_8722,N_8869);
nor U9106 (N_9106,N_8914,N_8973);
or U9107 (N_9107,N_8589,N_8726);
and U9108 (N_9108,N_8720,N_8572);
or U9109 (N_9109,N_8951,N_8848);
nor U9110 (N_9110,N_8676,N_8597);
or U9111 (N_9111,N_8580,N_8500);
and U9112 (N_9112,N_8831,N_8906);
nand U9113 (N_9113,N_8806,N_8573);
nor U9114 (N_9114,N_8544,N_8966);
xnor U9115 (N_9115,N_8654,N_8985);
nor U9116 (N_9116,N_8800,N_8533);
nor U9117 (N_9117,N_8877,N_8871);
nand U9118 (N_9118,N_8773,N_8811);
nand U9119 (N_9119,N_8547,N_8788);
xnor U9120 (N_9120,N_8643,N_8997);
and U9121 (N_9121,N_8517,N_8691);
and U9122 (N_9122,N_8632,N_8858);
and U9123 (N_9123,N_8958,N_8571);
or U9124 (N_9124,N_8975,N_8998);
nand U9125 (N_9125,N_8976,N_8521);
nor U9126 (N_9126,N_8627,N_8548);
and U9127 (N_9127,N_8881,N_8988);
or U9128 (N_9128,N_8542,N_8684);
nand U9129 (N_9129,N_8537,N_8925);
nor U9130 (N_9130,N_8794,N_8859);
nor U9131 (N_9131,N_8633,N_8543);
and U9132 (N_9132,N_8609,N_8736);
nand U9133 (N_9133,N_8783,N_8735);
nand U9134 (N_9134,N_8803,N_8699);
or U9135 (N_9135,N_8678,N_8702);
nand U9136 (N_9136,N_8775,N_8716);
nor U9137 (N_9137,N_8752,N_8801);
nor U9138 (N_9138,N_8661,N_8967);
and U9139 (N_9139,N_8989,N_8682);
or U9140 (N_9140,N_8552,N_8851);
xnor U9141 (N_9141,N_8977,N_8865);
and U9142 (N_9142,N_8972,N_8854);
nor U9143 (N_9143,N_8868,N_8771);
and U9144 (N_9144,N_8557,N_8737);
and U9145 (N_9145,N_8711,N_8536);
nand U9146 (N_9146,N_8920,N_8909);
nand U9147 (N_9147,N_8839,N_8979);
nand U9148 (N_9148,N_8516,N_8732);
and U9149 (N_9149,N_8680,N_8843);
and U9150 (N_9150,N_8814,N_8605);
and U9151 (N_9151,N_8980,N_8828);
nand U9152 (N_9152,N_8743,N_8921);
nor U9153 (N_9153,N_8719,N_8742);
nor U9154 (N_9154,N_8744,N_8934);
nor U9155 (N_9155,N_8791,N_8864);
and U9156 (N_9156,N_8710,N_8894);
nor U9157 (N_9157,N_8651,N_8690);
and U9158 (N_9158,N_8520,N_8917);
nand U9159 (N_9159,N_8655,N_8556);
and U9160 (N_9160,N_8992,N_8553);
and U9161 (N_9161,N_8841,N_8964);
and U9162 (N_9162,N_8891,N_8595);
and U9163 (N_9163,N_8637,N_8941);
nor U9164 (N_9164,N_8709,N_8890);
nand U9165 (N_9165,N_8945,N_8872);
and U9166 (N_9166,N_8969,N_8860);
and U9167 (N_9167,N_8758,N_8541);
nand U9168 (N_9168,N_8512,N_8786);
and U9169 (N_9169,N_8617,N_8776);
and U9170 (N_9170,N_8903,N_8708);
nand U9171 (N_9171,N_8849,N_8707);
and U9172 (N_9172,N_8787,N_8598);
or U9173 (N_9173,N_8511,N_8832);
and U9174 (N_9174,N_8613,N_8745);
and U9175 (N_9175,N_8777,N_8837);
nor U9176 (N_9176,N_8918,N_8808);
and U9177 (N_9177,N_8902,N_8845);
nand U9178 (N_9178,N_8824,N_8725);
nor U9179 (N_9179,N_8954,N_8638);
or U9180 (N_9180,N_8628,N_8892);
nand U9181 (N_9181,N_8785,N_8554);
and U9182 (N_9182,N_8668,N_8657);
or U9183 (N_9183,N_8956,N_8600);
nand U9184 (N_9184,N_8836,N_8695);
nand U9185 (N_9185,N_8584,N_8947);
and U9186 (N_9186,N_8990,N_8987);
and U9187 (N_9187,N_8948,N_8604);
nor U9188 (N_9188,N_8731,N_8721);
and U9189 (N_9189,N_8639,N_8965);
nor U9190 (N_9190,N_8937,N_8924);
nor U9191 (N_9191,N_8798,N_8986);
and U9192 (N_9192,N_8518,N_8870);
nand U9193 (N_9193,N_8982,N_8968);
or U9194 (N_9194,N_8807,N_8596);
or U9195 (N_9195,N_8728,N_8852);
nand U9196 (N_9196,N_8527,N_8574);
and U9197 (N_9197,N_8930,N_8588);
or U9198 (N_9198,N_8608,N_8623);
nor U9199 (N_9199,N_8622,N_8674);
nand U9200 (N_9200,N_8799,N_8822);
and U9201 (N_9201,N_8932,N_8873);
and U9202 (N_9202,N_8759,N_8825);
and U9203 (N_9203,N_8715,N_8899);
xnor U9204 (N_9204,N_8560,N_8531);
nand U9205 (N_9205,N_8523,N_8878);
nand U9206 (N_9206,N_8827,N_8578);
nand U9207 (N_9207,N_8659,N_8692);
nand U9208 (N_9208,N_8624,N_8626);
and U9209 (N_9209,N_8887,N_8660);
nand U9210 (N_9210,N_8823,N_8812);
or U9211 (N_9211,N_8926,N_8816);
or U9212 (N_9212,N_8983,N_8857);
nand U9213 (N_9213,N_8686,N_8583);
nor U9214 (N_9214,N_8570,N_8970);
or U9215 (N_9215,N_8898,N_8943);
or U9216 (N_9216,N_8582,N_8526);
and U9217 (N_9217,N_8910,N_8840);
nand U9218 (N_9218,N_8562,N_8515);
nor U9219 (N_9219,N_8688,N_8885);
nor U9220 (N_9220,N_8647,N_8946);
or U9221 (N_9221,N_8675,N_8750);
and U9222 (N_9222,N_8781,N_8534);
nand U9223 (N_9223,N_8905,N_8555);
and U9224 (N_9224,N_8763,N_8838);
nand U9225 (N_9225,N_8963,N_8635);
and U9226 (N_9226,N_8830,N_8539);
and U9227 (N_9227,N_8819,N_8590);
nor U9228 (N_9228,N_8503,N_8769);
and U9229 (N_9229,N_8936,N_8772);
nand U9230 (N_9230,N_8889,N_8581);
xnor U9231 (N_9231,N_8764,N_8672);
and U9232 (N_9232,N_8912,N_8529);
xor U9233 (N_9233,N_8549,N_8935);
or U9234 (N_9234,N_8508,N_8953);
nor U9235 (N_9235,N_8650,N_8683);
nand U9236 (N_9236,N_8501,N_8875);
and U9237 (N_9237,N_8522,N_8957);
and U9238 (N_9238,N_8618,N_8705);
and U9239 (N_9239,N_8765,N_8640);
and U9240 (N_9240,N_8510,N_8566);
and U9241 (N_9241,N_8862,N_8795);
nand U9242 (N_9242,N_8575,N_8569);
nor U9243 (N_9243,N_8540,N_8528);
or U9244 (N_9244,N_8706,N_8670);
nor U9245 (N_9245,N_8714,N_8502);
and U9246 (N_9246,N_8748,N_8796);
nor U9247 (N_9247,N_8856,N_8861);
and U9248 (N_9248,N_8505,N_8962);
nor U9249 (N_9249,N_8850,N_8734);
nor U9250 (N_9250,N_8509,N_8827);
xor U9251 (N_9251,N_8880,N_8545);
nand U9252 (N_9252,N_8749,N_8877);
nor U9253 (N_9253,N_8816,N_8916);
nand U9254 (N_9254,N_8906,N_8575);
nand U9255 (N_9255,N_8843,N_8796);
and U9256 (N_9256,N_8596,N_8554);
nor U9257 (N_9257,N_8901,N_8884);
or U9258 (N_9258,N_8579,N_8776);
nand U9259 (N_9259,N_8881,N_8870);
or U9260 (N_9260,N_8611,N_8991);
or U9261 (N_9261,N_8873,N_8756);
nand U9262 (N_9262,N_8511,N_8647);
or U9263 (N_9263,N_8720,N_8894);
nor U9264 (N_9264,N_8551,N_8531);
nor U9265 (N_9265,N_8859,N_8843);
nor U9266 (N_9266,N_8699,N_8725);
nand U9267 (N_9267,N_8527,N_8968);
nand U9268 (N_9268,N_8942,N_8819);
nand U9269 (N_9269,N_8964,N_8704);
and U9270 (N_9270,N_8526,N_8689);
nand U9271 (N_9271,N_8966,N_8708);
or U9272 (N_9272,N_8846,N_8654);
nand U9273 (N_9273,N_8957,N_8535);
nor U9274 (N_9274,N_8614,N_8760);
nor U9275 (N_9275,N_8836,N_8583);
nor U9276 (N_9276,N_8879,N_8640);
and U9277 (N_9277,N_8738,N_8940);
nor U9278 (N_9278,N_8983,N_8555);
nand U9279 (N_9279,N_8510,N_8732);
nand U9280 (N_9280,N_8729,N_8727);
and U9281 (N_9281,N_8583,N_8570);
nand U9282 (N_9282,N_8998,N_8955);
or U9283 (N_9283,N_8802,N_8576);
nor U9284 (N_9284,N_8526,N_8895);
nor U9285 (N_9285,N_8855,N_8534);
and U9286 (N_9286,N_8672,N_8724);
nand U9287 (N_9287,N_8700,N_8591);
and U9288 (N_9288,N_8625,N_8941);
xor U9289 (N_9289,N_8896,N_8841);
nand U9290 (N_9290,N_8958,N_8926);
nor U9291 (N_9291,N_8925,N_8909);
nand U9292 (N_9292,N_8725,N_8785);
or U9293 (N_9293,N_8760,N_8940);
xnor U9294 (N_9294,N_8770,N_8874);
or U9295 (N_9295,N_8803,N_8807);
nand U9296 (N_9296,N_8689,N_8502);
or U9297 (N_9297,N_8548,N_8681);
or U9298 (N_9298,N_8867,N_8534);
nand U9299 (N_9299,N_8571,N_8549);
and U9300 (N_9300,N_8523,N_8723);
and U9301 (N_9301,N_8707,N_8646);
or U9302 (N_9302,N_8562,N_8510);
and U9303 (N_9303,N_8864,N_8555);
nor U9304 (N_9304,N_8509,N_8936);
nor U9305 (N_9305,N_8525,N_8963);
xnor U9306 (N_9306,N_8882,N_8537);
or U9307 (N_9307,N_8962,N_8968);
and U9308 (N_9308,N_8832,N_8856);
nand U9309 (N_9309,N_8649,N_8581);
and U9310 (N_9310,N_8678,N_8872);
nor U9311 (N_9311,N_8632,N_8842);
nand U9312 (N_9312,N_8739,N_8552);
and U9313 (N_9313,N_8652,N_8501);
and U9314 (N_9314,N_8727,N_8903);
nand U9315 (N_9315,N_8826,N_8902);
nor U9316 (N_9316,N_8674,N_8724);
or U9317 (N_9317,N_8637,N_8522);
nand U9318 (N_9318,N_8781,N_8724);
nand U9319 (N_9319,N_8815,N_8824);
nand U9320 (N_9320,N_8828,N_8672);
or U9321 (N_9321,N_8895,N_8729);
and U9322 (N_9322,N_8597,N_8590);
nor U9323 (N_9323,N_8503,N_8876);
nor U9324 (N_9324,N_8863,N_8564);
nor U9325 (N_9325,N_8809,N_8600);
and U9326 (N_9326,N_8929,N_8615);
nor U9327 (N_9327,N_8682,N_8980);
xor U9328 (N_9328,N_8890,N_8608);
or U9329 (N_9329,N_8976,N_8717);
and U9330 (N_9330,N_8912,N_8936);
xnor U9331 (N_9331,N_8548,N_8974);
and U9332 (N_9332,N_8951,N_8585);
or U9333 (N_9333,N_8509,N_8600);
nor U9334 (N_9334,N_8566,N_8888);
and U9335 (N_9335,N_8802,N_8612);
nor U9336 (N_9336,N_8546,N_8700);
or U9337 (N_9337,N_8529,N_8841);
or U9338 (N_9338,N_8578,N_8539);
and U9339 (N_9339,N_8826,N_8567);
nor U9340 (N_9340,N_8980,N_8814);
and U9341 (N_9341,N_8954,N_8571);
or U9342 (N_9342,N_8808,N_8542);
and U9343 (N_9343,N_8710,N_8787);
nand U9344 (N_9344,N_8991,N_8603);
nor U9345 (N_9345,N_8567,N_8719);
nor U9346 (N_9346,N_8876,N_8644);
nor U9347 (N_9347,N_8920,N_8691);
nor U9348 (N_9348,N_8915,N_8589);
nand U9349 (N_9349,N_8907,N_8865);
nand U9350 (N_9350,N_8715,N_8946);
nor U9351 (N_9351,N_8976,N_8881);
nor U9352 (N_9352,N_8649,N_8950);
and U9353 (N_9353,N_8641,N_8506);
and U9354 (N_9354,N_8746,N_8519);
nor U9355 (N_9355,N_8910,N_8615);
or U9356 (N_9356,N_8556,N_8982);
or U9357 (N_9357,N_8504,N_8694);
or U9358 (N_9358,N_8960,N_8551);
nor U9359 (N_9359,N_8596,N_8666);
nand U9360 (N_9360,N_8911,N_8771);
nand U9361 (N_9361,N_8603,N_8821);
or U9362 (N_9362,N_8534,N_8887);
and U9363 (N_9363,N_8634,N_8754);
or U9364 (N_9364,N_8877,N_8991);
nand U9365 (N_9365,N_8957,N_8903);
or U9366 (N_9366,N_8667,N_8598);
nor U9367 (N_9367,N_8569,N_8725);
nor U9368 (N_9368,N_8809,N_8810);
nand U9369 (N_9369,N_8841,N_8998);
nor U9370 (N_9370,N_8852,N_8740);
nand U9371 (N_9371,N_8659,N_8905);
and U9372 (N_9372,N_8929,N_8882);
nand U9373 (N_9373,N_8959,N_8990);
nor U9374 (N_9374,N_8905,N_8906);
nor U9375 (N_9375,N_8955,N_8758);
or U9376 (N_9376,N_8512,N_8687);
or U9377 (N_9377,N_8607,N_8770);
or U9378 (N_9378,N_8870,N_8733);
or U9379 (N_9379,N_8880,N_8698);
or U9380 (N_9380,N_8688,N_8548);
nand U9381 (N_9381,N_8657,N_8938);
nand U9382 (N_9382,N_8669,N_8806);
or U9383 (N_9383,N_8700,N_8614);
nor U9384 (N_9384,N_8694,N_8989);
nand U9385 (N_9385,N_8918,N_8936);
or U9386 (N_9386,N_8694,N_8834);
and U9387 (N_9387,N_8552,N_8644);
and U9388 (N_9388,N_8787,N_8958);
and U9389 (N_9389,N_8731,N_8918);
or U9390 (N_9390,N_8895,N_8580);
nand U9391 (N_9391,N_8656,N_8686);
and U9392 (N_9392,N_8759,N_8643);
or U9393 (N_9393,N_8790,N_8505);
nand U9394 (N_9394,N_8508,N_8813);
or U9395 (N_9395,N_8707,N_8618);
nor U9396 (N_9396,N_8846,N_8912);
and U9397 (N_9397,N_8577,N_8707);
nand U9398 (N_9398,N_8646,N_8959);
nor U9399 (N_9399,N_8558,N_8513);
or U9400 (N_9400,N_8873,N_8684);
nor U9401 (N_9401,N_8990,N_8529);
and U9402 (N_9402,N_8788,N_8944);
nand U9403 (N_9403,N_8848,N_8600);
nor U9404 (N_9404,N_8563,N_8852);
and U9405 (N_9405,N_8825,N_8841);
nand U9406 (N_9406,N_8717,N_8603);
or U9407 (N_9407,N_8643,N_8939);
nor U9408 (N_9408,N_8888,N_8731);
nor U9409 (N_9409,N_8726,N_8757);
or U9410 (N_9410,N_8924,N_8518);
or U9411 (N_9411,N_8993,N_8593);
nand U9412 (N_9412,N_8652,N_8880);
nor U9413 (N_9413,N_8546,N_8833);
nor U9414 (N_9414,N_8809,N_8711);
and U9415 (N_9415,N_8910,N_8721);
nor U9416 (N_9416,N_8669,N_8678);
nor U9417 (N_9417,N_8641,N_8868);
nor U9418 (N_9418,N_8564,N_8891);
or U9419 (N_9419,N_8532,N_8855);
and U9420 (N_9420,N_8800,N_8599);
and U9421 (N_9421,N_8745,N_8714);
nand U9422 (N_9422,N_8945,N_8935);
or U9423 (N_9423,N_8908,N_8529);
or U9424 (N_9424,N_8557,N_8712);
nand U9425 (N_9425,N_8955,N_8819);
nor U9426 (N_9426,N_8995,N_8745);
nor U9427 (N_9427,N_8864,N_8850);
nor U9428 (N_9428,N_8789,N_8664);
nand U9429 (N_9429,N_8646,N_8770);
nand U9430 (N_9430,N_8699,N_8713);
and U9431 (N_9431,N_8686,N_8772);
or U9432 (N_9432,N_8750,N_8954);
nand U9433 (N_9433,N_8592,N_8596);
or U9434 (N_9434,N_8808,N_8853);
and U9435 (N_9435,N_8844,N_8846);
or U9436 (N_9436,N_8837,N_8891);
nand U9437 (N_9437,N_8604,N_8537);
nor U9438 (N_9438,N_8766,N_8748);
nor U9439 (N_9439,N_8790,N_8564);
and U9440 (N_9440,N_8685,N_8818);
nand U9441 (N_9441,N_8755,N_8909);
or U9442 (N_9442,N_8669,N_8559);
xor U9443 (N_9443,N_8564,N_8839);
or U9444 (N_9444,N_8504,N_8780);
nor U9445 (N_9445,N_8778,N_8532);
and U9446 (N_9446,N_8650,N_8541);
or U9447 (N_9447,N_8710,N_8942);
nor U9448 (N_9448,N_8706,N_8898);
or U9449 (N_9449,N_8979,N_8664);
and U9450 (N_9450,N_8595,N_8922);
and U9451 (N_9451,N_8898,N_8721);
nor U9452 (N_9452,N_8707,N_8953);
or U9453 (N_9453,N_8684,N_8589);
or U9454 (N_9454,N_8779,N_8876);
or U9455 (N_9455,N_8746,N_8751);
nor U9456 (N_9456,N_8808,N_8566);
nand U9457 (N_9457,N_8844,N_8845);
nor U9458 (N_9458,N_8531,N_8746);
and U9459 (N_9459,N_8803,N_8845);
nor U9460 (N_9460,N_8645,N_8525);
or U9461 (N_9461,N_8704,N_8955);
nor U9462 (N_9462,N_8894,N_8778);
and U9463 (N_9463,N_8618,N_8763);
xor U9464 (N_9464,N_8620,N_8686);
nand U9465 (N_9465,N_8626,N_8707);
nand U9466 (N_9466,N_8571,N_8525);
nor U9467 (N_9467,N_8696,N_8604);
or U9468 (N_9468,N_8829,N_8672);
and U9469 (N_9469,N_8768,N_8620);
and U9470 (N_9470,N_8707,N_8598);
or U9471 (N_9471,N_8650,N_8574);
nand U9472 (N_9472,N_8686,N_8829);
or U9473 (N_9473,N_8500,N_8862);
nand U9474 (N_9474,N_8685,N_8529);
nor U9475 (N_9475,N_8552,N_8961);
nor U9476 (N_9476,N_8612,N_8916);
and U9477 (N_9477,N_8704,N_8963);
and U9478 (N_9478,N_8669,N_8592);
nor U9479 (N_9479,N_8586,N_8767);
or U9480 (N_9480,N_8898,N_8602);
nand U9481 (N_9481,N_8725,N_8803);
nor U9482 (N_9482,N_8967,N_8779);
nand U9483 (N_9483,N_8677,N_8624);
xnor U9484 (N_9484,N_8684,N_8753);
nand U9485 (N_9485,N_8530,N_8679);
nand U9486 (N_9486,N_8646,N_8882);
and U9487 (N_9487,N_8597,N_8631);
and U9488 (N_9488,N_8733,N_8576);
nand U9489 (N_9489,N_8915,N_8993);
nor U9490 (N_9490,N_8583,N_8931);
nor U9491 (N_9491,N_8896,N_8955);
nor U9492 (N_9492,N_8958,N_8635);
and U9493 (N_9493,N_8786,N_8697);
and U9494 (N_9494,N_8624,N_8641);
or U9495 (N_9495,N_8567,N_8805);
and U9496 (N_9496,N_8945,N_8628);
or U9497 (N_9497,N_8619,N_8979);
and U9498 (N_9498,N_8691,N_8650);
or U9499 (N_9499,N_8844,N_8654);
nor U9500 (N_9500,N_9473,N_9412);
nand U9501 (N_9501,N_9116,N_9481);
nand U9502 (N_9502,N_9377,N_9199);
nand U9503 (N_9503,N_9156,N_9479);
and U9504 (N_9504,N_9222,N_9451);
nor U9505 (N_9505,N_9234,N_9410);
nor U9506 (N_9506,N_9297,N_9064);
nor U9507 (N_9507,N_9150,N_9106);
nand U9508 (N_9508,N_9491,N_9212);
nor U9509 (N_9509,N_9382,N_9147);
nand U9510 (N_9510,N_9185,N_9157);
nor U9511 (N_9511,N_9276,N_9302);
nand U9512 (N_9512,N_9260,N_9236);
or U9513 (N_9513,N_9361,N_9174);
or U9514 (N_9514,N_9172,N_9215);
and U9515 (N_9515,N_9312,N_9279);
or U9516 (N_9516,N_9207,N_9427);
nor U9517 (N_9517,N_9034,N_9430);
nand U9518 (N_9518,N_9233,N_9120);
or U9519 (N_9519,N_9329,N_9321);
nor U9520 (N_9520,N_9189,N_9243);
or U9521 (N_9521,N_9424,N_9470);
or U9522 (N_9522,N_9217,N_9494);
and U9523 (N_9523,N_9013,N_9265);
nand U9524 (N_9524,N_9250,N_9404);
and U9525 (N_9525,N_9453,N_9067);
nor U9526 (N_9526,N_9002,N_9488);
and U9527 (N_9527,N_9399,N_9240);
and U9528 (N_9528,N_9314,N_9208);
nand U9529 (N_9529,N_9228,N_9118);
nand U9530 (N_9530,N_9449,N_9105);
nand U9531 (N_9531,N_9082,N_9360);
nand U9532 (N_9532,N_9495,N_9176);
or U9533 (N_9533,N_9204,N_9299);
nor U9534 (N_9534,N_9091,N_9017);
xor U9535 (N_9535,N_9325,N_9306);
or U9536 (N_9536,N_9254,N_9261);
and U9537 (N_9537,N_9319,N_9139);
nor U9538 (N_9538,N_9249,N_9422);
nor U9539 (N_9539,N_9386,N_9363);
nand U9540 (N_9540,N_9489,N_9206);
and U9541 (N_9541,N_9478,N_9256);
and U9542 (N_9542,N_9127,N_9187);
nand U9543 (N_9543,N_9037,N_9493);
nor U9544 (N_9544,N_9378,N_9328);
nor U9545 (N_9545,N_9197,N_9179);
and U9546 (N_9546,N_9160,N_9462);
xnor U9547 (N_9547,N_9225,N_9447);
or U9548 (N_9548,N_9027,N_9200);
and U9549 (N_9549,N_9251,N_9330);
nor U9550 (N_9550,N_9242,N_9439);
nor U9551 (N_9551,N_9020,N_9280);
nand U9552 (N_9552,N_9272,N_9030);
and U9553 (N_9553,N_9050,N_9088);
and U9554 (N_9554,N_9262,N_9364);
nor U9555 (N_9555,N_9468,N_9218);
and U9556 (N_9556,N_9009,N_9496);
and U9557 (N_9557,N_9099,N_9372);
nand U9558 (N_9558,N_9390,N_9144);
or U9559 (N_9559,N_9008,N_9061);
xor U9560 (N_9560,N_9438,N_9487);
nor U9561 (N_9561,N_9352,N_9055);
or U9562 (N_9562,N_9431,N_9343);
or U9563 (N_9563,N_9201,N_9095);
nand U9564 (N_9564,N_9333,N_9413);
or U9565 (N_9565,N_9440,N_9283);
and U9566 (N_9566,N_9007,N_9205);
nor U9567 (N_9567,N_9474,N_9112);
nor U9568 (N_9568,N_9367,N_9133);
and U9569 (N_9569,N_9096,N_9429);
and U9570 (N_9570,N_9191,N_9497);
nor U9571 (N_9571,N_9196,N_9420);
and U9572 (N_9572,N_9264,N_9214);
or U9573 (N_9573,N_9137,N_9047);
nand U9574 (N_9574,N_9275,N_9351);
or U9575 (N_9575,N_9461,N_9340);
xor U9576 (N_9576,N_9128,N_9433);
and U9577 (N_9577,N_9428,N_9051);
nor U9578 (N_9578,N_9122,N_9166);
and U9579 (N_9579,N_9288,N_9045);
or U9580 (N_9580,N_9292,N_9031);
and U9581 (N_9581,N_9444,N_9245);
or U9582 (N_9582,N_9028,N_9407);
nand U9583 (N_9583,N_9266,N_9063);
xor U9584 (N_9584,N_9103,N_9130);
nand U9585 (N_9585,N_9350,N_9417);
nand U9586 (N_9586,N_9383,N_9000);
nor U9587 (N_9587,N_9075,N_9403);
nor U9588 (N_9588,N_9300,N_9175);
and U9589 (N_9589,N_9107,N_9224);
nand U9590 (N_9590,N_9258,N_9068);
nand U9591 (N_9591,N_9190,N_9238);
nor U9592 (N_9592,N_9322,N_9317);
xor U9593 (N_9593,N_9001,N_9011);
nor U9594 (N_9594,N_9062,N_9135);
xnor U9595 (N_9595,N_9094,N_9411);
or U9596 (N_9596,N_9347,N_9311);
and U9597 (N_9597,N_9016,N_9467);
or U9598 (N_9598,N_9355,N_9346);
or U9599 (N_9599,N_9257,N_9015);
nand U9600 (N_9600,N_9229,N_9296);
and U9601 (N_9601,N_9371,N_9277);
nand U9602 (N_9602,N_9286,N_9472);
nand U9603 (N_9603,N_9394,N_9337);
nor U9604 (N_9604,N_9216,N_9263);
and U9605 (N_9605,N_9273,N_9052);
and U9606 (N_9606,N_9387,N_9301);
and U9607 (N_9607,N_9396,N_9409);
nor U9608 (N_9608,N_9004,N_9080);
and U9609 (N_9609,N_9448,N_9129);
nor U9610 (N_9610,N_9246,N_9131);
nand U9611 (N_9611,N_9038,N_9101);
and U9612 (N_9612,N_9048,N_9359);
or U9613 (N_9613,N_9119,N_9146);
or U9614 (N_9614,N_9141,N_9056);
and U9615 (N_9615,N_9081,N_9419);
nand U9616 (N_9616,N_9161,N_9142);
and U9617 (N_9617,N_9353,N_9165);
and U9618 (N_9618,N_9108,N_9036);
and U9619 (N_9619,N_9071,N_9078);
and U9620 (N_9620,N_9148,N_9111);
or U9621 (N_9621,N_9385,N_9327);
and U9622 (N_9622,N_9338,N_9211);
nor U9623 (N_9623,N_9090,N_9282);
and U9624 (N_9624,N_9446,N_9092);
xor U9625 (N_9625,N_9425,N_9025);
nand U9626 (N_9626,N_9171,N_9397);
or U9627 (N_9627,N_9093,N_9269);
nand U9628 (N_9628,N_9485,N_9180);
nand U9629 (N_9629,N_9437,N_9332);
and U9630 (N_9630,N_9290,N_9073);
or U9631 (N_9631,N_9193,N_9209);
and U9632 (N_9632,N_9458,N_9226);
nor U9633 (N_9633,N_9158,N_9416);
and U9634 (N_9634,N_9138,N_9252);
or U9635 (N_9635,N_9358,N_9083);
or U9636 (N_9636,N_9298,N_9421);
and U9637 (N_9637,N_9121,N_9305);
or U9638 (N_9638,N_9384,N_9220);
nor U9639 (N_9639,N_9339,N_9356);
nand U9640 (N_9640,N_9046,N_9392);
and U9641 (N_9641,N_9499,N_9151);
nand U9642 (N_9642,N_9309,N_9436);
and U9643 (N_9643,N_9043,N_9369);
nand U9644 (N_9644,N_9365,N_9259);
or U9645 (N_9645,N_9477,N_9223);
nand U9646 (N_9646,N_9124,N_9284);
nand U9647 (N_9647,N_9021,N_9418);
nor U9648 (N_9648,N_9024,N_9460);
nor U9649 (N_9649,N_9401,N_9270);
nor U9650 (N_9650,N_9406,N_9132);
and U9651 (N_9651,N_9498,N_9098);
nand U9652 (N_9652,N_9060,N_9441);
nor U9653 (N_9653,N_9426,N_9086);
and U9654 (N_9654,N_9077,N_9005);
and U9655 (N_9655,N_9239,N_9195);
and U9656 (N_9656,N_9029,N_9408);
and U9657 (N_9657,N_9041,N_9054);
xor U9658 (N_9658,N_9456,N_9089);
nand U9659 (N_9659,N_9115,N_9023);
nor U9660 (N_9660,N_9181,N_9235);
and U9661 (N_9661,N_9295,N_9248);
or U9662 (N_9662,N_9388,N_9465);
and U9663 (N_9663,N_9085,N_9326);
nor U9664 (N_9664,N_9381,N_9318);
or U9665 (N_9665,N_9159,N_9308);
or U9666 (N_9666,N_9471,N_9402);
nand U9667 (N_9667,N_9152,N_9304);
nor U9668 (N_9668,N_9442,N_9227);
or U9669 (N_9669,N_9186,N_9274);
and U9670 (N_9670,N_9084,N_9188);
nand U9671 (N_9671,N_9315,N_9231);
and U9672 (N_9672,N_9357,N_9393);
or U9673 (N_9673,N_9348,N_9010);
nor U9674 (N_9674,N_9219,N_9323);
or U9675 (N_9675,N_9202,N_9482);
nor U9676 (N_9676,N_9278,N_9268);
and U9677 (N_9677,N_9154,N_9042);
or U9678 (N_9678,N_9221,N_9480);
nand U9679 (N_9679,N_9281,N_9345);
and U9680 (N_9680,N_9170,N_9484);
or U9681 (N_9681,N_9452,N_9153);
nor U9682 (N_9682,N_9287,N_9183);
nand U9683 (N_9683,N_9162,N_9102);
nand U9684 (N_9684,N_9395,N_9104);
and U9685 (N_9685,N_9293,N_9069);
nor U9686 (N_9686,N_9044,N_9012);
or U9687 (N_9687,N_9198,N_9033);
or U9688 (N_9688,N_9177,N_9344);
and U9689 (N_9689,N_9289,N_9113);
and U9690 (N_9690,N_9173,N_9167);
or U9691 (N_9691,N_9334,N_9079);
and U9692 (N_9692,N_9109,N_9379);
and U9693 (N_9693,N_9123,N_9059);
or U9694 (N_9694,N_9134,N_9140);
and U9695 (N_9695,N_9163,N_9423);
nand U9696 (N_9696,N_9483,N_9040);
nand U9697 (N_9697,N_9058,N_9398);
nand U9698 (N_9698,N_9271,N_9457);
and U9699 (N_9699,N_9169,N_9366);
or U9700 (N_9700,N_9232,N_9466);
nor U9701 (N_9701,N_9400,N_9267);
and U9702 (N_9702,N_9049,N_9294);
or U9703 (N_9703,N_9476,N_9014);
nor U9704 (N_9704,N_9255,N_9370);
nor U9705 (N_9705,N_9450,N_9168);
or U9706 (N_9706,N_9405,N_9389);
or U9707 (N_9707,N_9316,N_9155);
nand U9708 (N_9708,N_9194,N_9097);
and U9709 (N_9709,N_9039,N_9391);
and U9710 (N_9710,N_9336,N_9022);
nand U9711 (N_9711,N_9443,N_9469);
xnor U9712 (N_9712,N_9241,N_9459);
and U9713 (N_9713,N_9070,N_9237);
or U9714 (N_9714,N_9368,N_9331);
or U9715 (N_9715,N_9026,N_9285);
nand U9716 (N_9716,N_9455,N_9125);
nor U9717 (N_9717,N_9076,N_9303);
nor U9718 (N_9718,N_9486,N_9376);
nand U9719 (N_9719,N_9341,N_9053);
nor U9720 (N_9720,N_9164,N_9464);
nor U9721 (N_9721,N_9244,N_9490);
or U9722 (N_9722,N_9072,N_9324);
nand U9723 (N_9723,N_9230,N_9136);
nand U9724 (N_9724,N_9349,N_9006);
nand U9725 (N_9725,N_9320,N_9414);
xor U9726 (N_9726,N_9032,N_9342);
or U9727 (N_9727,N_9066,N_9475);
nor U9728 (N_9728,N_9380,N_9335);
and U9729 (N_9729,N_9100,N_9210);
nor U9730 (N_9730,N_9184,N_9362);
nand U9731 (N_9731,N_9003,N_9313);
nor U9732 (N_9732,N_9434,N_9114);
nor U9733 (N_9733,N_9463,N_9074);
and U9734 (N_9734,N_9149,N_9035);
nand U9735 (N_9735,N_9454,N_9126);
nand U9736 (N_9736,N_9018,N_9374);
or U9737 (N_9737,N_9145,N_9117);
xnor U9738 (N_9738,N_9373,N_9110);
and U9739 (N_9739,N_9432,N_9307);
nand U9740 (N_9740,N_9203,N_9087);
and U9741 (N_9741,N_9182,N_9057);
nand U9742 (N_9742,N_9065,N_9375);
nand U9743 (N_9743,N_9354,N_9247);
nor U9744 (N_9744,N_9019,N_9213);
nor U9745 (N_9745,N_9310,N_9192);
or U9746 (N_9746,N_9143,N_9492);
and U9747 (N_9747,N_9178,N_9291);
nand U9748 (N_9748,N_9435,N_9253);
nand U9749 (N_9749,N_9415,N_9445);
nand U9750 (N_9750,N_9260,N_9159);
nand U9751 (N_9751,N_9408,N_9296);
or U9752 (N_9752,N_9390,N_9412);
and U9753 (N_9753,N_9345,N_9341);
nand U9754 (N_9754,N_9230,N_9312);
and U9755 (N_9755,N_9453,N_9476);
and U9756 (N_9756,N_9385,N_9393);
and U9757 (N_9757,N_9340,N_9408);
nand U9758 (N_9758,N_9421,N_9063);
nor U9759 (N_9759,N_9481,N_9271);
nand U9760 (N_9760,N_9034,N_9178);
nor U9761 (N_9761,N_9101,N_9350);
and U9762 (N_9762,N_9410,N_9416);
or U9763 (N_9763,N_9208,N_9411);
nand U9764 (N_9764,N_9391,N_9021);
nor U9765 (N_9765,N_9151,N_9188);
nor U9766 (N_9766,N_9410,N_9296);
and U9767 (N_9767,N_9043,N_9093);
or U9768 (N_9768,N_9161,N_9080);
nor U9769 (N_9769,N_9285,N_9457);
nand U9770 (N_9770,N_9371,N_9093);
nand U9771 (N_9771,N_9167,N_9139);
nor U9772 (N_9772,N_9214,N_9015);
nor U9773 (N_9773,N_9171,N_9468);
and U9774 (N_9774,N_9273,N_9353);
or U9775 (N_9775,N_9152,N_9129);
nor U9776 (N_9776,N_9211,N_9057);
nand U9777 (N_9777,N_9267,N_9241);
nor U9778 (N_9778,N_9174,N_9057);
nor U9779 (N_9779,N_9195,N_9378);
nand U9780 (N_9780,N_9287,N_9299);
nor U9781 (N_9781,N_9401,N_9368);
xor U9782 (N_9782,N_9381,N_9205);
and U9783 (N_9783,N_9200,N_9453);
or U9784 (N_9784,N_9341,N_9163);
and U9785 (N_9785,N_9224,N_9361);
nor U9786 (N_9786,N_9276,N_9382);
and U9787 (N_9787,N_9126,N_9039);
or U9788 (N_9788,N_9063,N_9227);
nor U9789 (N_9789,N_9299,N_9279);
nand U9790 (N_9790,N_9323,N_9414);
or U9791 (N_9791,N_9461,N_9334);
and U9792 (N_9792,N_9400,N_9277);
and U9793 (N_9793,N_9100,N_9447);
xor U9794 (N_9794,N_9226,N_9170);
and U9795 (N_9795,N_9459,N_9463);
nand U9796 (N_9796,N_9379,N_9461);
xor U9797 (N_9797,N_9434,N_9263);
or U9798 (N_9798,N_9332,N_9405);
and U9799 (N_9799,N_9114,N_9247);
nand U9800 (N_9800,N_9347,N_9124);
nor U9801 (N_9801,N_9051,N_9150);
nand U9802 (N_9802,N_9029,N_9340);
nand U9803 (N_9803,N_9490,N_9464);
and U9804 (N_9804,N_9453,N_9234);
nand U9805 (N_9805,N_9423,N_9047);
nor U9806 (N_9806,N_9353,N_9115);
nor U9807 (N_9807,N_9227,N_9410);
or U9808 (N_9808,N_9100,N_9293);
nor U9809 (N_9809,N_9111,N_9181);
or U9810 (N_9810,N_9310,N_9138);
nand U9811 (N_9811,N_9271,N_9450);
nor U9812 (N_9812,N_9305,N_9197);
nor U9813 (N_9813,N_9063,N_9468);
nor U9814 (N_9814,N_9486,N_9426);
or U9815 (N_9815,N_9384,N_9150);
nand U9816 (N_9816,N_9328,N_9186);
nand U9817 (N_9817,N_9076,N_9155);
and U9818 (N_9818,N_9391,N_9358);
or U9819 (N_9819,N_9215,N_9368);
and U9820 (N_9820,N_9388,N_9268);
and U9821 (N_9821,N_9039,N_9203);
nor U9822 (N_9822,N_9491,N_9235);
and U9823 (N_9823,N_9023,N_9421);
nand U9824 (N_9824,N_9463,N_9076);
and U9825 (N_9825,N_9408,N_9237);
or U9826 (N_9826,N_9015,N_9494);
or U9827 (N_9827,N_9192,N_9116);
xnor U9828 (N_9828,N_9338,N_9082);
or U9829 (N_9829,N_9176,N_9165);
nor U9830 (N_9830,N_9321,N_9146);
or U9831 (N_9831,N_9383,N_9099);
nand U9832 (N_9832,N_9270,N_9177);
nand U9833 (N_9833,N_9349,N_9452);
nand U9834 (N_9834,N_9254,N_9126);
nand U9835 (N_9835,N_9131,N_9121);
nor U9836 (N_9836,N_9447,N_9326);
nand U9837 (N_9837,N_9173,N_9408);
xor U9838 (N_9838,N_9012,N_9021);
nor U9839 (N_9839,N_9004,N_9126);
nand U9840 (N_9840,N_9218,N_9317);
or U9841 (N_9841,N_9080,N_9307);
xnor U9842 (N_9842,N_9253,N_9405);
nor U9843 (N_9843,N_9134,N_9417);
nand U9844 (N_9844,N_9483,N_9141);
nor U9845 (N_9845,N_9483,N_9263);
and U9846 (N_9846,N_9092,N_9150);
or U9847 (N_9847,N_9469,N_9419);
xor U9848 (N_9848,N_9192,N_9168);
or U9849 (N_9849,N_9359,N_9038);
and U9850 (N_9850,N_9141,N_9276);
and U9851 (N_9851,N_9181,N_9344);
or U9852 (N_9852,N_9232,N_9058);
xnor U9853 (N_9853,N_9145,N_9386);
nor U9854 (N_9854,N_9488,N_9150);
or U9855 (N_9855,N_9339,N_9252);
nand U9856 (N_9856,N_9005,N_9416);
and U9857 (N_9857,N_9244,N_9173);
and U9858 (N_9858,N_9173,N_9479);
nand U9859 (N_9859,N_9371,N_9340);
or U9860 (N_9860,N_9274,N_9381);
xnor U9861 (N_9861,N_9448,N_9289);
and U9862 (N_9862,N_9395,N_9350);
and U9863 (N_9863,N_9260,N_9217);
nor U9864 (N_9864,N_9371,N_9155);
and U9865 (N_9865,N_9063,N_9090);
or U9866 (N_9866,N_9117,N_9018);
xor U9867 (N_9867,N_9159,N_9372);
nand U9868 (N_9868,N_9418,N_9055);
nor U9869 (N_9869,N_9114,N_9337);
and U9870 (N_9870,N_9369,N_9174);
nor U9871 (N_9871,N_9083,N_9413);
nand U9872 (N_9872,N_9464,N_9108);
and U9873 (N_9873,N_9363,N_9359);
nor U9874 (N_9874,N_9456,N_9235);
nor U9875 (N_9875,N_9411,N_9209);
or U9876 (N_9876,N_9172,N_9334);
or U9877 (N_9877,N_9004,N_9082);
or U9878 (N_9878,N_9401,N_9165);
nand U9879 (N_9879,N_9175,N_9072);
or U9880 (N_9880,N_9322,N_9234);
nand U9881 (N_9881,N_9469,N_9083);
nand U9882 (N_9882,N_9260,N_9258);
nor U9883 (N_9883,N_9073,N_9456);
nor U9884 (N_9884,N_9136,N_9354);
or U9885 (N_9885,N_9295,N_9237);
or U9886 (N_9886,N_9058,N_9444);
or U9887 (N_9887,N_9261,N_9250);
nor U9888 (N_9888,N_9059,N_9064);
and U9889 (N_9889,N_9453,N_9358);
nand U9890 (N_9890,N_9199,N_9134);
or U9891 (N_9891,N_9368,N_9015);
and U9892 (N_9892,N_9423,N_9466);
or U9893 (N_9893,N_9046,N_9001);
or U9894 (N_9894,N_9150,N_9457);
and U9895 (N_9895,N_9439,N_9460);
nand U9896 (N_9896,N_9295,N_9227);
or U9897 (N_9897,N_9163,N_9066);
nand U9898 (N_9898,N_9064,N_9191);
nor U9899 (N_9899,N_9191,N_9037);
or U9900 (N_9900,N_9093,N_9059);
nand U9901 (N_9901,N_9352,N_9100);
nand U9902 (N_9902,N_9227,N_9374);
and U9903 (N_9903,N_9375,N_9392);
nor U9904 (N_9904,N_9071,N_9111);
nand U9905 (N_9905,N_9084,N_9130);
nand U9906 (N_9906,N_9457,N_9043);
nor U9907 (N_9907,N_9403,N_9066);
and U9908 (N_9908,N_9083,N_9028);
nor U9909 (N_9909,N_9210,N_9393);
nor U9910 (N_9910,N_9155,N_9420);
nor U9911 (N_9911,N_9134,N_9458);
or U9912 (N_9912,N_9464,N_9167);
nor U9913 (N_9913,N_9005,N_9154);
and U9914 (N_9914,N_9026,N_9152);
nor U9915 (N_9915,N_9429,N_9380);
nand U9916 (N_9916,N_9112,N_9231);
nand U9917 (N_9917,N_9208,N_9234);
and U9918 (N_9918,N_9011,N_9394);
nor U9919 (N_9919,N_9077,N_9325);
nand U9920 (N_9920,N_9149,N_9156);
or U9921 (N_9921,N_9240,N_9472);
nand U9922 (N_9922,N_9308,N_9135);
and U9923 (N_9923,N_9156,N_9469);
and U9924 (N_9924,N_9468,N_9283);
xnor U9925 (N_9925,N_9112,N_9433);
and U9926 (N_9926,N_9271,N_9391);
nand U9927 (N_9927,N_9259,N_9182);
and U9928 (N_9928,N_9266,N_9469);
and U9929 (N_9929,N_9486,N_9389);
and U9930 (N_9930,N_9090,N_9439);
xnor U9931 (N_9931,N_9215,N_9150);
nand U9932 (N_9932,N_9301,N_9494);
nor U9933 (N_9933,N_9036,N_9444);
or U9934 (N_9934,N_9240,N_9436);
xor U9935 (N_9935,N_9156,N_9183);
or U9936 (N_9936,N_9098,N_9270);
nor U9937 (N_9937,N_9040,N_9301);
nor U9938 (N_9938,N_9425,N_9058);
and U9939 (N_9939,N_9059,N_9045);
or U9940 (N_9940,N_9228,N_9158);
and U9941 (N_9941,N_9480,N_9159);
or U9942 (N_9942,N_9170,N_9031);
nand U9943 (N_9943,N_9253,N_9475);
nand U9944 (N_9944,N_9020,N_9354);
nand U9945 (N_9945,N_9492,N_9376);
nor U9946 (N_9946,N_9058,N_9372);
nor U9947 (N_9947,N_9345,N_9086);
and U9948 (N_9948,N_9139,N_9485);
nand U9949 (N_9949,N_9158,N_9018);
nor U9950 (N_9950,N_9415,N_9410);
nor U9951 (N_9951,N_9337,N_9090);
nand U9952 (N_9952,N_9282,N_9302);
nor U9953 (N_9953,N_9383,N_9364);
or U9954 (N_9954,N_9265,N_9140);
nor U9955 (N_9955,N_9165,N_9344);
nand U9956 (N_9956,N_9130,N_9183);
and U9957 (N_9957,N_9240,N_9256);
and U9958 (N_9958,N_9315,N_9277);
or U9959 (N_9959,N_9438,N_9258);
and U9960 (N_9960,N_9257,N_9286);
or U9961 (N_9961,N_9066,N_9011);
nand U9962 (N_9962,N_9064,N_9165);
nor U9963 (N_9963,N_9272,N_9454);
nand U9964 (N_9964,N_9137,N_9395);
nor U9965 (N_9965,N_9052,N_9441);
nor U9966 (N_9966,N_9377,N_9102);
and U9967 (N_9967,N_9084,N_9193);
and U9968 (N_9968,N_9364,N_9293);
nor U9969 (N_9969,N_9112,N_9095);
and U9970 (N_9970,N_9207,N_9266);
nand U9971 (N_9971,N_9021,N_9449);
nor U9972 (N_9972,N_9026,N_9103);
nand U9973 (N_9973,N_9413,N_9012);
nor U9974 (N_9974,N_9095,N_9453);
or U9975 (N_9975,N_9042,N_9258);
nand U9976 (N_9976,N_9011,N_9151);
or U9977 (N_9977,N_9363,N_9042);
or U9978 (N_9978,N_9072,N_9361);
and U9979 (N_9979,N_9008,N_9125);
nand U9980 (N_9980,N_9282,N_9228);
nand U9981 (N_9981,N_9086,N_9420);
nand U9982 (N_9982,N_9085,N_9281);
nand U9983 (N_9983,N_9460,N_9031);
nand U9984 (N_9984,N_9250,N_9011);
nand U9985 (N_9985,N_9141,N_9271);
or U9986 (N_9986,N_9493,N_9238);
nand U9987 (N_9987,N_9082,N_9336);
nand U9988 (N_9988,N_9116,N_9406);
nand U9989 (N_9989,N_9304,N_9292);
nand U9990 (N_9990,N_9054,N_9433);
nor U9991 (N_9991,N_9194,N_9449);
nor U9992 (N_9992,N_9125,N_9442);
and U9993 (N_9993,N_9463,N_9178);
or U9994 (N_9994,N_9241,N_9399);
xor U9995 (N_9995,N_9071,N_9490);
nand U9996 (N_9996,N_9400,N_9084);
or U9997 (N_9997,N_9331,N_9322);
and U9998 (N_9998,N_9417,N_9314);
or U9999 (N_9999,N_9292,N_9075);
nor UO_0 (O_0,N_9824,N_9740);
nand UO_1 (O_1,N_9972,N_9817);
or UO_2 (O_2,N_9903,N_9505);
and UO_3 (O_3,N_9967,N_9850);
nor UO_4 (O_4,N_9602,N_9880);
nor UO_5 (O_5,N_9790,N_9653);
and UO_6 (O_6,N_9864,N_9714);
nand UO_7 (O_7,N_9552,N_9874);
nand UO_8 (O_8,N_9904,N_9726);
nand UO_9 (O_9,N_9551,N_9748);
xor UO_10 (O_10,N_9618,N_9854);
nor UO_11 (O_11,N_9562,N_9773);
and UO_12 (O_12,N_9796,N_9574);
nand UO_13 (O_13,N_9632,N_9544);
and UO_14 (O_14,N_9558,N_9553);
nor UO_15 (O_15,N_9929,N_9987);
and UO_16 (O_16,N_9828,N_9568);
and UO_17 (O_17,N_9986,N_9640);
nand UO_18 (O_18,N_9589,N_9570);
nand UO_19 (O_19,N_9948,N_9901);
and UO_20 (O_20,N_9722,N_9501);
or UO_21 (O_21,N_9756,N_9849);
nor UO_22 (O_22,N_9921,N_9692);
nand UO_23 (O_23,N_9662,N_9718);
nand UO_24 (O_24,N_9684,N_9971);
and UO_25 (O_25,N_9803,N_9584);
nand UO_26 (O_26,N_9676,N_9649);
nand UO_27 (O_27,N_9897,N_9833);
nor UO_28 (O_28,N_9869,N_9706);
and UO_29 (O_29,N_9541,N_9761);
nor UO_30 (O_30,N_9937,N_9703);
nor UO_31 (O_31,N_9882,N_9741);
and UO_32 (O_32,N_9563,N_9855);
or UO_33 (O_33,N_9910,N_9607);
nor UO_34 (O_34,N_9603,N_9680);
nor UO_35 (O_35,N_9786,N_9559);
nor UO_36 (O_36,N_9592,N_9908);
nor UO_37 (O_37,N_9531,N_9823);
nor UO_38 (O_38,N_9645,N_9567);
nor UO_39 (O_39,N_9715,N_9515);
nand UO_40 (O_40,N_9853,N_9927);
and UO_41 (O_41,N_9754,N_9815);
or UO_42 (O_42,N_9651,N_9524);
nor UO_43 (O_43,N_9711,N_9700);
nand UO_44 (O_44,N_9776,N_9890);
nor UO_45 (O_45,N_9822,N_9801);
nor UO_46 (O_46,N_9642,N_9737);
and UO_47 (O_47,N_9917,N_9941);
nand UO_48 (O_48,N_9628,N_9959);
or UO_49 (O_49,N_9652,N_9968);
and UO_50 (O_50,N_9919,N_9637);
xor UO_51 (O_51,N_9630,N_9569);
nand UO_52 (O_52,N_9634,N_9956);
or UO_53 (O_53,N_9591,N_9852);
or UO_54 (O_54,N_9902,N_9696);
and UO_55 (O_55,N_9557,N_9939);
nand UO_56 (O_56,N_9631,N_9673);
or UO_57 (O_57,N_9646,N_9510);
nor UO_58 (O_58,N_9808,N_9728);
or UO_59 (O_59,N_9845,N_9774);
nand UO_60 (O_60,N_9780,N_9738);
nor UO_61 (O_61,N_9935,N_9861);
nor UO_62 (O_62,N_9763,N_9647);
or UO_63 (O_63,N_9520,N_9605);
nor UO_64 (O_64,N_9606,N_9920);
nor UO_65 (O_65,N_9566,N_9907);
or UO_66 (O_66,N_9709,N_9678);
or UO_67 (O_67,N_9529,N_9835);
and UO_68 (O_68,N_9608,N_9648);
or UO_69 (O_69,N_9526,N_9571);
and UO_70 (O_70,N_9745,N_9858);
nand UO_71 (O_71,N_9821,N_9621);
nor UO_72 (O_72,N_9970,N_9781);
nand UO_73 (O_73,N_9791,N_9827);
nor UO_74 (O_74,N_9635,N_9554);
nand UO_75 (O_75,N_9543,N_9800);
or UO_76 (O_76,N_9712,N_9985);
and UO_77 (O_77,N_9946,N_9590);
nand UO_78 (O_78,N_9831,N_9926);
or UO_79 (O_79,N_9685,N_9725);
nor UO_80 (O_80,N_9577,N_9922);
nor UO_81 (O_81,N_9534,N_9832);
nor UO_82 (O_82,N_9744,N_9597);
or UO_83 (O_83,N_9930,N_9964);
and UO_84 (O_84,N_9810,N_9547);
and UO_85 (O_85,N_9913,N_9996);
nor UO_86 (O_86,N_9537,N_9578);
xnor UO_87 (O_87,N_9693,N_9743);
nand UO_88 (O_88,N_9719,N_9573);
and UO_89 (O_89,N_9953,N_9610);
and UO_90 (O_90,N_9699,N_9976);
and UO_91 (O_91,N_9538,N_9876);
nand UO_92 (O_92,N_9733,N_9825);
and UO_93 (O_93,N_9797,N_9936);
or UO_94 (O_94,N_9881,N_9670);
nor UO_95 (O_95,N_9951,N_9585);
or UO_96 (O_96,N_9812,N_9807);
or UO_97 (O_97,N_9883,N_9766);
nor UO_98 (O_98,N_9517,N_9896);
nand UO_99 (O_99,N_9504,N_9898);
nor UO_100 (O_100,N_9809,N_9717);
nor UO_101 (O_101,N_9995,N_9656);
or UO_102 (O_102,N_9928,N_9788);
and UO_103 (O_103,N_9530,N_9851);
nand UO_104 (O_104,N_9730,N_9514);
nor UO_105 (O_105,N_9620,N_9724);
nand UO_106 (O_106,N_9793,N_9508);
xnor UO_107 (O_107,N_9870,N_9871);
and UO_108 (O_108,N_9842,N_9594);
and UO_109 (O_109,N_9772,N_9931);
and UO_110 (O_110,N_9736,N_9636);
nand UO_111 (O_111,N_9616,N_9522);
nand UO_112 (O_112,N_9990,N_9701);
or UO_113 (O_113,N_9997,N_9688);
nand UO_114 (O_114,N_9866,N_9657);
nor UO_115 (O_115,N_9583,N_9775);
nor UO_116 (O_116,N_9671,N_9527);
nor UO_117 (O_117,N_9778,N_9731);
nor UO_118 (O_118,N_9844,N_9818);
or UO_119 (O_119,N_9945,N_9599);
nand UO_120 (O_120,N_9969,N_9598);
nor UO_121 (O_121,N_9965,N_9681);
nor UO_122 (O_122,N_9752,N_9750);
nand UO_123 (O_123,N_9804,N_9973);
nand UO_124 (O_124,N_9802,N_9723);
xnor UO_125 (O_125,N_9507,N_9708);
nor UO_126 (O_126,N_9887,N_9899);
nand UO_127 (O_127,N_9934,N_9694);
nand UO_128 (O_128,N_9713,N_9716);
or UO_129 (O_129,N_9665,N_9873);
nand UO_130 (O_130,N_9792,N_9848);
nor UO_131 (O_131,N_9669,N_9655);
nor UO_132 (O_132,N_9674,N_9998);
nor UO_133 (O_133,N_9843,N_9769);
or UO_134 (O_134,N_9698,N_9555);
and UO_135 (O_135,N_9867,N_9641);
and UO_136 (O_136,N_9727,N_9878);
and UO_137 (O_137,N_9675,N_9575);
nor UO_138 (O_138,N_9548,N_9952);
and UO_139 (O_139,N_9622,N_9747);
or UO_140 (O_140,N_9545,N_9872);
and UO_141 (O_141,N_9550,N_9734);
or UO_142 (O_142,N_9638,N_9729);
or UO_143 (O_143,N_9885,N_9512);
nand UO_144 (O_144,N_9954,N_9888);
and UO_145 (O_145,N_9863,N_9933);
and UO_146 (O_146,N_9923,N_9509);
and UO_147 (O_147,N_9771,N_9753);
or UO_148 (O_148,N_9629,N_9539);
nor UO_149 (O_149,N_9875,N_9837);
or UO_150 (O_150,N_9609,N_9667);
and UO_151 (O_151,N_9593,N_9565);
nor UO_152 (O_152,N_9588,N_9877);
or UO_153 (O_153,N_9991,N_9915);
and UO_154 (O_154,N_9798,N_9758);
nand UO_155 (O_155,N_9892,N_9770);
and UO_156 (O_156,N_9695,N_9556);
xor UO_157 (O_157,N_9579,N_9633);
nand UO_158 (O_158,N_9511,N_9962);
nor UO_159 (O_159,N_9742,N_9705);
or UO_160 (O_160,N_9978,N_9813);
and UO_161 (O_161,N_9572,N_9942);
nor UO_162 (O_162,N_9940,N_9513);
nor UO_163 (O_163,N_9966,N_9615);
nand UO_164 (O_164,N_9604,N_9523);
nor UO_165 (O_165,N_9977,N_9768);
nor UO_166 (O_166,N_9784,N_9687);
and UO_167 (O_167,N_9516,N_9884);
nand UO_168 (O_168,N_9980,N_9519);
xnor UO_169 (O_169,N_9658,N_9777);
nand UO_170 (O_170,N_9982,N_9889);
and UO_171 (O_171,N_9617,N_9785);
nand UO_172 (O_172,N_9668,N_9895);
and UO_173 (O_173,N_9746,N_9826);
and UO_174 (O_174,N_9625,N_9814);
nor UO_175 (O_175,N_9536,N_9533);
and UO_176 (O_176,N_9999,N_9672);
nand UO_177 (O_177,N_9664,N_9949);
nor UO_178 (O_178,N_9686,N_9830);
or UO_179 (O_179,N_9805,N_9542);
or UO_180 (O_180,N_9783,N_9834);
nor UO_181 (O_181,N_9794,N_9900);
nor UO_182 (O_182,N_9663,N_9535);
nand UO_183 (O_183,N_9587,N_9626);
xor UO_184 (O_184,N_9916,N_9912);
nand UO_185 (O_185,N_9650,N_9525);
nand UO_186 (O_186,N_9816,N_9984);
xnor UO_187 (O_187,N_9540,N_9576);
nor UO_188 (O_188,N_9613,N_9528);
nand UO_189 (O_189,N_9677,N_9865);
and UO_190 (O_190,N_9857,N_9732);
or UO_191 (O_191,N_9707,N_9721);
or UO_192 (O_192,N_9847,N_9679);
nand UO_193 (O_193,N_9979,N_9759);
nand UO_194 (O_194,N_9811,N_9581);
nand UO_195 (O_195,N_9683,N_9596);
nor UO_196 (O_196,N_9955,N_9600);
and UO_197 (O_197,N_9654,N_9503);
nand UO_198 (O_198,N_9947,N_9661);
nand UO_199 (O_199,N_9720,N_9893);
and UO_200 (O_200,N_9846,N_9521);
nand UO_201 (O_201,N_9739,N_9561);
nor UO_202 (O_202,N_9960,N_9838);
nor UO_203 (O_203,N_9697,N_9765);
nand UO_204 (O_204,N_9820,N_9840);
nand UO_205 (O_205,N_9690,N_9983);
nor UO_206 (O_206,N_9918,N_9619);
or UO_207 (O_207,N_9623,N_9611);
nor UO_208 (O_208,N_9764,N_9779);
and UO_209 (O_209,N_9806,N_9682);
nand UO_210 (O_210,N_9894,N_9659);
nand UO_211 (O_211,N_9924,N_9767);
and UO_212 (O_212,N_9839,N_9932);
or UO_213 (O_213,N_9549,N_9860);
nor UO_214 (O_214,N_9981,N_9958);
nor UO_215 (O_215,N_9612,N_9950);
and UO_216 (O_216,N_9974,N_9710);
nand UO_217 (O_217,N_9582,N_9819);
nor UO_218 (O_218,N_9944,N_9757);
nor UO_219 (O_219,N_9789,N_9595);
or UO_220 (O_220,N_9957,N_9782);
xor UO_221 (O_221,N_9643,N_9564);
xnor UO_222 (O_222,N_9886,N_9644);
nor UO_223 (O_223,N_9580,N_9601);
and UO_224 (O_224,N_9532,N_9502);
or UO_225 (O_225,N_9660,N_9500);
and UO_226 (O_226,N_9891,N_9994);
nor UO_227 (O_227,N_9879,N_9751);
or UO_228 (O_228,N_9735,N_9989);
nor UO_229 (O_229,N_9586,N_9506);
nor UO_230 (O_230,N_9914,N_9627);
or UO_231 (O_231,N_9988,N_9829);
nor UO_232 (O_232,N_9992,N_9560);
and UO_233 (O_233,N_9911,N_9749);
nor UO_234 (O_234,N_9925,N_9856);
or UO_235 (O_235,N_9799,N_9760);
and UO_236 (O_236,N_9762,N_9963);
nor UO_237 (O_237,N_9787,N_9906);
nand UO_238 (O_238,N_9943,N_9614);
and UO_239 (O_239,N_9639,N_9624);
or UO_240 (O_240,N_9859,N_9961);
or UO_241 (O_241,N_9905,N_9689);
nor UO_242 (O_242,N_9862,N_9795);
nor UO_243 (O_243,N_9938,N_9704);
or UO_244 (O_244,N_9868,N_9755);
or UO_245 (O_245,N_9702,N_9993);
or UO_246 (O_246,N_9975,N_9691);
nor UO_247 (O_247,N_9518,N_9909);
or UO_248 (O_248,N_9546,N_9841);
nor UO_249 (O_249,N_9836,N_9666);
nor UO_250 (O_250,N_9820,N_9898);
nor UO_251 (O_251,N_9856,N_9606);
nand UO_252 (O_252,N_9730,N_9962);
nor UO_253 (O_253,N_9620,N_9625);
nor UO_254 (O_254,N_9995,N_9820);
and UO_255 (O_255,N_9949,N_9607);
nor UO_256 (O_256,N_9850,N_9733);
and UO_257 (O_257,N_9948,N_9778);
nand UO_258 (O_258,N_9500,N_9664);
or UO_259 (O_259,N_9812,N_9553);
and UO_260 (O_260,N_9845,N_9926);
nor UO_261 (O_261,N_9589,N_9698);
and UO_262 (O_262,N_9726,N_9809);
and UO_263 (O_263,N_9926,N_9854);
nand UO_264 (O_264,N_9672,N_9862);
or UO_265 (O_265,N_9596,N_9648);
nor UO_266 (O_266,N_9610,N_9800);
or UO_267 (O_267,N_9778,N_9864);
and UO_268 (O_268,N_9578,N_9761);
nand UO_269 (O_269,N_9624,N_9758);
and UO_270 (O_270,N_9608,N_9986);
nand UO_271 (O_271,N_9511,N_9549);
and UO_272 (O_272,N_9713,N_9608);
nor UO_273 (O_273,N_9600,N_9756);
xnor UO_274 (O_274,N_9783,N_9529);
and UO_275 (O_275,N_9862,N_9542);
nor UO_276 (O_276,N_9738,N_9666);
nor UO_277 (O_277,N_9755,N_9621);
nor UO_278 (O_278,N_9775,N_9711);
nand UO_279 (O_279,N_9903,N_9738);
nand UO_280 (O_280,N_9878,N_9814);
nand UO_281 (O_281,N_9689,N_9568);
or UO_282 (O_282,N_9984,N_9973);
and UO_283 (O_283,N_9834,N_9612);
and UO_284 (O_284,N_9816,N_9843);
nor UO_285 (O_285,N_9908,N_9598);
nand UO_286 (O_286,N_9582,N_9959);
or UO_287 (O_287,N_9545,N_9976);
nand UO_288 (O_288,N_9570,N_9703);
nor UO_289 (O_289,N_9704,N_9906);
or UO_290 (O_290,N_9564,N_9827);
nand UO_291 (O_291,N_9873,N_9671);
and UO_292 (O_292,N_9992,N_9960);
or UO_293 (O_293,N_9549,N_9855);
nand UO_294 (O_294,N_9823,N_9884);
and UO_295 (O_295,N_9784,N_9755);
xor UO_296 (O_296,N_9658,N_9726);
nand UO_297 (O_297,N_9706,N_9723);
or UO_298 (O_298,N_9872,N_9726);
and UO_299 (O_299,N_9601,N_9581);
and UO_300 (O_300,N_9643,N_9642);
nor UO_301 (O_301,N_9897,N_9623);
and UO_302 (O_302,N_9965,N_9793);
and UO_303 (O_303,N_9711,N_9967);
and UO_304 (O_304,N_9564,N_9989);
nor UO_305 (O_305,N_9819,N_9856);
and UO_306 (O_306,N_9538,N_9577);
nor UO_307 (O_307,N_9743,N_9510);
or UO_308 (O_308,N_9780,N_9628);
nor UO_309 (O_309,N_9667,N_9913);
nand UO_310 (O_310,N_9883,N_9971);
and UO_311 (O_311,N_9697,N_9906);
nor UO_312 (O_312,N_9919,N_9871);
and UO_313 (O_313,N_9746,N_9876);
nand UO_314 (O_314,N_9786,N_9803);
nand UO_315 (O_315,N_9877,N_9914);
and UO_316 (O_316,N_9707,N_9821);
nand UO_317 (O_317,N_9689,N_9703);
nand UO_318 (O_318,N_9684,N_9990);
nand UO_319 (O_319,N_9890,N_9901);
nor UO_320 (O_320,N_9770,N_9525);
or UO_321 (O_321,N_9744,N_9790);
xnor UO_322 (O_322,N_9868,N_9896);
nand UO_323 (O_323,N_9602,N_9956);
xnor UO_324 (O_324,N_9594,N_9538);
or UO_325 (O_325,N_9507,N_9797);
and UO_326 (O_326,N_9619,N_9718);
nand UO_327 (O_327,N_9621,N_9690);
and UO_328 (O_328,N_9709,N_9746);
nand UO_329 (O_329,N_9737,N_9994);
or UO_330 (O_330,N_9760,N_9565);
nor UO_331 (O_331,N_9717,N_9637);
nand UO_332 (O_332,N_9533,N_9672);
or UO_333 (O_333,N_9537,N_9597);
nand UO_334 (O_334,N_9985,N_9683);
nor UO_335 (O_335,N_9869,N_9856);
nand UO_336 (O_336,N_9854,N_9998);
nand UO_337 (O_337,N_9510,N_9938);
and UO_338 (O_338,N_9641,N_9645);
or UO_339 (O_339,N_9657,N_9700);
or UO_340 (O_340,N_9785,N_9769);
or UO_341 (O_341,N_9574,N_9958);
nor UO_342 (O_342,N_9976,N_9990);
and UO_343 (O_343,N_9790,N_9566);
nand UO_344 (O_344,N_9896,N_9871);
or UO_345 (O_345,N_9772,N_9925);
or UO_346 (O_346,N_9607,N_9727);
nand UO_347 (O_347,N_9662,N_9609);
nor UO_348 (O_348,N_9599,N_9760);
and UO_349 (O_349,N_9770,N_9881);
nor UO_350 (O_350,N_9939,N_9573);
or UO_351 (O_351,N_9594,N_9781);
nor UO_352 (O_352,N_9872,N_9621);
nor UO_353 (O_353,N_9998,N_9556);
and UO_354 (O_354,N_9729,N_9846);
and UO_355 (O_355,N_9939,N_9850);
nor UO_356 (O_356,N_9564,N_9612);
or UO_357 (O_357,N_9651,N_9548);
and UO_358 (O_358,N_9546,N_9790);
xnor UO_359 (O_359,N_9839,N_9568);
nand UO_360 (O_360,N_9544,N_9652);
and UO_361 (O_361,N_9662,N_9936);
nor UO_362 (O_362,N_9808,N_9549);
and UO_363 (O_363,N_9973,N_9640);
nor UO_364 (O_364,N_9813,N_9727);
or UO_365 (O_365,N_9669,N_9810);
or UO_366 (O_366,N_9845,N_9874);
nand UO_367 (O_367,N_9696,N_9562);
nand UO_368 (O_368,N_9706,N_9762);
nand UO_369 (O_369,N_9772,N_9530);
or UO_370 (O_370,N_9809,N_9815);
nand UO_371 (O_371,N_9913,N_9972);
xor UO_372 (O_372,N_9794,N_9538);
nor UO_373 (O_373,N_9828,N_9590);
and UO_374 (O_374,N_9738,N_9700);
nor UO_375 (O_375,N_9707,N_9708);
nor UO_376 (O_376,N_9990,N_9857);
and UO_377 (O_377,N_9624,N_9842);
nand UO_378 (O_378,N_9702,N_9600);
nand UO_379 (O_379,N_9870,N_9925);
nor UO_380 (O_380,N_9634,N_9536);
nor UO_381 (O_381,N_9814,N_9549);
xnor UO_382 (O_382,N_9991,N_9629);
and UO_383 (O_383,N_9665,N_9995);
or UO_384 (O_384,N_9961,N_9995);
and UO_385 (O_385,N_9974,N_9752);
nor UO_386 (O_386,N_9653,N_9526);
or UO_387 (O_387,N_9983,N_9765);
and UO_388 (O_388,N_9502,N_9970);
or UO_389 (O_389,N_9778,N_9875);
nor UO_390 (O_390,N_9945,N_9503);
nor UO_391 (O_391,N_9511,N_9592);
nor UO_392 (O_392,N_9862,N_9847);
nand UO_393 (O_393,N_9822,N_9805);
nand UO_394 (O_394,N_9618,N_9533);
and UO_395 (O_395,N_9578,N_9534);
nor UO_396 (O_396,N_9644,N_9975);
or UO_397 (O_397,N_9911,N_9865);
or UO_398 (O_398,N_9590,N_9772);
and UO_399 (O_399,N_9616,N_9750);
xor UO_400 (O_400,N_9823,N_9755);
and UO_401 (O_401,N_9687,N_9838);
and UO_402 (O_402,N_9901,N_9979);
or UO_403 (O_403,N_9979,N_9795);
and UO_404 (O_404,N_9558,N_9685);
or UO_405 (O_405,N_9974,N_9992);
nand UO_406 (O_406,N_9857,N_9825);
or UO_407 (O_407,N_9891,N_9988);
nand UO_408 (O_408,N_9905,N_9789);
nor UO_409 (O_409,N_9550,N_9972);
or UO_410 (O_410,N_9592,N_9832);
or UO_411 (O_411,N_9520,N_9823);
xor UO_412 (O_412,N_9863,N_9575);
or UO_413 (O_413,N_9813,N_9514);
nand UO_414 (O_414,N_9779,N_9916);
nor UO_415 (O_415,N_9705,N_9525);
or UO_416 (O_416,N_9827,N_9883);
or UO_417 (O_417,N_9608,N_9889);
nor UO_418 (O_418,N_9700,N_9622);
and UO_419 (O_419,N_9590,N_9666);
nor UO_420 (O_420,N_9947,N_9557);
or UO_421 (O_421,N_9956,N_9726);
or UO_422 (O_422,N_9519,N_9543);
nand UO_423 (O_423,N_9872,N_9666);
nand UO_424 (O_424,N_9851,N_9988);
or UO_425 (O_425,N_9873,N_9761);
or UO_426 (O_426,N_9580,N_9642);
nand UO_427 (O_427,N_9940,N_9787);
nand UO_428 (O_428,N_9569,N_9720);
and UO_429 (O_429,N_9600,N_9543);
nor UO_430 (O_430,N_9668,N_9851);
nor UO_431 (O_431,N_9868,N_9922);
or UO_432 (O_432,N_9684,N_9657);
nand UO_433 (O_433,N_9961,N_9950);
nand UO_434 (O_434,N_9811,N_9907);
and UO_435 (O_435,N_9928,N_9643);
xor UO_436 (O_436,N_9590,N_9799);
and UO_437 (O_437,N_9730,N_9961);
or UO_438 (O_438,N_9767,N_9709);
xor UO_439 (O_439,N_9985,N_9656);
or UO_440 (O_440,N_9724,N_9662);
nor UO_441 (O_441,N_9801,N_9611);
and UO_442 (O_442,N_9589,N_9933);
xnor UO_443 (O_443,N_9880,N_9750);
or UO_444 (O_444,N_9508,N_9573);
and UO_445 (O_445,N_9663,N_9769);
nor UO_446 (O_446,N_9569,N_9825);
xnor UO_447 (O_447,N_9978,N_9616);
and UO_448 (O_448,N_9590,N_9855);
and UO_449 (O_449,N_9549,N_9888);
or UO_450 (O_450,N_9883,N_9525);
or UO_451 (O_451,N_9577,N_9976);
and UO_452 (O_452,N_9639,N_9965);
or UO_453 (O_453,N_9740,N_9554);
nand UO_454 (O_454,N_9660,N_9713);
nor UO_455 (O_455,N_9895,N_9743);
nand UO_456 (O_456,N_9765,N_9865);
nor UO_457 (O_457,N_9586,N_9750);
nand UO_458 (O_458,N_9668,N_9894);
or UO_459 (O_459,N_9540,N_9759);
and UO_460 (O_460,N_9618,N_9695);
or UO_461 (O_461,N_9958,N_9926);
or UO_462 (O_462,N_9690,N_9839);
or UO_463 (O_463,N_9672,N_9744);
nand UO_464 (O_464,N_9894,N_9553);
nand UO_465 (O_465,N_9505,N_9586);
nor UO_466 (O_466,N_9522,N_9737);
nand UO_467 (O_467,N_9607,N_9534);
nor UO_468 (O_468,N_9886,N_9894);
or UO_469 (O_469,N_9747,N_9942);
nor UO_470 (O_470,N_9728,N_9811);
or UO_471 (O_471,N_9797,N_9680);
nor UO_472 (O_472,N_9922,N_9712);
nor UO_473 (O_473,N_9758,N_9639);
nor UO_474 (O_474,N_9831,N_9746);
or UO_475 (O_475,N_9960,N_9685);
or UO_476 (O_476,N_9908,N_9775);
nor UO_477 (O_477,N_9581,N_9711);
nand UO_478 (O_478,N_9641,N_9913);
nand UO_479 (O_479,N_9993,N_9810);
nand UO_480 (O_480,N_9696,N_9525);
nand UO_481 (O_481,N_9630,N_9962);
nor UO_482 (O_482,N_9607,N_9749);
nand UO_483 (O_483,N_9898,N_9641);
or UO_484 (O_484,N_9772,N_9722);
and UO_485 (O_485,N_9554,N_9922);
or UO_486 (O_486,N_9776,N_9796);
xor UO_487 (O_487,N_9542,N_9902);
and UO_488 (O_488,N_9890,N_9822);
nand UO_489 (O_489,N_9729,N_9581);
nor UO_490 (O_490,N_9583,N_9862);
nand UO_491 (O_491,N_9818,N_9917);
nor UO_492 (O_492,N_9965,N_9910);
and UO_493 (O_493,N_9877,N_9748);
or UO_494 (O_494,N_9556,N_9883);
and UO_495 (O_495,N_9805,N_9889);
nand UO_496 (O_496,N_9899,N_9701);
nor UO_497 (O_497,N_9588,N_9952);
and UO_498 (O_498,N_9551,N_9926);
and UO_499 (O_499,N_9835,N_9832);
xor UO_500 (O_500,N_9771,N_9741);
nor UO_501 (O_501,N_9876,N_9815);
nand UO_502 (O_502,N_9652,N_9846);
nor UO_503 (O_503,N_9519,N_9649);
nor UO_504 (O_504,N_9778,N_9754);
or UO_505 (O_505,N_9982,N_9824);
nor UO_506 (O_506,N_9757,N_9749);
or UO_507 (O_507,N_9584,N_9683);
nor UO_508 (O_508,N_9986,N_9647);
and UO_509 (O_509,N_9940,N_9832);
nor UO_510 (O_510,N_9707,N_9685);
nor UO_511 (O_511,N_9825,N_9814);
or UO_512 (O_512,N_9766,N_9620);
and UO_513 (O_513,N_9889,N_9679);
nor UO_514 (O_514,N_9658,N_9973);
and UO_515 (O_515,N_9944,N_9646);
xor UO_516 (O_516,N_9532,N_9672);
or UO_517 (O_517,N_9670,N_9548);
nor UO_518 (O_518,N_9742,N_9568);
nand UO_519 (O_519,N_9704,N_9942);
or UO_520 (O_520,N_9545,N_9670);
nand UO_521 (O_521,N_9961,N_9933);
nand UO_522 (O_522,N_9540,N_9524);
nor UO_523 (O_523,N_9962,N_9603);
or UO_524 (O_524,N_9795,N_9928);
and UO_525 (O_525,N_9600,N_9781);
and UO_526 (O_526,N_9510,N_9921);
nor UO_527 (O_527,N_9663,N_9725);
and UO_528 (O_528,N_9830,N_9603);
or UO_529 (O_529,N_9823,N_9945);
and UO_530 (O_530,N_9536,N_9689);
or UO_531 (O_531,N_9960,N_9568);
and UO_532 (O_532,N_9981,N_9942);
and UO_533 (O_533,N_9740,N_9530);
or UO_534 (O_534,N_9501,N_9645);
nor UO_535 (O_535,N_9717,N_9519);
xor UO_536 (O_536,N_9558,N_9942);
or UO_537 (O_537,N_9571,N_9831);
or UO_538 (O_538,N_9568,N_9942);
nor UO_539 (O_539,N_9873,N_9603);
or UO_540 (O_540,N_9981,N_9615);
nor UO_541 (O_541,N_9504,N_9720);
nand UO_542 (O_542,N_9619,N_9507);
or UO_543 (O_543,N_9655,N_9762);
or UO_544 (O_544,N_9819,N_9767);
nand UO_545 (O_545,N_9724,N_9739);
or UO_546 (O_546,N_9767,N_9834);
nand UO_547 (O_547,N_9638,N_9877);
or UO_548 (O_548,N_9516,N_9504);
nand UO_549 (O_549,N_9723,N_9794);
and UO_550 (O_550,N_9682,N_9957);
nor UO_551 (O_551,N_9902,N_9517);
nand UO_552 (O_552,N_9812,N_9873);
nor UO_553 (O_553,N_9735,N_9894);
nand UO_554 (O_554,N_9633,N_9529);
nor UO_555 (O_555,N_9899,N_9845);
nand UO_556 (O_556,N_9877,N_9671);
xor UO_557 (O_557,N_9855,N_9655);
and UO_558 (O_558,N_9977,N_9883);
and UO_559 (O_559,N_9906,N_9882);
nor UO_560 (O_560,N_9891,N_9508);
nand UO_561 (O_561,N_9952,N_9783);
or UO_562 (O_562,N_9606,N_9931);
and UO_563 (O_563,N_9909,N_9979);
nand UO_564 (O_564,N_9700,N_9518);
nor UO_565 (O_565,N_9665,N_9834);
nor UO_566 (O_566,N_9739,N_9604);
and UO_567 (O_567,N_9794,N_9656);
nor UO_568 (O_568,N_9642,N_9817);
nor UO_569 (O_569,N_9811,N_9839);
nor UO_570 (O_570,N_9554,N_9994);
or UO_571 (O_571,N_9726,N_9659);
nand UO_572 (O_572,N_9782,N_9838);
nand UO_573 (O_573,N_9763,N_9660);
nor UO_574 (O_574,N_9901,N_9581);
and UO_575 (O_575,N_9530,N_9617);
nand UO_576 (O_576,N_9545,N_9643);
nor UO_577 (O_577,N_9903,N_9687);
nor UO_578 (O_578,N_9629,N_9548);
and UO_579 (O_579,N_9873,N_9736);
and UO_580 (O_580,N_9976,N_9878);
nand UO_581 (O_581,N_9756,N_9763);
nand UO_582 (O_582,N_9972,N_9885);
and UO_583 (O_583,N_9678,N_9928);
nor UO_584 (O_584,N_9567,N_9938);
and UO_585 (O_585,N_9729,N_9750);
nand UO_586 (O_586,N_9513,N_9871);
and UO_587 (O_587,N_9967,N_9761);
nor UO_588 (O_588,N_9764,N_9775);
nand UO_589 (O_589,N_9525,N_9549);
nor UO_590 (O_590,N_9666,N_9694);
or UO_591 (O_591,N_9955,N_9977);
nand UO_592 (O_592,N_9869,N_9827);
and UO_593 (O_593,N_9973,N_9766);
or UO_594 (O_594,N_9826,N_9674);
nand UO_595 (O_595,N_9964,N_9986);
and UO_596 (O_596,N_9528,N_9622);
nand UO_597 (O_597,N_9952,N_9876);
nand UO_598 (O_598,N_9608,N_9693);
or UO_599 (O_599,N_9532,N_9978);
nand UO_600 (O_600,N_9986,N_9967);
nand UO_601 (O_601,N_9818,N_9565);
nor UO_602 (O_602,N_9674,N_9916);
or UO_603 (O_603,N_9826,N_9662);
and UO_604 (O_604,N_9737,N_9751);
nor UO_605 (O_605,N_9810,N_9843);
nor UO_606 (O_606,N_9539,N_9509);
nor UO_607 (O_607,N_9629,N_9917);
and UO_608 (O_608,N_9629,N_9705);
or UO_609 (O_609,N_9662,N_9925);
nand UO_610 (O_610,N_9532,N_9610);
nand UO_611 (O_611,N_9879,N_9706);
nor UO_612 (O_612,N_9961,N_9973);
or UO_613 (O_613,N_9850,N_9772);
nor UO_614 (O_614,N_9703,N_9634);
nor UO_615 (O_615,N_9881,N_9987);
nand UO_616 (O_616,N_9543,N_9569);
nand UO_617 (O_617,N_9779,N_9920);
nand UO_618 (O_618,N_9743,N_9607);
and UO_619 (O_619,N_9982,N_9501);
nor UO_620 (O_620,N_9998,N_9947);
or UO_621 (O_621,N_9621,N_9954);
nand UO_622 (O_622,N_9924,N_9997);
nor UO_623 (O_623,N_9808,N_9897);
nand UO_624 (O_624,N_9619,N_9844);
nand UO_625 (O_625,N_9663,N_9592);
nor UO_626 (O_626,N_9832,N_9885);
and UO_627 (O_627,N_9605,N_9981);
or UO_628 (O_628,N_9882,N_9898);
nand UO_629 (O_629,N_9879,N_9538);
or UO_630 (O_630,N_9789,N_9801);
xnor UO_631 (O_631,N_9626,N_9692);
nand UO_632 (O_632,N_9774,N_9813);
or UO_633 (O_633,N_9798,N_9585);
and UO_634 (O_634,N_9865,N_9531);
nand UO_635 (O_635,N_9914,N_9917);
nand UO_636 (O_636,N_9892,N_9984);
nor UO_637 (O_637,N_9524,N_9869);
and UO_638 (O_638,N_9870,N_9717);
nand UO_639 (O_639,N_9527,N_9584);
nand UO_640 (O_640,N_9809,N_9509);
nor UO_641 (O_641,N_9706,N_9832);
or UO_642 (O_642,N_9859,N_9836);
or UO_643 (O_643,N_9942,N_9837);
and UO_644 (O_644,N_9952,N_9603);
and UO_645 (O_645,N_9869,N_9743);
nand UO_646 (O_646,N_9883,N_9554);
or UO_647 (O_647,N_9689,N_9692);
or UO_648 (O_648,N_9559,N_9896);
xnor UO_649 (O_649,N_9851,N_9524);
nand UO_650 (O_650,N_9921,N_9544);
and UO_651 (O_651,N_9521,N_9565);
nor UO_652 (O_652,N_9966,N_9974);
or UO_653 (O_653,N_9640,N_9902);
nor UO_654 (O_654,N_9850,N_9726);
nand UO_655 (O_655,N_9978,N_9565);
and UO_656 (O_656,N_9655,N_9698);
nor UO_657 (O_657,N_9748,N_9955);
or UO_658 (O_658,N_9982,N_9512);
and UO_659 (O_659,N_9538,N_9635);
nand UO_660 (O_660,N_9969,N_9757);
nand UO_661 (O_661,N_9973,N_9694);
and UO_662 (O_662,N_9595,N_9980);
nor UO_663 (O_663,N_9766,N_9636);
and UO_664 (O_664,N_9882,N_9521);
nand UO_665 (O_665,N_9578,N_9656);
or UO_666 (O_666,N_9823,N_9734);
or UO_667 (O_667,N_9586,N_9698);
nor UO_668 (O_668,N_9909,N_9919);
nor UO_669 (O_669,N_9681,N_9900);
or UO_670 (O_670,N_9774,N_9581);
nand UO_671 (O_671,N_9927,N_9507);
and UO_672 (O_672,N_9621,N_9514);
and UO_673 (O_673,N_9802,N_9509);
or UO_674 (O_674,N_9862,N_9685);
or UO_675 (O_675,N_9636,N_9533);
and UO_676 (O_676,N_9876,N_9591);
and UO_677 (O_677,N_9719,N_9553);
or UO_678 (O_678,N_9824,N_9609);
nor UO_679 (O_679,N_9698,N_9527);
or UO_680 (O_680,N_9850,N_9764);
nand UO_681 (O_681,N_9849,N_9588);
and UO_682 (O_682,N_9708,N_9970);
nand UO_683 (O_683,N_9551,N_9811);
or UO_684 (O_684,N_9843,N_9766);
nor UO_685 (O_685,N_9667,N_9809);
or UO_686 (O_686,N_9873,N_9705);
and UO_687 (O_687,N_9907,N_9738);
or UO_688 (O_688,N_9764,N_9777);
nor UO_689 (O_689,N_9992,N_9990);
nand UO_690 (O_690,N_9645,N_9890);
nand UO_691 (O_691,N_9622,N_9931);
and UO_692 (O_692,N_9999,N_9914);
nor UO_693 (O_693,N_9667,N_9540);
nand UO_694 (O_694,N_9775,N_9748);
and UO_695 (O_695,N_9850,N_9873);
or UO_696 (O_696,N_9974,N_9876);
nand UO_697 (O_697,N_9644,N_9776);
nor UO_698 (O_698,N_9559,N_9527);
and UO_699 (O_699,N_9644,N_9974);
and UO_700 (O_700,N_9728,N_9607);
nor UO_701 (O_701,N_9882,N_9615);
nand UO_702 (O_702,N_9760,N_9731);
or UO_703 (O_703,N_9947,N_9948);
nor UO_704 (O_704,N_9506,N_9981);
nand UO_705 (O_705,N_9955,N_9813);
nand UO_706 (O_706,N_9843,N_9515);
nand UO_707 (O_707,N_9796,N_9525);
and UO_708 (O_708,N_9691,N_9812);
or UO_709 (O_709,N_9551,N_9970);
xor UO_710 (O_710,N_9538,N_9870);
and UO_711 (O_711,N_9627,N_9954);
nand UO_712 (O_712,N_9949,N_9805);
nand UO_713 (O_713,N_9895,N_9774);
or UO_714 (O_714,N_9983,N_9940);
nor UO_715 (O_715,N_9963,N_9820);
nand UO_716 (O_716,N_9682,N_9949);
or UO_717 (O_717,N_9541,N_9703);
or UO_718 (O_718,N_9791,N_9883);
xor UO_719 (O_719,N_9934,N_9890);
nand UO_720 (O_720,N_9512,N_9746);
nand UO_721 (O_721,N_9530,N_9883);
nor UO_722 (O_722,N_9790,N_9614);
nand UO_723 (O_723,N_9555,N_9631);
or UO_724 (O_724,N_9877,N_9694);
nand UO_725 (O_725,N_9824,N_9555);
or UO_726 (O_726,N_9981,N_9918);
nor UO_727 (O_727,N_9673,N_9656);
nand UO_728 (O_728,N_9505,N_9829);
and UO_729 (O_729,N_9817,N_9827);
and UO_730 (O_730,N_9862,N_9921);
or UO_731 (O_731,N_9873,N_9687);
and UO_732 (O_732,N_9708,N_9839);
nor UO_733 (O_733,N_9675,N_9939);
xnor UO_734 (O_734,N_9968,N_9570);
nor UO_735 (O_735,N_9953,N_9926);
and UO_736 (O_736,N_9828,N_9972);
nand UO_737 (O_737,N_9854,N_9667);
nor UO_738 (O_738,N_9725,N_9835);
or UO_739 (O_739,N_9701,N_9583);
nor UO_740 (O_740,N_9747,N_9904);
and UO_741 (O_741,N_9790,N_9554);
nor UO_742 (O_742,N_9740,N_9579);
or UO_743 (O_743,N_9748,N_9619);
nand UO_744 (O_744,N_9504,N_9548);
nor UO_745 (O_745,N_9994,N_9513);
and UO_746 (O_746,N_9765,N_9863);
or UO_747 (O_747,N_9659,N_9830);
nand UO_748 (O_748,N_9943,N_9538);
nand UO_749 (O_749,N_9832,N_9961);
nor UO_750 (O_750,N_9815,N_9897);
and UO_751 (O_751,N_9676,N_9526);
nor UO_752 (O_752,N_9503,N_9888);
or UO_753 (O_753,N_9703,N_9933);
xor UO_754 (O_754,N_9744,N_9728);
nand UO_755 (O_755,N_9783,N_9970);
nor UO_756 (O_756,N_9957,N_9925);
nor UO_757 (O_757,N_9626,N_9739);
nand UO_758 (O_758,N_9570,N_9524);
nor UO_759 (O_759,N_9577,N_9512);
and UO_760 (O_760,N_9774,N_9745);
xnor UO_761 (O_761,N_9589,N_9927);
or UO_762 (O_762,N_9631,N_9999);
nand UO_763 (O_763,N_9605,N_9566);
and UO_764 (O_764,N_9944,N_9829);
and UO_765 (O_765,N_9512,N_9862);
and UO_766 (O_766,N_9905,N_9669);
nand UO_767 (O_767,N_9577,N_9610);
nand UO_768 (O_768,N_9707,N_9768);
xnor UO_769 (O_769,N_9945,N_9696);
nor UO_770 (O_770,N_9935,N_9681);
nor UO_771 (O_771,N_9883,N_9671);
and UO_772 (O_772,N_9995,N_9509);
or UO_773 (O_773,N_9559,N_9867);
or UO_774 (O_774,N_9657,N_9720);
or UO_775 (O_775,N_9975,N_9985);
nand UO_776 (O_776,N_9542,N_9885);
nand UO_777 (O_777,N_9981,N_9931);
xor UO_778 (O_778,N_9744,N_9601);
nor UO_779 (O_779,N_9907,N_9805);
or UO_780 (O_780,N_9899,N_9946);
nor UO_781 (O_781,N_9881,N_9729);
or UO_782 (O_782,N_9835,N_9729);
nor UO_783 (O_783,N_9778,N_9895);
or UO_784 (O_784,N_9633,N_9533);
nand UO_785 (O_785,N_9822,N_9522);
nand UO_786 (O_786,N_9656,N_9571);
nor UO_787 (O_787,N_9572,N_9786);
nand UO_788 (O_788,N_9961,N_9800);
or UO_789 (O_789,N_9931,N_9587);
or UO_790 (O_790,N_9781,N_9733);
nor UO_791 (O_791,N_9586,N_9548);
and UO_792 (O_792,N_9547,N_9943);
nor UO_793 (O_793,N_9687,N_9915);
or UO_794 (O_794,N_9626,N_9584);
nor UO_795 (O_795,N_9850,N_9631);
or UO_796 (O_796,N_9985,N_9516);
nor UO_797 (O_797,N_9541,N_9562);
and UO_798 (O_798,N_9767,N_9719);
or UO_799 (O_799,N_9605,N_9701);
nor UO_800 (O_800,N_9803,N_9833);
and UO_801 (O_801,N_9803,N_9796);
and UO_802 (O_802,N_9719,N_9638);
and UO_803 (O_803,N_9548,N_9817);
nor UO_804 (O_804,N_9889,N_9902);
nor UO_805 (O_805,N_9622,N_9826);
and UO_806 (O_806,N_9789,N_9995);
or UO_807 (O_807,N_9986,N_9985);
or UO_808 (O_808,N_9688,N_9894);
and UO_809 (O_809,N_9731,N_9637);
nor UO_810 (O_810,N_9974,N_9712);
and UO_811 (O_811,N_9928,N_9701);
and UO_812 (O_812,N_9997,N_9563);
and UO_813 (O_813,N_9916,N_9901);
or UO_814 (O_814,N_9862,N_9628);
nand UO_815 (O_815,N_9995,N_9887);
nand UO_816 (O_816,N_9622,N_9942);
and UO_817 (O_817,N_9614,N_9824);
nand UO_818 (O_818,N_9522,N_9587);
nor UO_819 (O_819,N_9664,N_9998);
nor UO_820 (O_820,N_9709,N_9934);
nor UO_821 (O_821,N_9774,N_9689);
and UO_822 (O_822,N_9663,N_9766);
nor UO_823 (O_823,N_9753,N_9716);
nor UO_824 (O_824,N_9577,N_9824);
nor UO_825 (O_825,N_9558,N_9639);
and UO_826 (O_826,N_9693,N_9907);
nor UO_827 (O_827,N_9982,N_9593);
nor UO_828 (O_828,N_9793,N_9648);
or UO_829 (O_829,N_9585,N_9544);
and UO_830 (O_830,N_9938,N_9719);
nor UO_831 (O_831,N_9580,N_9637);
or UO_832 (O_832,N_9802,N_9713);
nor UO_833 (O_833,N_9753,N_9831);
and UO_834 (O_834,N_9952,N_9825);
xor UO_835 (O_835,N_9502,N_9684);
nor UO_836 (O_836,N_9828,N_9645);
and UO_837 (O_837,N_9958,N_9738);
nand UO_838 (O_838,N_9963,N_9870);
and UO_839 (O_839,N_9989,N_9879);
or UO_840 (O_840,N_9941,N_9817);
or UO_841 (O_841,N_9803,N_9994);
and UO_842 (O_842,N_9501,N_9787);
nor UO_843 (O_843,N_9656,N_9663);
nor UO_844 (O_844,N_9792,N_9724);
or UO_845 (O_845,N_9782,N_9849);
or UO_846 (O_846,N_9761,N_9825);
nand UO_847 (O_847,N_9949,N_9988);
and UO_848 (O_848,N_9510,N_9844);
and UO_849 (O_849,N_9996,N_9735);
nand UO_850 (O_850,N_9679,N_9764);
xnor UO_851 (O_851,N_9710,N_9555);
nand UO_852 (O_852,N_9556,N_9791);
nor UO_853 (O_853,N_9849,N_9652);
nand UO_854 (O_854,N_9594,N_9839);
or UO_855 (O_855,N_9503,N_9779);
nor UO_856 (O_856,N_9569,N_9514);
nand UO_857 (O_857,N_9968,N_9996);
nor UO_858 (O_858,N_9692,N_9976);
nand UO_859 (O_859,N_9536,N_9911);
or UO_860 (O_860,N_9796,N_9559);
xnor UO_861 (O_861,N_9715,N_9860);
nor UO_862 (O_862,N_9739,N_9502);
nor UO_863 (O_863,N_9686,N_9827);
or UO_864 (O_864,N_9747,N_9518);
and UO_865 (O_865,N_9522,N_9708);
nor UO_866 (O_866,N_9971,N_9800);
or UO_867 (O_867,N_9932,N_9838);
nor UO_868 (O_868,N_9862,N_9632);
and UO_869 (O_869,N_9768,N_9807);
nand UO_870 (O_870,N_9789,N_9815);
or UO_871 (O_871,N_9648,N_9567);
nor UO_872 (O_872,N_9825,N_9702);
and UO_873 (O_873,N_9519,N_9742);
and UO_874 (O_874,N_9706,N_9781);
or UO_875 (O_875,N_9692,N_9853);
and UO_876 (O_876,N_9915,N_9662);
nand UO_877 (O_877,N_9956,N_9549);
xnor UO_878 (O_878,N_9900,N_9868);
and UO_879 (O_879,N_9573,N_9725);
xor UO_880 (O_880,N_9873,N_9684);
and UO_881 (O_881,N_9631,N_9560);
nand UO_882 (O_882,N_9811,N_9822);
nand UO_883 (O_883,N_9811,N_9876);
and UO_884 (O_884,N_9633,N_9884);
xor UO_885 (O_885,N_9514,N_9877);
nand UO_886 (O_886,N_9716,N_9894);
or UO_887 (O_887,N_9835,N_9982);
nor UO_888 (O_888,N_9578,N_9920);
nand UO_889 (O_889,N_9514,N_9703);
or UO_890 (O_890,N_9867,N_9898);
nand UO_891 (O_891,N_9874,N_9942);
or UO_892 (O_892,N_9951,N_9654);
or UO_893 (O_893,N_9583,N_9847);
xnor UO_894 (O_894,N_9894,N_9761);
nor UO_895 (O_895,N_9637,N_9516);
nor UO_896 (O_896,N_9503,N_9519);
or UO_897 (O_897,N_9665,N_9579);
and UO_898 (O_898,N_9645,N_9817);
nor UO_899 (O_899,N_9573,N_9522);
nor UO_900 (O_900,N_9706,N_9809);
or UO_901 (O_901,N_9778,N_9696);
nand UO_902 (O_902,N_9769,N_9859);
nand UO_903 (O_903,N_9520,N_9903);
nand UO_904 (O_904,N_9998,N_9662);
nand UO_905 (O_905,N_9859,N_9688);
nor UO_906 (O_906,N_9773,N_9735);
xnor UO_907 (O_907,N_9638,N_9843);
nand UO_908 (O_908,N_9693,N_9623);
or UO_909 (O_909,N_9679,N_9938);
nand UO_910 (O_910,N_9612,N_9896);
nand UO_911 (O_911,N_9953,N_9664);
nand UO_912 (O_912,N_9809,N_9880);
or UO_913 (O_913,N_9970,N_9895);
and UO_914 (O_914,N_9674,N_9694);
and UO_915 (O_915,N_9583,N_9921);
nand UO_916 (O_916,N_9602,N_9860);
nand UO_917 (O_917,N_9957,N_9768);
nor UO_918 (O_918,N_9862,N_9709);
xnor UO_919 (O_919,N_9851,N_9894);
nand UO_920 (O_920,N_9624,N_9686);
or UO_921 (O_921,N_9609,N_9595);
and UO_922 (O_922,N_9720,N_9886);
and UO_923 (O_923,N_9891,N_9509);
and UO_924 (O_924,N_9614,N_9985);
xor UO_925 (O_925,N_9725,N_9657);
nor UO_926 (O_926,N_9794,N_9578);
and UO_927 (O_927,N_9529,N_9672);
or UO_928 (O_928,N_9749,N_9890);
nand UO_929 (O_929,N_9834,N_9712);
and UO_930 (O_930,N_9908,N_9666);
and UO_931 (O_931,N_9975,N_9752);
nand UO_932 (O_932,N_9942,N_9978);
nor UO_933 (O_933,N_9582,N_9897);
or UO_934 (O_934,N_9668,N_9569);
and UO_935 (O_935,N_9534,N_9771);
and UO_936 (O_936,N_9937,N_9842);
and UO_937 (O_937,N_9615,N_9517);
nand UO_938 (O_938,N_9871,N_9805);
nor UO_939 (O_939,N_9552,N_9629);
and UO_940 (O_940,N_9974,N_9636);
or UO_941 (O_941,N_9738,N_9570);
nor UO_942 (O_942,N_9600,N_9880);
nand UO_943 (O_943,N_9540,N_9655);
nand UO_944 (O_944,N_9771,N_9698);
nand UO_945 (O_945,N_9996,N_9954);
or UO_946 (O_946,N_9595,N_9722);
or UO_947 (O_947,N_9927,N_9707);
and UO_948 (O_948,N_9514,N_9676);
or UO_949 (O_949,N_9912,N_9686);
and UO_950 (O_950,N_9523,N_9939);
nor UO_951 (O_951,N_9563,N_9691);
nor UO_952 (O_952,N_9996,N_9744);
and UO_953 (O_953,N_9570,N_9576);
nand UO_954 (O_954,N_9575,N_9635);
or UO_955 (O_955,N_9626,N_9545);
or UO_956 (O_956,N_9773,N_9503);
nor UO_957 (O_957,N_9558,N_9918);
nor UO_958 (O_958,N_9928,N_9710);
or UO_959 (O_959,N_9919,N_9518);
or UO_960 (O_960,N_9593,N_9763);
nor UO_961 (O_961,N_9599,N_9548);
nor UO_962 (O_962,N_9705,N_9993);
nand UO_963 (O_963,N_9907,N_9541);
nor UO_964 (O_964,N_9729,N_9889);
nor UO_965 (O_965,N_9908,N_9979);
nor UO_966 (O_966,N_9971,N_9780);
and UO_967 (O_967,N_9913,N_9977);
or UO_968 (O_968,N_9619,N_9798);
and UO_969 (O_969,N_9691,N_9753);
and UO_970 (O_970,N_9560,N_9674);
or UO_971 (O_971,N_9923,N_9812);
or UO_972 (O_972,N_9843,N_9906);
nand UO_973 (O_973,N_9622,N_9661);
nor UO_974 (O_974,N_9850,N_9544);
nor UO_975 (O_975,N_9571,N_9608);
nand UO_976 (O_976,N_9519,N_9893);
nand UO_977 (O_977,N_9763,N_9818);
nand UO_978 (O_978,N_9519,N_9747);
and UO_979 (O_979,N_9570,N_9648);
or UO_980 (O_980,N_9730,N_9954);
and UO_981 (O_981,N_9612,N_9943);
nor UO_982 (O_982,N_9945,N_9684);
or UO_983 (O_983,N_9562,N_9673);
nor UO_984 (O_984,N_9546,N_9655);
nor UO_985 (O_985,N_9621,N_9887);
or UO_986 (O_986,N_9682,N_9890);
and UO_987 (O_987,N_9639,N_9973);
and UO_988 (O_988,N_9833,N_9783);
or UO_989 (O_989,N_9686,N_9553);
nand UO_990 (O_990,N_9753,N_9906);
and UO_991 (O_991,N_9530,N_9662);
and UO_992 (O_992,N_9954,N_9856);
or UO_993 (O_993,N_9916,N_9923);
and UO_994 (O_994,N_9807,N_9518);
and UO_995 (O_995,N_9785,N_9903);
or UO_996 (O_996,N_9545,N_9797);
and UO_997 (O_997,N_9528,N_9931);
nand UO_998 (O_998,N_9649,N_9820);
and UO_999 (O_999,N_9946,N_9687);
or UO_1000 (O_1000,N_9569,N_9560);
nand UO_1001 (O_1001,N_9870,N_9628);
nor UO_1002 (O_1002,N_9502,N_9898);
or UO_1003 (O_1003,N_9851,N_9809);
and UO_1004 (O_1004,N_9514,N_9576);
nand UO_1005 (O_1005,N_9900,N_9556);
nand UO_1006 (O_1006,N_9820,N_9510);
nor UO_1007 (O_1007,N_9954,N_9869);
and UO_1008 (O_1008,N_9606,N_9781);
and UO_1009 (O_1009,N_9774,N_9848);
nor UO_1010 (O_1010,N_9990,N_9854);
nor UO_1011 (O_1011,N_9837,N_9931);
nor UO_1012 (O_1012,N_9648,N_9848);
nand UO_1013 (O_1013,N_9734,N_9868);
nand UO_1014 (O_1014,N_9560,N_9798);
and UO_1015 (O_1015,N_9649,N_9859);
nand UO_1016 (O_1016,N_9598,N_9616);
xnor UO_1017 (O_1017,N_9552,N_9957);
nand UO_1018 (O_1018,N_9794,N_9999);
nor UO_1019 (O_1019,N_9737,N_9673);
nor UO_1020 (O_1020,N_9737,N_9846);
and UO_1021 (O_1021,N_9751,N_9595);
xor UO_1022 (O_1022,N_9618,N_9506);
and UO_1023 (O_1023,N_9737,N_9732);
nor UO_1024 (O_1024,N_9876,N_9785);
nand UO_1025 (O_1025,N_9518,N_9931);
and UO_1026 (O_1026,N_9782,N_9866);
and UO_1027 (O_1027,N_9678,N_9852);
nand UO_1028 (O_1028,N_9582,N_9845);
nand UO_1029 (O_1029,N_9773,N_9972);
and UO_1030 (O_1030,N_9857,N_9704);
and UO_1031 (O_1031,N_9664,N_9840);
nand UO_1032 (O_1032,N_9879,N_9998);
and UO_1033 (O_1033,N_9853,N_9500);
or UO_1034 (O_1034,N_9937,N_9813);
and UO_1035 (O_1035,N_9654,N_9539);
nand UO_1036 (O_1036,N_9751,N_9606);
and UO_1037 (O_1037,N_9523,N_9618);
or UO_1038 (O_1038,N_9912,N_9887);
or UO_1039 (O_1039,N_9638,N_9916);
nor UO_1040 (O_1040,N_9791,N_9957);
nor UO_1041 (O_1041,N_9666,N_9507);
nand UO_1042 (O_1042,N_9511,N_9695);
nand UO_1043 (O_1043,N_9557,N_9711);
nor UO_1044 (O_1044,N_9972,N_9844);
nor UO_1045 (O_1045,N_9578,N_9692);
or UO_1046 (O_1046,N_9761,N_9688);
and UO_1047 (O_1047,N_9732,N_9657);
nor UO_1048 (O_1048,N_9777,N_9599);
nand UO_1049 (O_1049,N_9715,N_9944);
nand UO_1050 (O_1050,N_9515,N_9638);
and UO_1051 (O_1051,N_9721,N_9808);
nor UO_1052 (O_1052,N_9622,N_9989);
and UO_1053 (O_1053,N_9559,N_9902);
nor UO_1054 (O_1054,N_9520,N_9630);
nor UO_1055 (O_1055,N_9617,N_9768);
nor UO_1056 (O_1056,N_9637,N_9563);
nor UO_1057 (O_1057,N_9682,N_9558);
nand UO_1058 (O_1058,N_9545,N_9817);
or UO_1059 (O_1059,N_9665,N_9982);
nor UO_1060 (O_1060,N_9673,N_9964);
and UO_1061 (O_1061,N_9562,N_9909);
nor UO_1062 (O_1062,N_9636,N_9911);
or UO_1063 (O_1063,N_9589,N_9649);
or UO_1064 (O_1064,N_9521,N_9865);
nor UO_1065 (O_1065,N_9896,N_9621);
nor UO_1066 (O_1066,N_9756,N_9747);
or UO_1067 (O_1067,N_9604,N_9858);
or UO_1068 (O_1068,N_9720,N_9958);
nand UO_1069 (O_1069,N_9828,N_9970);
nand UO_1070 (O_1070,N_9947,N_9642);
xor UO_1071 (O_1071,N_9932,N_9721);
or UO_1072 (O_1072,N_9783,N_9591);
or UO_1073 (O_1073,N_9624,N_9566);
and UO_1074 (O_1074,N_9506,N_9754);
nand UO_1075 (O_1075,N_9784,N_9987);
or UO_1076 (O_1076,N_9559,N_9546);
nand UO_1077 (O_1077,N_9969,N_9895);
nor UO_1078 (O_1078,N_9800,N_9686);
and UO_1079 (O_1079,N_9954,N_9786);
and UO_1080 (O_1080,N_9701,N_9507);
or UO_1081 (O_1081,N_9874,N_9933);
nor UO_1082 (O_1082,N_9533,N_9860);
or UO_1083 (O_1083,N_9774,N_9585);
nand UO_1084 (O_1084,N_9896,N_9644);
and UO_1085 (O_1085,N_9745,N_9887);
nand UO_1086 (O_1086,N_9521,N_9958);
nand UO_1087 (O_1087,N_9921,N_9586);
or UO_1088 (O_1088,N_9685,N_9776);
nor UO_1089 (O_1089,N_9730,N_9690);
nand UO_1090 (O_1090,N_9997,N_9680);
or UO_1091 (O_1091,N_9860,N_9516);
and UO_1092 (O_1092,N_9572,N_9588);
or UO_1093 (O_1093,N_9622,N_9534);
or UO_1094 (O_1094,N_9624,N_9935);
nand UO_1095 (O_1095,N_9671,N_9614);
nand UO_1096 (O_1096,N_9634,N_9918);
or UO_1097 (O_1097,N_9638,N_9662);
or UO_1098 (O_1098,N_9505,N_9630);
and UO_1099 (O_1099,N_9884,N_9750);
and UO_1100 (O_1100,N_9895,N_9866);
nor UO_1101 (O_1101,N_9705,N_9843);
and UO_1102 (O_1102,N_9598,N_9573);
nand UO_1103 (O_1103,N_9543,N_9640);
or UO_1104 (O_1104,N_9999,N_9824);
nand UO_1105 (O_1105,N_9756,N_9883);
nand UO_1106 (O_1106,N_9550,N_9963);
nand UO_1107 (O_1107,N_9814,N_9850);
nor UO_1108 (O_1108,N_9505,N_9599);
nor UO_1109 (O_1109,N_9970,N_9660);
nand UO_1110 (O_1110,N_9804,N_9888);
and UO_1111 (O_1111,N_9557,N_9501);
nor UO_1112 (O_1112,N_9651,N_9517);
and UO_1113 (O_1113,N_9973,N_9888);
xor UO_1114 (O_1114,N_9659,N_9967);
or UO_1115 (O_1115,N_9902,N_9972);
or UO_1116 (O_1116,N_9536,N_9566);
or UO_1117 (O_1117,N_9960,N_9598);
nand UO_1118 (O_1118,N_9679,N_9832);
and UO_1119 (O_1119,N_9954,N_9736);
nand UO_1120 (O_1120,N_9784,N_9747);
nand UO_1121 (O_1121,N_9739,N_9734);
nand UO_1122 (O_1122,N_9883,N_9738);
nor UO_1123 (O_1123,N_9575,N_9651);
and UO_1124 (O_1124,N_9903,N_9631);
nor UO_1125 (O_1125,N_9779,N_9630);
nand UO_1126 (O_1126,N_9837,N_9976);
or UO_1127 (O_1127,N_9615,N_9771);
or UO_1128 (O_1128,N_9802,N_9769);
and UO_1129 (O_1129,N_9672,N_9957);
xnor UO_1130 (O_1130,N_9767,N_9595);
nand UO_1131 (O_1131,N_9804,N_9570);
and UO_1132 (O_1132,N_9985,N_9701);
or UO_1133 (O_1133,N_9642,N_9788);
and UO_1134 (O_1134,N_9898,N_9593);
and UO_1135 (O_1135,N_9601,N_9518);
nand UO_1136 (O_1136,N_9545,N_9983);
nor UO_1137 (O_1137,N_9997,N_9643);
and UO_1138 (O_1138,N_9705,N_9582);
or UO_1139 (O_1139,N_9981,N_9830);
nor UO_1140 (O_1140,N_9924,N_9737);
and UO_1141 (O_1141,N_9664,N_9686);
nor UO_1142 (O_1142,N_9883,N_9949);
nor UO_1143 (O_1143,N_9727,N_9882);
or UO_1144 (O_1144,N_9937,N_9762);
and UO_1145 (O_1145,N_9932,N_9517);
or UO_1146 (O_1146,N_9506,N_9998);
nor UO_1147 (O_1147,N_9871,N_9916);
xnor UO_1148 (O_1148,N_9523,N_9856);
or UO_1149 (O_1149,N_9561,N_9827);
or UO_1150 (O_1150,N_9831,N_9703);
nand UO_1151 (O_1151,N_9756,N_9931);
and UO_1152 (O_1152,N_9798,N_9952);
and UO_1153 (O_1153,N_9995,N_9996);
nand UO_1154 (O_1154,N_9667,N_9538);
or UO_1155 (O_1155,N_9501,N_9781);
nand UO_1156 (O_1156,N_9512,N_9670);
xnor UO_1157 (O_1157,N_9724,N_9925);
nor UO_1158 (O_1158,N_9553,N_9525);
nor UO_1159 (O_1159,N_9748,N_9526);
and UO_1160 (O_1160,N_9637,N_9632);
or UO_1161 (O_1161,N_9987,N_9915);
and UO_1162 (O_1162,N_9621,N_9789);
and UO_1163 (O_1163,N_9615,N_9996);
or UO_1164 (O_1164,N_9775,N_9938);
or UO_1165 (O_1165,N_9513,N_9634);
or UO_1166 (O_1166,N_9706,N_9512);
nand UO_1167 (O_1167,N_9770,N_9629);
nor UO_1168 (O_1168,N_9618,N_9663);
and UO_1169 (O_1169,N_9858,N_9643);
or UO_1170 (O_1170,N_9815,N_9811);
and UO_1171 (O_1171,N_9692,N_9500);
nor UO_1172 (O_1172,N_9681,N_9732);
and UO_1173 (O_1173,N_9891,N_9784);
and UO_1174 (O_1174,N_9625,N_9616);
nor UO_1175 (O_1175,N_9845,N_9504);
or UO_1176 (O_1176,N_9533,N_9996);
and UO_1177 (O_1177,N_9666,N_9746);
or UO_1178 (O_1178,N_9549,N_9691);
and UO_1179 (O_1179,N_9912,N_9609);
nor UO_1180 (O_1180,N_9793,N_9520);
and UO_1181 (O_1181,N_9541,N_9769);
nor UO_1182 (O_1182,N_9781,N_9960);
and UO_1183 (O_1183,N_9655,N_9828);
nor UO_1184 (O_1184,N_9795,N_9629);
nand UO_1185 (O_1185,N_9822,N_9657);
or UO_1186 (O_1186,N_9576,N_9754);
nor UO_1187 (O_1187,N_9882,N_9536);
and UO_1188 (O_1188,N_9942,N_9524);
and UO_1189 (O_1189,N_9784,N_9758);
nand UO_1190 (O_1190,N_9663,N_9910);
and UO_1191 (O_1191,N_9976,N_9537);
nand UO_1192 (O_1192,N_9625,N_9538);
and UO_1193 (O_1193,N_9815,N_9837);
nand UO_1194 (O_1194,N_9894,N_9546);
or UO_1195 (O_1195,N_9731,N_9516);
xnor UO_1196 (O_1196,N_9732,N_9714);
and UO_1197 (O_1197,N_9619,N_9912);
or UO_1198 (O_1198,N_9632,N_9966);
nand UO_1199 (O_1199,N_9982,N_9599);
xor UO_1200 (O_1200,N_9702,N_9669);
nand UO_1201 (O_1201,N_9761,N_9802);
nor UO_1202 (O_1202,N_9853,N_9767);
and UO_1203 (O_1203,N_9877,N_9770);
or UO_1204 (O_1204,N_9819,N_9579);
nor UO_1205 (O_1205,N_9539,N_9803);
nor UO_1206 (O_1206,N_9836,N_9744);
and UO_1207 (O_1207,N_9594,N_9912);
and UO_1208 (O_1208,N_9978,N_9619);
and UO_1209 (O_1209,N_9638,N_9692);
and UO_1210 (O_1210,N_9681,N_9837);
and UO_1211 (O_1211,N_9867,N_9505);
nand UO_1212 (O_1212,N_9623,N_9994);
nand UO_1213 (O_1213,N_9563,N_9551);
and UO_1214 (O_1214,N_9837,N_9842);
and UO_1215 (O_1215,N_9573,N_9949);
or UO_1216 (O_1216,N_9764,N_9883);
and UO_1217 (O_1217,N_9727,N_9916);
or UO_1218 (O_1218,N_9769,N_9685);
nor UO_1219 (O_1219,N_9743,N_9532);
nor UO_1220 (O_1220,N_9747,N_9659);
or UO_1221 (O_1221,N_9731,N_9912);
xnor UO_1222 (O_1222,N_9872,N_9584);
and UO_1223 (O_1223,N_9604,N_9927);
or UO_1224 (O_1224,N_9650,N_9871);
and UO_1225 (O_1225,N_9992,N_9750);
xor UO_1226 (O_1226,N_9805,N_9881);
and UO_1227 (O_1227,N_9600,N_9764);
nand UO_1228 (O_1228,N_9750,N_9742);
nand UO_1229 (O_1229,N_9708,N_9733);
or UO_1230 (O_1230,N_9950,N_9594);
or UO_1231 (O_1231,N_9641,N_9653);
and UO_1232 (O_1232,N_9704,N_9750);
or UO_1233 (O_1233,N_9672,N_9699);
or UO_1234 (O_1234,N_9910,N_9984);
nand UO_1235 (O_1235,N_9982,N_9639);
nand UO_1236 (O_1236,N_9517,N_9906);
nand UO_1237 (O_1237,N_9712,N_9964);
and UO_1238 (O_1238,N_9657,N_9521);
or UO_1239 (O_1239,N_9603,N_9535);
nor UO_1240 (O_1240,N_9862,N_9719);
or UO_1241 (O_1241,N_9816,N_9556);
or UO_1242 (O_1242,N_9575,N_9875);
and UO_1243 (O_1243,N_9582,N_9604);
nor UO_1244 (O_1244,N_9881,N_9565);
nor UO_1245 (O_1245,N_9894,N_9517);
nand UO_1246 (O_1246,N_9609,N_9957);
nor UO_1247 (O_1247,N_9625,N_9663);
nand UO_1248 (O_1248,N_9967,N_9526);
and UO_1249 (O_1249,N_9681,N_9809);
nand UO_1250 (O_1250,N_9972,N_9648);
nor UO_1251 (O_1251,N_9907,N_9850);
nor UO_1252 (O_1252,N_9583,N_9507);
and UO_1253 (O_1253,N_9944,N_9761);
and UO_1254 (O_1254,N_9608,N_9891);
or UO_1255 (O_1255,N_9737,N_9660);
or UO_1256 (O_1256,N_9942,N_9728);
nand UO_1257 (O_1257,N_9502,N_9825);
nor UO_1258 (O_1258,N_9887,N_9860);
nor UO_1259 (O_1259,N_9538,N_9741);
nor UO_1260 (O_1260,N_9966,N_9621);
nor UO_1261 (O_1261,N_9643,N_9995);
nor UO_1262 (O_1262,N_9556,N_9594);
nor UO_1263 (O_1263,N_9576,N_9531);
or UO_1264 (O_1264,N_9728,N_9673);
nand UO_1265 (O_1265,N_9743,N_9718);
and UO_1266 (O_1266,N_9670,N_9680);
nor UO_1267 (O_1267,N_9833,N_9575);
nor UO_1268 (O_1268,N_9997,N_9994);
or UO_1269 (O_1269,N_9516,N_9503);
nand UO_1270 (O_1270,N_9990,N_9790);
nand UO_1271 (O_1271,N_9950,N_9850);
nand UO_1272 (O_1272,N_9895,N_9636);
nand UO_1273 (O_1273,N_9575,N_9838);
nor UO_1274 (O_1274,N_9822,N_9774);
nand UO_1275 (O_1275,N_9782,N_9767);
or UO_1276 (O_1276,N_9645,N_9530);
nand UO_1277 (O_1277,N_9675,N_9904);
or UO_1278 (O_1278,N_9813,N_9583);
nor UO_1279 (O_1279,N_9597,N_9736);
nand UO_1280 (O_1280,N_9540,N_9677);
nand UO_1281 (O_1281,N_9648,N_9566);
nand UO_1282 (O_1282,N_9513,N_9923);
and UO_1283 (O_1283,N_9564,N_9983);
nor UO_1284 (O_1284,N_9971,N_9593);
nor UO_1285 (O_1285,N_9787,N_9897);
nor UO_1286 (O_1286,N_9772,N_9509);
and UO_1287 (O_1287,N_9808,N_9517);
nand UO_1288 (O_1288,N_9663,N_9751);
nand UO_1289 (O_1289,N_9857,N_9911);
nor UO_1290 (O_1290,N_9805,N_9585);
and UO_1291 (O_1291,N_9687,N_9847);
and UO_1292 (O_1292,N_9738,N_9927);
nor UO_1293 (O_1293,N_9982,N_9752);
or UO_1294 (O_1294,N_9886,N_9962);
and UO_1295 (O_1295,N_9690,N_9994);
or UO_1296 (O_1296,N_9783,N_9716);
nand UO_1297 (O_1297,N_9577,N_9533);
and UO_1298 (O_1298,N_9660,N_9632);
or UO_1299 (O_1299,N_9654,N_9927);
and UO_1300 (O_1300,N_9615,N_9902);
nand UO_1301 (O_1301,N_9800,N_9739);
or UO_1302 (O_1302,N_9676,N_9607);
or UO_1303 (O_1303,N_9644,N_9628);
and UO_1304 (O_1304,N_9781,N_9597);
nand UO_1305 (O_1305,N_9923,N_9811);
or UO_1306 (O_1306,N_9687,N_9775);
and UO_1307 (O_1307,N_9699,N_9501);
nand UO_1308 (O_1308,N_9901,N_9580);
and UO_1309 (O_1309,N_9946,N_9652);
nand UO_1310 (O_1310,N_9727,N_9583);
nor UO_1311 (O_1311,N_9713,N_9625);
nand UO_1312 (O_1312,N_9877,N_9964);
nor UO_1313 (O_1313,N_9952,N_9886);
nand UO_1314 (O_1314,N_9538,N_9504);
or UO_1315 (O_1315,N_9575,N_9583);
nand UO_1316 (O_1316,N_9537,N_9515);
nor UO_1317 (O_1317,N_9639,N_9900);
or UO_1318 (O_1318,N_9983,N_9980);
or UO_1319 (O_1319,N_9618,N_9592);
xnor UO_1320 (O_1320,N_9975,N_9504);
or UO_1321 (O_1321,N_9582,N_9932);
nor UO_1322 (O_1322,N_9972,N_9882);
or UO_1323 (O_1323,N_9705,N_9952);
nor UO_1324 (O_1324,N_9786,N_9711);
and UO_1325 (O_1325,N_9819,N_9933);
nand UO_1326 (O_1326,N_9552,N_9769);
nor UO_1327 (O_1327,N_9864,N_9859);
and UO_1328 (O_1328,N_9505,N_9677);
nand UO_1329 (O_1329,N_9657,N_9863);
nor UO_1330 (O_1330,N_9624,N_9868);
or UO_1331 (O_1331,N_9851,N_9791);
nor UO_1332 (O_1332,N_9664,N_9804);
nor UO_1333 (O_1333,N_9876,N_9970);
or UO_1334 (O_1334,N_9555,N_9950);
or UO_1335 (O_1335,N_9885,N_9690);
or UO_1336 (O_1336,N_9804,N_9886);
or UO_1337 (O_1337,N_9969,N_9797);
or UO_1338 (O_1338,N_9644,N_9742);
nor UO_1339 (O_1339,N_9711,N_9713);
or UO_1340 (O_1340,N_9704,N_9979);
and UO_1341 (O_1341,N_9662,N_9804);
or UO_1342 (O_1342,N_9639,N_9533);
or UO_1343 (O_1343,N_9766,N_9836);
nand UO_1344 (O_1344,N_9523,N_9934);
and UO_1345 (O_1345,N_9910,N_9504);
nand UO_1346 (O_1346,N_9929,N_9660);
nor UO_1347 (O_1347,N_9779,N_9820);
nand UO_1348 (O_1348,N_9777,N_9869);
nand UO_1349 (O_1349,N_9688,N_9635);
or UO_1350 (O_1350,N_9594,N_9828);
or UO_1351 (O_1351,N_9803,N_9515);
or UO_1352 (O_1352,N_9977,N_9878);
and UO_1353 (O_1353,N_9862,N_9873);
nand UO_1354 (O_1354,N_9883,N_9687);
nor UO_1355 (O_1355,N_9691,N_9865);
and UO_1356 (O_1356,N_9803,N_9501);
and UO_1357 (O_1357,N_9576,N_9877);
or UO_1358 (O_1358,N_9630,N_9944);
and UO_1359 (O_1359,N_9580,N_9969);
nor UO_1360 (O_1360,N_9683,N_9931);
and UO_1361 (O_1361,N_9951,N_9956);
nand UO_1362 (O_1362,N_9619,N_9797);
nor UO_1363 (O_1363,N_9638,N_9671);
and UO_1364 (O_1364,N_9874,N_9993);
and UO_1365 (O_1365,N_9925,N_9837);
and UO_1366 (O_1366,N_9992,N_9902);
nor UO_1367 (O_1367,N_9546,N_9742);
nand UO_1368 (O_1368,N_9627,N_9793);
nand UO_1369 (O_1369,N_9685,N_9991);
nor UO_1370 (O_1370,N_9700,N_9825);
nand UO_1371 (O_1371,N_9520,N_9542);
nand UO_1372 (O_1372,N_9604,N_9645);
and UO_1373 (O_1373,N_9993,N_9643);
and UO_1374 (O_1374,N_9554,N_9925);
nand UO_1375 (O_1375,N_9719,N_9702);
and UO_1376 (O_1376,N_9984,N_9669);
and UO_1377 (O_1377,N_9512,N_9810);
xor UO_1378 (O_1378,N_9977,N_9848);
nor UO_1379 (O_1379,N_9976,N_9814);
nand UO_1380 (O_1380,N_9837,N_9608);
nand UO_1381 (O_1381,N_9933,N_9666);
nand UO_1382 (O_1382,N_9680,N_9818);
nand UO_1383 (O_1383,N_9738,N_9554);
nand UO_1384 (O_1384,N_9703,N_9646);
xnor UO_1385 (O_1385,N_9892,N_9579);
nor UO_1386 (O_1386,N_9634,N_9558);
nor UO_1387 (O_1387,N_9758,N_9836);
and UO_1388 (O_1388,N_9620,N_9810);
nand UO_1389 (O_1389,N_9872,N_9810);
and UO_1390 (O_1390,N_9974,N_9952);
and UO_1391 (O_1391,N_9594,N_9792);
nor UO_1392 (O_1392,N_9681,N_9606);
xor UO_1393 (O_1393,N_9787,N_9772);
nand UO_1394 (O_1394,N_9624,N_9798);
xnor UO_1395 (O_1395,N_9945,N_9515);
nor UO_1396 (O_1396,N_9844,N_9624);
nand UO_1397 (O_1397,N_9674,N_9991);
nor UO_1398 (O_1398,N_9854,N_9515);
nor UO_1399 (O_1399,N_9916,N_9533);
and UO_1400 (O_1400,N_9710,N_9658);
or UO_1401 (O_1401,N_9760,N_9987);
or UO_1402 (O_1402,N_9537,N_9905);
and UO_1403 (O_1403,N_9546,N_9551);
and UO_1404 (O_1404,N_9555,N_9609);
and UO_1405 (O_1405,N_9915,N_9716);
nand UO_1406 (O_1406,N_9669,N_9620);
nand UO_1407 (O_1407,N_9625,N_9903);
and UO_1408 (O_1408,N_9586,N_9688);
or UO_1409 (O_1409,N_9741,N_9579);
nand UO_1410 (O_1410,N_9755,N_9920);
and UO_1411 (O_1411,N_9731,N_9568);
or UO_1412 (O_1412,N_9628,N_9807);
nor UO_1413 (O_1413,N_9832,N_9733);
nand UO_1414 (O_1414,N_9531,N_9820);
and UO_1415 (O_1415,N_9570,N_9753);
and UO_1416 (O_1416,N_9605,N_9875);
or UO_1417 (O_1417,N_9537,N_9614);
nor UO_1418 (O_1418,N_9622,N_9785);
or UO_1419 (O_1419,N_9892,N_9644);
and UO_1420 (O_1420,N_9577,N_9914);
and UO_1421 (O_1421,N_9743,N_9886);
nand UO_1422 (O_1422,N_9515,N_9987);
and UO_1423 (O_1423,N_9995,N_9688);
or UO_1424 (O_1424,N_9827,N_9778);
nand UO_1425 (O_1425,N_9824,N_9872);
nor UO_1426 (O_1426,N_9778,N_9721);
nand UO_1427 (O_1427,N_9942,N_9627);
and UO_1428 (O_1428,N_9961,N_9957);
nor UO_1429 (O_1429,N_9895,N_9938);
nor UO_1430 (O_1430,N_9703,N_9989);
or UO_1431 (O_1431,N_9638,N_9978);
and UO_1432 (O_1432,N_9913,N_9693);
nor UO_1433 (O_1433,N_9889,N_9528);
nor UO_1434 (O_1434,N_9617,N_9774);
nand UO_1435 (O_1435,N_9542,N_9796);
and UO_1436 (O_1436,N_9618,N_9884);
nor UO_1437 (O_1437,N_9734,N_9930);
nor UO_1438 (O_1438,N_9577,N_9695);
nor UO_1439 (O_1439,N_9849,N_9851);
or UO_1440 (O_1440,N_9676,N_9851);
and UO_1441 (O_1441,N_9999,N_9720);
or UO_1442 (O_1442,N_9892,N_9698);
nand UO_1443 (O_1443,N_9773,N_9757);
or UO_1444 (O_1444,N_9552,N_9900);
or UO_1445 (O_1445,N_9728,N_9510);
and UO_1446 (O_1446,N_9670,N_9672);
nor UO_1447 (O_1447,N_9770,N_9592);
and UO_1448 (O_1448,N_9694,N_9715);
nor UO_1449 (O_1449,N_9670,N_9696);
and UO_1450 (O_1450,N_9937,N_9747);
or UO_1451 (O_1451,N_9608,N_9580);
or UO_1452 (O_1452,N_9911,N_9776);
or UO_1453 (O_1453,N_9848,N_9916);
and UO_1454 (O_1454,N_9910,N_9732);
or UO_1455 (O_1455,N_9533,N_9597);
or UO_1456 (O_1456,N_9822,N_9636);
nand UO_1457 (O_1457,N_9608,N_9878);
and UO_1458 (O_1458,N_9513,N_9973);
or UO_1459 (O_1459,N_9699,N_9653);
nor UO_1460 (O_1460,N_9762,N_9666);
or UO_1461 (O_1461,N_9805,N_9547);
nand UO_1462 (O_1462,N_9746,N_9633);
and UO_1463 (O_1463,N_9707,N_9643);
nand UO_1464 (O_1464,N_9933,N_9939);
nand UO_1465 (O_1465,N_9667,N_9997);
and UO_1466 (O_1466,N_9989,N_9706);
nor UO_1467 (O_1467,N_9512,N_9545);
or UO_1468 (O_1468,N_9621,N_9993);
and UO_1469 (O_1469,N_9914,N_9916);
xor UO_1470 (O_1470,N_9542,N_9634);
nand UO_1471 (O_1471,N_9644,N_9725);
nand UO_1472 (O_1472,N_9705,N_9789);
nor UO_1473 (O_1473,N_9939,N_9998);
and UO_1474 (O_1474,N_9899,N_9572);
nor UO_1475 (O_1475,N_9679,N_9833);
nand UO_1476 (O_1476,N_9959,N_9916);
nor UO_1477 (O_1477,N_9572,N_9844);
nor UO_1478 (O_1478,N_9897,N_9921);
nor UO_1479 (O_1479,N_9542,N_9540);
xor UO_1480 (O_1480,N_9731,N_9903);
and UO_1481 (O_1481,N_9575,N_9980);
or UO_1482 (O_1482,N_9993,N_9973);
and UO_1483 (O_1483,N_9546,N_9964);
nand UO_1484 (O_1484,N_9532,N_9664);
nand UO_1485 (O_1485,N_9622,N_9666);
nor UO_1486 (O_1486,N_9727,N_9738);
nand UO_1487 (O_1487,N_9638,N_9564);
nor UO_1488 (O_1488,N_9615,N_9812);
nand UO_1489 (O_1489,N_9918,N_9723);
nor UO_1490 (O_1490,N_9995,N_9536);
nand UO_1491 (O_1491,N_9692,N_9858);
and UO_1492 (O_1492,N_9625,N_9613);
or UO_1493 (O_1493,N_9921,N_9585);
and UO_1494 (O_1494,N_9514,N_9807);
and UO_1495 (O_1495,N_9565,N_9706);
and UO_1496 (O_1496,N_9813,N_9926);
nand UO_1497 (O_1497,N_9907,N_9672);
nor UO_1498 (O_1498,N_9953,N_9698);
and UO_1499 (O_1499,N_9563,N_9842);
endmodule