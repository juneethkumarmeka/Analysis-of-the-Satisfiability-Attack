module basic_2500_25000_3000_25_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_205,In_624);
and U1 (N_1,In_1517,In_1806);
xor U2 (N_2,In_2137,In_1586);
and U3 (N_3,In_406,In_1005);
xor U4 (N_4,In_2128,In_1269);
xor U5 (N_5,In_1411,In_2294);
nor U6 (N_6,In_2317,In_1633);
or U7 (N_7,In_1379,In_1448);
and U8 (N_8,In_1964,In_1827);
nor U9 (N_9,In_1449,In_1898);
xor U10 (N_10,In_975,In_1290);
nand U11 (N_11,In_15,In_2447);
nor U12 (N_12,In_1690,In_452);
nand U13 (N_13,In_2487,In_1292);
nor U14 (N_14,In_2057,In_1276);
or U15 (N_15,In_374,In_203);
nand U16 (N_16,In_1091,In_1);
and U17 (N_17,In_2250,In_1667);
nand U18 (N_18,In_1535,In_1233);
or U19 (N_19,In_504,In_695);
nor U20 (N_20,In_653,In_1275);
nand U21 (N_21,In_332,In_2405);
xnor U22 (N_22,In_1482,In_1372);
nand U23 (N_23,In_1741,In_1953);
and U24 (N_24,In_1112,In_1610);
nor U25 (N_25,In_582,In_931);
or U26 (N_26,In_1573,In_1363);
nand U27 (N_27,In_2056,In_2013);
or U28 (N_28,In_1748,In_2088);
xor U29 (N_29,In_32,In_1859);
nand U30 (N_30,In_606,In_1049);
nand U31 (N_31,In_755,In_388);
nand U32 (N_32,In_1753,In_1862);
or U33 (N_33,In_1644,In_882);
nor U34 (N_34,In_1246,In_360);
nand U35 (N_35,In_1506,In_1696);
or U36 (N_36,In_2208,In_2174);
or U37 (N_37,In_736,In_1874);
and U38 (N_38,In_2467,In_1978);
nor U39 (N_39,In_18,In_111);
nor U40 (N_40,In_278,In_1801);
nand U41 (N_41,In_2380,In_1105);
xor U42 (N_42,In_2114,In_268);
and U43 (N_43,In_889,In_1918);
nand U44 (N_44,In_2358,In_145);
xor U45 (N_45,In_2162,In_2101);
nand U46 (N_46,In_1420,In_346);
nor U47 (N_47,In_1404,In_1832);
xor U48 (N_48,In_1323,In_1220);
or U49 (N_49,In_44,In_1103);
or U50 (N_50,In_2212,In_1254);
or U51 (N_51,In_901,In_52);
or U52 (N_52,In_2229,In_2366);
or U53 (N_53,In_1894,In_1400);
nor U54 (N_54,In_874,In_343);
xor U55 (N_55,In_519,In_2465);
nor U56 (N_56,In_982,In_1581);
and U57 (N_57,In_1468,In_1167);
nor U58 (N_58,In_2340,In_1587);
nand U59 (N_59,In_1324,In_2075);
or U60 (N_60,In_1052,In_867);
nand U61 (N_61,In_541,In_1346);
nor U62 (N_62,In_709,In_1523);
and U63 (N_63,In_121,In_2330);
or U64 (N_64,In_712,In_1335);
nand U65 (N_65,In_91,In_772);
nand U66 (N_66,In_546,In_985);
and U67 (N_67,In_2471,In_50);
or U68 (N_68,In_1933,In_2063);
xnor U69 (N_69,In_1516,In_1443);
nand U70 (N_70,In_796,In_1460);
and U71 (N_71,In_1129,In_478);
and U72 (N_72,In_690,In_2308);
xor U73 (N_73,In_1618,In_2233);
and U74 (N_74,In_1377,In_1202);
nand U75 (N_75,In_1939,In_1773);
xor U76 (N_76,In_1958,In_920);
or U77 (N_77,In_1344,In_960);
and U78 (N_78,In_253,In_1149);
nand U79 (N_79,In_1170,In_2018);
xor U80 (N_80,In_1847,In_669);
and U81 (N_81,In_34,In_1775);
and U82 (N_82,In_1876,In_2403);
or U83 (N_83,In_643,In_1023);
nor U84 (N_84,In_1382,In_2425);
nor U85 (N_85,In_2112,In_313);
nand U86 (N_86,In_2437,In_114);
or U87 (N_87,In_1118,In_1406);
nor U88 (N_88,In_2117,In_1555);
and U89 (N_89,In_836,In_2006);
or U90 (N_90,In_449,In_560);
and U91 (N_91,In_280,In_658);
and U92 (N_92,In_2498,In_498);
or U93 (N_93,In_547,In_2341);
nor U94 (N_94,In_551,In_1466);
xor U95 (N_95,In_959,In_14);
nand U96 (N_96,In_370,In_1788);
nor U97 (N_97,In_312,In_1484);
or U98 (N_98,In_688,In_1676);
nand U99 (N_99,In_414,In_1536);
and U100 (N_100,In_69,In_678);
nor U101 (N_101,In_2218,In_1194);
nor U102 (N_102,In_1424,In_1125);
xnor U103 (N_103,In_1279,In_2159);
xnor U104 (N_104,In_2352,In_711);
and U105 (N_105,In_0,In_1074);
nor U106 (N_106,In_1286,In_1139);
xor U107 (N_107,In_1645,In_774);
nor U108 (N_108,In_74,In_2316);
or U109 (N_109,In_824,In_1543);
nor U110 (N_110,In_1698,In_36);
nand U111 (N_111,In_1471,In_2066);
nor U112 (N_112,In_57,In_1765);
nor U113 (N_113,In_817,In_5);
xnor U114 (N_114,In_2153,In_483);
nand U115 (N_115,In_155,In_422);
or U116 (N_116,In_38,In_1650);
nor U117 (N_117,In_2313,In_1567);
nand U118 (N_118,In_88,In_637);
and U119 (N_119,In_123,In_2446);
or U120 (N_120,In_2043,In_1226);
nand U121 (N_121,In_1248,In_1266);
or U122 (N_122,In_380,In_101);
nor U123 (N_123,In_771,In_764);
xnor U124 (N_124,In_729,In_1879);
nand U125 (N_125,In_2203,In_1759);
xnor U126 (N_126,In_1895,In_251);
nand U127 (N_127,In_635,In_178);
nand U128 (N_128,In_375,In_1016);
nor U129 (N_129,In_1002,In_2123);
nand U130 (N_130,In_883,In_219);
xor U131 (N_131,In_2076,In_788);
nor U132 (N_132,In_130,In_1619);
xnor U133 (N_133,In_310,In_176);
xnor U134 (N_134,In_182,In_656);
and U135 (N_135,In_2016,In_1163);
and U136 (N_136,In_169,In_2111);
nand U137 (N_137,In_197,In_1176);
nand U138 (N_138,In_1467,In_2289);
nand U139 (N_139,In_1926,In_210);
or U140 (N_140,In_68,In_2125);
xnor U141 (N_141,In_1986,In_508);
nand U142 (N_142,In_723,In_2464);
nand U143 (N_143,In_1623,In_337);
nor U144 (N_144,In_282,In_2049);
or U145 (N_145,In_2299,In_2115);
xnor U146 (N_146,In_1841,In_1479);
or U147 (N_147,In_1577,In_206);
xnor U148 (N_148,In_1595,In_599);
xnor U149 (N_149,In_434,In_394);
nand U150 (N_150,In_1911,In_1080);
nand U151 (N_151,In_604,In_1844);
nor U152 (N_152,In_1205,In_1299);
nor U153 (N_153,In_482,In_953);
nor U154 (N_154,In_1602,In_1168);
nor U155 (N_155,In_2344,In_317);
and U156 (N_156,In_837,In_459);
nand U157 (N_157,In_1132,In_1849);
or U158 (N_158,In_1071,In_1124);
or U159 (N_159,In_1663,In_396);
xor U160 (N_160,In_307,In_513);
nand U161 (N_161,In_947,In_1368);
xnor U162 (N_162,In_99,In_1883);
or U163 (N_163,In_1831,In_299);
nor U164 (N_164,In_1743,In_1064);
or U165 (N_165,In_97,In_2170);
nor U166 (N_166,In_1944,In_497);
xor U167 (N_167,In_1502,In_2486);
or U168 (N_168,In_2482,In_196);
xnor U169 (N_169,In_783,In_446);
nand U170 (N_170,In_2354,In_1942);
nand U171 (N_171,In_1798,In_240);
and U172 (N_172,In_2278,In_803);
or U173 (N_173,In_2420,In_1309);
nand U174 (N_174,In_2382,In_1921);
nand U175 (N_175,In_1777,In_922);
nor U176 (N_176,In_1751,In_85);
and U177 (N_177,In_179,In_737);
and U178 (N_178,In_598,In_1902);
or U179 (N_179,In_86,In_1012);
xor U180 (N_180,In_1130,In_1814);
nand U181 (N_181,In_556,In_146);
and U182 (N_182,In_1735,In_1329);
nor U183 (N_183,In_2288,In_1558);
nand U184 (N_184,In_775,In_195);
or U185 (N_185,In_2267,In_1829);
nor U186 (N_186,In_1813,In_428);
xnor U187 (N_187,In_201,In_2182);
and U188 (N_188,In_495,In_1399);
or U189 (N_189,In_1733,In_1306);
or U190 (N_190,In_1745,In_440);
nand U191 (N_191,In_345,In_916);
xor U192 (N_192,In_42,In_1212);
and U193 (N_193,In_505,In_214);
xnor U194 (N_194,In_2244,In_2196);
or U195 (N_195,In_565,In_1004);
nand U196 (N_196,In_2434,In_1353);
and U197 (N_197,In_691,In_1010);
nand U198 (N_198,In_1960,In_1600);
xnor U199 (N_199,In_971,In_750);
nor U200 (N_200,In_651,In_1073);
nor U201 (N_201,In_256,In_2255);
xor U202 (N_202,In_1700,In_2302);
nor U203 (N_203,In_1744,In_2400);
and U204 (N_204,In_1819,In_2067);
and U205 (N_205,In_601,In_1235);
nor U206 (N_206,In_185,In_212);
and U207 (N_207,In_2413,In_2499);
or U208 (N_208,In_1247,In_1222);
xor U209 (N_209,In_190,In_144);
and U210 (N_210,In_1864,In_2161);
nand U211 (N_211,In_2284,In_825);
nand U212 (N_212,In_2239,In_1982);
xor U213 (N_213,In_1891,In_1906);
nand U214 (N_214,In_581,In_1432);
and U215 (N_215,In_2264,In_1111);
or U216 (N_216,In_1772,In_2320);
nor U217 (N_217,In_77,In_1845);
nand U218 (N_218,In_1405,In_1314);
nor U219 (N_219,In_1360,In_297);
xnor U220 (N_220,In_2453,In_1526);
nand U221 (N_221,In_827,In_262);
and U222 (N_222,In_2221,In_2107);
xnor U223 (N_223,In_7,In_845);
xnor U224 (N_224,In_1407,In_2458);
and U225 (N_225,In_1000,In_1199);
xnor U226 (N_226,In_2414,In_2324);
xnor U227 (N_227,In_1469,In_1598);
and U228 (N_228,In_671,In_104);
nand U229 (N_229,In_1626,In_1712);
or U230 (N_230,In_373,In_2444);
xnor U231 (N_231,In_910,In_2209);
nor U232 (N_232,In_743,In_1262);
nand U233 (N_233,In_237,In_131);
or U234 (N_234,In_425,In_2064);
xnor U235 (N_235,In_154,In_2065);
nand U236 (N_236,In_367,In_1380);
xor U237 (N_237,In_410,In_998);
or U238 (N_238,In_137,In_1179);
or U239 (N_239,In_892,In_1033);
nor U240 (N_240,In_2036,In_2496);
nor U241 (N_241,In_1336,In_2130);
nand U242 (N_242,In_435,In_1447);
nand U243 (N_243,In_1677,In_1968);
nand U244 (N_244,In_404,In_134);
nor U245 (N_245,In_65,In_315);
nor U246 (N_246,In_53,In_2214);
or U247 (N_247,In_2393,In_496);
xnor U248 (N_248,In_792,In_285);
nor U249 (N_249,In_879,In_1491);
nor U250 (N_250,In_600,In_23);
nand U251 (N_251,In_1983,In_1569);
and U252 (N_252,In_1590,In_1008);
and U253 (N_253,In_662,In_1685);
xor U254 (N_254,In_480,In_458);
or U255 (N_255,In_2298,In_2290);
or U256 (N_256,In_105,In_1711);
nand U257 (N_257,In_2491,In_2466);
xnor U258 (N_258,In_468,In_2004);
xnor U259 (N_259,In_1548,In_532);
nand U260 (N_260,In_2071,In_1808);
xnor U261 (N_261,In_306,In_2379);
xnor U262 (N_262,In_1823,In_1239);
or U263 (N_263,In_1320,In_1350);
nand U264 (N_264,In_1783,In_2273);
nand U265 (N_265,In_39,In_942);
and U266 (N_266,In_687,In_1349);
or U267 (N_267,In_438,In_431);
xnor U268 (N_268,In_2473,In_984);
nor U269 (N_269,In_1853,In_1617);
nor U270 (N_270,In_2483,In_1528);
nand U271 (N_271,In_194,In_925);
or U272 (N_272,In_1648,In_782);
nand U273 (N_273,In_621,In_550);
xnor U274 (N_274,In_1724,In_1295);
and U275 (N_275,In_2274,In_443);
nor U276 (N_276,In_558,In_2242);
or U277 (N_277,In_1966,In_2394);
and U278 (N_278,In_727,In_328);
nand U279 (N_279,In_1486,In_1758);
nor U280 (N_280,In_826,In_853);
or U281 (N_281,In_427,In_491);
or U282 (N_282,In_780,In_106);
xnor U283 (N_283,In_778,In_2493);
and U284 (N_284,In_2476,In_663);
nand U285 (N_285,In_1721,In_1672);
nand U286 (N_286,In_453,In_1252);
xnor U287 (N_287,In_2306,In_1452);
nand U288 (N_288,In_186,In_2178);
nand U289 (N_289,In_1385,In_6);
or U290 (N_290,In_9,In_619);
and U291 (N_291,In_56,In_1995);
xor U292 (N_292,In_2377,In_1270);
and U293 (N_293,In_433,In_1767);
or U294 (N_294,In_2364,In_1722);
nand U295 (N_295,In_2106,In_1340);
xor U296 (N_296,In_1790,In_2073);
xnor U297 (N_297,In_184,In_1305);
xor U298 (N_298,In_979,In_1422);
nand U299 (N_299,In_226,In_1375);
and U300 (N_300,In_3,In_1576);
nor U301 (N_301,In_110,In_1093);
and U302 (N_302,In_1739,In_161);
xnor U303 (N_303,In_852,In_913);
or U304 (N_304,In_2281,In_236);
or U305 (N_305,In_1734,In_2199);
nor U306 (N_306,In_704,In_76);
nor U307 (N_307,In_1531,In_151);
nor U308 (N_308,In_1656,In_1582);
and U309 (N_309,In_1583,In_1086);
xnor U310 (N_310,In_2426,In_615);
xor U311 (N_311,In_1373,In_1588);
xnor U312 (N_312,In_850,In_473);
nand U313 (N_313,In_1917,In_2353);
xnor U314 (N_314,In_518,In_2310);
xor U315 (N_315,In_2440,In_896);
nand U316 (N_316,In_230,In_397);
nor U317 (N_317,In_1024,In_109);
and U318 (N_318,In_1800,In_1161);
nand U319 (N_319,In_682,In_1760);
and U320 (N_320,In_385,In_1157);
or U321 (N_321,In_168,In_1668);
xor U322 (N_322,In_965,In_744);
or U323 (N_323,In_364,In_795);
and U324 (N_324,In_1888,In_320);
or U325 (N_325,In_1263,In_823);
nand U326 (N_326,In_1997,In_475);
nand U327 (N_327,In_2032,In_1365);
nor U328 (N_328,In_646,In_192);
xor U329 (N_329,In_2135,In_456);
or U330 (N_330,In_289,In_1723);
xor U331 (N_331,In_1857,In_1666);
and U332 (N_332,In_1768,In_1533);
nand U333 (N_333,In_1769,In_1402);
or U334 (N_334,In_1515,In_1341);
and U335 (N_335,In_1374,In_486);
nand U336 (N_336,In_333,In_2254);
nand U337 (N_337,In_1785,In_1538);
or U338 (N_338,In_2047,In_864);
xnor U339 (N_339,In_90,In_1265);
or U340 (N_340,In_1509,In_634);
nand U341 (N_341,In_1981,In_923);
xor U342 (N_342,In_542,In_2183);
nand U343 (N_343,In_1574,In_1187);
nand U344 (N_344,In_1088,In_1462);
and U345 (N_345,In_93,In_1454);
nand U346 (N_346,In_1699,In_697);
nand U347 (N_347,In_1348,In_2334);
nand U348 (N_348,In_748,In_1974);
nor U349 (N_349,In_885,In_2068);
and U350 (N_350,In_1897,In_2213);
nand U351 (N_351,In_1860,In_2042);
or U352 (N_352,In_464,In_1729);
xor U353 (N_353,In_351,In_1294);
and U354 (N_354,In_1611,In_930);
nand U355 (N_355,In_685,In_603);
nand U356 (N_356,In_1761,In_1647);
xor U357 (N_357,In_1705,In_1505);
or U358 (N_358,In_1638,In_302);
and U359 (N_359,In_1669,In_1549);
xnor U360 (N_360,In_2103,In_1090);
or U361 (N_361,In_1440,In_739);
nand U362 (N_362,In_1268,In_2205);
nand U363 (N_363,In_638,In_1094);
or U364 (N_364,In_1657,In_747);
nand U365 (N_365,In_1766,In_1629);
or U366 (N_366,In_2217,In_932);
or U367 (N_367,In_1866,In_2241);
nor U368 (N_368,In_2157,In_2030);
nor U369 (N_369,In_1027,In_602);
and U370 (N_370,In_2416,In_517);
or U371 (N_371,In_1381,In_342);
or U372 (N_372,In_978,In_399);
nor U373 (N_373,In_1909,In_1870);
nor U374 (N_374,In_2100,In_886);
or U375 (N_375,In_1259,In_1920);
nor U376 (N_376,In_2345,In_1863);
or U377 (N_377,In_158,In_200);
or U378 (N_378,In_2484,In_1355);
nand U379 (N_379,In_1654,In_862);
or U380 (N_380,In_758,In_1055);
or U381 (N_381,In_319,In_1786);
or U382 (N_382,In_2022,In_460);
xnor U383 (N_383,In_107,In_1106);
and U384 (N_384,In_2285,In_1726);
and U385 (N_385,In_2454,In_1334);
or U386 (N_386,In_1245,In_787);
xnor U387 (N_387,In_1352,In_1508);
and U388 (N_388,In_1674,In_1455);
xor U389 (N_389,In_330,In_376);
and U390 (N_390,In_790,In_501);
nand U391 (N_391,In_576,In_1433);
nor U392 (N_392,In_2045,In_605);
xor U393 (N_393,In_140,In_1316);
nand U394 (N_394,In_1196,In_187);
nor U395 (N_395,In_944,In_2169);
nor U396 (N_396,In_1211,In_1472);
xor U397 (N_397,In_2408,In_1994);
xnor U398 (N_398,In_676,In_848);
or U399 (N_399,In_171,In_325);
nor U400 (N_400,In_395,In_166);
or U401 (N_401,In_745,In_1951);
or U402 (N_402,In_991,In_1830);
and U403 (N_403,In_1755,In_1311);
or U404 (N_404,In_1571,In_2085);
nor U405 (N_405,In_4,In_2005);
xnor U406 (N_406,In_972,In_1051);
nand U407 (N_407,In_1584,In_390);
nor U408 (N_408,In_681,In_1216);
or U409 (N_409,In_2390,In_2238);
nand U410 (N_410,In_1564,In_596);
xnor U411 (N_411,In_479,In_689);
nor U412 (N_412,In_1042,In_1172);
and U413 (N_413,In_1865,In_1481);
xnor U414 (N_414,In_648,In_2488);
xor U415 (N_415,In_2104,In_647);
nor U416 (N_416,In_1274,In_1155);
xor U417 (N_417,In_1634,In_2108);
or U418 (N_418,In_846,In_2286);
nand U419 (N_419,In_629,In_820);
xor U420 (N_420,In_2146,In_1240);
nand U421 (N_421,In_1195,In_1181);
nand U422 (N_422,In_585,In_949);
and U423 (N_423,In_2432,In_350);
and U424 (N_424,In_562,In_1241);
xnor U425 (N_425,In_1703,In_1503);
and U426 (N_426,In_2227,In_1818);
nand U427 (N_427,In_2003,In_819);
or U428 (N_428,In_1347,In_437);
nand U429 (N_429,In_2410,In_21);
nand U430 (N_430,In_512,In_311);
or U431 (N_431,In_1089,In_1281);
nand U432 (N_432,In_1164,In_2185);
nand U433 (N_433,In_2094,In_272);
and U434 (N_434,In_1718,In_898);
and U435 (N_435,In_1804,In_847);
xor U436 (N_436,In_331,In_1796);
and U437 (N_437,In_1145,In_2201);
xnor U438 (N_438,In_2215,In_429);
nand U439 (N_439,In_1643,In_1512);
or U440 (N_440,In_768,In_2448);
and U441 (N_441,In_1924,In_242);
nor U442 (N_442,In_1518,In_1639);
and U443 (N_443,In_188,In_2309);
nand U444 (N_444,In_2445,In_1811);
and U445 (N_445,In_442,In_509);
xnor U446 (N_446,In_457,In_2369);
or U447 (N_447,In_1511,In_900);
or U448 (N_448,In_673,In_261);
and U449 (N_449,In_2142,In_1298);
xnor U450 (N_450,In_1458,In_421);
xor U451 (N_451,In_1585,In_2194);
xnor U452 (N_452,In_485,In_1756);
and U453 (N_453,In_379,In_674);
nor U454 (N_454,In_2198,In_2433);
nand U455 (N_455,In_564,In_450);
nor U456 (N_456,In_1122,In_415);
and U457 (N_457,In_1683,In_1500);
xnor U458 (N_458,In_1445,In_2261);
nand U459 (N_459,In_1036,In_2339);
nand U460 (N_460,In_2200,In_983);
xnor U461 (N_461,In_935,In_521);
nand U462 (N_462,In_1688,In_1364);
nand U463 (N_463,In_22,In_1257);
xor U464 (N_464,In_149,In_812);
and U465 (N_465,In_2335,In_1127);
xnor U466 (N_466,In_1489,In_2315);
xor U467 (N_467,In_1682,In_1169);
xor U468 (N_468,In_2083,In_1493);
or U469 (N_469,In_2026,In_1303);
nand U470 (N_470,In_163,In_1625);
and U471 (N_471,In_1680,In_1770);
xnor U472 (N_472,In_921,In_357);
nand U473 (N_473,In_70,In_2140);
and U474 (N_474,In_1366,In_816);
and U475 (N_475,In_153,In_1905);
nor U476 (N_476,In_1795,In_447);
and U477 (N_477,In_135,In_525);
xnor U478 (N_478,In_1872,In_2314);
nor U479 (N_479,In_2150,In_1037);
nand U480 (N_480,In_1473,In_940);
and U481 (N_481,In_1395,In_2177);
or U482 (N_482,In_1048,In_30);
or U483 (N_483,In_157,In_1868);
xor U484 (N_484,In_2109,In_528);
nor U485 (N_485,In_1728,In_402);
and U486 (N_486,In_1594,In_283);
nor U487 (N_487,In_365,In_2034);
and U488 (N_488,In_423,In_1457);
xor U489 (N_489,In_284,In_1313);
or U490 (N_490,In_811,In_2406);
nand U491 (N_491,In_636,In_1128);
nand U492 (N_492,In_1026,In_941);
or U493 (N_493,In_1253,In_1175);
nand U494 (N_494,In_666,In_1096);
nand U495 (N_495,In_511,In_1852);
xnor U496 (N_496,In_1507,In_2297);
or U497 (N_497,In_363,In_859);
xor U498 (N_498,In_1809,In_948);
or U499 (N_499,In_694,In_1427);
and U500 (N_500,In_1547,In_120);
or U501 (N_501,In_970,In_1732);
nor U502 (N_502,In_897,In_1030);
nor U503 (N_503,In_193,In_1925);
or U504 (N_504,In_804,In_1542);
or U505 (N_505,In_361,In_1747);
or U506 (N_506,In_1630,In_1017);
nor U507 (N_507,In_2388,In_2351);
nand U508 (N_508,In_1839,In_2291);
nand U509 (N_509,In_813,In_1361);
and U510 (N_510,In_1495,In_444);
and U511 (N_511,In_1114,In_2431);
nor U512 (N_512,In_1725,In_439);
or U513 (N_513,In_2019,In_152);
nor U514 (N_514,In_872,In_1702);
xnor U515 (N_515,In_865,In_286);
or U516 (N_516,In_175,In_1011);
nand U517 (N_517,In_641,In_448);
nand U518 (N_518,In_822,In_715);
xor U519 (N_519,In_866,In_1159);
and U520 (N_520,In_1223,In_1209);
xor U521 (N_521,In_1807,In_1560);
or U522 (N_522,In_2412,In_246);
and U523 (N_523,In_908,In_821);
xnor U524 (N_524,In_831,In_617);
nor U525 (N_525,In_1296,In_1300);
xnor U526 (N_526,In_2025,In_296);
and U527 (N_527,In_580,In_2474);
xor U528 (N_528,In_2051,In_1428);
or U529 (N_529,In_539,In_493);
xor U530 (N_530,In_1740,In_2328);
nand U531 (N_531,In_1686,In_391);
nor U532 (N_532,In_515,In_2462);
and U533 (N_533,In_1419,In_1015);
xor U534 (N_534,In_1050,In_372);
or U535 (N_535,In_1025,In_494);
nand U536 (N_536,In_2099,In_700);
or U537 (N_537,In_534,In_902);
and U538 (N_538,In_752,In_675);
and U539 (N_539,In_1237,In_668);
and U540 (N_540,In_527,In_191);
or U541 (N_541,In_974,In_522);
and U542 (N_542,In_37,In_122);
xnor U543 (N_543,In_281,In_2000);
nand U544 (N_544,In_2230,In_549);
nand U545 (N_545,In_1083,In_514);
nand U546 (N_546,In_1006,In_1731);
nor U547 (N_547,In_594,In_2287);
and U548 (N_548,In_112,In_392);
and U549 (N_549,In_2148,In_1836);
nand U550 (N_550,In_1072,In_150);
and U551 (N_551,In_524,In_1701);
or U552 (N_552,In_436,In_2074);
nor U553 (N_553,In_1100,In_1717);
nand U554 (N_554,In_8,In_1230);
xnor U555 (N_555,In_2300,In_911);
or U556 (N_556,In_502,In_2457);
or U557 (N_557,In_1068,In_2422);
xor U558 (N_558,In_2438,In_951);
nor U559 (N_559,In_1338,In_753);
nand U560 (N_560,In_2359,In_2391);
nand U561 (N_561,In_1180,In_316);
and U562 (N_562,In_1131,In_1362);
and U563 (N_563,In_1186,In_702);
nand U564 (N_564,In_173,In_1957);
or U565 (N_565,In_1488,In_344);
nor U566 (N_566,In_2452,In_628);
nor U567 (N_567,In_381,In_347);
xor U568 (N_568,In_2087,In_1062);
xor U569 (N_569,In_705,In_54);
or U570 (N_570,In_555,In_1962);
and U571 (N_571,In_1183,In_24);
or U572 (N_572,In_1359,In_1975);
xor U573 (N_573,In_573,In_119);
xor U574 (N_574,In_113,In_481);
and U575 (N_575,In_1142,In_1976);
nor U576 (N_576,In_1153,In_2450);
and U577 (N_577,In_2490,In_894);
nor U578 (N_578,In_25,In_1651);
and U579 (N_579,In_1221,In_786);
nand U580 (N_580,In_856,In_1875);
xnor U581 (N_581,In_2235,In_1301);
or U582 (N_582,In_245,In_170);
or U583 (N_583,In_291,In_1102);
nor U584 (N_584,In_1060,In_939);
and U585 (N_585,In_1671,In_1356);
or U586 (N_586,In_1007,In_2118);
and U587 (N_587,In_1204,In_751);
or U588 (N_588,In_2322,In_593);
nand U589 (N_589,In_2263,In_2143);
or U590 (N_590,In_757,In_917);
nor U591 (N_591,In_1412,In_1490);
nand U592 (N_592,In_1737,In_2243);
xor U593 (N_593,In_1085,In_1843);
or U594 (N_594,In_1855,In_2319);
or U595 (N_595,In_1655,In_577);
nor U596 (N_596,In_2389,In_2331);
or U597 (N_597,In_880,In_1636);
nand U598 (N_598,In_1283,In_1229);
or U599 (N_599,In_1236,In_2383);
and U600 (N_600,In_248,In_1430);
xnor U601 (N_601,In_1842,In_1126);
and U602 (N_602,In_1659,In_945);
or U603 (N_603,In_608,In_1403);
or U604 (N_604,In_2436,In_1927);
or U605 (N_605,In_794,In_1616);
xnor U606 (N_606,In_595,In_1946);
nand U607 (N_607,In_2193,In_797);
xor U608 (N_608,In_1288,In_765);
and U609 (N_609,In_721,In_1578);
and U610 (N_610,In_1392,In_1119);
nor U611 (N_611,In_1182,In_1799);
xnor U612 (N_612,In_1907,In_1084);
and U613 (N_613,In_572,In_1061);
nor U614 (N_614,In_929,In_2348);
or U615 (N_615,In_1456,In_568);
nor U616 (N_616,In_1173,In_1719);
xnor U617 (N_617,In_2280,In_2325);
nand U618 (N_618,In_1021,In_1949);
or U619 (N_619,In_633,In_966);
nand U620 (N_620,In_1637,In_2070);
nand U621 (N_621,In_1217,In_2347);
xor U622 (N_622,In_544,In_1692);
xnor U623 (N_623,In_1434,In_2301);
xor U624 (N_624,In_275,In_1463);
nand U625 (N_625,In_2014,In_419);
or U626 (N_626,In_1816,In_1140);
nand U627 (N_627,In_946,In_1150);
nand U628 (N_628,In_958,In_1207);
nor U629 (N_629,In_1020,In_2097);
nor U630 (N_630,In_1990,In_2470);
xnor U631 (N_631,In_1408,In_1261);
nor U632 (N_632,In_1442,In_258);
nor U633 (N_633,In_1076,In_1952);
xnor U634 (N_634,In_976,In_467);
xnor U635 (N_635,In_1444,In_339);
nor U636 (N_636,In_1562,In_2054);
xnor U637 (N_637,In_2258,In_58);
xnor U638 (N_638,In_116,In_368);
xor U639 (N_639,In_578,In_1736);
nand U640 (N_640,In_536,In_1589);
and U641 (N_641,In_996,In_234);
and U642 (N_642,In_1880,In_378);
or U643 (N_643,In_645,In_1774);
xnor U644 (N_644,In_1694,In_888);
or U645 (N_645,In_1504,In_2307);
nor U646 (N_646,In_890,In_1544);
and U647 (N_647,In_1961,In_2002);
xnor U648 (N_648,In_411,In_766);
nor U649 (N_649,In_2024,In_1928);
nand U650 (N_650,In_1660,In_1653);
and U651 (N_651,In_1691,In_588);
xor U652 (N_652,In_98,In_13);
nor U653 (N_653,In_1554,In_1522);
nand U654 (N_654,In_1613,In_273);
nor U655 (N_655,In_1550,In_125);
nand U656 (N_656,In_1837,In_2038);
nor U657 (N_657,In_997,In_1709);
or U658 (N_658,In_2417,In_73);
nand U659 (N_659,In_10,In_95);
xor U660 (N_660,In_740,In_2152);
xnor U661 (N_661,In_243,In_156);
xor U662 (N_662,In_1228,In_589);
nor U663 (N_663,In_430,In_1580);
nor U664 (N_664,In_686,In_499);
nand U665 (N_665,In_2495,In_408);
and U666 (N_666,In_180,In_400);
nand U667 (N_667,In_2260,In_584);
nand U668 (N_668,In_2131,In_2296);
nor U669 (N_669,In_2396,In_303);
nand U670 (N_670,In_838,In_1441);
nand U671 (N_671,In_1069,In_2384);
nor U672 (N_672,In_1826,In_1998);
and U673 (N_673,In_1154,In_1977);
nand U674 (N_674,In_586,In_1915);
nand U675 (N_675,In_1805,In_269);
nor U676 (N_676,In_1890,In_338);
nand U677 (N_677,In_554,In_2423);
and U678 (N_678,In_1596,In_336);
xnor U679 (N_679,In_147,In_398);
nand U680 (N_680,In_973,In_1117);
or U681 (N_681,In_1174,In_763);
xor U682 (N_682,In_1494,In_839);
xor U683 (N_683,In_854,In_416);
and U684 (N_684,In_2409,In_1987);
or U685 (N_685,In_569,In_2009);
and U686 (N_686,In_905,In_115);
and U687 (N_687,In_1201,In_1797);
nand U688 (N_688,In_791,In_1214);
nor U689 (N_689,In_1284,In_1307);
nand U690 (N_690,In_2077,In_2224);
nor U691 (N_691,In_1470,In_279);
nand U692 (N_692,In_19,In_1532);
and U693 (N_693,In_72,In_217);
nand U694 (N_694,In_1781,In_1792);
xnor U695 (N_695,In_2078,In_1243);
nor U696 (N_696,In_1714,In_693);
nor U697 (N_697,In_1191,In_477);
xor U698 (N_698,In_2356,In_858);
nand U699 (N_699,In_2210,In_1453);
nand U700 (N_700,In_79,In_2337);
or U701 (N_701,In_806,In_167);
and U702 (N_702,In_707,In_2228);
nor U703 (N_703,In_181,In_1646);
nand U704 (N_704,In_567,In_208);
and U705 (N_705,In_1206,In_2091);
xor U706 (N_706,In_2407,In_49);
nand U707 (N_707,In_2304,In_834);
or U708 (N_708,In_999,In_1120);
xnor U709 (N_709,In_1955,In_1867);
and U710 (N_710,In_724,In_124);
and U711 (N_711,In_650,In_207);
and U712 (N_712,In_2265,In_1658);
or U713 (N_713,In_1339,In_2132);
nand U714 (N_714,In_1152,In_1267);
xnor U715 (N_715,In_1746,In_1971);
and U716 (N_716,In_1825,In_1972);
nand U717 (N_717,In_2081,In_625);
or U718 (N_718,In_1615,In_510);
nand U719 (N_719,In_548,In_2472);
nand U720 (N_720,In_714,In_835);
or U721 (N_721,In_47,In_1019);
nor U722 (N_722,In_102,In_557);
xor U723 (N_723,In_798,In_472);
nand U724 (N_724,In_1092,In_1110);
xnor U725 (N_725,In_1628,In_861);
and U726 (N_726,In_2126,In_810);
or U727 (N_727,In_591,In_2165);
nor U728 (N_728,In_1916,In_1985);
and U729 (N_729,In_127,In_570);
and U730 (N_730,In_2144,In_1147);
nor U731 (N_731,In_1948,In_1383);
and U732 (N_732,In_2192,In_2375);
xnor U733 (N_733,In_455,In_746);
nor U734 (N_734,In_2021,In_1098);
nor U735 (N_735,In_912,In_1492);
xor U736 (N_736,In_274,In_784);
nor U737 (N_737,In_407,In_1815);
nor U738 (N_738,In_1687,In_1219);
xor U739 (N_739,In_1749,In_1652);
and U740 (N_740,In_1710,In_2181);
xor U741 (N_741,In_267,In_2202);
nand U742 (N_742,In_955,In_717);
and U743 (N_743,In_2478,In_2058);
nor U744 (N_744,In_937,In_614);
and U745 (N_745,In_209,In_1264);
and U746 (N_746,In_1561,In_654);
or U747 (N_747,In_667,In_907);
nor U748 (N_748,In_722,In_2098);
nand U749 (N_749,In_28,In_1794);
xor U750 (N_750,In_1597,In_1695);
xnor U751 (N_751,In_2342,In_1959);
xor U752 (N_752,In_579,In_215);
nor U753 (N_753,In_2028,In_927);
or U754 (N_754,In_863,In_1941);
xnor U755 (N_755,In_63,In_31);
xnor U756 (N_756,In_451,In_566);
or U757 (N_757,In_1078,In_2180);
nand U758 (N_758,In_703,In_293);
nor U759 (N_759,In_597,In_1258);
xor U760 (N_760,In_575,In_1932);
and U761 (N_761,In_1413,In_2485);
nand U762 (N_762,In_2475,In_1609);
nand U763 (N_763,In_309,In_961);
and U764 (N_764,In_683,In_1097);
and U765 (N_765,In_545,In_55);
nor U766 (N_766,In_432,In_2122);
xnor U767 (N_767,In_409,In_2404);
nand U768 (N_768,In_1409,In_2323);
nor U769 (N_769,In_298,In_2093);
and U770 (N_770,In_138,In_841);
and U771 (N_771,In_263,In_1936);
nor U772 (N_772,In_1136,In_1184);
nand U773 (N_773,In_96,In_2172);
and U774 (N_774,In_382,In_789);
and U775 (N_775,In_1133,In_799);
and U776 (N_776,In_2031,In_1640);
or U777 (N_777,In_1899,In_1082);
or U778 (N_778,In_770,In_1351);
nor U779 (N_779,In_334,In_733);
or U780 (N_780,In_851,In_1165);
and U781 (N_781,In_881,In_2129);
or U782 (N_782,In_1255,In_1973);
xnor U783 (N_783,In_1134,In_2418);
or U784 (N_784,In_1858,In_1606);
xnor U785 (N_785,In_1670,In_726);
and U786 (N_786,In_1431,In_1778);
nand U787 (N_787,In_2037,In_1081);
nor U788 (N_788,In_484,In_2350);
and U789 (N_789,In_148,In_1227);
or U790 (N_790,In_843,In_1041);
or U791 (N_791,In_1713,In_2187);
nand U792 (N_792,In_2141,In_304);
nand U793 (N_793,In_631,In_2363);
nand U794 (N_794,In_489,In_1771);
or U795 (N_795,In_957,In_1446);
nor U796 (N_796,In_1459,In_1166);
or U797 (N_797,In_356,In_118);
xor U798 (N_798,In_1903,In_1635);
nand U799 (N_799,In_873,In_1137);
or U800 (N_800,In_2050,In_471);
nand U801 (N_801,In_899,In_785);
nor U802 (N_802,In_1115,In_216);
xor U803 (N_803,In_767,In_2421);
and U804 (N_804,In_563,In_2121);
xor U805 (N_805,In_1527,In_2246);
nor U806 (N_806,In_871,In_1333);
and U807 (N_807,In_1218,In_2441);
and U808 (N_808,In_1930,In_969);
nand U809 (N_809,In_229,In_1641);
nor U810 (N_810,In_2124,In_661);
nor U811 (N_811,In_2386,In_2175);
xnor U812 (N_812,In_1480,In_1208);
nand U813 (N_813,In_696,In_1203);
nand U814 (N_814,In_1889,In_117);
xor U815 (N_815,In_1256,In_2173);
nor U816 (N_816,In_254,In_1330);
xnor U817 (N_817,In_1171,In_1546);
or U818 (N_818,In_1833,In_26);
nand U819 (N_819,In_418,In_620);
nand U820 (N_820,In_781,In_2259);
xnor U821 (N_821,In_1160,In_553);
nand U822 (N_822,In_1534,In_1107);
and U823 (N_823,In_132,In_340);
and U824 (N_824,In_830,In_2318);
and U825 (N_825,In_227,In_1162);
nand U826 (N_826,In_590,In_1116);
or U827 (N_827,In_607,In_2321);
xnor U828 (N_828,In_1840,In_2275);
and U829 (N_829,In_1886,In_815);
and U830 (N_830,In_725,In_2158);
nor U831 (N_831,In_1421,In_2295);
xnor U832 (N_832,In_2079,In_341);
and U833 (N_833,In_613,In_2017);
and U834 (N_834,In_1787,In_1896);
and U835 (N_835,In_2186,In_1497);
nor U836 (N_836,In_462,In_2376);
or U837 (N_837,In_321,In_204);
or U838 (N_838,In_17,In_100);
xor U839 (N_839,In_1429,In_571);
or U840 (N_840,In_1993,In_1620);
xor U841 (N_841,In_35,In_507);
nand U842 (N_842,In_2040,In_84);
xor U843 (N_843,In_1271,In_1013);
xnor U844 (N_844,In_2204,In_1067);
nand U845 (N_845,In_2357,In_2080);
nor U846 (N_846,In_1822,In_1437);
or U847 (N_847,In_1631,In_1664);
nor U848 (N_848,In_2371,In_1121);
and U849 (N_849,In_1135,In_1901);
and U850 (N_850,In_2044,In_1989);
nor U851 (N_851,In_1234,In_1869);
nand U852 (N_852,In_290,In_51);
or U853 (N_853,In_355,In_832);
nand U854 (N_854,In_369,In_143);
nor U855 (N_855,In_1332,In_94);
or U856 (N_856,In_45,In_1059);
nor U857 (N_857,In_611,In_1394);
nand U858 (N_858,In_389,In_233);
or U859 (N_859,In_857,In_1559);
nor U860 (N_860,In_906,In_2411);
nor U861 (N_861,In_670,In_1553);
nor U862 (N_862,In_809,In_655);
xor U863 (N_863,In_1848,In_1224);
xor U864 (N_864,In_1780,In_1095);
or U865 (N_865,In_1621,In_2249);
nand U866 (N_866,In_2035,In_2084);
or U867 (N_867,In_1540,In_198);
and U868 (N_868,In_1530,In_630);
xor U869 (N_869,In_887,In_639);
nor U870 (N_870,In_386,In_895);
and U871 (N_871,In_849,In_904);
or U872 (N_872,In_1337,In_1297);
and U873 (N_873,In_1282,In_1919);
or U874 (N_874,In_754,In_777);
and U875 (N_875,In_1940,In_943);
nor U876 (N_876,In_1752,In_2011);
xor U877 (N_877,In_1317,In_29);
nand U878 (N_878,In_249,In_352);
or U879 (N_879,In_2179,In_2195);
nor U880 (N_880,In_2155,In_640);
or U881 (N_881,In_2191,In_1675);
and U882 (N_882,In_807,In_1793);
and U883 (N_883,In_1038,In_876);
or U884 (N_884,In_2220,In_2252);
xnor U885 (N_885,In_387,In_2096);
nor U886 (N_886,In_1308,In_277);
xor U887 (N_887,In_164,In_909);
or U888 (N_888,In_1058,In_2329);
nor U889 (N_889,In_2355,In_1754);
nor U890 (N_890,In_1319,In_1963);
xor U891 (N_891,In_1885,In_160);
nor U892 (N_892,In_1101,In_878);
and U893 (N_893,In_1225,In_441);
nand U894 (N_894,In_260,In_1950);
xnor U895 (N_895,In_1113,In_1878);
or U896 (N_896,In_329,In_884);
nor U897 (N_897,In_1369,In_1393);
xnor U898 (N_898,In_2270,In_1358);
nand U899 (N_899,In_2029,In_2419);
xnor U900 (N_900,In_2282,In_1873);
xnor U901 (N_901,In_592,In_1934);
xor U902 (N_902,In_252,In_964);
nand U903 (N_903,In_1730,In_1367);
nor U904 (N_904,In_1956,In_1715);
nand U905 (N_905,In_718,In_642);
or U906 (N_906,In_684,In_1143);
nand U907 (N_907,In_2136,In_1851);
xnor U908 (N_908,In_1900,In_300);
or U909 (N_909,In_1566,In_2443);
or U910 (N_910,In_840,In_2269);
and U911 (N_911,In_1824,In_1464);
xnor U912 (N_912,In_2164,In_2401);
or U913 (N_913,In_1524,In_1200);
nand U914 (N_914,In_75,In_844);
nand U915 (N_915,In_1046,In_294);
nor U916 (N_916,In_1327,In_1077);
or U917 (N_917,In_326,In_2248);
nand U918 (N_918,In_992,In_1593);
xor U919 (N_919,In_914,In_2166);
nand U920 (N_920,In_2145,In_2039);
nor U921 (N_921,In_83,In_384);
or U922 (N_922,In_2189,In_2435);
nand U923 (N_923,In_2469,In_1416);
nor U924 (N_924,In_1075,In_933);
nand U925 (N_925,In_1520,In_413);
nor U926 (N_926,In_1250,In_2455);
xnor U927 (N_927,In_2052,In_1802);
and U928 (N_928,In_731,In_1396);
xor U929 (N_929,In_1465,In_2468);
and U930 (N_930,In_1720,In_1426);
and U931 (N_931,In_986,In_244);
or U932 (N_932,In_1996,In_11);
and U933 (N_933,In_994,In_2216);
or U934 (N_934,In_1414,In_1244);
xnor U935 (N_935,In_223,In_773);
nor U936 (N_936,In_713,In_1716);
nand U937 (N_937,In_1681,In_139);
nor U938 (N_938,In_814,In_78);
or U939 (N_939,In_1803,In_915);
xor U940 (N_940,In_1189,In_2268);
nor U941 (N_941,In_990,In_842);
nand U942 (N_942,In_1525,In_622);
xnor U943 (N_943,In_225,In_761);
and U944 (N_944,In_652,In_1912);
nand U945 (N_945,In_405,In_1539);
or U946 (N_946,In_232,In_1387);
nand U947 (N_947,In_1354,In_1861);
and U948 (N_948,In_1967,In_1579);
xnor U949 (N_949,In_1991,In_2160);
or U950 (N_950,In_1914,In_1938);
nor U951 (N_951,In_1193,In_222);
and U952 (N_952,In_2225,In_1791);
or U953 (N_953,In_89,In_224);
nand U954 (N_954,In_977,In_1328);
nand U955 (N_955,In_728,In_1782);
nor U956 (N_956,In_1044,In_954);
xnor U957 (N_957,In_2167,In_470);
nand U958 (N_958,In_561,In_2463);
and U959 (N_959,In_760,In_2171);
or U960 (N_960,In_1141,In_802);
and U961 (N_961,In_324,In_1476);
nand U962 (N_962,In_698,In_1499);
nand U963 (N_963,In_869,In_1661);
nand U964 (N_964,In_2480,In_1034);
nor U965 (N_965,In_2428,In_2211);
nor U966 (N_966,In_420,In_1887);
nor U967 (N_967,In_855,In_1451);
or U968 (N_968,In_2451,In_526);
xor U969 (N_969,In_2041,In_2207);
xor U970 (N_970,In_1984,In_2247);
nand U971 (N_971,In_33,In_829);
or U972 (N_972,In_2402,In_362);
or U973 (N_973,In_1622,In_609);
nand U974 (N_974,In_2015,In_2303);
nor U975 (N_975,In_1923,In_2008);
nand U976 (N_976,In_66,In_108);
xnor U977 (N_977,In_2338,In_46);
nor U978 (N_978,In_1706,In_936);
and U979 (N_979,In_1817,In_1001);
or U980 (N_980,In_129,In_530);
xnor U981 (N_981,In_1018,In_503);
xnor U982 (N_982,In_142,In_1401);
xor U983 (N_983,In_1552,In_967);
and U984 (N_984,In_1810,In_644);
or U985 (N_985,In_265,In_469);
nor U986 (N_986,In_1697,In_1231);
nor U987 (N_987,In_1679,In_2430);
and U988 (N_988,In_2279,In_2089);
nor U989 (N_989,In_276,In_2102);
or U990 (N_990,In_1557,In_529);
xor U991 (N_991,In_314,In_2368);
and U992 (N_992,In_424,In_213);
or U993 (N_993,In_241,In_266);
nor U994 (N_994,In_924,In_318);
xnor U995 (N_995,In_2397,In_1291);
xnor U996 (N_996,In_87,In_1391);
xnor U997 (N_997,In_1881,In_1929);
xnor U998 (N_998,In_2219,In_2360);
and U999 (N_999,In_1326,In_348);
nand U1000 (N_1000,N_366,N_749);
nor U1001 (N_1001,N_27,N_961);
nor U1002 (N_1002,N_537,N_80);
and U1003 (N_1003,N_29,N_535);
or U1004 (N_1004,N_626,In_2053);
nand U1005 (N_1005,N_41,N_980);
nor U1006 (N_1006,N_553,N_243);
xor U1007 (N_1007,In_270,N_276);
xor U1008 (N_1008,N_70,N_113);
or U1009 (N_1009,N_963,N_94);
or U1010 (N_1010,N_824,In_2);
or U1011 (N_1011,N_98,N_772);
xnor U1012 (N_1012,N_723,N_154);
or U1013 (N_1013,N_385,N_750);
or U1014 (N_1014,N_652,In_177);
and U1015 (N_1015,N_566,N_169);
and U1016 (N_1016,N_454,N_251);
nor U1017 (N_1017,N_704,N_559);
and U1018 (N_1018,N_856,N_229);
nor U1019 (N_1019,N_640,N_509);
nand U1020 (N_1020,N_710,In_1678);
nand U1021 (N_1021,In_1965,N_861);
nand U1022 (N_1022,N_12,N_711);
or U1023 (N_1023,N_122,N_754);
xnor U1024 (N_1024,N_307,N_193);
and U1025 (N_1025,N_205,In_288);
and U1026 (N_1026,N_787,N_436);
nor U1027 (N_1027,N_521,In_664);
and U1028 (N_1028,N_811,In_956);
xnor U1029 (N_1029,In_2343,N_77);
nor U1030 (N_1030,N_594,In_401);
and U1031 (N_1031,N_302,In_1521);
or U1032 (N_1032,N_679,N_547);
xor U1033 (N_1033,In_1318,N_548);
xnor U1034 (N_1034,N_792,In_2048);
or U1035 (N_1035,N_355,N_442);
or U1036 (N_1036,N_47,N_808);
nor U1037 (N_1037,N_266,N_242);
or U1038 (N_1038,In_1439,In_2381);
or U1039 (N_1039,N_650,In_730);
nand U1040 (N_1040,N_245,N_427);
xnor U1041 (N_1041,N_874,In_1325);
xor U1042 (N_1042,In_2429,In_162);
xor U1043 (N_1043,In_2163,N_877);
and U1044 (N_1044,N_727,In_1565);
or U1045 (N_1045,In_1260,N_317);
or U1046 (N_1046,N_136,N_76);
nor U1047 (N_1047,N_666,N_10);
nor U1048 (N_1048,N_83,N_479);
or U1049 (N_1049,N_492,N_876);
xnor U1050 (N_1050,N_948,In_1764);
and U1051 (N_1051,N_982,In_1931);
nand U1052 (N_1052,N_13,N_511);
and U1053 (N_1053,N_206,N_507);
xnor U1054 (N_1054,N_775,N_354);
xnor U1055 (N_1055,N_289,N_917);
xor U1056 (N_1056,N_984,In_2147);
xnor U1057 (N_1057,N_998,In_1992);
nand U1058 (N_1058,N_313,N_740);
xor U1059 (N_1059,In_2349,N_432);
or U1060 (N_1060,N_519,In_2398);
or U1061 (N_1061,N_167,N_579);
and U1062 (N_1062,N_560,N_437);
xor U1063 (N_1063,In_1979,N_873);
nand U1064 (N_1064,In_919,N_6);
nand U1065 (N_1065,N_709,N_486);
and U1066 (N_1066,N_830,N_1);
nand U1067 (N_1067,N_138,N_497);
nor U1068 (N_1068,N_204,N_938);
nand U1069 (N_1069,N_935,In_800);
nor U1070 (N_1070,In_2206,N_693);
nand U1071 (N_1071,N_272,N_870);
nand U1072 (N_1072,N_194,In_1376);
xor U1073 (N_1073,In_1757,N_778);
and U1074 (N_1074,N_880,N_678);
nand U1075 (N_1075,In_627,N_867);
and U1076 (N_1076,In_649,N_940);
nor U1077 (N_1077,N_165,N_149);
xnor U1078 (N_1078,N_600,N_34);
nand U1079 (N_1079,N_121,N_415);
nand U1080 (N_1080,N_869,N_786);
and U1081 (N_1081,N_155,In_1969);
nor U1082 (N_1082,N_717,N_196);
or U1083 (N_1083,N_120,In_1605);
nand U1084 (N_1084,N_326,N_655);
nor U1085 (N_1085,N_765,In_699);
or U1086 (N_1086,N_36,N_890);
nor U1087 (N_1087,N_224,N_662);
nor U1088 (N_1088,In_1293,N_841);
or U1089 (N_1089,N_103,N_612);
nor U1090 (N_1090,N_417,N_425);
nand U1091 (N_1091,N_258,N_45);
nor U1092 (N_1092,In_1146,N_728);
and U1093 (N_1093,In_706,N_915);
nand U1094 (N_1094,N_993,In_801);
and U1095 (N_1095,In_1599,N_449);
and U1096 (N_1096,N_905,N_541);
and U1097 (N_1097,N_857,N_803);
and U1098 (N_1098,N_32,N_677);
xnor U1099 (N_1099,N_340,N_247);
xnor U1100 (N_1100,In_1065,N_868);
xor U1101 (N_1101,In_2184,N_598);
nand U1102 (N_1102,N_974,N_275);
xor U1103 (N_1103,N_127,N_304);
nand U1104 (N_1104,N_766,N_249);
nand U1105 (N_1105,In_189,N_350);
nor U1106 (N_1106,In_1188,N_588);
xnor U1107 (N_1107,N_763,N_410);
and U1108 (N_1108,N_871,In_1384);
nor U1109 (N_1109,In_2116,N_48);
and U1110 (N_1110,In_1158,N_996);
or U1111 (N_1111,In_1280,N_450);
nand U1112 (N_1112,N_911,In_2292);
or U1113 (N_1113,N_327,In_71);
or U1114 (N_1114,In_128,In_1704);
and U1115 (N_1115,In_1871,N_746);
or U1116 (N_1116,N_733,N_922);
xor U1117 (N_1117,In_16,In_1980);
xnor U1118 (N_1118,N_458,N_226);
xor U1119 (N_1119,In_417,N_587);
or U1120 (N_1120,N_90,In_1031);
nor U1121 (N_1121,In_366,N_150);
nor U1122 (N_1122,N_471,N_718);
nand U1123 (N_1123,In_779,In_749);
nor U1124 (N_1124,In_2479,N_744);
nand U1125 (N_1125,In_1884,In_228);
xnor U1126 (N_1126,In_860,N_960);
nor U1127 (N_1127,N_375,In_1591);
xnor U1128 (N_1128,N_531,N_826);
nor U1129 (N_1129,In_2442,N_633);
and U1130 (N_1130,N_369,In_2395);
or U1131 (N_1131,N_109,N_310);
nand U1132 (N_1132,N_930,N_253);
xnor U1133 (N_1133,In_1910,In_2151);
nand U1134 (N_1134,N_296,In_1763);
nor U1135 (N_1135,N_696,N_398);
and U1136 (N_1136,N_360,In_1541);
nor U1137 (N_1137,N_517,N_762);
xor U1138 (N_1138,In_1487,In_2370);
nor U1139 (N_1139,In_2226,In_2105);
or U1140 (N_1140,In_2061,N_164);
and U1141 (N_1141,In_734,N_74);
nand U1142 (N_1142,N_664,In_2046);
nor U1143 (N_1143,N_828,In_1537);
or U1144 (N_1144,N_406,N_295);
and U1145 (N_1145,N_312,N_311);
or U1146 (N_1146,In_2373,N_706);
and U1147 (N_1147,N_502,N_314);
nor U1148 (N_1148,In_487,N_146);
nand U1149 (N_1149,In_2072,N_260);
and U1150 (N_1150,N_965,N_783);
xor U1151 (N_1151,N_75,In_531);
nor U1152 (N_1152,N_599,In_2133);
xor U1153 (N_1153,N_409,N_148);
nand U1154 (N_1154,In_1812,In_2092);
or U1155 (N_1155,In_1607,N_571);
and U1156 (N_1156,N_3,N_390);
xor U1157 (N_1157,In_2336,In_710);
and U1158 (N_1158,N_373,In_903);
and U1159 (N_1159,N_757,N_234);
nor U1160 (N_1160,N_86,In_1425);
nand U1161 (N_1161,In_769,N_331);
or U1162 (N_1162,N_202,N_575);
xor U1163 (N_1163,N_608,In_2362);
and U1164 (N_1164,N_708,In_891);
or U1165 (N_1165,N_144,N_837);
nand U1166 (N_1166,N_423,In_612);
xnor U1167 (N_1167,N_23,N_73);
xor U1168 (N_1168,N_823,In_1418);
nor U1169 (N_1169,N_203,In_926);
and U1170 (N_1170,N_208,N_741);
xnor U1171 (N_1171,N_512,N_816);
or U1172 (N_1172,In_1498,N_593);
xnor U1173 (N_1173,In_660,N_207);
or U1174 (N_1174,N_418,N_564);
or U1175 (N_1175,N_651,N_790);
nor U1176 (N_1176,In_221,N_49);
and U1177 (N_1177,N_761,N_707);
nand U1178 (N_1178,In_292,N_605);
and U1179 (N_1179,N_128,N_470);
or U1180 (N_1180,N_473,N_399);
nor U1181 (N_1181,N_428,N_35);
xnor U1182 (N_1182,N_15,N_294);
and U1183 (N_1183,In_1108,N_884);
or U1184 (N_1184,N_189,N_163);
and U1185 (N_1185,N_25,N_446);
and U1186 (N_1186,N_43,N_301);
or U1187 (N_1187,N_33,N_380);
xor U1188 (N_1188,N_606,In_1039);
and U1189 (N_1189,In_1834,N_453);
nand U1190 (N_1190,N_274,In_995);
xnor U1191 (N_1191,N_26,N_157);
or U1192 (N_1192,In_67,N_545);
nor U1193 (N_1193,N_456,N_279);
and U1194 (N_1194,N_957,N_526);
xnor U1195 (N_1195,N_420,In_103);
or U1196 (N_1196,In_218,N_215);
and U1197 (N_1197,In_1066,In_583);
nor U1198 (N_1198,In_1386,In_2139);
xnor U1199 (N_1199,N_508,N_506);
or U1200 (N_1200,N_720,In_454);
xnor U1201 (N_1201,N_618,N_851);
xnor U1202 (N_1202,N_269,N_63);
nor U1203 (N_1203,N_768,N_457);
nand U1204 (N_1204,N_889,N_953);
or U1205 (N_1205,N_668,N_695);
or U1206 (N_1206,N_863,N_2);
nand U1207 (N_1207,In_1370,In_2271);
xor U1208 (N_1208,In_1820,N_567);
xor U1209 (N_1209,N_110,N_694);
xnor U1210 (N_1210,N_186,N_178);
or U1211 (N_1211,In_708,N_287);
nand U1212 (N_1212,N_478,N_183);
xnor U1213 (N_1213,In_327,In_1835);
xnor U1214 (N_1214,N_382,N_795);
xnor U1215 (N_1215,N_151,In_2256);
and U1216 (N_1216,N_161,In_305);
or U1217 (N_1217,N_764,N_734);
nand U1218 (N_1218,In_1496,N_132);
or U1219 (N_1219,N_44,N_18);
nor U1220 (N_1220,N_576,N_839);
and U1221 (N_1221,In_793,N_732);
xor U1222 (N_1222,In_1029,N_627);
or U1223 (N_1223,N_461,N_5);
nor U1224 (N_1224,In_1138,N_177);
xor U1225 (N_1225,N_939,In_488);
or U1226 (N_1226,N_438,In_968);
and U1227 (N_1227,N_529,N_614);
nand U1228 (N_1228,N_218,N_495);
xor U1229 (N_1229,N_941,N_337);
nand U1230 (N_1230,N_983,N_909);
and U1231 (N_1231,N_849,In_808);
nand U1232 (N_1232,N_14,In_1935);
or U1233 (N_1233,N_752,In_2232);
nand U1234 (N_1234,N_28,N_219);
and U1235 (N_1235,In_2090,N_268);
xnor U1236 (N_1236,N_546,In_1877);
and U1237 (N_1237,N_67,N_630);
xnor U1238 (N_1238,In_610,N_555);
nor U1239 (N_1239,N_702,N_628);
xnor U1240 (N_1240,In_2276,N_966);
nor U1241 (N_1241,In_1151,N_166);
xor U1242 (N_1242,In_1846,N_568);
nand U1243 (N_1243,In_1398,In_805);
and U1244 (N_1244,N_291,N_407);
xor U1245 (N_1245,N_820,N_852);
nor U1246 (N_1246,N_888,N_345);
and U1247 (N_1247,In_183,N_435);
or U1248 (N_1248,N_241,In_1192);
nand U1249 (N_1249,In_82,N_788);
and U1250 (N_1250,N_179,In_1551);
or U1251 (N_1251,N_59,In_1056);
xor U1252 (N_1252,In_2231,In_818);
xor U1253 (N_1253,N_482,In_271);
or U1254 (N_1254,N_447,N_898);
nand U1255 (N_1255,In_1624,In_2456);
nand U1256 (N_1256,N_819,N_916);
and U1257 (N_1257,N_745,N_434);
or U1258 (N_1258,N_501,N_534);
nor U1259 (N_1259,N_848,In_500);
nand U1260 (N_1260,N_60,In_2082);
xnor U1261 (N_1261,N_596,N_714);
or U1262 (N_1262,N_332,In_989);
or U1263 (N_1263,N_156,In_1304);
xnor U1264 (N_1264,N_780,N_37);
nand U1265 (N_1265,In_1450,N_945);
or U1266 (N_1266,N_946,N_907);
xor U1267 (N_1267,N_283,In_2378);
nor U1268 (N_1268,In_1742,In_2367);
xnor U1269 (N_1269,N_971,In_1501);
nor U1270 (N_1270,N_221,In_1144);
nor U1271 (N_1271,N_958,N_514);
xor U1272 (N_1272,N_844,In_2427);
and U1273 (N_1273,N_691,N_141);
nor U1274 (N_1274,N_469,In_1063);
nand U1275 (N_1275,In_1053,N_46);
xnor U1276 (N_1276,N_855,N_227);
or U1277 (N_1277,N_680,In_403);
or U1278 (N_1278,In_136,N_364);
nand U1279 (N_1279,In_1436,In_1649);
nand U1280 (N_1280,N_956,N_902);
nand U1281 (N_1281,In_1397,In_1603);
xor U1282 (N_1282,In_1970,N_979);
xor U1283 (N_1283,N_441,N_271);
or U1284 (N_1284,In_520,N_235);
xnor U1285 (N_1285,N_969,N_671);
xor U1286 (N_1286,N_928,N_604);
nor U1287 (N_1287,N_338,In_2332);
xnor U1288 (N_1288,N_64,In_1210);
nand U1289 (N_1289,N_753,N_411);
xnor U1290 (N_1290,N_927,N_716);
xor U1291 (N_1291,N_254,In_426);
or U1292 (N_1292,N_321,N_270);
or U1293 (N_1293,N_368,In_463);
nor U1294 (N_1294,N_220,In_255);
and U1295 (N_1295,N_700,N_82);
or U1296 (N_1296,N_949,N_987);
nor U1297 (N_1297,N_527,N_51);
nor U1298 (N_1298,N_475,In_833);
xnor U1299 (N_1299,N_383,N_817);
and U1300 (N_1300,N_107,N_284);
nand U1301 (N_1301,N_617,N_439);
and U1302 (N_1302,N_638,N_16);
nor U1303 (N_1303,N_543,In_1592);
xnor U1304 (N_1304,N_601,N_954);
nor U1305 (N_1305,N_288,N_991);
nand U1306 (N_1306,N_17,N_522);
and U1307 (N_1307,In_62,In_1302);
xor U1308 (N_1308,N_463,N_257);
or U1309 (N_1309,N_65,N_391);
nand U1310 (N_1310,In_1474,N_342);
xnor U1311 (N_1311,N_675,N_324);
and U1312 (N_1312,In_1821,In_43);
and U1313 (N_1313,N_228,N_562);
xor U1314 (N_1314,N_858,In_1087);
nand U1315 (N_1315,N_920,In_2119);
nand U1316 (N_1316,N_670,In_2326);
or U1317 (N_1317,N_607,N_467);
and U1318 (N_1318,N_92,N_866);
and U1319 (N_1319,N_850,N_168);
and U1320 (N_1320,N_20,In_323);
nor U1321 (N_1321,N_431,N_656);
or U1322 (N_1322,N_145,N_0);
and U1323 (N_1323,N_238,N_395);
nor U1324 (N_1324,N_815,N_133);
nand U1325 (N_1325,N_616,N_703);
nor U1326 (N_1326,N_119,In_231);
or U1327 (N_1327,In_701,N_947);
and U1328 (N_1328,N_644,N_101);
nor U1329 (N_1329,N_147,In_988);
nand U1330 (N_1330,N_376,N_936);
nor U1331 (N_1331,N_343,N_333);
nand U1332 (N_1332,In_1632,N_569);
and U1333 (N_1333,N_756,In_1665);
xor U1334 (N_1334,In_626,In_735);
and U1335 (N_1335,N_267,N_912);
and U1336 (N_1336,In_1693,N_676);
and U1337 (N_1337,In_1388,N_216);
nand U1338 (N_1338,N_899,N_794);
xor U1339 (N_1339,N_209,N_225);
nand U1340 (N_1340,N_505,In_126);
nand U1341 (N_1341,N_451,In_2477);
and U1342 (N_1342,N_900,N_827);
nand U1343 (N_1343,In_81,In_1009);
nor U1344 (N_1344,N_481,In_535);
nand U1345 (N_1345,In_1322,N_838);
and U1346 (N_1346,N_440,N_213);
and U1347 (N_1347,In_1483,N_933);
nor U1348 (N_1348,N_636,N_951);
nor U1349 (N_1349,In_1099,N_22);
or U1350 (N_1350,In_868,In_301);
and U1351 (N_1351,N_865,In_1570);
nor U1352 (N_1352,In_875,In_1892);
or U1353 (N_1353,N_747,N_712);
nor U1354 (N_1354,N_658,N_152);
and U1355 (N_1355,N_31,In_1310);
nand U1356 (N_1356,In_165,N_8);
nor U1357 (N_1357,N_879,In_680);
or U1358 (N_1358,N_344,In_2149);
xor U1359 (N_1359,N_480,N_445);
nand U1360 (N_1360,N_386,N_277);
nand U1361 (N_1361,N_172,N_525);
and U1362 (N_1362,N_800,N_544);
nand U1363 (N_1363,In_259,N_443);
nand U1364 (N_1364,N_860,N_494);
nand U1365 (N_1365,N_755,N_619);
nor U1366 (N_1366,N_893,In_2156);
xor U1367 (N_1367,In_538,N_730);
and U1368 (N_1368,N_796,In_574);
xnor U1369 (N_1369,In_1123,In_1342);
nand U1370 (N_1370,In_1054,In_2138);
nand U1371 (N_1371,In_1908,N_847);
nor U1372 (N_1372,In_756,N_955);
nand U1373 (N_1373,In_516,N_959);
and U1374 (N_1374,N_118,N_129);
or U1375 (N_1375,In_1708,N_906);
nand U1376 (N_1376,In_159,N_182);
and U1377 (N_1377,N_484,N_833);
nand U1378 (N_1378,N_743,N_188);
nor U1379 (N_1379,N_914,N_532);
xor U1380 (N_1380,In_2424,N_685);
or U1381 (N_1381,N_643,N_985);
and U1382 (N_1382,In_1435,N_782);
and U1383 (N_1383,In_2365,N_715);
or U1384 (N_1384,N_97,N_705);
and U1385 (N_1385,In_1148,N_503);
nor U1386 (N_1386,In_2188,N_625);
nand U1387 (N_1387,N_214,N_358);
and U1388 (N_1388,N_822,N_190);
nand U1389 (N_1389,N_319,N_595);
and U1390 (N_1390,In_1238,In_2283);
nand U1391 (N_1391,In_938,In_2127);
xor U1392 (N_1392,N_185,N_318);
nor U1393 (N_1393,In_199,N_924);
nor U1394 (N_1394,N_690,In_762);
nor U1395 (N_1395,In_238,In_2346);
xnor U1396 (N_1396,N_498,In_1371);
xnor U1397 (N_1397,N_329,In_1389);
nand U1398 (N_1398,In_2253,In_1278);
nand U1399 (N_1399,N_773,N_973);
nor U1400 (N_1400,In_64,N_160);
xnor U1401 (N_1401,N_986,N_736);
nand U1402 (N_1402,In_2439,N_646);
nor U1403 (N_1403,N_309,In_1762);
and U1404 (N_1404,N_389,N_779);
or U1405 (N_1405,N_923,In_250);
or U1406 (N_1406,N_388,N_171);
nand U1407 (N_1407,In_2333,N_353);
and U1408 (N_1408,N_404,N_950);
nand U1409 (N_1409,N_729,N_341);
nor U1410 (N_1410,In_1689,N_197);
or U1411 (N_1411,N_66,N_444);
nand U1412 (N_1412,N_465,N_552);
and U1413 (N_1413,N_845,In_1197);
nor U1414 (N_1414,N_175,N_57);
nor U1415 (N_1415,N_367,N_490);
nor U1416 (N_1416,N_981,N_499);
nand U1417 (N_1417,In_1572,N_299);
xnor U1418 (N_1418,N_894,In_41);
xnor U1419 (N_1419,N_162,N_95);
nor U1420 (N_1420,In_1215,In_828);
nand U1421 (N_1421,N_223,In_371);
nand U1422 (N_1422,In_92,In_2312);
nand U1423 (N_1423,N_102,N_233);
nor U1424 (N_1424,N_530,In_1035);
xor U1425 (N_1425,N_89,N_806);
nand U1426 (N_1426,N_114,In_1922);
nand U1427 (N_1427,In_1856,In_1277);
and U1428 (N_1428,In_540,N_58);
nand U1429 (N_1429,N_854,N_661);
nand U1430 (N_1430,In_1477,In_133);
xor U1431 (N_1431,N_230,In_1510);
or U1432 (N_1432,N_131,N_212);
nor U1433 (N_1433,N_903,N_797);
xor U1434 (N_1434,N_290,In_2059);
xnor U1435 (N_1435,In_523,N_262);
and U1436 (N_1436,In_2095,N_524);
or U1437 (N_1437,N_19,N_292);
nand U1438 (N_1438,In_2449,In_1057);
and U1439 (N_1439,N_846,N_777);
nand U1440 (N_1440,N_789,In_1904);
or U1441 (N_1441,N_843,N_416);
xnor U1442 (N_1442,In_61,N_256);
nand U1443 (N_1443,N_572,N_721);
or U1444 (N_1444,N_580,N_24);
nor U1445 (N_1445,N_615,N_809);
xor U1446 (N_1446,N_306,In_1417);
xnor U1447 (N_1447,In_1273,N_85);
nand U1448 (N_1448,N_335,N_265);
xor U1449 (N_1449,In_27,In_1028);
or U1450 (N_1450,N_105,In_1662);
nand U1451 (N_1451,In_1529,N_738);
xor U1452 (N_1452,N_859,N_760);
xor U1453 (N_1453,In_2113,N_645);
nor U1454 (N_1454,N_71,N_831);
or U1455 (N_1455,In_2399,N_518);
nor U1456 (N_1456,N_187,N_584);
or U1457 (N_1457,N_539,N_834);
nor U1458 (N_1458,N_813,N_170);
nor U1459 (N_1459,N_378,In_1673);
nor U1460 (N_1460,N_278,In_2062);
xor U1461 (N_1461,N_42,N_591);
nand U1462 (N_1462,In_476,In_2374);
and U1463 (N_1463,N_139,In_1601);
and U1464 (N_1464,N_937,In_962);
and U1465 (N_1465,N_400,N_972);
xnor U1466 (N_1466,N_7,N_356);
xor U1467 (N_1467,N_943,In_1475);
and U1468 (N_1468,N_913,In_1070);
or U1469 (N_1469,N_829,In_893);
and U1470 (N_1470,N_426,N_520);
nand U1471 (N_1471,N_143,N_682);
nor U1472 (N_1472,N_142,N_774);
xnor U1473 (N_1473,N_408,N_261);
nand U1474 (N_1474,N_647,In_172);
nor U1475 (N_1475,N_130,N_952);
nand U1476 (N_1476,In_2110,N_466);
xor U1477 (N_1477,N_513,N_597);
nor U1478 (N_1478,N_840,N_252);
nor U1479 (N_1479,N_123,In_980);
nor U1480 (N_1480,N_336,In_1249);
and U1481 (N_1481,N_975,N_54);
and U1482 (N_1482,N_55,In_1289);
xor U1483 (N_1483,In_349,N_237);
nand U1484 (N_1484,In_308,N_394);
xnor U1485 (N_1485,In_393,N_759);
xnor U1486 (N_1486,N_583,N_392);
xor U1487 (N_1487,N_106,N_832);
nand U1488 (N_1488,In_2481,In_202);
or U1489 (N_1489,N_72,N_489);
and U1490 (N_1490,N_681,In_987);
nand U1491 (N_1491,In_2134,N_201);
xnor U1492 (N_1492,N_488,In_1109);
and U1493 (N_1493,In_672,N_784);
nor U1494 (N_1494,In_2387,N_582);
nor U1495 (N_1495,In_1321,In_981);
and U1496 (N_1496,In_1357,N_672);
xnor U1497 (N_1497,N_232,N_791);
or U1498 (N_1498,In_877,In_1943);
nand U1499 (N_1499,In_2001,In_2010);
and U1500 (N_1500,N_610,In_759);
or U1501 (N_1501,In_353,N_673);
nand U1502 (N_1502,In_2277,N_115);
and U1503 (N_1503,In_738,N_565);
xnor U1504 (N_1504,N_496,N_153);
nor U1505 (N_1505,N_236,In_1177);
xor U1506 (N_1506,N_421,In_543);
and U1507 (N_1507,In_1415,In_80);
and U1508 (N_1508,N_192,N_362);
nand U1509 (N_1509,In_950,In_461);
and U1510 (N_1510,N_613,N_402);
and U1511 (N_1511,N_231,N_632);
nor U1512 (N_1512,N_69,In_2222);
xnor U1513 (N_1513,N_448,In_2033);
and U1514 (N_1514,In_1988,N_504);
nand U1515 (N_1515,N_533,In_1410);
nand U1516 (N_1516,N_550,N_305);
nor U1517 (N_1517,N_663,N_528);
or U1518 (N_1518,N_648,N_722);
and U1519 (N_1519,In_2237,N_887);
nor U1520 (N_1520,N_649,In_1014);
nand U1521 (N_1521,N_191,N_798);
xnor U1522 (N_1522,N_735,N_248);
or U1523 (N_1523,N_556,In_2120);
nor U1524 (N_1524,In_1945,N_91);
xor U1525 (N_1525,N_477,N_126);
nor U1526 (N_1526,N_642,In_322);
nand U1527 (N_1527,N_882,N_396);
xnor U1528 (N_1528,N_405,N_282);
nor U1529 (N_1529,N_117,N_96);
or U1530 (N_1530,In_1893,N_944);
xnor U1531 (N_1531,N_464,N_976);
or U1532 (N_1532,N_422,N_100);
or U1533 (N_1533,N_500,In_2272);
nand U1534 (N_1534,N_771,In_1345);
xor U1535 (N_1535,N_687,N_563);
and U1536 (N_1536,N_11,N_574);
and U1537 (N_1537,N_39,N_483);
nor U1538 (N_1538,In_1285,N_629);
and U1539 (N_1539,N_322,N_540);
nand U1540 (N_1540,In_60,N_918);
xnor U1541 (N_1541,In_2060,In_1738);
xnor U1542 (N_1542,N_999,N_578);
nor U1543 (N_1543,N_240,In_12);
nor U1544 (N_1544,N_412,In_2023);
or U1545 (N_1545,In_677,In_1612);
or U1546 (N_1546,In_1556,In_1913);
and U1547 (N_1547,N_112,N_99);
or U1548 (N_1548,In_587,N_239);
or U1549 (N_1549,In_1604,In_2266);
nand U1550 (N_1550,N_472,N_429);
xnor U1551 (N_1551,N_853,In_2007);
nor U1552 (N_1552,In_1287,In_716);
nand U1553 (N_1553,N_9,N_637);
nor U1554 (N_1554,N_801,In_466);
nor U1555 (N_1555,N_586,In_1937);
xor U1556 (N_1556,N_878,N_688);
nand U1557 (N_1557,N_724,N_308);
xor U1558 (N_1558,In_335,N_536);
nand U1559 (N_1559,N_62,In_2020);
and U1560 (N_1560,In_1707,In_2190);
and U1561 (N_1561,N_802,In_1779);
and U1562 (N_1562,N_908,N_897);
nand U1563 (N_1563,N_419,In_2257);
nand U1564 (N_1564,N_4,N_919);
xor U1565 (N_1565,N_403,N_654);
and U1566 (N_1566,In_2415,N_38);
nor U1567 (N_1567,N_134,In_2012);
nor U1568 (N_1568,In_2305,In_1828);
nor U1569 (N_1569,In_2154,N_104);
and U1570 (N_1570,N_697,In_1003);
xor U1571 (N_1571,N_825,N_557);
and U1572 (N_1572,In_1040,N_686);
xnor U1573 (N_1573,N_297,N_199);
xnor U1574 (N_1574,N_211,N_452);
or U1575 (N_1575,N_281,N_468);
or U1576 (N_1576,N_52,N_348);
and U1577 (N_1577,N_684,In_2055);
or U1578 (N_1578,N_864,N_767);
nand U1579 (N_1579,N_731,In_1947);
or U1580 (N_1580,N_931,N_589);
xnor U1581 (N_1581,In_2069,In_632);
nor U1582 (N_1582,N_891,N_50);
nor U1583 (N_1583,In_1104,N_217);
xor U1584 (N_1584,N_570,N_929);
xnor U1585 (N_1585,N_669,N_365);
and U1586 (N_1586,In_1438,In_1331);
xnor U1587 (N_1587,In_1032,N_901);
xnor U1588 (N_1588,N_30,N_379);
nand U1589 (N_1589,N_180,In_2461);
nand U1590 (N_1590,N_804,In_1568);
nor U1591 (N_1591,In_1079,N_719);
nor U1592 (N_1592,N_493,N_424);
xnor U1593 (N_1593,In_2385,N_476);
or U1594 (N_1594,N_692,N_523);
nand U1595 (N_1595,N_325,N_176);
nor U1596 (N_1596,N_300,In_1022);
nand U1597 (N_1597,N_173,N_111);
xnor U1598 (N_1598,N_286,N_184);
and U1599 (N_1599,N_315,In_2459);
nand U1600 (N_1600,N_590,In_2327);
or U1601 (N_1601,In_1043,N_621);
nand U1602 (N_1602,N_140,N_84);
and U1603 (N_1603,N_818,N_997);
or U1604 (N_1604,In_59,In_1485);
or U1605 (N_1605,N_56,N_751);
and U1606 (N_1606,In_359,N_725);
and U1607 (N_1607,N_895,N_769);
xor U1608 (N_1608,N_515,In_1999);
nor U1609 (N_1609,N_455,N_934);
nand U1610 (N_1610,N_896,In_1242);
xor U1611 (N_1611,N_78,N_538);
nand U1612 (N_1612,N_81,In_2372);
nor U1613 (N_1613,In_235,N_926);
xnor U1614 (N_1614,In_742,In_993);
and U1615 (N_1615,In_506,N_558);
nand U1616 (N_1616,N_263,In_719);
and U1617 (N_1617,N_970,N_807);
nor U1618 (N_1618,In_659,N_181);
and U1619 (N_1619,In_1563,N_904);
or U1620 (N_1620,In_2240,N_886);
nor U1621 (N_1621,N_835,N_748);
nand U1622 (N_1622,N_942,In_2497);
xnor U1623 (N_1623,In_692,N_698);
or U1624 (N_1624,N_137,In_1047);
and U1625 (N_1625,In_1478,N_40);
and U1626 (N_1626,N_881,N_430);
nand U1627 (N_1627,In_1545,In_533);
nor U1628 (N_1628,N_372,N_603);
or U1629 (N_1629,N_799,In_732);
or U1630 (N_1630,N_93,In_1954);
nor U1631 (N_1631,N_61,N_159);
xnor U1632 (N_1632,N_910,In_618);
xnor U1633 (N_1633,N_921,In_679);
xor U1634 (N_1634,In_623,N_487);
nor U1635 (N_1635,In_377,N_875);
or U1636 (N_1636,In_934,N_200);
xor U1637 (N_1637,N_108,In_1343);
and U1638 (N_1638,In_1251,N_116);
nor U1639 (N_1639,In_1789,N_320);
xor U1640 (N_1640,N_198,N_491);
xor U1641 (N_1641,In_776,In_2311);
or U1642 (N_1642,N_293,N_577);
nor U1643 (N_1643,N_657,N_255);
and U1644 (N_1644,In_1519,N_334);
xnor U1645 (N_1645,N_561,N_770);
or U1646 (N_1646,N_551,N_978);
nand U1647 (N_1647,N_932,N_885);
and U1648 (N_1648,In_1185,In_1727);
nand U1649 (N_1649,In_665,In_1514);
xnor U1650 (N_1650,N_374,In_1178);
or U1651 (N_1651,N_872,N_631);
nor U1652 (N_1652,N_280,In_928);
nor U1653 (N_1653,N_359,In_741);
nand U1654 (N_1654,N_510,In_264);
or U1655 (N_1655,N_805,In_354);
nor U1656 (N_1656,In_2489,In_963);
nor U1657 (N_1657,N_964,N_346);
nand U1658 (N_1658,N_285,N_370);
nand U1659 (N_1659,N_381,In_720);
or U1660 (N_1660,In_412,N_689);
nor U1661 (N_1661,N_814,N_836);
and U1662 (N_1662,In_1232,N_883);
xor U1663 (N_1663,In_220,In_657);
or U1664 (N_1664,N_363,N_812);
nand U1665 (N_1665,N_387,N_992);
nor U1666 (N_1666,N_667,N_674);
nor U1667 (N_1667,N_726,N_810);
nor U1668 (N_1668,N_758,N_303);
nand U1669 (N_1669,In_1378,N_330);
or U1670 (N_1670,N_977,N_371);
and U1671 (N_1671,N_88,N_713);
xnor U1672 (N_1672,In_1784,N_393);
nor U1673 (N_1673,N_892,N_516);
xor U1674 (N_1674,N_842,N_660);
or U1675 (N_1675,N_776,In_2086);
and U1676 (N_1676,N_641,N_995);
or U1677 (N_1677,N_862,N_361);
nand U1678 (N_1678,N_397,N_622);
nor U1679 (N_1679,N_135,N_87);
and U1680 (N_1680,N_124,N_990);
xnor U1681 (N_1681,In_465,In_616);
xor U1682 (N_1682,In_2361,In_1156);
nor U1683 (N_1683,In_1390,In_2262);
xor U1684 (N_1684,In_1684,N_210);
and U1685 (N_1685,N_967,N_328);
nor U1686 (N_1686,N_581,N_793);
nor U1687 (N_1687,N_347,In_1642);
nor U1688 (N_1688,In_2245,In_490);
xnor U1689 (N_1689,In_247,N_549);
and U1690 (N_1690,N_602,In_1213);
nor U1691 (N_1691,N_701,In_20);
or U1692 (N_1692,N_414,In_1854);
or U1693 (N_1693,N_665,In_918);
xnor U1694 (N_1694,N_683,In_2293);
and U1695 (N_1695,In_2236,In_1627);
xnor U1696 (N_1696,N_174,In_2494);
and U1697 (N_1697,N_462,In_1608);
or U1698 (N_1698,N_433,N_79);
nand U1699 (N_1699,In_239,In_1750);
xnor U1700 (N_1700,N_573,In_2234);
nor U1701 (N_1701,N_611,In_1614);
and U1702 (N_1702,N_653,N_620);
nand U1703 (N_1703,In_48,N_962);
nand U1704 (N_1704,In_1045,In_2492);
or U1705 (N_1705,N_250,N_554);
nor U1706 (N_1706,In_2168,N_988);
or U1707 (N_1707,In_1312,In_1198);
xor U1708 (N_1708,N_968,N_925);
nand U1709 (N_1709,N_739,In_295);
and U1710 (N_1710,N_609,In_2176);
xnor U1711 (N_1711,N_195,N_349);
xor U1712 (N_1712,In_2392,N_273);
or U1713 (N_1713,N_542,N_624);
and U1714 (N_1714,N_635,N_125);
nor U1715 (N_1715,N_737,N_742);
or U1716 (N_1716,N_244,In_40);
xnor U1717 (N_1717,N_377,N_459);
xor U1718 (N_1718,N_699,N_158);
or U1719 (N_1719,In_1776,In_445);
xor U1720 (N_1720,N_485,In_1315);
and U1721 (N_1721,N_994,In_1575);
or U1722 (N_1722,N_264,In_1850);
nand U1723 (N_1723,N_246,In_2223);
xnor U1724 (N_1724,In_1838,N_785);
or U1725 (N_1725,N_781,N_351);
xor U1726 (N_1726,N_384,In_1423);
or U1727 (N_1727,N_659,In_2197);
xor U1728 (N_1728,In_1882,N_222);
xor U1729 (N_1729,N_357,N_323);
nand U1730 (N_1730,In_257,N_821);
or U1731 (N_1731,In_287,N_460);
nor U1732 (N_1732,N_339,In_358);
or U1733 (N_1733,N_298,N_413);
xor U1734 (N_1734,In_1513,In_2027);
nor U1735 (N_1735,In_952,N_68);
and U1736 (N_1736,N_259,In_559);
nand U1737 (N_1737,In_870,In_174);
xor U1738 (N_1738,In_474,In_1272);
and U1739 (N_1739,N_592,In_492);
and U1740 (N_1740,N_474,N_53);
nor U1741 (N_1741,N_401,N_585);
or U1742 (N_1742,In_2460,N_352);
nor U1743 (N_1743,In_1190,N_989);
xnor U1744 (N_1744,In_552,N_634);
xnor U1745 (N_1745,In_141,N_639);
xnor U1746 (N_1746,N_623,In_2251);
nand U1747 (N_1747,In_383,In_1461);
nor U1748 (N_1748,N_316,N_21);
nor U1749 (N_1749,In_211,In_537);
and U1750 (N_1750,N_286,In_928);
xnor U1751 (N_1751,In_2333,N_957);
xnor U1752 (N_1752,N_134,N_650);
nand U1753 (N_1753,N_214,N_299);
nand U1754 (N_1754,N_436,In_1969);
xnor U1755 (N_1755,N_883,N_673);
nand U1756 (N_1756,N_271,N_356);
xnor U1757 (N_1757,N_538,N_937);
or U1758 (N_1758,N_518,N_453);
nand U1759 (N_1759,N_87,N_701);
and U1760 (N_1760,N_764,N_578);
and U1761 (N_1761,In_1607,N_216);
or U1762 (N_1762,N_399,In_657);
and U1763 (N_1763,In_708,N_847);
xnor U1764 (N_1764,In_2374,N_264);
nand U1765 (N_1765,N_771,N_955);
nor U1766 (N_1766,In_1980,In_719);
xor U1767 (N_1767,N_344,N_231);
nand U1768 (N_1768,In_1461,N_214);
nor U1769 (N_1769,N_504,In_202);
and U1770 (N_1770,In_818,N_832);
or U1771 (N_1771,In_1662,N_839);
nand U1772 (N_1772,N_812,N_671);
or U1773 (N_1773,In_2110,In_623);
nand U1774 (N_1774,N_241,In_2154);
nand U1775 (N_1775,N_754,N_549);
xor U1776 (N_1776,In_2055,N_14);
nand U1777 (N_1777,In_1293,In_1513);
xor U1778 (N_1778,In_2385,N_668);
and U1779 (N_1779,In_1014,In_2);
xor U1780 (N_1780,N_49,N_923);
or U1781 (N_1781,In_2007,N_220);
xor U1782 (N_1782,N_891,N_452);
and U1783 (N_1783,N_542,In_2459);
nor U1784 (N_1784,N_690,In_988);
or U1785 (N_1785,In_81,N_582);
nand U1786 (N_1786,N_142,In_1232);
and U1787 (N_1787,N_139,N_692);
xor U1788 (N_1788,N_100,In_2429);
and U1789 (N_1789,In_1066,N_539);
and U1790 (N_1790,N_334,In_950);
or U1791 (N_1791,N_580,N_531);
nor U1792 (N_1792,N_845,In_1965);
xnor U1793 (N_1793,N_954,In_891);
xor U1794 (N_1794,In_1910,N_332);
and U1795 (N_1795,In_1087,N_387);
nor U1796 (N_1796,N_886,N_529);
nor U1797 (N_1797,N_858,N_464);
and U1798 (N_1798,N_974,N_824);
or U1799 (N_1799,N_532,N_625);
nor U1800 (N_1800,In_366,N_366);
xor U1801 (N_1801,N_612,In_2147);
or U1802 (N_1802,N_298,N_579);
and U1803 (N_1803,N_148,N_666);
xnor U1804 (N_1804,N_882,N_243);
nand U1805 (N_1805,N_105,N_744);
and U1806 (N_1806,N_345,N_341);
xnor U1807 (N_1807,In_2459,N_217);
nor U1808 (N_1808,In_2190,N_780);
and U1809 (N_1809,N_268,N_205);
nor U1810 (N_1810,In_335,N_98);
xor U1811 (N_1811,N_638,In_2);
or U1812 (N_1812,In_2059,N_462);
and U1813 (N_1813,N_50,In_2139);
nand U1814 (N_1814,N_691,N_593);
xnor U1815 (N_1815,N_962,In_2256);
nor U1816 (N_1816,N_271,N_179);
xnor U1817 (N_1817,In_1665,In_1197);
nand U1818 (N_1818,N_729,N_278);
nand U1819 (N_1819,N_684,N_683);
nand U1820 (N_1820,In_250,N_75);
and U1821 (N_1821,N_577,N_706);
nand U1822 (N_1822,N_902,In_988);
nand U1823 (N_1823,In_868,N_904);
or U1824 (N_1824,N_202,N_322);
nor U1825 (N_1825,N_642,N_836);
nand U1826 (N_1826,N_307,In_963);
or U1827 (N_1827,In_1188,N_669);
xor U1828 (N_1828,N_17,N_85);
or U1829 (N_1829,N_904,N_888);
or U1830 (N_1830,In_2477,In_2113);
and U1831 (N_1831,N_714,N_499);
or U1832 (N_1832,N_513,N_440);
nand U1833 (N_1833,N_719,In_665);
nor U1834 (N_1834,In_1342,N_819);
nand U1835 (N_1835,N_869,N_908);
and U1836 (N_1836,N_487,N_24);
and U1837 (N_1837,N_932,N_877);
and U1838 (N_1838,N_586,N_50);
xor U1839 (N_1839,N_183,N_477);
xnor U1840 (N_1840,N_850,In_62);
and U1841 (N_1841,N_816,N_390);
xor U1842 (N_1842,N_755,In_2082);
and U1843 (N_1843,N_716,N_132);
nor U1844 (N_1844,In_1607,In_1285);
nand U1845 (N_1845,N_428,In_1592);
and U1846 (N_1846,N_99,N_185);
nand U1847 (N_1847,N_681,N_984);
or U1848 (N_1848,N_869,N_683);
nand U1849 (N_1849,N_866,In_552);
or U1850 (N_1850,N_326,N_567);
nor U1851 (N_1851,In_918,N_550);
and U1852 (N_1852,In_1519,In_618);
and U1853 (N_1853,N_51,N_474);
or U1854 (N_1854,N_916,N_874);
nand U1855 (N_1855,N_670,N_254);
xnor U1856 (N_1856,N_492,N_691);
nor U1857 (N_1857,In_264,N_148);
nor U1858 (N_1858,N_684,N_118);
and U1859 (N_1859,N_64,N_636);
nand U1860 (N_1860,N_49,N_868);
xor U1861 (N_1861,In_126,N_946);
nor U1862 (N_1862,N_826,N_65);
nor U1863 (N_1863,In_1197,In_1784);
nor U1864 (N_1864,N_610,In_247);
or U1865 (N_1865,In_1461,N_232);
or U1866 (N_1866,N_747,N_734);
or U1867 (N_1867,In_735,N_564);
nand U1868 (N_1868,In_1273,N_797);
nand U1869 (N_1869,N_664,N_853);
nor U1870 (N_1870,N_434,N_724);
or U1871 (N_1871,N_939,N_221);
xor U1872 (N_1872,N_192,In_1871);
or U1873 (N_1873,N_756,In_12);
and U1874 (N_1874,In_1487,N_922);
and U1875 (N_1875,N_321,N_289);
nor U1876 (N_1876,In_1947,N_923);
or U1877 (N_1877,In_133,In_454);
or U1878 (N_1878,N_513,N_966);
or U1879 (N_1879,N_739,In_59);
and U1880 (N_1880,N_161,N_908);
xor U1881 (N_1881,In_2494,In_2277);
nand U1882 (N_1882,N_325,In_1045);
or U1883 (N_1883,In_877,In_2333);
nand U1884 (N_1884,In_680,N_419);
nand U1885 (N_1885,In_1325,In_2168);
or U1886 (N_1886,In_172,N_980);
nand U1887 (N_1887,In_474,In_808);
xnor U1888 (N_1888,N_525,In_2134);
xnor U1889 (N_1889,In_2333,In_540);
nor U1890 (N_1890,N_460,N_261);
or U1891 (N_1891,N_575,N_304);
nor U1892 (N_1892,N_64,N_248);
nor U1893 (N_1893,In_1043,N_829);
or U1894 (N_1894,N_481,In_239);
nor U1895 (N_1895,N_419,N_4);
or U1896 (N_1896,N_507,N_676);
nor U1897 (N_1897,In_2120,N_701);
nor U1898 (N_1898,N_655,N_267);
nand U1899 (N_1899,N_147,In_583);
xor U1900 (N_1900,In_875,In_952);
and U1901 (N_1901,N_551,N_953);
or U1902 (N_1902,N_661,N_715);
and U1903 (N_1903,N_480,N_892);
or U1904 (N_1904,In_81,N_371);
or U1905 (N_1905,N_399,In_2188);
and U1906 (N_1906,In_1537,N_286);
xnor U1907 (N_1907,N_502,In_2277);
and U1908 (N_1908,N_142,In_1892);
nand U1909 (N_1909,In_2251,N_734);
nor U1910 (N_1910,In_264,In_950);
nor U1911 (N_1911,N_475,In_1592);
and U1912 (N_1912,In_1242,In_174);
or U1913 (N_1913,N_43,In_2256);
xor U1914 (N_1914,N_704,In_1627);
xnor U1915 (N_1915,In_1185,N_974);
nand U1916 (N_1916,N_946,N_62);
nor U1917 (N_1917,In_60,N_929);
or U1918 (N_1918,N_869,N_634);
or U1919 (N_1919,N_947,In_1884);
nor U1920 (N_1920,N_22,N_631);
or U1921 (N_1921,N_888,N_807);
nor U1922 (N_1922,In_870,N_15);
and U1923 (N_1923,N_576,N_903);
nand U1924 (N_1924,N_76,N_939);
xnor U1925 (N_1925,N_323,N_709);
or U1926 (N_1926,In_2092,In_535);
nand U1927 (N_1927,N_734,In_523);
or U1928 (N_1928,N_277,N_248);
nand U1929 (N_1929,N_465,N_43);
nor U1930 (N_1930,N_720,N_476);
or U1931 (N_1931,N_969,N_749);
xnor U1932 (N_1932,N_16,N_123);
xnor U1933 (N_1933,N_10,N_483);
xnor U1934 (N_1934,N_755,In_2069);
nand U1935 (N_1935,N_909,N_278);
nor U1936 (N_1936,N_358,N_515);
nor U1937 (N_1937,N_739,N_734);
nand U1938 (N_1938,N_2,N_960);
nor U1939 (N_1939,N_396,N_241);
xnor U1940 (N_1940,N_243,N_18);
or U1941 (N_1941,N_363,N_496);
or U1942 (N_1942,N_633,N_916);
nor U1943 (N_1943,N_615,N_43);
nor U1944 (N_1944,N_444,N_767);
xnor U1945 (N_1945,In_20,In_2367);
xnor U1946 (N_1946,N_511,N_111);
xnor U1947 (N_1947,N_980,N_220);
nor U1948 (N_1948,N_536,In_1109);
xnor U1949 (N_1949,N_228,N_892);
nor U1950 (N_1950,In_1397,N_377);
or U1951 (N_1951,N_395,N_3);
and U1952 (N_1952,In_1570,N_487);
or U1953 (N_1953,N_670,N_580);
nor U1954 (N_1954,In_800,In_1704);
and U1955 (N_1955,N_955,In_934);
nor U1956 (N_1956,In_2134,N_280);
or U1957 (N_1957,N_519,N_195);
nand U1958 (N_1958,N_333,N_468);
nor U1959 (N_1959,N_45,N_662);
or U1960 (N_1960,N_136,N_87);
and U1961 (N_1961,N_7,N_207);
or U1962 (N_1962,N_384,In_1063);
or U1963 (N_1963,In_952,N_494);
xnor U1964 (N_1964,In_1123,N_463);
and U1965 (N_1965,N_70,N_509);
nor U1966 (N_1966,N_88,In_490);
xnor U1967 (N_1967,N_636,N_696);
nand U1968 (N_1968,In_1325,N_398);
or U1969 (N_1969,In_762,N_459);
xor U1970 (N_1970,N_971,N_459);
nand U1971 (N_1971,N_958,N_333);
and U1972 (N_1972,In_1079,N_549);
or U1973 (N_1973,N_840,In_1376);
nor U1974 (N_1974,N_909,N_598);
xnor U1975 (N_1975,In_177,N_534);
or U1976 (N_1976,N_771,N_226);
or U1977 (N_1977,N_806,N_715);
nor U1978 (N_1978,In_2095,N_173);
and U1979 (N_1979,N_645,In_2061);
xnor U1980 (N_1980,In_308,N_414);
or U1981 (N_1981,N_798,N_500);
nand U1982 (N_1982,N_257,In_2);
nor U1983 (N_1983,N_630,In_2489);
and U1984 (N_1984,In_1009,N_600);
nor U1985 (N_1985,N_209,N_315);
nand U1986 (N_1986,In_1185,N_931);
xor U1987 (N_1987,N_301,In_818);
xor U1988 (N_1988,N_423,N_63);
nor U1989 (N_1989,N_545,N_60);
xor U1990 (N_1990,N_741,N_436);
or U1991 (N_1991,In_1784,N_172);
xor U1992 (N_1992,N_684,N_103);
nor U1993 (N_1993,In_2062,N_476);
or U1994 (N_1994,N_714,N_336);
and U1995 (N_1995,N_755,N_557);
nand U1996 (N_1996,N_528,N_374);
or U1997 (N_1997,N_878,N_213);
xor U1998 (N_1998,N_217,N_268);
or U1999 (N_1999,In_1665,In_574);
or U2000 (N_2000,N_1052,N_1050);
or U2001 (N_2001,N_1143,N_1276);
xnor U2002 (N_2002,N_1381,N_1077);
or U2003 (N_2003,N_1378,N_1010);
nor U2004 (N_2004,N_1836,N_1533);
nand U2005 (N_2005,N_1066,N_1762);
nand U2006 (N_2006,N_1815,N_1142);
or U2007 (N_2007,N_1277,N_1203);
nand U2008 (N_2008,N_1095,N_1356);
or U2009 (N_2009,N_1526,N_1910);
xnor U2010 (N_2010,N_1907,N_1484);
or U2011 (N_2011,N_1185,N_1508);
or U2012 (N_2012,N_1574,N_1666);
nand U2013 (N_2013,N_1956,N_1531);
or U2014 (N_2014,N_1818,N_1935);
nand U2015 (N_2015,N_1544,N_1013);
nor U2016 (N_2016,N_1228,N_1237);
nor U2017 (N_2017,N_1596,N_1992);
xnor U2018 (N_2018,N_1546,N_1780);
and U2019 (N_2019,N_1857,N_1254);
nand U2020 (N_2020,N_1941,N_1957);
nand U2021 (N_2021,N_1012,N_1991);
or U2022 (N_2022,N_1832,N_1045);
and U2023 (N_2023,N_1986,N_1248);
and U2024 (N_2024,N_1782,N_1459);
xnor U2025 (N_2025,N_1244,N_1483);
and U2026 (N_2026,N_1668,N_1914);
nor U2027 (N_2027,N_1583,N_1690);
nand U2028 (N_2028,N_1336,N_1498);
and U2029 (N_2029,N_1979,N_1220);
or U2030 (N_2030,N_1494,N_1427);
and U2031 (N_2031,N_1132,N_1809);
and U2032 (N_2032,N_1232,N_1698);
or U2033 (N_2033,N_1094,N_1783);
nand U2034 (N_2034,N_1672,N_1161);
xnor U2035 (N_2035,N_1437,N_1333);
xnor U2036 (N_2036,N_1263,N_1478);
nor U2037 (N_2037,N_1100,N_1730);
or U2038 (N_2038,N_1476,N_1577);
and U2039 (N_2039,N_1227,N_1694);
nor U2040 (N_2040,N_1485,N_1587);
and U2041 (N_2041,N_1075,N_1453);
nand U2042 (N_2042,N_1300,N_1819);
nand U2043 (N_2043,N_1324,N_1491);
and U2044 (N_2044,N_1908,N_1864);
or U2045 (N_2045,N_1404,N_1977);
nand U2046 (N_2046,N_1684,N_1497);
or U2047 (N_2047,N_1359,N_1616);
nand U2048 (N_2048,N_1482,N_1353);
and U2049 (N_2049,N_1656,N_1887);
xor U2050 (N_2050,N_1791,N_1880);
nand U2051 (N_2051,N_1322,N_1234);
nor U2052 (N_2052,N_1190,N_1868);
xnor U2053 (N_2053,N_1273,N_1924);
nand U2054 (N_2054,N_1997,N_1499);
xnor U2055 (N_2055,N_1509,N_1090);
nor U2056 (N_2056,N_1905,N_1942);
nor U2057 (N_2057,N_1446,N_1029);
and U2058 (N_2058,N_1529,N_1993);
and U2059 (N_2059,N_1795,N_1397);
and U2060 (N_2060,N_1319,N_1418);
nor U2061 (N_2061,N_1629,N_1267);
nand U2062 (N_2062,N_1704,N_1054);
or U2063 (N_2063,N_1842,N_1088);
and U2064 (N_2064,N_1944,N_1586);
or U2065 (N_2065,N_1206,N_1843);
nand U2066 (N_2066,N_1584,N_1189);
nor U2067 (N_2067,N_1712,N_1387);
nor U2068 (N_2068,N_1652,N_1466);
nand U2069 (N_2069,N_1834,N_1999);
or U2070 (N_2070,N_1802,N_1970);
nand U2071 (N_2071,N_1817,N_1022);
nor U2072 (N_2072,N_1810,N_1166);
nor U2073 (N_2073,N_1108,N_1624);
or U2074 (N_2074,N_1049,N_1718);
nand U2075 (N_2075,N_1384,N_1511);
nand U2076 (N_2076,N_1737,N_1726);
xor U2077 (N_2077,N_1673,N_1686);
nor U2078 (N_2078,N_1229,N_1177);
nor U2079 (N_2079,N_1891,N_1106);
xnor U2080 (N_2080,N_1148,N_1713);
or U2081 (N_2081,N_1146,N_1444);
nor U2082 (N_2082,N_1565,N_1931);
or U2083 (N_2083,N_1503,N_1197);
nor U2084 (N_2084,N_1110,N_1119);
or U2085 (N_2085,N_1994,N_1948);
xor U2086 (N_2086,N_1937,N_1352);
xnor U2087 (N_2087,N_1055,N_1566);
nor U2088 (N_2088,N_1501,N_1240);
nor U2089 (N_2089,N_1530,N_1245);
xnor U2090 (N_2090,N_1572,N_1215);
or U2091 (N_2091,N_1424,N_1136);
nor U2092 (N_2092,N_1304,N_1609);
or U2093 (N_2093,N_1893,N_1377);
or U2094 (N_2094,N_1047,N_1770);
and U2095 (N_2095,N_1123,N_1109);
nor U2096 (N_2096,N_1676,N_1920);
nor U2097 (N_2097,N_1663,N_1811);
nand U2098 (N_2098,N_1379,N_1084);
xnor U2099 (N_2099,N_1514,N_1329);
nand U2100 (N_2100,N_1440,N_1293);
xor U2101 (N_2101,N_1207,N_1939);
nor U2102 (N_2102,N_1775,N_1291);
nand U2103 (N_2103,N_1350,N_1214);
nand U2104 (N_2104,N_1985,N_1035);
and U2105 (N_2105,N_1854,N_1168);
nand U2106 (N_2106,N_1925,N_1724);
xor U2107 (N_2107,N_1205,N_1496);
xor U2108 (N_2108,N_1432,N_1470);
and U2109 (N_2109,N_1703,N_1820);
xnor U2110 (N_2110,N_1442,N_1978);
xor U2111 (N_2111,N_1890,N_1705);
xor U2112 (N_2112,N_1246,N_1238);
xnor U2113 (N_2113,N_1830,N_1431);
nand U2114 (N_2114,N_1539,N_1328);
nor U2115 (N_2115,N_1112,N_1623);
nor U2116 (N_2116,N_1715,N_1471);
nor U2117 (N_2117,N_1990,N_1492);
nor U2118 (N_2118,N_1315,N_1043);
xnor U2119 (N_2119,N_1848,N_1216);
nand U2120 (N_2120,N_1631,N_1635);
and U2121 (N_2121,N_1252,N_1493);
or U2122 (N_2122,N_1430,N_1294);
and U2123 (N_2123,N_1633,N_1875);
nand U2124 (N_2124,N_1621,N_1217);
and U2125 (N_2125,N_1688,N_1695);
and U2126 (N_2126,N_1464,N_1318);
or U2127 (N_2127,N_1786,N_1561);
xor U2128 (N_2128,N_1973,N_1534);
xnor U2129 (N_2129,N_1133,N_1756);
or U2130 (N_2130,N_1524,N_1916);
and U2131 (N_2131,N_1736,N_1398);
nand U2132 (N_2132,N_1428,N_1570);
and U2133 (N_2133,N_1522,N_1996);
and U2134 (N_2134,N_1439,N_1846);
nor U2135 (N_2135,N_1327,N_1323);
nor U2136 (N_2136,N_1760,N_1982);
xnor U2137 (N_2137,N_1212,N_1460);
or U2138 (N_2138,N_1821,N_1900);
xnor U2139 (N_2139,N_1989,N_1056);
xnor U2140 (N_2140,N_1950,N_1487);
nor U2141 (N_2141,N_1320,N_1373);
nand U2142 (N_2142,N_1800,N_1241);
and U2143 (N_2143,N_1946,N_1061);
xor U2144 (N_2144,N_1157,N_1902);
and U2145 (N_2145,N_1287,N_1627);
nand U2146 (N_2146,N_1193,N_1505);
xor U2147 (N_2147,N_1375,N_1002);
nor U2148 (N_2148,N_1284,N_1257);
or U2149 (N_2149,N_1311,N_1003);
nand U2150 (N_2150,N_1763,N_1341);
xnor U2151 (N_2151,N_1733,N_1648);
or U2152 (N_2152,N_1417,N_1018);
or U2153 (N_2153,N_1844,N_1401);
or U2154 (N_2154,N_1292,N_1568);
or U2155 (N_2155,N_1281,N_1500);
xnor U2156 (N_2156,N_1051,N_1681);
nand U2157 (N_2157,N_1380,N_1269);
xor U2158 (N_2158,N_1007,N_1934);
and U2159 (N_2159,N_1863,N_1972);
nor U2160 (N_2160,N_1741,N_1364);
and U2161 (N_2161,N_1664,N_1504);
and U2162 (N_2162,N_1735,N_1171);
nor U2163 (N_2163,N_1537,N_1877);
xnor U2164 (N_2164,N_1553,N_1144);
nand U2165 (N_2165,N_1567,N_1366);
and U2166 (N_2166,N_1610,N_1048);
and U2167 (N_2167,N_1831,N_1167);
or U2168 (N_2168,N_1871,N_1789);
xnor U2169 (N_2169,N_1679,N_1474);
and U2170 (N_2170,N_1159,N_1141);
nand U2171 (N_2171,N_1345,N_1951);
xnor U2172 (N_2172,N_1779,N_1469);
nand U2173 (N_2173,N_1298,N_1776);
nand U2174 (N_2174,N_1701,N_1727);
or U2175 (N_2175,N_1837,N_1289);
nor U2176 (N_2176,N_1005,N_1600);
nand U2177 (N_2177,N_1130,N_1646);
xor U2178 (N_2178,N_1608,N_1001);
and U2179 (N_2179,N_1243,N_1117);
nor U2180 (N_2180,N_1351,N_1344);
or U2181 (N_2181,N_1016,N_1078);
nor U2182 (N_2182,N_1115,N_1137);
or U2183 (N_2183,N_1231,N_1236);
nor U2184 (N_2184,N_1034,N_1552);
or U2185 (N_2185,N_1467,N_1588);
and U2186 (N_2186,N_1649,N_1692);
and U2187 (N_2187,N_1156,N_1172);
nand U2188 (N_2188,N_1677,N_1784);
and U2189 (N_2189,N_1625,N_1067);
nand U2190 (N_2190,N_1962,N_1771);
nor U2191 (N_2191,N_1725,N_1873);
or U2192 (N_2192,N_1974,N_1180);
nor U2193 (N_2193,N_1481,N_1472);
or U2194 (N_2194,N_1279,N_1098);
nor U2195 (N_2195,N_1268,N_1886);
xor U2196 (N_2196,N_1987,N_1798);
or U2197 (N_2197,N_1731,N_1285);
nor U2198 (N_2198,N_1423,N_1706);
or U2199 (N_2199,N_1976,N_1402);
nand U2200 (N_2200,N_1879,N_1461);
nand U2201 (N_2201,N_1255,N_1295);
and U2202 (N_2202,N_1420,N_1175);
or U2203 (N_2203,N_1126,N_1599);
and U2204 (N_2204,N_1326,N_1097);
or U2205 (N_2205,N_1995,N_1198);
nor U2206 (N_2206,N_1302,N_1611);
xor U2207 (N_2207,N_1564,N_1580);
xnor U2208 (N_2208,N_1286,N_1169);
nor U2209 (N_2209,N_1393,N_1516);
and U2210 (N_2210,N_1918,N_1980);
nor U2211 (N_2211,N_1274,N_1219);
nand U2212 (N_2212,N_1452,N_1921);
and U2213 (N_2213,N_1260,N_1363);
nor U2214 (N_2214,N_1801,N_1058);
nand U2215 (N_2215,N_1806,N_1194);
and U2216 (N_2216,N_1099,N_1540);
and U2217 (N_2217,N_1340,N_1549);
or U2218 (N_2218,N_1201,N_1176);
nand U2219 (N_2219,N_1573,N_1693);
xnor U2220 (N_2220,N_1885,N_1707);
nand U2221 (N_2221,N_1181,N_1096);
xnor U2222 (N_2222,N_1738,N_1256);
or U2223 (N_2223,N_1264,N_1657);
or U2224 (N_2224,N_1755,N_1745);
nor U2225 (N_2225,N_1338,N_1647);
nor U2226 (N_2226,N_1342,N_1556);
and U2227 (N_2227,N_1637,N_1395);
and U2228 (N_2228,N_1039,N_1129);
and U2229 (N_2229,N_1932,N_1278);
xor U2230 (N_2230,N_1547,N_1523);
nand U2231 (N_2231,N_1445,N_1369);
xnor U2232 (N_2232,N_1060,N_1032);
or U2233 (N_2233,N_1774,N_1486);
nand U2234 (N_2234,N_1334,N_1984);
and U2235 (N_2235,N_1744,N_1532);
or U2236 (N_2236,N_1262,N_1845);
and U2237 (N_2237,N_1799,N_1113);
or U2238 (N_2238,N_1027,N_1408);
or U2239 (N_2239,N_1301,N_1772);
or U2240 (N_2240,N_1081,N_1926);
nor U2241 (N_2241,N_1165,N_1680);
and U2242 (N_2242,N_1697,N_1915);
xnor U2243 (N_2243,N_1714,N_1665);
or U2244 (N_2244,N_1785,N_1952);
or U2245 (N_2245,N_1917,N_1923);
and U2246 (N_2246,N_1768,N_1020);
xor U2247 (N_2247,N_1959,N_1696);
nor U2248 (N_2248,N_1101,N_1019);
nor U2249 (N_2249,N_1904,N_1033);
nor U2250 (N_2250,N_1813,N_1797);
or U2251 (N_2251,N_1150,N_1740);
nand U2252 (N_2252,N_1839,N_1669);
xor U2253 (N_2253,N_1147,N_1451);
nand U2254 (N_2254,N_1441,N_1971);
and U2255 (N_2255,N_1218,N_1938);
and U2256 (N_2256,N_1030,N_1897);
nor U2257 (N_2257,N_1475,N_1325);
nand U2258 (N_2258,N_1860,N_1687);
and U2259 (N_2259,N_1662,N_1009);
nor U2260 (N_2260,N_1296,N_1722);
and U2261 (N_2261,N_1211,N_1757);
and U2262 (N_2262,N_1548,N_1089);
and U2263 (N_2263,N_1747,N_1833);
xor U2264 (N_2264,N_1729,N_1140);
xor U2265 (N_2265,N_1913,N_1660);
or U2266 (N_2266,N_1513,N_1793);
and U2267 (N_2267,N_1188,N_1601);
nor U2268 (N_2268,N_1275,N_1495);
nor U2269 (N_2269,N_1415,N_1645);
and U2270 (N_2270,N_1856,N_1360);
nor U2271 (N_2271,N_1015,N_1391);
xor U2272 (N_2272,N_1357,N_1655);
and U2273 (N_2273,N_1116,N_1138);
and U2274 (N_2274,N_1909,N_1752);
or U2275 (N_2275,N_1355,N_1271);
nor U2276 (N_2276,N_1571,N_1720);
xnor U2277 (N_2277,N_1781,N_1878);
xor U2278 (N_2278,N_1557,N_1603);
xor U2279 (N_2279,N_1807,N_1865);
nor U2280 (N_2280,N_1683,N_1210);
and U2281 (N_2281,N_1554,N_1396);
xnor U2282 (N_2282,N_1414,N_1576);
nand U2283 (N_2283,N_1528,N_1195);
xor U2284 (N_2284,N_1105,N_1826);
or U2285 (N_2285,N_1164,N_1685);
nand U2286 (N_2286,N_1111,N_1899);
nand U2287 (N_2287,N_1024,N_1390);
or U2288 (N_2288,N_1889,N_1847);
nor U2289 (N_2289,N_1896,N_1881);
xnor U2290 (N_2290,N_1450,N_1827);
or U2291 (N_2291,N_1983,N_1183);
nor U2292 (N_2292,N_1882,N_1765);
and U2293 (N_2293,N_1796,N_1717);
or U2294 (N_2294,N_1125,N_1367);
and U2295 (N_2295,N_1410,N_1225);
and U2296 (N_2296,N_1372,N_1949);
and U2297 (N_2297,N_1739,N_1804);
nor U2298 (N_2298,N_1803,N_1604);
nand U2299 (N_2299,N_1041,N_1409);
nor U2300 (N_2300,N_1894,N_1605);
xor U2301 (N_2301,N_1788,N_1011);
or U2302 (N_2302,N_1331,N_1640);
and U2303 (N_2303,N_1025,N_1426);
and U2304 (N_2304,N_1922,N_1134);
or U2305 (N_2305,N_1407,N_1063);
xnor U2306 (N_2306,N_1967,N_1163);
nor U2307 (N_2307,N_1242,N_1912);
nand U2308 (N_2308,N_1966,N_1700);
or U2309 (N_2309,N_1307,N_1152);
or U2310 (N_2310,N_1006,N_1859);
nor U2311 (N_2311,N_1591,N_1139);
or U2312 (N_2312,N_1840,N_1449);
nor U2313 (N_2313,N_1512,N_1658);
or U2314 (N_2314,N_1749,N_1422);
nand U2315 (N_2315,N_1614,N_1230);
nor U2316 (N_2316,N_1585,N_1044);
nor U2317 (N_2317,N_1767,N_1065);
xor U2318 (N_2318,N_1038,N_1149);
xnor U2319 (N_2319,N_1928,N_1288);
or U2320 (N_2320,N_1639,N_1456);
nor U2321 (N_2321,N_1200,N_1617);
xor U2322 (N_2322,N_1028,N_1728);
and U2323 (N_2323,N_1644,N_1187);
or U2324 (N_2324,N_1515,N_1064);
nor U2325 (N_2325,N_1874,N_1317);
nand U2326 (N_2326,N_1435,N_1308);
nand U2327 (N_2327,N_1135,N_1947);
or U2328 (N_2328,N_1702,N_1343);
nand U2329 (N_2329,N_1869,N_1400);
nand U2330 (N_2330,N_1154,N_1208);
nor U2331 (N_2331,N_1835,N_1790);
nor U2332 (N_2332,N_1930,N_1622);
and U2333 (N_2333,N_1578,N_1936);
and U2334 (N_2334,N_1371,N_1719);
or U2335 (N_2335,N_1259,N_1732);
nand U2336 (N_2336,N_1607,N_1517);
xor U2337 (N_2337,N_1209,N_1634);
nand U2338 (N_2338,N_1661,N_1121);
and U2339 (N_2339,N_1734,N_1448);
xor U2340 (N_2340,N_1087,N_1862);
or U2341 (N_2341,N_1822,N_1076);
xor U2342 (N_2342,N_1870,N_1433);
and U2343 (N_2343,N_1222,N_1825);
nand U2344 (N_2344,N_1419,N_1678);
or U2345 (N_2345,N_1346,N_1828);
and U2346 (N_2346,N_1093,N_1838);
xor U2347 (N_2347,N_1309,N_1266);
or U2348 (N_2348,N_1754,N_1592);
and U2349 (N_2349,N_1155,N_1017);
and U2350 (N_2350,N_1455,N_1674);
xnor U2351 (N_2351,N_1849,N_1330);
xor U2352 (N_2352,N_1250,N_1861);
or U2353 (N_2353,N_1597,N_1883);
and U2354 (N_2354,N_1965,N_1794);
and U2355 (N_2355,N_1858,N_1429);
xnor U2356 (N_2356,N_1290,N_1316);
xor U2357 (N_2357,N_1312,N_1385);
xnor U2358 (N_2358,N_1969,N_1299);
nand U2359 (N_2359,N_1283,N_1462);
nor U2360 (N_2360,N_1955,N_1204);
nor U2361 (N_2361,N_1083,N_1223);
nand U2362 (N_2362,N_1743,N_1510);
and U2363 (N_2363,N_1620,N_1349);
or U2364 (N_2364,N_1542,N_1746);
and U2365 (N_2365,N_1068,N_1598);
or U2366 (N_2366,N_1479,N_1691);
xor U2367 (N_2367,N_1590,N_1521);
xor U2368 (N_2368,N_1394,N_1280);
xor U2369 (N_2369,N_1911,N_1436);
nand U2370 (N_2370,N_1368,N_1468);
nand U2371 (N_2371,N_1416,N_1235);
nor U2372 (N_2372,N_1708,N_1008);
or U2373 (N_2373,N_1758,N_1569);
nor U2374 (N_2374,N_1853,N_1773);
or U2375 (N_2375,N_1122,N_1642);
nand U2376 (N_2376,N_1618,N_1748);
nor U2377 (N_2377,N_1619,N_1406);
or U2378 (N_2378,N_1411,N_1816);
nor U2379 (N_2379,N_1104,N_1761);
nand U2380 (N_2380,N_1575,N_1502);
and U2381 (N_2381,N_1382,N_1593);
xor U2382 (N_2382,N_1927,N_1270);
or U2383 (N_2383,N_1091,N_1388);
and U2384 (N_2384,N_1901,N_1626);
nor U2385 (N_2385,N_1551,N_1457);
nor U2386 (N_2386,N_1425,N_1852);
or U2387 (N_2387,N_1124,N_1589);
and U2388 (N_2388,N_1153,N_1310);
and U2389 (N_2389,N_1536,N_1594);
nor U2390 (N_2390,N_1313,N_1906);
nand U2391 (N_2391,N_1612,N_1337);
and U2392 (N_2392,N_1438,N_1253);
xnor U2393 (N_2393,N_1667,N_1777);
and U2394 (N_2394,N_1872,N_1651);
nand U2395 (N_2395,N_1145,N_1102);
xor U2396 (N_2396,N_1563,N_1160);
nor U2397 (N_2397,N_1389,N_1919);
nor U2398 (N_2398,N_1332,N_1092);
nor U2399 (N_2399,N_1057,N_1792);
and U2400 (N_2400,N_1710,N_1042);
nor U2401 (N_2401,N_1477,N_1850);
nor U2402 (N_2402,N_1347,N_1659);
and U2403 (N_2403,N_1233,N_1202);
xnor U2404 (N_2404,N_1374,N_1151);
nand U2405 (N_2405,N_1463,N_1829);
xor U2406 (N_2406,N_1898,N_1615);
and U2407 (N_2407,N_1582,N_1014);
and U2408 (N_2408,N_1953,N_1321);
and U2409 (N_2409,N_1545,N_1753);
and U2410 (N_2410,N_1670,N_1370);
and U2411 (N_2411,N_1386,N_1335);
or U2412 (N_2412,N_1541,N_1527);
and U2413 (N_2413,N_1682,N_1812);
nor U2414 (N_2414,N_1412,N_1535);
xor U2415 (N_2415,N_1559,N_1399);
or U2416 (N_2416,N_1162,N_1787);
nand U2417 (N_2417,N_1689,N_1128);
and U2418 (N_2418,N_1653,N_1506);
xnor U2419 (N_2419,N_1628,N_1488);
xor U2420 (N_2420,N_1037,N_1630);
nor U2421 (N_2421,N_1884,N_1723);
xor U2422 (N_2422,N_1403,N_1000);
nor U2423 (N_2423,N_1489,N_1766);
or U2424 (N_2424,N_1383,N_1595);
or U2425 (N_2425,N_1179,N_1158);
or U2426 (N_2426,N_1004,N_1173);
xnor U2427 (N_2427,N_1988,N_1750);
nand U2428 (N_2428,N_1114,N_1876);
and U2429 (N_2429,N_1447,N_1954);
nor U2430 (N_2430,N_1348,N_1251);
and U2431 (N_2431,N_1888,N_1711);
xnor U2432 (N_2432,N_1841,N_1303);
or U2433 (N_2433,N_1520,N_1103);
or U2434 (N_2434,N_1632,N_1434);
nand U2435 (N_2435,N_1354,N_1072);
and U2436 (N_2436,N_1558,N_1361);
nand U2437 (N_2437,N_1074,N_1960);
nand U2438 (N_2438,N_1080,N_1261);
or U2439 (N_2439,N_1602,N_1855);
nor U2440 (N_2440,N_1036,N_1062);
and U2441 (N_2441,N_1636,N_1555);
or U2442 (N_2442,N_1454,N_1606);
nand U2443 (N_2443,N_1525,N_1507);
nor U2444 (N_2444,N_1823,N_1943);
nor U2445 (N_2445,N_1265,N_1824);
nor U2446 (N_2446,N_1131,N_1413);
nand U2447 (N_2447,N_1107,N_1339);
xor U2448 (N_2448,N_1895,N_1769);
nor U2449 (N_2449,N_1358,N_1085);
or U2450 (N_2450,N_1643,N_1282);
xor U2451 (N_2451,N_1073,N_1239);
and U2452 (N_2452,N_1945,N_1082);
or U2453 (N_2453,N_1675,N_1069);
nor U2454 (N_2454,N_1026,N_1405);
nor U2455 (N_2455,N_1964,N_1981);
or U2456 (N_2456,N_1805,N_1184);
xnor U2457 (N_2457,N_1550,N_1751);
or U2458 (N_2458,N_1851,N_1314);
or U2459 (N_2459,N_1046,N_1581);
nand U2460 (N_2460,N_1272,N_1053);
or U2461 (N_2461,N_1305,N_1473);
or U2462 (N_2462,N_1178,N_1023);
nor U2463 (N_2463,N_1903,N_1808);
or U2464 (N_2464,N_1716,N_1968);
nand U2465 (N_2465,N_1306,N_1086);
or U2466 (N_2466,N_1070,N_1196);
or U2467 (N_2467,N_1933,N_1031);
nand U2468 (N_2468,N_1249,N_1365);
and U2469 (N_2469,N_1699,N_1543);
and U2470 (N_2470,N_1654,N_1940);
xor U2471 (N_2471,N_1538,N_1465);
or U2472 (N_2472,N_1079,N_1579);
or U2473 (N_2473,N_1224,N_1226);
nor U2474 (N_2474,N_1998,N_1421);
nand U2475 (N_2475,N_1120,N_1458);
xor U2476 (N_2476,N_1519,N_1021);
and U2477 (N_2477,N_1170,N_1186);
xnor U2478 (N_2478,N_1759,N_1192);
nor U2479 (N_2479,N_1778,N_1127);
xnor U2480 (N_2480,N_1867,N_1480);
or U2481 (N_2481,N_1059,N_1376);
nor U2482 (N_2482,N_1742,N_1199);
or U2483 (N_2483,N_1764,N_1392);
nand U2484 (N_2484,N_1650,N_1040);
and U2485 (N_2485,N_1975,N_1518);
or U2486 (N_2486,N_1958,N_1297);
nand U2487 (N_2487,N_1641,N_1613);
xnor U2488 (N_2488,N_1671,N_1638);
nor U2489 (N_2489,N_1191,N_1247);
xor U2490 (N_2490,N_1221,N_1362);
and U2491 (N_2491,N_1961,N_1560);
nand U2492 (N_2492,N_1443,N_1963);
nor U2493 (N_2493,N_1258,N_1174);
nand U2494 (N_2494,N_1929,N_1866);
and U2495 (N_2495,N_1490,N_1562);
xnor U2496 (N_2496,N_1118,N_1213);
xor U2497 (N_2497,N_1182,N_1709);
xor U2498 (N_2498,N_1721,N_1071);
nand U2499 (N_2499,N_1892,N_1814);
or U2500 (N_2500,N_1462,N_1311);
and U2501 (N_2501,N_1377,N_1468);
nor U2502 (N_2502,N_1665,N_1482);
nor U2503 (N_2503,N_1889,N_1065);
nand U2504 (N_2504,N_1346,N_1339);
and U2505 (N_2505,N_1187,N_1354);
xnor U2506 (N_2506,N_1558,N_1511);
xor U2507 (N_2507,N_1724,N_1289);
nor U2508 (N_2508,N_1893,N_1653);
or U2509 (N_2509,N_1282,N_1782);
and U2510 (N_2510,N_1744,N_1055);
xor U2511 (N_2511,N_1505,N_1083);
nand U2512 (N_2512,N_1519,N_1601);
or U2513 (N_2513,N_1867,N_1074);
nand U2514 (N_2514,N_1989,N_1489);
nand U2515 (N_2515,N_1855,N_1659);
and U2516 (N_2516,N_1442,N_1689);
nand U2517 (N_2517,N_1744,N_1544);
or U2518 (N_2518,N_1385,N_1216);
nand U2519 (N_2519,N_1314,N_1036);
xor U2520 (N_2520,N_1884,N_1166);
and U2521 (N_2521,N_1833,N_1920);
xor U2522 (N_2522,N_1927,N_1654);
or U2523 (N_2523,N_1422,N_1591);
and U2524 (N_2524,N_1244,N_1669);
nor U2525 (N_2525,N_1109,N_1276);
or U2526 (N_2526,N_1322,N_1899);
nand U2527 (N_2527,N_1923,N_1648);
and U2528 (N_2528,N_1269,N_1475);
xor U2529 (N_2529,N_1867,N_1700);
nand U2530 (N_2530,N_1522,N_1651);
nand U2531 (N_2531,N_1428,N_1288);
and U2532 (N_2532,N_1086,N_1071);
xor U2533 (N_2533,N_1376,N_1573);
or U2534 (N_2534,N_1625,N_1621);
or U2535 (N_2535,N_1111,N_1536);
nor U2536 (N_2536,N_1781,N_1147);
nor U2537 (N_2537,N_1099,N_1393);
xor U2538 (N_2538,N_1725,N_1743);
or U2539 (N_2539,N_1730,N_1622);
or U2540 (N_2540,N_1971,N_1144);
or U2541 (N_2541,N_1182,N_1980);
nor U2542 (N_2542,N_1056,N_1370);
xor U2543 (N_2543,N_1587,N_1136);
nor U2544 (N_2544,N_1948,N_1029);
nand U2545 (N_2545,N_1402,N_1059);
nor U2546 (N_2546,N_1394,N_1120);
xnor U2547 (N_2547,N_1471,N_1943);
and U2548 (N_2548,N_1496,N_1436);
nand U2549 (N_2549,N_1915,N_1898);
and U2550 (N_2550,N_1490,N_1097);
xor U2551 (N_2551,N_1641,N_1592);
or U2552 (N_2552,N_1624,N_1481);
xor U2553 (N_2553,N_1135,N_1972);
xor U2554 (N_2554,N_1101,N_1111);
nor U2555 (N_2555,N_1056,N_1395);
nor U2556 (N_2556,N_1638,N_1409);
or U2557 (N_2557,N_1182,N_1874);
and U2558 (N_2558,N_1049,N_1088);
nand U2559 (N_2559,N_1102,N_1507);
nand U2560 (N_2560,N_1270,N_1875);
nand U2561 (N_2561,N_1874,N_1927);
or U2562 (N_2562,N_1222,N_1016);
and U2563 (N_2563,N_1022,N_1748);
or U2564 (N_2564,N_1838,N_1104);
xor U2565 (N_2565,N_1636,N_1305);
xor U2566 (N_2566,N_1637,N_1856);
nand U2567 (N_2567,N_1462,N_1294);
nor U2568 (N_2568,N_1583,N_1333);
nor U2569 (N_2569,N_1733,N_1203);
and U2570 (N_2570,N_1145,N_1808);
nand U2571 (N_2571,N_1027,N_1431);
nor U2572 (N_2572,N_1227,N_1204);
xnor U2573 (N_2573,N_1152,N_1500);
nor U2574 (N_2574,N_1520,N_1151);
and U2575 (N_2575,N_1505,N_1006);
nor U2576 (N_2576,N_1486,N_1206);
nor U2577 (N_2577,N_1394,N_1699);
nor U2578 (N_2578,N_1162,N_1977);
nor U2579 (N_2579,N_1053,N_1522);
or U2580 (N_2580,N_1463,N_1442);
nand U2581 (N_2581,N_1541,N_1837);
xnor U2582 (N_2582,N_1731,N_1164);
nand U2583 (N_2583,N_1979,N_1559);
nor U2584 (N_2584,N_1984,N_1753);
and U2585 (N_2585,N_1649,N_1043);
and U2586 (N_2586,N_1087,N_1067);
nand U2587 (N_2587,N_1218,N_1867);
or U2588 (N_2588,N_1761,N_1833);
nand U2589 (N_2589,N_1702,N_1686);
xnor U2590 (N_2590,N_1638,N_1985);
nor U2591 (N_2591,N_1893,N_1746);
nor U2592 (N_2592,N_1939,N_1977);
nand U2593 (N_2593,N_1097,N_1926);
or U2594 (N_2594,N_1869,N_1478);
xnor U2595 (N_2595,N_1813,N_1399);
nand U2596 (N_2596,N_1178,N_1666);
xnor U2597 (N_2597,N_1722,N_1140);
nand U2598 (N_2598,N_1344,N_1626);
or U2599 (N_2599,N_1386,N_1423);
nand U2600 (N_2600,N_1509,N_1739);
xnor U2601 (N_2601,N_1744,N_1184);
and U2602 (N_2602,N_1846,N_1689);
xnor U2603 (N_2603,N_1012,N_1872);
nand U2604 (N_2604,N_1236,N_1234);
or U2605 (N_2605,N_1771,N_1591);
nor U2606 (N_2606,N_1604,N_1311);
nor U2607 (N_2607,N_1374,N_1396);
nor U2608 (N_2608,N_1000,N_1279);
nand U2609 (N_2609,N_1029,N_1166);
and U2610 (N_2610,N_1928,N_1905);
nand U2611 (N_2611,N_1798,N_1302);
nand U2612 (N_2612,N_1215,N_1267);
and U2613 (N_2613,N_1264,N_1857);
and U2614 (N_2614,N_1870,N_1517);
and U2615 (N_2615,N_1959,N_1160);
or U2616 (N_2616,N_1669,N_1784);
xor U2617 (N_2617,N_1960,N_1710);
nand U2618 (N_2618,N_1268,N_1221);
nor U2619 (N_2619,N_1497,N_1505);
xor U2620 (N_2620,N_1827,N_1334);
xnor U2621 (N_2621,N_1803,N_1387);
or U2622 (N_2622,N_1216,N_1708);
nand U2623 (N_2623,N_1528,N_1096);
xor U2624 (N_2624,N_1766,N_1191);
nand U2625 (N_2625,N_1892,N_1063);
nand U2626 (N_2626,N_1566,N_1045);
xor U2627 (N_2627,N_1278,N_1377);
or U2628 (N_2628,N_1389,N_1066);
nor U2629 (N_2629,N_1571,N_1380);
nor U2630 (N_2630,N_1222,N_1057);
nor U2631 (N_2631,N_1020,N_1752);
and U2632 (N_2632,N_1531,N_1775);
xnor U2633 (N_2633,N_1023,N_1667);
xnor U2634 (N_2634,N_1224,N_1298);
xnor U2635 (N_2635,N_1796,N_1433);
nand U2636 (N_2636,N_1971,N_1238);
nand U2637 (N_2637,N_1893,N_1894);
and U2638 (N_2638,N_1992,N_1134);
xor U2639 (N_2639,N_1635,N_1509);
nor U2640 (N_2640,N_1073,N_1017);
or U2641 (N_2641,N_1754,N_1059);
nor U2642 (N_2642,N_1713,N_1205);
nand U2643 (N_2643,N_1289,N_1317);
or U2644 (N_2644,N_1965,N_1998);
and U2645 (N_2645,N_1019,N_1134);
or U2646 (N_2646,N_1462,N_1892);
nand U2647 (N_2647,N_1993,N_1392);
or U2648 (N_2648,N_1318,N_1358);
xor U2649 (N_2649,N_1114,N_1849);
and U2650 (N_2650,N_1076,N_1419);
nor U2651 (N_2651,N_1883,N_1143);
nor U2652 (N_2652,N_1708,N_1189);
or U2653 (N_2653,N_1611,N_1357);
nand U2654 (N_2654,N_1545,N_1739);
or U2655 (N_2655,N_1215,N_1037);
and U2656 (N_2656,N_1778,N_1636);
or U2657 (N_2657,N_1866,N_1554);
xnor U2658 (N_2658,N_1288,N_1084);
nand U2659 (N_2659,N_1311,N_1615);
nor U2660 (N_2660,N_1725,N_1405);
xor U2661 (N_2661,N_1034,N_1020);
nor U2662 (N_2662,N_1748,N_1211);
xor U2663 (N_2663,N_1666,N_1366);
nand U2664 (N_2664,N_1637,N_1158);
and U2665 (N_2665,N_1085,N_1297);
nor U2666 (N_2666,N_1343,N_1164);
and U2667 (N_2667,N_1636,N_1566);
nor U2668 (N_2668,N_1864,N_1388);
nor U2669 (N_2669,N_1148,N_1316);
xnor U2670 (N_2670,N_1537,N_1913);
nand U2671 (N_2671,N_1520,N_1830);
nand U2672 (N_2672,N_1041,N_1722);
nand U2673 (N_2673,N_1244,N_1867);
xnor U2674 (N_2674,N_1941,N_1014);
nor U2675 (N_2675,N_1429,N_1884);
nor U2676 (N_2676,N_1820,N_1545);
nor U2677 (N_2677,N_1876,N_1808);
xor U2678 (N_2678,N_1271,N_1458);
nand U2679 (N_2679,N_1233,N_1008);
and U2680 (N_2680,N_1582,N_1397);
nand U2681 (N_2681,N_1935,N_1986);
nor U2682 (N_2682,N_1591,N_1440);
and U2683 (N_2683,N_1593,N_1641);
xor U2684 (N_2684,N_1456,N_1191);
nor U2685 (N_2685,N_1120,N_1091);
and U2686 (N_2686,N_1326,N_1370);
nand U2687 (N_2687,N_1135,N_1999);
nand U2688 (N_2688,N_1805,N_1385);
and U2689 (N_2689,N_1229,N_1759);
and U2690 (N_2690,N_1927,N_1326);
nor U2691 (N_2691,N_1090,N_1913);
nor U2692 (N_2692,N_1226,N_1038);
nand U2693 (N_2693,N_1716,N_1616);
nand U2694 (N_2694,N_1304,N_1275);
or U2695 (N_2695,N_1541,N_1638);
nor U2696 (N_2696,N_1043,N_1470);
nor U2697 (N_2697,N_1330,N_1004);
nor U2698 (N_2698,N_1149,N_1441);
nand U2699 (N_2699,N_1987,N_1834);
xor U2700 (N_2700,N_1201,N_1906);
and U2701 (N_2701,N_1259,N_1091);
or U2702 (N_2702,N_1798,N_1905);
or U2703 (N_2703,N_1060,N_1884);
and U2704 (N_2704,N_1681,N_1235);
and U2705 (N_2705,N_1970,N_1395);
nor U2706 (N_2706,N_1996,N_1947);
or U2707 (N_2707,N_1724,N_1884);
nor U2708 (N_2708,N_1011,N_1507);
xor U2709 (N_2709,N_1043,N_1945);
nor U2710 (N_2710,N_1796,N_1898);
xor U2711 (N_2711,N_1742,N_1714);
nor U2712 (N_2712,N_1137,N_1227);
or U2713 (N_2713,N_1393,N_1086);
or U2714 (N_2714,N_1932,N_1943);
or U2715 (N_2715,N_1131,N_1439);
nand U2716 (N_2716,N_1458,N_1744);
nand U2717 (N_2717,N_1346,N_1982);
or U2718 (N_2718,N_1271,N_1980);
and U2719 (N_2719,N_1833,N_1112);
nor U2720 (N_2720,N_1043,N_1398);
xor U2721 (N_2721,N_1809,N_1975);
nor U2722 (N_2722,N_1332,N_1916);
or U2723 (N_2723,N_1749,N_1717);
and U2724 (N_2724,N_1135,N_1043);
nor U2725 (N_2725,N_1645,N_1123);
and U2726 (N_2726,N_1561,N_1798);
nand U2727 (N_2727,N_1589,N_1968);
xnor U2728 (N_2728,N_1367,N_1580);
xor U2729 (N_2729,N_1123,N_1001);
nand U2730 (N_2730,N_1880,N_1574);
nor U2731 (N_2731,N_1839,N_1493);
nand U2732 (N_2732,N_1954,N_1985);
or U2733 (N_2733,N_1073,N_1512);
nor U2734 (N_2734,N_1727,N_1511);
or U2735 (N_2735,N_1245,N_1386);
or U2736 (N_2736,N_1849,N_1171);
xor U2737 (N_2737,N_1490,N_1818);
nand U2738 (N_2738,N_1560,N_1216);
nand U2739 (N_2739,N_1598,N_1544);
xor U2740 (N_2740,N_1887,N_1326);
xor U2741 (N_2741,N_1203,N_1056);
nor U2742 (N_2742,N_1710,N_1215);
nor U2743 (N_2743,N_1390,N_1169);
and U2744 (N_2744,N_1609,N_1782);
nor U2745 (N_2745,N_1025,N_1950);
nand U2746 (N_2746,N_1321,N_1109);
and U2747 (N_2747,N_1934,N_1084);
xnor U2748 (N_2748,N_1313,N_1252);
xnor U2749 (N_2749,N_1343,N_1956);
nor U2750 (N_2750,N_1685,N_1582);
or U2751 (N_2751,N_1595,N_1220);
and U2752 (N_2752,N_1638,N_1702);
nand U2753 (N_2753,N_1550,N_1087);
nor U2754 (N_2754,N_1387,N_1961);
xor U2755 (N_2755,N_1162,N_1057);
nand U2756 (N_2756,N_1942,N_1748);
xnor U2757 (N_2757,N_1222,N_1845);
nor U2758 (N_2758,N_1199,N_1770);
xnor U2759 (N_2759,N_1074,N_1741);
or U2760 (N_2760,N_1125,N_1009);
nand U2761 (N_2761,N_1922,N_1313);
xnor U2762 (N_2762,N_1044,N_1443);
nor U2763 (N_2763,N_1445,N_1693);
nand U2764 (N_2764,N_1746,N_1391);
nand U2765 (N_2765,N_1018,N_1215);
xor U2766 (N_2766,N_1151,N_1941);
xnor U2767 (N_2767,N_1692,N_1705);
nor U2768 (N_2768,N_1368,N_1904);
nand U2769 (N_2769,N_1303,N_1489);
nand U2770 (N_2770,N_1621,N_1927);
and U2771 (N_2771,N_1280,N_1997);
or U2772 (N_2772,N_1379,N_1817);
nand U2773 (N_2773,N_1503,N_1903);
nor U2774 (N_2774,N_1030,N_1674);
xor U2775 (N_2775,N_1602,N_1706);
and U2776 (N_2776,N_1791,N_1915);
nor U2777 (N_2777,N_1389,N_1406);
nor U2778 (N_2778,N_1677,N_1539);
nand U2779 (N_2779,N_1692,N_1019);
or U2780 (N_2780,N_1728,N_1093);
or U2781 (N_2781,N_1375,N_1779);
or U2782 (N_2782,N_1601,N_1716);
nand U2783 (N_2783,N_1617,N_1868);
xor U2784 (N_2784,N_1954,N_1020);
or U2785 (N_2785,N_1126,N_1297);
or U2786 (N_2786,N_1003,N_1791);
nand U2787 (N_2787,N_1879,N_1031);
and U2788 (N_2788,N_1294,N_1160);
nand U2789 (N_2789,N_1116,N_1045);
and U2790 (N_2790,N_1396,N_1871);
nand U2791 (N_2791,N_1033,N_1354);
or U2792 (N_2792,N_1799,N_1934);
and U2793 (N_2793,N_1806,N_1049);
nand U2794 (N_2794,N_1730,N_1230);
nand U2795 (N_2795,N_1981,N_1680);
or U2796 (N_2796,N_1753,N_1152);
or U2797 (N_2797,N_1457,N_1056);
nand U2798 (N_2798,N_1112,N_1061);
and U2799 (N_2799,N_1814,N_1348);
or U2800 (N_2800,N_1406,N_1107);
xor U2801 (N_2801,N_1076,N_1933);
or U2802 (N_2802,N_1184,N_1953);
nand U2803 (N_2803,N_1740,N_1786);
xor U2804 (N_2804,N_1288,N_1101);
nand U2805 (N_2805,N_1547,N_1747);
nor U2806 (N_2806,N_1395,N_1154);
or U2807 (N_2807,N_1869,N_1879);
nand U2808 (N_2808,N_1945,N_1907);
xnor U2809 (N_2809,N_1479,N_1500);
or U2810 (N_2810,N_1317,N_1550);
or U2811 (N_2811,N_1391,N_1413);
or U2812 (N_2812,N_1775,N_1652);
nor U2813 (N_2813,N_1546,N_1928);
or U2814 (N_2814,N_1939,N_1029);
xnor U2815 (N_2815,N_1723,N_1510);
nor U2816 (N_2816,N_1302,N_1230);
xor U2817 (N_2817,N_1417,N_1321);
nand U2818 (N_2818,N_1491,N_1564);
or U2819 (N_2819,N_1270,N_1822);
nand U2820 (N_2820,N_1792,N_1327);
and U2821 (N_2821,N_1339,N_1764);
and U2822 (N_2822,N_1291,N_1880);
xnor U2823 (N_2823,N_1833,N_1250);
nand U2824 (N_2824,N_1438,N_1032);
and U2825 (N_2825,N_1852,N_1531);
and U2826 (N_2826,N_1992,N_1074);
xor U2827 (N_2827,N_1175,N_1127);
nand U2828 (N_2828,N_1048,N_1777);
xnor U2829 (N_2829,N_1999,N_1664);
and U2830 (N_2830,N_1723,N_1475);
and U2831 (N_2831,N_1949,N_1936);
and U2832 (N_2832,N_1262,N_1821);
nor U2833 (N_2833,N_1679,N_1190);
and U2834 (N_2834,N_1519,N_1457);
nand U2835 (N_2835,N_1723,N_1436);
or U2836 (N_2836,N_1437,N_1567);
and U2837 (N_2837,N_1830,N_1701);
nand U2838 (N_2838,N_1956,N_1124);
nor U2839 (N_2839,N_1257,N_1957);
or U2840 (N_2840,N_1536,N_1911);
or U2841 (N_2841,N_1590,N_1496);
or U2842 (N_2842,N_1267,N_1210);
nand U2843 (N_2843,N_1141,N_1184);
or U2844 (N_2844,N_1799,N_1059);
or U2845 (N_2845,N_1830,N_1206);
nor U2846 (N_2846,N_1323,N_1269);
or U2847 (N_2847,N_1129,N_1131);
nor U2848 (N_2848,N_1884,N_1818);
xor U2849 (N_2849,N_1340,N_1291);
nor U2850 (N_2850,N_1831,N_1889);
and U2851 (N_2851,N_1651,N_1513);
nand U2852 (N_2852,N_1270,N_1372);
and U2853 (N_2853,N_1905,N_1384);
nor U2854 (N_2854,N_1981,N_1907);
nor U2855 (N_2855,N_1639,N_1325);
xnor U2856 (N_2856,N_1363,N_1961);
nand U2857 (N_2857,N_1585,N_1945);
or U2858 (N_2858,N_1088,N_1454);
xnor U2859 (N_2859,N_1900,N_1936);
nor U2860 (N_2860,N_1442,N_1924);
or U2861 (N_2861,N_1963,N_1065);
nor U2862 (N_2862,N_1108,N_1334);
nor U2863 (N_2863,N_1919,N_1511);
nor U2864 (N_2864,N_1884,N_1510);
nor U2865 (N_2865,N_1361,N_1975);
xnor U2866 (N_2866,N_1906,N_1729);
and U2867 (N_2867,N_1286,N_1058);
xnor U2868 (N_2868,N_1460,N_1147);
and U2869 (N_2869,N_1970,N_1872);
xor U2870 (N_2870,N_1844,N_1747);
and U2871 (N_2871,N_1505,N_1709);
nor U2872 (N_2872,N_1018,N_1290);
nand U2873 (N_2873,N_1696,N_1264);
xor U2874 (N_2874,N_1651,N_1207);
nand U2875 (N_2875,N_1476,N_1355);
nor U2876 (N_2876,N_1841,N_1949);
or U2877 (N_2877,N_1556,N_1574);
and U2878 (N_2878,N_1949,N_1114);
and U2879 (N_2879,N_1736,N_1628);
or U2880 (N_2880,N_1812,N_1329);
nor U2881 (N_2881,N_1766,N_1916);
nand U2882 (N_2882,N_1284,N_1415);
xor U2883 (N_2883,N_1283,N_1588);
xor U2884 (N_2884,N_1592,N_1360);
and U2885 (N_2885,N_1366,N_1628);
nand U2886 (N_2886,N_1236,N_1603);
nor U2887 (N_2887,N_1632,N_1943);
nand U2888 (N_2888,N_1080,N_1367);
nor U2889 (N_2889,N_1000,N_1523);
xor U2890 (N_2890,N_1895,N_1339);
xnor U2891 (N_2891,N_1407,N_1816);
xnor U2892 (N_2892,N_1504,N_1290);
nand U2893 (N_2893,N_1419,N_1630);
xor U2894 (N_2894,N_1542,N_1873);
and U2895 (N_2895,N_1853,N_1157);
and U2896 (N_2896,N_1963,N_1908);
nor U2897 (N_2897,N_1370,N_1721);
and U2898 (N_2898,N_1679,N_1328);
or U2899 (N_2899,N_1870,N_1554);
nand U2900 (N_2900,N_1342,N_1196);
or U2901 (N_2901,N_1382,N_1231);
nand U2902 (N_2902,N_1524,N_1717);
xnor U2903 (N_2903,N_1319,N_1267);
nand U2904 (N_2904,N_1715,N_1565);
and U2905 (N_2905,N_1752,N_1411);
nand U2906 (N_2906,N_1162,N_1803);
or U2907 (N_2907,N_1724,N_1002);
or U2908 (N_2908,N_1094,N_1370);
nor U2909 (N_2909,N_1311,N_1487);
and U2910 (N_2910,N_1945,N_1354);
nor U2911 (N_2911,N_1972,N_1787);
and U2912 (N_2912,N_1945,N_1370);
nor U2913 (N_2913,N_1409,N_1091);
and U2914 (N_2914,N_1853,N_1138);
and U2915 (N_2915,N_1718,N_1370);
or U2916 (N_2916,N_1735,N_1986);
nor U2917 (N_2917,N_1368,N_1676);
and U2918 (N_2918,N_1757,N_1257);
or U2919 (N_2919,N_1031,N_1488);
and U2920 (N_2920,N_1157,N_1610);
or U2921 (N_2921,N_1687,N_1632);
nor U2922 (N_2922,N_1181,N_1453);
nand U2923 (N_2923,N_1101,N_1409);
xor U2924 (N_2924,N_1790,N_1014);
nand U2925 (N_2925,N_1076,N_1724);
nand U2926 (N_2926,N_1782,N_1621);
or U2927 (N_2927,N_1130,N_1620);
or U2928 (N_2928,N_1172,N_1085);
and U2929 (N_2929,N_1444,N_1324);
nand U2930 (N_2930,N_1420,N_1747);
nor U2931 (N_2931,N_1811,N_1278);
nand U2932 (N_2932,N_1332,N_1406);
xnor U2933 (N_2933,N_1764,N_1654);
xnor U2934 (N_2934,N_1145,N_1764);
and U2935 (N_2935,N_1127,N_1818);
and U2936 (N_2936,N_1670,N_1285);
xor U2937 (N_2937,N_1306,N_1786);
and U2938 (N_2938,N_1733,N_1483);
xnor U2939 (N_2939,N_1136,N_1383);
nand U2940 (N_2940,N_1099,N_1139);
xor U2941 (N_2941,N_1766,N_1385);
nand U2942 (N_2942,N_1925,N_1619);
nand U2943 (N_2943,N_1760,N_1570);
nor U2944 (N_2944,N_1393,N_1439);
and U2945 (N_2945,N_1704,N_1201);
xnor U2946 (N_2946,N_1708,N_1336);
xor U2947 (N_2947,N_1268,N_1891);
and U2948 (N_2948,N_1383,N_1478);
nand U2949 (N_2949,N_1564,N_1868);
or U2950 (N_2950,N_1177,N_1537);
or U2951 (N_2951,N_1114,N_1751);
and U2952 (N_2952,N_1335,N_1079);
or U2953 (N_2953,N_1933,N_1902);
nor U2954 (N_2954,N_1957,N_1414);
xor U2955 (N_2955,N_1241,N_1001);
or U2956 (N_2956,N_1632,N_1261);
nand U2957 (N_2957,N_1318,N_1644);
or U2958 (N_2958,N_1746,N_1244);
and U2959 (N_2959,N_1672,N_1310);
nand U2960 (N_2960,N_1043,N_1205);
nand U2961 (N_2961,N_1356,N_1964);
or U2962 (N_2962,N_1740,N_1047);
xor U2963 (N_2963,N_1551,N_1419);
nor U2964 (N_2964,N_1744,N_1767);
nor U2965 (N_2965,N_1541,N_1862);
nand U2966 (N_2966,N_1659,N_1082);
nor U2967 (N_2967,N_1678,N_1298);
and U2968 (N_2968,N_1471,N_1843);
and U2969 (N_2969,N_1293,N_1334);
xor U2970 (N_2970,N_1207,N_1196);
xnor U2971 (N_2971,N_1179,N_1291);
and U2972 (N_2972,N_1866,N_1113);
xor U2973 (N_2973,N_1955,N_1108);
nand U2974 (N_2974,N_1002,N_1864);
nand U2975 (N_2975,N_1465,N_1855);
and U2976 (N_2976,N_1235,N_1429);
nand U2977 (N_2977,N_1478,N_1075);
xnor U2978 (N_2978,N_1553,N_1860);
and U2979 (N_2979,N_1294,N_1834);
and U2980 (N_2980,N_1776,N_1215);
nand U2981 (N_2981,N_1406,N_1737);
xor U2982 (N_2982,N_1786,N_1612);
xor U2983 (N_2983,N_1991,N_1412);
nor U2984 (N_2984,N_1115,N_1356);
xnor U2985 (N_2985,N_1199,N_1016);
or U2986 (N_2986,N_1784,N_1859);
nand U2987 (N_2987,N_1951,N_1746);
nor U2988 (N_2988,N_1789,N_1185);
and U2989 (N_2989,N_1009,N_1184);
nand U2990 (N_2990,N_1969,N_1488);
xnor U2991 (N_2991,N_1702,N_1206);
nand U2992 (N_2992,N_1230,N_1324);
and U2993 (N_2993,N_1021,N_1471);
xnor U2994 (N_2994,N_1770,N_1782);
nor U2995 (N_2995,N_1068,N_1586);
and U2996 (N_2996,N_1642,N_1309);
or U2997 (N_2997,N_1828,N_1697);
and U2998 (N_2998,N_1988,N_1104);
or U2999 (N_2999,N_1042,N_1072);
xor U3000 (N_3000,N_2458,N_2519);
or U3001 (N_3001,N_2858,N_2233);
nand U3002 (N_3002,N_2943,N_2487);
nand U3003 (N_3003,N_2777,N_2823);
xnor U3004 (N_3004,N_2963,N_2450);
nand U3005 (N_3005,N_2689,N_2786);
nand U3006 (N_3006,N_2043,N_2162);
nor U3007 (N_3007,N_2948,N_2238);
xnor U3008 (N_3008,N_2835,N_2330);
nand U3009 (N_3009,N_2815,N_2701);
or U3010 (N_3010,N_2505,N_2181);
and U3011 (N_3011,N_2308,N_2876);
or U3012 (N_3012,N_2604,N_2580);
or U3013 (N_3013,N_2406,N_2925);
or U3014 (N_3014,N_2376,N_2237);
xnor U3015 (N_3015,N_2543,N_2071);
nand U3016 (N_3016,N_2540,N_2704);
nand U3017 (N_3017,N_2561,N_2537);
or U3018 (N_3018,N_2807,N_2620);
nor U3019 (N_3019,N_2502,N_2816);
xor U3020 (N_3020,N_2247,N_2562);
or U3021 (N_3021,N_2437,N_2080);
xor U3022 (N_3022,N_2892,N_2365);
nor U3023 (N_3023,N_2426,N_2115);
and U3024 (N_3024,N_2705,N_2186);
or U3025 (N_3025,N_2433,N_2718);
and U3026 (N_3026,N_2479,N_2851);
or U3027 (N_3027,N_2837,N_2668);
and U3028 (N_3028,N_2574,N_2964);
nor U3029 (N_3029,N_2383,N_2163);
xnor U3030 (N_3030,N_2370,N_2098);
nor U3031 (N_3031,N_2530,N_2239);
and U3032 (N_3032,N_2885,N_2691);
xnor U3033 (N_3033,N_2926,N_2256);
nor U3034 (N_3034,N_2398,N_2386);
nor U3035 (N_3035,N_2494,N_2980);
nand U3036 (N_3036,N_2898,N_2659);
and U3037 (N_3037,N_2297,N_2836);
nand U3038 (N_3038,N_2860,N_2595);
nor U3039 (N_3039,N_2912,N_2687);
xnor U3040 (N_3040,N_2766,N_2351);
nor U3041 (N_3041,N_2000,N_2552);
or U3042 (N_3042,N_2591,N_2294);
or U3043 (N_3043,N_2920,N_2944);
nand U3044 (N_3044,N_2734,N_2024);
and U3045 (N_3045,N_2295,N_2198);
xnor U3046 (N_3046,N_2594,N_2063);
xor U3047 (N_3047,N_2189,N_2306);
nor U3048 (N_3048,N_2439,N_2656);
or U3049 (N_3049,N_2817,N_2371);
and U3050 (N_3050,N_2125,N_2628);
and U3051 (N_3051,N_2087,N_2631);
xnor U3052 (N_3052,N_2206,N_2831);
xor U3053 (N_3053,N_2970,N_2464);
nand U3054 (N_3054,N_2467,N_2062);
nand U3055 (N_3055,N_2870,N_2289);
or U3056 (N_3056,N_2958,N_2429);
and U3057 (N_3057,N_2379,N_2723);
nor U3058 (N_3058,N_2217,N_2149);
and U3059 (N_3059,N_2548,N_2966);
xnor U3060 (N_3060,N_2515,N_2418);
or U3061 (N_3061,N_2927,N_2449);
xnor U3062 (N_3062,N_2410,N_2536);
xor U3063 (N_3063,N_2269,N_2216);
xor U3064 (N_3064,N_2446,N_2753);
nand U3065 (N_3065,N_2324,N_2174);
and U3066 (N_3066,N_2250,N_2385);
nand U3067 (N_3067,N_2872,N_2973);
or U3068 (N_3068,N_2647,N_2378);
nor U3069 (N_3069,N_2034,N_2882);
nand U3070 (N_3070,N_2696,N_2585);
and U3071 (N_3071,N_2048,N_2147);
xnor U3072 (N_3072,N_2611,N_2353);
or U3073 (N_3073,N_2188,N_2278);
and U3074 (N_3074,N_2928,N_2259);
nor U3075 (N_3075,N_2806,N_2660);
xnor U3076 (N_3076,N_2171,N_2305);
nand U3077 (N_3077,N_2771,N_2686);
and U3078 (N_3078,N_2751,N_2599);
or U3079 (N_3079,N_2785,N_2824);
xor U3080 (N_3080,N_2945,N_2225);
nand U3081 (N_3081,N_2669,N_2682);
nor U3082 (N_3082,N_2972,N_2867);
or U3083 (N_3083,N_2531,N_2018);
nand U3084 (N_3084,N_2637,N_2170);
and U3085 (N_3085,N_2922,N_2135);
and U3086 (N_3086,N_2729,N_2626);
nor U3087 (N_3087,N_2110,N_2275);
xor U3088 (N_3088,N_2648,N_2150);
xor U3089 (N_3089,N_2005,N_2372);
nor U3090 (N_3090,N_2608,N_2903);
nor U3091 (N_3091,N_2838,N_2231);
xor U3092 (N_3092,N_2445,N_2169);
nor U3093 (N_3093,N_2442,N_2456);
nor U3094 (N_3094,N_2588,N_2763);
or U3095 (N_3095,N_2347,N_2553);
xor U3096 (N_3096,N_2214,N_2857);
nor U3097 (N_3097,N_2544,N_2525);
or U3098 (N_3098,N_2335,N_2740);
and U3099 (N_3099,N_2513,N_2451);
or U3100 (N_3100,N_2025,N_2008);
and U3101 (N_3101,N_2440,N_2953);
nand U3102 (N_3102,N_2469,N_2853);
xnor U3103 (N_3103,N_2360,N_2829);
xnor U3104 (N_3104,N_2855,N_2050);
xor U3105 (N_3105,N_2127,N_2760);
nor U3106 (N_3106,N_2232,N_2055);
and U3107 (N_3107,N_2399,N_2327);
and U3108 (N_3108,N_2597,N_2322);
and U3109 (N_3109,N_2741,N_2182);
or U3110 (N_3110,N_2719,N_2253);
xor U3111 (N_3111,N_2340,N_2567);
nor U3112 (N_3112,N_2454,N_2218);
nor U3113 (N_3113,N_2605,N_2013);
and U3114 (N_3114,N_2747,N_2804);
nand U3115 (N_3115,N_2263,N_2489);
nand U3116 (N_3116,N_2998,N_2971);
or U3117 (N_3117,N_2276,N_2821);
nor U3118 (N_3118,N_2653,N_2550);
or U3119 (N_3119,N_2713,N_2685);
and U3120 (N_3120,N_2392,N_2140);
nor U3121 (N_3121,N_2332,N_2508);
xnor U3122 (N_3122,N_2600,N_2665);
xor U3123 (N_3123,N_2257,N_2711);
or U3124 (N_3124,N_2354,N_2714);
and U3125 (N_3125,N_2077,N_2795);
xor U3126 (N_3126,N_2623,N_2158);
nor U3127 (N_3127,N_2678,N_2731);
and U3128 (N_3128,N_2111,N_2681);
nor U3129 (N_3129,N_2148,N_2888);
nor U3130 (N_3130,N_2936,N_2046);
and U3131 (N_3131,N_2905,N_2296);
nor U3132 (N_3132,N_2667,N_2862);
nor U3133 (N_3133,N_2160,N_2066);
nand U3134 (N_3134,N_2547,N_2315);
or U3135 (N_3135,N_2987,N_2526);
nand U3136 (N_3136,N_2044,N_2880);
nand U3137 (N_3137,N_2030,N_2907);
nand U3138 (N_3138,N_2377,N_2956);
xnor U3139 (N_3139,N_2828,N_2997);
and U3140 (N_3140,N_2655,N_2509);
nand U3141 (N_3141,N_2798,N_2106);
nor U3142 (N_3142,N_2323,N_2617);
or U3143 (N_3143,N_2221,N_2921);
nand U3144 (N_3144,N_2395,N_2792);
xnor U3145 (N_3145,N_2499,N_2841);
nand U3146 (N_3146,N_2251,N_2664);
nand U3147 (N_3147,N_2675,N_2299);
and U3148 (N_3148,N_2176,N_2028);
or U3149 (N_3149,N_2116,N_2725);
nand U3150 (N_3150,N_2493,N_2707);
nor U3151 (N_3151,N_2465,N_2739);
xor U3152 (N_3152,N_2461,N_2863);
or U3153 (N_3153,N_2443,N_2274);
xnor U3154 (N_3154,N_2281,N_2690);
and U3155 (N_3155,N_2428,N_2783);
or U3156 (N_3156,N_2721,N_2425);
xor U3157 (N_3157,N_2624,N_2965);
xor U3158 (N_3158,N_2931,N_2390);
nor U3159 (N_3159,N_2078,N_2284);
xnor U3160 (N_3160,N_2645,N_2706);
nand U3161 (N_3161,N_2015,N_2897);
or U3162 (N_3162,N_2503,N_2033);
or U3163 (N_3163,N_2640,N_2618);
nand U3164 (N_3164,N_2038,N_2568);
nor U3165 (N_3165,N_2118,N_2932);
and U3166 (N_3166,N_2962,N_2343);
nor U3167 (N_3167,N_2615,N_2081);
and U3168 (N_3168,N_2128,N_2420);
xnor U3169 (N_3169,N_2243,N_2144);
or U3170 (N_3170,N_2758,N_2727);
or U3171 (N_3171,N_2448,N_2325);
nand U3172 (N_3172,N_2844,N_2268);
xnor U3173 (N_3173,N_2344,N_2213);
nor U3174 (N_3174,N_2491,N_2381);
or U3175 (N_3175,N_2840,N_2793);
nand U3176 (N_3176,N_2934,N_2812);
xnor U3177 (N_3177,N_2180,N_2722);
or U3178 (N_3178,N_2400,N_2004);
and U3179 (N_3179,N_2782,N_2363);
xor U3180 (N_3180,N_2569,N_2396);
xnor U3181 (N_3181,N_2166,N_2416);
nand U3182 (N_3182,N_2389,N_2133);
nand U3183 (N_3183,N_2661,N_2303);
nand U3184 (N_3184,N_2463,N_2167);
or U3185 (N_3185,N_2930,N_2079);
nand U3186 (N_3186,N_2603,N_2288);
xor U3187 (N_3187,N_2053,N_2610);
nand U3188 (N_3188,N_2107,N_2658);
xnor U3189 (N_3189,N_2680,N_2036);
xor U3190 (N_3190,N_2146,N_2411);
or U3191 (N_3191,N_2103,N_2510);
xnor U3192 (N_3192,N_2279,N_2674);
nand U3193 (N_3193,N_2843,N_2468);
or U3194 (N_3194,N_2693,N_2482);
nand U3195 (N_3195,N_2156,N_2616);
and U3196 (N_3196,N_2177,N_2878);
nor U3197 (N_3197,N_2310,N_2480);
nor U3198 (N_3198,N_2999,N_2151);
nor U3199 (N_3199,N_2326,N_2141);
nand U3200 (N_3200,N_2102,N_2316);
xnor U3201 (N_3201,N_2412,N_2991);
or U3202 (N_3202,N_2527,N_2587);
or U3203 (N_3203,N_2774,N_2096);
nor U3204 (N_3204,N_2590,N_2649);
or U3205 (N_3205,N_2496,N_2120);
nor U3206 (N_3206,N_2121,N_2803);
and U3207 (N_3207,N_2545,N_2961);
xnor U3208 (N_3208,N_2935,N_2614);
nand U3209 (N_3209,N_2780,N_2471);
xnor U3210 (N_3210,N_2336,N_2388);
nor U3211 (N_3211,N_2374,N_2357);
and U3212 (N_3212,N_2052,N_2341);
nor U3213 (N_3213,N_2134,N_2229);
nor U3214 (N_3214,N_2248,N_2300);
or U3215 (N_3215,N_2960,N_2947);
xor U3216 (N_3216,N_2775,N_2483);
and U3217 (N_3217,N_2265,N_2227);
nand U3218 (N_3218,N_2772,N_2241);
nor U3219 (N_3219,N_2498,N_2159);
xnor U3220 (N_3220,N_2799,N_2283);
nor U3221 (N_3221,N_2695,N_2466);
or U3222 (N_3222,N_2427,N_2067);
and U3223 (N_3223,N_2039,N_2684);
and U3224 (N_3224,N_2700,N_2161);
nor U3225 (N_3225,N_2114,N_2403);
or U3226 (N_3226,N_2260,N_2976);
nor U3227 (N_3227,N_2031,N_2058);
and U3228 (N_3228,N_2348,N_2254);
and U3229 (N_3229,N_2318,N_2712);
and U3230 (N_3230,N_2756,N_2040);
nor U3231 (N_3231,N_2084,N_2869);
xnor U3232 (N_3232,N_2978,N_2663);
nor U3233 (N_3233,N_2601,N_2003);
and U3234 (N_3234,N_2258,N_2549);
nand U3235 (N_3235,N_2175,N_2621);
xor U3236 (N_3236,N_2282,N_2069);
xnor U3237 (N_3237,N_2950,N_2421);
nor U3238 (N_3238,N_2773,N_2850);
xor U3239 (N_3239,N_2100,N_2195);
nor U3240 (N_3240,N_2190,N_2317);
or U3241 (N_3241,N_2082,N_2968);
nand U3242 (N_3242,N_2236,N_2994);
and U3243 (N_3243,N_2890,N_2262);
and U3244 (N_3244,N_2035,N_2800);
xnor U3245 (N_3245,N_2452,N_2313);
nor U3246 (N_3246,N_2209,N_2949);
or U3247 (N_3247,N_2811,N_2724);
xnor U3248 (N_3248,N_2635,N_2431);
or U3249 (N_3249,N_2564,N_2413);
or U3250 (N_3250,N_2524,N_2622);
nor U3251 (N_3251,N_2813,N_2632);
nor U3252 (N_3252,N_2277,N_2405);
xor U3253 (N_3253,N_2534,N_2894);
or U3254 (N_3254,N_2364,N_2809);
or U3255 (N_3255,N_2923,N_2280);
nand U3256 (N_3256,N_2022,N_2818);
nor U3257 (N_3257,N_2764,N_2027);
and U3258 (N_3258,N_2959,N_2203);
xor U3259 (N_3259,N_2345,N_2730);
or U3260 (N_3260,N_2019,N_2839);
or U3261 (N_3261,N_2650,N_2742);
and U3262 (N_3262,N_2808,N_2155);
and U3263 (N_3263,N_2520,N_2884);
nand U3264 (N_3264,N_2954,N_2387);
or U3265 (N_3265,N_2228,N_2613);
xnor U3266 (N_3266,N_2485,N_2814);
xnor U3267 (N_3267,N_2287,N_2602);
nand U3268 (N_3268,N_2293,N_2091);
nand U3269 (N_3269,N_2791,N_2652);
or U3270 (N_3270,N_2679,N_2619);
nor U3271 (N_3271,N_2021,N_2459);
nand U3272 (N_3272,N_2995,N_2132);
xor U3273 (N_3273,N_2319,N_2506);
nand U3274 (N_3274,N_2057,N_2641);
nor U3275 (N_3275,N_2767,N_2715);
and U3276 (N_3276,N_2202,N_2474);
nand U3277 (N_3277,N_2676,N_2754);
nand U3278 (N_3278,N_2745,N_2447);
xor U3279 (N_3279,N_2797,N_2165);
nor U3280 (N_3280,N_2436,N_2752);
nor U3281 (N_3281,N_2460,N_2204);
and U3282 (N_3282,N_2551,N_2886);
or U3283 (N_3283,N_2801,N_2432);
or U3284 (N_3284,N_2988,N_2009);
nor U3285 (N_3285,N_2252,N_2117);
nor U3286 (N_3286,N_2235,N_2779);
and U3287 (N_3287,N_2909,N_2919);
nor U3288 (N_3288,N_2736,N_2422);
and U3289 (N_3289,N_2255,N_2606);
xor U3290 (N_3290,N_2845,N_2511);
xnor U3291 (N_3291,N_2761,N_2023);
nor U3292 (N_3292,N_2556,N_2827);
nor U3293 (N_3293,N_2504,N_2895);
nand U3294 (N_3294,N_2220,N_2153);
xor U3295 (N_3295,N_2143,N_2402);
nand U3296 (N_3296,N_2291,N_2794);
or U3297 (N_3297,N_2952,N_2307);
and U3298 (N_3298,N_2861,N_2982);
xnor U3299 (N_3299,N_2875,N_2942);
and U3300 (N_3300,N_2933,N_2352);
xor U3301 (N_3301,N_2266,N_2735);
nand U3302 (N_3302,N_2984,N_2532);
xnor U3303 (N_3303,N_2789,N_2394);
xor U3304 (N_3304,N_2865,N_2555);
nand U3305 (N_3305,N_2369,N_2393);
nor U3306 (N_3306,N_2646,N_2271);
or U3307 (N_3307,N_2673,N_2311);
nor U3308 (N_3308,N_2638,N_2802);
xnor U3309 (N_3309,N_2967,N_2846);
xnor U3310 (N_3310,N_2554,N_2717);
nor U3311 (N_3311,N_2037,N_2085);
xnor U3312 (N_3312,N_2486,N_2191);
xor U3313 (N_3313,N_2273,N_2629);
nand U3314 (N_3314,N_2075,N_2946);
or U3315 (N_3315,N_2083,N_2901);
xnor U3316 (N_3316,N_2744,N_2002);
nand U3317 (N_3317,N_2434,N_2709);
xor U3318 (N_3318,N_2208,N_2415);
and U3319 (N_3319,N_2112,N_2157);
or U3320 (N_3320,N_2748,N_2697);
and U3321 (N_3321,N_2570,N_2993);
xor U3322 (N_3322,N_2914,N_2516);
nor U3323 (N_3323,N_2197,N_2755);
nand U3324 (N_3324,N_2732,N_2488);
or U3325 (N_3325,N_2362,N_2918);
or U3326 (N_3326,N_2879,N_2407);
xnor U3327 (N_3327,N_2331,N_2401);
nand U3328 (N_3328,N_2579,N_2196);
nand U3329 (N_3329,N_2981,N_2654);
and U3330 (N_3330,N_2762,N_2571);
and U3331 (N_3331,N_2129,N_2598);
nand U3332 (N_3332,N_2578,N_2941);
xnor U3333 (N_3333,N_2834,N_2086);
or U3334 (N_3334,N_2020,N_2910);
and U3335 (N_3335,N_2337,N_2737);
xnor U3336 (N_3336,N_2651,N_2226);
and U3337 (N_3337,N_2874,N_2832);
nand U3338 (N_3338,N_2051,N_2856);
nor U3339 (N_3339,N_2868,N_2728);
nand U3340 (N_3340,N_2951,N_2957);
nand U3341 (N_3341,N_2507,N_2924);
xor U3342 (N_3342,N_2059,N_2566);
xnor U3343 (N_3343,N_2917,N_2974);
or U3344 (N_3344,N_2887,N_2164);
xor U3345 (N_3345,N_2193,N_2788);
nor U3346 (N_3346,N_2285,N_2639);
xnor U3347 (N_3347,N_2708,N_2154);
and U3348 (N_3348,N_2969,N_2358);
xnor U3349 (N_3349,N_2738,N_2123);
xnor U3350 (N_3350,N_2359,N_2750);
nor U3351 (N_3351,N_2979,N_2430);
nand U3352 (N_3352,N_2384,N_2475);
nand U3353 (N_3353,N_2242,N_2893);
xnor U3354 (N_3354,N_2528,N_2866);
or U3355 (N_3355,N_2017,N_2350);
xnor U3356 (N_3356,N_2417,N_2007);
xnor U3357 (N_3357,N_2047,N_2261);
or U3358 (N_3358,N_2983,N_2090);
and U3359 (N_3359,N_2314,N_2136);
xnor U3360 (N_3360,N_2312,N_2996);
nor U3361 (N_3361,N_2060,N_2356);
or U3362 (N_3362,N_2557,N_2630);
nand U3363 (N_3363,N_2523,N_2877);
and U3364 (N_3364,N_2896,N_2414);
or U3365 (N_3365,N_2710,N_2184);
nand U3366 (N_3366,N_2746,N_2073);
nand U3367 (N_3367,N_2847,N_2986);
xor U3368 (N_3368,N_2938,N_2716);
nand U3369 (N_3369,N_2848,N_2940);
nand U3370 (N_3370,N_2576,N_2301);
xor U3371 (N_3371,N_2435,N_2457);
xor U3372 (N_3372,N_2219,N_2194);
xnor U3373 (N_3373,N_2726,N_2264);
or U3374 (N_3374,N_2484,N_2581);
nor U3375 (N_3375,N_2929,N_2759);
nand U3376 (N_3376,N_2346,N_2492);
nor U3377 (N_3377,N_2391,N_2230);
or U3378 (N_3378,N_2212,N_2093);
nor U3379 (N_3379,N_2224,N_2056);
and U3380 (N_3380,N_2596,N_2477);
nor U3381 (N_3381,N_2068,N_2699);
and U3382 (N_3382,N_2249,N_2329);
or U3383 (N_3383,N_2563,N_2521);
nand U3384 (N_3384,N_2992,N_2011);
xor U3385 (N_3385,N_2419,N_2852);
xnor U3386 (N_3386,N_2559,N_2881);
or U3387 (N_3387,N_2769,N_2694);
and U3388 (N_3388,N_2573,N_2683);
nand U3389 (N_3389,N_2286,N_2070);
xor U3390 (N_3390,N_2634,N_2104);
xnor U3391 (N_3391,N_2522,N_2572);
and U3392 (N_3392,N_2201,N_2309);
nand U3393 (N_3393,N_2627,N_2138);
xnor U3394 (N_3394,N_2349,N_2854);
nor U3395 (N_3395,N_2533,N_2582);
nor U3396 (N_3396,N_2272,N_2334);
or U3397 (N_3397,N_2408,N_2476);
and U3398 (N_3398,N_2560,N_2558);
nor U3399 (N_3399,N_2200,N_2733);
or U3400 (N_3400,N_2065,N_2985);
nand U3401 (N_3401,N_2500,N_2438);
nor U3402 (N_3402,N_2215,N_2382);
and U3403 (N_3403,N_2054,N_2913);
nand U3404 (N_3404,N_2178,N_2061);
nor U3405 (N_3405,N_2074,N_2207);
xor U3406 (N_3406,N_2045,N_2749);
xor U3407 (N_3407,N_2546,N_2805);
and U3408 (N_3408,N_2826,N_2472);
xor U3409 (N_3409,N_2899,N_2139);
nand U3410 (N_3410,N_2001,N_2101);
or U3411 (N_3411,N_2333,N_2302);
xnor U3412 (N_3412,N_2906,N_2172);
and U3413 (N_3413,N_2270,N_2183);
nor U3414 (N_3414,N_2320,N_2757);
xor U3415 (N_3415,N_2517,N_2240);
nor U3416 (N_3416,N_2790,N_2016);
and U3417 (N_3417,N_2478,N_2010);
or U3418 (N_3418,N_2644,N_2124);
or U3419 (N_3419,N_2677,N_2538);
and U3420 (N_3420,N_2849,N_2234);
and U3421 (N_3421,N_2088,N_2720);
xor U3422 (N_3422,N_2702,N_2137);
xnor U3423 (N_3423,N_2397,N_2368);
nand U3424 (N_3424,N_2355,N_2453);
xnor U3425 (N_3425,N_2592,N_2819);
nor U3426 (N_3426,N_2495,N_2409);
and U3427 (N_3427,N_2404,N_2891);
nor U3428 (N_3428,N_2338,N_2776);
xor U3429 (N_3429,N_2671,N_2049);
or U3430 (N_3430,N_2328,N_2900);
xnor U3431 (N_3431,N_2481,N_2784);
xor U3432 (N_3432,N_2529,N_2089);
nand U3433 (N_3433,N_2032,N_2042);
or U3434 (N_3434,N_2444,N_2575);
or U3435 (N_3435,N_2670,N_2099);
and U3436 (N_3436,N_2367,N_2512);
or U3437 (N_3437,N_2642,N_2883);
or U3438 (N_3438,N_2244,N_2542);
nor U3439 (N_3439,N_2119,N_2168);
and U3440 (N_3440,N_2122,N_2825);
nor U3441 (N_3441,N_2179,N_2339);
and U3442 (N_3442,N_2873,N_2076);
xor U3443 (N_3443,N_2583,N_2541);
xnor U3444 (N_3444,N_2373,N_2908);
xor U3445 (N_3445,N_2006,N_2937);
nand U3446 (N_3446,N_2361,N_2424);
nor U3447 (N_3447,N_2113,N_2904);
nor U3448 (N_3448,N_2108,N_2094);
xor U3449 (N_3449,N_2152,N_2666);
nor U3450 (N_3450,N_2455,N_2612);
or U3451 (N_3451,N_2565,N_2130);
or U3452 (N_3452,N_2321,N_2211);
nand U3453 (N_3453,N_2939,N_2131);
nand U3454 (N_3454,N_2187,N_2911);
and U3455 (N_3455,N_2497,N_2366);
nand U3456 (N_3456,N_2095,N_2185);
nor U3457 (N_3457,N_2026,N_2955);
nor U3458 (N_3458,N_2633,N_2625);
nor U3459 (N_3459,N_2072,N_2842);
nand U3460 (N_3460,N_2109,N_2342);
or U3461 (N_3461,N_2770,N_2796);
or U3462 (N_3462,N_2657,N_2859);
nand U3463 (N_3463,N_2743,N_2977);
xor U3464 (N_3464,N_2787,N_2820);
xnor U3465 (N_3465,N_2535,N_2292);
nor U3466 (N_3466,N_2643,N_2205);
or U3467 (N_3467,N_2223,N_2830);
or U3468 (N_3468,N_2304,N_2990);
and U3469 (N_3469,N_2473,N_2380);
nor U3470 (N_3470,N_2539,N_2267);
or U3471 (N_3471,N_2810,N_2871);
nor U3472 (N_3472,N_2298,N_2778);
xnor U3473 (N_3473,N_2097,N_2423);
nand U3474 (N_3474,N_2672,N_2902);
nor U3475 (N_3475,N_2290,N_2518);
xor U3476 (N_3476,N_2589,N_2245);
nand U3477 (N_3477,N_2889,N_2636);
xor U3478 (N_3478,N_2698,N_2514);
nand U3479 (N_3479,N_2441,N_2864);
and U3480 (N_3480,N_2916,N_2105);
nor U3481 (N_3481,N_2012,N_2014);
or U3482 (N_3482,N_2501,N_2703);
nor U3483 (N_3483,N_2092,N_2584);
xnor U3484 (N_3484,N_2222,N_2490);
and U3485 (N_3485,N_2375,N_2199);
nor U3486 (N_3486,N_2822,N_2577);
nor U3487 (N_3487,N_2662,N_2781);
xnor U3488 (N_3488,N_2173,N_2989);
nor U3489 (N_3489,N_2765,N_2192);
xnor U3490 (N_3490,N_2915,N_2607);
xor U3491 (N_3491,N_2609,N_2142);
nand U3492 (N_3492,N_2688,N_2246);
nand U3493 (N_3493,N_2593,N_2029);
xor U3494 (N_3494,N_2692,N_2041);
nor U3495 (N_3495,N_2145,N_2462);
or U3496 (N_3496,N_2833,N_2064);
nor U3497 (N_3497,N_2126,N_2210);
xor U3498 (N_3498,N_2586,N_2470);
nor U3499 (N_3499,N_2975,N_2768);
nand U3500 (N_3500,N_2232,N_2943);
xor U3501 (N_3501,N_2460,N_2682);
and U3502 (N_3502,N_2330,N_2081);
and U3503 (N_3503,N_2366,N_2468);
xor U3504 (N_3504,N_2770,N_2668);
nor U3505 (N_3505,N_2707,N_2940);
and U3506 (N_3506,N_2649,N_2207);
xnor U3507 (N_3507,N_2065,N_2367);
xnor U3508 (N_3508,N_2029,N_2436);
nor U3509 (N_3509,N_2765,N_2478);
nand U3510 (N_3510,N_2227,N_2277);
and U3511 (N_3511,N_2045,N_2762);
xor U3512 (N_3512,N_2651,N_2932);
and U3513 (N_3513,N_2864,N_2190);
nand U3514 (N_3514,N_2969,N_2088);
nand U3515 (N_3515,N_2040,N_2188);
nand U3516 (N_3516,N_2254,N_2721);
nand U3517 (N_3517,N_2644,N_2223);
nor U3518 (N_3518,N_2710,N_2613);
and U3519 (N_3519,N_2006,N_2369);
xnor U3520 (N_3520,N_2207,N_2119);
and U3521 (N_3521,N_2969,N_2340);
xnor U3522 (N_3522,N_2302,N_2071);
xor U3523 (N_3523,N_2062,N_2543);
xor U3524 (N_3524,N_2708,N_2008);
nor U3525 (N_3525,N_2916,N_2552);
nand U3526 (N_3526,N_2650,N_2329);
xor U3527 (N_3527,N_2798,N_2031);
or U3528 (N_3528,N_2489,N_2652);
or U3529 (N_3529,N_2060,N_2767);
and U3530 (N_3530,N_2329,N_2060);
xnor U3531 (N_3531,N_2895,N_2903);
xor U3532 (N_3532,N_2270,N_2984);
and U3533 (N_3533,N_2103,N_2470);
nand U3534 (N_3534,N_2678,N_2030);
or U3535 (N_3535,N_2629,N_2285);
and U3536 (N_3536,N_2368,N_2396);
or U3537 (N_3537,N_2589,N_2900);
nand U3538 (N_3538,N_2119,N_2822);
or U3539 (N_3539,N_2039,N_2574);
nand U3540 (N_3540,N_2633,N_2234);
or U3541 (N_3541,N_2150,N_2679);
or U3542 (N_3542,N_2916,N_2756);
or U3543 (N_3543,N_2884,N_2602);
and U3544 (N_3544,N_2304,N_2081);
xnor U3545 (N_3545,N_2287,N_2713);
xnor U3546 (N_3546,N_2847,N_2444);
and U3547 (N_3547,N_2862,N_2684);
nor U3548 (N_3548,N_2628,N_2038);
or U3549 (N_3549,N_2386,N_2681);
and U3550 (N_3550,N_2672,N_2823);
xnor U3551 (N_3551,N_2896,N_2425);
nor U3552 (N_3552,N_2533,N_2144);
nand U3553 (N_3553,N_2743,N_2563);
and U3554 (N_3554,N_2914,N_2038);
nor U3555 (N_3555,N_2010,N_2333);
and U3556 (N_3556,N_2992,N_2286);
xor U3557 (N_3557,N_2981,N_2429);
and U3558 (N_3558,N_2268,N_2205);
nand U3559 (N_3559,N_2919,N_2403);
xor U3560 (N_3560,N_2304,N_2637);
xor U3561 (N_3561,N_2017,N_2234);
nand U3562 (N_3562,N_2851,N_2825);
nor U3563 (N_3563,N_2708,N_2486);
nand U3564 (N_3564,N_2476,N_2919);
nand U3565 (N_3565,N_2436,N_2714);
or U3566 (N_3566,N_2357,N_2057);
nor U3567 (N_3567,N_2784,N_2605);
xor U3568 (N_3568,N_2146,N_2526);
nand U3569 (N_3569,N_2873,N_2984);
xnor U3570 (N_3570,N_2206,N_2841);
nand U3571 (N_3571,N_2230,N_2263);
or U3572 (N_3572,N_2962,N_2375);
xor U3573 (N_3573,N_2920,N_2220);
and U3574 (N_3574,N_2055,N_2469);
and U3575 (N_3575,N_2138,N_2488);
or U3576 (N_3576,N_2377,N_2288);
and U3577 (N_3577,N_2369,N_2207);
or U3578 (N_3578,N_2341,N_2065);
and U3579 (N_3579,N_2427,N_2529);
nand U3580 (N_3580,N_2662,N_2151);
and U3581 (N_3581,N_2091,N_2386);
xor U3582 (N_3582,N_2758,N_2811);
nor U3583 (N_3583,N_2089,N_2380);
xor U3584 (N_3584,N_2173,N_2268);
or U3585 (N_3585,N_2683,N_2734);
or U3586 (N_3586,N_2210,N_2901);
and U3587 (N_3587,N_2296,N_2282);
nand U3588 (N_3588,N_2622,N_2397);
and U3589 (N_3589,N_2001,N_2216);
xor U3590 (N_3590,N_2565,N_2587);
and U3591 (N_3591,N_2175,N_2179);
nand U3592 (N_3592,N_2906,N_2355);
and U3593 (N_3593,N_2555,N_2361);
nor U3594 (N_3594,N_2100,N_2594);
and U3595 (N_3595,N_2591,N_2867);
xnor U3596 (N_3596,N_2446,N_2537);
nor U3597 (N_3597,N_2164,N_2651);
nand U3598 (N_3598,N_2246,N_2605);
nor U3599 (N_3599,N_2228,N_2103);
xnor U3600 (N_3600,N_2819,N_2199);
xor U3601 (N_3601,N_2435,N_2867);
xnor U3602 (N_3602,N_2906,N_2251);
nor U3603 (N_3603,N_2919,N_2267);
nand U3604 (N_3604,N_2704,N_2622);
xnor U3605 (N_3605,N_2026,N_2229);
xnor U3606 (N_3606,N_2801,N_2695);
nor U3607 (N_3607,N_2687,N_2286);
and U3608 (N_3608,N_2315,N_2391);
or U3609 (N_3609,N_2844,N_2172);
xnor U3610 (N_3610,N_2646,N_2160);
or U3611 (N_3611,N_2895,N_2846);
or U3612 (N_3612,N_2687,N_2712);
and U3613 (N_3613,N_2098,N_2659);
or U3614 (N_3614,N_2616,N_2452);
or U3615 (N_3615,N_2315,N_2168);
nor U3616 (N_3616,N_2700,N_2795);
and U3617 (N_3617,N_2605,N_2624);
or U3618 (N_3618,N_2351,N_2211);
and U3619 (N_3619,N_2175,N_2779);
or U3620 (N_3620,N_2691,N_2511);
nand U3621 (N_3621,N_2875,N_2614);
and U3622 (N_3622,N_2147,N_2373);
or U3623 (N_3623,N_2298,N_2912);
and U3624 (N_3624,N_2144,N_2692);
nor U3625 (N_3625,N_2687,N_2019);
or U3626 (N_3626,N_2267,N_2910);
or U3627 (N_3627,N_2803,N_2854);
nand U3628 (N_3628,N_2877,N_2950);
and U3629 (N_3629,N_2484,N_2742);
and U3630 (N_3630,N_2795,N_2550);
nor U3631 (N_3631,N_2114,N_2155);
and U3632 (N_3632,N_2759,N_2852);
and U3633 (N_3633,N_2327,N_2096);
nand U3634 (N_3634,N_2078,N_2059);
and U3635 (N_3635,N_2762,N_2842);
or U3636 (N_3636,N_2545,N_2233);
or U3637 (N_3637,N_2097,N_2597);
xnor U3638 (N_3638,N_2227,N_2707);
xnor U3639 (N_3639,N_2335,N_2969);
nor U3640 (N_3640,N_2663,N_2113);
and U3641 (N_3641,N_2781,N_2106);
or U3642 (N_3642,N_2289,N_2344);
and U3643 (N_3643,N_2617,N_2685);
xnor U3644 (N_3644,N_2899,N_2723);
or U3645 (N_3645,N_2922,N_2780);
or U3646 (N_3646,N_2796,N_2982);
or U3647 (N_3647,N_2365,N_2987);
or U3648 (N_3648,N_2664,N_2299);
nand U3649 (N_3649,N_2030,N_2949);
or U3650 (N_3650,N_2857,N_2751);
nor U3651 (N_3651,N_2782,N_2127);
and U3652 (N_3652,N_2484,N_2476);
nand U3653 (N_3653,N_2392,N_2646);
or U3654 (N_3654,N_2928,N_2641);
or U3655 (N_3655,N_2570,N_2561);
xnor U3656 (N_3656,N_2048,N_2114);
or U3657 (N_3657,N_2205,N_2339);
or U3658 (N_3658,N_2534,N_2290);
xor U3659 (N_3659,N_2666,N_2209);
xnor U3660 (N_3660,N_2979,N_2614);
and U3661 (N_3661,N_2289,N_2069);
and U3662 (N_3662,N_2486,N_2764);
and U3663 (N_3663,N_2132,N_2467);
or U3664 (N_3664,N_2077,N_2379);
nor U3665 (N_3665,N_2225,N_2057);
nand U3666 (N_3666,N_2240,N_2580);
and U3667 (N_3667,N_2750,N_2345);
nor U3668 (N_3668,N_2382,N_2578);
nand U3669 (N_3669,N_2023,N_2252);
and U3670 (N_3670,N_2887,N_2232);
xnor U3671 (N_3671,N_2857,N_2701);
nand U3672 (N_3672,N_2851,N_2580);
nor U3673 (N_3673,N_2387,N_2806);
xor U3674 (N_3674,N_2726,N_2009);
and U3675 (N_3675,N_2872,N_2771);
and U3676 (N_3676,N_2879,N_2090);
nor U3677 (N_3677,N_2078,N_2221);
nand U3678 (N_3678,N_2079,N_2359);
nor U3679 (N_3679,N_2268,N_2434);
nand U3680 (N_3680,N_2646,N_2816);
or U3681 (N_3681,N_2686,N_2493);
and U3682 (N_3682,N_2381,N_2710);
and U3683 (N_3683,N_2241,N_2389);
and U3684 (N_3684,N_2383,N_2575);
xor U3685 (N_3685,N_2986,N_2837);
nor U3686 (N_3686,N_2723,N_2292);
or U3687 (N_3687,N_2673,N_2744);
or U3688 (N_3688,N_2671,N_2965);
nor U3689 (N_3689,N_2758,N_2200);
or U3690 (N_3690,N_2286,N_2956);
or U3691 (N_3691,N_2959,N_2865);
nand U3692 (N_3692,N_2857,N_2470);
and U3693 (N_3693,N_2304,N_2395);
nand U3694 (N_3694,N_2537,N_2771);
nand U3695 (N_3695,N_2971,N_2883);
or U3696 (N_3696,N_2944,N_2725);
or U3697 (N_3697,N_2524,N_2199);
nor U3698 (N_3698,N_2281,N_2884);
or U3699 (N_3699,N_2551,N_2389);
or U3700 (N_3700,N_2970,N_2104);
xnor U3701 (N_3701,N_2433,N_2462);
or U3702 (N_3702,N_2759,N_2463);
nor U3703 (N_3703,N_2852,N_2287);
and U3704 (N_3704,N_2236,N_2523);
nor U3705 (N_3705,N_2504,N_2728);
nor U3706 (N_3706,N_2048,N_2867);
or U3707 (N_3707,N_2325,N_2131);
and U3708 (N_3708,N_2583,N_2845);
and U3709 (N_3709,N_2824,N_2830);
and U3710 (N_3710,N_2457,N_2020);
and U3711 (N_3711,N_2890,N_2537);
nand U3712 (N_3712,N_2216,N_2525);
and U3713 (N_3713,N_2394,N_2537);
and U3714 (N_3714,N_2634,N_2481);
xor U3715 (N_3715,N_2654,N_2165);
nor U3716 (N_3716,N_2218,N_2732);
and U3717 (N_3717,N_2820,N_2164);
and U3718 (N_3718,N_2611,N_2927);
and U3719 (N_3719,N_2036,N_2273);
nor U3720 (N_3720,N_2998,N_2111);
and U3721 (N_3721,N_2968,N_2525);
and U3722 (N_3722,N_2135,N_2072);
nor U3723 (N_3723,N_2936,N_2389);
and U3724 (N_3724,N_2074,N_2261);
nand U3725 (N_3725,N_2178,N_2835);
or U3726 (N_3726,N_2160,N_2164);
xnor U3727 (N_3727,N_2363,N_2687);
or U3728 (N_3728,N_2129,N_2345);
nor U3729 (N_3729,N_2231,N_2861);
nor U3730 (N_3730,N_2431,N_2306);
xor U3731 (N_3731,N_2463,N_2815);
or U3732 (N_3732,N_2817,N_2421);
nor U3733 (N_3733,N_2101,N_2461);
nor U3734 (N_3734,N_2999,N_2540);
xnor U3735 (N_3735,N_2543,N_2022);
nand U3736 (N_3736,N_2791,N_2431);
and U3737 (N_3737,N_2125,N_2731);
nor U3738 (N_3738,N_2414,N_2962);
and U3739 (N_3739,N_2443,N_2854);
xor U3740 (N_3740,N_2672,N_2109);
xor U3741 (N_3741,N_2156,N_2535);
and U3742 (N_3742,N_2437,N_2829);
xnor U3743 (N_3743,N_2803,N_2677);
nor U3744 (N_3744,N_2009,N_2288);
xor U3745 (N_3745,N_2383,N_2952);
nand U3746 (N_3746,N_2762,N_2684);
nand U3747 (N_3747,N_2359,N_2865);
xnor U3748 (N_3748,N_2217,N_2525);
and U3749 (N_3749,N_2891,N_2270);
nor U3750 (N_3750,N_2843,N_2180);
xnor U3751 (N_3751,N_2447,N_2526);
and U3752 (N_3752,N_2329,N_2691);
nand U3753 (N_3753,N_2843,N_2587);
xnor U3754 (N_3754,N_2915,N_2090);
nand U3755 (N_3755,N_2517,N_2296);
and U3756 (N_3756,N_2649,N_2900);
or U3757 (N_3757,N_2237,N_2496);
and U3758 (N_3758,N_2596,N_2606);
nor U3759 (N_3759,N_2062,N_2271);
nand U3760 (N_3760,N_2381,N_2688);
nand U3761 (N_3761,N_2830,N_2661);
and U3762 (N_3762,N_2536,N_2956);
or U3763 (N_3763,N_2714,N_2400);
nand U3764 (N_3764,N_2094,N_2907);
or U3765 (N_3765,N_2563,N_2500);
nand U3766 (N_3766,N_2465,N_2116);
and U3767 (N_3767,N_2132,N_2779);
or U3768 (N_3768,N_2752,N_2649);
xor U3769 (N_3769,N_2151,N_2686);
nor U3770 (N_3770,N_2718,N_2352);
and U3771 (N_3771,N_2953,N_2751);
nand U3772 (N_3772,N_2445,N_2545);
and U3773 (N_3773,N_2210,N_2601);
or U3774 (N_3774,N_2350,N_2196);
nor U3775 (N_3775,N_2593,N_2256);
nor U3776 (N_3776,N_2255,N_2468);
and U3777 (N_3777,N_2072,N_2119);
nor U3778 (N_3778,N_2902,N_2164);
nand U3779 (N_3779,N_2944,N_2810);
nor U3780 (N_3780,N_2359,N_2456);
xnor U3781 (N_3781,N_2554,N_2386);
and U3782 (N_3782,N_2433,N_2954);
or U3783 (N_3783,N_2907,N_2932);
xnor U3784 (N_3784,N_2574,N_2000);
and U3785 (N_3785,N_2142,N_2178);
nor U3786 (N_3786,N_2407,N_2878);
or U3787 (N_3787,N_2925,N_2211);
xor U3788 (N_3788,N_2519,N_2036);
nor U3789 (N_3789,N_2427,N_2081);
nand U3790 (N_3790,N_2076,N_2306);
nand U3791 (N_3791,N_2514,N_2133);
nor U3792 (N_3792,N_2894,N_2650);
and U3793 (N_3793,N_2424,N_2672);
and U3794 (N_3794,N_2450,N_2265);
or U3795 (N_3795,N_2856,N_2115);
xnor U3796 (N_3796,N_2317,N_2200);
nand U3797 (N_3797,N_2576,N_2718);
or U3798 (N_3798,N_2327,N_2635);
or U3799 (N_3799,N_2402,N_2375);
xnor U3800 (N_3800,N_2650,N_2125);
nand U3801 (N_3801,N_2259,N_2967);
nand U3802 (N_3802,N_2490,N_2657);
and U3803 (N_3803,N_2847,N_2492);
xor U3804 (N_3804,N_2644,N_2332);
nand U3805 (N_3805,N_2803,N_2829);
or U3806 (N_3806,N_2696,N_2490);
and U3807 (N_3807,N_2380,N_2902);
nor U3808 (N_3808,N_2309,N_2390);
or U3809 (N_3809,N_2186,N_2706);
nor U3810 (N_3810,N_2744,N_2612);
or U3811 (N_3811,N_2088,N_2758);
nor U3812 (N_3812,N_2226,N_2539);
nor U3813 (N_3813,N_2122,N_2005);
nand U3814 (N_3814,N_2493,N_2833);
nand U3815 (N_3815,N_2458,N_2678);
nor U3816 (N_3816,N_2205,N_2951);
xnor U3817 (N_3817,N_2205,N_2381);
nor U3818 (N_3818,N_2035,N_2307);
and U3819 (N_3819,N_2444,N_2845);
nand U3820 (N_3820,N_2367,N_2641);
nand U3821 (N_3821,N_2990,N_2408);
nor U3822 (N_3822,N_2261,N_2358);
nor U3823 (N_3823,N_2423,N_2031);
and U3824 (N_3824,N_2128,N_2498);
or U3825 (N_3825,N_2905,N_2763);
and U3826 (N_3826,N_2230,N_2701);
xnor U3827 (N_3827,N_2365,N_2715);
xnor U3828 (N_3828,N_2010,N_2582);
or U3829 (N_3829,N_2027,N_2750);
and U3830 (N_3830,N_2518,N_2736);
nand U3831 (N_3831,N_2654,N_2710);
nand U3832 (N_3832,N_2017,N_2387);
or U3833 (N_3833,N_2458,N_2707);
nand U3834 (N_3834,N_2579,N_2608);
xor U3835 (N_3835,N_2470,N_2288);
nor U3836 (N_3836,N_2335,N_2227);
or U3837 (N_3837,N_2921,N_2226);
and U3838 (N_3838,N_2062,N_2682);
xnor U3839 (N_3839,N_2025,N_2926);
nand U3840 (N_3840,N_2395,N_2250);
nand U3841 (N_3841,N_2032,N_2121);
xnor U3842 (N_3842,N_2323,N_2441);
xor U3843 (N_3843,N_2919,N_2445);
xnor U3844 (N_3844,N_2266,N_2642);
or U3845 (N_3845,N_2410,N_2871);
nand U3846 (N_3846,N_2538,N_2842);
and U3847 (N_3847,N_2318,N_2886);
xnor U3848 (N_3848,N_2736,N_2369);
and U3849 (N_3849,N_2254,N_2438);
xor U3850 (N_3850,N_2368,N_2231);
nand U3851 (N_3851,N_2373,N_2125);
nand U3852 (N_3852,N_2691,N_2953);
xor U3853 (N_3853,N_2351,N_2792);
or U3854 (N_3854,N_2928,N_2450);
xor U3855 (N_3855,N_2229,N_2598);
and U3856 (N_3856,N_2405,N_2369);
xor U3857 (N_3857,N_2026,N_2029);
xnor U3858 (N_3858,N_2439,N_2965);
and U3859 (N_3859,N_2285,N_2155);
or U3860 (N_3860,N_2127,N_2972);
nand U3861 (N_3861,N_2285,N_2622);
nand U3862 (N_3862,N_2147,N_2364);
xnor U3863 (N_3863,N_2407,N_2460);
nand U3864 (N_3864,N_2985,N_2673);
nand U3865 (N_3865,N_2289,N_2857);
nand U3866 (N_3866,N_2951,N_2657);
nor U3867 (N_3867,N_2286,N_2765);
nor U3868 (N_3868,N_2747,N_2691);
and U3869 (N_3869,N_2646,N_2479);
and U3870 (N_3870,N_2593,N_2539);
xnor U3871 (N_3871,N_2157,N_2116);
and U3872 (N_3872,N_2101,N_2429);
and U3873 (N_3873,N_2698,N_2309);
xor U3874 (N_3874,N_2096,N_2047);
or U3875 (N_3875,N_2977,N_2401);
and U3876 (N_3876,N_2451,N_2222);
nand U3877 (N_3877,N_2693,N_2525);
and U3878 (N_3878,N_2577,N_2876);
xor U3879 (N_3879,N_2710,N_2382);
nor U3880 (N_3880,N_2222,N_2491);
and U3881 (N_3881,N_2329,N_2297);
or U3882 (N_3882,N_2427,N_2562);
nand U3883 (N_3883,N_2335,N_2591);
xnor U3884 (N_3884,N_2564,N_2119);
nand U3885 (N_3885,N_2593,N_2217);
and U3886 (N_3886,N_2133,N_2070);
and U3887 (N_3887,N_2531,N_2453);
nor U3888 (N_3888,N_2179,N_2103);
nand U3889 (N_3889,N_2510,N_2501);
and U3890 (N_3890,N_2067,N_2571);
xnor U3891 (N_3891,N_2104,N_2566);
or U3892 (N_3892,N_2269,N_2027);
nand U3893 (N_3893,N_2697,N_2351);
and U3894 (N_3894,N_2056,N_2401);
nand U3895 (N_3895,N_2251,N_2429);
nor U3896 (N_3896,N_2732,N_2427);
nand U3897 (N_3897,N_2553,N_2110);
nand U3898 (N_3898,N_2627,N_2914);
or U3899 (N_3899,N_2816,N_2927);
nor U3900 (N_3900,N_2792,N_2090);
nor U3901 (N_3901,N_2518,N_2789);
xnor U3902 (N_3902,N_2852,N_2301);
xor U3903 (N_3903,N_2643,N_2979);
nor U3904 (N_3904,N_2920,N_2734);
nand U3905 (N_3905,N_2956,N_2090);
xor U3906 (N_3906,N_2820,N_2932);
and U3907 (N_3907,N_2229,N_2729);
or U3908 (N_3908,N_2700,N_2584);
nand U3909 (N_3909,N_2203,N_2435);
xnor U3910 (N_3910,N_2396,N_2018);
nor U3911 (N_3911,N_2471,N_2629);
xor U3912 (N_3912,N_2264,N_2901);
or U3913 (N_3913,N_2338,N_2664);
or U3914 (N_3914,N_2621,N_2209);
and U3915 (N_3915,N_2156,N_2971);
or U3916 (N_3916,N_2275,N_2757);
nor U3917 (N_3917,N_2458,N_2054);
nor U3918 (N_3918,N_2230,N_2053);
xor U3919 (N_3919,N_2073,N_2829);
nand U3920 (N_3920,N_2903,N_2869);
or U3921 (N_3921,N_2039,N_2757);
or U3922 (N_3922,N_2829,N_2787);
nand U3923 (N_3923,N_2857,N_2341);
nand U3924 (N_3924,N_2929,N_2603);
xor U3925 (N_3925,N_2644,N_2943);
nand U3926 (N_3926,N_2847,N_2887);
nand U3927 (N_3927,N_2556,N_2041);
xnor U3928 (N_3928,N_2316,N_2597);
nand U3929 (N_3929,N_2939,N_2613);
nand U3930 (N_3930,N_2282,N_2537);
nand U3931 (N_3931,N_2507,N_2607);
nor U3932 (N_3932,N_2958,N_2903);
xor U3933 (N_3933,N_2510,N_2831);
or U3934 (N_3934,N_2525,N_2319);
nor U3935 (N_3935,N_2572,N_2209);
and U3936 (N_3936,N_2939,N_2748);
and U3937 (N_3937,N_2859,N_2182);
nor U3938 (N_3938,N_2301,N_2506);
and U3939 (N_3939,N_2526,N_2353);
xnor U3940 (N_3940,N_2859,N_2617);
xnor U3941 (N_3941,N_2135,N_2742);
xor U3942 (N_3942,N_2483,N_2689);
and U3943 (N_3943,N_2150,N_2256);
nand U3944 (N_3944,N_2628,N_2238);
or U3945 (N_3945,N_2923,N_2513);
xnor U3946 (N_3946,N_2786,N_2420);
xnor U3947 (N_3947,N_2834,N_2518);
nor U3948 (N_3948,N_2714,N_2198);
nor U3949 (N_3949,N_2728,N_2161);
or U3950 (N_3950,N_2494,N_2620);
and U3951 (N_3951,N_2308,N_2983);
and U3952 (N_3952,N_2322,N_2682);
nor U3953 (N_3953,N_2541,N_2560);
xnor U3954 (N_3954,N_2489,N_2852);
nor U3955 (N_3955,N_2970,N_2570);
or U3956 (N_3956,N_2782,N_2349);
nand U3957 (N_3957,N_2329,N_2045);
xor U3958 (N_3958,N_2500,N_2494);
and U3959 (N_3959,N_2563,N_2840);
and U3960 (N_3960,N_2610,N_2832);
and U3961 (N_3961,N_2209,N_2352);
nor U3962 (N_3962,N_2835,N_2239);
or U3963 (N_3963,N_2848,N_2840);
and U3964 (N_3964,N_2301,N_2347);
or U3965 (N_3965,N_2607,N_2983);
and U3966 (N_3966,N_2104,N_2998);
or U3967 (N_3967,N_2475,N_2822);
nor U3968 (N_3968,N_2557,N_2592);
nor U3969 (N_3969,N_2029,N_2008);
nor U3970 (N_3970,N_2365,N_2361);
and U3971 (N_3971,N_2388,N_2756);
nand U3972 (N_3972,N_2039,N_2207);
nand U3973 (N_3973,N_2649,N_2675);
and U3974 (N_3974,N_2994,N_2840);
nor U3975 (N_3975,N_2526,N_2791);
and U3976 (N_3976,N_2379,N_2847);
xnor U3977 (N_3977,N_2599,N_2958);
or U3978 (N_3978,N_2973,N_2573);
nor U3979 (N_3979,N_2453,N_2795);
xor U3980 (N_3980,N_2036,N_2809);
nand U3981 (N_3981,N_2568,N_2118);
nand U3982 (N_3982,N_2269,N_2671);
nor U3983 (N_3983,N_2303,N_2723);
nor U3984 (N_3984,N_2576,N_2903);
xnor U3985 (N_3985,N_2934,N_2322);
and U3986 (N_3986,N_2990,N_2993);
xor U3987 (N_3987,N_2915,N_2288);
or U3988 (N_3988,N_2345,N_2825);
xor U3989 (N_3989,N_2305,N_2119);
xnor U3990 (N_3990,N_2987,N_2210);
and U3991 (N_3991,N_2147,N_2133);
or U3992 (N_3992,N_2206,N_2518);
and U3993 (N_3993,N_2798,N_2775);
or U3994 (N_3994,N_2207,N_2455);
xor U3995 (N_3995,N_2781,N_2698);
and U3996 (N_3996,N_2525,N_2196);
xor U3997 (N_3997,N_2668,N_2234);
nor U3998 (N_3998,N_2731,N_2909);
nor U3999 (N_3999,N_2209,N_2516);
nand U4000 (N_4000,N_3496,N_3463);
or U4001 (N_4001,N_3744,N_3650);
and U4002 (N_4002,N_3702,N_3751);
nand U4003 (N_4003,N_3003,N_3637);
xnor U4004 (N_4004,N_3665,N_3449);
or U4005 (N_4005,N_3500,N_3270);
nor U4006 (N_4006,N_3492,N_3838);
nor U4007 (N_4007,N_3269,N_3551);
xnor U4008 (N_4008,N_3651,N_3135);
nor U4009 (N_4009,N_3849,N_3935);
nand U4010 (N_4010,N_3450,N_3214);
or U4011 (N_4011,N_3313,N_3262);
xnor U4012 (N_4012,N_3824,N_3795);
and U4013 (N_4013,N_3895,N_3932);
nor U4014 (N_4014,N_3167,N_3521);
or U4015 (N_4015,N_3805,N_3557);
or U4016 (N_4016,N_3616,N_3470);
nand U4017 (N_4017,N_3993,N_3754);
and U4018 (N_4018,N_3326,N_3640);
xnor U4019 (N_4019,N_3355,N_3857);
or U4020 (N_4020,N_3042,N_3632);
and U4021 (N_4021,N_3462,N_3584);
xor U4022 (N_4022,N_3976,N_3447);
nor U4023 (N_4023,N_3207,N_3208);
nand U4024 (N_4024,N_3036,N_3051);
or U4025 (N_4025,N_3622,N_3002);
nand U4026 (N_4026,N_3115,N_3394);
nor U4027 (N_4027,N_3922,N_3393);
nand U4028 (N_4028,N_3337,N_3340);
or U4029 (N_4029,N_3310,N_3009);
xor U4030 (N_4030,N_3093,N_3037);
and U4031 (N_4031,N_3639,N_3627);
nor U4032 (N_4032,N_3726,N_3290);
and U4033 (N_4033,N_3113,N_3257);
nand U4034 (N_4034,N_3284,N_3690);
nand U4035 (N_4035,N_3867,N_3148);
nand U4036 (N_4036,N_3101,N_3728);
xor U4037 (N_4037,N_3069,N_3731);
and U4038 (N_4038,N_3593,N_3831);
xor U4039 (N_4039,N_3094,N_3634);
and U4040 (N_4040,N_3747,N_3397);
and U4041 (N_4041,N_3578,N_3966);
nand U4042 (N_4042,N_3890,N_3926);
and U4043 (N_4043,N_3095,N_3872);
and U4044 (N_4044,N_3717,N_3729);
nor U4045 (N_4045,N_3066,N_3361);
or U4046 (N_4046,N_3959,N_3794);
nand U4047 (N_4047,N_3373,N_3892);
or U4048 (N_4048,N_3352,N_3635);
nor U4049 (N_4049,N_3621,N_3230);
or U4050 (N_4050,N_3429,N_3520);
or U4051 (N_4051,N_3392,N_3772);
or U4052 (N_4052,N_3014,N_3955);
nand U4053 (N_4053,N_3711,N_3279);
nand U4054 (N_4054,N_3739,N_3811);
nand U4055 (N_4055,N_3797,N_3197);
nand U4056 (N_4056,N_3833,N_3385);
or U4057 (N_4057,N_3497,N_3885);
nand U4058 (N_4058,N_3937,N_3203);
nor U4059 (N_4059,N_3556,N_3212);
nand U4060 (N_4060,N_3855,N_3254);
nand U4061 (N_4061,N_3567,N_3399);
xnor U4062 (N_4062,N_3607,N_3939);
or U4063 (N_4063,N_3472,N_3043);
xor U4064 (N_4064,N_3952,N_3564);
nand U4065 (N_4065,N_3527,N_3765);
nand U4066 (N_4066,N_3968,N_3334);
or U4067 (N_4067,N_3341,N_3599);
nand U4068 (N_4068,N_3245,N_3484);
nor U4069 (N_4069,N_3327,N_3265);
and U4070 (N_4070,N_3718,N_3431);
nand U4071 (N_4071,N_3884,N_3495);
nand U4072 (N_4072,N_3998,N_3874);
nor U4073 (N_4073,N_3930,N_3630);
nand U4074 (N_4074,N_3905,N_3321);
nor U4075 (N_4075,N_3915,N_3151);
nand U4076 (N_4076,N_3682,N_3163);
nor U4077 (N_4077,N_3019,N_3364);
xnor U4078 (N_4078,N_3073,N_3901);
and U4079 (N_4079,N_3071,N_3818);
xnor U4080 (N_4080,N_3840,N_3445);
or U4081 (N_4081,N_3425,N_3878);
nand U4082 (N_4082,N_3129,N_3192);
nor U4083 (N_4083,N_3819,N_3376);
or U4084 (N_4084,N_3722,N_3238);
and U4085 (N_4085,N_3598,N_3343);
and U4086 (N_4086,N_3519,N_3542);
and U4087 (N_4087,N_3735,N_3414);
or U4088 (N_4088,N_3416,N_3807);
or U4089 (N_4089,N_3064,N_3684);
nand U4090 (N_4090,N_3098,N_3780);
nand U4091 (N_4091,N_3044,N_3286);
and U4092 (N_4092,N_3137,N_3736);
and U4093 (N_4093,N_3276,N_3015);
nor U4094 (N_4094,N_3712,N_3963);
nor U4095 (N_4095,N_3215,N_3329);
or U4096 (N_4096,N_3038,N_3268);
nor U4097 (N_4097,N_3832,N_3891);
and U4098 (N_4098,N_3443,N_3454);
xnor U4099 (N_4099,N_3177,N_3703);
and U4100 (N_4100,N_3132,N_3530);
xor U4101 (N_4101,N_3881,N_3656);
or U4102 (N_4102,N_3107,N_3048);
or U4103 (N_4103,N_3689,N_3304);
xor U4104 (N_4104,N_3802,N_3216);
xnor U4105 (N_4105,N_3017,N_3829);
nand U4106 (N_4106,N_3349,N_3750);
or U4107 (N_4107,N_3478,N_3150);
and U4108 (N_4108,N_3827,N_3408);
or U4109 (N_4109,N_3236,N_3675);
and U4110 (N_4110,N_3390,N_3025);
or U4111 (N_4111,N_3929,N_3446);
nand U4112 (N_4112,N_3138,N_3468);
nor U4113 (N_4113,N_3263,N_3790);
nor U4114 (N_4114,N_3547,N_3130);
and U4115 (N_4115,N_3152,N_3055);
or U4116 (N_4116,N_3205,N_3474);
or U4117 (N_4117,N_3652,N_3219);
or U4118 (N_4118,N_3610,N_3312);
xnor U4119 (N_4119,N_3237,N_3260);
xor U4120 (N_4120,N_3725,N_3285);
nor U4121 (N_4121,N_3283,N_3879);
nand U4122 (N_4122,N_3620,N_3605);
xnor U4123 (N_4123,N_3169,N_3866);
nand U4124 (N_4124,N_3302,N_3916);
nor U4125 (N_4125,N_3843,N_3409);
and U4126 (N_4126,N_3767,N_3836);
or U4127 (N_4127,N_3110,N_3581);
nand U4128 (N_4128,N_3781,N_3315);
nor U4129 (N_4129,N_3332,N_3004);
xnor U4130 (N_4130,N_3774,N_3104);
nand U4131 (N_4131,N_3858,N_3515);
or U4132 (N_4132,N_3602,N_3835);
and U4133 (N_4133,N_3041,N_3424);
xnor U4134 (N_4134,N_3995,N_3295);
nor U4135 (N_4135,N_3422,N_3360);
xor U4136 (N_4136,N_3507,N_3733);
or U4137 (N_4137,N_3075,N_3821);
or U4138 (N_4138,N_3126,N_3058);
nand U4139 (N_4139,N_3940,N_3411);
nand U4140 (N_4140,N_3097,N_3938);
nor U4141 (N_4141,N_3145,N_3924);
nor U4142 (N_4142,N_3413,N_3859);
or U4143 (N_4143,N_3034,N_3758);
xnor U4144 (N_4144,N_3994,N_3860);
nor U4145 (N_4145,N_3643,N_3812);
nand U4146 (N_4146,N_3681,N_3603);
and U4147 (N_4147,N_3168,N_3294);
nand U4148 (N_4148,N_3080,N_3172);
nor U4149 (N_4149,N_3190,N_3089);
or U4150 (N_4150,N_3655,N_3629);
nand U4151 (N_4151,N_3691,N_3856);
nand U4152 (N_4152,N_3708,N_3421);
nand U4153 (N_4153,N_3165,N_3367);
or U4154 (N_4154,N_3473,N_3768);
nor U4155 (N_4155,N_3287,N_3776);
xor U4156 (N_4156,N_3377,N_3523);
nor U4157 (N_4157,N_3442,N_3218);
and U4158 (N_4158,N_3911,N_3773);
and U4159 (N_4159,N_3186,N_3088);
nand U4160 (N_4160,N_3202,N_3518);
xnor U4161 (N_4161,N_3756,N_3585);
or U4162 (N_4162,N_3980,N_3432);
or U4163 (N_4163,N_3488,N_3252);
xnor U4164 (N_4164,N_3986,N_3510);
or U4165 (N_4165,N_3160,N_3699);
and U4166 (N_4166,N_3301,N_3128);
or U4167 (N_4167,N_3996,N_3391);
nand U4168 (N_4168,N_3091,N_3382);
nor U4169 (N_4169,N_3493,N_3734);
nand U4170 (N_4170,N_3970,N_3694);
xor U4171 (N_4171,N_3589,N_3346);
nand U4172 (N_4172,N_3083,N_3925);
xnor U4173 (N_4173,N_3062,N_3412);
and U4174 (N_4174,N_3224,N_3727);
and U4175 (N_4175,N_3330,N_3513);
nand U4176 (N_4176,N_3876,N_3792);
and U4177 (N_4177,N_3503,N_3297);
nand U4178 (N_4178,N_3577,N_3828);
nor U4179 (N_4179,N_3181,N_3716);
nand U4180 (N_4180,N_3668,N_3457);
or U4181 (N_4181,N_3992,N_3369);
xnor U4182 (N_4182,N_3389,N_3316);
xor U4183 (N_4183,N_3788,N_3809);
and U4184 (N_4184,N_3264,N_3914);
and U4185 (N_4185,N_3806,N_3875);
xor U4186 (N_4186,N_3842,N_3331);
nor U4187 (N_4187,N_3526,N_3789);
nor U4188 (N_4188,N_3056,N_3837);
or U4189 (N_4189,N_3125,N_3335);
or U4190 (N_4190,N_3933,N_3653);
and U4191 (N_4191,N_3345,N_3848);
nor U4192 (N_4192,N_3082,N_3841);
and U4193 (N_4193,N_3498,N_3235);
nor U4194 (N_4194,N_3005,N_3396);
or U4195 (N_4195,N_3199,N_3437);
nand U4196 (N_4196,N_3453,N_3477);
xnor U4197 (N_4197,N_3149,N_3823);
or U4198 (N_4198,N_3957,N_3719);
and U4199 (N_4199,N_3989,N_3491);
and U4200 (N_4200,N_3763,N_3969);
nand U4201 (N_4201,N_3886,N_3775);
or U4202 (N_4202,N_3375,N_3371);
nor U4203 (N_4203,N_3956,N_3291);
nand U4204 (N_4204,N_3024,N_3325);
and U4205 (N_4205,N_3196,N_3779);
xor U4206 (N_4206,N_3534,N_3971);
nor U4207 (N_4207,N_3535,N_3626);
or U4208 (N_4208,N_3580,N_3464);
and U4209 (N_4209,N_3545,N_3814);
or U4210 (N_4210,N_3942,N_3870);
xnor U4211 (N_4211,N_3465,N_3839);
nor U4212 (N_4212,N_3673,N_3380);
nor U4213 (N_4213,N_3180,N_3723);
xor U4214 (N_4214,N_3067,N_3174);
and U4215 (N_4215,N_3973,N_3808);
and U4216 (N_4216,N_3524,N_3121);
xnor U4217 (N_4217,N_3710,N_3919);
xnor U4218 (N_4218,N_3090,N_3271);
xnor U4219 (N_4219,N_3013,N_3509);
or U4220 (N_4220,N_3060,N_3695);
or U4221 (N_4221,N_3553,N_3575);
xnor U4222 (N_4222,N_3221,N_3793);
or U4223 (N_4223,N_3123,N_3894);
xor U4224 (N_4224,N_3501,N_3749);
nand U4225 (N_4225,N_3240,N_3983);
or U4226 (N_4226,N_3601,N_3008);
nor U4227 (N_4227,N_3517,N_3537);
nand U4228 (N_4228,N_3381,N_3225);
xor U4229 (N_4229,N_3687,N_3825);
and U4230 (N_4230,N_3159,N_3011);
nand U4231 (N_4231,N_3877,N_3666);
and U4232 (N_4232,N_3210,N_3554);
and U4233 (N_4233,N_3247,N_3906);
or U4234 (N_4234,N_3579,N_3228);
or U4235 (N_4235,N_3344,N_3303);
and U4236 (N_4236,N_3696,N_3991);
and U4237 (N_4237,N_3158,N_3587);
and U4238 (N_4238,N_3931,N_3372);
nand U4239 (N_4239,N_3012,N_3977);
nor U4240 (N_4240,N_3748,N_3538);
nand U4241 (N_4241,N_3006,N_3568);
and U4242 (N_4242,N_3489,N_3786);
nor U4243 (N_4243,N_3198,N_3118);
xnor U4244 (N_4244,N_3461,N_3647);
xor U4245 (N_4245,N_3040,N_3280);
nand U4246 (N_4246,N_3423,N_3282);
or U4247 (N_4247,N_3189,N_3570);
nor U4248 (N_4248,N_3179,N_3760);
nand U4249 (N_4249,N_3573,N_3713);
xor U4250 (N_4250,N_3398,N_3374);
and U4251 (N_4251,N_3288,N_3810);
and U4252 (N_4252,N_3033,N_3541);
nand U4253 (N_4253,N_3106,N_3532);
nor U4254 (N_4254,N_3771,N_3596);
and U4255 (N_4255,N_3074,N_3417);
nand U4256 (N_4256,N_3927,N_3904);
nor U4257 (N_4257,N_3613,N_3427);
nor U4258 (N_4258,N_3117,N_3709);
and U4259 (N_4259,N_3897,N_3333);
nor U4260 (N_4260,N_3267,N_3920);
xnor U4261 (N_4261,N_3997,N_3528);
nand U4262 (N_4262,N_3102,N_3657);
and U4263 (N_4263,N_3258,N_3898);
and U4264 (N_4264,N_3582,N_3428);
nand U4265 (N_4265,N_3363,N_3590);
nor U4266 (N_4266,N_3544,N_3173);
xor U4267 (N_4267,N_3761,N_3045);
nor U4268 (N_4268,N_3863,N_3595);
nor U4269 (N_4269,N_3241,N_3830);
nor U4270 (N_4270,N_3155,N_3027);
and U4271 (N_4271,N_3623,N_3184);
and U4272 (N_4272,N_3949,N_3307);
nand U4273 (N_4273,N_3063,N_3274);
and U4274 (N_4274,N_3299,N_3248);
or U4275 (N_4275,N_3109,N_3944);
xnor U4276 (N_4276,N_3693,N_3068);
nor U4277 (N_4277,N_3338,N_3705);
and U4278 (N_4278,N_3234,N_3049);
and U4279 (N_4279,N_3482,N_3441);
and U4280 (N_4280,N_3921,N_3686);
or U4281 (N_4281,N_3813,N_3958);
or U4282 (N_4282,N_3249,N_3318);
and U4283 (N_4283,N_3434,N_3746);
nor U4284 (N_4284,N_3420,N_3146);
or U4285 (N_4285,N_3591,N_3801);
nand U4286 (N_4286,N_3592,N_3559);
nor U4287 (N_4287,N_3999,N_3153);
xnor U4288 (N_4288,N_3663,N_3784);
xor U4289 (N_4289,N_3239,N_3383);
xnor U4290 (N_4290,N_3755,N_3231);
nor U4291 (N_4291,N_3990,N_3913);
and U4292 (N_4292,N_3444,N_3365);
nand U4293 (N_4293,N_3139,N_3026);
nor U4294 (N_4294,N_3426,N_3182);
nor U4295 (N_4295,N_3743,N_3514);
and U4296 (N_4296,N_3679,N_3311);
nand U4297 (N_4297,N_3759,N_3671);
or U4298 (N_4298,N_3609,N_3982);
nor U4299 (N_4299,N_3936,N_3079);
nand U4300 (N_4300,N_3688,N_3407);
nand U4301 (N_4301,N_3851,N_3220);
nor U4302 (N_4302,N_3753,N_3550);
xor U4303 (N_4303,N_3256,N_3644);
xnor U4304 (N_4304,N_3834,N_3571);
and U4305 (N_4305,N_3010,N_3529);
nor U4306 (N_4306,N_3560,N_3979);
nand U4307 (N_4307,N_3471,N_3084);
or U4308 (N_4308,N_3386,N_3868);
or U4309 (N_4309,N_3661,N_3370);
or U4310 (N_4310,N_3029,N_3406);
or U4311 (N_4311,N_3562,N_3880);
nand U4312 (N_4312,N_3531,N_3378);
or U4313 (N_4313,N_3309,N_3972);
nand U4314 (N_4314,N_3561,N_3960);
nand U4315 (N_4315,N_3078,N_3511);
nor U4316 (N_4316,N_3401,N_3193);
nor U4317 (N_4317,N_3762,N_3116);
xor U4318 (N_4318,N_3604,N_3777);
nand U4319 (N_4319,N_3853,N_3065);
nand U4320 (N_4320,N_3854,N_3120);
and U4321 (N_4321,N_3483,N_3502);
nand U4322 (N_4322,N_3804,N_3893);
xnor U4323 (N_4323,N_3251,N_3978);
nor U4324 (N_4324,N_3147,N_3485);
nor U4325 (N_4325,N_3730,N_3667);
and U4326 (N_4326,N_3233,N_3188);
nor U4327 (N_4327,N_3354,N_3617);
or U4328 (N_4328,N_3574,N_3171);
xor U4329 (N_4329,N_3720,N_3206);
nor U4330 (N_4330,N_3273,N_3974);
and U4331 (N_4331,N_3319,N_3862);
and U4332 (N_4332,N_3259,N_3817);
xnor U4333 (N_4333,N_3964,N_3481);
xor U4334 (N_4334,N_3266,N_3648);
or U4335 (N_4335,N_3050,N_3016);
nand U4336 (N_4336,N_3096,N_3296);
xor U4337 (N_4337,N_3244,N_3070);
nand U4338 (N_4338,N_3882,N_3680);
and U4339 (N_4339,N_3324,N_3742);
nor U4340 (N_4340,N_3451,N_3685);
or U4341 (N_4341,N_3466,N_3250);
and U4342 (N_4342,N_3323,N_3984);
nor U4343 (N_4343,N_3628,N_3134);
nand U4344 (N_4344,N_3111,N_3918);
xor U4345 (N_4345,N_3764,N_3439);
xor U4346 (N_4346,N_3030,N_3700);
xnor U4347 (N_4347,N_3458,N_3945);
and U4348 (N_4348,N_3692,N_3320);
nor U4349 (N_4349,N_3778,N_3486);
xnor U4350 (N_4350,N_3131,N_3490);
or U4351 (N_4351,N_3908,N_3606);
xor U4352 (N_4352,N_3664,N_3348);
and U4353 (N_4353,N_3583,N_3480);
nand U4354 (N_4354,N_3624,N_3187);
nand U4355 (N_4355,N_3194,N_3555);
and U4356 (N_4356,N_3766,N_3087);
or U4357 (N_4357,N_3112,N_3847);
and U4358 (N_4358,N_3092,N_3907);
nor U4359 (N_4359,N_3714,N_3298);
and U4360 (N_4360,N_3275,N_3127);
and U4361 (N_4361,N_3119,N_3563);
and U4362 (N_4362,N_3770,N_3917);
nand U4363 (N_4363,N_3405,N_3715);
and U4364 (N_4364,N_3888,N_3232);
xnor U4365 (N_4365,N_3217,N_3223);
nor U4366 (N_4366,N_3438,N_3704);
nand U4367 (N_4367,N_3072,N_3469);
xor U4368 (N_4368,N_3645,N_3951);
nor U4369 (N_4369,N_3176,N_3353);
nand U4370 (N_4370,N_3494,N_3799);
nor U4371 (N_4371,N_3674,N_3950);
xor U4372 (N_4372,N_3435,N_3359);
nand U4373 (N_4373,N_3740,N_3572);
nor U4374 (N_4374,N_3183,N_3954);
nand U4375 (N_4375,N_3614,N_3512);
or U4376 (N_4376,N_3649,N_3156);
nor U4377 (N_4377,N_3081,N_3631);
and U4378 (N_4378,N_3314,N_3300);
or U4379 (N_4379,N_3430,N_3379);
or U4380 (N_4380,N_3387,N_3455);
nor U4381 (N_4381,N_3659,N_3946);
or U4382 (N_4382,N_3076,N_3195);
nand U4383 (N_4383,N_3419,N_3204);
xor U4384 (N_4384,N_3021,N_3873);
nand U4385 (N_4385,N_3633,N_3404);
nand U4386 (N_4386,N_3328,N_3549);
and U4387 (N_4387,N_3738,N_3525);
xor U4388 (N_4388,N_3981,N_3077);
xor U4389 (N_4389,N_3253,N_3909);
xnor U4390 (N_4390,N_3962,N_3141);
or U4391 (N_4391,N_3900,N_3707);
and U4392 (N_4392,N_3162,N_3400);
nand U4393 (N_4393,N_3820,N_3122);
xor U4394 (N_4394,N_3059,N_3516);
nor U4395 (N_4395,N_3105,N_3366);
xnor U4396 (N_4396,N_3887,N_3698);
xor U4397 (N_4397,N_3899,N_3351);
nor U4398 (N_4398,N_3229,N_3757);
and U4399 (N_4399,N_3611,N_3683);
nand U4400 (N_4400,N_3987,N_3099);
nand U4401 (N_4401,N_3277,N_3305);
or U4402 (N_4402,N_3053,N_3796);
and U4403 (N_4403,N_3732,N_3865);
and U4404 (N_4404,N_3124,N_3467);
nand U4405 (N_4405,N_3787,N_3456);
xnor U4406 (N_4406,N_3178,N_3846);
or U4407 (N_4407,N_3154,N_3869);
nor U4408 (N_4408,N_3782,N_3800);
nor U4409 (N_4409,N_3415,N_3928);
xor U4410 (N_4410,N_3368,N_3504);
xnor U4411 (N_4411,N_3741,N_3350);
or U4412 (N_4412,N_3289,N_3646);
and U4413 (N_4413,N_3803,N_3020);
or U4414 (N_4414,N_3246,N_3031);
and U4415 (N_4415,N_3961,N_3844);
nand U4416 (N_4416,N_3499,N_3902);
nand U4417 (N_4417,N_3001,N_3676);
or U4418 (N_4418,N_3508,N_3227);
xnor U4419 (N_4419,N_3032,N_3903);
nand U4420 (N_4420,N_3752,N_3308);
xor U4421 (N_4421,N_3185,N_3845);
nor U4422 (N_4422,N_3452,N_3543);
or U4423 (N_4423,N_3669,N_3597);
nand U4424 (N_4424,N_3861,N_3826);
nor U4425 (N_4425,N_3170,N_3166);
or U4426 (N_4426,N_3670,N_3487);
nor U4427 (N_4427,N_3850,N_3815);
nor U4428 (N_4428,N_3114,N_3548);
nor U4429 (N_4429,N_3975,N_3594);
xnor U4430 (N_4430,N_3586,N_3242);
nor U4431 (N_4431,N_3852,N_3061);
or U4432 (N_4432,N_3783,N_3086);
and U4433 (N_4433,N_3943,N_3057);
nor U4434 (N_4434,N_3965,N_3322);
nand U4435 (N_4435,N_3459,N_3213);
or U4436 (N_4436,N_3342,N_3745);
or U4437 (N_4437,N_3724,N_3947);
nand U4438 (N_4438,N_3967,N_3636);
or U4439 (N_4439,N_3505,N_3460);
nand U4440 (N_4440,N_3046,N_3362);
or U4441 (N_4441,N_3281,N_3654);
xnor U4442 (N_4442,N_3347,N_3357);
or U4443 (N_4443,N_3448,N_3007);
xor U4444 (N_4444,N_3039,N_3822);
nor U4445 (N_4445,N_3161,N_3871);
nor U4446 (N_4446,N_3769,N_3103);
nor U4447 (N_4447,N_3261,N_3660);
xnor U4448 (N_4448,N_3641,N_3576);
or U4449 (N_4449,N_3910,N_3336);
or U4450 (N_4450,N_3565,N_3608);
xnor U4451 (N_4451,N_3384,N_3028);
xnor U4452 (N_4452,N_3278,N_3018);
or U4453 (N_4453,N_3136,N_3306);
xnor U4454 (N_4454,N_3164,N_3953);
nor U4455 (N_4455,N_3395,N_3619);
nand U4456 (N_4456,N_3292,N_3923);
nand U4457 (N_4457,N_3142,N_3243);
xor U4458 (N_4458,N_3402,N_3226);
xor U4459 (N_4459,N_3791,N_3540);
nor U4460 (N_4460,N_3211,N_3615);
and U4461 (N_4461,N_3816,N_3785);
nand U4462 (N_4462,N_3476,N_3418);
nor U4463 (N_4463,N_3864,N_3356);
and U4464 (N_4464,N_3618,N_3638);
and U4465 (N_4465,N_3479,N_3317);
xnor U4466 (N_4466,N_3896,N_3737);
nor U4467 (N_4467,N_3588,N_3475);
nand U4468 (N_4468,N_3536,N_3625);
nor U4469 (N_4469,N_3358,N_3200);
and U4470 (N_4470,N_3533,N_3912);
nor U4471 (N_4471,N_3552,N_3721);
nor U4472 (N_4472,N_3209,N_3272);
or U4473 (N_4473,N_3140,N_3255);
xor U4474 (N_4474,N_3035,N_3889);
nor U4475 (N_4475,N_3662,N_3934);
xnor U4476 (N_4476,N_3388,N_3191);
or U4477 (N_4477,N_3000,N_3697);
nand U4478 (N_4478,N_3558,N_3440);
xnor U4479 (N_4479,N_3706,N_3433);
and U4480 (N_4480,N_3201,N_3157);
or U4481 (N_4481,N_3539,N_3600);
and U4482 (N_4482,N_3985,N_3677);
nand U4483 (N_4483,N_3403,N_3052);
xor U4484 (N_4484,N_3023,N_3672);
nor U4485 (N_4485,N_3988,N_3883);
nand U4486 (N_4486,N_3546,N_3436);
nor U4487 (N_4487,N_3798,N_3100);
xor U4488 (N_4488,N_3108,N_3222);
nor U4489 (N_4489,N_3047,N_3658);
nor U4490 (N_4490,N_3054,N_3143);
xnor U4491 (N_4491,N_3522,N_3948);
nor U4492 (N_4492,N_3175,N_3293);
nand U4493 (N_4493,N_3506,N_3144);
nand U4494 (N_4494,N_3569,N_3133);
and U4495 (N_4495,N_3678,N_3410);
nor U4496 (N_4496,N_3642,N_3612);
nand U4497 (N_4497,N_3566,N_3022);
and U4498 (N_4498,N_3085,N_3701);
or U4499 (N_4499,N_3339,N_3941);
nor U4500 (N_4500,N_3498,N_3672);
and U4501 (N_4501,N_3916,N_3239);
xnor U4502 (N_4502,N_3712,N_3492);
nor U4503 (N_4503,N_3617,N_3386);
and U4504 (N_4504,N_3606,N_3369);
and U4505 (N_4505,N_3775,N_3339);
xor U4506 (N_4506,N_3670,N_3076);
or U4507 (N_4507,N_3084,N_3798);
xnor U4508 (N_4508,N_3582,N_3541);
nor U4509 (N_4509,N_3604,N_3627);
nor U4510 (N_4510,N_3629,N_3792);
nand U4511 (N_4511,N_3355,N_3165);
or U4512 (N_4512,N_3505,N_3537);
nand U4513 (N_4513,N_3149,N_3712);
nor U4514 (N_4514,N_3582,N_3975);
nand U4515 (N_4515,N_3234,N_3098);
and U4516 (N_4516,N_3991,N_3442);
nor U4517 (N_4517,N_3293,N_3281);
or U4518 (N_4518,N_3045,N_3845);
nand U4519 (N_4519,N_3115,N_3416);
nor U4520 (N_4520,N_3591,N_3628);
or U4521 (N_4521,N_3588,N_3469);
nand U4522 (N_4522,N_3418,N_3946);
and U4523 (N_4523,N_3572,N_3270);
or U4524 (N_4524,N_3871,N_3271);
and U4525 (N_4525,N_3364,N_3961);
nor U4526 (N_4526,N_3711,N_3347);
xnor U4527 (N_4527,N_3499,N_3527);
or U4528 (N_4528,N_3777,N_3957);
and U4529 (N_4529,N_3772,N_3099);
nand U4530 (N_4530,N_3448,N_3186);
or U4531 (N_4531,N_3319,N_3629);
nand U4532 (N_4532,N_3250,N_3574);
nor U4533 (N_4533,N_3661,N_3780);
or U4534 (N_4534,N_3454,N_3786);
or U4535 (N_4535,N_3127,N_3932);
xnor U4536 (N_4536,N_3993,N_3970);
nand U4537 (N_4537,N_3791,N_3756);
nand U4538 (N_4538,N_3288,N_3088);
xor U4539 (N_4539,N_3848,N_3128);
xor U4540 (N_4540,N_3663,N_3764);
xor U4541 (N_4541,N_3998,N_3321);
nand U4542 (N_4542,N_3867,N_3689);
and U4543 (N_4543,N_3260,N_3635);
xnor U4544 (N_4544,N_3312,N_3317);
and U4545 (N_4545,N_3154,N_3029);
nand U4546 (N_4546,N_3771,N_3315);
or U4547 (N_4547,N_3200,N_3115);
nor U4548 (N_4548,N_3840,N_3572);
and U4549 (N_4549,N_3575,N_3651);
nand U4550 (N_4550,N_3212,N_3904);
nand U4551 (N_4551,N_3585,N_3467);
or U4552 (N_4552,N_3606,N_3957);
xnor U4553 (N_4553,N_3414,N_3682);
or U4554 (N_4554,N_3201,N_3296);
xor U4555 (N_4555,N_3107,N_3452);
nand U4556 (N_4556,N_3033,N_3113);
nor U4557 (N_4557,N_3741,N_3738);
nor U4558 (N_4558,N_3701,N_3140);
nor U4559 (N_4559,N_3571,N_3608);
nand U4560 (N_4560,N_3539,N_3174);
or U4561 (N_4561,N_3140,N_3315);
and U4562 (N_4562,N_3044,N_3574);
or U4563 (N_4563,N_3919,N_3184);
nand U4564 (N_4564,N_3509,N_3842);
xor U4565 (N_4565,N_3788,N_3191);
xnor U4566 (N_4566,N_3961,N_3187);
or U4567 (N_4567,N_3189,N_3041);
xnor U4568 (N_4568,N_3136,N_3816);
nor U4569 (N_4569,N_3638,N_3641);
or U4570 (N_4570,N_3850,N_3553);
or U4571 (N_4571,N_3971,N_3577);
xnor U4572 (N_4572,N_3340,N_3415);
or U4573 (N_4573,N_3387,N_3779);
or U4574 (N_4574,N_3501,N_3254);
xor U4575 (N_4575,N_3629,N_3839);
nor U4576 (N_4576,N_3266,N_3751);
nor U4577 (N_4577,N_3952,N_3002);
xnor U4578 (N_4578,N_3417,N_3694);
nor U4579 (N_4579,N_3495,N_3918);
and U4580 (N_4580,N_3815,N_3164);
and U4581 (N_4581,N_3239,N_3468);
and U4582 (N_4582,N_3550,N_3152);
xnor U4583 (N_4583,N_3917,N_3553);
nand U4584 (N_4584,N_3607,N_3842);
nand U4585 (N_4585,N_3996,N_3296);
and U4586 (N_4586,N_3791,N_3807);
xor U4587 (N_4587,N_3526,N_3881);
nor U4588 (N_4588,N_3040,N_3460);
or U4589 (N_4589,N_3524,N_3124);
and U4590 (N_4590,N_3554,N_3789);
nand U4591 (N_4591,N_3509,N_3089);
xor U4592 (N_4592,N_3268,N_3676);
nor U4593 (N_4593,N_3680,N_3927);
or U4594 (N_4594,N_3977,N_3732);
and U4595 (N_4595,N_3977,N_3274);
xor U4596 (N_4596,N_3111,N_3083);
nor U4597 (N_4597,N_3527,N_3238);
and U4598 (N_4598,N_3094,N_3646);
and U4599 (N_4599,N_3321,N_3310);
nor U4600 (N_4600,N_3992,N_3399);
nand U4601 (N_4601,N_3637,N_3708);
and U4602 (N_4602,N_3479,N_3603);
xor U4603 (N_4603,N_3614,N_3359);
and U4604 (N_4604,N_3931,N_3458);
nor U4605 (N_4605,N_3319,N_3488);
nand U4606 (N_4606,N_3516,N_3257);
xnor U4607 (N_4607,N_3124,N_3606);
or U4608 (N_4608,N_3393,N_3737);
xnor U4609 (N_4609,N_3086,N_3530);
nor U4610 (N_4610,N_3235,N_3604);
nand U4611 (N_4611,N_3125,N_3684);
or U4612 (N_4612,N_3358,N_3727);
nand U4613 (N_4613,N_3313,N_3564);
or U4614 (N_4614,N_3008,N_3403);
nor U4615 (N_4615,N_3973,N_3828);
xnor U4616 (N_4616,N_3518,N_3216);
nor U4617 (N_4617,N_3763,N_3381);
or U4618 (N_4618,N_3111,N_3865);
and U4619 (N_4619,N_3158,N_3083);
xnor U4620 (N_4620,N_3980,N_3617);
xnor U4621 (N_4621,N_3865,N_3684);
xnor U4622 (N_4622,N_3624,N_3271);
or U4623 (N_4623,N_3839,N_3610);
nand U4624 (N_4624,N_3248,N_3167);
and U4625 (N_4625,N_3374,N_3289);
and U4626 (N_4626,N_3983,N_3837);
and U4627 (N_4627,N_3188,N_3135);
nand U4628 (N_4628,N_3353,N_3941);
and U4629 (N_4629,N_3963,N_3012);
and U4630 (N_4630,N_3586,N_3813);
and U4631 (N_4631,N_3854,N_3981);
xnor U4632 (N_4632,N_3485,N_3444);
xnor U4633 (N_4633,N_3102,N_3211);
nor U4634 (N_4634,N_3122,N_3749);
nand U4635 (N_4635,N_3633,N_3564);
nand U4636 (N_4636,N_3946,N_3986);
and U4637 (N_4637,N_3095,N_3662);
and U4638 (N_4638,N_3157,N_3763);
or U4639 (N_4639,N_3105,N_3850);
nor U4640 (N_4640,N_3950,N_3456);
xnor U4641 (N_4641,N_3596,N_3311);
xor U4642 (N_4642,N_3448,N_3423);
nor U4643 (N_4643,N_3913,N_3809);
nand U4644 (N_4644,N_3385,N_3183);
xnor U4645 (N_4645,N_3616,N_3163);
or U4646 (N_4646,N_3338,N_3340);
or U4647 (N_4647,N_3422,N_3397);
or U4648 (N_4648,N_3870,N_3439);
or U4649 (N_4649,N_3292,N_3891);
xnor U4650 (N_4650,N_3444,N_3982);
nand U4651 (N_4651,N_3635,N_3426);
nand U4652 (N_4652,N_3094,N_3493);
nor U4653 (N_4653,N_3701,N_3493);
nor U4654 (N_4654,N_3880,N_3931);
and U4655 (N_4655,N_3717,N_3796);
or U4656 (N_4656,N_3068,N_3339);
nor U4657 (N_4657,N_3325,N_3311);
nand U4658 (N_4658,N_3800,N_3375);
xnor U4659 (N_4659,N_3499,N_3242);
nand U4660 (N_4660,N_3065,N_3217);
xor U4661 (N_4661,N_3333,N_3217);
nand U4662 (N_4662,N_3664,N_3642);
and U4663 (N_4663,N_3269,N_3919);
or U4664 (N_4664,N_3626,N_3740);
nand U4665 (N_4665,N_3983,N_3010);
xor U4666 (N_4666,N_3138,N_3418);
nor U4667 (N_4667,N_3067,N_3923);
and U4668 (N_4668,N_3509,N_3497);
and U4669 (N_4669,N_3655,N_3658);
nor U4670 (N_4670,N_3229,N_3301);
or U4671 (N_4671,N_3491,N_3219);
or U4672 (N_4672,N_3418,N_3896);
xnor U4673 (N_4673,N_3625,N_3400);
or U4674 (N_4674,N_3913,N_3298);
nand U4675 (N_4675,N_3589,N_3919);
or U4676 (N_4676,N_3250,N_3936);
nor U4677 (N_4677,N_3234,N_3984);
and U4678 (N_4678,N_3303,N_3150);
and U4679 (N_4679,N_3598,N_3835);
nand U4680 (N_4680,N_3946,N_3172);
nor U4681 (N_4681,N_3637,N_3664);
and U4682 (N_4682,N_3702,N_3271);
nand U4683 (N_4683,N_3865,N_3782);
nor U4684 (N_4684,N_3078,N_3185);
nand U4685 (N_4685,N_3281,N_3198);
nor U4686 (N_4686,N_3518,N_3122);
nor U4687 (N_4687,N_3052,N_3244);
or U4688 (N_4688,N_3659,N_3440);
nand U4689 (N_4689,N_3887,N_3620);
and U4690 (N_4690,N_3874,N_3250);
nor U4691 (N_4691,N_3233,N_3779);
and U4692 (N_4692,N_3955,N_3683);
nand U4693 (N_4693,N_3592,N_3939);
nor U4694 (N_4694,N_3844,N_3126);
nor U4695 (N_4695,N_3369,N_3168);
or U4696 (N_4696,N_3624,N_3839);
xor U4697 (N_4697,N_3422,N_3083);
and U4698 (N_4698,N_3618,N_3647);
nor U4699 (N_4699,N_3966,N_3152);
or U4700 (N_4700,N_3787,N_3413);
and U4701 (N_4701,N_3519,N_3080);
nand U4702 (N_4702,N_3026,N_3472);
nor U4703 (N_4703,N_3920,N_3168);
or U4704 (N_4704,N_3788,N_3458);
and U4705 (N_4705,N_3836,N_3175);
xor U4706 (N_4706,N_3513,N_3262);
and U4707 (N_4707,N_3182,N_3395);
and U4708 (N_4708,N_3950,N_3701);
nand U4709 (N_4709,N_3450,N_3239);
or U4710 (N_4710,N_3773,N_3770);
xor U4711 (N_4711,N_3547,N_3210);
xnor U4712 (N_4712,N_3048,N_3187);
nor U4713 (N_4713,N_3903,N_3447);
or U4714 (N_4714,N_3559,N_3638);
nor U4715 (N_4715,N_3178,N_3858);
or U4716 (N_4716,N_3212,N_3925);
or U4717 (N_4717,N_3666,N_3482);
nand U4718 (N_4718,N_3429,N_3378);
nand U4719 (N_4719,N_3480,N_3595);
nor U4720 (N_4720,N_3954,N_3408);
nand U4721 (N_4721,N_3691,N_3500);
nand U4722 (N_4722,N_3144,N_3236);
nor U4723 (N_4723,N_3507,N_3826);
and U4724 (N_4724,N_3757,N_3832);
and U4725 (N_4725,N_3197,N_3693);
nor U4726 (N_4726,N_3512,N_3032);
nand U4727 (N_4727,N_3562,N_3863);
nor U4728 (N_4728,N_3905,N_3752);
nand U4729 (N_4729,N_3400,N_3940);
and U4730 (N_4730,N_3733,N_3518);
nand U4731 (N_4731,N_3880,N_3128);
xnor U4732 (N_4732,N_3599,N_3193);
nand U4733 (N_4733,N_3693,N_3940);
and U4734 (N_4734,N_3413,N_3168);
nand U4735 (N_4735,N_3295,N_3827);
xor U4736 (N_4736,N_3982,N_3798);
nand U4737 (N_4737,N_3442,N_3107);
or U4738 (N_4738,N_3236,N_3806);
xnor U4739 (N_4739,N_3559,N_3978);
nor U4740 (N_4740,N_3698,N_3170);
and U4741 (N_4741,N_3279,N_3486);
and U4742 (N_4742,N_3949,N_3237);
or U4743 (N_4743,N_3407,N_3193);
and U4744 (N_4744,N_3230,N_3847);
or U4745 (N_4745,N_3857,N_3847);
and U4746 (N_4746,N_3658,N_3996);
xor U4747 (N_4747,N_3813,N_3854);
xnor U4748 (N_4748,N_3884,N_3551);
nand U4749 (N_4749,N_3871,N_3796);
and U4750 (N_4750,N_3645,N_3774);
xor U4751 (N_4751,N_3523,N_3120);
nand U4752 (N_4752,N_3367,N_3414);
and U4753 (N_4753,N_3624,N_3575);
xor U4754 (N_4754,N_3945,N_3757);
and U4755 (N_4755,N_3311,N_3100);
and U4756 (N_4756,N_3172,N_3907);
nand U4757 (N_4757,N_3784,N_3115);
or U4758 (N_4758,N_3100,N_3642);
nor U4759 (N_4759,N_3981,N_3087);
xnor U4760 (N_4760,N_3812,N_3209);
xnor U4761 (N_4761,N_3303,N_3734);
nor U4762 (N_4762,N_3758,N_3898);
nor U4763 (N_4763,N_3892,N_3702);
nand U4764 (N_4764,N_3667,N_3526);
nand U4765 (N_4765,N_3263,N_3695);
nand U4766 (N_4766,N_3093,N_3378);
xnor U4767 (N_4767,N_3774,N_3474);
nand U4768 (N_4768,N_3000,N_3866);
xor U4769 (N_4769,N_3894,N_3320);
nor U4770 (N_4770,N_3886,N_3654);
nand U4771 (N_4771,N_3904,N_3065);
xnor U4772 (N_4772,N_3227,N_3582);
and U4773 (N_4773,N_3854,N_3616);
xnor U4774 (N_4774,N_3518,N_3745);
or U4775 (N_4775,N_3877,N_3733);
nor U4776 (N_4776,N_3500,N_3832);
nand U4777 (N_4777,N_3375,N_3920);
or U4778 (N_4778,N_3971,N_3666);
xor U4779 (N_4779,N_3273,N_3080);
nand U4780 (N_4780,N_3682,N_3565);
xnor U4781 (N_4781,N_3734,N_3234);
and U4782 (N_4782,N_3412,N_3466);
and U4783 (N_4783,N_3053,N_3588);
xnor U4784 (N_4784,N_3141,N_3545);
nand U4785 (N_4785,N_3692,N_3777);
nand U4786 (N_4786,N_3579,N_3102);
nand U4787 (N_4787,N_3735,N_3197);
and U4788 (N_4788,N_3771,N_3835);
or U4789 (N_4789,N_3487,N_3325);
and U4790 (N_4790,N_3950,N_3578);
nor U4791 (N_4791,N_3252,N_3485);
or U4792 (N_4792,N_3460,N_3077);
or U4793 (N_4793,N_3672,N_3952);
xor U4794 (N_4794,N_3411,N_3598);
and U4795 (N_4795,N_3361,N_3540);
nand U4796 (N_4796,N_3844,N_3903);
nand U4797 (N_4797,N_3642,N_3814);
nand U4798 (N_4798,N_3832,N_3696);
and U4799 (N_4799,N_3111,N_3158);
and U4800 (N_4800,N_3988,N_3004);
xor U4801 (N_4801,N_3904,N_3726);
xnor U4802 (N_4802,N_3174,N_3882);
nor U4803 (N_4803,N_3005,N_3750);
nor U4804 (N_4804,N_3763,N_3987);
nand U4805 (N_4805,N_3558,N_3109);
xnor U4806 (N_4806,N_3060,N_3085);
or U4807 (N_4807,N_3393,N_3360);
nor U4808 (N_4808,N_3696,N_3916);
and U4809 (N_4809,N_3352,N_3134);
and U4810 (N_4810,N_3299,N_3148);
nor U4811 (N_4811,N_3372,N_3215);
nand U4812 (N_4812,N_3103,N_3640);
and U4813 (N_4813,N_3351,N_3443);
xnor U4814 (N_4814,N_3753,N_3785);
or U4815 (N_4815,N_3711,N_3340);
xor U4816 (N_4816,N_3387,N_3440);
and U4817 (N_4817,N_3671,N_3201);
or U4818 (N_4818,N_3077,N_3119);
nor U4819 (N_4819,N_3896,N_3505);
nor U4820 (N_4820,N_3205,N_3634);
nor U4821 (N_4821,N_3869,N_3341);
nor U4822 (N_4822,N_3544,N_3608);
nand U4823 (N_4823,N_3016,N_3110);
and U4824 (N_4824,N_3600,N_3496);
nor U4825 (N_4825,N_3695,N_3765);
nand U4826 (N_4826,N_3565,N_3674);
nor U4827 (N_4827,N_3429,N_3778);
nand U4828 (N_4828,N_3828,N_3071);
or U4829 (N_4829,N_3475,N_3034);
and U4830 (N_4830,N_3912,N_3282);
or U4831 (N_4831,N_3116,N_3794);
and U4832 (N_4832,N_3174,N_3508);
xor U4833 (N_4833,N_3142,N_3479);
nor U4834 (N_4834,N_3160,N_3873);
nand U4835 (N_4835,N_3316,N_3337);
and U4836 (N_4836,N_3245,N_3164);
and U4837 (N_4837,N_3980,N_3131);
and U4838 (N_4838,N_3351,N_3754);
xnor U4839 (N_4839,N_3668,N_3839);
xor U4840 (N_4840,N_3968,N_3976);
nor U4841 (N_4841,N_3940,N_3184);
nor U4842 (N_4842,N_3852,N_3029);
and U4843 (N_4843,N_3734,N_3208);
or U4844 (N_4844,N_3055,N_3512);
or U4845 (N_4845,N_3598,N_3775);
and U4846 (N_4846,N_3806,N_3708);
or U4847 (N_4847,N_3186,N_3370);
or U4848 (N_4848,N_3111,N_3549);
or U4849 (N_4849,N_3171,N_3828);
or U4850 (N_4850,N_3422,N_3849);
or U4851 (N_4851,N_3040,N_3372);
nand U4852 (N_4852,N_3756,N_3574);
and U4853 (N_4853,N_3371,N_3512);
or U4854 (N_4854,N_3439,N_3721);
nor U4855 (N_4855,N_3191,N_3928);
xor U4856 (N_4856,N_3090,N_3741);
and U4857 (N_4857,N_3744,N_3015);
and U4858 (N_4858,N_3280,N_3548);
xor U4859 (N_4859,N_3815,N_3684);
xnor U4860 (N_4860,N_3169,N_3828);
and U4861 (N_4861,N_3702,N_3768);
nand U4862 (N_4862,N_3451,N_3472);
or U4863 (N_4863,N_3451,N_3210);
nand U4864 (N_4864,N_3402,N_3801);
and U4865 (N_4865,N_3330,N_3227);
nor U4866 (N_4866,N_3579,N_3050);
nand U4867 (N_4867,N_3449,N_3601);
nand U4868 (N_4868,N_3761,N_3423);
nor U4869 (N_4869,N_3810,N_3078);
nand U4870 (N_4870,N_3707,N_3070);
and U4871 (N_4871,N_3084,N_3445);
nor U4872 (N_4872,N_3919,N_3731);
nor U4873 (N_4873,N_3972,N_3534);
xor U4874 (N_4874,N_3254,N_3363);
xor U4875 (N_4875,N_3700,N_3088);
xnor U4876 (N_4876,N_3326,N_3649);
xnor U4877 (N_4877,N_3747,N_3569);
nor U4878 (N_4878,N_3975,N_3632);
xnor U4879 (N_4879,N_3435,N_3559);
nor U4880 (N_4880,N_3377,N_3252);
xnor U4881 (N_4881,N_3872,N_3690);
or U4882 (N_4882,N_3389,N_3394);
xnor U4883 (N_4883,N_3987,N_3602);
xnor U4884 (N_4884,N_3779,N_3308);
or U4885 (N_4885,N_3750,N_3525);
nor U4886 (N_4886,N_3920,N_3112);
nor U4887 (N_4887,N_3374,N_3353);
and U4888 (N_4888,N_3296,N_3208);
or U4889 (N_4889,N_3263,N_3338);
nor U4890 (N_4890,N_3574,N_3127);
and U4891 (N_4891,N_3693,N_3894);
xnor U4892 (N_4892,N_3055,N_3167);
or U4893 (N_4893,N_3166,N_3206);
and U4894 (N_4894,N_3586,N_3915);
or U4895 (N_4895,N_3156,N_3004);
xnor U4896 (N_4896,N_3502,N_3381);
nand U4897 (N_4897,N_3234,N_3175);
nor U4898 (N_4898,N_3503,N_3756);
nand U4899 (N_4899,N_3563,N_3376);
or U4900 (N_4900,N_3495,N_3048);
nand U4901 (N_4901,N_3875,N_3251);
xnor U4902 (N_4902,N_3693,N_3835);
xor U4903 (N_4903,N_3740,N_3610);
and U4904 (N_4904,N_3443,N_3896);
or U4905 (N_4905,N_3439,N_3893);
and U4906 (N_4906,N_3242,N_3598);
xor U4907 (N_4907,N_3828,N_3275);
and U4908 (N_4908,N_3456,N_3110);
nor U4909 (N_4909,N_3463,N_3623);
or U4910 (N_4910,N_3056,N_3551);
or U4911 (N_4911,N_3685,N_3211);
xor U4912 (N_4912,N_3101,N_3238);
nand U4913 (N_4913,N_3770,N_3504);
nor U4914 (N_4914,N_3890,N_3337);
and U4915 (N_4915,N_3787,N_3808);
nand U4916 (N_4916,N_3284,N_3235);
or U4917 (N_4917,N_3638,N_3577);
and U4918 (N_4918,N_3910,N_3036);
nor U4919 (N_4919,N_3329,N_3446);
xor U4920 (N_4920,N_3267,N_3883);
nor U4921 (N_4921,N_3802,N_3351);
nor U4922 (N_4922,N_3729,N_3368);
nor U4923 (N_4923,N_3975,N_3686);
or U4924 (N_4924,N_3028,N_3231);
nand U4925 (N_4925,N_3196,N_3371);
or U4926 (N_4926,N_3598,N_3858);
or U4927 (N_4927,N_3954,N_3779);
and U4928 (N_4928,N_3007,N_3193);
or U4929 (N_4929,N_3175,N_3263);
nor U4930 (N_4930,N_3724,N_3092);
xor U4931 (N_4931,N_3926,N_3215);
or U4932 (N_4932,N_3482,N_3009);
or U4933 (N_4933,N_3909,N_3394);
or U4934 (N_4934,N_3450,N_3894);
nor U4935 (N_4935,N_3593,N_3742);
and U4936 (N_4936,N_3847,N_3047);
nor U4937 (N_4937,N_3012,N_3156);
xor U4938 (N_4938,N_3302,N_3652);
xor U4939 (N_4939,N_3415,N_3216);
nand U4940 (N_4940,N_3002,N_3930);
nor U4941 (N_4941,N_3770,N_3808);
or U4942 (N_4942,N_3319,N_3158);
nor U4943 (N_4943,N_3860,N_3343);
xor U4944 (N_4944,N_3565,N_3238);
and U4945 (N_4945,N_3691,N_3095);
xnor U4946 (N_4946,N_3094,N_3072);
xnor U4947 (N_4947,N_3299,N_3472);
and U4948 (N_4948,N_3019,N_3587);
nand U4949 (N_4949,N_3322,N_3952);
nor U4950 (N_4950,N_3009,N_3682);
nor U4951 (N_4951,N_3958,N_3752);
nand U4952 (N_4952,N_3469,N_3392);
nor U4953 (N_4953,N_3564,N_3237);
xor U4954 (N_4954,N_3765,N_3748);
nand U4955 (N_4955,N_3022,N_3405);
and U4956 (N_4956,N_3713,N_3279);
xnor U4957 (N_4957,N_3919,N_3909);
xor U4958 (N_4958,N_3369,N_3390);
or U4959 (N_4959,N_3949,N_3588);
xor U4960 (N_4960,N_3766,N_3689);
or U4961 (N_4961,N_3525,N_3085);
xnor U4962 (N_4962,N_3084,N_3400);
nor U4963 (N_4963,N_3764,N_3364);
xnor U4964 (N_4964,N_3712,N_3387);
nand U4965 (N_4965,N_3004,N_3652);
and U4966 (N_4966,N_3045,N_3973);
nand U4967 (N_4967,N_3528,N_3418);
or U4968 (N_4968,N_3835,N_3767);
or U4969 (N_4969,N_3930,N_3488);
nor U4970 (N_4970,N_3397,N_3328);
nand U4971 (N_4971,N_3395,N_3481);
nand U4972 (N_4972,N_3975,N_3647);
or U4973 (N_4973,N_3357,N_3855);
nand U4974 (N_4974,N_3008,N_3871);
or U4975 (N_4975,N_3894,N_3015);
nor U4976 (N_4976,N_3379,N_3578);
xnor U4977 (N_4977,N_3913,N_3794);
nand U4978 (N_4978,N_3727,N_3254);
xor U4979 (N_4979,N_3174,N_3808);
and U4980 (N_4980,N_3888,N_3447);
xor U4981 (N_4981,N_3576,N_3130);
nor U4982 (N_4982,N_3195,N_3697);
or U4983 (N_4983,N_3320,N_3717);
xnor U4984 (N_4984,N_3081,N_3148);
or U4985 (N_4985,N_3803,N_3173);
nor U4986 (N_4986,N_3200,N_3481);
nor U4987 (N_4987,N_3598,N_3328);
and U4988 (N_4988,N_3082,N_3479);
nand U4989 (N_4989,N_3400,N_3403);
or U4990 (N_4990,N_3307,N_3860);
xor U4991 (N_4991,N_3615,N_3899);
nor U4992 (N_4992,N_3884,N_3296);
nand U4993 (N_4993,N_3374,N_3451);
nand U4994 (N_4994,N_3420,N_3075);
or U4995 (N_4995,N_3106,N_3535);
nand U4996 (N_4996,N_3875,N_3168);
and U4997 (N_4997,N_3701,N_3832);
nor U4998 (N_4998,N_3364,N_3401);
nor U4999 (N_4999,N_3427,N_3998);
or U5000 (N_5000,N_4105,N_4810);
and U5001 (N_5001,N_4012,N_4997);
and U5002 (N_5002,N_4566,N_4995);
nor U5003 (N_5003,N_4272,N_4956);
xnor U5004 (N_5004,N_4660,N_4923);
and U5005 (N_5005,N_4268,N_4366);
or U5006 (N_5006,N_4223,N_4982);
or U5007 (N_5007,N_4229,N_4665);
xor U5008 (N_5008,N_4168,N_4432);
nor U5009 (N_5009,N_4795,N_4263);
xnor U5010 (N_5010,N_4902,N_4716);
nor U5011 (N_5011,N_4865,N_4221);
or U5012 (N_5012,N_4637,N_4866);
and U5013 (N_5013,N_4149,N_4319);
xnor U5014 (N_5014,N_4226,N_4671);
nor U5015 (N_5015,N_4050,N_4393);
or U5016 (N_5016,N_4843,N_4502);
nor U5017 (N_5017,N_4893,N_4008);
nor U5018 (N_5018,N_4046,N_4495);
nor U5019 (N_5019,N_4531,N_4610);
nor U5020 (N_5020,N_4621,N_4792);
and U5021 (N_5021,N_4453,N_4853);
nor U5022 (N_5022,N_4498,N_4636);
nor U5023 (N_5023,N_4712,N_4753);
xnor U5024 (N_5024,N_4897,N_4697);
xor U5025 (N_5025,N_4499,N_4294);
xor U5026 (N_5026,N_4324,N_4891);
or U5027 (N_5027,N_4929,N_4405);
nand U5028 (N_5028,N_4835,N_4051);
nor U5029 (N_5029,N_4774,N_4447);
nor U5030 (N_5030,N_4337,N_4348);
nand U5031 (N_5031,N_4979,N_4068);
or U5032 (N_5032,N_4501,N_4157);
and U5033 (N_5033,N_4336,N_4900);
xor U5034 (N_5034,N_4738,N_4202);
xor U5035 (N_5035,N_4609,N_4555);
nand U5036 (N_5036,N_4536,N_4957);
nand U5037 (N_5037,N_4075,N_4988);
nand U5038 (N_5038,N_4392,N_4074);
and U5039 (N_5039,N_4854,N_4707);
xor U5040 (N_5040,N_4573,N_4399);
nand U5041 (N_5041,N_4426,N_4276);
nand U5042 (N_5042,N_4408,N_4641);
nor U5043 (N_5043,N_4187,N_4062);
nand U5044 (N_5044,N_4483,N_4986);
nor U5045 (N_5045,N_4166,N_4941);
or U5046 (N_5046,N_4819,N_4984);
or U5047 (N_5047,N_4106,N_4603);
nand U5048 (N_5048,N_4242,N_4706);
nand U5049 (N_5049,N_4072,N_4925);
xor U5050 (N_5050,N_4734,N_4703);
xor U5051 (N_5051,N_4846,N_4670);
xnor U5052 (N_5052,N_4653,N_4232);
nor U5053 (N_5053,N_4812,N_4701);
nor U5054 (N_5054,N_4484,N_4086);
and U5055 (N_5055,N_4595,N_4264);
xnor U5056 (N_5056,N_4092,N_4119);
and U5057 (N_5057,N_4506,N_4873);
and U5058 (N_5058,N_4145,N_4201);
nand U5059 (N_5059,N_4411,N_4369);
and U5060 (N_5060,N_4427,N_4619);
or U5061 (N_5061,N_4236,N_4698);
nand U5062 (N_5062,N_4615,N_4761);
and U5063 (N_5063,N_4919,N_4554);
or U5064 (N_5064,N_4347,N_4474);
xnor U5065 (N_5065,N_4765,N_4974);
nand U5066 (N_5066,N_4602,N_4546);
and U5067 (N_5067,N_4173,N_4401);
and U5068 (N_5068,N_4255,N_4332);
nor U5069 (N_5069,N_4262,N_4683);
nor U5070 (N_5070,N_4564,N_4446);
or U5071 (N_5071,N_4133,N_4815);
or U5072 (N_5072,N_4083,N_4917);
or U5073 (N_5073,N_4890,N_4633);
and U5074 (N_5074,N_4673,N_4420);
and U5075 (N_5075,N_4850,N_4174);
nand U5076 (N_5076,N_4104,N_4384);
nor U5077 (N_5077,N_4151,N_4318);
or U5078 (N_5078,N_4482,N_4307);
xnor U5079 (N_5079,N_4936,N_4958);
xor U5080 (N_5080,N_4030,N_4049);
nand U5081 (N_5081,N_4311,N_4213);
or U5082 (N_5082,N_4584,N_4343);
xor U5083 (N_5083,N_4487,N_4711);
or U5084 (N_5084,N_4772,N_4274);
xor U5085 (N_5085,N_4693,N_4129);
xnor U5086 (N_5086,N_4597,N_4436);
nand U5087 (N_5087,N_4461,N_4558);
or U5088 (N_5088,N_4358,N_4857);
and U5089 (N_5089,N_4305,N_4212);
nor U5090 (N_5090,N_4723,N_4414);
or U5091 (N_5091,N_4052,N_4048);
nor U5092 (N_5092,N_4109,N_4991);
nor U5093 (N_5093,N_4450,N_4136);
xnor U5094 (N_5094,N_4870,N_4651);
nand U5095 (N_5095,N_4728,N_4493);
nor U5096 (N_5096,N_4837,N_4375);
nand U5097 (N_5097,N_4422,N_4057);
and U5098 (N_5098,N_4704,N_4019);
nand U5099 (N_5099,N_4198,N_4605);
or U5100 (N_5100,N_4195,N_4515);
or U5101 (N_5101,N_4926,N_4672);
nor U5102 (N_5102,N_4472,N_4530);
and U5103 (N_5103,N_4029,N_4100);
and U5104 (N_5104,N_4516,N_4117);
nand U5105 (N_5105,N_4503,N_4282);
nor U5106 (N_5106,N_4994,N_4175);
xnor U5107 (N_5107,N_4244,N_4519);
nor U5108 (N_5108,N_4759,N_4060);
nand U5109 (N_5109,N_4070,N_4120);
or U5110 (N_5110,N_4055,N_4667);
nor U5111 (N_5111,N_4628,N_4940);
and U5112 (N_5112,N_4257,N_4203);
xor U5113 (N_5113,N_4218,N_4485);
nand U5114 (N_5114,N_4512,N_4038);
or U5115 (N_5115,N_4763,N_4180);
nand U5116 (N_5116,N_4581,N_4700);
and U5117 (N_5117,N_4959,N_4888);
nand U5118 (N_5118,N_4007,N_4549);
or U5119 (N_5119,N_4669,N_4658);
nor U5120 (N_5120,N_4248,N_4177);
and U5121 (N_5121,N_4833,N_4981);
or U5122 (N_5122,N_4002,N_4334);
or U5123 (N_5123,N_4063,N_4799);
and U5124 (N_5124,N_4785,N_4088);
xnor U5125 (N_5125,N_4924,N_4190);
and U5126 (N_5126,N_4378,N_4783);
nor U5127 (N_5127,N_4879,N_4517);
and U5128 (N_5128,N_4552,N_4126);
or U5129 (N_5129,N_4421,N_4178);
and U5130 (N_5130,N_4372,N_4972);
and U5131 (N_5131,N_4323,N_4845);
nor U5132 (N_5132,N_4777,N_4804);
nand U5133 (N_5133,N_4277,N_4301);
or U5134 (N_5134,N_4451,N_4035);
nand U5135 (N_5135,N_4026,N_4599);
nand U5136 (N_5136,N_4877,N_4389);
nor U5137 (N_5137,N_4524,N_4749);
nand U5138 (N_5138,N_4113,N_4322);
and U5139 (N_5139,N_4831,N_4655);
nor U5140 (N_5140,N_4607,N_4067);
and U5141 (N_5141,N_4526,N_4565);
xnor U5142 (N_5142,N_4497,N_4782);
xor U5143 (N_5143,N_4338,N_4954);
nand U5144 (N_5144,N_4085,N_4488);
nand U5145 (N_5145,N_4541,N_4842);
or U5146 (N_5146,N_4130,N_4741);
or U5147 (N_5147,N_4646,N_4945);
nand U5148 (N_5148,N_4886,N_4153);
or U5149 (N_5149,N_4027,N_4654);
and U5150 (N_5150,N_4752,N_4754);
nand U5151 (N_5151,N_4718,N_4054);
nand U5152 (N_5152,N_4793,N_4736);
nand U5153 (N_5153,N_4556,N_4714);
xor U5154 (N_5154,N_4836,N_4989);
or U5155 (N_5155,N_4234,N_4569);
or U5156 (N_5156,N_4813,N_4118);
nor U5157 (N_5157,N_4943,N_4518);
xor U5158 (N_5158,N_4477,N_4528);
nand U5159 (N_5159,N_4587,N_4437);
and U5160 (N_5160,N_4222,N_4289);
nor U5161 (N_5161,N_4797,N_4321);
xnor U5162 (N_5162,N_4768,N_4912);
nand U5163 (N_5163,N_4508,N_4589);
xnor U5164 (N_5164,N_4814,N_4454);
nand U5165 (N_5165,N_4056,N_4790);
nand U5166 (N_5166,N_4639,N_4333);
and U5167 (N_5167,N_4844,N_4791);
nand U5168 (N_5168,N_4722,N_4416);
or U5169 (N_5169,N_4039,N_4542);
nor U5170 (N_5170,N_4152,N_4364);
or U5171 (N_5171,N_4380,N_4439);
and U5172 (N_5172,N_4598,N_4291);
nand U5173 (N_5173,N_4486,N_4457);
and U5174 (N_5174,N_4823,N_4143);
or U5175 (N_5175,N_4188,N_4681);
xnor U5176 (N_5176,N_4987,N_4847);
or U5177 (N_5177,N_4458,N_4720);
and U5178 (N_5178,N_4928,N_4871);
xor U5179 (N_5179,N_4832,N_4801);
nor U5180 (N_5180,N_4861,N_4095);
or U5181 (N_5181,N_4424,N_4579);
or U5182 (N_5182,N_4544,N_4182);
nor U5183 (N_5183,N_4507,N_4043);
and U5184 (N_5184,N_4135,N_4583);
nand U5185 (N_5185,N_4121,N_4227);
xnor U5186 (N_5186,N_4976,N_4748);
or U5187 (N_5187,N_4971,N_4396);
nor U5188 (N_5188,N_4356,N_4031);
nor U5189 (N_5189,N_4370,N_4675);
or U5190 (N_5190,N_4826,N_4586);
and U5191 (N_5191,N_4538,N_4894);
or U5192 (N_5192,N_4081,N_4076);
nor U5193 (N_5193,N_4381,N_4059);
and U5194 (N_5194,N_4295,N_4429);
and U5195 (N_5195,N_4539,N_4725);
and U5196 (N_5196,N_4390,N_4361);
xnor U5197 (N_5197,N_4668,N_4529);
and U5198 (N_5198,N_4445,N_4091);
nand U5199 (N_5199,N_4908,N_4317);
or U5200 (N_5200,N_4192,N_4131);
and U5201 (N_5201,N_4946,N_4612);
xor U5202 (N_5202,N_4443,N_4339);
xor U5203 (N_5203,N_4470,N_4617);
nand U5204 (N_5204,N_4200,N_4535);
or U5205 (N_5205,N_4138,N_4514);
xor U5206 (N_5206,N_4596,N_4025);
or U5207 (N_5207,N_4137,N_4985);
nand U5208 (N_5208,N_4481,N_4721);
or U5209 (N_5209,N_4601,N_4841);
xnor U5210 (N_5210,N_4652,N_4727);
and U5211 (N_5211,N_4090,N_4839);
and U5212 (N_5212,N_4998,N_4073);
nor U5213 (N_5213,N_4357,N_4112);
nor U5214 (N_5214,N_4314,N_4116);
xnor U5215 (N_5215,N_4139,N_4872);
nor U5216 (N_5216,N_4860,N_4513);
and U5217 (N_5217,N_4868,N_4690);
or U5218 (N_5218,N_4699,N_4309);
nand U5219 (N_5219,N_4648,N_4071);
xnor U5220 (N_5220,N_4563,N_4330);
and U5221 (N_5221,N_4258,N_4694);
nand U5222 (N_5222,N_4623,N_4293);
and U5223 (N_5223,N_4830,N_4757);
nand U5224 (N_5224,N_4363,N_4160);
xor U5225 (N_5225,N_4983,N_4822);
or U5226 (N_5226,N_4036,N_4476);
nor U5227 (N_5227,N_4540,N_4292);
nand U5228 (N_5228,N_4433,N_4775);
and U5229 (N_5229,N_4124,N_4034);
nor U5230 (N_5230,N_4183,N_4903);
and U5231 (N_5231,N_4467,N_4764);
and U5232 (N_5232,N_4883,N_4313);
nand U5233 (N_5233,N_4172,N_4942);
and U5234 (N_5234,N_4875,N_4933);
xor U5235 (N_5235,N_4395,N_4550);
nor U5236 (N_5236,N_4171,N_4354);
and U5237 (N_5237,N_4820,N_4779);
and U5238 (N_5238,N_4993,N_4614);
xnor U5239 (N_5239,N_4093,N_4110);
xor U5240 (N_5240,N_4645,N_4918);
xor U5241 (N_5241,N_4448,N_4931);
nand U5242 (N_5242,N_4144,N_4053);
or U5243 (N_5243,N_4280,N_4922);
or U5244 (N_5244,N_4527,N_4973);
xor U5245 (N_5245,N_4838,N_4352);
or U5246 (N_5246,N_4570,N_4297);
or U5247 (N_5247,N_4000,N_4613);
or U5248 (N_5248,N_4388,N_4800);
and U5249 (N_5249,N_4409,N_4927);
nand U5250 (N_5250,N_4456,N_4691);
xor U5251 (N_5251,N_4231,N_4150);
nand U5252 (N_5252,N_4729,N_4878);
and U5253 (N_5253,N_4909,N_4705);
xnor U5254 (N_5254,N_4626,N_4308);
nand U5255 (N_5255,N_4310,N_4266);
or U5256 (N_5256,N_4784,N_4325);
nor U5257 (N_5257,N_4851,N_4629);
nand U5258 (N_5258,N_4215,N_4967);
or U5259 (N_5259,N_4678,N_4193);
and U5260 (N_5260,N_4045,N_4125);
and U5261 (N_5261,N_4904,N_4089);
nor U5262 (N_5262,N_4913,N_4096);
nor U5263 (N_5263,N_4661,N_4164);
nor U5264 (N_5264,N_4638,N_4811);
or U5265 (N_5265,N_4199,N_4440);
or U5266 (N_5266,N_4733,N_4462);
xnor U5267 (N_5267,N_4735,N_4802);
nand U5268 (N_5268,N_4312,N_4907);
or U5269 (N_5269,N_4270,N_4999);
xor U5270 (N_5270,N_4786,N_4147);
or U5271 (N_5271,N_4859,N_4659);
xor U5272 (N_5272,N_4134,N_4079);
nand U5273 (N_5273,N_4058,N_4666);
nand U5274 (N_5274,N_4141,N_4478);
nand U5275 (N_5275,N_4047,N_4480);
and U5276 (N_5276,N_4769,N_4186);
xor U5277 (N_5277,N_4568,N_4162);
nor U5278 (N_5278,N_4750,N_4037);
or U5279 (N_5279,N_4575,N_4024);
nor U5280 (N_5280,N_4856,N_4934);
nor U5281 (N_5281,N_4821,N_4377);
nand U5282 (N_5282,N_4961,N_4600);
or U5283 (N_5283,N_4287,N_4858);
nor U5284 (N_5284,N_4567,N_4340);
nand U5285 (N_5285,N_4680,N_4169);
nor U5286 (N_5286,N_4158,N_4015);
or U5287 (N_5287,N_4737,N_4165);
nor U5288 (N_5288,N_4402,N_4867);
nor U5289 (N_5289,N_4417,N_4385);
or U5290 (N_5290,N_4726,N_4335);
xnor U5291 (N_5291,N_4228,N_4884);
and U5292 (N_5292,N_4649,N_4852);
nand U5293 (N_5293,N_4561,N_4241);
nor U5294 (N_5294,N_4465,N_4816);
and U5295 (N_5295,N_4953,N_4018);
nor U5296 (N_5296,N_4630,N_4968);
nor U5297 (N_5297,N_4044,N_4916);
xnor U5298 (N_5298,N_4747,N_4397);
xor U5299 (N_5299,N_4643,N_4434);
and U5300 (N_5300,N_4625,N_4689);
or U5301 (N_5301,N_4876,N_4349);
and U5302 (N_5302,N_4582,N_4041);
xnor U5303 (N_5303,N_4829,N_4604);
xnor U5304 (N_5304,N_4685,N_4881);
nand U5305 (N_5305,N_4892,N_4848);
nand U5306 (N_5306,N_4901,N_4809);
nor U5307 (N_5307,N_4365,N_4123);
or U5308 (N_5308,N_4306,N_4154);
and U5309 (N_5309,N_4430,N_4220);
nand U5310 (N_5310,N_4955,N_4895);
and U5311 (N_5311,N_4492,N_4013);
nand U5312 (N_5312,N_4115,N_4368);
or U5313 (N_5313,N_4444,N_4920);
xor U5314 (N_5314,N_4744,N_4887);
xnor U5315 (N_5315,N_4082,N_4345);
nand U5316 (N_5316,N_4194,N_4914);
and U5317 (N_5317,N_4534,N_4246);
nand U5318 (N_5318,N_4864,N_4647);
xnor U5319 (N_5319,N_4780,N_4404);
or U5320 (N_5320,N_4403,N_4862);
nand U5321 (N_5321,N_4874,N_4284);
xnor U5322 (N_5322,N_4585,N_4696);
xnor U5323 (N_5323,N_4009,N_4464);
xor U5324 (N_5324,N_4398,N_4679);
and U5325 (N_5325,N_4373,N_4743);
nor U5326 (N_5326,N_4731,N_4935);
nand U5327 (N_5327,N_4006,N_4910);
or U5328 (N_5328,N_4281,N_4618);
nor U5329 (N_5329,N_4371,N_4899);
and U5330 (N_5330,N_4423,N_4217);
or U5331 (N_5331,N_4692,N_4064);
xor U5332 (N_5332,N_4253,N_4479);
nor U5333 (N_5333,N_4709,N_4407);
nor U5334 (N_5334,N_4606,N_4634);
or U5335 (N_5335,N_4562,N_4329);
xnor U5336 (N_5336,N_4156,N_4966);
xnor U5337 (N_5337,N_4551,N_4611);
or U5338 (N_5338,N_4400,N_4921);
nor U5339 (N_5339,N_4205,N_4475);
nand U5340 (N_5340,N_4882,N_4504);
xnor U5341 (N_5341,N_4449,N_4500);
xor U5342 (N_5342,N_4885,N_4715);
nand U5343 (N_5343,N_4017,N_4435);
nand U5344 (N_5344,N_4616,N_4644);
and U5345 (N_5345,N_4824,N_4828);
nor U5346 (N_5346,N_4155,N_4631);
xnor U5347 (N_5347,N_4951,N_4033);
and U5348 (N_5348,N_4014,N_4418);
and U5349 (N_5349,N_4163,N_4094);
and U5350 (N_5350,N_4494,N_4290);
and U5351 (N_5351,N_4346,N_4328);
xor U5352 (N_5352,N_4146,N_4469);
nand U5353 (N_5353,N_4243,N_4066);
xor U5354 (N_5354,N_4965,N_4207);
xor U5355 (N_5355,N_4572,N_4932);
nand U5356 (N_5356,N_4591,N_4939);
or U5357 (N_5357,N_4196,N_4185);
or U5358 (N_5358,N_4216,N_4303);
xor U5359 (N_5359,N_4710,N_4950);
and U5360 (N_5360,N_4732,N_4717);
or U5361 (N_5361,N_4355,N_4412);
xor U5362 (N_5362,N_4557,N_4594);
nand U5363 (N_5363,N_4635,N_4442);
xnor U5364 (N_5364,N_4003,N_4580);
xnor U5365 (N_5365,N_4419,N_4320);
nor U5366 (N_5366,N_4394,N_4204);
nor U5367 (N_5367,N_4148,N_4010);
nor U5368 (N_5368,N_4627,N_4273);
or U5369 (N_5369,N_4898,N_4578);
xor U5370 (N_5370,N_4560,N_4084);
and U5371 (N_5371,N_4949,N_4344);
nor U5372 (N_5372,N_4510,N_4316);
or U5373 (N_5373,N_4379,N_4778);
xnor U5374 (N_5374,N_4767,N_4632);
xor U5375 (N_5375,N_4537,N_4342);
nand U5376 (N_5376,N_4751,N_4278);
nor U5377 (N_5377,N_4520,N_4592);
nand U5378 (N_5378,N_4252,N_4249);
nand U5379 (N_5379,N_4863,N_4896);
nand U5380 (N_5380,N_4571,N_4740);
or U5381 (N_5381,N_4376,N_4758);
and U5382 (N_5382,N_4739,N_4331);
and U5383 (N_5383,N_4708,N_4840);
or U5384 (N_5384,N_4099,N_4576);
xor U5385 (N_5385,N_4776,N_4992);
nor U5386 (N_5386,N_4794,N_4413);
xor U5387 (N_5387,N_4490,N_4496);
or U5388 (N_5388,N_4102,N_4713);
nand U5389 (N_5389,N_4525,N_4179);
or U5390 (N_5390,N_4286,N_4210);
and U5391 (N_5391,N_4028,N_4001);
xnor U5392 (N_5392,N_4937,N_4107);
xor U5393 (N_5393,N_4762,N_4265);
xor U5394 (N_5394,N_4251,N_4111);
nand U5395 (N_5395,N_4745,N_4771);
xor U5396 (N_5396,N_4553,N_4807);
nand U5397 (N_5397,N_4122,N_4543);
xnor U5398 (N_5398,N_4880,N_4834);
or U5399 (N_5399,N_4952,N_4425);
nand U5400 (N_5400,N_4522,N_4415);
xnor U5401 (N_5401,N_4161,N_4978);
nand U5402 (N_5402,N_4011,N_4127);
nand U5403 (N_5403,N_4230,N_4237);
or U5404 (N_5404,N_4719,N_4386);
or U5405 (N_5405,N_4906,N_4608);
nand U5406 (N_5406,N_4970,N_4463);
and U5407 (N_5407,N_4097,N_4730);
and U5408 (N_5408,N_4428,N_4327);
nand U5409 (N_5409,N_4022,N_4548);
or U5410 (N_5410,N_4825,N_4990);
xor U5411 (N_5411,N_4359,N_4948);
nand U5412 (N_5412,N_4855,N_4300);
nor U5413 (N_5413,N_4657,N_4593);
or U5414 (N_5414,N_4818,N_4686);
xnor U5415 (N_5415,N_4211,N_4233);
and U5416 (N_5416,N_4267,N_4960);
or U5417 (N_5417,N_4078,N_4299);
nand U5418 (N_5418,N_4214,N_4770);
and U5419 (N_5419,N_4042,N_4167);
nor U5420 (N_5420,N_4781,N_4020);
and U5421 (N_5421,N_4466,N_4590);
nor U5422 (N_5422,N_4460,N_4760);
xor U5423 (N_5423,N_4240,N_4963);
xor U5424 (N_5424,N_4468,N_4969);
nor U5425 (N_5425,N_4441,N_4259);
nor U5426 (N_5426,N_4219,N_4206);
nand U5427 (N_5427,N_4915,N_4269);
xnor U5428 (N_5428,N_4746,N_4650);
nor U5429 (N_5429,N_4523,N_4040);
xnor U5430 (N_5430,N_4471,N_4315);
nand U5431 (N_5431,N_4624,N_4656);
xor U5432 (N_5432,N_4664,N_4261);
nand U5433 (N_5433,N_4964,N_4473);
nor U5434 (N_5434,N_4004,N_4620);
and U5435 (N_5435,N_4947,N_4197);
or U5436 (N_5436,N_4574,N_4021);
nor U5437 (N_5437,N_4235,N_4061);
nand U5438 (N_5438,N_4455,N_4170);
nor U5439 (N_5439,N_4275,N_4254);
xnor U5440 (N_5440,N_4766,N_4509);
nor U5441 (N_5441,N_4695,N_4245);
xor U5442 (N_5442,N_4805,N_4353);
or U5443 (N_5443,N_4930,N_4406);
nor U5444 (N_5444,N_4374,N_4756);
and U5445 (N_5445,N_4796,N_4005);
nor U5446 (N_5446,N_4383,N_4431);
nor U5447 (N_5447,N_4225,N_4452);
or U5448 (N_5448,N_4016,N_4087);
nor U5449 (N_5449,N_4209,N_4849);
nor U5450 (N_5450,N_4533,N_4755);
and U5451 (N_5451,N_4367,N_4351);
nor U5452 (N_5452,N_4250,N_4382);
nor U5453 (N_5453,N_4132,N_4980);
or U5454 (N_5454,N_4975,N_4676);
nor U5455 (N_5455,N_4080,N_4489);
and U5456 (N_5456,N_4302,N_4911);
and U5457 (N_5457,N_4588,N_4640);
nor U5458 (N_5458,N_4459,N_4288);
xnor U5459 (N_5459,N_4682,N_4101);
xor U5460 (N_5460,N_4069,N_4789);
xnor U5461 (N_5461,N_4023,N_4128);
and U5462 (N_5462,N_4140,N_4521);
and U5463 (N_5463,N_4511,N_4577);
nor U5464 (N_5464,N_4362,N_4360);
and U5465 (N_5465,N_4247,N_4742);
or U5466 (N_5466,N_4962,N_4977);
or U5467 (N_5467,N_4798,N_4532);
or U5468 (N_5468,N_4350,N_4279);
nand U5469 (N_5469,N_4238,N_4817);
and U5470 (N_5470,N_4505,N_4889);
xor U5471 (N_5471,N_4298,N_4905);
nand U5472 (N_5472,N_4285,N_4224);
nand U5473 (N_5473,N_4808,N_4674);
xor U5474 (N_5474,N_4181,N_4239);
and U5475 (N_5475,N_4326,N_4184);
nor U5476 (N_5476,N_4827,N_4176);
nand U5477 (N_5477,N_4341,N_4491);
or U5478 (N_5478,N_4662,N_4687);
and U5479 (N_5479,N_4387,N_4787);
nor U5480 (N_5480,N_4869,N_4702);
nand U5481 (N_5481,N_4547,N_4788);
xor U5482 (N_5482,N_4410,N_4724);
nor U5483 (N_5483,N_4642,N_4773);
or U5484 (N_5484,N_4677,N_4108);
or U5485 (N_5485,N_4065,N_4077);
and U5486 (N_5486,N_4191,N_4304);
nor U5487 (N_5487,N_4159,N_4545);
and U5488 (N_5488,N_4806,N_4098);
nor U5489 (N_5489,N_4256,N_4688);
xnor U5490 (N_5490,N_4938,N_4622);
xnor U5491 (N_5491,N_4559,N_4189);
nand U5492 (N_5492,N_4803,N_4663);
nand U5493 (N_5493,N_4260,N_4296);
nor U5494 (N_5494,N_4208,N_4114);
xnor U5495 (N_5495,N_4684,N_4391);
and U5496 (N_5496,N_4142,N_4944);
or U5497 (N_5497,N_4271,N_4438);
or U5498 (N_5498,N_4032,N_4996);
xnor U5499 (N_5499,N_4283,N_4103);
and U5500 (N_5500,N_4567,N_4503);
or U5501 (N_5501,N_4321,N_4253);
xor U5502 (N_5502,N_4483,N_4119);
nor U5503 (N_5503,N_4150,N_4019);
nand U5504 (N_5504,N_4967,N_4353);
nor U5505 (N_5505,N_4984,N_4372);
nand U5506 (N_5506,N_4838,N_4269);
nor U5507 (N_5507,N_4208,N_4782);
and U5508 (N_5508,N_4646,N_4373);
nand U5509 (N_5509,N_4913,N_4691);
and U5510 (N_5510,N_4488,N_4164);
nor U5511 (N_5511,N_4063,N_4605);
xor U5512 (N_5512,N_4621,N_4831);
xnor U5513 (N_5513,N_4544,N_4407);
nand U5514 (N_5514,N_4198,N_4130);
nand U5515 (N_5515,N_4425,N_4157);
xor U5516 (N_5516,N_4690,N_4114);
nor U5517 (N_5517,N_4718,N_4217);
or U5518 (N_5518,N_4921,N_4860);
nand U5519 (N_5519,N_4638,N_4307);
nor U5520 (N_5520,N_4850,N_4900);
nand U5521 (N_5521,N_4964,N_4199);
nand U5522 (N_5522,N_4202,N_4544);
or U5523 (N_5523,N_4308,N_4074);
nor U5524 (N_5524,N_4826,N_4245);
or U5525 (N_5525,N_4377,N_4374);
and U5526 (N_5526,N_4771,N_4617);
nand U5527 (N_5527,N_4697,N_4828);
and U5528 (N_5528,N_4321,N_4894);
or U5529 (N_5529,N_4566,N_4502);
and U5530 (N_5530,N_4769,N_4561);
nand U5531 (N_5531,N_4168,N_4732);
nand U5532 (N_5532,N_4620,N_4179);
nand U5533 (N_5533,N_4104,N_4020);
and U5534 (N_5534,N_4871,N_4603);
and U5535 (N_5535,N_4559,N_4694);
or U5536 (N_5536,N_4659,N_4164);
nor U5537 (N_5537,N_4170,N_4701);
or U5538 (N_5538,N_4771,N_4795);
and U5539 (N_5539,N_4057,N_4975);
and U5540 (N_5540,N_4965,N_4455);
xor U5541 (N_5541,N_4365,N_4720);
xnor U5542 (N_5542,N_4125,N_4720);
xor U5543 (N_5543,N_4063,N_4082);
nor U5544 (N_5544,N_4109,N_4010);
and U5545 (N_5545,N_4245,N_4662);
and U5546 (N_5546,N_4473,N_4005);
nor U5547 (N_5547,N_4416,N_4421);
nor U5548 (N_5548,N_4799,N_4508);
xnor U5549 (N_5549,N_4847,N_4127);
nand U5550 (N_5550,N_4567,N_4806);
xnor U5551 (N_5551,N_4296,N_4427);
nor U5552 (N_5552,N_4723,N_4606);
xor U5553 (N_5553,N_4803,N_4668);
nor U5554 (N_5554,N_4292,N_4828);
nor U5555 (N_5555,N_4391,N_4733);
nor U5556 (N_5556,N_4194,N_4519);
nand U5557 (N_5557,N_4057,N_4986);
nor U5558 (N_5558,N_4791,N_4471);
xor U5559 (N_5559,N_4108,N_4268);
and U5560 (N_5560,N_4527,N_4358);
or U5561 (N_5561,N_4991,N_4556);
and U5562 (N_5562,N_4391,N_4424);
xor U5563 (N_5563,N_4764,N_4074);
or U5564 (N_5564,N_4772,N_4265);
nand U5565 (N_5565,N_4409,N_4293);
or U5566 (N_5566,N_4495,N_4876);
xnor U5567 (N_5567,N_4396,N_4588);
nor U5568 (N_5568,N_4685,N_4189);
and U5569 (N_5569,N_4366,N_4039);
and U5570 (N_5570,N_4309,N_4437);
nor U5571 (N_5571,N_4937,N_4972);
or U5572 (N_5572,N_4181,N_4642);
nor U5573 (N_5573,N_4812,N_4158);
nand U5574 (N_5574,N_4001,N_4873);
nor U5575 (N_5575,N_4627,N_4798);
and U5576 (N_5576,N_4615,N_4824);
nand U5577 (N_5577,N_4708,N_4276);
and U5578 (N_5578,N_4083,N_4467);
nand U5579 (N_5579,N_4621,N_4524);
and U5580 (N_5580,N_4191,N_4508);
and U5581 (N_5581,N_4714,N_4861);
nand U5582 (N_5582,N_4201,N_4195);
nor U5583 (N_5583,N_4191,N_4529);
nand U5584 (N_5584,N_4230,N_4529);
nand U5585 (N_5585,N_4311,N_4227);
or U5586 (N_5586,N_4494,N_4287);
xnor U5587 (N_5587,N_4182,N_4651);
nand U5588 (N_5588,N_4509,N_4831);
xor U5589 (N_5589,N_4544,N_4035);
xnor U5590 (N_5590,N_4268,N_4713);
xor U5591 (N_5591,N_4003,N_4731);
xnor U5592 (N_5592,N_4945,N_4924);
or U5593 (N_5593,N_4759,N_4740);
xnor U5594 (N_5594,N_4556,N_4581);
nor U5595 (N_5595,N_4969,N_4305);
and U5596 (N_5596,N_4467,N_4407);
or U5597 (N_5597,N_4398,N_4014);
nor U5598 (N_5598,N_4763,N_4497);
and U5599 (N_5599,N_4963,N_4057);
or U5600 (N_5600,N_4056,N_4572);
or U5601 (N_5601,N_4242,N_4223);
xnor U5602 (N_5602,N_4312,N_4895);
or U5603 (N_5603,N_4295,N_4144);
and U5604 (N_5604,N_4586,N_4226);
nor U5605 (N_5605,N_4178,N_4227);
nor U5606 (N_5606,N_4184,N_4495);
or U5607 (N_5607,N_4991,N_4910);
xor U5608 (N_5608,N_4179,N_4836);
and U5609 (N_5609,N_4741,N_4307);
or U5610 (N_5610,N_4179,N_4665);
nor U5611 (N_5611,N_4858,N_4683);
nor U5612 (N_5612,N_4803,N_4169);
nor U5613 (N_5613,N_4927,N_4877);
xnor U5614 (N_5614,N_4404,N_4758);
and U5615 (N_5615,N_4237,N_4326);
xor U5616 (N_5616,N_4691,N_4254);
nor U5617 (N_5617,N_4881,N_4997);
nand U5618 (N_5618,N_4302,N_4966);
nand U5619 (N_5619,N_4067,N_4398);
nor U5620 (N_5620,N_4265,N_4273);
nand U5621 (N_5621,N_4379,N_4217);
and U5622 (N_5622,N_4420,N_4398);
or U5623 (N_5623,N_4125,N_4987);
xor U5624 (N_5624,N_4697,N_4895);
nor U5625 (N_5625,N_4525,N_4069);
and U5626 (N_5626,N_4440,N_4095);
nor U5627 (N_5627,N_4186,N_4611);
or U5628 (N_5628,N_4359,N_4086);
or U5629 (N_5629,N_4054,N_4248);
or U5630 (N_5630,N_4845,N_4002);
nand U5631 (N_5631,N_4648,N_4823);
and U5632 (N_5632,N_4085,N_4450);
xnor U5633 (N_5633,N_4363,N_4226);
nand U5634 (N_5634,N_4551,N_4759);
nand U5635 (N_5635,N_4301,N_4230);
xnor U5636 (N_5636,N_4615,N_4850);
xor U5637 (N_5637,N_4066,N_4395);
nor U5638 (N_5638,N_4010,N_4243);
nand U5639 (N_5639,N_4307,N_4850);
xor U5640 (N_5640,N_4640,N_4722);
nor U5641 (N_5641,N_4536,N_4990);
nand U5642 (N_5642,N_4215,N_4957);
xnor U5643 (N_5643,N_4951,N_4338);
or U5644 (N_5644,N_4894,N_4644);
nand U5645 (N_5645,N_4122,N_4374);
or U5646 (N_5646,N_4225,N_4537);
xnor U5647 (N_5647,N_4244,N_4898);
nor U5648 (N_5648,N_4486,N_4477);
or U5649 (N_5649,N_4020,N_4844);
nor U5650 (N_5650,N_4273,N_4908);
or U5651 (N_5651,N_4290,N_4377);
xnor U5652 (N_5652,N_4106,N_4714);
nand U5653 (N_5653,N_4846,N_4770);
nand U5654 (N_5654,N_4406,N_4221);
or U5655 (N_5655,N_4797,N_4857);
and U5656 (N_5656,N_4041,N_4652);
or U5657 (N_5657,N_4881,N_4193);
and U5658 (N_5658,N_4968,N_4815);
xnor U5659 (N_5659,N_4638,N_4964);
and U5660 (N_5660,N_4969,N_4282);
or U5661 (N_5661,N_4033,N_4433);
xor U5662 (N_5662,N_4722,N_4609);
nor U5663 (N_5663,N_4579,N_4804);
xnor U5664 (N_5664,N_4538,N_4134);
nand U5665 (N_5665,N_4261,N_4115);
or U5666 (N_5666,N_4870,N_4429);
nand U5667 (N_5667,N_4669,N_4259);
and U5668 (N_5668,N_4193,N_4649);
xnor U5669 (N_5669,N_4403,N_4934);
nor U5670 (N_5670,N_4738,N_4967);
nand U5671 (N_5671,N_4894,N_4850);
or U5672 (N_5672,N_4591,N_4434);
nand U5673 (N_5673,N_4079,N_4680);
and U5674 (N_5674,N_4661,N_4206);
and U5675 (N_5675,N_4506,N_4694);
and U5676 (N_5676,N_4343,N_4261);
or U5677 (N_5677,N_4546,N_4037);
and U5678 (N_5678,N_4110,N_4894);
and U5679 (N_5679,N_4602,N_4479);
nand U5680 (N_5680,N_4710,N_4001);
nand U5681 (N_5681,N_4669,N_4176);
xor U5682 (N_5682,N_4046,N_4607);
and U5683 (N_5683,N_4936,N_4886);
or U5684 (N_5684,N_4635,N_4064);
nor U5685 (N_5685,N_4909,N_4413);
or U5686 (N_5686,N_4724,N_4788);
nor U5687 (N_5687,N_4038,N_4252);
nor U5688 (N_5688,N_4260,N_4579);
and U5689 (N_5689,N_4950,N_4092);
and U5690 (N_5690,N_4817,N_4952);
nor U5691 (N_5691,N_4381,N_4517);
xor U5692 (N_5692,N_4278,N_4789);
xnor U5693 (N_5693,N_4472,N_4804);
nand U5694 (N_5694,N_4866,N_4609);
nor U5695 (N_5695,N_4355,N_4220);
nand U5696 (N_5696,N_4216,N_4535);
xnor U5697 (N_5697,N_4410,N_4661);
or U5698 (N_5698,N_4149,N_4352);
or U5699 (N_5699,N_4386,N_4599);
nor U5700 (N_5700,N_4305,N_4538);
or U5701 (N_5701,N_4842,N_4245);
nor U5702 (N_5702,N_4767,N_4184);
or U5703 (N_5703,N_4584,N_4492);
nand U5704 (N_5704,N_4272,N_4534);
or U5705 (N_5705,N_4691,N_4169);
xnor U5706 (N_5706,N_4199,N_4113);
xor U5707 (N_5707,N_4712,N_4373);
xor U5708 (N_5708,N_4508,N_4004);
nor U5709 (N_5709,N_4956,N_4228);
nand U5710 (N_5710,N_4874,N_4495);
nor U5711 (N_5711,N_4125,N_4305);
and U5712 (N_5712,N_4073,N_4631);
and U5713 (N_5713,N_4008,N_4891);
xor U5714 (N_5714,N_4142,N_4201);
xor U5715 (N_5715,N_4784,N_4512);
nand U5716 (N_5716,N_4316,N_4573);
and U5717 (N_5717,N_4469,N_4169);
nor U5718 (N_5718,N_4946,N_4739);
nand U5719 (N_5719,N_4433,N_4766);
nor U5720 (N_5720,N_4914,N_4430);
and U5721 (N_5721,N_4334,N_4111);
nand U5722 (N_5722,N_4761,N_4377);
and U5723 (N_5723,N_4356,N_4618);
or U5724 (N_5724,N_4904,N_4060);
nor U5725 (N_5725,N_4355,N_4940);
nor U5726 (N_5726,N_4746,N_4598);
and U5727 (N_5727,N_4814,N_4350);
or U5728 (N_5728,N_4453,N_4998);
and U5729 (N_5729,N_4784,N_4294);
nor U5730 (N_5730,N_4303,N_4298);
or U5731 (N_5731,N_4903,N_4654);
nand U5732 (N_5732,N_4430,N_4146);
nor U5733 (N_5733,N_4838,N_4172);
xor U5734 (N_5734,N_4763,N_4991);
nand U5735 (N_5735,N_4519,N_4105);
nor U5736 (N_5736,N_4711,N_4840);
xor U5737 (N_5737,N_4725,N_4744);
nor U5738 (N_5738,N_4110,N_4990);
and U5739 (N_5739,N_4825,N_4742);
and U5740 (N_5740,N_4466,N_4074);
and U5741 (N_5741,N_4753,N_4689);
nand U5742 (N_5742,N_4981,N_4189);
xnor U5743 (N_5743,N_4849,N_4546);
xor U5744 (N_5744,N_4609,N_4532);
nand U5745 (N_5745,N_4527,N_4741);
nand U5746 (N_5746,N_4263,N_4729);
and U5747 (N_5747,N_4261,N_4903);
nand U5748 (N_5748,N_4595,N_4715);
or U5749 (N_5749,N_4788,N_4941);
and U5750 (N_5750,N_4288,N_4990);
nand U5751 (N_5751,N_4880,N_4492);
xor U5752 (N_5752,N_4923,N_4712);
nor U5753 (N_5753,N_4583,N_4943);
nand U5754 (N_5754,N_4031,N_4528);
xor U5755 (N_5755,N_4966,N_4215);
nand U5756 (N_5756,N_4642,N_4884);
xnor U5757 (N_5757,N_4805,N_4234);
xor U5758 (N_5758,N_4806,N_4226);
and U5759 (N_5759,N_4868,N_4024);
nand U5760 (N_5760,N_4291,N_4656);
and U5761 (N_5761,N_4737,N_4050);
nand U5762 (N_5762,N_4265,N_4340);
and U5763 (N_5763,N_4357,N_4819);
or U5764 (N_5764,N_4600,N_4453);
or U5765 (N_5765,N_4739,N_4146);
xnor U5766 (N_5766,N_4098,N_4672);
and U5767 (N_5767,N_4462,N_4431);
xor U5768 (N_5768,N_4959,N_4829);
xor U5769 (N_5769,N_4524,N_4398);
or U5770 (N_5770,N_4995,N_4520);
or U5771 (N_5771,N_4888,N_4193);
and U5772 (N_5772,N_4634,N_4888);
nand U5773 (N_5773,N_4512,N_4070);
nor U5774 (N_5774,N_4767,N_4032);
and U5775 (N_5775,N_4909,N_4484);
nand U5776 (N_5776,N_4125,N_4594);
xnor U5777 (N_5777,N_4004,N_4298);
or U5778 (N_5778,N_4797,N_4754);
and U5779 (N_5779,N_4439,N_4307);
or U5780 (N_5780,N_4875,N_4164);
and U5781 (N_5781,N_4093,N_4277);
nor U5782 (N_5782,N_4085,N_4694);
nand U5783 (N_5783,N_4321,N_4108);
nor U5784 (N_5784,N_4474,N_4512);
and U5785 (N_5785,N_4401,N_4232);
xnor U5786 (N_5786,N_4120,N_4551);
and U5787 (N_5787,N_4909,N_4553);
and U5788 (N_5788,N_4068,N_4565);
xor U5789 (N_5789,N_4797,N_4107);
and U5790 (N_5790,N_4295,N_4487);
nor U5791 (N_5791,N_4337,N_4400);
or U5792 (N_5792,N_4034,N_4930);
nor U5793 (N_5793,N_4455,N_4266);
or U5794 (N_5794,N_4465,N_4034);
nor U5795 (N_5795,N_4847,N_4785);
or U5796 (N_5796,N_4602,N_4088);
or U5797 (N_5797,N_4244,N_4576);
nor U5798 (N_5798,N_4577,N_4605);
nor U5799 (N_5799,N_4924,N_4076);
nand U5800 (N_5800,N_4523,N_4097);
nor U5801 (N_5801,N_4523,N_4943);
xor U5802 (N_5802,N_4550,N_4275);
nor U5803 (N_5803,N_4014,N_4839);
and U5804 (N_5804,N_4315,N_4526);
nand U5805 (N_5805,N_4865,N_4250);
or U5806 (N_5806,N_4004,N_4475);
and U5807 (N_5807,N_4890,N_4406);
and U5808 (N_5808,N_4022,N_4240);
or U5809 (N_5809,N_4756,N_4873);
nand U5810 (N_5810,N_4098,N_4286);
and U5811 (N_5811,N_4143,N_4792);
and U5812 (N_5812,N_4609,N_4668);
nor U5813 (N_5813,N_4098,N_4103);
nor U5814 (N_5814,N_4848,N_4697);
nor U5815 (N_5815,N_4226,N_4479);
nand U5816 (N_5816,N_4968,N_4371);
xnor U5817 (N_5817,N_4331,N_4622);
nor U5818 (N_5818,N_4216,N_4006);
nand U5819 (N_5819,N_4050,N_4053);
or U5820 (N_5820,N_4706,N_4540);
and U5821 (N_5821,N_4668,N_4986);
or U5822 (N_5822,N_4554,N_4531);
or U5823 (N_5823,N_4475,N_4996);
and U5824 (N_5824,N_4612,N_4759);
or U5825 (N_5825,N_4612,N_4650);
xnor U5826 (N_5826,N_4229,N_4895);
or U5827 (N_5827,N_4996,N_4245);
nor U5828 (N_5828,N_4201,N_4217);
or U5829 (N_5829,N_4297,N_4266);
xnor U5830 (N_5830,N_4674,N_4835);
xor U5831 (N_5831,N_4469,N_4223);
nand U5832 (N_5832,N_4464,N_4215);
nand U5833 (N_5833,N_4028,N_4893);
and U5834 (N_5834,N_4328,N_4828);
nand U5835 (N_5835,N_4849,N_4353);
nor U5836 (N_5836,N_4272,N_4451);
nand U5837 (N_5837,N_4134,N_4428);
nand U5838 (N_5838,N_4026,N_4448);
and U5839 (N_5839,N_4430,N_4078);
or U5840 (N_5840,N_4276,N_4071);
and U5841 (N_5841,N_4155,N_4757);
nor U5842 (N_5842,N_4513,N_4906);
and U5843 (N_5843,N_4744,N_4842);
or U5844 (N_5844,N_4909,N_4243);
and U5845 (N_5845,N_4629,N_4952);
nor U5846 (N_5846,N_4746,N_4658);
nand U5847 (N_5847,N_4493,N_4891);
or U5848 (N_5848,N_4455,N_4569);
xnor U5849 (N_5849,N_4570,N_4017);
or U5850 (N_5850,N_4425,N_4998);
and U5851 (N_5851,N_4136,N_4823);
nand U5852 (N_5852,N_4375,N_4918);
nor U5853 (N_5853,N_4359,N_4223);
xnor U5854 (N_5854,N_4011,N_4950);
xnor U5855 (N_5855,N_4547,N_4838);
nor U5856 (N_5856,N_4454,N_4790);
xor U5857 (N_5857,N_4267,N_4330);
nand U5858 (N_5858,N_4638,N_4596);
nor U5859 (N_5859,N_4219,N_4410);
and U5860 (N_5860,N_4900,N_4413);
and U5861 (N_5861,N_4518,N_4690);
or U5862 (N_5862,N_4748,N_4185);
nor U5863 (N_5863,N_4781,N_4829);
or U5864 (N_5864,N_4227,N_4395);
or U5865 (N_5865,N_4534,N_4329);
and U5866 (N_5866,N_4296,N_4339);
xor U5867 (N_5867,N_4788,N_4930);
or U5868 (N_5868,N_4131,N_4596);
nand U5869 (N_5869,N_4939,N_4607);
nor U5870 (N_5870,N_4871,N_4060);
and U5871 (N_5871,N_4803,N_4624);
and U5872 (N_5872,N_4648,N_4842);
or U5873 (N_5873,N_4636,N_4547);
or U5874 (N_5874,N_4070,N_4212);
and U5875 (N_5875,N_4458,N_4983);
xor U5876 (N_5876,N_4017,N_4382);
nor U5877 (N_5877,N_4232,N_4302);
xnor U5878 (N_5878,N_4954,N_4039);
nor U5879 (N_5879,N_4771,N_4003);
xor U5880 (N_5880,N_4260,N_4307);
nor U5881 (N_5881,N_4553,N_4515);
nand U5882 (N_5882,N_4679,N_4648);
nand U5883 (N_5883,N_4515,N_4747);
nor U5884 (N_5884,N_4173,N_4282);
nand U5885 (N_5885,N_4034,N_4460);
nor U5886 (N_5886,N_4109,N_4642);
nand U5887 (N_5887,N_4811,N_4032);
or U5888 (N_5888,N_4445,N_4593);
or U5889 (N_5889,N_4669,N_4662);
xor U5890 (N_5890,N_4955,N_4406);
nor U5891 (N_5891,N_4130,N_4357);
nand U5892 (N_5892,N_4870,N_4895);
xnor U5893 (N_5893,N_4192,N_4364);
nand U5894 (N_5894,N_4159,N_4052);
nor U5895 (N_5895,N_4489,N_4933);
or U5896 (N_5896,N_4061,N_4391);
nor U5897 (N_5897,N_4584,N_4359);
nand U5898 (N_5898,N_4419,N_4196);
nand U5899 (N_5899,N_4461,N_4258);
and U5900 (N_5900,N_4326,N_4080);
and U5901 (N_5901,N_4421,N_4924);
nor U5902 (N_5902,N_4574,N_4298);
xnor U5903 (N_5903,N_4604,N_4944);
nand U5904 (N_5904,N_4986,N_4408);
nand U5905 (N_5905,N_4022,N_4765);
nand U5906 (N_5906,N_4646,N_4872);
and U5907 (N_5907,N_4628,N_4781);
and U5908 (N_5908,N_4344,N_4755);
xor U5909 (N_5909,N_4919,N_4639);
xor U5910 (N_5910,N_4777,N_4946);
nand U5911 (N_5911,N_4545,N_4475);
xor U5912 (N_5912,N_4087,N_4891);
nor U5913 (N_5913,N_4472,N_4768);
xnor U5914 (N_5914,N_4328,N_4570);
or U5915 (N_5915,N_4282,N_4368);
nor U5916 (N_5916,N_4716,N_4781);
nor U5917 (N_5917,N_4261,N_4262);
xnor U5918 (N_5918,N_4964,N_4197);
nand U5919 (N_5919,N_4754,N_4258);
or U5920 (N_5920,N_4393,N_4858);
xnor U5921 (N_5921,N_4159,N_4913);
and U5922 (N_5922,N_4143,N_4800);
or U5923 (N_5923,N_4044,N_4088);
or U5924 (N_5924,N_4319,N_4741);
xor U5925 (N_5925,N_4093,N_4242);
nor U5926 (N_5926,N_4633,N_4493);
nor U5927 (N_5927,N_4323,N_4171);
nor U5928 (N_5928,N_4107,N_4566);
and U5929 (N_5929,N_4004,N_4968);
nor U5930 (N_5930,N_4435,N_4308);
or U5931 (N_5931,N_4231,N_4037);
nand U5932 (N_5932,N_4710,N_4626);
nor U5933 (N_5933,N_4124,N_4256);
and U5934 (N_5934,N_4267,N_4947);
or U5935 (N_5935,N_4167,N_4745);
xor U5936 (N_5936,N_4978,N_4392);
or U5937 (N_5937,N_4348,N_4982);
and U5938 (N_5938,N_4444,N_4961);
nor U5939 (N_5939,N_4087,N_4101);
xnor U5940 (N_5940,N_4288,N_4007);
and U5941 (N_5941,N_4179,N_4870);
or U5942 (N_5942,N_4950,N_4738);
xor U5943 (N_5943,N_4416,N_4027);
or U5944 (N_5944,N_4551,N_4179);
nor U5945 (N_5945,N_4492,N_4668);
nand U5946 (N_5946,N_4329,N_4472);
and U5947 (N_5947,N_4501,N_4008);
nor U5948 (N_5948,N_4386,N_4752);
nor U5949 (N_5949,N_4784,N_4276);
nand U5950 (N_5950,N_4029,N_4593);
or U5951 (N_5951,N_4887,N_4455);
or U5952 (N_5952,N_4955,N_4202);
nor U5953 (N_5953,N_4160,N_4639);
xnor U5954 (N_5954,N_4784,N_4499);
and U5955 (N_5955,N_4993,N_4744);
or U5956 (N_5956,N_4972,N_4689);
nand U5957 (N_5957,N_4428,N_4776);
xnor U5958 (N_5958,N_4223,N_4832);
xor U5959 (N_5959,N_4424,N_4852);
xnor U5960 (N_5960,N_4165,N_4767);
or U5961 (N_5961,N_4340,N_4379);
nor U5962 (N_5962,N_4371,N_4362);
xnor U5963 (N_5963,N_4177,N_4509);
xnor U5964 (N_5964,N_4453,N_4335);
or U5965 (N_5965,N_4947,N_4788);
and U5966 (N_5966,N_4776,N_4634);
and U5967 (N_5967,N_4865,N_4768);
or U5968 (N_5968,N_4924,N_4950);
or U5969 (N_5969,N_4786,N_4092);
and U5970 (N_5970,N_4016,N_4555);
nand U5971 (N_5971,N_4094,N_4445);
nor U5972 (N_5972,N_4302,N_4827);
nand U5973 (N_5973,N_4001,N_4410);
nand U5974 (N_5974,N_4108,N_4838);
or U5975 (N_5975,N_4241,N_4590);
xnor U5976 (N_5976,N_4152,N_4856);
and U5977 (N_5977,N_4709,N_4942);
nor U5978 (N_5978,N_4777,N_4873);
nand U5979 (N_5979,N_4047,N_4170);
xor U5980 (N_5980,N_4196,N_4364);
nor U5981 (N_5981,N_4259,N_4418);
nand U5982 (N_5982,N_4308,N_4120);
nor U5983 (N_5983,N_4717,N_4695);
nand U5984 (N_5984,N_4154,N_4066);
nand U5985 (N_5985,N_4304,N_4883);
and U5986 (N_5986,N_4427,N_4990);
xor U5987 (N_5987,N_4417,N_4378);
nand U5988 (N_5988,N_4758,N_4721);
nor U5989 (N_5989,N_4923,N_4683);
nand U5990 (N_5990,N_4597,N_4191);
nor U5991 (N_5991,N_4652,N_4658);
nand U5992 (N_5992,N_4559,N_4851);
and U5993 (N_5993,N_4166,N_4685);
and U5994 (N_5994,N_4949,N_4071);
xnor U5995 (N_5995,N_4298,N_4739);
and U5996 (N_5996,N_4505,N_4391);
and U5997 (N_5997,N_4760,N_4819);
xnor U5998 (N_5998,N_4772,N_4753);
or U5999 (N_5999,N_4771,N_4100);
xor U6000 (N_6000,N_5458,N_5279);
and U6001 (N_6001,N_5796,N_5445);
and U6002 (N_6002,N_5207,N_5942);
nand U6003 (N_6003,N_5679,N_5506);
or U6004 (N_6004,N_5593,N_5031);
nor U6005 (N_6005,N_5700,N_5763);
xor U6006 (N_6006,N_5660,N_5632);
xor U6007 (N_6007,N_5200,N_5585);
or U6008 (N_6008,N_5893,N_5193);
and U6009 (N_6009,N_5344,N_5244);
xor U6010 (N_6010,N_5802,N_5111);
and U6011 (N_6011,N_5347,N_5994);
and U6012 (N_6012,N_5661,N_5842);
nand U6013 (N_6013,N_5823,N_5190);
xnor U6014 (N_6014,N_5872,N_5595);
or U6015 (N_6015,N_5248,N_5432);
xor U6016 (N_6016,N_5156,N_5274);
or U6017 (N_6017,N_5051,N_5170);
xnor U6018 (N_6018,N_5501,N_5012);
xor U6019 (N_6019,N_5684,N_5007);
nand U6020 (N_6020,N_5371,N_5058);
and U6021 (N_6021,N_5927,N_5982);
and U6022 (N_6022,N_5097,N_5681);
nand U6023 (N_6023,N_5389,N_5416);
nand U6024 (N_6024,N_5333,N_5728);
nand U6025 (N_6025,N_5052,N_5537);
nor U6026 (N_6026,N_5492,N_5809);
nand U6027 (N_6027,N_5509,N_5615);
nor U6028 (N_6028,N_5125,N_5308);
xnor U6029 (N_6029,N_5486,N_5450);
and U6030 (N_6030,N_5461,N_5337);
nor U6031 (N_6031,N_5663,N_5730);
nor U6032 (N_6032,N_5890,N_5251);
nor U6033 (N_6033,N_5570,N_5104);
nor U6034 (N_6034,N_5664,N_5600);
and U6035 (N_6035,N_5522,N_5993);
or U6036 (N_6036,N_5448,N_5855);
xor U6037 (N_6037,N_5873,N_5519);
or U6038 (N_6038,N_5082,N_5395);
nor U6039 (N_6039,N_5704,N_5628);
nand U6040 (N_6040,N_5422,N_5294);
xor U6041 (N_6041,N_5240,N_5971);
xor U6042 (N_6042,N_5306,N_5036);
xor U6043 (N_6043,N_5933,N_5760);
nand U6044 (N_6044,N_5277,N_5215);
nand U6045 (N_6045,N_5310,N_5493);
nor U6046 (N_6046,N_5881,N_5188);
nand U6047 (N_6047,N_5192,N_5008);
and U6048 (N_6048,N_5987,N_5559);
and U6049 (N_6049,N_5099,N_5633);
nor U6050 (N_6050,N_5382,N_5604);
nand U6051 (N_6051,N_5405,N_5617);
and U6052 (N_6052,N_5153,N_5652);
xor U6053 (N_6053,N_5981,N_5388);
and U6054 (N_6054,N_5943,N_5568);
or U6055 (N_6055,N_5410,N_5980);
nand U6056 (N_6056,N_5949,N_5607);
nand U6057 (N_6057,N_5752,N_5683);
or U6058 (N_6058,N_5466,N_5169);
xor U6059 (N_6059,N_5092,N_5489);
nand U6060 (N_6060,N_5123,N_5619);
xnor U6061 (N_6061,N_5019,N_5204);
and U6062 (N_6062,N_5222,N_5849);
and U6063 (N_6063,N_5866,N_5363);
or U6064 (N_6064,N_5290,N_5361);
nor U6065 (N_6065,N_5733,N_5920);
xor U6066 (N_6066,N_5673,N_5187);
nor U6067 (N_6067,N_5707,N_5770);
xnor U6068 (N_6068,N_5546,N_5912);
and U6069 (N_6069,N_5136,N_5198);
or U6070 (N_6070,N_5751,N_5321);
xor U6071 (N_6071,N_5236,N_5780);
nor U6072 (N_6072,N_5721,N_5374);
and U6073 (N_6073,N_5483,N_5699);
xor U6074 (N_6074,N_5861,N_5490);
nand U6075 (N_6075,N_5259,N_5112);
or U6076 (N_6076,N_5938,N_5762);
nor U6077 (N_6077,N_5576,N_5850);
nor U6078 (N_6078,N_5117,N_5747);
nand U6079 (N_6079,N_5909,N_5364);
xnor U6080 (N_6080,N_5426,N_5494);
nor U6081 (N_6081,N_5984,N_5391);
nand U6082 (N_6082,N_5063,N_5709);
nand U6083 (N_6083,N_5022,N_5465);
nor U6084 (N_6084,N_5841,N_5015);
xor U6085 (N_6085,N_5075,N_5275);
and U6086 (N_6086,N_5788,N_5667);
nand U6087 (N_6087,N_5696,N_5803);
xor U6088 (N_6088,N_5285,N_5379);
nor U6089 (N_6089,N_5503,N_5550);
and U6090 (N_6090,N_5918,N_5009);
xor U6091 (N_6091,N_5393,N_5038);
nand U6092 (N_6092,N_5655,N_5280);
xnor U6093 (N_6093,N_5304,N_5901);
or U6094 (N_6094,N_5074,N_5767);
xor U6095 (N_6095,N_5342,N_5247);
nor U6096 (N_6096,N_5487,N_5032);
nand U6097 (N_6097,N_5710,N_5228);
nand U6098 (N_6098,N_5394,N_5078);
or U6099 (N_6099,N_5232,N_5133);
or U6100 (N_6100,N_5851,N_5556);
nand U6101 (N_6101,N_5557,N_5161);
nor U6102 (N_6102,N_5772,N_5206);
and U6103 (N_6103,N_5879,N_5497);
and U6104 (N_6104,N_5553,N_5723);
nor U6105 (N_6105,N_5962,N_5138);
or U6106 (N_6106,N_5406,N_5440);
and U6107 (N_6107,N_5902,N_5155);
and U6108 (N_6108,N_5249,N_5857);
or U6109 (N_6109,N_5241,N_5053);
or U6110 (N_6110,N_5965,N_5224);
xnor U6111 (N_6111,N_5287,N_5647);
xnor U6112 (N_6112,N_5024,N_5846);
nor U6113 (N_6113,N_5442,N_5402);
xor U6114 (N_6114,N_5336,N_5544);
nor U6115 (N_6115,N_5985,N_5941);
nor U6116 (N_6116,N_5343,N_5047);
nor U6117 (N_6117,N_5675,N_5531);
and U6118 (N_6118,N_5330,N_5184);
or U6119 (N_6119,N_5037,N_5590);
or U6120 (N_6120,N_5460,N_5937);
nand U6121 (N_6121,N_5844,N_5334);
xor U6122 (N_6122,N_5835,N_5495);
nor U6123 (N_6123,N_5609,N_5635);
nand U6124 (N_6124,N_5441,N_5484);
nor U6125 (N_6125,N_5235,N_5423);
nor U6126 (N_6126,N_5740,N_5404);
and U6127 (N_6127,N_5346,N_5976);
and U6128 (N_6128,N_5739,N_5479);
xnor U6129 (N_6129,N_5477,N_5087);
nand U6130 (N_6130,N_5071,N_5292);
nand U6131 (N_6131,N_5606,N_5716);
and U6132 (N_6132,N_5457,N_5164);
and U6133 (N_6133,N_5515,N_5952);
and U6134 (N_6134,N_5476,N_5620);
and U6135 (N_6135,N_5118,N_5973);
and U6136 (N_6136,N_5313,N_5961);
nand U6137 (N_6137,N_5676,N_5282);
nor U6138 (N_6138,N_5877,N_5349);
xnor U6139 (N_6139,N_5613,N_5250);
or U6140 (N_6140,N_5725,N_5482);
and U6141 (N_6141,N_5666,N_5623);
or U6142 (N_6142,N_5350,N_5936);
or U6143 (N_6143,N_5535,N_5209);
xnor U6144 (N_6144,N_5843,N_5002);
or U6145 (N_6145,N_5812,N_5614);
xnor U6146 (N_6146,N_5447,N_5540);
or U6147 (N_6147,N_5376,N_5714);
nor U6148 (N_6148,N_5425,N_5372);
or U6149 (N_6149,N_5814,N_5318);
or U6150 (N_6150,N_5171,N_5565);
and U6151 (N_6151,N_5791,N_5265);
and U6152 (N_6152,N_5654,N_5194);
or U6153 (N_6153,N_5094,N_5778);
and U6154 (N_6154,N_5252,N_5335);
xnor U6155 (N_6155,N_5820,N_5945);
or U6156 (N_6156,N_5642,N_5705);
and U6157 (N_6157,N_5419,N_5225);
nor U6158 (N_6158,N_5929,N_5889);
or U6159 (N_6159,N_5883,N_5512);
nand U6160 (N_6160,N_5946,N_5745);
or U6161 (N_6161,N_5473,N_5256);
and U6162 (N_6162,N_5758,N_5650);
nor U6163 (N_6163,N_5988,N_5935);
xnor U6164 (N_6164,N_5491,N_5924);
nand U6165 (N_6165,N_5808,N_5178);
or U6166 (N_6166,N_5864,N_5689);
or U6167 (N_6167,N_5862,N_5817);
and U6168 (N_6168,N_5514,N_5320);
or U6169 (N_6169,N_5338,N_5355);
or U6170 (N_6170,N_5102,N_5880);
and U6171 (N_6171,N_5197,N_5746);
or U6172 (N_6172,N_5401,N_5795);
or U6173 (N_6173,N_5828,N_5212);
nand U6174 (N_6174,N_5339,N_5692);
or U6175 (N_6175,N_5970,N_5034);
xor U6176 (N_6176,N_5827,N_5884);
nand U6177 (N_6177,N_5967,N_5000);
or U6178 (N_6178,N_5646,N_5124);
xnor U6179 (N_6179,N_5056,N_5627);
nor U6180 (N_6180,N_5621,N_5602);
xor U6181 (N_6181,N_5975,N_5631);
nor U6182 (N_6182,N_5387,N_5288);
or U6183 (N_6183,N_5694,N_5738);
nand U6184 (N_6184,N_5083,N_5048);
and U6185 (N_6185,N_5831,N_5734);
nor U6186 (N_6186,N_5854,N_5947);
and U6187 (N_6187,N_5765,N_5014);
or U6188 (N_6188,N_5977,N_5407);
or U6189 (N_6189,N_5129,N_5160);
or U6190 (N_6190,N_5311,N_5584);
nor U6191 (N_6191,N_5324,N_5090);
and U6192 (N_6192,N_5594,N_5412);
nand U6193 (N_6193,N_5640,N_5260);
nand U6194 (N_6194,N_5016,N_5582);
nor U6195 (N_6195,N_5166,N_5549);
xor U6196 (N_6196,N_5586,N_5253);
and U6197 (N_6197,N_5792,N_5701);
and U6198 (N_6198,N_5291,N_5325);
or U6199 (N_6199,N_5378,N_5892);
nand U6200 (N_6200,N_5896,N_5305);
and U6201 (N_6201,N_5498,N_5470);
xor U6202 (N_6202,N_5688,N_5216);
and U6203 (N_6203,N_5598,N_5181);
nor U6204 (N_6204,N_5695,N_5579);
or U6205 (N_6205,N_5352,N_5648);
and U6206 (N_6206,N_5932,N_5370);
nand U6207 (N_6207,N_5951,N_5906);
nor U6208 (N_6208,N_5934,N_5830);
and U6209 (N_6209,N_5567,N_5543);
xnor U6210 (N_6210,N_5532,N_5233);
xnor U6211 (N_6211,N_5541,N_5524);
or U6212 (N_6212,N_5496,N_5528);
nor U6213 (N_6213,N_5757,N_5079);
xor U6214 (N_6214,N_5454,N_5298);
nand U6215 (N_6215,N_5399,N_5774);
or U6216 (N_6216,N_5042,N_5044);
and U6217 (N_6217,N_5357,N_5122);
nor U6218 (N_6218,N_5536,N_5601);
and U6219 (N_6219,N_5173,N_5213);
nor U6220 (N_6220,N_5467,N_5891);
and U6221 (N_6221,N_5756,N_5319);
nand U6222 (N_6222,N_5560,N_5061);
nor U6223 (N_6223,N_5070,N_5469);
xnor U6224 (N_6224,N_5326,N_5574);
and U6225 (N_6225,N_5089,N_5886);
xnor U6226 (N_6226,N_5972,N_5383);
nor U6227 (N_6227,N_5203,N_5182);
and U6228 (N_6228,N_5358,N_5997);
xnor U6229 (N_6229,N_5919,N_5622);
xor U6230 (N_6230,N_5651,N_5869);
xor U6231 (N_6231,N_5093,N_5353);
nor U6232 (N_6232,N_5775,N_5013);
or U6233 (N_6233,N_5750,N_5858);
xnor U6234 (N_6234,N_5086,N_5508);
nor U6235 (N_6235,N_5793,N_5020);
and U6236 (N_6236,N_5159,N_5452);
nor U6237 (N_6237,N_5996,N_5800);
nand U6238 (N_6238,N_5922,N_5668);
nor U6239 (N_6239,N_5715,N_5429);
nor U6240 (N_6240,N_5871,N_5766);
and U6241 (N_6241,N_5659,N_5882);
nand U6242 (N_6242,N_5424,N_5433);
and U6243 (N_6243,N_5764,N_5327);
xnor U6244 (N_6244,N_5768,N_5107);
nand U6245 (N_6245,N_5045,N_5787);
nand U6246 (N_6246,N_5572,N_5255);
nand U6247 (N_6247,N_5773,N_5183);
nor U6248 (N_6248,N_5273,N_5816);
nand U6249 (N_6249,N_5526,N_5966);
or U6250 (N_6250,N_5571,N_5995);
and U6251 (N_6251,N_5834,N_5340);
nor U6252 (N_6252,N_5610,N_5103);
nand U6253 (N_6253,N_5776,N_5026);
nor U6254 (N_6254,N_5296,N_5040);
and U6255 (N_6255,N_5521,N_5811);
nand U6256 (N_6256,N_5234,N_5077);
or U6257 (N_6257,N_5096,N_5067);
xnor U6258 (N_6258,N_5113,N_5120);
nor U6259 (N_6259,N_5630,N_5964);
nand U6260 (N_6260,N_5525,N_5989);
nand U6261 (N_6261,N_5926,N_5438);
or U6262 (N_6262,N_5106,N_5175);
and U6263 (N_6263,N_5345,N_5185);
nor U6264 (N_6264,N_5639,N_5281);
and U6265 (N_6265,N_5069,N_5580);
xnor U6266 (N_6266,N_5848,N_5208);
and U6267 (N_6267,N_5930,N_5210);
xnor U6268 (N_6268,N_5436,N_5231);
nor U6269 (N_6269,N_5904,N_5748);
nor U6270 (N_6270,N_5687,N_5561);
or U6271 (N_6271,N_5144,N_5202);
and U6272 (N_6272,N_5832,N_5468);
or U6273 (N_6273,N_5146,N_5944);
or U6274 (N_6274,N_5218,N_5948);
nor U6275 (N_6275,N_5242,N_5505);
nand U6276 (N_6276,N_5868,N_5779);
nor U6277 (N_6277,N_5332,N_5769);
nor U6278 (N_6278,N_5307,N_5786);
xor U6279 (N_6279,N_5035,N_5511);
and U6280 (N_6280,N_5867,N_5471);
xor U6281 (N_6281,N_5270,N_5819);
xnor U6282 (N_6282,N_5785,N_5520);
and U6283 (N_6283,N_5366,N_5805);
nand U6284 (N_6284,N_5116,N_5076);
xnor U6285 (N_6285,N_5907,N_5421);
nor U6286 (N_6286,N_5916,N_5711);
and U6287 (N_6287,N_5434,N_5480);
and U6288 (N_6288,N_5720,N_5727);
nor U6289 (N_6289,N_5804,N_5749);
xor U6290 (N_6290,N_5417,N_5529);
and U6291 (N_6291,N_5088,N_5824);
nand U6292 (N_6292,N_5697,N_5518);
or U6293 (N_6293,N_5799,N_5592);
and U6294 (N_6294,N_5027,N_5736);
nor U6295 (N_6295,N_5428,N_5563);
or U6296 (N_6296,N_5140,N_5073);
nand U6297 (N_6297,N_5878,N_5744);
or U6298 (N_6298,N_5743,N_5612);
and U6299 (N_6299,N_5176,N_5322);
nor U6300 (N_6300,N_5978,N_5196);
or U6301 (N_6301,N_5564,N_5794);
xnor U6302 (N_6302,N_5569,N_5653);
and U6303 (N_6303,N_5057,N_5264);
and U6304 (N_6304,N_5829,N_5547);
nand U6305 (N_6305,N_5085,N_5152);
or U6306 (N_6306,N_5205,N_5380);
or U6307 (N_6307,N_5128,N_5925);
nand U6308 (N_6308,N_5712,N_5685);
nand U6309 (N_6309,N_5478,N_5825);
nand U6310 (N_6310,N_5006,N_5451);
and U6311 (N_6311,N_5999,N_5453);
and U6312 (N_6312,N_5992,N_5297);
xor U6313 (N_6313,N_5905,N_5545);
xor U6314 (N_6314,N_5023,N_5810);
nand U6315 (N_6315,N_5356,N_5017);
xor U6316 (N_6316,N_5254,N_5789);
and U6317 (N_6317,N_5777,N_5645);
nand U6318 (N_6318,N_5151,N_5554);
or U6319 (N_6319,N_5735,N_5286);
nand U6320 (N_6320,N_5657,N_5068);
nor U6321 (N_6321,N_5656,N_5258);
nand U6322 (N_6322,N_5269,N_5143);
or U6323 (N_6323,N_5761,N_5921);
or U6324 (N_6324,N_5499,N_5134);
nor U6325 (N_6325,N_5899,N_5797);
and U6326 (N_6326,N_5029,N_5360);
or U6327 (N_6327,N_5616,N_5940);
nor U6328 (N_6328,N_5162,N_5859);
nor U6329 (N_6329,N_5900,N_5227);
and U6330 (N_6330,N_5534,N_5672);
and U6331 (N_6331,N_5163,N_5367);
and U6332 (N_6332,N_5516,N_5986);
xnor U6333 (N_6333,N_5003,N_5806);
nand U6334 (N_6334,N_5312,N_5953);
and U6335 (N_6335,N_5180,N_5158);
nor U6336 (N_6336,N_5662,N_5888);
or U6337 (N_6337,N_5599,N_5548);
or U6338 (N_6338,N_5132,N_5413);
nor U6339 (N_6339,N_5538,N_5605);
and U6340 (N_6340,N_5121,N_5510);
nor U6341 (N_6341,N_5010,N_5875);
nand U6342 (N_6342,N_5135,N_5475);
nor U6343 (N_6343,N_5507,N_5415);
xor U6344 (N_6344,N_5137,N_5481);
or U6345 (N_6345,N_5649,N_5098);
or U6346 (N_6346,N_5865,N_5959);
or U6347 (N_6347,N_5046,N_5573);
and U6348 (N_6348,N_5359,N_5464);
and U6349 (N_6349,N_5798,N_5969);
nor U6350 (N_6350,N_5018,N_5065);
xor U6351 (N_6351,N_5392,N_5243);
or U6352 (N_6352,N_5950,N_5983);
xor U6353 (N_6353,N_5502,N_5317);
nand U6354 (N_6354,N_5894,N_5271);
or U6355 (N_6355,N_5539,N_5062);
nand U6356 (N_6356,N_5011,N_5130);
nor U6357 (N_6357,N_5221,N_5638);
nand U6358 (N_6358,N_5643,N_5914);
nor U6359 (N_6359,N_5119,N_5462);
and U6360 (N_6360,N_5669,N_5726);
and U6361 (N_6361,N_5753,N_5431);
and U6362 (N_6362,N_5276,N_5691);
and U6363 (N_6363,N_5245,N_5084);
or U6364 (N_6364,N_5368,N_5837);
or U6365 (N_6365,N_5049,N_5703);
xor U6366 (N_6366,N_5958,N_5239);
or U6367 (N_6367,N_5398,N_5729);
nor U6368 (N_6368,N_5303,N_5558);
nor U6369 (N_6369,N_5080,N_5870);
and U6370 (N_6370,N_5028,N_5913);
and U6371 (N_6371,N_5853,N_5001);
nor U6372 (N_6372,N_5167,N_5437);
nor U6373 (N_6373,N_5636,N_5755);
or U6374 (N_6374,N_5737,N_5267);
or U6375 (N_6375,N_5066,N_5004);
xnor U6376 (N_6376,N_5742,N_5148);
xnor U6377 (N_6377,N_5390,N_5377);
or U6378 (N_6378,N_5211,N_5634);
xnor U6379 (N_6379,N_5724,N_5229);
xnor U6380 (N_6380,N_5990,N_5172);
and U6381 (N_6381,N_5408,N_5637);
nor U6382 (N_6382,N_5455,N_5095);
or U6383 (N_6383,N_5690,N_5575);
xor U6384 (N_6384,N_5386,N_5149);
xor U6385 (N_6385,N_5939,N_5081);
nand U6386 (N_6386,N_5513,N_5845);
xnor U6387 (N_6387,N_5385,N_5677);
xnor U6388 (N_6388,N_5555,N_5456);
nor U6389 (N_6389,N_5472,N_5551);
and U6390 (N_6390,N_5754,N_5396);
nor U6391 (N_6391,N_5674,N_5917);
xor U6392 (N_6392,N_5329,N_5856);
xor U6393 (N_6393,N_5446,N_5847);
and U6394 (N_6394,N_5177,N_5956);
xor U6395 (N_6395,N_5141,N_5246);
or U6396 (N_6396,N_5562,N_5384);
or U6397 (N_6397,N_5566,N_5315);
xor U6398 (N_6398,N_5801,N_5400);
and U6399 (N_6399,N_5860,N_5109);
nand U6400 (N_6400,N_5373,N_5108);
or U6401 (N_6401,N_5488,N_5238);
or U6402 (N_6402,N_5348,N_5409);
or U6403 (N_6403,N_5459,N_5781);
and U6404 (N_6404,N_5091,N_5100);
xnor U6405 (N_6405,N_5443,N_5043);
xnor U6406 (N_6406,N_5186,N_5836);
nor U6407 (N_6407,N_5289,N_5527);
nand U6408 (N_6408,N_5702,N_5449);
or U6409 (N_6409,N_5299,N_5991);
xnor U6410 (N_6410,N_5105,N_5272);
nor U6411 (N_6411,N_5583,N_5577);
and U6412 (N_6412,N_5369,N_5552);
or U6413 (N_6413,N_5974,N_5603);
and U6414 (N_6414,N_5041,N_5915);
nand U6415 (N_6415,N_5807,N_5581);
nor U6416 (N_6416,N_5826,N_5782);
or U6417 (N_6417,N_5191,N_5790);
nor U6418 (N_6418,N_5517,N_5686);
and U6419 (N_6419,N_5230,N_5126);
nor U6420 (N_6420,N_5223,N_5055);
nand U6421 (N_6421,N_5365,N_5608);
nor U6422 (N_6422,N_5874,N_5968);
xor U6423 (N_6423,N_5427,N_5611);
xnor U6424 (N_6424,N_5833,N_5059);
xor U6425 (N_6425,N_5852,N_5025);
and U6426 (N_6426,N_5375,N_5226);
and U6427 (N_6427,N_5114,N_5911);
nand U6428 (N_6428,N_5179,N_5718);
nand U6429 (N_6429,N_5033,N_5219);
and U6430 (N_6430,N_5439,N_5923);
or U6431 (N_6431,N_5821,N_5403);
nor U6432 (N_6432,N_5813,N_5054);
and U6433 (N_6433,N_5485,N_5713);
or U6434 (N_6434,N_5698,N_5931);
and U6435 (N_6435,N_5381,N_5876);
nand U6436 (N_6436,N_5597,N_5641);
nor U6437 (N_6437,N_5463,N_5717);
or U6438 (N_6438,N_5237,N_5895);
nor U6439 (N_6439,N_5266,N_5110);
xor U6440 (N_6440,N_5295,N_5131);
nand U6441 (N_6441,N_5261,N_5588);
nor U6442 (N_6442,N_5351,N_5822);
nor U6443 (N_6443,N_5005,N_5618);
nand U6444 (N_6444,N_5928,N_5523);
nand U6445 (N_6445,N_5587,N_5199);
or U6446 (N_6446,N_5154,N_5021);
or U6447 (N_6447,N_5629,N_5771);
and U6448 (N_6448,N_5474,N_5397);
and U6449 (N_6449,N_5220,N_5957);
and U6450 (N_6450,N_5435,N_5127);
and U6451 (N_6451,N_5839,N_5411);
nor U6452 (N_6452,N_5139,N_5217);
nor U6453 (N_6453,N_5101,N_5626);
xnor U6454 (N_6454,N_5840,N_5578);
nand U6455 (N_6455,N_5072,N_5998);
or U6456 (N_6456,N_5644,N_5362);
or U6457 (N_6457,N_5284,N_5838);
nand U6458 (N_6458,N_5354,N_5418);
nand U6459 (N_6459,N_5624,N_5979);
nand U6460 (N_6460,N_5504,N_5189);
nand U6461 (N_6461,N_5145,N_5328);
nor U6462 (N_6462,N_5300,N_5314);
nor U6463 (N_6463,N_5731,N_5309);
or U6464 (N_6464,N_5910,N_5706);
nand U6465 (N_6465,N_5030,N_5165);
and U6466 (N_6466,N_5262,N_5050);
and U6467 (N_6467,N_5708,N_5671);
nor U6468 (N_6468,N_5784,N_5625);
nand U6469 (N_6469,N_5283,N_5783);
or U6470 (N_6470,N_5908,N_5500);
nor U6471 (N_6471,N_5887,N_5670);
nor U6472 (N_6472,N_5530,N_5060);
and U6473 (N_6473,N_5064,N_5682);
or U6474 (N_6474,N_5542,N_5039);
and U6475 (N_6475,N_5722,N_5142);
nor U6476 (N_6476,N_5195,N_5963);
and U6477 (N_6477,N_5960,N_5818);
or U6478 (N_6478,N_5759,N_5414);
xor U6479 (N_6479,N_5863,N_5903);
nand U6480 (N_6480,N_5897,N_5658);
xnor U6481 (N_6481,N_5533,N_5693);
nand U6482 (N_6482,N_5323,N_5591);
or U6483 (N_6483,N_5293,N_5898);
and U6484 (N_6484,N_5214,N_5147);
xor U6485 (N_6485,N_5150,N_5815);
nand U6486 (N_6486,N_5268,N_5430);
xor U6487 (N_6487,N_5278,N_5301);
nand U6488 (N_6488,N_5741,N_5665);
nand U6489 (N_6489,N_5316,N_5589);
nor U6490 (N_6490,N_5420,N_5257);
nand U6491 (N_6491,N_5174,N_5678);
nand U6492 (N_6492,N_5331,N_5719);
and U6493 (N_6493,N_5302,N_5954);
and U6494 (N_6494,N_5263,N_5201);
or U6495 (N_6495,N_5341,N_5168);
or U6496 (N_6496,N_5955,N_5157);
xnor U6497 (N_6497,N_5680,N_5115);
nand U6498 (N_6498,N_5444,N_5885);
nand U6499 (N_6499,N_5596,N_5732);
nor U6500 (N_6500,N_5455,N_5713);
nand U6501 (N_6501,N_5322,N_5342);
and U6502 (N_6502,N_5094,N_5727);
and U6503 (N_6503,N_5439,N_5496);
or U6504 (N_6504,N_5568,N_5926);
or U6505 (N_6505,N_5669,N_5933);
xnor U6506 (N_6506,N_5393,N_5239);
xor U6507 (N_6507,N_5062,N_5498);
nand U6508 (N_6508,N_5638,N_5401);
nor U6509 (N_6509,N_5969,N_5431);
or U6510 (N_6510,N_5905,N_5383);
xor U6511 (N_6511,N_5253,N_5060);
xor U6512 (N_6512,N_5585,N_5119);
xnor U6513 (N_6513,N_5155,N_5936);
nand U6514 (N_6514,N_5055,N_5126);
xor U6515 (N_6515,N_5284,N_5678);
xnor U6516 (N_6516,N_5838,N_5055);
xnor U6517 (N_6517,N_5593,N_5806);
nor U6518 (N_6518,N_5108,N_5735);
nand U6519 (N_6519,N_5073,N_5324);
xor U6520 (N_6520,N_5505,N_5620);
xnor U6521 (N_6521,N_5960,N_5697);
nor U6522 (N_6522,N_5381,N_5501);
and U6523 (N_6523,N_5588,N_5556);
xor U6524 (N_6524,N_5270,N_5565);
nor U6525 (N_6525,N_5938,N_5096);
or U6526 (N_6526,N_5246,N_5438);
xnor U6527 (N_6527,N_5227,N_5370);
nand U6528 (N_6528,N_5980,N_5994);
nand U6529 (N_6529,N_5305,N_5467);
and U6530 (N_6530,N_5878,N_5953);
nor U6531 (N_6531,N_5551,N_5883);
or U6532 (N_6532,N_5076,N_5659);
xnor U6533 (N_6533,N_5974,N_5820);
or U6534 (N_6534,N_5696,N_5860);
nor U6535 (N_6535,N_5115,N_5622);
nor U6536 (N_6536,N_5671,N_5712);
nor U6537 (N_6537,N_5952,N_5386);
xor U6538 (N_6538,N_5658,N_5462);
and U6539 (N_6539,N_5858,N_5991);
nand U6540 (N_6540,N_5572,N_5616);
nor U6541 (N_6541,N_5020,N_5953);
or U6542 (N_6542,N_5952,N_5533);
nor U6543 (N_6543,N_5834,N_5226);
nor U6544 (N_6544,N_5938,N_5185);
xnor U6545 (N_6545,N_5647,N_5160);
or U6546 (N_6546,N_5186,N_5440);
nand U6547 (N_6547,N_5859,N_5214);
nand U6548 (N_6548,N_5862,N_5624);
nor U6549 (N_6549,N_5195,N_5466);
nand U6550 (N_6550,N_5668,N_5901);
and U6551 (N_6551,N_5307,N_5768);
and U6552 (N_6552,N_5797,N_5746);
and U6553 (N_6553,N_5195,N_5307);
or U6554 (N_6554,N_5527,N_5680);
nand U6555 (N_6555,N_5908,N_5564);
or U6556 (N_6556,N_5845,N_5156);
or U6557 (N_6557,N_5424,N_5331);
or U6558 (N_6558,N_5939,N_5348);
xor U6559 (N_6559,N_5199,N_5283);
xnor U6560 (N_6560,N_5024,N_5900);
xor U6561 (N_6561,N_5955,N_5144);
xor U6562 (N_6562,N_5002,N_5982);
and U6563 (N_6563,N_5482,N_5860);
nor U6564 (N_6564,N_5159,N_5588);
xnor U6565 (N_6565,N_5394,N_5102);
or U6566 (N_6566,N_5914,N_5634);
nand U6567 (N_6567,N_5192,N_5073);
nor U6568 (N_6568,N_5157,N_5911);
nand U6569 (N_6569,N_5208,N_5967);
nand U6570 (N_6570,N_5477,N_5611);
nor U6571 (N_6571,N_5803,N_5336);
nand U6572 (N_6572,N_5054,N_5080);
nor U6573 (N_6573,N_5989,N_5826);
and U6574 (N_6574,N_5829,N_5563);
xnor U6575 (N_6575,N_5951,N_5845);
nand U6576 (N_6576,N_5641,N_5062);
or U6577 (N_6577,N_5731,N_5440);
and U6578 (N_6578,N_5709,N_5225);
nor U6579 (N_6579,N_5365,N_5683);
or U6580 (N_6580,N_5451,N_5160);
and U6581 (N_6581,N_5529,N_5005);
and U6582 (N_6582,N_5817,N_5143);
xor U6583 (N_6583,N_5156,N_5381);
and U6584 (N_6584,N_5727,N_5168);
or U6585 (N_6585,N_5309,N_5654);
nand U6586 (N_6586,N_5116,N_5236);
and U6587 (N_6587,N_5162,N_5026);
and U6588 (N_6588,N_5668,N_5857);
xor U6589 (N_6589,N_5150,N_5498);
nand U6590 (N_6590,N_5720,N_5833);
nor U6591 (N_6591,N_5412,N_5161);
and U6592 (N_6592,N_5325,N_5983);
nor U6593 (N_6593,N_5785,N_5939);
and U6594 (N_6594,N_5980,N_5959);
xor U6595 (N_6595,N_5783,N_5826);
nor U6596 (N_6596,N_5445,N_5749);
xnor U6597 (N_6597,N_5297,N_5021);
nor U6598 (N_6598,N_5698,N_5298);
nor U6599 (N_6599,N_5548,N_5508);
or U6600 (N_6600,N_5646,N_5117);
nor U6601 (N_6601,N_5374,N_5348);
nor U6602 (N_6602,N_5915,N_5695);
or U6603 (N_6603,N_5448,N_5188);
nand U6604 (N_6604,N_5774,N_5223);
and U6605 (N_6605,N_5106,N_5062);
nand U6606 (N_6606,N_5026,N_5441);
xnor U6607 (N_6607,N_5869,N_5935);
or U6608 (N_6608,N_5085,N_5015);
nand U6609 (N_6609,N_5487,N_5991);
and U6610 (N_6610,N_5165,N_5796);
nand U6611 (N_6611,N_5690,N_5060);
nor U6612 (N_6612,N_5269,N_5023);
nand U6613 (N_6613,N_5647,N_5517);
nand U6614 (N_6614,N_5250,N_5983);
nor U6615 (N_6615,N_5642,N_5809);
xor U6616 (N_6616,N_5625,N_5481);
or U6617 (N_6617,N_5043,N_5392);
nor U6618 (N_6618,N_5868,N_5008);
or U6619 (N_6619,N_5005,N_5396);
nor U6620 (N_6620,N_5649,N_5349);
and U6621 (N_6621,N_5780,N_5071);
nand U6622 (N_6622,N_5793,N_5149);
nand U6623 (N_6623,N_5784,N_5226);
nand U6624 (N_6624,N_5991,N_5282);
nor U6625 (N_6625,N_5905,N_5591);
nand U6626 (N_6626,N_5396,N_5427);
nand U6627 (N_6627,N_5900,N_5813);
nand U6628 (N_6628,N_5711,N_5027);
xnor U6629 (N_6629,N_5973,N_5465);
nand U6630 (N_6630,N_5323,N_5393);
nor U6631 (N_6631,N_5154,N_5935);
xnor U6632 (N_6632,N_5896,N_5443);
and U6633 (N_6633,N_5960,N_5952);
nor U6634 (N_6634,N_5845,N_5656);
or U6635 (N_6635,N_5269,N_5939);
nand U6636 (N_6636,N_5697,N_5103);
nor U6637 (N_6637,N_5835,N_5262);
or U6638 (N_6638,N_5831,N_5409);
and U6639 (N_6639,N_5053,N_5057);
nor U6640 (N_6640,N_5869,N_5245);
nand U6641 (N_6641,N_5976,N_5592);
xor U6642 (N_6642,N_5040,N_5597);
or U6643 (N_6643,N_5106,N_5790);
nor U6644 (N_6644,N_5156,N_5565);
nor U6645 (N_6645,N_5925,N_5032);
xor U6646 (N_6646,N_5788,N_5750);
and U6647 (N_6647,N_5215,N_5073);
nand U6648 (N_6648,N_5061,N_5746);
nand U6649 (N_6649,N_5828,N_5520);
nand U6650 (N_6650,N_5647,N_5434);
or U6651 (N_6651,N_5397,N_5582);
nand U6652 (N_6652,N_5497,N_5116);
xor U6653 (N_6653,N_5138,N_5733);
nor U6654 (N_6654,N_5879,N_5323);
nand U6655 (N_6655,N_5961,N_5911);
and U6656 (N_6656,N_5325,N_5264);
and U6657 (N_6657,N_5404,N_5729);
nand U6658 (N_6658,N_5830,N_5676);
nor U6659 (N_6659,N_5162,N_5172);
or U6660 (N_6660,N_5355,N_5897);
xnor U6661 (N_6661,N_5703,N_5063);
xor U6662 (N_6662,N_5476,N_5379);
and U6663 (N_6663,N_5309,N_5944);
nor U6664 (N_6664,N_5241,N_5174);
or U6665 (N_6665,N_5008,N_5021);
and U6666 (N_6666,N_5506,N_5999);
or U6667 (N_6667,N_5728,N_5780);
nand U6668 (N_6668,N_5856,N_5004);
xor U6669 (N_6669,N_5804,N_5289);
nand U6670 (N_6670,N_5981,N_5365);
nor U6671 (N_6671,N_5802,N_5511);
nand U6672 (N_6672,N_5608,N_5827);
and U6673 (N_6673,N_5510,N_5890);
nand U6674 (N_6674,N_5147,N_5690);
and U6675 (N_6675,N_5719,N_5956);
xnor U6676 (N_6676,N_5420,N_5806);
nand U6677 (N_6677,N_5909,N_5725);
nor U6678 (N_6678,N_5524,N_5216);
nor U6679 (N_6679,N_5185,N_5339);
xor U6680 (N_6680,N_5496,N_5206);
xnor U6681 (N_6681,N_5737,N_5429);
xnor U6682 (N_6682,N_5966,N_5554);
nand U6683 (N_6683,N_5358,N_5592);
or U6684 (N_6684,N_5789,N_5596);
nand U6685 (N_6685,N_5779,N_5547);
nand U6686 (N_6686,N_5239,N_5773);
and U6687 (N_6687,N_5124,N_5500);
and U6688 (N_6688,N_5359,N_5452);
and U6689 (N_6689,N_5584,N_5686);
or U6690 (N_6690,N_5126,N_5019);
or U6691 (N_6691,N_5838,N_5107);
nor U6692 (N_6692,N_5947,N_5743);
and U6693 (N_6693,N_5290,N_5278);
xnor U6694 (N_6694,N_5475,N_5825);
or U6695 (N_6695,N_5334,N_5788);
nand U6696 (N_6696,N_5111,N_5065);
nand U6697 (N_6697,N_5523,N_5627);
and U6698 (N_6698,N_5684,N_5432);
and U6699 (N_6699,N_5313,N_5318);
or U6700 (N_6700,N_5312,N_5581);
or U6701 (N_6701,N_5778,N_5007);
or U6702 (N_6702,N_5641,N_5240);
and U6703 (N_6703,N_5144,N_5727);
nand U6704 (N_6704,N_5568,N_5482);
or U6705 (N_6705,N_5737,N_5102);
nand U6706 (N_6706,N_5698,N_5452);
or U6707 (N_6707,N_5328,N_5999);
or U6708 (N_6708,N_5341,N_5361);
xor U6709 (N_6709,N_5919,N_5831);
xnor U6710 (N_6710,N_5715,N_5064);
and U6711 (N_6711,N_5849,N_5256);
nand U6712 (N_6712,N_5699,N_5551);
and U6713 (N_6713,N_5294,N_5405);
nand U6714 (N_6714,N_5260,N_5975);
nor U6715 (N_6715,N_5566,N_5506);
xnor U6716 (N_6716,N_5518,N_5567);
or U6717 (N_6717,N_5450,N_5780);
or U6718 (N_6718,N_5769,N_5547);
nand U6719 (N_6719,N_5997,N_5749);
or U6720 (N_6720,N_5747,N_5751);
nand U6721 (N_6721,N_5737,N_5647);
nand U6722 (N_6722,N_5827,N_5136);
xnor U6723 (N_6723,N_5992,N_5951);
xnor U6724 (N_6724,N_5297,N_5966);
nand U6725 (N_6725,N_5638,N_5452);
and U6726 (N_6726,N_5413,N_5248);
xor U6727 (N_6727,N_5179,N_5598);
nor U6728 (N_6728,N_5967,N_5730);
nor U6729 (N_6729,N_5809,N_5050);
nor U6730 (N_6730,N_5433,N_5305);
nand U6731 (N_6731,N_5989,N_5099);
xnor U6732 (N_6732,N_5866,N_5003);
xor U6733 (N_6733,N_5945,N_5554);
nor U6734 (N_6734,N_5083,N_5218);
and U6735 (N_6735,N_5270,N_5185);
and U6736 (N_6736,N_5132,N_5266);
xor U6737 (N_6737,N_5210,N_5367);
and U6738 (N_6738,N_5112,N_5354);
and U6739 (N_6739,N_5307,N_5220);
nand U6740 (N_6740,N_5017,N_5396);
xnor U6741 (N_6741,N_5699,N_5713);
nor U6742 (N_6742,N_5269,N_5926);
and U6743 (N_6743,N_5726,N_5299);
xor U6744 (N_6744,N_5812,N_5118);
and U6745 (N_6745,N_5127,N_5779);
or U6746 (N_6746,N_5252,N_5269);
or U6747 (N_6747,N_5004,N_5900);
xnor U6748 (N_6748,N_5511,N_5419);
nand U6749 (N_6749,N_5279,N_5917);
or U6750 (N_6750,N_5383,N_5635);
or U6751 (N_6751,N_5520,N_5330);
nor U6752 (N_6752,N_5137,N_5745);
nor U6753 (N_6753,N_5053,N_5022);
nand U6754 (N_6754,N_5772,N_5590);
nand U6755 (N_6755,N_5409,N_5116);
nand U6756 (N_6756,N_5373,N_5198);
xnor U6757 (N_6757,N_5121,N_5682);
or U6758 (N_6758,N_5794,N_5012);
and U6759 (N_6759,N_5892,N_5724);
or U6760 (N_6760,N_5516,N_5494);
nor U6761 (N_6761,N_5365,N_5926);
nor U6762 (N_6762,N_5979,N_5517);
nand U6763 (N_6763,N_5496,N_5508);
nand U6764 (N_6764,N_5005,N_5573);
xnor U6765 (N_6765,N_5425,N_5283);
nand U6766 (N_6766,N_5313,N_5422);
nor U6767 (N_6767,N_5059,N_5208);
nand U6768 (N_6768,N_5113,N_5827);
or U6769 (N_6769,N_5709,N_5505);
or U6770 (N_6770,N_5722,N_5499);
xnor U6771 (N_6771,N_5674,N_5314);
and U6772 (N_6772,N_5755,N_5109);
or U6773 (N_6773,N_5538,N_5440);
or U6774 (N_6774,N_5054,N_5062);
or U6775 (N_6775,N_5558,N_5629);
xor U6776 (N_6776,N_5097,N_5516);
nor U6777 (N_6777,N_5679,N_5934);
nand U6778 (N_6778,N_5071,N_5719);
nor U6779 (N_6779,N_5361,N_5399);
nor U6780 (N_6780,N_5821,N_5921);
or U6781 (N_6781,N_5245,N_5264);
nand U6782 (N_6782,N_5800,N_5412);
and U6783 (N_6783,N_5222,N_5201);
and U6784 (N_6784,N_5696,N_5018);
nand U6785 (N_6785,N_5076,N_5474);
xor U6786 (N_6786,N_5364,N_5368);
xnor U6787 (N_6787,N_5229,N_5156);
or U6788 (N_6788,N_5648,N_5747);
nand U6789 (N_6789,N_5283,N_5276);
nor U6790 (N_6790,N_5666,N_5444);
xnor U6791 (N_6791,N_5628,N_5705);
and U6792 (N_6792,N_5283,N_5439);
nand U6793 (N_6793,N_5982,N_5539);
nor U6794 (N_6794,N_5095,N_5273);
xnor U6795 (N_6795,N_5728,N_5650);
nand U6796 (N_6796,N_5721,N_5931);
nand U6797 (N_6797,N_5628,N_5744);
or U6798 (N_6798,N_5397,N_5423);
xnor U6799 (N_6799,N_5976,N_5174);
or U6800 (N_6800,N_5231,N_5982);
nand U6801 (N_6801,N_5965,N_5120);
or U6802 (N_6802,N_5406,N_5235);
or U6803 (N_6803,N_5613,N_5570);
and U6804 (N_6804,N_5063,N_5873);
or U6805 (N_6805,N_5834,N_5375);
and U6806 (N_6806,N_5287,N_5022);
xor U6807 (N_6807,N_5050,N_5207);
nor U6808 (N_6808,N_5934,N_5935);
xor U6809 (N_6809,N_5009,N_5099);
or U6810 (N_6810,N_5860,N_5602);
or U6811 (N_6811,N_5790,N_5337);
nor U6812 (N_6812,N_5246,N_5717);
xor U6813 (N_6813,N_5636,N_5202);
nand U6814 (N_6814,N_5850,N_5016);
and U6815 (N_6815,N_5415,N_5087);
nor U6816 (N_6816,N_5032,N_5231);
nand U6817 (N_6817,N_5897,N_5681);
nor U6818 (N_6818,N_5581,N_5643);
or U6819 (N_6819,N_5989,N_5196);
or U6820 (N_6820,N_5896,N_5528);
or U6821 (N_6821,N_5194,N_5131);
nor U6822 (N_6822,N_5553,N_5011);
xor U6823 (N_6823,N_5428,N_5633);
nand U6824 (N_6824,N_5289,N_5020);
or U6825 (N_6825,N_5430,N_5306);
or U6826 (N_6826,N_5326,N_5231);
nor U6827 (N_6827,N_5981,N_5875);
or U6828 (N_6828,N_5062,N_5789);
or U6829 (N_6829,N_5510,N_5541);
nand U6830 (N_6830,N_5580,N_5407);
nand U6831 (N_6831,N_5410,N_5698);
or U6832 (N_6832,N_5022,N_5187);
or U6833 (N_6833,N_5441,N_5855);
nor U6834 (N_6834,N_5036,N_5084);
nand U6835 (N_6835,N_5720,N_5881);
xnor U6836 (N_6836,N_5513,N_5581);
nand U6837 (N_6837,N_5789,N_5158);
nand U6838 (N_6838,N_5517,N_5020);
nand U6839 (N_6839,N_5677,N_5974);
nor U6840 (N_6840,N_5918,N_5876);
and U6841 (N_6841,N_5887,N_5174);
or U6842 (N_6842,N_5388,N_5320);
xnor U6843 (N_6843,N_5332,N_5473);
and U6844 (N_6844,N_5894,N_5548);
xor U6845 (N_6845,N_5342,N_5909);
nand U6846 (N_6846,N_5839,N_5058);
and U6847 (N_6847,N_5055,N_5925);
xnor U6848 (N_6848,N_5749,N_5813);
and U6849 (N_6849,N_5896,N_5599);
nand U6850 (N_6850,N_5360,N_5195);
nor U6851 (N_6851,N_5675,N_5718);
xor U6852 (N_6852,N_5540,N_5020);
nor U6853 (N_6853,N_5335,N_5639);
nor U6854 (N_6854,N_5672,N_5653);
nor U6855 (N_6855,N_5118,N_5426);
xnor U6856 (N_6856,N_5938,N_5684);
or U6857 (N_6857,N_5726,N_5884);
nand U6858 (N_6858,N_5199,N_5150);
nor U6859 (N_6859,N_5739,N_5160);
xor U6860 (N_6860,N_5423,N_5336);
or U6861 (N_6861,N_5335,N_5108);
or U6862 (N_6862,N_5087,N_5753);
nor U6863 (N_6863,N_5721,N_5362);
and U6864 (N_6864,N_5274,N_5905);
and U6865 (N_6865,N_5434,N_5072);
xnor U6866 (N_6866,N_5815,N_5198);
xor U6867 (N_6867,N_5585,N_5509);
and U6868 (N_6868,N_5479,N_5610);
nand U6869 (N_6869,N_5095,N_5768);
nor U6870 (N_6870,N_5405,N_5743);
xor U6871 (N_6871,N_5408,N_5777);
nor U6872 (N_6872,N_5394,N_5510);
or U6873 (N_6873,N_5116,N_5085);
or U6874 (N_6874,N_5376,N_5118);
or U6875 (N_6875,N_5051,N_5260);
nor U6876 (N_6876,N_5961,N_5514);
and U6877 (N_6877,N_5728,N_5135);
nand U6878 (N_6878,N_5613,N_5688);
nand U6879 (N_6879,N_5736,N_5213);
xor U6880 (N_6880,N_5346,N_5225);
nand U6881 (N_6881,N_5378,N_5123);
or U6882 (N_6882,N_5518,N_5841);
xnor U6883 (N_6883,N_5147,N_5072);
and U6884 (N_6884,N_5478,N_5048);
xor U6885 (N_6885,N_5232,N_5073);
xor U6886 (N_6886,N_5743,N_5382);
nand U6887 (N_6887,N_5168,N_5368);
nor U6888 (N_6888,N_5196,N_5568);
nand U6889 (N_6889,N_5383,N_5300);
nor U6890 (N_6890,N_5214,N_5661);
and U6891 (N_6891,N_5819,N_5305);
nand U6892 (N_6892,N_5078,N_5451);
and U6893 (N_6893,N_5055,N_5437);
xnor U6894 (N_6894,N_5888,N_5292);
nor U6895 (N_6895,N_5303,N_5014);
xnor U6896 (N_6896,N_5405,N_5589);
xor U6897 (N_6897,N_5959,N_5331);
or U6898 (N_6898,N_5929,N_5281);
and U6899 (N_6899,N_5309,N_5849);
nand U6900 (N_6900,N_5778,N_5709);
xor U6901 (N_6901,N_5563,N_5545);
and U6902 (N_6902,N_5251,N_5888);
nor U6903 (N_6903,N_5278,N_5420);
and U6904 (N_6904,N_5401,N_5569);
nor U6905 (N_6905,N_5204,N_5891);
nor U6906 (N_6906,N_5718,N_5846);
nand U6907 (N_6907,N_5726,N_5034);
xnor U6908 (N_6908,N_5531,N_5213);
nor U6909 (N_6909,N_5916,N_5704);
xor U6910 (N_6910,N_5990,N_5774);
nor U6911 (N_6911,N_5030,N_5683);
or U6912 (N_6912,N_5962,N_5411);
xnor U6913 (N_6913,N_5330,N_5017);
xnor U6914 (N_6914,N_5648,N_5112);
and U6915 (N_6915,N_5794,N_5975);
and U6916 (N_6916,N_5862,N_5584);
and U6917 (N_6917,N_5707,N_5844);
xnor U6918 (N_6918,N_5083,N_5858);
nor U6919 (N_6919,N_5345,N_5836);
nor U6920 (N_6920,N_5289,N_5901);
nor U6921 (N_6921,N_5160,N_5826);
and U6922 (N_6922,N_5670,N_5278);
xor U6923 (N_6923,N_5851,N_5876);
and U6924 (N_6924,N_5061,N_5694);
nor U6925 (N_6925,N_5203,N_5202);
or U6926 (N_6926,N_5388,N_5073);
nor U6927 (N_6927,N_5229,N_5507);
xor U6928 (N_6928,N_5904,N_5993);
nor U6929 (N_6929,N_5879,N_5068);
nand U6930 (N_6930,N_5861,N_5976);
nor U6931 (N_6931,N_5268,N_5283);
or U6932 (N_6932,N_5344,N_5054);
or U6933 (N_6933,N_5417,N_5275);
and U6934 (N_6934,N_5423,N_5539);
or U6935 (N_6935,N_5691,N_5726);
and U6936 (N_6936,N_5244,N_5385);
xor U6937 (N_6937,N_5157,N_5403);
xnor U6938 (N_6938,N_5091,N_5563);
xor U6939 (N_6939,N_5574,N_5460);
or U6940 (N_6940,N_5154,N_5020);
and U6941 (N_6941,N_5958,N_5224);
or U6942 (N_6942,N_5811,N_5579);
nand U6943 (N_6943,N_5309,N_5816);
and U6944 (N_6944,N_5428,N_5256);
and U6945 (N_6945,N_5966,N_5011);
nand U6946 (N_6946,N_5993,N_5180);
xnor U6947 (N_6947,N_5989,N_5239);
nor U6948 (N_6948,N_5700,N_5060);
nand U6949 (N_6949,N_5034,N_5011);
xnor U6950 (N_6950,N_5549,N_5922);
nand U6951 (N_6951,N_5863,N_5112);
and U6952 (N_6952,N_5447,N_5375);
or U6953 (N_6953,N_5775,N_5464);
or U6954 (N_6954,N_5721,N_5602);
nor U6955 (N_6955,N_5745,N_5538);
xnor U6956 (N_6956,N_5853,N_5560);
and U6957 (N_6957,N_5659,N_5707);
nor U6958 (N_6958,N_5835,N_5390);
xor U6959 (N_6959,N_5298,N_5681);
and U6960 (N_6960,N_5191,N_5889);
xnor U6961 (N_6961,N_5489,N_5967);
or U6962 (N_6962,N_5995,N_5014);
or U6963 (N_6963,N_5369,N_5921);
xnor U6964 (N_6964,N_5854,N_5183);
or U6965 (N_6965,N_5565,N_5759);
or U6966 (N_6966,N_5038,N_5668);
and U6967 (N_6967,N_5154,N_5274);
or U6968 (N_6968,N_5962,N_5234);
or U6969 (N_6969,N_5249,N_5415);
or U6970 (N_6970,N_5442,N_5058);
xnor U6971 (N_6971,N_5013,N_5328);
nand U6972 (N_6972,N_5338,N_5819);
xnor U6973 (N_6973,N_5566,N_5191);
nand U6974 (N_6974,N_5014,N_5273);
or U6975 (N_6975,N_5986,N_5905);
nor U6976 (N_6976,N_5361,N_5384);
and U6977 (N_6977,N_5238,N_5710);
nand U6978 (N_6978,N_5464,N_5442);
nor U6979 (N_6979,N_5618,N_5075);
nor U6980 (N_6980,N_5339,N_5881);
and U6981 (N_6981,N_5867,N_5952);
or U6982 (N_6982,N_5129,N_5608);
nor U6983 (N_6983,N_5115,N_5686);
nand U6984 (N_6984,N_5943,N_5761);
and U6985 (N_6985,N_5039,N_5116);
xnor U6986 (N_6986,N_5250,N_5350);
xor U6987 (N_6987,N_5421,N_5490);
xnor U6988 (N_6988,N_5124,N_5879);
nor U6989 (N_6989,N_5952,N_5255);
or U6990 (N_6990,N_5586,N_5557);
and U6991 (N_6991,N_5157,N_5631);
nand U6992 (N_6992,N_5208,N_5178);
nor U6993 (N_6993,N_5801,N_5777);
xor U6994 (N_6994,N_5150,N_5889);
xor U6995 (N_6995,N_5800,N_5198);
xor U6996 (N_6996,N_5731,N_5552);
xnor U6997 (N_6997,N_5532,N_5870);
or U6998 (N_6998,N_5063,N_5489);
xor U6999 (N_6999,N_5872,N_5558);
nor U7000 (N_7000,N_6220,N_6041);
xnor U7001 (N_7001,N_6540,N_6029);
and U7002 (N_7002,N_6557,N_6727);
nor U7003 (N_7003,N_6454,N_6021);
xnor U7004 (N_7004,N_6067,N_6235);
xnor U7005 (N_7005,N_6955,N_6660);
nor U7006 (N_7006,N_6700,N_6891);
nor U7007 (N_7007,N_6569,N_6825);
xnor U7008 (N_7008,N_6225,N_6365);
or U7009 (N_7009,N_6059,N_6732);
nand U7010 (N_7010,N_6736,N_6315);
and U7011 (N_7011,N_6232,N_6508);
and U7012 (N_7012,N_6299,N_6722);
and U7013 (N_7013,N_6723,N_6184);
or U7014 (N_7014,N_6410,N_6885);
and U7015 (N_7015,N_6575,N_6134);
nand U7016 (N_7016,N_6491,N_6471);
or U7017 (N_7017,N_6519,N_6153);
nand U7018 (N_7018,N_6164,N_6149);
or U7019 (N_7019,N_6151,N_6439);
xnor U7020 (N_7020,N_6774,N_6800);
or U7021 (N_7021,N_6999,N_6820);
nand U7022 (N_7022,N_6387,N_6193);
and U7023 (N_7023,N_6422,N_6648);
xor U7024 (N_7024,N_6452,N_6168);
nor U7025 (N_7025,N_6547,N_6453);
and U7026 (N_7026,N_6297,N_6495);
xnor U7027 (N_7027,N_6699,N_6518);
or U7028 (N_7028,N_6636,N_6864);
and U7029 (N_7029,N_6412,N_6009);
or U7030 (N_7030,N_6393,N_6243);
xor U7031 (N_7031,N_6620,N_6244);
nand U7032 (N_7032,N_6320,N_6106);
xnor U7033 (N_7033,N_6857,N_6119);
or U7034 (N_7034,N_6994,N_6192);
nand U7035 (N_7035,N_6592,N_6687);
nor U7036 (N_7036,N_6381,N_6094);
xor U7037 (N_7037,N_6643,N_6350);
xor U7038 (N_7038,N_6429,N_6444);
nor U7039 (N_7039,N_6406,N_6582);
nor U7040 (N_7040,N_6023,N_6658);
xor U7041 (N_7041,N_6497,N_6222);
xor U7042 (N_7042,N_6421,N_6216);
nand U7043 (N_7043,N_6652,N_6664);
or U7044 (N_7044,N_6534,N_6420);
or U7045 (N_7045,N_6418,N_6672);
xor U7046 (N_7046,N_6487,N_6738);
xnor U7047 (N_7047,N_6536,N_6383);
and U7048 (N_7048,N_6959,N_6115);
nand U7049 (N_7049,N_6758,N_6018);
or U7050 (N_7050,N_6697,N_6177);
nor U7051 (N_7051,N_6572,N_6596);
nor U7052 (N_7052,N_6267,N_6550);
or U7053 (N_7053,N_6924,N_6032);
xnor U7054 (N_7054,N_6897,N_6101);
nand U7055 (N_7055,N_6522,N_6366);
nor U7056 (N_7056,N_6436,N_6790);
nand U7057 (N_7057,N_6348,N_6413);
xor U7058 (N_7058,N_6679,N_6868);
xnor U7059 (N_7059,N_6795,N_6245);
or U7060 (N_7060,N_6754,N_6208);
or U7061 (N_7061,N_6000,N_6206);
nand U7062 (N_7062,N_6887,N_6064);
nand U7063 (N_7063,N_6476,N_6185);
nand U7064 (N_7064,N_6593,N_6740);
nor U7065 (N_7065,N_6603,N_6640);
nand U7066 (N_7066,N_6947,N_6678);
nand U7067 (N_7067,N_6416,N_6645);
and U7068 (N_7068,N_6969,N_6797);
or U7069 (N_7069,N_6538,N_6323);
nor U7070 (N_7070,N_6580,N_6874);
nand U7071 (N_7071,N_6762,N_6621);
or U7072 (N_7072,N_6928,N_6120);
and U7073 (N_7073,N_6945,N_6667);
nor U7074 (N_7074,N_6057,N_6772);
nand U7075 (N_7075,N_6895,N_6015);
nand U7076 (N_7076,N_6458,N_6583);
and U7077 (N_7077,N_6711,N_6319);
and U7078 (N_7078,N_6211,N_6574);
xnor U7079 (N_7079,N_6637,N_6089);
or U7080 (N_7080,N_6663,N_6005);
and U7081 (N_7081,N_6174,N_6460);
nor U7082 (N_7082,N_6619,N_6338);
nand U7083 (N_7083,N_6719,N_6730);
nand U7084 (N_7084,N_6869,N_6777);
xor U7085 (N_7085,N_6257,N_6317);
xor U7086 (N_7086,N_6769,N_6759);
nand U7087 (N_7087,N_6913,N_6889);
nand U7088 (N_7088,N_6814,N_6570);
nand U7089 (N_7089,N_6539,N_6258);
or U7090 (N_7090,N_6720,N_6828);
and U7091 (N_7091,N_6349,N_6241);
xnor U7092 (N_7092,N_6311,N_6405);
nand U7093 (N_7093,N_6266,N_6563);
nor U7094 (N_7094,N_6052,N_6294);
or U7095 (N_7095,N_6501,N_6705);
and U7096 (N_7096,N_6129,N_6346);
xor U7097 (N_7097,N_6635,N_6038);
xor U7098 (N_7098,N_6933,N_6447);
and U7099 (N_7099,N_6143,N_6749);
nor U7100 (N_7100,N_6974,N_6287);
nor U7101 (N_7101,N_6489,N_6028);
nor U7102 (N_7102,N_6624,N_6859);
nand U7103 (N_7103,N_6541,N_6992);
nand U7104 (N_7104,N_6404,N_6104);
or U7105 (N_7105,N_6710,N_6062);
nand U7106 (N_7106,N_6839,N_6303);
or U7107 (N_7107,N_6816,N_6829);
or U7108 (N_7108,N_6466,N_6163);
or U7109 (N_7109,N_6837,N_6930);
xor U7110 (N_7110,N_6097,N_6778);
nand U7111 (N_7111,N_6801,N_6763);
or U7112 (N_7112,N_6110,N_6233);
xnor U7113 (N_7113,N_6262,N_6647);
and U7114 (N_7114,N_6701,N_6111);
xor U7115 (N_7115,N_6074,N_6884);
xor U7116 (N_7116,N_6483,N_6506);
nor U7117 (N_7117,N_6627,N_6296);
xor U7118 (N_7118,N_6558,N_6988);
nand U7119 (N_7119,N_6069,N_6157);
or U7120 (N_7120,N_6911,N_6438);
and U7121 (N_7121,N_6917,N_6448);
or U7122 (N_7122,N_6920,N_6165);
xnor U7123 (N_7123,N_6813,N_6626);
xor U7124 (N_7124,N_6354,N_6597);
and U7125 (N_7125,N_6983,N_6330);
and U7126 (N_7126,N_6646,N_6161);
and U7127 (N_7127,N_6671,N_6760);
nor U7128 (N_7128,N_6113,N_6733);
xor U7129 (N_7129,N_6980,N_6461);
nand U7130 (N_7130,N_6352,N_6811);
nor U7131 (N_7131,N_6644,N_6782);
and U7132 (N_7132,N_6159,N_6326);
xor U7133 (N_7133,N_6043,N_6934);
and U7134 (N_7134,N_6083,N_6707);
nor U7135 (N_7135,N_6601,N_6309);
xor U7136 (N_7136,N_6831,N_6375);
nand U7137 (N_7137,N_6382,N_6526);
xor U7138 (N_7138,N_6669,N_6271);
and U7139 (N_7139,N_6914,N_6929);
and U7140 (N_7140,N_6351,N_6888);
nand U7141 (N_7141,N_6553,N_6567);
nand U7142 (N_7142,N_6953,N_6316);
or U7143 (N_7143,N_6552,N_6450);
or U7144 (N_7144,N_6250,N_6084);
and U7145 (N_7145,N_6688,N_6171);
or U7146 (N_7146,N_6230,N_6610);
xor U7147 (N_7147,N_6044,N_6103);
nand U7148 (N_7148,N_6036,N_6715);
and U7149 (N_7149,N_6449,N_6657);
or U7150 (N_7150,N_6949,N_6872);
xor U7151 (N_7151,N_6086,N_6815);
nand U7152 (N_7152,N_6773,N_6982);
or U7153 (N_7153,N_6984,N_6692);
or U7154 (N_7154,N_6053,N_6173);
nor U7155 (N_7155,N_6154,N_6823);
or U7156 (N_7156,N_6817,N_6729);
xnor U7157 (N_7157,N_6842,N_6144);
xnor U7158 (N_7158,N_6175,N_6473);
xnor U7159 (N_7159,N_6957,N_6785);
or U7160 (N_7160,N_6904,N_6373);
xnor U7161 (N_7161,N_6581,N_6131);
or U7162 (N_7162,N_6200,N_6863);
nand U7163 (N_7163,N_6750,N_6076);
nor U7164 (N_7164,N_6105,N_6408);
or U7165 (N_7165,N_6457,N_6465);
and U7166 (N_7166,N_6588,N_6475);
or U7167 (N_7167,N_6283,N_6288);
nor U7168 (N_7168,N_6630,N_6302);
and U7169 (N_7169,N_6456,N_6555);
xnor U7170 (N_7170,N_6551,N_6632);
or U7171 (N_7171,N_6851,N_6724);
nand U7172 (N_7172,N_6870,N_6493);
nor U7173 (N_7173,N_6007,N_6136);
xor U7174 (N_7174,N_6910,N_6251);
nand U7175 (N_7175,N_6589,N_6617);
or U7176 (N_7176,N_6606,N_6977);
and U7177 (N_7177,N_6198,N_6060);
nor U7178 (N_7178,N_6395,N_6231);
or U7179 (N_7179,N_6649,N_6591);
and U7180 (N_7180,N_6178,N_6135);
nand U7181 (N_7181,N_6298,N_6203);
or U7182 (N_7182,N_6484,N_6363);
nor U7183 (N_7183,N_6826,N_6873);
and U7184 (N_7184,N_6042,N_6860);
or U7185 (N_7185,N_6432,N_6242);
nor U7186 (N_7186,N_6818,N_6639);
nor U7187 (N_7187,N_6162,N_6892);
nor U7188 (N_7188,N_6331,N_6051);
xnor U7189 (N_7189,N_6045,N_6409);
and U7190 (N_7190,N_6995,N_6686);
nor U7191 (N_7191,N_6150,N_6716);
xor U7192 (N_7192,N_6335,N_6158);
nand U7193 (N_7193,N_6215,N_6407);
nand U7194 (N_7194,N_6342,N_6071);
nand U7195 (N_7195,N_6771,N_6921);
and U7196 (N_7196,N_6279,N_6682);
or U7197 (N_7197,N_6332,N_6962);
xor U7198 (N_7198,N_6830,N_6399);
and U7199 (N_7199,N_6204,N_6369);
nor U7200 (N_7200,N_6708,N_6088);
nor U7201 (N_7201,N_6940,N_6605);
or U7202 (N_7202,N_6166,N_6846);
and U7203 (N_7203,N_6295,N_6238);
and U7204 (N_7204,N_6445,N_6952);
nand U7205 (N_7205,N_6079,N_6040);
xnor U7206 (N_7206,N_6077,N_6525);
nand U7207 (N_7207,N_6879,N_6145);
and U7208 (N_7208,N_6004,N_6998);
and U7209 (N_7209,N_6673,N_6430);
and U7210 (N_7210,N_6991,N_6584);
nor U7211 (N_7211,N_6030,N_6061);
nor U7212 (N_7212,N_6305,N_6919);
xor U7213 (N_7213,N_6195,N_6946);
and U7214 (N_7214,N_6753,N_6306);
nand U7215 (N_7215,N_6625,N_6341);
xnor U7216 (N_7216,N_6236,N_6100);
and U7217 (N_7217,N_6254,N_6390);
or U7218 (N_7218,N_6132,N_6609);
or U7219 (N_7219,N_6549,N_6034);
and U7220 (N_7220,N_6344,N_6020);
or U7221 (N_7221,N_6081,N_6396);
and U7222 (N_7222,N_6065,N_6883);
nand U7223 (N_7223,N_6560,N_6993);
nand U7224 (N_7224,N_6237,N_6668);
or U7225 (N_7225,N_6424,N_6109);
xor U7226 (N_7226,N_6260,N_6310);
and U7227 (N_7227,N_6082,N_6691);
nor U7228 (N_7228,N_6116,N_6922);
nor U7229 (N_7229,N_6702,N_6093);
nand U7230 (N_7230,N_6099,N_6265);
or U7231 (N_7231,N_6505,N_6985);
nand U7232 (N_7232,N_6474,N_6056);
nor U7233 (N_7233,N_6598,N_6415);
xor U7234 (N_7234,N_6741,N_6339);
nor U7235 (N_7235,N_6511,N_6284);
or U7236 (N_7236,N_6803,N_6936);
nor U7237 (N_7237,N_6514,N_6205);
nand U7238 (N_7238,N_6507,N_6973);
nor U7239 (N_7239,N_6717,N_6943);
nor U7240 (N_7240,N_6942,N_6285);
or U7241 (N_7241,N_6893,N_6345);
xnor U7242 (N_7242,N_6167,N_6950);
and U7243 (N_7243,N_6123,N_6014);
nand U7244 (N_7244,N_6440,N_6472);
nand U7245 (N_7245,N_6270,N_6967);
and U7246 (N_7246,N_6228,N_6901);
and U7247 (N_7247,N_6768,N_6427);
nor U7248 (N_7248,N_6935,N_6796);
xnor U7249 (N_7249,N_6480,N_6389);
and U7250 (N_7250,N_6329,N_6488);
xnor U7251 (N_7251,N_6358,N_6926);
nor U7252 (N_7252,N_6090,N_6559);
and U7253 (N_7253,N_6989,N_6651);
xnor U7254 (N_7254,N_6812,N_6026);
nand U7255 (N_7255,N_6903,N_6356);
or U7256 (N_7256,N_6479,N_6118);
or U7257 (N_7257,N_6531,N_6304);
nand U7258 (N_7258,N_6862,N_6226);
xor U7259 (N_7259,N_6755,N_6912);
or U7260 (N_7260,N_6391,N_6397);
nand U7261 (N_7261,N_6655,N_6209);
nor U7262 (N_7262,N_6152,N_6709);
or U7263 (N_7263,N_6960,N_6607);
and U7264 (N_7264,N_6054,N_6462);
nor U7265 (N_7265,N_6804,N_6737);
and U7266 (N_7266,N_6680,N_6576);
nand U7267 (N_7267,N_6325,N_6114);
xor U7268 (N_7268,N_6779,N_6140);
xor U7269 (N_7269,N_6336,N_6742);
nor U7270 (N_7270,N_6739,N_6963);
or U7271 (N_7271,N_6047,N_6761);
nor U7272 (N_7272,N_6791,N_6923);
or U7273 (N_7273,N_6512,N_6401);
and U7274 (N_7274,N_6517,N_6698);
nor U7275 (N_7275,N_6971,N_6039);
nand U7276 (N_7276,N_6898,N_6292);
nand U7277 (N_7277,N_6684,N_6757);
nand U7278 (N_7278,N_6359,N_6641);
nand U7279 (N_7279,N_6808,N_6308);
nand U7280 (N_7280,N_6524,N_6661);
nor U7281 (N_7281,N_6180,N_6470);
xnor U7282 (N_7282,N_6642,N_6681);
or U7283 (N_7283,N_6835,N_6091);
and U7284 (N_7284,N_6234,N_6377);
xnor U7285 (N_7285,N_6075,N_6728);
nor U7286 (N_7286,N_6033,N_6246);
or U7287 (N_7287,N_6908,N_6824);
and U7288 (N_7288,N_6419,N_6871);
xnor U7289 (N_7289,N_6931,N_6148);
nand U7290 (N_7290,N_6916,N_6016);
nor U7291 (N_7291,N_6735,N_6533);
nor U7292 (N_7292,N_6256,N_6756);
nor U7293 (N_7293,N_6746,N_6146);
xnor U7294 (N_7294,N_6822,N_6585);
nor U7295 (N_7295,N_6918,N_6496);
nand U7296 (N_7296,N_6503,N_6314);
xnor U7297 (N_7297,N_6527,N_6747);
or U7298 (N_7298,N_6063,N_6293);
nand U7299 (N_7299,N_6788,N_6941);
nor U7300 (N_7300,N_6455,N_6035);
or U7301 (N_7301,N_6147,N_6564);
or U7302 (N_7302,N_6194,N_6855);
nand U7303 (N_7303,N_6227,N_6012);
nand U7304 (N_7304,N_6944,N_6532);
and U7305 (N_7305,N_6008,N_6400);
or U7306 (N_7306,N_6670,N_6578);
or U7307 (N_7307,N_6137,N_6384);
nand U7308 (N_7308,N_6614,N_6770);
xnor U7309 (N_7309,N_6628,N_6544);
and U7310 (N_7310,N_6378,N_6181);
or U7311 (N_7311,N_6282,N_6277);
and U7312 (N_7312,N_6169,N_6938);
xor U7313 (N_7313,N_6223,N_6858);
xor U7314 (N_7314,N_6834,N_6182);
nand U7315 (N_7315,N_6442,N_6662);
nor U7316 (N_7316,N_6612,N_6490);
or U7317 (N_7317,N_6392,N_6676);
or U7318 (N_7318,N_6275,N_6434);
xor U7319 (N_7319,N_6433,N_6172);
nand U7320 (N_7320,N_6852,N_6838);
nor U7321 (N_7321,N_6902,N_6398);
nor U7322 (N_7322,N_6080,N_6191);
or U7323 (N_7323,N_6713,N_6229);
xnor U7324 (N_7324,N_6725,N_6677);
and U7325 (N_7325,N_6896,N_6721);
nor U7326 (N_7326,N_6968,N_6685);
nor U7327 (N_7327,N_6556,N_6502);
nand U7328 (N_7328,N_6899,N_6031);
nand U7329 (N_7329,N_6900,N_6765);
nand U7330 (N_7330,N_6854,N_6312);
nor U7331 (N_7331,N_6805,N_6190);
xnor U7332 (N_7332,N_6613,N_6714);
nor U7333 (N_7333,N_6767,N_6545);
or U7334 (N_7334,N_6376,N_6878);
nand U7335 (N_7335,N_6978,N_6849);
xor U7336 (N_7336,N_6446,N_6122);
xnor U7337 (N_7337,N_6876,N_6217);
and U7338 (N_7338,N_6752,N_6554);
and U7339 (N_7339,N_6261,N_6125);
xnor U7340 (N_7340,N_6504,N_6964);
xnor U7341 (N_7341,N_6718,N_6482);
or U7342 (N_7342,N_6590,N_6499);
xor U7343 (N_7343,N_6290,N_6050);
nor U7344 (N_7344,N_6783,N_6510);
xor U7345 (N_7345,N_6515,N_6521);
nor U7346 (N_7346,N_6078,N_6961);
and U7347 (N_7347,N_6469,N_6529);
or U7348 (N_7348,N_6986,N_6599);
nand U7349 (N_7349,N_6112,N_6500);
nand U7350 (N_7350,N_6520,N_6807);
nor U7351 (N_7351,N_6478,N_6970);
or U7352 (N_7352,N_6107,N_6731);
xor U7353 (N_7353,N_6255,N_6594);
or U7354 (N_7354,N_6058,N_6095);
and U7355 (N_7355,N_6987,N_6353);
and U7356 (N_7356,N_6695,N_6139);
xnor U7357 (N_7357,N_6611,N_6321);
xor U7358 (N_7358,N_6799,N_6070);
xnor U7359 (N_7359,N_6179,N_6881);
nand U7360 (N_7360,N_6543,N_6046);
nor U7361 (N_7361,N_6748,N_6128);
nand U7362 (N_7362,N_6650,N_6343);
nand U7363 (N_7363,N_6806,N_6201);
nand U7364 (N_7364,N_6049,N_6126);
and U7365 (N_7365,N_6017,N_6633);
and U7366 (N_7366,N_6653,N_6367);
nor U7367 (N_7367,N_6186,N_6827);
or U7368 (N_7368,N_6966,N_6385);
xnor U7369 (N_7369,N_6787,N_6467);
nor U7370 (N_7370,N_6027,N_6734);
xor U7371 (N_7371,N_6498,N_6568);
nor U7372 (N_7372,N_6751,N_6333);
xor U7373 (N_7373,N_6357,N_6975);
nor U7374 (N_7374,N_6587,N_6997);
or U7375 (N_7375,N_6802,N_6096);
and U7376 (N_7376,N_6214,N_6792);
nand U7377 (N_7377,N_6219,N_6890);
nor U7378 (N_7378,N_6882,N_6481);
nor U7379 (N_7379,N_6210,N_6766);
or U7380 (N_7380,N_6608,N_6334);
and U7381 (N_7381,N_6127,N_6011);
and U7382 (N_7382,N_6509,N_6066);
or U7383 (N_7383,N_6130,N_6615);
xor U7384 (N_7384,N_6459,N_6108);
or U7385 (N_7385,N_6623,N_6068);
nor U7386 (N_7386,N_6542,N_6425);
or U7387 (N_7387,N_6280,N_6102);
nor U7388 (N_7388,N_6877,N_6979);
or U7389 (N_7389,N_6318,N_6809);
xor U7390 (N_7390,N_6417,N_6745);
and U7391 (N_7391,N_6704,N_6301);
nor U7392 (N_7392,N_6798,N_6530);
nor U7393 (N_7393,N_6784,N_6665);
xnor U7394 (N_7394,N_6259,N_6431);
nand U7395 (N_7395,N_6240,N_6024);
nor U7396 (N_7396,N_6786,N_6337);
xor U7397 (N_7397,N_6965,N_6142);
xnor U7398 (N_7398,N_6264,N_6932);
xor U7399 (N_7399,N_6278,N_6138);
xor U7400 (N_7400,N_6291,N_6819);
xnor U7401 (N_7401,N_6616,N_6866);
and U7402 (N_7402,N_6022,N_6213);
or U7403 (N_7403,N_6477,N_6402);
nor U7404 (N_7404,N_6845,N_6037);
nand U7405 (N_7405,N_6492,N_6972);
nor U7406 (N_7406,N_6380,N_6388);
and U7407 (N_7407,N_6327,N_6516);
nor U7408 (N_7408,N_6300,N_6844);
xnor U7409 (N_7409,N_6703,N_6072);
nand U7410 (N_7410,N_6656,N_6781);
nand U7411 (N_7411,N_6428,N_6252);
or U7412 (N_7412,N_6124,N_6437);
nand U7413 (N_7413,N_6372,N_6622);
nor U7414 (N_7414,N_6602,N_6764);
and U7415 (N_7415,N_6189,N_6836);
nand U7416 (N_7416,N_6573,N_6571);
or U7417 (N_7417,N_6239,N_6631);
and U7418 (N_7418,N_6861,N_6843);
nor U7419 (N_7419,N_6019,N_6322);
nor U7420 (N_7420,N_6324,N_6411);
nor U7421 (N_7421,N_6810,N_6435);
or U7422 (N_7422,N_6155,N_6562);
nor U7423 (N_7423,N_6187,N_6535);
and U7424 (N_7424,N_6451,N_6666);
nor U7425 (N_7425,N_6013,N_6875);
nor U7426 (N_7426,N_6586,N_6025);
nand U7427 (N_7427,N_6659,N_6976);
and U7428 (N_7428,N_6954,N_6276);
xnor U7429 (N_7429,N_6133,N_6561);
and U7430 (N_7430,N_6577,N_6548);
or U7431 (N_7431,N_6360,N_6832);
xor U7432 (N_7432,N_6907,N_6618);
or U7433 (N_7433,N_6909,N_6990);
or U7434 (N_7434,N_6464,N_6156);
or U7435 (N_7435,N_6712,N_6629);
xor U7436 (N_7436,N_6207,N_6833);
xor U7437 (N_7437,N_6981,N_6347);
xor U7438 (N_7438,N_6566,N_6821);
and U7439 (N_7439,N_6002,N_6414);
and U7440 (N_7440,N_6307,N_6361);
or U7441 (N_7441,N_6386,N_6170);
nor U7442 (N_7442,N_6513,N_6092);
or U7443 (N_7443,N_6370,N_6654);
or U7444 (N_7444,N_6689,N_6674);
nor U7445 (N_7445,N_6379,N_6055);
nor U7446 (N_7446,N_6218,N_6188);
and U7447 (N_7447,N_6604,N_6371);
nand U7448 (N_7448,N_6865,N_6906);
nor U7449 (N_7449,N_6085,N_6794);
or U7450 (N_7450,N_6726,N_6867);
or U7451 (N_7451,N_6634,N_6263);
nor U7452 (N_7452,N_6776,N_6696);
nor U7453 (N_7453,N_6197,N_6523);
or U7454 (N_7454,N_6048,N_6249);
nand U7455 (N_7455,N_6247,N_6394);
xnor U7456 (N_7456,N_6253,N_6956);
nand U7457 (N_7457,N_6693,N_6328);
nor U7458 (N_7458,N_6364,N_6925);
nor U7459 (N_7459,N_6468,N_6403);
nand U7460 (N_7460,N_6951,N_6362);
xor U7461 (N_7461,N_6098,N_6274);
and U7462 (N_7462,N_6486,N_6905);
xor U7463 (N_7463,N_6780,N_6268);
nand U7464 (N_7464,N_6638,N_6537);
nand U7465 (N_7465,N_6579,N_6340);
and U7466 (N_7466,N_6775,N_6528);
xor U7467 (N_7467,N_6937,N_6600);
nand U7468 (N_7468,N_6939,N_6199);
xnor U7469 (N_7469,N_6886,N_6847);
or U7470 (N_7470,N_6840,N_6286);
and U7471 (N_7471,N_6224,N_6423);
xnor U7472 (N_7472,N_6281,N_6176);
and U7473 (N_7473,N_6690,N_6141);
nand U7474 (N_7474,N_6958,N_6073);
xor U7475 (N_7475,N_6196,N_6272);
and U7476 (N_7476,N_6248,N_6565);
or U7477 (N_7477,N_6001,N_6744);
nor U7478 (N_7478,N_6441,N_6374);
xnor U7479 (N_7479,N_6269,N_6212);
nand U7480 (N_7480,N_6183,N_6675);
nor U7481 (N_7481,N_6485,N_6494);
nor U7482 (N_7482,N_6443,N_6121);
and U7483 (N_7483,N_6202,N_6880);
nand U7484 (N_7484,N_6743,N_6853);
and U7485 (N_7485,N_6221,N_6006);
nor U7486 (N_7486,N_6694,N_6426);
nor U7487 (N_7487,N_6355,N_6848);
and U7488 (N_7488,N_6273,N_6117);
or U7489 (N_7489,N_6789,N_6087);
xor U7490 (N_7490,N_6856,N_6010);
nand U7491 (N_7491,N_6683,N_6915);
xnor U7492 (N_7492,N_6289,N_6793);
xor U7493 (N_7493,N_6160,N_6463);
nor U7494 (N_7494,N_6996,N_6850);
or U7495 (N_7495,N_6706,N_6368);
and U7496 (N_7496,N_6003,N_6927);
nand U7497 (N_7497,N_6948,N_6841);
xnor U7498 (N_7498,N_6313,N_6894);
nor U7499 (N_7499,N_6595,N_6546);
or U7500 (N_7500,N_6148,N_6528);
nand U7501 (N_7501,N_6537,N_6104);
nand U7502 (N_7502,N_6594,N_6761);
nand U7503 (N_7503,N_6036,N_6280);
and U7504 (N_7504,N_6930,N_6800);
and U7505 (N_7505,N_6236,N_6170);
xnor U7506 (N_7506,N_6904,N_6297);
nor U7507 (N_7507,N_6806,N_6428);
and U7508 (N_7508,N_6206,N_6330);
or U7509 (N_7509,N_6820,N_6139);
nand U7510 (N_7510,N_6065,N_6436);
xnor U7511 (N_7511,N_6293,N_6279);
xor U7512 (N_7512,N_6034,N_6422);
nand U7513 (N_7513,N_6743,N_6136);
nand U7514 (N_7514,N_6375,N_6189);
or U7515 (N_7515,N_6525,N_6296);
and U7516 (N_7516,N_6534,N_6067);
or U7517 (N_7517,N_6055,N_6752);
and U7518 (N_7518,N_6172,N_6942);
and U7519 (N_7519,N_6556,N_6816);
or U7520 (N_7520,N_6524,N_6437);
or U7521 (N_7521,N_6427,N_6497);
nor U7522 (N_7522,N_6312,N_6765);
and U7523 (N_7523,N_6264,N_6221);
nor U7524 (N_7524,N_6715,N_6954);
nand U7525 (N_7525,N_6540,N_6207);
nor U7526 (N_7526,N_6079,N_6850);
xnor U7527 (N_7527,N_6335,N_6860);
nor U7528 (N_7528,N_6320,N_6928);
or U7529 (N_7529,N_6309,N_6514);
nand U7530 (N_7530,N_6535,N_6126);
and U7531 (N_7531,N_6221,N_6064);
nand U7532 (N_7532,N_6461,N_6996);
or U7533 (N_7533,N_6096,N_6930);
or U7534 (N_7534,N_6429,N_6748);
or U7535 (N_7535,N_6258,N_6982);
xor U7536 (N_7536,N_6965,N_6637);
or U7537 (N_7537,N_6479,N_6693);
or U7538 (N_7538,N_6862,N_6075);
or U7539 (N_7539,N_6093,N_6695);
nand U7540 (N_7540,N_6368,N_6623);
or U7541 (N_7541,N_6964,N_6450);
or U7542 (N_7542,N_6377,N_6085);
or U7543 (N_7543,N_6729,N_6676);
nor U7544 (N_7544,N_6122,N_6598);
or U7545 (N_7545,N_6558,N_6798);
nand U7546 (N_7546,N_6968,N_6669);
nor U7547 (N_7547,N_6423,N_6613);
or U7548 (N_7548,N_6241,N_6713);
xnor U7549 (N_7549,N_6303,N_6658);
and U7550 (N_7550,N_6573,N_6676);
and U7551 (N_7551,N_6996,N_6818);
or U7552 (N_7552,N_6174,N_6955);
or U7553 (N_7553,N_6379,N_6664);
and U7554 (N_7554,N_6182,N_6451);
nand U7555 (N_7555,N_6051,N_6413);
and U7556 (N_7556,N_6694,N_6117);
nand U7557 (N_7557,N_6324,N_6875);
nor U7558 (N_7558,N_6143,N_6064);
nor U7559 (N_7559,N_6220,N_6326);
xnor U7560 (N_7560,N_6818,N_6082);
and U7561 (N_7561,N_6254,N_6628);
and U7562 (N_7562,N_6975,N_6114);
nor U7563 (N_7563,N_6369,N_6349);
or U7564 (N_7564,N_6108,N_6009);
nand U7565 (N_7565,N_6655,N_6067);
and U7566 (N_7566,N_6502,N_6212);
xnor U7567 (N_7567,N_6153,N_6025);
or U7568 (N_7568,N_6969,N_6626);
nor U7569 (N_7569,N_6740,N_6023);
and U7570 (N_7570,N_6482,N_6043);
nand U7571 (N_7571,N_6861,N_6190);
nand U7572 (N_7572,N_6139,N_6271);
and U7573 (N_7573,N_6683,N_6157);
or U7574 (N_7574,N_6530,N_6549);
and U7575 (N_7575,N_6616,N_6532);
xor U7576 (N_7576,N_6325,N_6290);
or U7577 (N_7577,N_6699,N_6478);
and U7578 (N_7578,N_6640,N_6327);
and U7579 (N_7579,N_6100,N_6782);
or U7580 (N_7580,N_6630,N_6328);
xor U7581 (N_7581,N_6294,N_6613);
xor U7582 (N_7582,N_6167,N_6544);
and U7583 (N_7583,N_6312,N_6910);
nand U7584 (N_7584,N_6928,N_6347);
nor U7585 (N_7585,N_6372,N_6117);
xor U7586 (N_7586,N_6475,N_6780);
and U7587 (N_7587,N_6405,N_6981);
and U7588 (N_7588,N_6121,N_6843);
xor U7589 (N_7589,N_6893,N_6776);
and U7590 (N_7590,N_6364,N_6985);
nand U7591 (N_7591,N_6649,N_6979);
or U7592 (N_7592,N_6331,N_6435);
and U7593 (N_7593,N_6969,N_6589);
and U7594 (N_7594,N_6908,N_6186);
nand U7595 (N_7595,N_6130,N_6542);
nand U7596 (N_7596,N_6424,N_6135);
xor U7597 (N_7597,N_6168,N_6528);
xnor U7598 (N_7598,N_6830,N_6527);
xnor U7599 (N_7599,N_6849,N_6065);
xnor U7600 (N_7600,N_6704,N_6694);
nor U7601 (N_7601,N_6485,N_6536);
or U7602 (N_7602,N_6860,N_6655);
or U7603 (N_7603,N_6117,N_6637);
nor U7604 (N_7604,N_6091,N_6585);
or U7605 (N_7605,N_6267,N_6888);
nor U7606 (N_7606,N_6217,N_6849);
or U7607 (N_7607,N_6326,N_6059);
nand U7608 (N_7608,N_6921,N_6946);
nor U7609 (N_7609,N_6396,N_6960);
and U7610 (N_7610,N_6711,N_6971);
and U7611 (N_7611,N_6042,N_6288);
and U7612 (N_7612,N_6401,N_6004);
or U7613 (N_7613,N_6327,N_6711);
nand U7614 (N_7614,N_6015,N_6399);
and U7615 (N_7615,N_6325,N_6909);
nor U7616 (N_7616,N_6354,N_6412);
nor U7617 (N_7617,N_6069,N_6530);
nor U7618 (N_7618,N_6845,N_6461);
and U7619 (N_7619,N_6319,N_6334);
nor U7620 (N_7620,N_6865,N_6436);
or U7621 (N_7621,N_6204,N_6993);
and U7622 (N_7622,N_6615,N_6355);
nand U7623 (N_7623,N_6693,N_6175);
nor U7624 (N_7624,N_6467,N_6852);
nand U7625 (N_7625,N_6682,N_6275);
nand U7626 (N_7626,N_6929,N_6865);
nor U7627 (N_7627,N_6835,N_6743);
and U7628 (N_7628,N_6876,N_6634);
and U7629 (N_7629,N_6887,N_6055);
and U7630 (N_7630,N_6022,N_6988);
and U7631 (N_7631,N_6879,N_6730);
nand U7632 (N_7632,N_6062,N_6358);
nor U7633 (N_7633,N_6959,N_6954);
or U7634 (N_7634,N_6928,N_6646);
or U7635 (N_7635,N_6146,N_6728);
nand U7636 (N_7636,N_6552,N_6838);
nor U7637 (N_7637,N_6276,N_6620);
and U7638 (N_7638,N_6542,N_6988);
or U7639 (N_7639,N_6157,N_6335);
nand U7640 (N_7640,N_6618,N_6350);
nand U7641 (N_7641,N_6469,N_6356);
xor U7642 (N_7642,N_6750,N_6133);
nand U7643 (N_7643,N_6077,N_6749);
xnor U7644 (N_7644,N_6535,N_6713);
or U7645 (N_7645,N_6561,N_6899);
xor U7646 (N_7646,N_6344,N_6067);
xor U7647 (N_7647,N_6470,N_6780);
nor U7648 (N_7648,N_6430,N_6277);
nor U7649 (N_7649,N_6514,N_6339);
nor U7650 (N_7650,N_6620,N_6313);
and U7651 (N_7651,N_6816,N_6871);
and U7652 (N_7652,N_6657,N_6417);
xnor U7653 (N_7653,N_6554,N_6193);
and U7654 (N_7654,N_6326,N_6600);
and U7655 (N_7655,N_6154,N_6704);
and U7656 (N_7656,N_6880,N_6566);
nand U7657 (N_7657,N_6017,N_6010);
or U7658 (N_7658,N_6294,N_6185);
nand U7659 (N_7659,N_6649,N_6837);
and U7660 (N_7660,N_6107,N_6828);
xnor U7661 (N_7661,N_6705,N_6920);
and U7662 (N_7662,N_6642,N_6196);
xor U7663 (N_7663,N_6667,N_6118);
xor U7664 (N_7664,N_6779,N_6889);
or U7665 (N_7665,N_6277,N_6372);
xor U7666 (N_7666,N_6326,N_6175);
nand U7667 (N_7667,N_6945,N_6747);
or U7668 (N_7668,N_6231,N_6232);
or U7669 (N_7669,N_6330,N_6977);
or U7670 (N_7670,N_6694,N_6233);
nand U7671 (N_7671,N_6594,N_6035);
xor U7672 (N_7672,N_6517,N_6283);
or U7673 (N_7673,N_6080,N_6043);
and U7674 (N_7674,N_6134,N_6147);
and U7675 (N_7675,N_6848,N_6171);
xnor U7676 (N_7676,N_6368,N_6852);
nor U7677 (N_7677,N_6120,N_6165);
and U7678 (N_7678,N_6740,N_6783);
xor U7679 (N_7679,N_6768,N_6566);
nand U7680 (N_7680,N_6477,N_6938);
or U7681 (N_7681,N_6712,N_6877);
nor U7682 (N_7682,N_6666,N_6039);
nand U7683 (N_7683,N_6738,N_6096);
or U7684 (N_7684,N_6299,N_6209);
nor U7685 (N_7685,N_6498,N_6094);
nor U7686 (N_7686,N_6763,N_6280);
xor U7687 (N_7687,N_6664,N_6781);
and U7688 (N_7688,N_6588,N_6811);
and U7689 (N_7689,N_6536,N_6542);
nand U7690 (N_7690,N_6080,N_6916);
or U7691 (N_7691,N_6620,N_6330);
and U7692 (N_7692,N_6258,N_6996);
and U7693 (N_7693,N_6872,N_6624);
and U7694 (N_7694,N_6195,N_6102);
nand U7695 (N_7695,N_6684,N_6106);
and U7696 (N_7696,N_6056,N_6639);
or U7697 (N_7697,N_6111,N_6758);
xor U7698 (N_7698,N_6806,N_6401);
and U7699 (N_7699,N_6506,N_6585);
nor U7700 (N_7700,N_6743,N_6068);
nor U7701 (N_7701,N_6171,N_6097);
or U7702 (N_7702,N_6924,N_6273);
xor U7703 (N_7703,N_6942,N_6954);
xor U7704 (N_7704,N_6954,N_6331);
nor U7705 (N_7705,N_6351,N_6396);
and U7706 (N_7706,N_6327,N_6757);
nor U7707 (N_7707,N_6822,N_6054);
or U7708 (N_7708,N_6319,N_6702);
and U7709 (N_7709,N_6674,N_6128);
or U7710 (N_7710,N_6618,N_6160);
xnor U7711 (N_7711,N_6988,N_6476);
xor U7712 (N_7712,N_6374,N_6185);
or U7713 (N_7713,N_6485,N_6742);
and U7714 (N_7714,N_6024,N_6268);
nor U7715 (N_7715,N_6848,N_6498);
nand U7716 (N_7716,N_6421,N_6240);
nand U7717 (N_7717,N_6611,N_6129);
nand U7718 (N_7718,N_6442,N_6510);
nor U7719 (N_7719,N_6606,N_6014);
and U7720 (N_7720,N_6898,N_6689);
xor U7721 (N_7721,N_6000,N_6372);
or U7722 (N_7722,N_6283,N_6432);
nor U7723 (N_7723,N_6172,N_6693);
and U7724 (N_7724,N_6045,N_6035);
and U7725 (N_7725,N_6665,N_6502);
nand U7726 (N_7726,N_6845,N_6838);
or U7727 (N_7727,N_6017,N_6437);
or U7728 (N_7728,N_6650,N_6782);
nor U7729 (N_7729,N_6766,N_6640);
or U7730 (N_7730,N_6908,N_6880);
nand U7731 (N_7731,N_6221,N_6249);
xor U7732 (N_7732,N_6526,N_6344);
or U7733 (N_7733,N_6064,N_6721);
and U7734 (N_7734,N_6706,N_6272);
xnor U7735 (N_7735,N_6820,N_6308);
or U7736 (N_7736,N_6321,N_6080);
nor U7737 (N_7737,N_6931,N_6911);
and U7738 (N_7738,N_6069,N_6260);
xnor U7739 (N_7739,N_6714,N_6543);
nor U7740 (N_7740,N_6981,N_6643);
nand U7741 (N_7741,N_6817,N_6389);
xnor U7742 (N_7742,N_6010,N_6979);
xor U7743 (N_7743,N_6165,N_6181);
nor U7744 (N_7744,N_6426,N_6524);
and U7745 (N_7745,N_6926,N_6261);
or U7746 (N_7746,N_6263,N_6405);
or U7747 (N_7747,N_6197,N_6150);
and U7748 (N_7748,N_6012,N_6106);
nor U7749 (N_7749,N_6845,N_6310);
nor U7750 (N_7750,N_6468,N_6899);
and U7751 (N_7751,N_6671,N_6100);
xor U7752 (N_7752,N_6918,N_6726);
and U7753 (N_7753,N_6136,N_6849);
or U7754 (N_7754,N_6615,N_6485);
xor U7755 (N_7755,N_6553,N_6876);
nor U7756 (N_7756,N_6689,N_6266);
nand U7757 (N_7757,N_6167,N_6240);
nand U7758 (N_7758,N_6854,N_6445);
nor U7759 (N_7759,N_6298,N_6364);
nor U7760 (N_7760,N_6817,N_6737);
nor U7761 (N_7761,N_6201,N_6779);
xor U7762 (N_7762,N_6257,N_6829);
nand U7763 (N_7763,N_6936,N_6311);
or U7764 (N_7764,N_6058,N_6803);
nor U7765 (N_7765,N_6185,N_6620);
or U7766 (N_7766,N_6954,N_6874);
or U7767 (N_7767,N_6643,N_6897);
nor U7768 (N_7768,N_6414,N_6904);
and U7769 (N_7769,N_6086,N_6674);
nand U7770 (N_7770,N_6586,N_6302);
xnor U7771 (N_7771,N_6196,N_6369);
xnor U7772 (N_7772,N_6339,N_6459);
nor U7773 (N_7773,N_6442,N_6151);
xnor U7774 (N_7774,N_6791,N_6954);
nor U7775 (N_7775,N_6112,N_6890);
xnor U7776 (N_7776,N_6982,N_6632);
nand U7777 (N_7777,N_6253,N_6070);
nor U7778 (N_7778,N_6249,N_6981);
xnor U7779 (N_7779,N_6058,N_6812);
nor U7780 (N_7780,N_6434,N_6650);
xor U7781 (N_7781,N_6458,N_6885);
and U7782 (N_7782,N_6550,N_6825);
and U7783 (N_7783,N_6387,N_6942);
nand U7784 (N_7784,N_6879,N_6152);
or U7785 (N_7785,N_6521,N_6261);
nor U7786 (N_7786,N_6015,N_6067);
nor U7787 (N_7787,N_6746,N_6869);
nor U7788 (N_7788,N_6540,N_6964);
and U7789 (N_7789,N_6931,N_6561);
or U7790 (N_7790,N_6728,N_6870);
xnor U7791 (N_7791,N_6037,N_6710);
and U7792 (N_7792,N_6125,N_6840);
nand U7793 (N_7793,N_6092,N_6808);
nand U7794 (N_7794,N_6470,N_6526);
or U7795 (N_7795,N_6677,N_6074);
nand U7796 (N_7796,N_6683,N_6628);
nor U7797 (N_7797,N_6235,N_6357);
and U7798 (N_7798,N_6345,N_6659);
nor U7799 (N_7799,N_6650,N_6159);
nand U7800 (N_7800,N_6408,N_6957);
and U7801 (N_7801,N_6324,N_6909);
and U7802 (N_7802,N_6919,N_6439);
xor U7803 (N_7803,N_6254,N_6695);
and U7804 (N_7804,N_6709,N_6859);
or U7805 (N_7805,N_6735,N_6285);
or U7806 (N_7806,N_6445,N_6317);
nand U7807 (N_7807,N_6946,N_6289);
nand U7808 (N_7808,N_6770,N_6989);
nor U7809 (N_7809,N_6680,N_6510);
xnor U7810 (N_7810,N_6548,N_6150);
xor U7811 (N_7811,N_6630,N_6127);
nand U7812 (N_7812,N_6224,N_6494);
and U7813 (N_7813,N_6489,N_6233);
or U7814 (N_7814,N_6859,N_6731);
xnor U7815 (N_7815,N_6672,N_6589);
and U7816 (N_7816,N_6934,N_6026);
nand U7817 (N_7817,N_6356,N_6369);
nand U7818 (N_7818,N_6976,N_6800);
or U7819 (N_7819,N_6946,N_6830);
or U7820 (N_7820,N_6576,N_6616);
or U7821 (N_7821,N_6208,N_6852);
and U7822 (N_7822,N_6469,N_6382);
nor U7823 (N_7823,N_6157,N_6429);
and U7824 (N_7824,N_6455,N_6328);
nand U7825 (N_7825,N_6047,N_6015);
or U7826 (N_7826,N_6795,N_6999);
xor U7827 (N_7827,N_6027,N_6583);
xnor U7828 (N_7828,N_6087,N_6377);
and U7829 (N_7829,N_6931,N_6000);
or U7830 (N_7830,N_6721,N_6920);
and U7831 (N_7831,N_6221,N_6070);
and U7832 (N_7832,N_6865,N_6251);
xnor U7833 (N_7833,N_6446,N_6514);
and U7834 (N_7834,N_6102,N_6350);
xor U7835 (N_7835,N_6468,N_6091);
nand U7836 (N_7836,N_6680,N_6571);
nand U7837 (N_7837,N_6081,N_6476);
and U7838 (N_7838,N_6833,N_6125);
and U7839 (N_7839,N_6436,N_6983);
nor U7840 (N_7840,N_6390,N_6050);
xor U7841 (N_7841,N_6283,N_6412);
nand U7842 (N_7842,N_6797,N_6661);
nand U7843 (N_7843,N_6174,N_6519);
xor U7844 (N_7844,N_6815,N_6638);
nand U7845 (N_7845,N_6677,N_6893);
or U7846 (N_7846,N_6167,N_6732);
or U7847 (N_7847,N_6229,N_6670);
and U7848 (N_7848,N_6694,N_6589);
or U7849 (N_7849,N_6198,N_6005);
nand U7850 (N_7850,N_6954,N_6474);
nor U7851 (N_7851,N_6954,N_6130);
xnor U7852 (N_7852,N_6728,N_6479);
nor U7853 (N_7853,N_6954,N_6350);
or U7854 (N_7854,N_6084,N_6387);
and U7855 (N_7855,N_6861,N_6410);
xor U7856 (N_7856,N_6406,N_6578);
and U7857 (N_7857,N_6581,N_6091);
xor U7858 (N_7858,N_6451,N_6207);
and U7859 (N_7859,N_6534,N_6394);
nand U7860 (N_7860,N_6443,N_6399);
xor U7861 (N_7861,N_6611,N_6081);
nand U7862 (N_7862,N_6898,N_6325);
nor U7863 (N_7863,N_6832,N_6727);
and U7864 (N_7864,N_6383,N_6410);
and U7865 (N_7865,N_6126,N_6966);
nand U7866 (N_7866,N_6958,N_6119);
nand U7867 (N_7867,N_6534,N_6594);
xor U7868 (N_7868,N_6033,N_6037);
nand U7869 (N_7869,N_6484,N_6468);
xor U7870 (N_7870,N_6498,N_6860);
xor U7871 (N_7871,N_6221,N_6323);
nor U7872 (N_7872,N_6665,N_6470);
nor U7873 (N_7873,N_6311,N_6431);
nor U7874 (N_7874,N_6885,N_6031);
nand U7875 (N_7875,N_6125,N_6735);
or U7876 (N_7876,N_6272,N_6368);
nor U7877 (N_7877,N_6326,N_6947);
and U7878 (N_7878,N_6015,N_6995);
nand U7879 (N_7879,N_6284,N_6098);
nand U7880 (N_7880,N_6258,N_6016);
and U7881 (N_7881,N_6048,N_6031);
nor U7882 (N_7882,N_6640,N_6669);
and U7883 (N_7883,N_6275,N_6522);
or U7884 (N_7884,N_6768,N_6287);
nand U7885 (N_7885,N_6275,N_6131);
xnor U7886 (N_7886,N_6209,N_6454);
and U7887 (N_7887,N_6370,N_6980);
nor U7888 (N_7888,N_6373,N_6734);
or U7889 (N_7889,N_6874,N_6161);
or U7890 (N_7890,N_6724,N_6105);
nand U7891 (N_7891,N_6350,N_6275);
and U7892 (N_7892,N_6884,N_6684);
nor U7893 (N_7893,N_6583,N_6485);
nor U7894 (N_7894,N_6340,N_6540);
and U7895 (N_7895,N_6161,N_6918);
xor U7896 (N_7896,N_6087,N_6763);
xor U7897 (N_7897,N_6786,N_6227);
and U7898 (N_7898,N_6911,N_6712);
nand U7899 (N_7899,N_6773,N_6095);
or U7900 (N_7900,N_6232,N_6347);
xor U7901 (N_7901,N_6242,N_6639);
nand U7902 (N_7902,N_6017,N_6053);
nor U7903 (N_7903,N_6378,N_6747);
xnor U7904 (N_7904,N_6136,N_6282);
or U7905 (N_7905,N_6442,N_6933);
nand U7906 (N_7906,N_6125,N_6353);
or U7907 (N_7907,N_6043,N_6763);
xor U7908 (N_7908,N_6700,N_6273);
xnor U7909 (N_7909,N_6102,N_6587);
xor U7910 (N_7910,N_6664,N_6412);
and U7911 (N_7911,N_6957,N_6657);
xnor U7912 (N_7912,N_6910,N_6425);
xor U7913 (N_7913,N_6949,N_6543);
nand U7914 (N_7914,N_6930,N_6030);
nand U7915 (N_7915,N_6334,N_6414);
nor U7916 (N_7916,N_6843,N_6510);
nand U7917 (N_7917,N_6973,N_6310);
nand U7918 (N_7918,N_6115,N_6493);
xnor U7919 (N_7919,N_6298,N_6825);
nand U7920 (N_7920,N_6081,N_6888);
xnor U7921 (N_7921,N_6985,N_6288);
nand U7922 (N_7922,N_6985,N_6247);
xnor U7923 (N_7923,N_6717,N_6973);
or U7924 (N_7924,N_6971,N_6453);
and U7925 (N_7925,N_6411,N_6302);
nand U7926 (N_7926,N_6880,N_6690);
and U7927 (N_7927,N_6815,N_6391);
nand U7928 (N_7928,N_6810,N_6421);
xor U7929 (N_7929,N_6286,N_6158);
nand U7930 (N_7930,N_6670,N_6314);
xnor U7931 (N_7931,N_6013,N_6734);
nor U7932 (N_7932,N_6890,N_6126);
and U7933 (N_7933,N_6878,N_6711);
nand U7934 (N_7934,N_6132,N_6546);
or U7935 (N_7935,N_6724,N_6959);
nand U7936 (N_7936,N_6472,N_6885);
and U7937 (N_7937,N_6503,N_6818);
and U7938 (N_7938,N_6121,N_6442);
or U7939 (N_7939,N_6983,N_6445);
nor U7940 (N_7940,N_6083,N_6595);
nand U7941 (N_7941,N_6612,N_6004);
and U7942 (N_7942,N_6018,N_6501);
xnor U7943 (N_7943,N_6578,N_6313);
xnor U7944 (N_7944,N_6113,N_6470);
nor U7945 (N_7945,N_6873,N_6493);
and U7946 (N_7946,N_6222,N_6506);
nor U7947 (N_7947,N_6789,N_6707);
and U7948 (N_7948,N_6791,N_6268);
nor U7949 (N_7949,N_6170,N_6553);
xor U7950 (N_7950,N_6445,N_6027);
nor U7951 (N_7951,N_6217,N_6596);
nand U7952 (N_7952,N_6525,N_6393);
nand U7953 (N_7953,N_6155,N_6619);
or U7954 (N_7954,N_6864,N_6776);
xor U7955 (N_7955,N_6070,N_6282);
and U7956 (N_7956,N_6099,N_6501);
nand U7957 (N_7957,N_6096,N_6436);
nand U7958 (N_7958,N_6298,N_6823);
xnor U7959 (N_7959,N_6930,N_6510);
or U7960 (N_7960,N_6897,N_6890);
or U7961 (N_7961,N_6020,N_6870);
nand U7962 (N_7962,N_6612,N_6379);
xor U7963 (N_7963,N_6714,N_6460);
and U7964 (N_7964,N_6029,N_6917);
nand U7965 (N_7965,N_6894,N_6622);
nand U7966 (N_7966,N_6618,N_6577);
nand U7967 (N_7967,N_6964,N_6982);
nor U7968 (N_7968,N_6514,N_6336);
xor U7969 (N_7969,N_6285,N_6140);
xnor U7970 (N_7970,N_6341,N_6322);
and U7971 (N_7971,N_6124,N_6259);
xor U7972 (N_7972,N_6348,N_6691);
nor U7973 (N_7973,N_6128,N_6086);
or U7974 (N_7974,N_6416,N_6989);
nor U7975 (N_7975,N_6160,N_6827);
and U7976 (N_7976,N_6872,N_6731);
xnor U7977 (N_7977,N_6661,N_6636);
or U7978 (N_7978,N_6250,N_6858);
and U7979 (N_7979,N_6765,N_6146);
and U7980 (N_7980,N_6190,N_6292);
and U7981 (N_7981,N_6950,N_6689);
and U7982 (N_7982,N_6959,N_6624);
nand U7983 (N_7983,N_6843,N_6787);
nor U7984 (N_7984,N_6033,N_6645);
nor U7985 (N_7985,N_6412,N_6685);
nor U7986 (N_7986,N_6929,N_6003);
xnor U7987 (N_7987,N_6340,N_6620);
and U7988 (N_7988,N_6725,N_6165);
xnor U7989 (N_7989,N_6737,N_6846);
or U7990 (N_7990,N_6769,N_6534);
nor U7991 (N_7991,N_6035,N_6311);
xor U7992 (N_7992,N_6815,N_6101);
nand U7993 (N_7993,N_6991,N_6568);
or U7994 (N_7994,N_6248,N_6491);
nor U7995 (N_7995,N_6070,N_6663);
nor U7996 (N_7996,N_6852,N_6676);
or U7997 (N_7997,N_6121,N_6382);
and U7998 (N_7998,N_6274,N_6032);
xor U7999 (N_7999,N_6652,N_6621);
xnor U8000 (N_8000,N_7689,N_7168);
or U8001 (N_8001,N_7761,N_7909);
or U8002 (N_8002,N_7192,N_7637);
xor U8003 (N_8003,N_7634,N_7413);
nor U8004 (N_8004,N_7996,N_7845);
nor U8005 (N_8005,N_7812,N_7514);
nor U8006 (N_8006,N_7276,N_7862);
nand U8007 (N_8007,N_7341,N_7694);
or U8008 (N_8008,N_7542,N_7858);
nor U8009 (N_8009,N_7839,N_7199);
nor U8010 (N_8010,N_7834,N_7850);
nand U8011 (N_8011,N_7213,N_7553);
or U8012 (N_8012,N_7280,N_7063);
and U8013 (N_8013,N_7976,N_7952);
and U8014 (N_8014,N_7030,N_7823);
nand U8015 (N_8015,N_7773,N_7581);
nor U8016 (N_8016,N_7854,N_7136);
and U8017 (N_8017,N_7599,N_7535);
xor U8018 (N_8018,N_7086,N_7620);
and U8019 (N_8019,N_7264,N_7505);
xor U8020 (N_8020,N_7272,N_7093);
or U8021 (N_8021,N_7540,N_7965);
or U8022 (N_8022,N_7920,N_7071);
xor U8023 (N_8023,N_7519,N_7717);
nor U8024 (N_8024,N_7632,N_7495);
and U8025 (N_8025,N_7431,N_7922);
nor U8026 (N_8026,N_7309,N_7810);
or U8027 (N_8027,N_7859,N_7066);
nor U8028 (N_8028,N_7225,N_7851);
and U8029 (N_8029,N_7143,N_7270);
xnor U8030 (N_8030,N_7550,N_7869);
nand U8031 (N_8031,N_7630,N_7307);
nor U8032 (N_8032,N_7652,N_7334);
nor U8033 (N_8033,N_7158,N_7041);
xnor U8034 (N_8034,N_7017,N_7035);
or U8035 (N_8035,N_7575,N_7001);
nand U8036 (N_8036,N_7663,N_7008);
xnor U8037 (N_8037,N_7672,N_7662);
or U8038 (N_8038,N_7464,N_7569);
nand U8039 (N_8039,N_7322,N_7527);
xnor U8040 (N_8040,N_7200,N_7275);
nor U8041 (N_8041,N_7049,N_7462);
xor U8042 (N_8042,N_7215,N_7872);
or U8043 (N_8043,N_7292,N_7233);
or U8044 (N_8044,N_7410,N_7353);
and U8045 (N_8045,N_7139,N_7611);
xnor U8046 (N_8046,N_7053,N_7202);
nor U8047 (N_8047,N_7148,N_7586);
xor U8048 (N_8048,N_7301,N_7019);
xor U8049 (N_8049,N_7696,N_7926);
nand U8050 (N_8050,N_7616,N_7991);
nor U8051 (N_8051,N_7409,N_7172);
nor U8052 (N_8052,N_7837,N_7546);
xnor U8053 (N_8053,N_7428,N_7325);
or U8054 (N_8054,N_7956,N_7140);
nand U8055 (N_8055,N_7848,N_7348);
or U8056 (N_8056,N_7960,N_7508);
and U8057 (N_8057,N_7877,N_7828);
nor U8058 (N_8058,N_7981,N_7602);
or U8059 (N_8059,N_7479,N_7510);
xnor U8060 (N_8060,N_7782,N_7561);
nand U8061 (N_8061,N_7890,N_7282);
and U8062 (N_8062,N_7372,N_7310);
or U8063 (N_8063,N_7523,N_7031);
xor U8064 (N_8064,N_7627,N_7929);
xnor U8065 (N_8065,N_7499,N_7695);
xor U8066 (N_8066,N_7313,N_7798);
nand U8067 (N_8067,N_7600,N_7359);
or U8068 (N_8068,N_7246,N_7084);
nor U8069 (N_8069,N_7911,N_7622);
nand U8070 (N_8070,N_7398,N_7323);
nor U8071 (N_8071,N_7746,N_7385);
and U8072 (N_8072,N_7285,N_7430);
xnor U8073 (N_8073,N_7653,N_7152);
or U8074 (N_8074,N_7950,N_7161);
or U8075 (N_8075,N_7463,N_7432);
nand U8076 (N_8076,N_7389,N_7083);
and U8077 (N_8077,N_7393,N_7394);
and U8078 (N_8078,N_7978,N_7186);
nand U8079 (N_8079,N_7294,N_7601);
xor U8080 (N_8080,N_7524,N_7931);
and U8081 (N_8081,N_7791,N_7090);
xnor U8082 (N_8082,N_7688,N_7603);
and U8083 (N_8083,N_7496,N_7594);
or U8084 (N_8084,N_7466,N_7554);
nor U8085 (N_8085,N_7818,N_7414);
xor U8086 (N_8086,N_7806,N_7450);
or U8087 (N_8087,N_7335,N_7261);
nor U8088 (N_8088,N_7932,N_7787);
and U8089 (N_8089,N_7470,N_7649);
nand U8090 (N_8090,N_7291,N_7945);
nand U8091 (N_8091,N_7918,N_7075);
and U8092 (N_8092,N_7775,N_7238);
or U8093 (N_8093,N_7897,N_7260);
nand U8094 (N_8094,N_7975,N_7296);
and U8095 (N_8095,N_7091,N_7486);
or U8096 (N_8096,N_7942,N_7183);
nand U8097 (N_8097,N_7244,N_7390);
and U8098 (N_8098,N_7191,N_7580);
nand U8099 (N_8099,N_7420,N_7239);
xnor U8100 (N_8100,N_7661,N_7752);
xor U8101 (N_8101,N_7279,N_7631);
and U8102 (N_8102,N_7471,N_7165);
or U8103 (N_8103,N_7009,N_7706);
or U8104 (N_8104,N_7194,N_7311);
nand U8105 (N_8105,N_7779,N_7357);
nor U8106 (N_8106,N_7465,N_7349);
xnor U8107 (N_8107,N_7740,N_7843);
nor U8108 (N_8108,N_7832,N_7125);
xnor U8109 (N_8109,N_7317,N_7059);
and U8110 (N_8110,N_7175,N_7456);
xor U8111 (N_8111,N_7055,N_7884);
nand U8112 (N_8112,N_7720,N_7380);
nor U8113 (N_8113,N_7392,N_7182);
nand U8114 (N_8114,N_7644,N_7697);
nand U8115 (N_8115,N_7951,N_7217);
and U8116 (N_8116,N_7343,N_7972);
nor U8117 (N_8117,N_7331,N_7724);
or U8118 (N_8118,N_7185,N_7676);
or U8119 (N_8119,N_7370,N_7794);
xor U8120 (N_8120,N_7024,N_7683);
nand U8121 (N_8121,N_7081,N_7352);
xor U8122 (N_8122,N_7014,N_7536);
nand U8123 (N_8123,N_7351,N_7226);
and U8124 (N_8124,N_7153,N_7783);
or U8125 (N_8125,N_7994,N_7937);
nand U8126 (N_8126,N_7589,N_7028);
and U8127 (N_8127,N_7820,N_7895);
and U8128 (N_8128,N_7485,N_7765);
nand U8129 (N_8129,N_7003,N_7670);
nand U8130 (N_8130,N_7615,N_7484);
and U8131 (N_8131,N_7777,N_7566);
or U8132 (N_8132,N_7189,N_7145);
nand U8133 (N_8133,N_7367,N_7381);
xnor U8134 (N_8134,N_7814,N_7660);
nand U8135 (N_8135,N_7744,N_7767);
nor U8136 (N_8136,N_7668,N_7618);
and U8137 (N_8137,N_7416,N_7210);
xor U8138 (N_8138,N_7598,N_7736);
xor U8139 (N_8139,N_7907,N_7224);
nor U8140 (N_8140,N_7005,N_7501);
or U8141 (N_8141,N_7048,N_7924);
nand U8142 (N_8142,N_7474,N_7707);
or U8143 (N_8143,N_7747,N_7541);
and U8144 (N_8144,N_7915,N_7154);
or U8145 (N_8145,N_7328,N_7312);
xnor U8146 (N_8146,N_7570,N_7281);
xnor U8147 (N_8147,N_7849,N_7982);
and U8148 (N_8148,N_7841,N_7677);
or U8149 (N_8149,N_7080,N_7129);
nand U8150 (N_8150,N_7111,N_7026);
or U8151 (N_8151,N_7399,N_7231);
nand U8152 (N_8152,N_7229,N_7050);
or U8153 (N_8153,N_7565,N_7072);
and U8154 (N_8154,N_7476,N_7838);
or U8155 (N_8155,N_7784,N_7891);
xor U8156 (N_8156,N_7875,N_7032);
and U8157 (N_8157,N_7273,N_7101);
or U8158 (N_8158,N_7252,N_7815);
xnor U8159 (N_8159,N_7330,N_7711);
nand U8160 (N_8160,N_7408,N_7308);
nand U8161 (N_8161,N_7984,N_7864);
nand U8162 (N_8162,N_7971,N_7641);
nor U8163 (N_8163,N_7625,N_7218);
xor U8164 (N_8164,N_7811,N_7443);
xor U8165 (N_8165,N_7852,N_7135);
nand U8166 (N_8166,N_7214,N_7504);
nand U8167 (N_8167,N_7481,N_7137);
nand U8168 (N_8168,N_7657,N_7089);
and U8169 (N_8169,N_7977,N_7721);
xnor U8170 (N_8170,N_7648,N_7656);
xnor U8171 (N_8171,N_7898,N_7962);
and U8172 (N_8172,N_7572,N_7954);
or U8173 (N_8173,N_7776,N_7635);
and U8174 (N_8174,N_7303,N_7650);
or U8175 (N_8175,N_7769,N_7167);
or U8176 (N_8176,N_7449,N_7438);
and U8177 (N_8177,N_7442,N_7404);
or U8178 (N_8178,N_7680,N_7057);
or U8179 (N_8179,N_7219,N_7873);
and U8180 (N_8180,N_7012,N_7521);
and U8181 (N_8181,N_7755,N_7813);
and U8182 (N_8182,N_7423,N_7262);
and U8183 (N_8183,N_7468,N_7989);
nand U8184 (N_8184,N_7729,N_7847);
and U8185 (N_8185,N_7560,N_7558);
nand U8186 (N_8186,N_7265,N_7062);
and U8187 (N_8187,N_7685,N_7100);
or U8188 (N_8188,N_7467,N_7245);
xor U8189 (N_8189,N_7665,N_7120);
nor U8190 (N_8190,N_7636,N_7318);
nand U8191 (N_8191,N_7029,N_7056);
and U8192 (N_8192,N_7251,N_7248);
nand U8193 (N_8193,N_7610,N_7574);
xnor U8194 (N_8194,N_7065,N_7157);
xor U8195 (N_8195,N_7402,N_7118);
xnor U8196 (N_8196,N_7206,N_7444);
and U8197 (N_8197,N_7520,N_7039);
nand U8198 (N_8198,N_7439,N_7133);
or U8199 (N_8199,N_7726,N_7347);
and U8200 (N_8200,N_7958,N_7534);
and U8201 (N_8201,N_7860,N_7802);
xor U8202 (N_8202,N_7435,N_7959);
and U8203 (N_8203,N_7743,N_7916);
nor U8204 (N_8204,N_7617,N_7461);
and U8205 (N_8205,N_7293,N_7588);
nand U8206 (N_8206,N_7104,N_7362);
nand U8207 (N_8207,N_7819,N_7422);
nor U8208 (N_8208,N_7412,N_7447);
xnor U8209 (N_8209,N_7543,N_7758);
and U8210 (N_8210,N_7336,N_7259);
or U8211 (N_8211,N_7830,N_7078);
and U8212 (N_8212,N_7639,N_7342);
xnor U8213 (N_8213,N_7522,N_7095);
or U8214 (N_8214,N_7256,N_7786);
and U8215 (N_8215,N_7337,N_7940);
or U8216 (N_8216,N_7705,N_7608);
and U8217 (N_8217,N_7356,N_7770);
or U8218 (N_8218,N_7419,N_7446);
nand U8219 (N_8219,N_7400,N_7421);
nand U8220 (N_8220,N_7228,N_7223);
and U8221 (N_8221,N_7516,N_7320);
nor U8222 (N_8222,N_7856,N_7271);
nor U8223 (N_8223,N_7339,N_7730);
and U8224 (N_8224,N_7824,N_7562);
or U8225 (N_8225,N_7868,N_7816);
xnor U8226 (N_8226,N_7759,N_7160);
nor U8227 (N_8227,N_7910,N_7299);
nor U8228 (N_8228,N_7426,N_7240);
nand U8229 (N_8229,N_7905,N_7295);
nand U8230 (N_8230,N_7013,N_7193);
or U8231 (N_8231,N_7124,N_7314);
xnor U8232 (N_8232,N_7757,N_7497);
nor U8233 (N_8233,N_7427,N_7908);
or U8234 (N_8234,N_7332,N_7621);
and U8235 (N_8235,N_7941,N_7258);
xnor U8236 (N_8236,N_7097,N_7300);
or U8237 (N_8237,N_7025,N_7038);
and U8238 (N_8238,N_7483,N_7712);
xor U8239 (N_8239,N_7804,N_7764);
nor U8240 (N_8240,N_7725,N_7582);
nor U8241 (N_8241,N_7990,N_7876);
xnor U8242 (N_8242,N_7731,N_7007);
nand U8243 (N_8243,N_7209,N_7079);
or U8244 (N_8244,N_7691,N_7604);
nor U8245 (N_8245,N_7774,N_7045);
and U8246 (N_8246,N_7887,N_7762);
and U8247 (N_8247,N_7983,N_7267);
and U8248 (N_8248,N_7568,N_7119);
xnor U8249 (N_8249,N_7623,N_7173);
xnor U8250 (N_8250,N_7290,N_7452);
nor U8251 (N_8251,N_7405,N_7675);
or U8252 (N_8252,N_7187,N_7638);
nand U8253 (N_8253,N_7808,N_7022);
and U8254 (N_8254,N_7042,N_7664);
nand U8255 (N_8255,N_7064,N_7344);
nand U8256 (N_8256,N_7987,N_7211);
xnor U8257 (N_8257,N_7180,N_7809);
and U8258 (N_8258,N_7247,N_7387);
xor U8259 (N_8259,N_7948,N_7571);
nand U8260 (N_8260,N_7943,N_7181);
xnor U8261 (N_8261,N_7678,N_7236);
and U8262 (N_8262,N_7242,N_7122);
and U8263 (N_8263,N_7197,N_7878);
nand U8264 (N_8264,N_7533,N_7130);
nor U8265 (N_8265,N_7174,N_7624);
xnor U8266 (N_8266,N_7961,N_7988);
nor U8267 (N_8267,N_7805,N_7741);
and U8268 (N_8268,N_7366,N_7365);
xnor U8269 (N_8269,N_7052,N_7844);
and U8270 (N_8270,N_7684,N_7425);
or U8271 (N_8271,N_7278,N_7556);
xor U8272 (N_8272,N_7107,N_7980);
xor U8273 (N_8273,N_7377,N_7358);
or U8274 (N_8274,N_7376,N_7583);
nand U8275 (N_8275,N_7885,N_7096);
xor U8276 (N_8276,N_7609,N_7208);
or U8277 (N_8277,N_7861,N_7249);
nand U8278 (N_8278,N_7973,N_7492);
nor U8279 (N_8279,N_7115,N_7526);
or U8280 (N_8280,N_7698,N_7826);
and U8281 (N_8281,N_7350,N_7947);
xnor U8282 (N_8282,N_7306,N_7188);
and U8283 (N_8283,N_7595,N_7445);
and U8284 (N_8284,N_7667,N_7298);
or U8285 (N_8285,N_7645,N_7169);
xnor U8286 (N_8286,N_7138,N_7655);
or U8287 (N_8287,N_7482,N_7727);
nand U8288 (N_8288,N_7195,N_7424);
nand U8289 (N_8289,N_7459,N_7997);
or U8290 (N_8290,N_7530,N_7551);
nand U8291 (N_8291,N_7612,N_7379);
and U8292 (N_8292,N_7255,N_7333);
nor U8293 (N_8293,N_7509,N_7305);
xnor U8294 (N_8294,N_7383,N_7478);
nand U8295 (N_8295,N_7870,N_7538);
or U8296 (N_8296,N_7525,N_7647);
and U8297 (N_8297,N_7099,N_7204);
xor U8298 (N_8298,N_7375,N_7319);
xnor U8299 (N_8299,N_7156,N_7790);
nor U8300 (N_8300,N_7894,N_7857);
and U8301 (N_8301,N_7781,N_7092);
or U8302 (N_8302,N_7709,N_7957);
nand U8303 (N_8303,N_7585,N_7250);
or U8304 (N_8304,N_7529,N_7407);
xor U8305 (N_8305,N_7498,N_7728);
nand U8306 (N_8306,N_7114,N_7701);
xnor U8307 (N_8307,N_7106,N_7513);
nand U8308 (N_8308,N_7902,N_7555);
nor U8309 (N_8309,N_7640,N_7102);
nand U8310 (N_8310,N_7666,N_7455);
nor U8311 (N_8311,N_7360,N_7179);
xor U8312 (N_8312,N_7734,N_7437);
or U8313 (N_8313,N_7141,N_7171);
or U8314 (N_8314,N_7692,N_7198);
nand U8315 (N_8315,N_7888,N_7998);
and U8316 (N_8316,N_7719,N_7490);
nand U8317 (N_8317,N_7355,N_7077);
nand U8318 (N_8318,N_7596,N_7220);
and U8319 (N_8319,N_7605,N_7853);
nand U8320 (N_8320,N_7833,N_7472);
nor U8321 (N_8321,N_7087,N_7900);
and U8322 (N_8322,N_7682,N_7715);
or U8323 (N_8323,N_7531,N_7708);
nand U8324 (N_8324,N_7874,N_7807);
and U8325 (N_8325,N_7286,N_7302);
nor U8326 (N_8326,N_7563,N_7283);
or U8327 (N_8327,N_7263,N_7934);
nor U8328 (N_8328,N_7974,N_7345);
and U8329 (N_8329,N_7879,N_7713);
or U8330 (N_8330,N_7254,N_7723);
and U8331 (N_8331,N_7234,N_7243);
nand U8332 (N_8332,N_7027,N_7034);
nand U8333 (N_8333,N_7166,N_7502);
nor U8334 (N_8334,N_7544,N_7257);
nand U8335 (N_8335,N_7069,N_7315);
nand U8336 (N_8336,N_7939,N_7127);
nand U8337 (N_8337,N_7590,N_7871);
and U8338 (N_8338,N_7722,N_7793);
nor U8339 (N_8339,N_7458,N_7411);
and U8340 (N_8340,N_7364,N_7576);
or U8341 (N_8341,N_7216,N_7235);
or U8342 (N_8342,N_7768,N_7018);
nor U8343 (N_8343,N_7919,N_7037);
nor U8344 (N_8344,N_7241,N_7528);
xor U8345 (N_8345,N_7789,N_7651);
or U8346 (N_8346,N_7825,N_7395);
nor U8347 (N_8347,N_7201,N_7477);
and U8348 (N_8348,N_7796,N_7454);
nor U8349 (N_8349,N_7134,N_7548);
nor U8350 (N_8350,N_7113,N_7488);
nor U8351 (N_8351,N_7170,N_7763);
xnor U8352 (N_8352,N_7440,N_7797);
nor U8353 (N_8353,N_7396,N_7326);
xnor U8354 (N_8354,N_7840,N_7274);
nor U8355 (N_8355,N_7040,N_7354);
and U8356 (N_8356,N_7591,N_7184);
nor U8357 (N_8357,N_7044,N_7659);
or U8358 (N_8358,N_7033,N_7906);
xnor U8359 (N_8359,N_7110,N_7517);
xnor U8360 (N_8360,N_7493,N_7710);
and U8361 (N_8361,N_7142,N_7817);
nand U8362 (N_8362,N_7094,N_7923);
nor U8363 (N_8363,N_7964,N_7889);
or U8364 (N_8364,N_7995,N_7117);
nor U8365 (N_8365,N_7015,N_7147);
nand U8366 (N_8366,N_7384,N_7549);
or U8367 (N_8367,N_7737,N_7867);
or U8368 (N_8368,N_7803,N_7968);
or U8369 (N_8369,N_7748,N_7979);
xor U8370 (N_8370,N_7732,N_7966);
nand U8371 (N_8371,N_7883,N_7654);
nor U8372 (N_8372,N_7785,N_7011);
nor U8373 (N_8373,N_7992,N_7999);
xor U8374 (N_8374,N_7382,N_7406);
and U8375 (N_8375,N_7739,N_7150);
nor U8376 (N_8376,N_7938,N_7606);
xnor U8377 (N_8377,N_7503,N_7512);
nor U8378 (N_8378,N_7750,N_7700);
and U8379 (N_8379,N_7196,N_7237);
or U8380 (N_8380,N_7917,N_7340);
or U8381 (N_8381,N_7453,N_7567);
xnor U8382 (N_8382,N_7855,N_7088);
and U8383 (N_8383,N_7500,N_7587);
xnor U8384 (N_8384,N_7842,N_7036);
xnor U8385 (N_8385,N_7674,N_7579);
and U8386 (N_8386,N_7105,N_7103);
xnor U8387 (N_8387,N_7388,N_7614);
nand U8388 (N_8388,N_7949,N_7827);
nand U8389 (N_8389,N_7953,N_7266);
xnor U8390 (N_8390,N_7441,N_7061);
xnor U8391 (N_8391,N_7108,N_7778);
nor U8392 (N_8392,N_7821,N_7899);
or U8393 (N_8393,N_7268,N_7159);
nand U8394 (N_8394,N_7829,N_7021);
xnor U8395 (N_8395,N_7002,N_7232);
nor U8396 (N_8396,N_7658,N_7151);
nor U8397 (N_8397,N_7507,N_7368);
or U8398 (N_8398,N_7126,N_7970);
and U8399 (N_8399,N_7491,N_7836);
xnor U8400 (N_8400,N_7799,N_7116);
nor U8401 (N_8401,N_7760,N_7936);
nand U8402 (N_8402,N_7112,N_7448);
nand U8403 (N_8403,N_7363,N_7155);
and U8404 (N_8404,N_7163,N_7628);
or U8405 (N_8405,N_7304,N_7986);
nand U8406 (N_8406,N_7955,N_7434);
nor U8407 (N_8407,N_7054,N_7573);
nor U8408 (N_8408,N_7020,N_7880);
and U8409 (N_8409,N_7288,N_7903);
xnor U8410 (N_8410,N_7532,N_7000);
nor U8411 (N_8411,N_7597,N_7329);
or U8412 (N_8412,N_7967,N_7010);
nand U8413 (N_8413,N_7742,N_7754);
nor U8414 (N_8414,N_7494,N_7378);
or U8415 (N_8415,N_7515,N_7386);
xnor U8416 (N_8416,N_7128,N_7073);
nand U8417 (N_8417,N_7074,N_7969);
nor U8418 (N_8418,N_7703,N_7222);
xor U8419 (N_8419,N_7993,N_7480);
and U8420 (N_8420,N_7646,N_7607);
nand U8421 (N_8421,N_7792,N_7082);
xor U8422 (N_8422,N_7109,N_7207);
nor U8423 (N_8423,N_7946,N_7369);
nor U8424 (N_8424,N_7780,N_7085);
nand U8425 (N_8425,N_7846,N_7788);
nor U8426 (N_8426,N_7702,N_7060);
or U8427 (N_8427,N_7051,N_7253);
or U8428 (N_8428,N_7230,N_7756);
and U8429 (N_8429,N_7417,N_7559);
nand U8430 (N_8430,N_7863,N_7487);
xor U8431 (N_8431,N_7518,N_7578);
nor U8432 (N_8432,N_7429,N_7149);
and U8433 (N_8433,N_7327,N_7047);
and U8434 (N_8434,N_7738,N_7324);
or U8435 (N_8435,N_7436,N_7506);
xnor U8436 (N_8436,N_7391,N_7227);
nand U8437 (N_8437,N_7346,N_7489);
or U8438 (N_8438,N_7552,N_7930);
and U8439 (N_8439,N_7933,N_7537);
nand U8440 (N_8440,N_7212,N_7985);
nand U8441 (N_8441,N_7004,N_7795);
nor U8442 (N_8442,N_7671,N_7433);
nand U8443 (N_8443,N_7800,N_7123);
or U8444 (N_8444,N_7669,N_7178);
or U8445 (N_8445,N_7771,N_7068);
and U8446 (N_8446,N_7475,N_7203);
xnor U8447 (N_8447,N_7944,N_7686);
nand U8448 (N_8448,N_7866,N_7882);
nor U8449 (N_8449,N_7460,N_7374);
xor U8450 (N_8450,N_7629,N_7321);
and U8451 (N_8451,N_7619,N_7690);
nand U8452 (N_8452,N_7023,N_7338);
nor U8453 (N_8453,N_7131,N_7642);
or U8454 (N_8454,N_7892,N_7749);
or U8455 (N_8455,N_7613,N_7545);
and U8456 (N_8456,N_7927,N_7626);
and U8457 (N_8457,N_7896,N_7144);
nor U8458 (N_8458,N_7006,N_7718);
and U8459 (N_8459,N_7557,N_7205);
nor U8460 (N_8460,N_7098,N_7371);
nor U8461 (N_8461,N_7164,N_7162);
xnor U8462 (N_8462,N_7584,N_7733);
nor U8463 (N_8463,N_7177,N_7592);
or U8464 (N_8464,N_7963,N_7146);
nand U8465 (N_8465,N_7067,N_7289);
nand U8466 (N_8466,N_7451,N_7865);
and U8467 (N_8467,N_7547,N_7418);
nand U8468 (N_8468,N_7176,N_7287);
or U8469 (N_8469,N_7886,N_7766);
nor U8470 (N_8470,N_7914,N_7835);
xor U8471 (N_8471,N_7801,N_7046);
nand U8472 (N_8472,N_7673,N_7457);
nor U8473 (N_8473,N_7681,N_7511);
xnor U8474 (N_8474,N_7284,N_7881);
xnor U8475 (N_8475,N_7753,N_7893);
or U8476 (N_8476,N_7132,N_7714);
xor U8477 (N_8477,N_7745,N_7269);
nor U8478 (N_8478,N_7373,N_7577);
nor U8479 (N_8479,N_7822,N_7277);
xor U8480 (N_8480,N_7121,N_7469);
nor U8481 (N_8481,N_7316,N_7901);
nor U8482 (N_8482,N_7564,N_7070);
or U8483 (N_8483,N_7593,N_7735);
xor U8484 (N_8484,N_7058,N_7925);
nor U8485 (N_8485,N_7704,N_7043);
nor U8486 (N_8486,N_7539,N_7190);
nand U8487 (N_8487,N_7687,N_7221);
xor U8488 (N_8488,N_7693,N_7716);
xor U8489 (N_8489,N_7679,N_7928);
or U8490 (N_8490,N_7473,N_7403);
xor U8491 (N_8491,N_7699,N_7935);
or U8492 (N_8492,N_7904,N_7751);
and U8493 (N_8493,N_7831,N_7361);
nand U8494 (N_8494,N_7633,N_7415);
and U8495 (N_8495,N_7397,N_7076);
xor U8496 (N_8496,N_7912,N_7297);
and U8497 (N_8497,N_7016,N_7401);
xnor U8498 (N_8498,N_7772,N_7643);
xor U8499 (N_8499,N_7913,N_7921);
nand U8500 (N_8500,N_7543,N_7154);
nand U8501 (N_8501,N_7891,N_7895);
or U8502 (N_8502,N_7069,N_7890);
nor U8503 (N_8503,N_7118,N_7858);
or U8504 (N_8504,N_7133,N_7813);
or U8505 (N_8505,N_7856,N_7841);
and U8506 (N_8506,N_7859,N_7478);
and U8507 (N_8507,N_7022,N_7245);
nor U8508 (N_8508,N_7591,N_7752);
and U8509 (N_8509,N_7992,N_7844);
and U8510 (N_8510,N_7838,N_7263);
nor U8511 (N_8511,N_7246,N_7985);
xnor U8512 (N_8512,N_7749,N_7012);
nand U8513 (N_8513,N_7923,N_7192);
nor U8514 (N_8514,N_7344,N_7067);
or U8515 (N_8515,N_7280,N_7195);
and U8516 (N_8516,N_7835,N_7321);
xor U8517 (N_8517,N_7782,N_7045);
and U8518 (N_8518,N_7674,N_7410);
nor U8519 (N_8519,N_7575,N_7618);
nor U8520 (N_8520,N_7099,N_7400);
or U8521 (N_8521,N_7645,N_7751);
xnor U8522 (N_8522,N_7452,N_7116);
xnor U8523 (N_8523,N_7466,N_7523);
or U8524 (N_8524,N_7378,N_7273);
or U8525 (N_8525,N_7363,N_7255);
nand U8526 (N_8526,N_7422,N_7345);
nor U8527 (N_8527,N_7874,N_7205);
nor U8528 (N_8528,N_7745,N_7807);
nor U8529 (N_8529,N_7881,N_7733);
nand U8530 (N_8530,N_7939,N_7620);
nor U8531 (N_8531,N_7158,N_7063);
nor U8532 (N_8532,N_7351,N_7208);
xor U8533 (N_8533,N_7970,N_7701);
nor U8534 (N_8534,N_7692,N_7402);
and U8535 (N_8535,N_7506,N_7336);
xnor U8536 (N_8536,N_7827,N_7862);
or U8537 (N_8537,N_7054,N_7440);
xnor U8538 (N_8538,N_7303,N_7440);
nand U8539 (N_8539,N_7589,N_7954);
and U8540 (N_8540,N_7240,N_7165);
nor U8541 (N_8541,N_7793,N_7194);
xnor U8542 (N_8542,N_7391,N_7659);
and U8543 (N_8543,N_7362,N_7698);
and U8544 (N_8544,N_7621,N_7456);
and U8545 (N_8545,N_7512,N_7712);
and U8546 (N_8546,N_7591,N_7799);
or U8547 (N_8547,N_7143,N_7140);
or U8548 (N_8548,N_7597,N_7599);
xor U8549 (N_8549,N_7287,N_7836);
and U8550 (N_8550,N_7469,N_7880);
or U8551 (N_8551,N_7878,N_7184);
and U8552 (N_8552,N_7268,N_7488);
and U8553 (N_8553,N_7101,N_7104);
xnor U8554 (N_8554,N_7487,N_7372);
or U8555 (N_8555,N_7234,N_7227);
nand U8556 (N_8556,N_7802,N_7063);
xor U8557 (N_8557,N_7944,N_7470);
nand U8558 (N_8558,N_7150,N_7078);
and U8559 (N_8559,N_7490,N_7020);
or U8560 (N_8560,N_7078,N_7584);
xor U8561 (N_8561,N_7621,N_7044);
and U8562 (N_8562,N_7357,N_7335);
and U8563 (N_8563,N_7975,N_7372);
nand U8564 (N_8564,N_7758,N_7093);
xor U8565 (N_8565,N_7151,N_7877);
or U8566 (N_8566,N_7211,N_7245);
xnor U8567 (N_8567,N_7973,N_7334);
nor U8568 (N_8568,N_7952,N_7039);
nor U8569 (N_8569,N_7288,N_7513);
and U8570 (N_8570,N_7400,N_7904);
and U8571 (N_8571,N_7990,N_7776);
xnor U8572 (N_8572,N_7301,N_7934);
nand U8573 (N_8573,N_7014,N_7104);
xnor U8574 (N_8574,N_7328,N_7062);
and U8575 (N_8575,N_7322,N_7013);
nor U8576 (N_8576,N_7079,N_7712);
and U8577 (N_8577,N_7436,N_7327);
xnor U8578 (N_8578,N_7455,N_7261);
nor U8579 (N_8579,N_7788,N_7684);
or U8580 (N_8580,N_7954,N_7884);
xor U8581 (N_8581,N_7016,N_7286);
nor U8582 (N_8582,N_7886,N_7232);
nand U8583 (N_8583,N_7146,N_7617);
xor U8584 (N_8584,N_7906,N_7899);
nand U8585 (N_8585,N_7885,N_7545);
or U8586 (N_8586,N_7021,N_7067);
nor U8587 (N_8587,N_7041,N_7766);
and U8588 (N_8588,N_7648,N_7316);
xor U8589 (N_8589,N_7369,N_7210);
nand U8590 (N_8590,N_7221,N_7621);
nor U8591 (N_8591,N_7024,N_7800);
or U8592 (N_8592,N_7992,N_7875);
nand U8593 (N_8593,N_7546,N_7488);
nor U8594 (N_8594,N_7398,N_7220);
xor U8595 (N_8595,N_7515,N_7283);
or U8596 (N_8596,N_7524,N_7496);
or U8597 (N_8597,N_7059,N_7218);
or U8598 (N_8598,N_7985,N_7271);
or U8599 (N_8599,N_7883,N_7810);
or U8600 (N_8600,N_7266,N_7247);
or U8601 (N_8601,N_7168,N_7374);
or U8602 (N_8602,N_7020,N_7723);
or U8603 (N_8603,N_7520,N_7215);
xor U8604 (N_8604,N_7176,N_7869);
nor U8605 (N_8605,N_7948,N_7113);
nand U8606 (N_8606,N_7219,N_7385);
and U8607 (N_8607,N_7090,N_7059);
nand U8608 (N_8608,N_7063,N_7804);
nand U8609 (N_8609,N_7497,N_7950);
and U8610 (N_8610,N_7588,N_7236);
nor U8611 (N_8611,N_7331,N_7302);
and U8612 (N_8612,N_7564,N_7071);
nor U8613 (N_8613,N_7683,N_7112);
and U8614 (N_8614,N_7049,N_7095);
nor U8615 (N_8615,N_7015,N_7877);
and U8616 (N_8616,N_7789,N_7674);
xnor U8617 (N_8617,N_7718,N_7906);
and U8618 (N_8618,N_7994,N_7974);
xnor U8619 (N_8619,N_7710,N_7464);
nand U8620 (N_8620,N_7077,N_7198);
and U8621 (N_8621,N_7102,N_7427);
or U8622 (N_8622,N_7573,N_7475);
nand U8623 (N_8623,N_7809,N_7989);
xor U8624 (N_8624,N_7804,N_7592);
or U8625 (N_8625,N_7606,N_7414);
xor U8626 (N_8626,N_7743,N_7963);
or U8627 (N_8627,N_7005,N_7263);
nand U8628 (N_8628,N_7639,N_7774);
xnor U8629 (N_8629,N_7478,N_7334);
xnor U8630 (N_8630,N_7093,N_7712);
and U8631 (N_8631,N_7282,N_7877);
and U8632 (N_8632,N_7893,N_7435);
and U8633 (N_8633,N_7918,N_7838);
nor U8634 (N_8634,N_7911,N_7638);
xnor U8635 (N_8635,N_7304,N_7055);
and U8636 (N_8636,N_7535,N_7053);
or U8637 (N_8637,N_7687,N_7108);
or U8638 (N_8638,N_7913,N_7460);
or U8639 (N_8639,N_7538,N_7932);
and U8640 (N_8640,N_7006,N_7815);
nand U8641 (N_8641,N_7417,N_7505);
xnor U8642 (N_8642,N_7322,N_7589);
and U8643 (N_8643,N_7555,N_7907);
nand U8644 (N_8644,N_7789,N_7821);
nand U8645 (N_8645,N_7172,N_7695);
nand U8646 (N_8646,N_7126,N_7835);
or U8647 (N_8647,N_7717,N_7816);
xnor U8648 (N_8648,N_7734,N_7930);
nor U8649 (N_8649,N_7008,N_7904);
nor U8650 (N_8650,N_7156,N_7830);
nand U8651 (N_8651,N_7757,N_7431);
nand U8652 (N_8652,N_7710,N_7371);
nor U8653 (N_8653,N_7241,N_7129);
xnor U8654 (N_8654,N_7840,N_7153);
nor U8655 (N_8655,N_7062,N_7782);
or U8656 (N_8656,N_7316,N_7889);
xor U8657 (N_8657,N_7642,N_7528);
and U8658 (N_8658,N_7031,N_7350);
and U8659 (N_8659,N_7175,N_7154);
nand U8660 (N_8660,N_7027,N_7687);
or U8661 (N_8661,N_7038,N_7301);
nand U8662 (N_8662,N_7954,N_7973);
nor U8663 (N_8663,N_7233,N_7742);
nor U8664 (N_8664,N_7609,N_7886);
nor U8665 (N_8665,N_7709,N_7772);
xor U8666 (N_8666,N_7100,N_7148);
xnor U8667 (N_8667,N_7258,N_7335);
or U8668 (N_8668,N_7414,N_7392);
nor U8669 (N_8669,N_7627,N_7744);
or U8670 (N_8670,N_7282,N_7291);
or U8671 (N_8671,N_7491,N_7711);
nand U8672 (N_8672,N_7112,N_7758);
nand U8673 (N_8673,N_7246,N_7700);
or U8674 (N_8674,N_7585,N_7763);
or U8675 (N_8675,N_7433,N_7789);
xor U8676 (N_8676,N_7236,N_7762);
and U8677 (N_8677,N_7044,N_7278);
and U8678 (N_8678,N_7538,N_7710);
nand U8679 (N_8679,N_7149,N_7231);
nand U8680 (N_8680,N_7418,N_7824);
xnor U8681 (N_8681,N_7457,N_7063);
and U8682 (N_8682,N_7308,N_7205);
or U8683 (N_8683,N_7575,N_7352);
nand U8684 (N_8684,N_7146,N_7578);
and U8685 (N_8685,N_7299,N_7732);
nor U8686 (N_8686,N_7420,N_7403);
nor U8687 (N_8687,N_7176,N_7962);
nand U8688 (N_8688,N_7981,N_7324);
or U8689 (N_8689,N_7884,N_7721);
nor U8690 (N_8690,N_7026,N_7930);
nand U8691 (N_8691,N_7756,N_7502);
nand U8692 (N_8692,N_7849,N_7701);
nor U8693 (N_8693,N_7414,N_7165);
and U8694 (N_8694,N_7951,N_7468);
and U8695 (N_8695,N_7312,N_7281);
and U8696 (N_8696,N_7571,N_7450);
and U8697 (N_8697,N_7803,N_7077);
nand U8698 (N_8698,N_7282,N_7520);
nand U8699 (N_8699,N_7129,N_7271);
and U8700 (N_8700,N_7674,N_7287);
or U8701 (N_8701,N_7695,N_7333);
nor U8702 (N_8702,N_7244,N_7698);
xor U8703 (N_8703,N_7100,N_7212);
nor U8704 (N_8704,N_7954,N_7710);
nand U8705 (N_8705,N_7523,N_7956);
nand U8706 (N_8706,N_7442,N_7381);
nor U8707 (N_8707,N_7668,N_7609);
xor U8708 (N_8708,N_7013,N_7749);
nand U8709 (N_8709,N_7304,N_7499);
xor U8710 (N_8710,N_7170,N_7816);
or U8711 (N_8711,N_7376,N_7849);
nand U8712 (N_8712,N_7202,N_7811);
or U8713 (N_8713,N_7509,N_7700);
nand U8714 (N_8714,N_7117,N_7470);
and U8715 (N_8715,N_7725,N_7938);
and U8716 (N_8716,N_7114,N_7150);
nand U8717 (N_8717,N_7878,N_7725);
and U8718 (N_8718,N_7747,N_7860);
and U8719 (N_8719,N_7392,N_7922);
xor U8720 (N_8720,N_7402,N_7806);
xnor U8721 (N_8721,N_7296,N_7082);
xnor U8722 (N_8722,N_7749,N_7328);
nand U8723 (N_8723,N_7027,N_7526);
nand U8724 (N_8724,N_7214,N_7958);
nand U8725 (N_8725,N_7831,N_7002);
nor U8726 (N_8726,N_7113,N_7806);
xor U8727 (N_8727,N_7788,N_7014);
or U8728 (N_8728,N_7273,N_7702);
or U8729 (N_8729,N_7869,N_7763);
nor U8730 (N_8730,N_7454,N_7368);
or U8731 (N_8731,N_7927,N_7897);
nand U8732 (N_8732,N_7969,N_7204);
and U8733 (N_8733,N_7237,N_7123);
and U8734 (N_8734,N_7438,N_7282);
xnor U8735 (N_8735,N_7353,N_7486);
nor U8736 (N_8736,N_7041,N_7841);
xor U8737 (N_8737,N_7364,N_7149);
nor U8738 (N_8738,N_7812,N_7393);
nand U8739 (N_8739,N_7614,N_7926);
nand U8740 (N_8740,N_7133,N_7444);
nand U8741 (N_8741,N_7751,N_7308);
nor U8742 (N_8742,N_7121,N_7441);
nand U8743 (N_8743,N_7868,N_7555);
xnor U8744 (N_8744,N_7962,N_7250);
nor U8745 (N_8745,N_7173,N_7146);
xor U8746 (N_8746,N_7397,N_7673);
xor U8747 (N_8747,N_7924,N_7115);
and U8748 (N_8748,N_7644,N_7530);
and U8749 (N_8749,N_7915,N_7782);
and U8750 (N_8750,N_7548,N_7572);
nor U8751 (N_8751,N_7972,N_7046);
nand U8752 (N_8752,N_7474,N_7625);
nand U8753 (N_8753,N_7051,N_7610);
nand U8754 (N_8754,N_7448,N_7213);
or U8755 (N_8755,N_7554,N_7212);
and U8756 (N_8756,N_7501,N_7321);
nor U8757 (N_8757,N_7472,N_7254);
or U8758 (N_8758,N_7355,N_7850);
nand U8759 (N_8759,N_7518,N_7736);
nor U8760 (N_8760,N_7571,N_7797);
and U8761 (N_8761,N_7279,N_7319);
and U8762 (N_8762,N_7752,N_7149);
nor U8763 (N_8763,N_7489,N_7298);
nor U8764 (N_8764,N_7925,N_7619);
and U8765 (N_8765,N_7087,N_7448);
xnor U8766 (N_8766,N_7135,N_7146);
and U8767 (N_8767,N_7740,N_7106);
and U8768 (N_8768,N_7505,N_7919);
nor U8769 (N_8769,N_7974,N_7473);
xnor U8770 (N_8770,N_7882,N_7501);
xor U8771 (N_8771,N_7992,N_7519);
or U8772 (N_8772,N_7100,N_7863);
and U8773 (N_8773,N_7606,N_7743);
and U8774 (N_8774,N_7026,N_7966);
or U8775 (N_8775,N_7144,N_7172);
and U8776 (N_8776,N_7761,N_7270);
nor U8777 (N_8777,N_7951,N_7404);
nand U8778 (N_8778,N_7749,N_7044);
nand U8779 (N_8779,N_7061,N_7507);
or U8780 (N_8780,N_7588,N_7088);
nor U8781 (N_8781,N_7475,N_7146);
and U8782 (N_8782,N_7127,N_7999);
and U8783 (N_8783,N_7951,N_7471);
nand U8784 (N_8784,N_7257,N_7003);
nor U8785 (N_8785,N_7400,N_7037);
nor U8786 (N_8786,N_7011,N_7485);
or U8787 (N_8787,N_7648,N_7117);
xnor U8788 (N_8788,N_7373,N_7948);
nand U8789 (N_8789,N_7682,N_7155);
or U8790 (N_8790,N_7148,N_7692);
and U8791 (N_8791,N_7904,N_7990);
nor U8792 (N_8792,N_7189,N_7233);
or U8793 (N_8793,N_7278,N_7180);
or U8794 (N_8794,N_7092,N_7581);
nand U8795 (N_8795,N_7119,N_7713);
nor U8796 (N_8796,N_7150,N_7442);
xnor U8797 (N_8797,N_7799,N_7311);
or U8798 (N_8798,N_7772,N_7830);
or U8799 (N_8799,N_7784,N_7699);
and U8800 (N_8800,N_7269,N_7790);
or U8801 (N_8801,N_7638,N_7632);
xnor U8802 (N_8802,N_7375,N_7540);
xor U8803 (N_8803,N_7298,N_7267);
xor U8804 (N_8804,N_7292,N_7403);
xnor U8805 (N_8805,N_7260,N_7264);
and U8806 (N_8806,N_7210,N_7924);
nand U8807 (N_8807,N_7345,N_7488);
nor U8808 (N_8808,N_7126,N_7584);
or U8809 (N_8809,N_7623,N_7931);
nor U8810 (N_8810,N_7662,N_7432);
xor U8811 (N_8811,N_7702,N_7215);
and U8812 (N_8812,N_7040,N_7445);
or U8813 (N_8813,N_7979,N_7045);
nand U8814 (N_8814,N_7480,N_7165);
nor U8815 (N_8815,N_7577,N_7687);
xnor U8816 (N_8816,N_7905,N_7269);
and U8817 (N_8817,N_7205,N_7103);
or U8818 (N_8818,N_7446,N_7028);
nor U8819 (N_8819,N_7280,N_7673);
xnor U8820 (N_8820,N_7714,N_7193);
nand U8821 (N_8821,N_7485,N_7466);
nor U8822 (N_8822,N_7646,N_7759);
or U8823 (N_8823,N_7990,N_7115);
or U8824 (N_8824,N_7370,N_7133);
nand U8825 (N_8825,N_7938,N_7808);
nand U8826 (N_8826,N_7541,N_7486);
nand U8827 (N_8827,N_7079,N_7750);
nand U8828 (N_8828,N_7907,N_7374);
nor U8829 (N_8829,N_7352,N_7690);
xor U8830 (N_8830,N_7355,N_7230);
nor U8831 (N_8831,N_7033,N_7184);
nor U8832 (N_8832,N_7948,N_7979);
nor U8833 (N_8833,N_7778,N_7461);
and U8834 (N_8834,N_7155,N_7150);
nor U8835 (N_8835,N_7537,N_7823);
and U8836 (N_8836,N_7767,N_7939);
and U8837 (N_8837,N_7862,N_7724);
or U8838 (N_8838,N_7896,N_7458);
or U8839 (N_8839,N_7112,N_7145);
nand U8840 (N_8840,N_7647,N_7325);
nor U8841 (N_8841,N_7097,N_7942);
and U8842 (N_8842,N_7556,N_7460);
and U8843 (N_8843,N_7192,N_7797);
and U8844 (N_8844,N_7877,N_7978);
nor U8845 (N_8845,N_7205,N_7373);
xor U8846 (N_8846,N_7175,N_7749);
xnor U8847 (N_8847,N_7768,N_7394);
xnor U8848 (N_8848,N_7717,N_7780);
nor U8849 (N_8849,N_7928,N_7178);
nor U8850 (N_8850,N_7523,N_7068);
or U8851 (N_8851,N_7461,N_7833);
and U8852 (N_8852,N_7074,N_7805);
nand U8853 (N_8853,N_7549,N_7999);
nor U8854 (N_8854,N_7541,N_7967);
nand U8855 (N_8855,N_7434,N_7352);
xnor U8856 (N_8856,N_7207,N_7482);
and U8857 (N_8857,N_7582,N_7079);
or U8858 (N_8858,N_7061,N_7730);
xnor U8859 (N_8859,N_7483,N_7274);
or U8860 (N_8860,N_7945,N_7967);
or U8861 (N_8861,N_7762,N_7427);
nand U8862 (N_8862,N_7425,N_7066);
or U8863 (N_8863,N_7520,N_7905);
and U8864 (N_8864,N_7890,N_7018);
nor U8865 (N_8865,N_7677,N_7930);
nand U8866 (N_8866,N_7425,N_7119);
nor U8867 (N_8867,N_7101,N_7673);
and U8868 (N_8868,N_7697,N_7465);
xor U8869 (N_8869,N_7008,N_7093);
or U8870 (N_8870,N_7111,N_7298);
or U8871 (N_8871,N_7536,N_7927);
nor U8872 (N_8872,N_7947,N_7923);
or U8873 (N_8873,N_7733,N_7807);
xnor U8874 (N_8874,N_7697,N_7143);
xor U8875 (N_8875,N_7675,N_7578);
nor U8876 (N_8876,N_7766,N_7818);
xnor U8877 (N_8877,N_7956,N_7886);
or U8878 (N_8878,N_7433,N_7005);
or U8879 (N_8879,N_7695,N_7619);
and U8880 (N_8880,N_7542,N_7575);
or U8881 (N_8881,N_7847,N_7459);
and U8882 (N_8882,N_7558,N_7181);
or U8883 (N_8883,N_7204,N_7853);
nor U8884 (N_8884,N_7290,N_7936);
or U8885 (N_8885,N_7937,N_7404);
and U8886 (N_8886,N_7318,N_7207);
nor U8887 (N_8887,N_7642,N_7645);
and U8888 (N_8888,N_7219,N_7418);
and U8889 (N_8889,N_7747,N_7490);
nor U8890 (N_8890,N_7069,N_7127);
or U8891 (N_8891,N_7566,N_7577);
and U8892 (N_8892,N_7529,N_7681);
and U8893 (N_8893,N_7306,N_7283);
nand U8894 (N_8894,N_7339,N_7100);
xor U8895 (N_8895,N_7309,N_7938);
and U8896 (N_8896,N_7741,N_7094);
or U8897 (N_8897,N_7259,N_7006);
nor U8898 (N_8898,N_7141,N_7968);
nor U8899 (N_8899,N_7142,N_7826);
nand U8900 (N_8900,N_7098,N_7765);
and U8901 (N_8901,N_7324,N_7532);
xor U8902 (N_8902,N_7085,N_7511);
nand U8903 (N_8903,N_7084,N_7372);
or U8904 (N_8904,N_7234,N_7921);
nand U8905 (N_8905,N_7799,N_7231);
and U8906 (N_8906,N_7300,N_7992);
xor U8907 (N_8907,N_7271,N_7237);
nor U8908 (N_8908,N_7785,N_7393);
or U8909 (N_8909,N_7837,N_7324);
xnor U8910 (N_8910,N_7128,N_7122);
nand U8911 (N_8911,N_7229,N_7605);
xor U8912 (N_8912,N_7285,N_7160);
nor U8913 (N_8913,N_7176,N_7291);
xnor U8914 (N_8914,N_7017,N_7830);
nor U8915 (N_8915,N_7074,N_7511);
and U8916 (N_8916,N_7359,N_7718);
and U8917 (N_8917,N_7100,N_7460);
or U8918 (N_8918,N_7660,N_7408);
or U8919 (N_8919,N_7224,N_7802);
or U8920 (N_8920,N_7405,N_7699);
and U8921 (N_8921,N_7933,N_7718);
or U8922 (N_8922,N_7877,N_7145);
nand U8923 (N_8923,N_7082,N_7314);
and U8924 (N_8924,N_7544,N_7174);
nor U8925 (N_8925,N_7493,N_7495);
nand U8926 (N_8926,N_7773,N_7118);
xor U8927 (N_8927,N_7812,N_7922);
nor U8928 (N_8928,N_7272,N_7294);
or U8929 (N_8929,N_7258,N_7894);
and U8930 (N_8930,N_7430,N_7169);
nor U8931 (N_8931,N_7689,N_7335);
nor U8932 (N_8932,N_7682,N_7288);
xnor U8933 (N_8933,N_7864,N_7457);
nor U8934 (N_8934,N_7400,N_7760);
and U8935 (N_8935,N_7849,N_7147);
or U8936 (N_8936,N_7640,N_7507);
xor U8937 (N_8937,N_7853,N_7703);
nand U8938 (N_8938,N_7641,N_7130);
nor U8939 (N_8939,N_7749,N_7702);
or U8940 (N_8940,N_7590,N_7614);
nor U8941 (N_8941,N_7931,N_7082);
nor U8942 (N_8942,N_7358,N_7872);
or U8943 (N_8943,N_7883,N_7375);
xor U8944 (N_8944,N_7974,N_7198);
or U8945 (N_8945,N_7552,N_7752);
and U8946 (N_8946,N_7148,N_7199);
nor U8947 (N_8947,N_7865,N_7376);
nor U8948 (N_8948,N_7552,N_7828);
nor U8949 (N_8949,N_7995,N_7335);
nand U8950 (N_8950,N_7792,N_7640);
nor U8951 (N_8951,N_7721,N_7195);
and U8952 (N_8952,N_7429,N_7146);
nor U8953 (N_8953,N_7686,N_7295);
or U8954 (N_8954,N_7612,N_7556);
and U8955 (N_8955,N_7929,N_7219);
nand U8956 (N_8956,N_7218,N_7717);
xor U8957 (N_8957,N_7541,N_7564);
nand U8958 (N_8958,N_7476,N_7510);
or U8959 (N_8959,N_7294,N_7461);
nand U8960 (N_8960,N_7006,N_7896);
nor U8961 (N_8961,N_7673,N_7017);
nor U8962 (N_8962,N_7440,N_7851);
and U8963 (N_8963,N_7202,N_7978);
or U8964 (N_8964,N_7680,N_7376);
nand U8965 (N_8965,N_7280,N_7521);
nor U8966 (N_8966,N_7096,N_7668);
and U8967 (N_8967,N_7166,N_7888);
xnor U8968 (N_8968,N_7716,N_7912);
or U8969 (N_8969,N_7170,N_7218);
or U8970 (N_8970,N_7742,N_7783);
and U8971 (N_8971,N_7368,N_7223);
or U8972 (N_8972,N_7506,N_7006);
nor U8973 (N_8973,N_7295,N_7276);
nor U8974 (N_8974,N_7042,N_7383);
or U8975 (N_8975,N_7773,N_7385);
nand U8976 (N_8976,N_7797,N_7351);
nand U8977 (N_8977,N_7387,N_7841);
and U8978 (N_8978,N_7806,N_7253);
or U8979 (N_8979,N_7486,N_7001);
and U8980 (N_8980,N_7077,N_7423);
nand U8981 (N_8981,N_7658,N_7654);
nand U8982 (N_8982,N_7725,N_7850);
and U8983 (N_8983,N_7091,N_7911);
nand U8984 (N_8984,N_7037,N_7899);
xnor U8985 (N_8985,N_7091,N_7310);
and U8986 (N_8986,N_7789,N_7166);
xnor U8987 (N_8987,N_7761,N_7806);
nor U8988 (N_8988,N_7491,N_7614);
or U8989 (N_8989,N_7729,N_7022);
nand U8990 (N_8990,N_7074,N_7629);
or U8991 (N_8991,N_7661,N_7238);
and U8992 (N_8992,N_7348,N_7488);
and U8993 (N_8993,N_7073,N_7982);
or U8994 (N_8994,N_7686,N_7018);
and U8995 (N_8995,N_7773,N_7398);
nand U8996 (N_8996,N_7906,N_7186);
or U8997 (N_8997,N_7714,N_7772);
nor U8998 (N_8998,N_7893,N_7654);
nand U8999 (N_8999,N_7404,N_7686);
xor U9000 (N_9000,N_8749,N_8358);
nor U9001 (N_9001,N_8039,N_8559);
or U9002 (N_9002,N_8769,N_8154);
nor U9003 (N_9003,N_8227,N_8915);
nor U9004 (N_9004,N_8340,N_8804);
and U9005 (N_9005,N_8996,N_8320);
nor U9006 (N_9006,N_8888,N_8676);
nand U9007 (N_9007,N_8525,N_8818);
xnor U9008 (N_9008,N_8071,N_8902);
xor U9009 (N_9009,N_8314,N_8136);
or U9010 (N_9010,N_8206,N_8354);
or U9011 (N_9011,N_8838,N_8107);
nand U9012 (N_9012,N_8569,N_8268);
nand U9013 (N_9013,N_8950,N_8586);
xnor U9014 (N_9014,N_8020,N_8670);
and U9015 (N_9015,N_8775,N_8948);
xor U9016 (N_9016,N_8587,N_8351);
xor U9017 (N_9017,N_8372,N_8729);
nor U9018 (N_9018,N_8700,N_8390);
or U9019 (N_9019,N_8632,N_8829);
xor U9020 (N_9020,N_8188,N_8633);
nand U9021 (N_9021,N_8190,N_8487);
or U9022 (N_9022,N_8044,N_8345);
nor U9023 (N_9023,N_8475,N_8477);
or U9024 (N_9024,N_8271,N_8016);
and U9025 (N_9025,N_8877,N_8984);
nand U9026 (N_9026,N_8885,N_8090);
and U9027 (N_9027,N_8100,N_8725);
xor U9028 (N_9028,N_8341,N_8108);
or U9029 (N_9029,N_8863,N_8373);
nand U9030 (N_9030,N_8425,N_8874);
xnor U9031 (N_9031,N_8097,N_8741);
or U9032 (N_9032,N_8618,N_8195);
and U9033 (N_9033,N_8791,N_8716);
nor U9034 (N_9034,N_8520,N_8544);
nor U9035 (N_9035,N_8878,N_8258);
or U9036 (N_9036,N_8147,N_8795);
and U9037 (N_9037,N_8709,N_8472);
and U9038 (N_9038,N_8199,N_8106);
xor U9039 (N_9039,N_8457,N_8708);
nand U9040 (N_9040,N_8453,N_8078);
and U9041 (N_9041,N_8242,N_8703);
or U9042 (N_9042,N_8507,N_8463);
nor U9043 (N_9043,N_8880,N_8419);
nor U9044 (N_9044,N_8380,N_8076);
xor U9045 (N_9045,N_8062,N_8461);
or U9046 (N_9046,N_8796,N_8201);
nand U9047 (N_9047,N_8790,N_8920);
nand U9048 (N_9048,N_8285,N_8315);
and U9049 (N_9049,N_8068,N_8157);
or U9050 (N_9050,N_8640,N_8911);
nor U9051 (N_9051,N_8261,N_8712);
and U9052 (N_9052,N_8462,N_8596);
xnor U9053 (N_9053,N_8698,N_8327);
and U9054 (N_9054,N_8947,N_8269);
nor U9055 (N_9055,N_8223,N_8822);
and U9056 (N_9056,N_8163,N_8659);
nor U9057 (N_9057,N_8115,N_8850);
nor U9058 (N_9058,N_8655,N_8980);
xnor U9059 (N_9059,N_8251,N_8089);
nor U9060 (N_9060,N_8515,N_8627);
xnor U9061 (N_9061,N_8392,N_8176);
and U9062 (N_9062,N_8502,N_8134);
and U9063 (N_9063,N_8198,N_8921);
nand U9064 (N_9064,N_8324,N_8069);
nor U9065 (N_9065,N_8526,N_8254);
nor U9066 (N_9066,N_8871,N_8932);
and U9067 (N_9067,N_8244,N_8181);
and U9068 (N_9068,N_8866,N_8672);
and U9069 (N_9069,N_8303,N_8930);
nor U9070 (N_9070,N_8872,N_8585);
and U9071 (N_9071,N_8479,N_8843);
and U9072 (N_9072,N_8070,N_8521);
and U9073 (N_9073,N_8578,N_8879);
nand U9074 (N_9074,N_8504,N_8143);
nor U9075 (N_9075,N_8631,N_8896);
xor U9076 (N_9076,N_8971,N_8421);
or U9077 (N_9077,N_8382,N_8882);
and U9078 (N_9078,N_8156,N_8292);
nor U9079 (N_9079,N_8000,N_8167);
nor U9080 (N_9080,N_8174,N_8083);
and U9081 (N_9081,N_8486,N_8404);
or U9082 (N_9082,N_8464,N_8045);
nor U9083 (N_9083,N_8812,N_8450);
and U9084 (N_9084,N_8636,N_8634);
nor U9085 (N_9085,N_8954,N_8538);
or U9086 (N_9086,N_8349,N_8770);
and U9087 (N_9087,N_8056,N_8756);
xnor U9088 (N_9088,N_8279,N_8801);
nor U9089 (N_9089,N_8609,N_8600);
nor U9090 (N_9090,N_8074,N_8131);
and U9091 (N_9091,N_8798,N_8958);
nor U9092 (N_9092,N_8498,N_8931);
and U9093 (N_9093,N_8506,N_8033);
or U9094 (N_9094,N_8029,N_8666);
and U9095 (N_9095,N_8912,N_8855);
and U9096 (N_9096,N_8316,N_8620);
or U9097 (N_9097,N_8658,N_8510);
and U9098 (N_9098,N_8063,N_8644);
xnor U9099 (N_9099,N_8519,N_8683);
xnor U9100 (N_9100,N_8706,N_8953);
nor U9101 (N_9101,N_8438,N_8601);
nand U9102 (N_9102,N_8868,N_8318);
and U9103 (N_9103,N_8326,N_8170);
and U9104 (N_9104,N_8629,N_8217);
nand U9105 (N_9105,N_8821,N_8919);
and U9106 (N_9106,N_8084,N_8649);
nand U9107 (N_9107,N_8577,N_8312);
xnor U9108 (N_9108,N_8323,N_8993);
and U9109 (N_9109,N_8375,N_8021);
and U9110 (N_9110,N_8210,N_8650);
xor U9111 (N_9111,N_8886,N_8053);
nand U9112 (N_9112,N_8619,N_8806);
or U9113 (N_9113,N_8309,N_8148);
xor U9114 (N_9114,N_8707,N_8408);
xnor U9115 (N_9115,N_8119,N_8359);
nor U9116 (N_9116,N_8196,N_8305);
nor U9117 (N_9117,N_8848,N_8881);
or U9118 (N_9118,N_8325,N_8155);
nand U9119 (N_9119,N_8678,N_8208);
or U9120 (N_9120,N_8200,N_8398);
and U9121 (N_9121,N_8718,N_8793);
nor U9122 (N_9122,N_8903,N_8471);
or U9123 (N_9123,N_8965,N_8307);
nor U9124 (N_9124,N_8481,N_8876);
or U9125 (N_9125,N_8832,N_8939);
nand U9126 (N_9126,N_8048,N_8681);
and U9127 (N_9127,N_8151,N_8745);
xor U9128 (N_9128,N_8413,N_8861);
nand U9129 (N_9129,N_8371,N_8758);
xor U9130 (N_9130,N_8165,N_8820);
nand U9131 (N_9131,N_8152,N_8067);
and U9132 (N_9132,N_8374,N_8897);
and U9133 (N_9133,N_8197,N_8228);
xor U9134 (N_9134,N_8643,N_8957);
nand U9135 (N_9135,N_8802,N_8813);
xnor U9136 (N_9136,N_8356,N_8355);
and U9137 (N_9137,N_8466,N_8517);
nand U9138 (N_9138,N_8081,N_8815);
and U9139 (N_9139,N_8563,N_8918);
or U9140 (N_9140,N_8975,N_8570);
nand U9141 (N_9141,N_8986,N_8998);
xnor U9142 (N_9142,N_8997,N_8335);
nand U9143 (N_9143,N_8465,N_8669);
or U9144 (N_9144,N_8590,N_8144);
and U9145 (N_9145,N_8289,N_8192);
or U9146 (N_9146,N_8782,N_8059);
or U9147 (N_9147,N_8027,N_8916);
xnor U9148 (N_9148,N_8278,N_8352);
and U9149 (N_9149,N_8330,N_8595);
nand U9150 (N_9150,N_8639,N_8853);
nand U9151 (N_9151,N_8524,N_8265);
nor U9152 (N_9152,N_8647,N_8982);
nor U9153 (N_9153,N_8873,N_8015);
or U9154 (N_9154,N_8987,N_8474);
nor U9155 (N_9155,N_8290,N_8075);
or U9156 (N_9156,N_8778,N_8363);
and U9157 (N_9157,N_8834,N_8328);
or U9158 (N_9158,N_8693,N_8929);
or U9159 (N_9159,N_8364,N_8792);
xor U9160 (N_9160,N_8414,N_8938);
nor U9161 (N_9161,N_8789,N_8742);
nand U9162 (N_9162,N_8146,N_8728);
nand U9163 (N_9163,N_8469,N_8376);
and U9164 (N_9164,N_8257,N_8281);
xnor U9165 (N_9165,N_8941,N_8560);
or U9166 (N_9166,N_8934,N_8186);
or U9167 (N_9167,N_8914,N_8434);
or U9168 (N_9168,N_8766,N_8495);
and U9169 (N_9169,N_8406,N_8130);
xnor U9170 (N_9170,N_8024,N_8992);
and U9171 (N_9171,N_8777,N_8999);
or U9172 (N_9172,N_8488,N_8531);
and U9173 (N_9173,N_8169,N_8500);
nand U9174 (N_9174,N_8420,N_8182);
nand U9175 (N_9175,N_8851,N_8910);
nand U9176 (N_9176,N_8150,N_8191);
nor U9177 (N_9177,N_8605,N_8123);
and U9178 (N_9178,N_8177,N_8956);
xor U9179 (N_9179,N_8091,N_8173);
nor U9180 (N_9180,N_8162,N_8933);
xnor U9181 (N_9181,N_8936,N_8602);
and U9182 (N_9182,N_8142,N_8411);
xor U9183 (N_9183,N_8892,N_8572);
nand U9184 (N_9184,N_8967,N_8779);
or U9185 (N_9185,N_8294,N_8653);
or U9186 (N_9186,N_8960,N_8484);
or U9187 (N_9187,N_8113,N_8386);
nand U9188 (N_9188,N_8125,N_8811);
nor U9189 (N_9189,N_8194,N_8893);
xor U9190 (N_9190,N_8651,N_8460);
or U9191 (N_9191,N_8109,N_8094);
nor U9192 (N_9192,N_8754,N_8935);
nor U9193 (N_9193,N_8383,N_8396);
and U9194 (N_9194,N_8235,N_8161);
nor U9195 (N_9195,N_8704,N_8731);
and U9196 (N_9196,N_8035,N_8267);
or U9197 (N_9197,N_8503,N_8567);
xor U9198 (N_9198,N_8682,N_8207);
nor U9199 (N_9199,N_8767,N_8166);
nor U9200 (N_9200,N_8193,N_8579);
nor U9201 (N_9201,N_8830,N_8613);
nand U9202 (N_9202,N_8378,N_8837);
nand U9203 (N_9203,N_8010,N_8737);
xnor U9204 (N_9204,N_8615,N_8339);
xor U9205 (N_9205,N_8007,N_8751);
nor U9206 (N_9206,N_8849,N_8665);
nand U9207 (N_9207,N_8606,N_8357);
or U9208 (N_9208,N_8895,N_8518);
nand U9209 (N_9209,N_8253,N_8485);
xnor U9210 (N_9210,N_8883,N_8072);
or U9211 (N_9211,N_8275,N_8141);
and U9212 (N_9212,N_8720,N_8400);
and U9213 (N_9213,N_8446,N_8299);
or U9214 (N_9214,N_8429,N_8512);
and U9215 (N_9215,N_8430,N_8394);
xor U9216 (N_9216,N_8426,N_8274);
nand U9217 (N_9217,N_8928,N_8179);
nand U9218 (N_9218,N_8648,N_8448);
nand U9219 (N_9219,N_8654,N_8291);
nand U9220 (N_9220,N_8841,N_8573);
nand U9221 (N_9221,N_8963,N_8001);
or U9222 (N_9222,N_8540,N_8370);
nor U9223 (N_9223,N_8679,N_8132);
nor U9224 (N_9224,N_8329,N_8722);
and U9225 (N_9225,N_8765,N_8610);
or U9226 (N_9226,N_8533,N_8857);
or U9227 (N_9227,N_8505,N_8427);
or U9228 (N_9228,N_8331,N_8899);
or U9229 (N_9229,N_8865,N_8974);
nand U9230 (N_9230,N_8819,N_8839);
nand U9231 (N_9231,N_8835,N_8065);
nand U9232 (N_9232,N_8828,N_8733);
or U9233 (N_9233,N_8388,N_8313);
xnor U9234 (N_9234,N_8671,N_8213);
and U9235 (N_9235,N_8012,N_8250);
or U9236 (N_9236,N_8657,N_8031);
nor U9237 (N_9237,N_8041,N_8444);
xnor U9238 (N_9238,N_8991,N_8407);
nor U9239 (N_9239,N_8183,N_8805);
nor U9240 (N_9240,N_8379,N_8467);
or U9241 (N_9241,N_8476,N_8255);
xor U9242 (N_9242,N_8638,N_8645);
and U9243 (N_9243,N_8454,N_8771);
nor U9244 (N_9244,N_8635,N_8551);
nor U9245 (N_9245,N_8064,N_8402);
nand U9246 (N_9246,N_8624,N_8087);
or U9247 (N_9247,N_8825,N_8491);
and U9248 (N_9248,N_8277,N_8616);
nand U9249 (N_9249,N_8565,N_8297);
nor U9250 (N_9250,N_8675,N_8336);
and U9251 (N_9251,N_8013,N_8715);
nand U9252 (N_9252,N_8478,N_8831);
nand U9253 (N_9253,N_8705,N_8922);
nand U9254 (N_9254,N_8668,N_8901);
and U9255 (N_9255,N_8387,N_8546);
nand U9256 (N_9256,N_8232,N_8612);
xor U9257 (N_9257,N_8234,N_8350);
nor U9258 (N_9258,N_8322,N_8236);
and U9259 (N_9259,N_8968,N_8311);
and U9260 (N_9260,N_8342,N_8810);
xor U9261 (N_9261,N_8739,N_8529);
and U9262 (N_9262,N_8721,N_8032);
and U9263 (N_9263,N_8717,N_8926);
nand U9264 (N_9264,N_8237,N_8497);
or U9265 (N_9265,N_8799,N_8293);
nand U9266 (N_9266,N_8367,N_8774);
nor U9267 (N_9267,N_8833,N_8827);
nor U9268 (N_9268,N_8262,N_8284);
nor U9269 (N_9269,N_8989,N_8036);
nand U9270 (N_9270,N_8889,N_8412);
xnor U9271 (N_9271,N_8913,N_8684);
nor U9272 (N_9272,N_8549,N_8691);
and U9273 (N_9273,N_8231,N_8887);
and U9274 (N_9274,N_8661,N_8149);
nor U9275 (N_9275,N_8875,N_8040);
xnor U9276 (N_9276,N_8058,N_8937);
xor U9277 (N_9277,N_8437,N_8384);
nor U9278 (N_9278,N_8334,N_8599);
xor U9279 (N_9279,N_8547,N_8701);
nand U9280 (N_9280,N_8270,N_8713);
and U9281 (N_9281,N_8447,N_8694);
xnor U9282 (N_9282,N_8302,N_8160);
xor U9283 (N_9283,N_8869,N_8854);
and U9284 (N_9284,N_8983,N_8088);
and U9285 (N_9285,N_8574,N_8321);
nor U9286 (N_9286,N_8308,N_8050);
and U9287 (N_9287,N_8501,N_8126);
nand U9288 (N_9288,N_8688,N_8272);
xnor U9289 (N_9289,N_8459,N_8099);
xnor U9290 (N_9290,N_8891,N_8924);
and U9291 (N_9291,N_8702,N_8019);
xor U9292 (N_9292,N_8159,N_8852);
and U9293 (N_9293,N_8381,N_8051);
nor U9294 (N_9294,N_8757,N_8976);
nor U9295 (N_9295,N_8391,N_8660);
xor U9296 (N_9296,N_8844,N_8224);
and U9297 (N_9297,N_8139,N_8562);
nand U9298 (N_9298,N_8823,N_8256);
nor U9299 (N_9299,N_8583,N_8296);
xnor U9300 (N_9300,N_8410,N_8499);
or U9301 (N_9301,N_8603,N_8755);
nand U9302 (N_9302,N_8780,N_8180);
or U9303 (N_9303,N_8752,N_8537);
nor U9304 (N_9304,N_8952,N_8128);
nand U9305 (N_9305,N_8856,N_8338);
xor U9306 (N_9306,N_8994,N_8319);
or U9307 (N_9307,N_8121,N_8061);
and U9308 (N_9308,N_8608,N_8022);
xnor U9309 (N_9309,N_8047,N_8079);
or U9310 (N_9310,N_8859,N_8216);
xor U9311 (N_9311,N_8252,N_8046);
nor U9312 (N_9312,N_8105,N_8781);
xnor U9313 (N_9313,N_8532,N_8263);
and U9314 (N_9314,N_8158,N_8699);
nand U9315 (N_9315,N_8772,N_8202);
or U9316 (N_9316,N_8824,N_8168);
nand U9317 (N_9317,N_8642,N_8346);
and U9318 (N_9318,N_8301,N_8424);
xnor U9319 (N_9319,N_8558,N_8037);
nor U9320 (N_9320,N_8028,N_8052);
and U9321 (N_9321,N_8451,N_8656);
nand U9322 (N_9322,N_8489,N_8995);
and U9323 (N_9323,N_8175,N_8748);
nor U9324 (N_9324,N_8082,N_8576);
and U9325 (N_9325,N_8542,N_8692);
nand U9326 (N_9326,N_8203,N_8005);
nand U9327 (N_9327,N_8862,N_8621);
or U9328 (N_9328,N_8724,N_8422);
xnor U9329 (N_9329,N_8456,N_8184);
nor U9330 (N_9330,N_8554,N_8528);
and U9331 (N_9331,N_8164,N_8840);
or U9332 (N_9332,N_8439,N_8759);
or U9333 (N_9333,N_8347,N_8055);
nand U9334 (N_9334,N_8496,N_8522);
nand U9335 (N_9335,N_8979,N_8401);
or U9336 (N_9336,N_8295,N_8222);
or U9337 (N_9337,N_8727,N_8317);
or U9338 (N_9338,N_8580,N_8575);
nor U9339 (N_9339,N_8508,N_8397);
and U9340 (N_9340,N_8416,N_8807);
nand U9341 (N_9341,N_8240,N_8153);
nand U9342 (N_9342,N_8761,N_8393);
xnor U9343 (N_9343,N_8981,N_8816);
and U9344 (N_9344,N_8204,N_8847);
xnor U9345 (N_9345,N_8137,N_8923);
xor U9346 (N_9346,N_8768,N_8259);
or U9347 (N_9347,N_8836,N_8095);
or U9348 (N_9348,N_8940,N_8455);
and U9349 (N_9349,N_8470,N_8212);
and U9350 (N_9350,N_8011,N_8622);
and U9351 (N_9351,N_8276,N_8905);
nor U9352 (N_9352,N_8145,N_8185);
or U9353 (N_9353,N_8740,N_8025);
xnor U9354 (N_9354,N_8955,N_8788);
xnor U9355 (N_9355,N_8114,N_8049);
xor U9356 (N_9356,N_8054,N_8568);
or U9357 (N_9357,N_8445,N_8909);
nor U9358 (N_9358,N_8431,N_8626);
and U9359 (N_9359,N_8399,N_8589);
xnor U9360 (N_9360,N_8026,N_8409);
nor U9361 (N_9361,N_8490,N_8764);
and U9362 (N_9362,N_8135,N_8870);
nand U9363 (N_9363,N_8978,N_8405);
nor U9364 (N_9364,N_8440,N_8743);
xnor U9365 (N_9365,N_8432,N_8593);
nor U9366 (N_9366,N_8218,N_8803);
nand U9367 (N_9367,N_8673,N_8494);
or U9368 (N_9368,N_8264,N_8073);
nand U9369 (N_9369,N_8030,N_8417);
or U9370 (N_9370,N_8038,N_8365);
or U9371 (N_9371,N_8187,N_8561);
and U9372 (N_9372,N_8077,N_8710);
or U9373 (N_9373,N_8233,N_8617);
nand U9374 (N_9374,N_8248,N_8864);
nor U9375 (N_9375,N_8369,N_8867);
and U9376 (N_9376,N_8990,N_8286);
and U9377 (N_9377,N_8641,N_8687);
or U9378 (N_9378,N_8066,N_8908);
or U9379 (N_9379,N_8623,N_8110);
xnor U9380 (N_9380,N_8680,N_8101);
nor U9381 (N_9381,N_8564,N_8458);
nor U9382 (N_9382,N_8723,N_8966);
and U9383 (N_9383,N_8898,N_8808);
nand U9384 (N_9384,N_8884,N_8018);
nand U9385 (N_9385,N_8760,N_8773);
and U9386 (N_9386,N_8189,N_8220);
xnor U9387 (N_9387,N_8415,N_8353);
nor U9388 (N_9388,N_8961,N_8423);
or U9389 (N_9389,N_8085,N_8753);
and U9390 (N_9390,N_8776,N_8266);
xnor U9391 (N_9391,N_8535,N_8973);
nand U9392 (N_9392,N_8566,N_8003);
nor U9393 (N_9393,N_8628,N_8133);
or U9394 (N_9394,N_8238,N_8418);
xnor U9395 (N_9395,N_8098,N_8797);
and U9396 (N_9396,N_8273,N_8241);
xnor U9397 (N_9397,N_8553,N_8591);
xor U9398 (N_9398,N_8625,N_8845);
nand U9399 (N_9399,N_8043,N_8171);
xor U9400 (N_9400,N_8280,N_8366);
and U9401 (N_9401,N_8215,N_8962);
nand U9402 (N_9402,N_8906,N_8536);
or U9403 (N_9403,N_8900,N_8787);
nand U9404 (N_9404,N_8664,N_8786);
nor U9405 (N_9405,N_8102,N_8118);
xnor U9406 (N_9406,N_8588,N_8744);
or U9407 (N_9407,N_8817,N_8763);
or U9408 (N_9408,N_8719,N_8970);
xnor U9409 (N_9409,N_8907,N_8172);
xor U9410 (N_9410,N_8221,N_8557);
xnor U9411 (N_9411,N_8904,N_8738);
nand U9412 (N_9412,N_8057,N_8300);
xor U9413 (N_9413,N_8129,N_8034);
or U9414 (N_9414,N_8138,N_8695);
and U9415 (N_9415,N_8677,N_8543);
xnor U9416 (N_9416,N_8604,N_8730);
and U9417 (N_9417,N_8945,N_8361);
or U9418 (N_9418,N_8711,N_8385);
or U9419 (N_9419,N_8433,N_8306);
or U9420 (N_9420,N_8229,N_8571);
and U9421 (N_9421,N_8493,N_8685);
nand U9422 (N_9422,N_8686,N_8959);
nor U9423 (N_9423,N_8548,N_8735);
nor U9424 (N_9424,N_8607,N_8023);
nand U9425 (N_9425,N_8435,N_8584);
nand U9426 (N_9426,N_8014,N_8509);
xnor U9427 (N_9427,N_8714,N_8927);
and U9428 (N_9428,N_8246,N_8667);
or U9429 (N_9429,N_8545,N_8245);
or U9430 (N_9430,N_8377,N_8582);
nand U9431 (N_9431,N_8287,N_8332);
and U9432 (N_9432,N_8794,N_8942);
or U9433 (N_9433,N_8663,N_8750);
nand U9434 (N_9434,N_8288,N_8178);
xnor U9435 (N_9435,N_8112,N_8482);
and U9436 (N_9436,N_8951,N_8513);
and U9437 (N_9437,N_8211,N_8225);
xor U9438 (N_9438,N_8826,N_8511);
nand U9439 (N_9439,N_8646,N_8080);
or U9440 (N_9440,N_8890,N_8747);
or U9441 (N_9441,N_8348,N_8483);
nand U9442 (N_9442,N_8333,N_8337);
nor U9443 (N_9443,N_8117,N_8697);
xnor U9444 (N_9444,N_8611,N_8592);
or U9445 (N_9445,N_8949,N_8403);
nand U9446 (N_9446,N_8310,N_8304);
nor U9447 (N_9447,N_8527,N_8004);
nand U9448 (N_9448,N_8539,N_8726);
nand U9449 (N_9449,N_8614,N_8002);
and U9450 (N_9450,N_8516,N_8783);
or U9451 (N_9451,N_8598,N_8042);
nor U9452 (N_9452,N_8111,N_8534);
or U9453 (N_9453,N_8243,N_8096);
or U9454 (N_9454,N_8086,N_8917);
xor U9455 (N_9455,N_8449,N_8122);
xnor U9456 (N_9456,N_8226,N_8630);
nor U9457 (N_9457,N_8556,N_8637);
or U9458 (N_9458,N_8943,N_8282);
nand U9459 (N_9459,N_8452,N_8581);
and U9460 (N_9460,N_8597,N_8977);
xnor U9461 (N_9461,N_8674,N_8436);
nor U9462 (N_9462,N_8480,N_8140);
xor U9463 (N_9463,N_8925,N_8814);
or U9464 (N_9464,N_8230,N_8652);
nand U9465 (N_9465,N_8944,N_8127);
xnor U9466 (N_9466,N_8809,N_8008);
xnor U9467 (N_9467,N_8492,N_8442);
xor U9468 (N_9468,N_8732,N_8060);
nand U9469 (N_9469,N_8468,N_8969);
nand U9470 (N_9470,N_8552,N_8009);
nor U9471 (N_9471,N_8784,N_8785);
xor U9472 (N_9472,N_8092,N_8360);
nor U9473 (N_9473,N_8964,N_8858);
or U9474 (N_9474,N_8988,N_8103);
and U9475 (N_9475,N_8734,N_8736);
and U9476 (N_9476,N_8846,N_8124);
xor U9477 (N_9477,N_8260,N_8443);
or U9478 (N_9478,N_8116,N_8219);
or U9479 (N_9479,N_8441,N_8550);
nand U9480 (N_9480,N_8017,N_8239);
xnor U9481 (N_9481,N_8594,N_8205);
nand U9482 (N_9482,N_8690,N_8104);
xor U9483 (N_9483,N_8762,N_8249);
xor U9484 (N_9484,N_8283,N_8214);
nor U9485 (N_9485,N_8946,N_8696);
or U9486 (N_9486,N_8746,N_8473);
xnor U9487 (N_9487,N_8972,N_8541);
nor U9488 (N_9488,N_8247,N_8800);
nand U9489 (N_9489,N_8555,N_8662);
nand U9490 (N_9490,N_8344,N_8368);
nand U9491 (N_9491,N_8298,N_8389);
nor U9492 (N_9492,N_8006,N_8395);
nor U9493 (N_9493,N_8523,N_8120);
nor U9494 (N_9494,N_8842,N_8093);
nor U9495 (N_9495,N_8530,N_8514);
or U9496 (N_9496,N_8428,N_8894);
or U9497 (N_9497,N_8860,N_8689);
nand U9498 (N_9498,N_8985,N_8209);
nor U9499 (N_9499,N_8362,N_8343);
xnor U9500 (N_9500,N_8137,N_8982);
nor U9501 (N_9501,N_8281,N_8189);
or U9502 (N_9502,N_8710,N_8066);
nand U9503 (N_9503,N_8702,N_8557);
or U9504 (N_9504,N_8351,N_8231);
nand U9505 (N_9505,N_8337,N_8402);
or U9506 (N_9506,N_8112,N_8996);
or U9507 (N_9507,N_8309,N_8779);
and U9508 (N_9508,N_8338,N_8357);
and U9509 (N_9509,N_8942,N_8763);
and U9510 (N_9510,N_8034,N_8989);
and U9511 (N_9511,N_8683,N_8076);
xor U9512 (N_9512,N_8791,N_8660);
xnor U9513 (N_9513,N_8813,N_8071);
xnor U9514 (N_9514,N_8051,N_8926);
nor U9515 (N_9515,N_8967,N_8349);
nand U9516 (N_9516,N_8920,N_8396);
nor U9517 (N_9517,N_8648,N_8695);
nand U9518 (N_9518,N_8709,N_8681);
nor U9519 (N_9519,N_8534,N_8632);
or U9520 (N_9520,N_8418,N_8375);
nor U9521 (N_9521,N_8994,N_8700);
or U9522 (N_9522,N_8246,N_8189);
or U9523 (N_9523,N_8006,N_8857);
xor U9524 (N_9524,N_8093,N_8614);
or U9525 (N_9525,N_8655,N_8354);
or U9526 (N_9526,N_8075,N_8115);
and U9527 (N_9527,N_8665,N_8568);
nor U9528 (N_9528,N_8210,N_8755);
nand U9529 (N_9529,N_8287,N_8971);
xor U9530 (N_9530,N_8843,N_8834);
xnor U9531 (N_9531,N_8175,N_8002);
and U9532 (N_9532,N_8866,N_8825);
or U9533 (N_9533,N_8442,N_8449);
or U9534 (N_9534,N_8898,N_8111);
nor U9535 (N_9535,N_8820,N_8722);
nor U9536 (N_9536,N_8637,N_8163);
nand U9537 (N_9537,N_8158,N_8127);
nand U9538 (N_9538,N_8830,N_8851);
or U9539 (N_9539,N_8050,N_8743);
or U9540 (N_9540,N_8611,N_8478);
xor U9541 (N_9541,N_8606,N_8327);
or U9542 (N_9542,N_8216,N_8567);
and U9543 (N_9543,N_8244,N_8380);
nor U9544 (N_9544,N_8315,N_8655);
and U9545 (N_9545,N_8778,N_8957);
nor U9546 (N_9546,N_8294,N_8572);
xnor U9547 (N_9547,N_8953,N_8928);
nand U9548 (N_9548,N_8376,N_8228);
or U9549 (N_9549,N_8998,N_8109);
and U9550 (N_9550,N_8932,N_8708);
and U9551 (N_9551,N_8875,N_8254);
xor U9552 (N_9552,N_8063,N_8990);
and U9553 (N_9553,N_8004,N_8473);
or U9554 (N_9554,N_8549,N_8353);
xor U9555 (N_9555,N_8833,N_8424);
nand U9556 (N_9556,N_8308,N_8514);
nand U9557 (N_9557,N_8540,N_8934);
and U9558 (N_9558,N_8515,N_8761);
and U9559 (N_9559,N_8358,N_8312);
nor U9560 (N_9560,N_8147,N_8334);
nor U9561 (N_9561,N_8199,N_8507);
nor U9562 (N_9562,N_8220,N_8088);
nor U9563 (N_9563,N_8002,N_8904);
and U9564 (N_9564,N_8606,N_8334);
nand U9565 (N_9565,N_8857,N_8431);
xnor U9566 (N_9566,N_8788,N_8633);
and U9567 (N_9567,N_8326,N_8057);
and U9568 (N_9568,N_8162,N_8127);
xor U9569 (N_9569,N_8137,N_8983);
and U9570 (N_9570,N_8112,N_8024);
and U9571 (N_9571,N_8031,N_8894);
nor U9572 (N_9572,N_8816,N_8349);
nand U9573 (N_9573,N_8010,N_8144);
xor U9574 (N_9574,N_8140,N_8255);
nand U9575 (N_9575,N_8055,N_8960);
or U9576 (N_9576,N_8992,N_8920);
nand U9577 (N_9577,N_8944,N_8756);
and U9578 (N_9578,N_8900,N_8004);
and U9579 (N_9579,N_8610,N_8464);
and U9580 (N_9580,N_8827,N_8043);
nand U9581 (N_9581,N_8901,N_8174);
or U9582 (N_9582,N_8325,N_8746);
and U9583 (N_9583,N_8769,N_8725);
or U9584 (N_9584,N_8506,N_8642);
nand U9585 (N_9585,N_8489,N_8018);
nand U9586 (N_9586,N_8896,N_8646);
and U9587 (N_9587,N_8936,N_8383);
nor U9588 (N_9588,N_8447,N_8796);
xnor U9589 (N_9589,N_8021,N_8436);
or U9590 (N_9590,N_8533,N_8983);
and U9591 (N_9591,N_8913,N_8355);
or U9592 (N_9592,N_8634,N_8016);
nor U9593 (N_9593,N_8538,N_8076);
nor U9594 (N_9594,N_8253,N_8358);
or U9595 (N_9595,N_8599,N_8632);
and U9596 (N_9596,N_8019,N_8293);
xnor U9597 (N_9597,N_8831,N_8745);
nand U9598 (N_9598,N_8177,N_8235);
or U9599 (N_9599,N_8939,N_8427);
xor U9600 (N_9600,N_8319,N_8264);
nand U9601 (N_9601,N_8797,N_8444);
and U9602 (N_9602,N_8695,N_8692);
nor U9603 (N_9603,N_8876,N_8077);
or U9604 (N_9604,N_8569,N_8079);
and U9605 (N_9605,N_8520,N_8139);
nor U9606 (N_9606,N_8285,N_8337);
nor U9607 (N_9607,N_8859,N_8404);
nor U9608 (N_9608,N_8797,N_8057);
xnor U9609 (N_9609,N_8058,N_8392);
nor U9610 (N_9610,N_8622,N_8349);
or U9611 (N_9611,N_8659,N_8452);
or U9612 (N_9612,N_8528,N_8832);
and U9613 (N_9613,N_8274,N_8658);
or U9614 (N_9614,N_8853,N_8732);
xnor U9615 (N_9615,N_8861,N_8633);
nor U9616 (N_9616,N_8272,N_8918);
nor U9617 (N_9617,N_8728,N_8295);
or U9618 (N_9618,N_8062,N_8356);
nand U9619 (N_9619,N_8601,N_8626);
xnor U9620 (N_9620,N_8323,N_8752);
xor U9621 (N_9621,N_8351,N_8278);
and U9622 (N_9622,N_8433,N_8864);
and U9623 (N_9623,N_8054,N_8497);
or U9624 (N_9624,N_8269,N_8061);
nand U9625 (N_9625,N_8380,N_8479);
or U9626 (N_9626,N_8126,N_8803);
and U9627 (N_9627,N_8800,N_8307);
or U9628 (N_9628,N_8197,N_8641);
nand U9629 (N_9629,N_8915,N_8997);
nor U9630 (N_9630,N_8804,N_8849);
or U9631 (N_9631,N_8094,N_8415);
xor U9632 (N_9632,N_8232,N_8069);
or U9633 (N_9633,N_8676,N_8236);
nor U9634 (N_9634,N_8731,N_8186);
nand U9635 (N_9635,N_8672,N_8934);
xor U9636 (N_9636,N_8940,N_8913);
or U9637 (N_9637,N_8720,N_8194);
or U9638 (N_9638,N_8477,N_8110);
xor U9639 (N_9639,N_8747,N_8675);
and U9640 (N_9640,N_8303,N_8712);
and U9641 (N_9641,N_8037,N_8883);
nor U9642 (N_9642,N_8513,N_8070);
xnor U9643 (N_9643,N_8914,N_8592);
xor U9644 (N_9644,N_8196,N_8588);
nand U9645 (N_9645,N_8532,N_8740);
or U9646 (N_9646,N_8785,N_8683);
nand U9647 (N_9647,N_8303,N_8996);
xnor U9648 (N_9648,N_8893,N_8269);
xor U9649 (N_9649,N_8769,N_8569);
or U9650 (N_9650,N_8342,N_8749);
nand U9651 (N_9651,N_8157,N_8856);
nand U9652 (N_9652,N_8862,N_8915);
or U9653 (N_9653,N_8984,N_8252);
and U9654 (N_9654,N_8989,N_8349);
nand U9655 (N_9655,N_8763,N_8649);
nor U9656 (N_9656,N_8568,N_8827);
nor U9657 (N_9657,N_8717,N_8985);
or U9658 (N_9658,N_8679,N_8280);
and U9659 (N_9659,N_8991,N_8118);
or U9660 (N_9660,N_8063,N_8855);
xnor U9661 (N_9661,N_8786,N_8253);
nor U9662 (N_9662,N_8300,N_8086);
xor U9663 (N_9663,N_8686,N_8038);
xor U9664 (N_9664,N_8942,N_8800);
nand U9665 (N_9665,N_8166,N_8736);
xnor U9666 (N_9666,N_8266,N_8747);
and U9667 (N_9667,N_8624,N_8931);
and U9668 (N_9668,N_8792,N_8712);
and U9669 (N_9669,N_8039,N_8099);
or U9670 (N_9670,N_8303,N_8741);
xor U9671 (N_9671,N_8589,N_8033);
or U9672 (N_9672,N_8343,N_8613);
xnor U9673 (N_9673,N_8839,N_8621);
and U9674 (N_9674,N_8764,N_8923);
or U9675 (N_9675,N_8083,N_8418);
and U9676 (N_9676,N_8282,N_8140);
nand U9677 (N_9677,N_8922,N_8051);
nor U9678 (N_9678,N_8533,N_8232);
nand U9679 (N_9679,N_8917,N_8808);
nor U9680 (N_9680,N_8738,N_8235);
and U9681 (N_9681,N_8172,N_8879);
nand U9682 (N_9682,N_8298,N_8803);
and U9683 (N_9683,N_8535,N_8514);
or U9684 (N_9684,N_8231,N_8716);
xor U9685 (N_9685,N_8543,N_8253);
xor U9686 (N_9686,N_8222,N_8442);
nand U9687 (N_9687,N_8562,N_8902);
and U9688 (N_9688,N_8904,N_8941);
nand U9689 (N_9689,N_8208,N_8655);
or U9690 (N_9690,N_8263,N_8635);
xor U9691 (N_9691,N_8785,N_8493);
nand U9692 (N_9692,N_8371,N_8181);
nand U9693 (N_9693,N_8827,N_8002);
and U9694 (N_9694,N_8700,N_8244);
and U9695 (N_9695,N_8682,N_8003);
xnor U9696 (N_9696,N_8142,N_8197);
xnor U9697 (N_9697,N_8769,N_8547);
nor U9698 (N_9698,N_8074,N_8521);
nand U9699 (N_9699,N_8236,N_8487);
xor U9700 (N_9700,N_8753,N_8951);
or U9701 (N_9701,N_8154,N_8705);
nor U9702 (N_9702,N_8040,N_8887);
or U9703 (N_9703,N_8327,N_8028);
nor U9704 (N_9704,N_8790,N_8101);
nand U9705 (N_9705,N_8199,N_8466);
nand U9706 (N_9706,N_8491,N_8069);
nor U9707 (N_9707,N_8141,N_8143);
xor U9708 (N_9708,N_8463,N_8157);
and U9709 (N_9709,N_8268,N_8382);
xnor U9710 (N_9710,N_8088,N_8770);
and U9711 (N_9711,N_8595,N_8304);
xor U9712 (N_9712,N_8829,N_8188);
xnor U9713 (N_9713,N_8088,N_8025);
nand U9714 (N_9714,N_8776,N_8766);
and U9715 (N_9715,N_8748,N_8491);
and U9716 (N_9716,N_8229,N_8845);
xnor U9717 (N_9717,N_8060,N_8404);
and U9718 (N_9718,N_8839,N_8476);
xor U9719 (N_9719,N_8230,N_8958);
and U9720 (N_9720,N_8912,N_8881);
xnor U9721 (N_9721,N_8553,N_8387);
nor U9722 (N_9722,N_8275,N_8352);
or U9723 (N_9723,N_8171,N_8656);
xor U9724 (N_9724,N_8341,N_8759);
and U9725 (N_9725,N_8845,N_8169);
nand U9726 (N_9726,N_8966,N_8732);
xor U9727 (N_9727,N_8857,N_8607);
xor U9728 (N_9728,N_8806,N_8564);
nor U9729 (N_9729,N_8152,N_8083);
xnor U9730 (N_9730,N_8291,N_8287);
and U9731 (N_9731,N_8877,N_8436);
and U9732 (N_9732,N_8836,N_8908);
nor U9733 (N_9733,N_8381,N_8316);
or U9734 (N_9734,N_8798,N_8292);
and U9735 (N_9735,N_8975,N_8362);
nor U9736 (N_9736,N_8540,N_8797);
nor U9737 (N_9737,N_8401,N_8945);
nor U9738 (N_9738,N_8509,N_8598);
xnor U9739 (N_9739,N_8981,N_8492);
or U9740 (N_9740,N_8776,N_8445);
and U9741 (N_9741,N_8229,N_8253);
nand U9742 (N_9742,N_8776,N_8466);
and U9743 (N_9743,N_8323,N_8045);
and U9744 (N_9744,N_8972,N_8594);
xor U9745 (N_9745,N_8169,N_8955);
nor U9746 (N_9746,N_8258,N_8221);
nand U9747 (N_9747,N_8313,N_8775);
and U9748 (N_9748,N_8703,N_8717);
xnor U9749 (N_9749,N_8017,N_8417);
nand U9750 (N_9750,N_8163,N_8886);
and U9751 (N_9751,N_8285,N_8830);
nand U9752 (N_9752,N_8310,N_8804);
and U9753 (N_9753,N_8617,N_8446);
nor U9754 (N_9754,N_8326,N_8690);
xor U9755 (N_9755,N_8915,N_8995);
xor U9756 (N_9756,N_8932,N_8219);
and U9757 (N_9757,N_8908,N_8941);
or U9758 (N_9758,N_8372,N_8918);
nand U9759 (N_9759,N_8625,N_8866);
nor U9760 (N_9760,N_8360,N_8616);
nor U9761 (N_9761,N_8232,N_8920);
nand U9762 (N_9762,N_8231,N_8721);
xnor U9763 (N_9763,N_8280,N_8413);
nor U9764 (N_9764,N_8724,N_8132);
nor U9765 (N_9765,N_8703,N_8017);
and U9766 (N_9766,N_8930,N_8244);
or U9767 (N_9767,N_8708,N_8337);
nor U9768 (N_9768,N_8256,N_8521);
or U9769 (N_9769,N_8233,N_8481);
and U9770 (N_9770,N_8121,N_8004);
nor U9771 (N_9771,N_8053,N_8320);
and U9772 (N_9772,N_8850,N_8312);
xor U9773 (N_9773,N_8798,N_8016);
nand U9774 (N_9774,N_8233,N_8645);
xor U9775 (N_9775,N_8623,N_8771);
nor U9776 (N_9776,N_8509,N_8234);
or U9777 (N_9777,N_8793,N_8995);
nor U9778 (N_9778,N_8812,N_8492);
xnor U9779 (N_9779,N_8439,N_8960);
xnor U9780 (N_9780,N_8232,N_8718);
and U9781 (N_9781,N_8397,N_8609);
and U9782 (N_9782,N_8365,N_8377);
and U9783 (N_9783,N_8269,N_8916);
xor U9784 (N_9784,N_8686,N_8404);
nor U9785 (N_9785,N_8493,N_8556);
or U9786 (N_9786,N_8488,N_8837);
nand U9787 (N_9787,N_8138,N_8858);
nor U9788 (N_9788,N_8547,N_8643);
nor U9789 (N_9789,N_8172,N_8388);
nor U9790 (N_9790,N_8022,N_8703);
nand U9791 (N_9791,N_8384,N_8271);
nand U9792 (N_9792,N_8305,N_8926);
xnor U9793 (N_9793,N_8337,N_8408);
nand U9794 (N_9794,N_8086,N_8152);
or U9795 (N_9795,N_8400,N_8950);
xor U9796 (N_9796,N_8968,N_8483);
nor U9797 (N_9797,N_8280,N_8704);
or U9798 (N_9798,N_8385,N_8853);
nor U9799 (N_9799,N_8265,N_8294);
and U9800 (N_9800,N_8679,N_8194);
xnor U9801 (N_9801,N_8416,N_8967);
and U9802 (N_9802,N_8741,N_8364);
xor U9803 (N_9803,N_8675,N_8652);
and U9804 (N_9804,N_8351,N_8834);
xor U9805 (N_9805,N_8452,N_8407);
and U9806 (N_9806,N_8894,N_8904);
and U9807 (N_9807,N_8259,N_8690);
or U9808 (N_9808,N_8462,N_8464);
nor U9809 (N_9809,N_8834,N_8551);
nor U9810 (N_9810,N_8253,N_8218);
nand U9811 (N_9811,N_8462,N_8148);
xor U9812 (N_9812,N_8074,N_8972);
nand U9813 (N_9813,N_8077,N_8990);
or U9814 (N_9814,N_8632,N_8479);
and U9815 (N_9815,N_8829,N_8473);
nor U9816 (N_9816,N_8004,N_8989);
nor U9817 (N_9817,N_8412,N_8843);
nor U9818 (N_9818,N_8236,N_8099);
nor U9819 (N_9819,N_8106,N_8624);
xnor U9820 (N_9820,N_8331,N_8976);
and U9821 (N_9821,N_8677,N_8100);
and U9822 (N_9822,N_8309,N_8506);
nor U9823 (N_9823,N_8980,N_8621);
or U9824 (N_9824,N_8578,N_8636);
nand U9825 (N_9825,N_8962,N_8854);
nor U9826 (N_9826,N_8361,N_8870);
or U9827 (N_9827,N_8015,N_8101);
or U9828 (N_9828,N_8191,N_8615);
and U9829 (N_9829,N_8900,N_8868);
and U9830 (N_9830,N_8506,N_8785);
nor U9831 (N_9831,N_8627,N_8601);
or U9832 (N_9832,N_8518,N_8419);
or U9833 (N_9833,N_8311,N_8180);
xnor U9834 (N_9834,N_8743,N_8830);
xnor U9835 (N_9835,N_8836,N_8463);
xnor U9836 (N_9836,N_8003,N_8757);
nor U9837 (N_9837,N_8431,N_8650);
and U9838 (N_9838,N_8658,N_8212);
xnor U9839 (N_9839,N_8571,N_8564);
nor U9840 (N_9840,N_8275,N_8570);
nand U9841 (N_9841,N_8007,N_8406);
nand U9842 (N_9842,N_8818,N_8402);
nor U9843 (N_9843,N_8476,N_8635);
and U9844 (N_9844,N_8787,N_8106);
or U9845 (N_9845,N_8287,N_8243);
xnor U9846 (N_9846,N_8015,N_8099);
or U9847 (N_9847,N_8853,N_8553);
nand U9848 (N_9848,N_8574,N_8567);
nand U9849 (N_9849,N_8184,N_8874);
nand U9850 (N_9850,N_8342,N_8157);
nand U9851 (N_9851,N_8109,N_8634);
or U9852 (N_9852,N_8738,N_8391);
nand U9853 (N_9853,N_8429,N_8275);
nand U9854 (N_9854,N_8758,N_8300);
nand U9855 (N_9855,N_8822,N_8766);
or U9856 (N_9856,N_8818,N_8309);
or U9857 (N_9857,N_8632,N_8984);
xnor U9858 (N_9858,N_8064,N_8183);
and U9859 (N_9859,N_8941,N_8019);
and U9860 (N_9860,N_8766,N_8080);
xor U9861 (N_9861,N_8347,N_8945);
nor U9862 (N_9862,N_8523,N_8945);
xor U9863 (N_9863,N_8210,N_8050);
and U9864 (N_9864,N_8316,N_8732);
and U9865 (N_9865,N_8092,N_8874);
nand U9866 (N_9866,N_8084,N_8469);
nand U9867 (N_9867,N_8818,N_8417);
or U9868 (N_9868,N_8312,N_8686);
or U9869 (N_9869,N_8785,N_8372);
nand U9870 (N_9870,N_8187,N_8227);
and U9871 (N_9871,N_8264,N_8642);
xor U9872 (N_9872,N_8081,N_8556);
and U9873 (N_9873,N_8523,N_8326);
and U9874 (N_9874,N_8895,N_8702);
nand U9875 (N_9875,N_8899,N_8021);
nand U9876 (N_9876,N_8869,N_8462);
nand U9877 (N_9877,N_8408,N_8945);
and U9878 (N_9878,N_8020,N_8409);
xor U9879 (N_9879,N_8759,N_8583);
or U9880 (N_9880,N_8303,N_8415);
and U9881 (N_9881,N_8015,N_8265);
and U9882 (N_9882,N_8588,N_8112);
or U9883 (N_9883,N_8236,N_8378);
nor U9884 (N_9884,N_8097,N_8337);
or U9885 (N_9885,N_8170,N_8244);
nand U9886 (N_9886,N_8787,N_8915);
nor U9887 (N_9887,N_8988,N_8800);
xnor U9888 (N_9888,N_8424,N_8942);
nand U9889 (N_9889,N_8469,N_8359);
or U9890 (N_9890,N_8731,N_8151);
nor U9891 (N_9891,N_8272,N_8588);
and U9892 (N_9892,N_8251,N_8199);
or U9893 (N_9893,N_8019,N_8189);
nor U9894 (N_9894,N_8644,N_8164);
xor U9895 (N_9895,N_8502,N_8557);
xnor U9896 (N_9896,N_8127,N_8438);
nand U9897 (N_9897,N_8038,N_8198);
nor U9898 (N_9898,N_8891,N_8441);
and U9899 (N_9899,N_8647,N_8418);
nor U9900 (N_9900,N_8880,N_8998);
xor U9901 (N_9901,N_8906,N_8853);
nor U9902 (N_9902,N_8911,N_8257);
and U9903 (N_9903,N_8155,N_8931);
nand U9904 (N_9904,N_8702,N_8161);
nand U9905 (N_9905,N_8051,N_8603);
and U9906 (N_9906,N_8925,N_8830);
nor U9907 (N_9907,N_8531,N_8959);
or U9908 (N_9908,N_8443,N_8810);
xor U9909 (N_9909,N_8097,N_8685);
nand U9910 (N_9910,N_8772,N_8044);
and U9911 (N_9911,N_8995,N_8674);
or U9912 (N_9912,N_8290,N_8708);
nor U9913 (N_9913,N_8302,N_8525);
nor U9914 (N_9914,N_8410,N_8947);
nand U9915 (N_9915,N_8715,N_8864);
nor U9916 (N_9916,N_8017,N_8618);
nor U9917 (N_9917,N_8870,N_8269);
or U9918 (N_9918,N_8879,N_8909);
xor U9919 (N_9919,N_8623,N_8958);
xor U9920 (N_9920,N_8673,N_8328);
or U9921 (N_9921,N_8267,N_8130);
and U9922 (N_9922,N_8213,N_8026);
xor U9923 (N_9923,N_8905,N_8790);
or U9924 (N_9924,N_8976,N_8222);
and U9925 (N_9925,N_8276,N_8350);
nor U9926 (N_9926,N_8874,N_8990);
nand U9927 (N_9927,N_8649,N_8500);
or U9928 (N_9928,N_8387,N_8256);
nand U9929 (N_9929,N_8041,N_8936);
nand U9930 (N_9930,N_8719,N_8714);
xor U9931 (N_9931,N_8239,N_8098);
or U9932 (N_9932,N_8795,N_8437);
or U9933 (N_9933,N_8274,N_8375);
and U9934 (N_9934,N_8851,N_8218);
nand U9935 (N_9935,N_8225,N_8687);
or U9936 (N_9936,N_8399,N_8354);
nand U9937 (N_9937,N_8293,N_8518);
xnor U9938 (N_9938,N_8750,N_8542);
or U9939 (N_9939,N_8890,N_8411);
nor U9940 (N_9940,N_8294,N_8371);
xor U9941 (N_9941,N_8674,N_8319);
and U9942 (N_9942,N_8105,N_8972);
xnor U9943 (N_9943,N_8065,N_8302);
xor U9944 (N_9944,N_8033,N_8694);
xor U9945 (N_9945,N_8362,N_8582);
and U9946 (N_9946,N_8948,N_8624);
and U9947 (N_9947,N_8655,N_8971);
nor U9948 (N_9948,N_8286,N_8290);
nand U9949 (N_9949,N_8963,N_8381);
xor U9950 (N_9950,N_8986,N_8127);
nor U9951 (N_9951,N_8262,N_8724);
nand U9952 (N_9952,N_8965,N_8009);
xnor U9953 (N_9953,N_8815,N_8485);
or U9954 (N_9954,N_8083,N_8044);
and U9955 (N_9955,N_8547,N_8937);
or U9956 (N_9956,N_8909,N_8793);
xor U9957 (N_9957,N_8622,N_8591);
nand U9958 (N_9958,N_8063,N_8882);
or U9959 (N_9959,N_8993,N_8176);
xor U9960 (N_9960,N_8110,N_8224);
xor U9961 (N_9961,N_8006,N_8495);
or U9962 (N_9962,N_8600,N_8744);
and U9963 (N_9963,N_8341,N_8006);
or U9964 (N_9964,N_8498,N_8358);
and U9965 (N_9965,N_8016,N_8024);
nand U9966 (N_9966,N_8524,N_8429);
xnor U9967 (N_9967,N_8037,N_8797);
and U9968 (N_9968,N_8144,N_8253);
nand U9969 (N_9969,N_8047,N_8736);
nor U9970 (N_9970,N_8645,N_8351);
nand U9971 (N_9971,N_8351,N_8325);
nor U9972 (N_9972,N_8513,N_8869);
nand U9973 (N_9973,N_8799,N_8041);
and U9974 (N_9974,N_8955,N_8775);
nor U9975 (N_9975,N_8922,N_8059);
xor U9976 (N_9976,N_8608,N_8493);
nand U9977 (N_9977,N_8654,N_8937);
nor U9978 (N_9978,N_8031,N_8471);
nor U9979 (N_9979,N_8195,N_8621);
and U9980 (N_9980,N_8214,N_8247);
and U9981 (N_9981,N_8603,N_8772);
nand U9982 (N_9982,N_8328,N_8768);
xnor U9983 (N_9983,N_8369,N_8356);
or U9984 (N_9984,N_8628,N_8324);
and U9985 (N_9985,N_8133,N_8501);
nand U9986 (N_9986,N_8889,N_8553);
nand U9987 (N_9987,N_8926,N_8053);
xnor U9988 (N_9988,N_8494,N_8256);
xnor U9989 (N_9989,N_8164,N_8280);
nand U9990 (N_9990,N_8899,N_8084);
nand U9991 (N_9991,N_8524,N_8994);
xnor U9992 (N_9992,N_8100,N_8198);
xor U9993 (N_9993,N_8741,N_8194);
or U9994 (N_9994,N_8487,N_8510);
and U9995 (N_9995,N_8274,N_8808);
xor U9996 (N_9996,N_8532,N_8568);
nor U9997 (N_9997,N_8378,N_8175);
and U9998 (N_9998,N_8716,N_8341);
nor U9999 (N_9999,N_8037,N_8084);
or U10000 (N_10000,N_9373,N_9291);
xnor U10001 (N_10001,N_9238,N_9931);
nand U10002 (N_10002,N_9885,N_9316);
or U10003 (N_10003,N_9494,N_9767);
nor U10004 (N_10004,N_9429,N_9173);
and U10005 (N_10005,N_9024,N_9439);
nor U10006 (N_10006,N_9865,N_9692);
nor U10007 (N_10007,N_9334,N_9691);
nand U10008 (N_10008,N_9405,N_9641);
xnor U10009 (N_10009,N_9739,N_9356);
and U10010 (N_10010,N_9218,N_9107);
nor U10011 (N_10011,N_9760,N_9999);
nor U10012 (N_10012,N_9797,N_9202);
xnor U10013 (N_10013,N_9050,N_9086);
nor U10014 (N_10014,N_9615,N_9069);
or U10015 (N_10015,N_9794,N_9390);
and U10016 (N_10016,N_9876,N_9526);
xor U10017 (N_10017,N_9795,N_9658);
xor U10018 (N_10018,N_9052,N_9700);
and U10019 (N_10019,N_9610,N_9905);
xor U10020 (N_10020,N_9210,N_9997);
and U10021 (N_10021,N_9869,N_9681);
or U10022 (N_10022,N_9828,N_9256);
nand U10023 (N_10023,N_9561,N_9467);
nor U10024 (N_10024,N_9542,N_9891);
xnor U10025 (N_10025,N_9490,N_9713);
nand U10026 (N_10026,N_9567,N_9226);
or U10027 (N_10027,N_9988,N_9991);
nor U10028 (N_10028,N_9637,N_9483);
and U10029 (N_10029,N_9604,N_9303);
xor U10030 (N_10030,N_9493,N_9234);
xor U10031 (N_10031,N_9856,N_9792);
nand U10032 (N_10032,N_9079,N_9450);
and U10033 (N_10033,N_9308,N_9621);
nor U10034 (N_10034,N_9309,N_9447);
and U10035 (N_10035,N_9881,N_9001);
or U10036 (N_10036,N_9694,N_9357);
nand U10037 (N_10037,N_9520,N_9258);
xor U10038 (N_10038,N_9227,N_9067);
and U10039 (N_10039,N_9082,N_9744);
or U10040 (N_10040,N_9386,N_9057);
nor U10041 (N_10041,N_9193,N_9593);
and U10042 (N_10042,N_9064,N_9034);
nand U10043 (N_10043,N_9338,N_9928);
and U10044 (N_10044,N_9573,N_9081);
and U10045 (N_10045,N_9867,N_9530);
xor U10046 (N_10046,N_9233,N_9804);
or U10047 (N_10047,N_9693,N_9206);
or U10048 (N_10048,N_9205,N_9484);
and U10049 (N_10049,N_9471,N_9720);
nor U10050 (N_10050,N_9640,N_9370);
or U10051 (N_10051,N_9848,N_9088);
nand U10052 (N_10052,N_9260,N_9464);
xnor U10053 (N_10053,N_9973,N_9643);
xor U10054 (N_10054,N_9457,N_9910);
and U10055 (N_10055,N_9400,N_9648);
nand U10056 (N_10056,N_9126,N_9280);
xor U10057 (N_10057,N_9441,N_9552);
and U10058 (N_10058,N_9159,N_9372);
xnor U10059 (N_10059,N_9476,N_9076);
nand U10060 (N_10060,N_9862,N_9754);
nand U10061 (N_10061,N_9903,N_9409);
nor U10062 (N_10062,N_9654,N_9055);
nand U10063 (N_10063,N_9111,N_9671);
nor U10064 (N_10064,N_9116,N_9385);
xor U10065 (N_10065,N_9866,N_9169);
nor U10066 (N_10066,N_9197,N_9897);
and U10067 (N_10067,N_9533,N_9304);
xnor U10068 (N_10068,N_9263,N_9004);
nor U10069 (N_10069,N_9732,N_9294);
and U10070 (N_10070,N_9051,N_9607);
nor U10071 (N_10071,N_9039,N_9564);
nor U10072 (N_10072,N_9266,N_9228);
nand U10073 (N_10073,N_9244,N_9300);
and U10074 (N_10074,N_9247,N_9054);
nand U10075 (N_10075,N_9305,N_9678);
and U10076 (N_10076,N_9726,N_9673);
nor U10077 (N_10077,N_9199,N_9670);
or U10078 (N_10078,N_9320,N_9783);
xnor U10079 (N_10079,N_9435,N_9524);
nand U10080 (N_10080,N_9818,N_9938);
xnor U10081 (N_10081,N_9463,N_9131);
or U10082 (N_10082,N_9666,N_9699);
and U10083 (N_10083,N_9185,N_9299);
and U10084 (N_10084,N_9874,N_9401);
nor U10085 (N_10085,N_9438,N_9838);
or U10086 (N_10086,N_9179,N_9870);
and U10087 (N_10087,N_9337,N_9675);
or U10088 (N_10088,N_9717,N_9295);
xnor U10089 (N_10089,N_9801,N_9889);
nor U10090 (N_10090,N_9198,N_9877);
and U10091 (N_10091,N_9029,N_9336);
or U10092 (N_10092,N_9736,N_9119);
nand U10093 (N_10093,N_9209,N_9926);
nand U10094 (N_10094,N_9620,N_9375);
and U10095 (N_10095,N_9721,N_9231);
xor U10096 (N_10096,N_9752,N_9301);
xor U10097 (N_10097,N_9410,N_9787);
nor U10098 (N_10098,N_9985,N_9940);
and U10099 (N_10099,N_9201,N_9384);
nor U10100 (N_10100,N_9239,N_9443);
nand U10101 (N_10101,N_9695,N_9200);
or U10102 (N_10102,N_9765,N_9243);
nor U10103 (N_10103,N_9017,N_9072);
or U10104 (N_10104,N_9237,N_9745);
or U10105 (N_10105,N_9106,N_9606);
nor U10106 (N_10106,N_9381,N_9275);
or U10107 (N_10107,N_9398,N_9759);
and U10108 (N_10108,N_9784,N_9424);
nor U10109 (N_10109,N_9909,N_9922);
and U10110 (N_10110,N_9407,N_9513);
nor U10111 (N_10111,N_9474,N_9556);
xnor U10112 (N_10112,N_9462,N_9093);
and U10113 (N_10113,N_9849,N_9269);
or U10114 (N_10114,N_9261,N_9432);
xnor U10115 (N_10115,N_9845,N_9329);
or U10116 (N_10116,N_9351,N_9078);
or U10117 (N_10117,N_9661,N_9453);
and U10118 (N_10118,N_9422,N_9125);
nand U10119 (N_10119,N_9104,N_9558);
or U10120 (N_10120,N_9177,N_9781);
nor U10121 (N_10121,N_9430,N_9684);
or U10122 (N_10122,N_9192,N_9006);
and U10123 (N_10123,N_9053,N_9742);
and U10124 (N_10124,N_9872,N_9811);
nor U10125 (N_10125,N_9598,N_9092);
nand U10126 (N_10126,N_9915,N_9639);
nand U10127 (N_10127,N_9049,N_9630);
and U10128 (N_10128,N_9778,N_9032);
nand U10129 (N_10129,N_9154,N_9182);
nand U10130 (N_10130,N_9954,N_9377);
or U10131 (N_10131,N_9124,N_9762);
nand U10132 (N_10132,N_9251,N_9584);
nand U10133 (N_10133,N_9028,N_9449);
nand U10134 (N_10134,N_9652,N_9802);
and U10135 (N_10135,N_9625,N_9293);
nand U10136 (N_10136,N_9286,N_9095);
or U10137 (N_10137,N_9901,N_9148);
or U10138 (N_10138,N_9688,N_9911);
or U10139 (N_10139,N_9701,N_9644);
and U10140 (N_10140,N_9216,N_9068);
or U10141 (N_10141,N_9623,N_9217);
xor U10142 (N_10142,N_9011,N_9091);
and U10143 (N_10143,N_9782,N_9576);
and U10144 (N_10144,N_9171,N_9989);
and U10145 (N_10145,N_9506,N_9097);
or U10146 (N_10146,N_9517,N_9510);
nor U10147 (N_10147,N_9757,N_9902);
or U10148 (N_10148,N_9307,N_9884);
nand U10149 (N_10149,N_9923,N_9735);
and U10150 (N_10150,N_9521,N_9037);
nand U10151 (N_10151,N_9033,N_9557);
nand U10152 (N_10152,N_9427,N_9488);
nand U10153 (N_10153,N_9824,N_9027);
and U10154 (N_10154,N_9858,N_9907);
and U10155 (N_10155,N_9821,N_9495);
or U10156 (N_10156,N_9588,N_9822);
or U10157 (N_10157,N_9916,N_9906);
nor U10158 (N_10158,N_9809,N_9519);
nor U10159 (N_10159,N_9737,N_9603);
xor U10160 (N_10160,N_9486,N_9344);
nor U10161 (N_10161,N_9974,N_9270);
xnor U10162 (N_10162,N_9135,N_9966);
nand U10163 (N_10163,N_9842,N_9761);
nand U10164 (N_10164,N_9843,N_9514);
nor U10165 (N_10165,N_9408,N_9340);
xnor U10166 (N_10166,N_9339,N_9317);
and U10167 (N_10167,N_9958,N_9235);
nor U10168 (N_10168,N_9361,N_9190);
nand U10169 (N_10169,N_9541,N_9302);
nor U10170 (N_10170,N_9707,N_9383);
and U10171 (N_10171,N_9937,N_9109);
and U10172 (N_10172,N_9272,N_9194);
or U10173 (N_10173,N_9609,N_9832);
and U10174 (N_10174,N_9850,N_9975);
or U10175 (N_10175,N_9946,N_9953);
or U10176 (N_10176,N_9016,N_9864);
nand U10177 (N_10177,N_9632,N_9428);
nand U10178 (N_10178,N_9914,N_9246);
nor U10179 (N_10179,N_9022,N_9245);
nand U10180 (N_10180,N_9306,N_9448);
or U10181 (N_10181,N_9793,N_9469);
and U10182 (N_10182,N_9638,N_9108);
nor U10183 (N_10183,N_9144,N_9477);
and U10184 (N_10184,N_9010,N_9747);
or U10185 (N_10185,N_9882,N_9536);
and U10186 (N_10186,N_9491,N_9933);
or U10187 (N_10187,N_9221,N_9013);
nor U10188 (N_10188,N_9844,N_9803);
or U10189 (N_10189,N_9583,N_9018);
or U10190 (N_10190,N_9129,N_9114);
or U10191 (N_10191,N_9267,N_9690);
xor U10192 (N_10192,N_9602,N_9712);
xor U10193 (N_10193,N_9616,N_9746);
xnor U10194 (N_10194,N_9330,N_9417);
nor U10195 (N_10195,N_9854,N_9825);
or U10196 (N_10196,N_9731,N_9359);
or U10197 (N_10197,N_9733,N_9472);
nor U10198 (N_10198,N_9976,N_9977);
nand U10199 (N_10199,N_9475,N_9364);
xnor U10200 (N_10200,N_9392,N_9815);
nor U10201 (N_10201,N_9133,N_9993);
or U10202 (N_10202,N_9855,N_9163);
nand U10203 (N_10203,N_9380,N_9348);
nor U10204 (N_10204,N_9478,N_9629);
xor U10205 (N_10205,N_9768,N_9503);
xnor U10206 (N_10206,N_9810,N_9662);
xor U10207 (N_10207,N_9705,N_9682);
nor U10208 (N_10208,N_9164,N_9137);
or U10209 (N_10209,N_9220,N_9442);
and U10210 (N_10210,N_9509,N_9113);
or U10211 (N_10211,N_9096,N_9539);
xnor U10212 (N_10212,N_9461,N_9618);
or U10213 (N_10213,N_9323,N_9659);
or U10214 (N_10214,N_9240,N_9635);
or U10215 (N_10215,N_9566,N_9956);
xnor U10216 (N_10216,N_9970,N_9951);
xnor U10217 (N_10217,N_9551,N_9389);
or U10218 (N_10218,N_9697,N_9020);
nor U10219 (N_10219,N_9987,N_9161);
nor U10220 (N_10220,N_9404,N_9813);
xor U10221 (N_10221,N_9395,N_9586);
nand U10222 (N_10222,N_9175,N_9957);
xor U10223 (N_10223,N_9741,N_9979);
xor U10224 (N_10224,N_9518,N_9262);
or U10225 (N_10225,N_9538,N_9574);
nand U10226 (N_10226,N_9722,N_9685);
nand U10227 (N_10227,N_9773,N_9667);
nor U10228 (N_10228,N_9780,N_9589);
nand U10229 (N_10229,N_9264,N_9590);
xnor U10230 (N_10230,N_9788,N_9656);
nand U10231 (N_10231,N_9689,N_9288);
nand U10232 (N_10232,N_9917,N_9531);
or U10233 (N_10233,N_9134,N_9799);
nand U10234 (N_10234,N_9073,N_9470);
xnor U10235 (N_10235,N_9204,N_9770);
nor U10236 (N_10236,N_9366,N_9995);
nor U10237 (N_10237,N_9327,N_9942);
or U10238 (N_10238,N_9485,N_9924);
xor U10239 (N_10239,N_9099,N_9645);
and U10240 (N_10240,N_9753,N_9600);
or U10241 (N_10241,N_9000,N_9203);
nor U10242 (N_10242,N_9649,N_9626);
nor U10243 (N_10243,N_9160,N_9873);
or U10244 (N_10244,N_9614,N_9687);
xor U10245 (N_10245,N_9172,N_9063);
nand U10246 (N_10246,N_9147,N_9298);
nand U10247 (N_10247,N_9962,N_9501);
nand U10248 (N_10248,N_9242,N_9894);
nor U10249 (N_10249,N_9335,N_9056);
or U10250 (N_10250,N_9837,N_9935);
nand U10251 (N_10251,N_9433,N_9676);
nor U10252 (N_10252,N_9343,N_9499);
nor U10253 (N_10253,N_9779,N_9756);
nor U10254 (N_10254,N_9543,N_9248);
xnor U10255 (N_10255,N_9080,N_9719);
nor U10256 (N_10256,N_9492,N_9898);
nand U10257 (N_10257,N_9311,N_9259);
xor U10258 (N_10258,N_9345,N_9886);
xnor U10259 (N_10259,N_9711,N_9515);
xnor U10260 (N_10260,N_9045,N_9893);
nor U10261 (N_10261,N_9165,N_9030);
and U10262 (N_10262,N_9347,N_9121);
and U10263 (N_10263,N_9504,N_9085);
and U10264 (N_10264,N_9149,N_9718);
or U10265 (N_10265,N_9419,N_9857);
or U10266 (N_10266,N_9315,N_9313);
nor U10267 (N_10267,N_9378,N_9101);
nand U10268 (N_10268,N_9679,N_9554);
nand U10269 (N_10269,N_9704,N_9749);
or U10270 (N_10270,N_9145,N_9505);
or U10271 (N_10271,N_9139,N_9672);
nor U10272 (N_10272,N_9727,N_9892);
or U10273 (N_10273,N_9277,N_9151);
or U10274 (N_10274,N_9814,N_9283);
nand U10275 (N_10275,N_9498,N_9015);
xor U10276 (N_10276,N_9599,N_9349);
and U10277 (N_10277,N_9657,N_9230);
xnor U10278 (N_10278,N_9900,N_9075);
nand U10279 (N_10279,N_9540,N_9066);
nor U10280 (N_10280,N_9391,N_9601);
nor U10281 (N_10281,N_9806,N_9785);
xor U10282 (N_10282,N_9978,N_9326);
xor U10283 (N_10283,N_9141,N_9211);
or U10284 (N_10284,N_9249,N_9547);
or U10285 (N_10285,N_9831,N_9367);
nor U10286 (N_10286,N_9038,N_9730);
or U10287 (N_10287,N_9331,N_9127);
and U10288 (N_10288,N_9094,N_9952);
xor U10289 (N_10289,N_9660,N_9103);
and U10290 (N_10290,N_9932,N_9333);
or U10291 (N_10291,N_9250,N_9612);
nand U10292 (N_10292,N_9466,N_9459);
and U10293 (N_10293,N_9580,N_9947);
nand U10294 (N_10294,N_9835,N_9955);
and U10295 (N_10295,N_9980,N_9964);
and U10296 (N_10296,N_9031,N_9310);
nor U10297 (N_10297,N_9553,N_9572);
nand U10298 (N_10298,N_9522,N_9983);
nand U10299 (N_10299,N_9142,N_9416);
or U10300 (N_10300,N_9534,N_9455);
nor U10301 (N_10301,N_9451,N_9456);
nand U10302 (N_10302,N_9512,N_9406);
xnor U10303 (N_10303,N_9930,N_9596);
or U10304 (N_10304,N_9847,N_9817);
or U10305 (N_10305,N_9986,N_9710);
or U10306 (N_10306,N_9423,N_9152);
nand U10307 (N_10307,N_9669,N_9665);
nand U10308 (N_10308,N_9290,N_9544);
and U10309 (N_10309,N_9786,N_9706);
nor U10310 (N_10310,N_9968,N_9841);
or U10311 (N_10311,N_9883,N_9215);
or U10312 (N_10312,N_9156,N_9362);
nor U10313 (N_10313,N_9895,N_9569);
or U10314 (N_10314,N_9207,N_9887);
and U10315 (N_10315,N_9703,N_9546);
nor U10316 (N_10316,N_9776,N_9436);
nor U10317 (N_10317,N_9943,N_9253);
and U10318 (N_10318,N_9140,N_9823);
nor U10319 (N_10319,N_9077,N_9166);
or U10320 (N_10320,N_9771,N_9473);
nor U10321 (N_10321,N_9425,N_9281);
xor U10322 (N_10322,N_9219,N_9899);
nand U10323 (N_10323,N_9002,N_9110);
xnor U10324 (N_10324,N_9146,N_9959);
and U10325 (N_10325,N_9545,N_9289);
nor U10326 (N_10326,N_9715,N_9322);
or U10327 (N_10327,N_9920,N_9945);
and U10328 (N_10328,N_9969,N_9388);
xor U10329 (N_10329,N_9664,N_9468);
nand U10330 (N_10330,N_9507,N_9851);
and U10331 (N_10331,N_9371,N_9826);
and U10332 (N_10332,N_9570,N_9830);
xnor U10333 (N_10333,N_9686,N_9296);
xor U10334 (N_10334,N_9846,N_9363);
nand U10335 (N_10335,N_9122,N_9724);
xor U10336 (N_10336,N_9071,N_9624);
and U10337 (N_10337,N_9655,N_9611);
nand U10338 (N_10338,N_9413,N_9585);
and U10339 (N_10339,N_9619,N_9668);
and U10340 (N_10340,N_9723,N_9994);
or U10341 (N_10341,N_9680,N_9229);
nor U10342 (N_10342,N_9941,N_9187);
xnor U10343 (N_10343,N_9734,N_9382);
or U10344 (N_10344,N_9790,N_9268);
nor U10345 (N_10345,N_9376,N_9508);
nand U10346 (N_10346,N_9496,N_9426);
xnor U10347 (N_10347,N_9368,N_9984);
nand U10348 (N_10348,N_9379,N_9083);
and U10349 (N_10349,N_9581,N_9170);
nor U10350 (N_10350,N_9683,N_9550);
xnor U10351 (N_10351,N_9112,N_9936);
nand U10352 (N_10352,N_9738,N_9729);
and U10353 (N_10353,N_9748,N_9403);
or U10354 (N_10354,N_9579,N_9992);
nand U10355 (N_10355,N_9186,N_9040);
xnor U10356 (N_10356,N_9279,N_9180);
nand U10357 (N_10357,N_9213,N_9879);
and U10358 (N_10358,N_9431,N_9608);
and U10359 (N_10359,N_9489,N_9816);
nor U10360 (N_10360,N_9025,N_9650);
nor U10361 (N_10361,N_9117,N_9374);
and U10362 (N_10362,N_9048,N_9089);
or U10363 (N_10363,N_9402,N_9312);
nand U10364 (N_10364,N_9653,N_9254);
nand U10365 (N_10365,N_9223,N_9829);
nor U10366 (N_10366,N_9714,N_9393);
xor U10367 (N_10367,N_9123,N_9440);
and U10368 (N_10368,N_9578,N_9257);
nor U10369 (N_10369,N_9224,N_9355);
and U10370 (N_10370,N_9852,N_9341);
and U10371 (N_10371,N_9225,N_9132);
and U10372 (N_10372,N_9274,N_9948);
or U10373 (N_10373,N_9434,N_9138);
or U10374 (N_10374,N_9528,N_9021);
nand U10375 (N_10375,N_9525,N_9549);
xnor U10376 (N_10376,N_9766,N_9325);
or U10377 (N_10377,N_9036,N_9919);
or U10378 (N_10378,N_9497,N_9728);
nor U10379 (N_10379,N_9314,N_9130);
and U10380 (N_10380,N_9062,N_9319);
xnor U10381 (N_10381,N_9880,N_9807);
nand U10382 (N_10382,N_9839,N_9888);
and U10383 (N_10383,N_9740,N_9005);
xnor U10384 (N_10384,N_9252,N_9763);
nand U10385 (N_10385,N_9421,N_9481);
xor U10386 (N_10386,N_9042,N_9044);
or U10387 (N_10387,N_9827,N_9871);
or U10388 (N_10388,N_9812,N_9796);
or U10389 (N_10389,N_9157,N_9232);
nand U10390 (N_10390,N_9353,N_9677);
and U10391 (N_10391,N_9155,N_9411);
or U10392 (N_10392,N_9758,N_9921);
xnor U10393 (N_10393,N_9860,N_9136);
and U10394 (N_10394,N_9532,N_9090);
xnor U10395 (N_10395,N_9646,N_9458);
nor U10396 (N_10396,N_9791,N_9582);
nor U10397 (N_10397,N_9058,N_9743);
xnor U10398 (N_10398,N_9500,N_9663);
or U10399 (N_10399,N_9352,N_9634);
nand U10400 (N_10400,N_9944,N_9415);
or U10401 (N_10401,N_9412,N_9420);
and U10402 (N_10402,N_9890,N_9102);
xnor U10403 (N_10403,N_9925,N_9878);
nor U10404 (N_10404,N_9287,N_9158);
nand U10405 (N_10405,N_9418,N_9961);
xnor U10406 (N_10406,N_9755,N_9444);
nor U10407 (N_10407,N_9592,N_9918);
or U10408 (N_10408,N_9360,N_9115);
xor U10409 (N_10409,N_9208,N_9949);
xnor U10410 (N_10410,N_9798,N_9009);
or U10411 (N_10411,N_9502,N_9853);
nand U10412 (N_10412,N_9061,N_9934);
or U10413 (N_10413,N_9452,N_9805);
xor U10414 (N_10414,N_9591,N_9571);
nand U10415 (N_10415,N_9358,N_9084);
nor U10416 (N_10416,N_9460,N_9184);
nand U10417 (N_10417,N_9982,N_9271);
and U10418 (N_10418,N_9196,N_9168);
or U10419 (N_10419,N_9482,N_9527);
xor U10420 (N_10420,N_9098,N_9631);
nand U10421 (N_10421,N_9750,N_9913);
nor U10422 (N_10422,N_9222,N_9696);
nor U10423 (N_10423,N_9575,N_9285);
nor U10424 (N_10424,N_9365,N_9176);
and U10425 (N_10425,N_9560,N_9725);
nor U10426 (N_10426,N_9511,N_9967);
and U10427 (N_10427,N_9394,N_9868);
or U10428 (N_10428,N_9998,N_9188);
xnor U10429 (N_10429,N_9808,N_9074);
or U10430 (N_10430,N_9278,N_9167);
and U10431 (N_10431,N_9181,N_9939);
or U10432 (N_10432,N_9284,N_9834);
nor U10433 (N_10433,N_9065,N_9627);
and U10434 (N_10434,N_9100,N_9772);
and U10435 (N_10435,N_9003,N_9060);
nand U10436 (N_10436,N_9789,N_9446);
and U10437 (N_10437,N_9342,N_9929);
nand U10438 (N_10438,N_9708,N_9800);
xor U10439 (N_10439,N_9698,N_9950);
nand U10440 (N_10440,N_9105,N_9118);
and U10441 (N_10441,N_9537,N_9622);
nand U10442 (N_10442,N_9613,N_9555);
nand U10443 (N_10443,N_9174,N_9354);
and U10444 (N_10444,N_9026,N_9143);
or U10445 (N_10445,N_9445,N_9764);
and U10446 (N_10446,N_9577,N_9605);
nor U10447 (N_10447,N_9189,N_9236);
and U10448 (N_10448,N_9059,N_9595);
or U10449 (N_10449,N_9387,N_9214);
nor U10450 (N_10450,N_9820,N_9162);
or U10451 (N_10451,N_9297,N_9014);
and U10452 (N_10452,N_9861,N_9328);
nor U10453 (N_10453,N_9041,N_9775);
and U10454 (N_10454,N_9647,N_9981);
nor U10455 (N_10455,N_9819,N_9047);
xnor U10456 (N_10456,N_9480,N_9332);
nor U10457 (N_10457,N_9963,N_9255);
xnor U10458 (N_10458,N_9465,N_9396);
nand U10459 (N_10459,N_9035,N_9971);
nor U10460 (N_10460,N_9265,N_9960);
nand U10461 (N_10461,N_9972,N_9023);
xnor U10462 (N_10462,N_9769,N_9548);
nand U10463 (N_10463,N_9008,N_9007);
xor U10464 (N_10464,N_9617,N_9702);
or U10465 (N_10465,N_9965,N_9195);
xnor U10466 (N_10466,N_9594,N_9183);
nand U10467 (N_10467,N_9716,N_9777);
nand U10468 (N_10468,N_9628,N_9516);
nor U10469 (N_10469,N_9642,N_9292);
xor U10470 (N_10470,N_9636,N_9568);
or U10471 (N_10471,N_9369,N_9321);
and U10472 (N_10472,N_9535,N_9414);
nor U10473 (N_10473,N_9128,N_9120);
or U10474 (N_10474,N_9043,N_9523);
and U10475 (N_10475,N_9487,N_9996);
xnor U10476 (N_10476,N_9346,N_9840);
nor U10477 (N_10477,N_9990,N_9833);
xor U10478 (N_10478,N_9191,N_9150);
xor U10479 (N_10479,N_9908,N_9529);
and U10480 (N_10480,N_9153,N_9241);
nor U10481 (N_10481,N_9904,N_9859);
or U10482 (N_10482,N_9651,N_9282);
and U10483 (N_10483,N_9276,N_9046);
and U10484 (N_10484,N_9273,N_9399);
or U10485 (N_10485,N_9674,N_9709);
nor U10486 (N_10486,N_9836,N_9454);
nand U10487 (N_10487,N_9559,N_9178);
or U10488 (N_10488,N_9875,N_9479);
or U10489 (N_10489,N_9633,N_9927);
xor U10490 (N_10490,N_9912,N_9863);
xor U10491 (N_10491,N_9212,N_9318);
or U10492 (N_10492,N_9019,N_9774);
nor U10493 (N_10493,N_9350,N_9896);
nand U10494 (N_10494,N_9397,N_9087);
nor U10495 (N_10495,N_9751,N_9012);
or U10496 (N_10496,N_9587,N_9070);
nand U10497 (N_10497,N_9437,N_9563);
nand U10498 (N_10498,N_9597,N_9562);
or U10499 (N_10499,N_9565,N_9324);
xnor U10500 (N_10500,N_9921,N_9041);
and U10501 (N_10501,N_9844,N_9345);
and U10502 (N_10502,N_9336,N_9123);
or U10503 (N_10503,N_9364,N_9685);
nor U10504 (N_10504,N_9218,N_9938);
xnor U10505 (N_10505,N_9921,N_9275);
and U10506 (N_10506,N_9892,N_9761);
nor U10507 (N_10507,N_9406,N_9263);
and U10508 (N_10508,N_9162,N_9107);
nand U10509 (N_10509,N_9457,N_9025);
or U10510 (N_10510,N_9635,N_9040);
and U10511 (N_10511,N_9663,N_9190);
nor U10512 (N_10512,N_9098,N_9025);
nor U10513 (N_10513,N_9940,N_9774);
or U10514 (N_10514,N_9757,N_9824);
nor U10515 (N_10515,N_9657,N_9551);
or U10516 (N_10516,N_9980,N_9845);
nand U10517 (N_10517,N_9693,N_9397);
nand U10518 (N_10518,N_9743,N_9397);
xor U10519 (N_10519,N_9244,N_9218);
nor U10520 (N_10520,N_9935,N_9280);
or U10521 (N_10521,N_9705,N_9676);
xnor U10522 (N_10522,N_9358,N_9616);
or U10523 (N_10523,N_9635,N_9310);
nand U10524 (N_10524,N_9157,N_9352);
nand U10525 (N_10525,N_9307,N_9389);
and U10526 (N_10526,N_9037,N_9998);
nor U10527 (N_10527,N_9803,N_9654);
nor U10528 (N_10528,N_9716,N_9883);
xnor U10529 (N_10529,N_9738,N_9042);
xnor U10530 (N_10530,N_9883,N_9148);
nand U10531 (N_10531,N_9453,N_9883);
or U10532 (N_10532,N_9096,N_9926);
or U10533 (N_10533,N_9149,N_9345);
and U10534 (N_10534,N_9997,N_9141);
nor U10535 (N_10535,N_9996,N_9280);
nor U10536 (N_10536,N_9067,N_9248);
and U10537 (N_10537,N_9178,N_9364);
nor U10538 (N_10538,N_9916,N_9296);
nor U10539 (N_10539,N_9382,N_9233);
and U10540 (N_10540,N_9378,N_9497);
xnor U10541 (N_10541,N_9006,N_9885);
or U10542 (N_10542,N_9607,N_9283);
nand U10543 (N_10543,N_9177,N_9547);
nand U10544 (N_10544,N_9936,N_9655);
xnor U10545 (N_10545,N_9916,N_9731);
nand U10546 (N_10546,N_9903,N_9999);
nand U10547 (N_10547,N_9360,N_9324);
nand U10548 (N_10548,N_9639,N_9951);
xor U10549 (N_10549,N_9612,N_9783);
nor U10550 (N_10550,N_9248,N_9283);
xor U10551 (N_10551,N_9723,N_9543);
xor U10552 (N_10552,N_9008,N_9090);
and U10553 (N_10553,N_9225,N_9482);
nand U10554 (N_10554,N_9120,N_9147);
and U10555 (N_10555,N_9099,N_9818);
xnor U10556 (N_10556,N_9964,N_9833);
xnor U10557 (N_10557,N_9162,N_9609);
nand U10558 (N_10558,N_9848,N_9943);
nor U10559 (N_10559,N_9097,N_9629);
nand U10560 (N_10560,N_9010,N_9561);
and U10561 (N_10561,N_9371,N_9916);
or U10562 (N_10562,N_9102,N_9278);
xor U10563 (N_10563,N_9620,N_9451);
or U10564 (N_10564,N_9426,N_9430);
xnor U10565 (N_10565,N_9639,N_9403);
nand U10566 (N_10566,N_9318,N_9710);
or U10567 (N_10567,N_9889,N_9342);
or U10568 (N_10568,N_9907,N_9529);
xnor U10569 (N_10569,N_9024,N_9511);
and U10570 (N_10570,N_9400,N_9406);
or U10571 (N_10571,N_9587,N_9320);
nand U10572 (N_10572,N_9468,N_9141);
nor U10573 (N_10573,N_9692,N_9406);
nand U10574 (N_10574,N_9543,N_9160);
nor U10575 (N_10575,N_9280,N_9464);
nand U10576 (N_10576,N_9249,N_9141);
xnor U10577 (N_10577,N_9506,N_9838);
or U10578 (N_10578,N_9295,N_9061);
or U10579 (N_10579,N_9410,N_9207);
nand U10580 (N_10580,N_9573,N_9499);
nor U10581 (N_10581,N_9252,N_9349);
nor U10582 (N_10582,N_9073,N_9854);
and U10583 (N_10583,N_9861,N_9330);
or U10584 (N_10584,N_9115,N_9419);
and U10585 (N_10585,N_9978,N_9757);
and U10586 (N_10586,N_9112,N_9700);
nand U10587 (N_10587,N_9183,N_9221);
nor U10588 (N_10588,N_9549,N_9260);
nand U10589 (N_10589,N_9322,N_9488);
xor U10590 (N_10590,N_9901,N_9135);
nand U10591 (N_10591,N_9397,N_9823);
and U10592 (N_10592,N_9294,N_9823);
xor U10593 (N_10593,N_9494,N_9330);
or U10594 (N_10594,N_9016,N_9350);
or U10595 (N_10595,N_9110,N_9827);
or U10596 (N_10596,N_9777,N_9465);
or U10597 (N_10597,N_9437,N_9819);
nand U10598 (N_10598,N_9988,N_9727);
or U10599 (N_10599,N_9556,N_9954);
xnor U10600 (N_10600,N_9113,N_9915);
xnor U10601 (N_10601,N_9711,N_9477);
xnor U10602 (N_10602,N_9491,N_9375);
and U10603 (N_10603,N_9362,N_9040);
and U10604 (N_10604,N_9148,N_9809);
and U10605 (N_10605,N_9939,N_9408);
nor U10606 (N_10606,N_9558,N_9663);
nor U10607 (N_10607,N_9936,N_9842);
xor U10608 (N_10608,N_9535,N_9969);
nand U10609 (N_10609,N_9738,N_9866);
nor U10610 (N_10610,N_9913,N_9049);
and U10611 (N_10611,N_9547,N_9414);
nor U10612 (N_10612,N_9393,N_9834);
nand U10613 (N_10613,N_9272,N_9088);
and U10614 (N_10614,N_9495,N_9021);
nand U10615 (N_10615,N_9459,N_9140);
or U10616 (N_10616,N_9371,N_9968);
nor U10617 (N_10617,N_9231,N_9317);
or U10618 (N_10618,N_9475,N_9803);
nand U10619 (N_10619,N_9362,N_9123);
nand U10620 (N_10620,N_9879,N_9470);
nor U10621 (N_10621,N_9956,N_9858);
nand U10622 (N_10622,N_9884,N_9278);
or U10623 (N_10623,N_9897,N_9592);
nor U10624 (N_10624,N_9610,N_9355);
and U10625 (N_10625,N_9852,N_9394);
nor U10626 (N_10626,N_9131,N_9579);
xnor U10627 (N_10627,N_9237,N_9886);
xor U10628 (N_10628,N_9189,N_9866);
xor U10629 (N_10629,N_9335,N_9899);
or U10630 (N_10630,N_9172,N_9529);
nor U10631 (N_10631,N_9140,N_9728);
nand U10632 (N_10632,N_9012,N_9329);
and U10633 (N_10633,N_9739,N_9537);
nand U10634 (N_10634,N_9966,N_9042);
and U10635 (N_10635,N_9331,N_9941);
nor U10636 (N_10636,N_9644,N_9290);
xor U10637 (N_10637,N_9022,N_9524);
xor U10638 (N_10638,N_9822,N_9729);
nand U10639 (N_10639,N_9039,N_9698);
nand U10640 (N_10640,N_9353,N_9307);
nor U10641 (N_10641,N_9976,N_9507);
nor U10642 (N_10642,N_9168,N_9656);
or U10643 (N_10643,N_9644,N_9587);
xnor U10644 (N_10644,N_9596,N_9359);
nand U10645 (N_10645,N_9738,N_9004);
xnor U10646 (N_10646,N_9804,N_9903);
xor U10647 (N_10647,N_9811,N_9723);
or U10648 (N_10648,N_9639,N_9836);
or U10649 (N_10649,N_9120,N_9477);
xor U10650 (N_10650,N_9696,N_9399);
nand U10651 (N_10651,N_9122,N_9772);
xor U10652 (N_10652,N_9141,N_9269);
and U10653 (N_10653,N_9165,N_9859);
nand U10654 (N_10654,N_9768,N_9323);
and U10655 (N_10655,N_9047,N_9603);
or U10656 (N_10656,N_9304,N_9327);
xnor U10657 (N_10657,N_9111,N_9115);
nand U10658 (N_10658,N_9251,N_9099);
nor U10659 (N_10659,N_9685,N_9151);
nor U10660 (N_10660,N_9623,N_9349);
xnor U10661 (N_10661,N_9421,N_9049);
xor U10662 (N_10662,N_9747,N_9800);
and U10663 (N_10663,N_9390,N_9340);
or U10664 (N_10664,N_9430,N_9557);
nor U10665 (N_10665,N_9491,N_9448);
nor U10666 (N_10666,N_9019,N_9010);
and U10667 (N_10667,N_9361,N_9220);
and U10668 (N_10668,N_9567,N_9669);
nand U10669 (N_10669,N_9080,N_9804);
nand U10670 (N_10670,N_9782,N_9180);
nand U10671 (N_10671,N_9152,N_9524);
nand U10672 (N_10672,N_9178,N_9902);
or U10673 (N_10673,N_9701,N_9155);
nor U10674 (N_10674,N_9568,N_9709);
xnor U10675 (N_10675,N_9777,N_9679);
nor U10676 (N_10676,N_9608,N_9584);
nor U10677 (N_10677,N_9119,N_9122);
nand U10678 (N_10678,N_9943,N_9600);
nor U10679 (N_10679,N_9420,N_9144);
nand U10680 (N_10680,N_9930,N_9307);
nor U10681 (N_10681,N_9217,N_9577);
nor U10682 (N_10682,N_9517,N_9588);
xnor U10683 (N_10683,N_9288,N_9331);
or U10684 (N_10684,N_9082,N_9719);
nor U10685 (N_10685,N_9306,N_9916);
nand U10686 (N_10686,N_9166,N_9628);
or U10687 (N_10687,N_9366,N_9350);
nor U10688 (N_10688,N_9244,N_9673);
and U10689 (N_10689,N_9690,N_9971);
and U10690 (N_10690,N_9570,N_9683);
and U10691 (N_10691,N_9219,N_9403);
or U10692 (N_10692,N_9070,N_9959);
nor U10693 (N_10693,N_9066,N_9605);
nand U10694 (N_10694,N_9040,N_9862);
and U10695 (N_10695,N_9744,N_9959);
and U10696 (N_10696,N_9317,N_9921);
or U10697 (N_10697,N_9332,N_9295);
xor U10698 (N_10698,N_9494,N_9655);
nand U10699 (N_10699,N_9613,N_9655);
nand U10700 (N_10700,N_9850,N_9102);
nand U10701 (N_10701,N_9841,N_9035);
xor U10702 (N_10702,N_9154,N_9210);
xor U10703 (N_10703,N_9148,N_9662);
xor U10704 (N_10704,N_9132,N_9555);
nand U10705 (N_10705,N_9000,N_9434);
xor U10706 (N_10706,N_9832,N_9354);
nand U10707 (N_10707,N_9152,N_9571);
nand U10708 (N_10708,N_9705,N_9152);
nor U10709 (N_10709,N_9056,N_9445);
or U10710 (N_10710,N_9334,N_9270);
xor U10711 (N_10711,N_9064,N_9997);
nand U10712 (N_10712,N_9738,N_9896);
xor U10713 (N_10713,N_9614,N_9268);
and U10714 (N_10714,N_9913,N_9423);
nand U10715 (N_10715,N_9952,N_9445);
and U10716 (N_10716,N_9739,N_9070);
xnor U10717 (N_10717,N_9275,N_9052);
nand U10718 (N_10718,N_9223,N_9315);
nor U10719 (N_10719,N_9391,N_9173);
and U10720 (N_10720,N_9459,N_9234);
and U10721 (N_10721,N_9981,N_9241);
or U10722 (N_10722,N_9746,N_9971);
or U10723 (N_10723,N_9704,N_9656);
and U10724 (N_10724,N_9849,N_9893);
nor U10725 (N_10725,N_9681,N_9996);
xor U10726 (N_10726,N_9516,N_9406);
nand U10727 (N_10727,N_9611,N_9763);
xor U10728 (N_10728,N_9013,N_9515);
nor U10729 (N_10729,N_9787,N_9663);
nand U10730 (N_10730,N_9167,N_9916);
or U10731 (N_10731,N_9345,N_9680);
and U10732 (N_10732,N_9125,N_9232);
xnor U10733 (N_10733,N_9735,N_9359);
nor U10734 (N_10734,N_9178,N_9152);
xor U10735 (N_10735,N_9977,N_9424);
nor U10736 (N_10736,N_9621,N_9220);
nor U10737 (N_10737,N_9145,N_9161);
or U10738 (N_10738,N_9908,N_9518);
or U10739 (N_10739,N_9268,N_9743);
nor U10740 (N_10740,N_9798,N_9265);
or U10741 (N_10741,N_9886,N_9209);
xor U10742 (N_10742,N_9202,N_9204);
nand U10743 (N_10743,N_9495,N_9644);
xor U10744 (N_10744,N_9372,N_9565);
xor U10745 (N_10745,N_9071,N_9174);
xnor U10746 (N_10746,N_9837,N_9132);
or U10747 (N_10747,N_9149,N_9119);
xnor U10748 (N_10748,N_9533,N_9032);
and U10749 (N_10749,N_9538,N_9191);
xnor U10750 (N_10750,N_9544,N_9033);
or U10751 (N_10751,N_9601,N_9847);
nor U10752 (N_10752,N_9751,N_9417);
xnor U10753 (N_10753,N_9974,N_9176);
or U10754 (N_10754,N_9651,N_9183);
or U10755 (N_10755,N_9435,N_9787);
or U10756 (N_10756,N_9504,N_9989);
or U10757 (N_10757,N_9977,N_9187);
xnor U10758 (N_10758,N_9726,N_9332);
or U10759 (N_10759,N_9751,N_9431);
xor U10760 (N_10760,N_9089,N_9254);
nor U10761 (N_10761,N_9926,N_9606);
nor U10762 (N_10762,N_9255,N_9304);
or U10763 (N_10763,N_9790,N_9733);
nor U10764 (N_10764,N_9397,N_9473);
and U10765 (N_10765,N_9386,N_9143);
xnor U10766 (N_10766,N_9908,N_9080);
xnor U10767 (N_10767,N_9046,N_9320);
xor U10768 (N_10768,N_9523,N_9922);
and U10769 (N_10769,N_9485,N_9458);
and U10770 (N_10770,N_9662,N_9756);
and U10771 (N_10771,N_9647,N_9893);
xnor U10772 (N_10772,N_9360,N_9993);
xnor U10773 (N_10773,N_9279,N_9355);
xor U10774 (N_10774,N_9694,N_9312);
and U10775 (N_10775,N_9673,N_9908);
xnor U10776 (N_10776,N_9092,N_9178);
and U10777 (N_10777,N_9636,N_9762);
xnor U10778 (N_10778,N_9887,N_9774);
nand U10779 (N_10779,N_9169,N_9554);
nand U10780 (N_10780,N_9621,N_9640);
nor U10781 (N_10781,N_9573,N_9253);
nor U10782 (N_10782,N_9069,N_9381);
or U10783 (N_10783,N_9006,N_9252);
or U10784 (N_10784,N_9754,N_9319);
xor U10785 (N_10785,N_9253,N_9076);
xor U10786 (N_10786,N_9372,N_9657);
xor U10787 (N_10787,N_9056,N_9456);
nand U10788 (N_10788,N_9940,N_9522);
and U10789 (N_10789,N_9016,N_9100);
nand U10790 (N_10790,N_9366,N_9763);
or U10791 (N_10791,N_9619,N_9294);
or U10792 (N_10792,N_9464,N_9071);
and U10793 (N_10793,N_9828,N_9921);
and U10794 (N_10794,N_9210,N_9955);
nor U10795 (N_10795,N_9154,N_9542);
nor U10796 (N_10796,N_9724,N_9898);
nand U10797 (N_10797,N_9969,N_9632);
xor U10798 (N_10798,N_9994,N_9239);
xnor U10799 (N_10799,N_9243,N_9322);
nor U10800 (N_10800,N_9829,N_9563);
nor U10801 (N_10801,N_9561,N_9437);
or U10802 (N_10802,N_9687,N_9297);
and U10803 (N_10803,N_9598,N_9440);
xnor U10804 (N_10804,N_9447,N_9778);
or U10805 (N_10805,N_9593,N_9725);
nor U10806 (N_10806,N_9945,N_9855);
or U10807 (N_10807,N_9419,N_9240);
xnor U10808 (N_10808,N_9316,N_9670);
xor U10809 (N_10809,N_9268,N_9365);
nand U10810 (N_10810,N_9531,N_9594);
or U10811 (N_10811,N_9734,N_9159);
or U10812 (N_10812,N_9435,N_9557);
nor U10813 (N_10813,N_9580,N_9671);
nor U10814 (N_10814,N_9162,N_9588);
and U10815 (N_10815,N_9436,N_9313);
and U10816 (N_10816,N_9259,N_9002);
nor U10817 (N_10817,N_9322,N_9593);
and U10818 (N_10818,N_9385,N_9767);
nand U10819 (N_10819,N_9888,N_9061);
xnor U10820 (N_10820,N_9691,N_9687);
nor U10821 (N_10821,N_9137,N_9659);
nand U10822 (N_10822,N_9591,N_9577);
and U10823 (N_10823,N_9098,N_9660);
or U10824 (N_10824,N_9728,N_9621);
xor U10825 (N_10825,N_9267,N_9568);
nor U10826 (N_10826,N_9604,N_9125);
or U10827 (N_10827,N_9724,N_9024);
xnor U10828 (N_10828,N_9885,N_9431);
or U10829 (N_10829,N_9265,N_9040);
nor U10830 (N_10830,N_9452,N_9027);
or U10831 (N_10831,N_9843,N_9494);
and U10832 (N_10832,N_9414,N_9995);
nor U10833 (N_10833,N_9995,N_9656);
nand U10834 (N_10834,N_9275,N_9830);
nor U10835 (N_10835,N_9357,N_9345);
and U10836 (N_10836,N_9260,N_9370);
nand U10837 (N_10837,N_9422,N_9214);
nand U10838 (N_10838,N_9114,N_9298);
xor U10839 (N_10839,N_9186,N_9928);
xnor U10840 (N_10840,N_9625,N_9745);
nor U10841 (N_10841,N_9760,N_9597);
and U10842 (N_10842,N_9650,N_9876);
or U10843 (N_10843,N_9101,N_9512);
nor U10844 (N_10844,N_9682,N_9108);
or U10845 (N_10845,N_9018,N_9263);
and U10846 (N_10846,N_9881,N_9157);
and U10847 (N_10847,N_9636,N_9603);
nor U10848 (N_10848,N_9243,N_9258);
and U10849 (N_10849,N_9752,N_9420);
xor U10850 (N_10850,N_9900,N_9778);
xor U10851 (N_10851,N_9529,N_9978);
and U10852 (N_10852,N_9250,N_9293);
xnor U10853 (N_10853,N_9996,N_9855);
nor U10854 (N_10854,N_9963,N_9813);
xnor U10855 (N_10855,N_9467,N_9689);
and U10856 (N_10856,N_9771,N_9205);
xor U10857 (N_10857,N_9522,N_9520);
nor U10858 (N_10858,N_9338,N_9044);
nand U10859 (N_10859,N_9434,N_9041);
nand U10860 (N_10860,N_9821,N_9233);
or U10861 (N_10861,N_9318,N_9034);
xnor U10862 (N_10862,N_9739,N_9672);
or U10863 (N_10863,N_9581,N_9844);
and U10864 (N_10864,N_9867,N_9161);
nor U10865 (N_10865,N_9754,N_9828);
or U10866 (N_10866,N_9253,N_9144);
or U10867 (N_10867,N_9407,N_9606);
nor U10868 (N_10868,N_9170,N_9103);
xnor U10869 (N_10869,N_9061,N_9177);
nor U10870 (N_10870,N_9362,N_9476);
nand U10871 (N_10871,N_9398,N_9527);
nor U10872 (N_10872,N_9608,N_9654);
and U10873 (N_10873,N_9711,N_9365);
nor U10874 (N_10874,N_9164,N_9067);
xnor U10875 (N_10875,N_9502,N_9810);
nor U10876 (N_10876,N_9679,N_9410);
nor U10877 (N_10877,N_9301,N_9394);
and U10878 (N_10878,N_9080,N_9281);
nand U10879 (N_10879,N_9020,N_9062);
xor U10880 (N_10880,N_9698,N_9463);
or U10881 (N_10881,N_9832,N_9705);
nor U10882 (N_10882,N_9273,N_9951);
or U10883 (N_10883,N_9560,N_9131);
xor U10884 (N_10884,N_9661,N_9758);
nor U10885 (N_10885,N_9363,N_9879);
xor U10886 (N_10886,N_9985,N_9713);
nor U10887 (N_10887,N_9325,N_9291);
and U10888 (N_10888,N_9952,N_9271);
or U10889 (N_10889,N_9666,N_9842);
nand U10890 (N_10890,N_9484,N_9596);
xor U10891 (N_10891,N_9778,N_9925);
nor U10892 (N_10892,N_9077,N_9648);
or U10893 (N_10893,N_9840,N_9549);
nor U10894 (N_10894,N_9182,N_9579);
and U10895 (N_10895,N_9824,N_9680);
nor U10896 (N_10896,N_9284,N_9810);
and U10897 (N_10897,N_9618,N_9377);
nand U10898 (N_10898,N_9917,N_9957);
or U10899 (N_10899,N_9641,N_9591);
nand U10900 (N_10900,N_9858,N_9851);
or U10901 (N_10901,N_9725,N_9521);
or U10902 (N_10902,N_9115,N_9906);
nor U10903 (N_10903,N_9983,N_9068);
nand U10904 (N_10904,N_9876,N_9210);
nand U10905 (N_10905,N_9512,N_9404);
nor U10906 (N_10906,N_9525,N_9166);
nand U10907 (N_10907,N_9041,N_9003);
nand U10908 (N_10908,N_9889,N_9431);
nor U10909 (N_10909,N_9677,N_9701);
nand U10910 (N_10910,N_9530,N_9200);
and U10911 (N_10911,N_9099,N_9939);
xor U10912 (N_10912,N_9819,N_9000);
nor U10913 (N_10913,N_9758,N_9286);
nor U10914 (N_10914,N_9309,N_9670);
nor U10915 (N_10915,N_9956,N_9253);
nor U10916 (N_10916,N_9777,N_9904);
nand U10917 (N_10917,N_9446,N_9230);
nor U10918 (N_10918,N_9346,N_9960);
nor U10919 (N_10919,N_9822,N_9634);
and U10920 (N_10920,N_9028,N_9143);
nor U10921 (N_10921,N_9242,N_9936);
xnor U10922 (N_10922,N_9967,N_9703);
or U10923 (N_10923,N_9158,N_9564);
and U10924 (N_10924,N_9367,N_9477);
xor U10925 (N_10925,N_9685,N_9505);
xor U10926 (N_10926,N_9119,N_9751);
xor U10927 (N_10927,N_9351,N_9111);
nand U10928 (N_10928,N_9486,N_9803);
nand U10929 (N_10929,N_9206,N_9999);
xnor U10930 (N_10930,N_9880,N_9686);
nor U10931 (N_10931,N_9270,N_9876);
nand U10932 (N_10932,N_9271,N_9061);
nand U10933 (N_10933,N_9489,N_9702);
xnor U10934 (N_10934,N_9069,N_9629);
xnor U10935 (N_10935,N_9436,N_9626);
xor U10936 (N_10936,N_9023,N_9028);
and U10937 (N_10937,N_9388,N_9624);
nor U10938 (N_10938,N_9719,N_9750);
xor U10939 (N_10939,N_9257,N_9786);
and U10940 (N_10940,N_9568,N_9920);
xnor U10941 (N_10941,N_9073,N_9503);
and U10942 (N_10942,N_9744,N_9986);
xnor U10943 (N_10943,N_9617,N_9686);
nand U10944 (N_10944,N_9496,N_9653);
nand U10945 (N_10945,N_9942,N_9946);
and U10946 (N_10946,N_9415,N_9029);
nand U10947 (N_10947,N_9175,N_9152);
nor U10948 (N_10948,N_9053,N_9072);
xnor U10949 (N_10949,N_9360,N_9779);
nor U10950 (N_10950,N_9285,N_9594);
or U10951 (N_10951,N_9312,N_9017);
or U10952 (N_10952,N_9929,N_9203);
or U10953 (N_10953,N_9256,N_9191);
nand U10954 (N_10954,N_9317,N_9008);
nor U10955 (N_10955,N_9293,N_9995);
and U10956 (N_10956,N_9601,N_9256);
and U10957 (N_10957,N_9507,N_9402);
xnor U10958 (N_10958,N_9589,N_9499);
or U10959 (N_10959,N_9324,N_9401);
xnor U10960 (N_10960,N_9237,N_9743);
nor U10961 (N_10961,N_9781,N_9721);
and U10962 (N_10962,N_9869,N_9383);
nand U10963 (N_10963,N_9035,N_9598);
xnor U10964 (N_10964,N_9518,N_9007);
nand U10965 (N_10965,N_9757,N_9727);
and U10966 (N_10966,N_9004,N_9034);
xnor U10967 (N_10967,N_9534,N_9842);
xnor U10968 (N_10968,N_9608,N_9509);
nand U10969 (N_10969,N_9671,N_9481);
nor U10970 (N_10970,N_9561,N_9656);
nor U10971 (N_10971,N_9443,N_9431);
and U10972 (N_10972,N_9606,N_9099);
and U10973 (N_10973,N_9627,N_9791);
or U10974 (N_10974,N_9255,N_9817);
and U10975 (N_10975,N_9694,N_9791);
or U10976 (N_10976,N_9043,N_9923);
nor U10977 (N_10977,N_9239,N_9430);
and U10978 (N_10978,N_9483,N_9749);
or U10979 (N_10979,N_9734,N_9141);
nor U10980 (N_10980,N_9989,N_9506);
nand U10981 (N_10981,N_9356,N_9816);
xor U10982 (N_10982,N_9352,N_9411);
nor U10983 (N_10983,N_9254,N_9835);
nand U10984 (N_10984,N_9504,N_9916);
xnor U10985 (N_10985,N_9419,N_9207);
and U10986 (N_10986,N_9381,N_9146);
nand U10987 (N_10987,N_9864,N_9333);
nand U10988 (N_10988,N_9242,N_9873);
and U10989 (N_10989,N_9724,N_9008);
and U10990 (N_10990,N_9442,N_9668);
xor U10991 (N_10991,N_9801,N_9778);
xnor U10992 (N_10992,N_9743,N_9440);
nand U10993 (N_10993,N_9338,N_9286);
or U10994 (N_10994,N_9026,N_9937);
nor U10995 (N_10995,N_9391,N_9710);
or U10996 (N_10996,N_9189,N_9519);
or U10997 (N_10997,N_9443,N_9246);
and U10998 (N_10998,N_9748,N_9325);
nand U10999 (N_10999,N_9428,N_9812);
nand U11000 (N_11000,N_10290,N_10144);
xnor U11001 (N_11001,N_10641,N_10998);
and U11002 (N_11002,N_10441,N_10390);
and U11003 (N_11003,N_10025,N_10425);
or U11004 (N_11004,N_10659,N_10191);
and U11005 (N_11005,N_10119,N_10525);
or U11006 (N_11006,N_10005,N_10829);
nand U11007 (N_11007,N_10939,N_10646);
xnor U11008 (N_11008,N_10462,N_10899);
xnor U11009 (N_11009,N_10850,N_10677);
nor U11010 (N_11010,N_10093,N_10698);
xor U11011 (N_11011,N_10630,N_10297);
nor U11012 (N_11012,N_10758,N_10350);
xor U11013 (N_11013,N_10812,N_10178);
nand U11014 (N_11014,N_10721,N_10931);
or U11015 (N_11015,N_10426,N_10387);
or U11016 (N_11016,N_10320,N_10354);
nand U11017 (N_11017,N_10436,N_10953);
or U11018 (N_11018,N_10832,N_10226);
or U11019 (N_11019,N_10032,N_10273);
nand U11020 (N_11020,N_10415,N_10193);
xor U11021 (N_11021,N_10932,N_10607);
and U11022 (N_11022,N_10835,N_10469);
nor U11023 (N_11023,N_10448,N_10565);
and U11024 (N_11024,N_10388,N_10050);
or U11025 (N_11025,N_10443,N_10514);
and U11026 (N_11026,N_10516,N_10192);
nand U11027 (N_11027,N_10082,N_10530);
xor U11028 (N_11028,N_10976,N_10960);
and U11029 (N_11029,N_10456,N_10055);
nand U11030 (N_11030,N_10317,N_10541);
and U11031 (N_11031,N_10464,N_10275);
xor U11032 (N_11032,N_10620,N_10311);
and U11033 (N_11033,N_10246,N_10162);
and U11034 (N_11034,N_10805,N_10625);
nand U11035 (N_11035,N_10225,N_10575);
nand U11036 (N_11036,N_10289,N_10324);
nor U11037 (N_11037,N_10858,N_10653);
and U11038 (N_11038,N_10529,N_10983);
nand U11039 (N_11039,N_10382,N_10654);
nand U11040 (N_11040,N_10287,N_10558);
nor U11041 (N_11041,N_10774,N_10295);
or U11042 (N_11042,N_10864,N_10474);
nand U11043 (N_11043,N_10458,N_10509);
and U11044 (N_11044,N_10680,N_10455);
or U11045 (N_11045,N_10650,N_10810);
nand U11046 (N_11046,N_10011,N_10971);
and U11047 (N_11047,N_10566,N_10229);
and U11048 (N_11048,N_10033,N_10645);
and U11049 (N_11049,N_10172,N_10555);
nor U11050 (N_11050,N_10635,N_10498);
nand U11051 (N_11051,N_10803,N_10522);
and U11052 (N_11052,N_10149,N_10790);
nor U11053 (N_11053,N_10450,N_10663);
or U11054 (N_11054,N_10793,N_10277);
nand U11055 (N_11055,N_10466,N_10628);
xnor U11056 (N_11056,N_10985,N_10940);
xor U11057 (N_11057,N_10293,N_10465);
and U11058 (N_11058,N_10769,N_10763);
nand U11059 (N_11059,N_10184,N_10512);
nand U11060 (N_11060,N_10696,N_10434);
nor U11061 (N_11061,N_10708,N_10956);
and U11062 (N_11062,N_10014,N_10564);
nor U11063 (N_11063,N_10261,N_10389);
or U11064 (N_11064,N_10271,N_10400);
nor U11065 (N_11065,N_10328,N_10705);
or U11066 (N_11066,N_10232,N_10840);
xor U11067 (N_11067,N_10775,N_10923);
nor U11068 (N_11068,N_10692,N_10737);
xnor U11069 (N_11069,N_10283,N_10588);
or U11070 (N_11070,N_10594,N_10164);
and U11071 (N_11071,N_10207,N_10276);
nor U11072 (N_11072,N_10726,N_10583);
or U11073 (N_11073,N_10623,N_10199);
nand U11074 (N_11074,N_10823,N_10347);
xor U11075 (N_11075,N_10013,N_10064);
nand U11076 (N_11076,N_10286,N_10930);
and U11077 (N_11077,N_10561,N_10539);
or U11078 (N_11078,N_10743,N_10560);
nor U11079 (N_11079,N_10242,N_10422);
and U11080 (N_11080,N_10490,N_10893);
or U11081 (N_11081,N_10127,N_10581);
nand U11082 (N_11082,N_10665,N_10611);
nand U11083 (N_11083,N_10818,N_10613);
and U11084 (N_11084,N_10385,N_10167);
xor U11085 (N_11085,N_10878,N_10402);
xor U11086 (N_11086,N_10264,N_10314);
nor U11087 (N_11087,N_10118,N_10648);
nor U11088 (N_11088,N_10221,N_10768);
nor U11089 (N_11089,N_10223,N_10218);
and U11090 (N_11090,N_10622,N_10727);
nand U11091 (N_11091,N_10955,N_10346);
nand U11092 (N_11092,N_10568,N_10690);
and U11093 (N_11093,N_10278,N_10291);
nor U11094 (N_11094,N_10305,N_10247);
and U11095 (N_11095,N_10656,N_10671);
nor U11096 (N_11096,N_10559,N_10517);
xor U11097 (N_11097,N_10703,N_10991);
or U11098 (N_11098,N_10492,N_10508);
xor U11099 (N_11099,N_10567,N_10658);
or U11100 (N_11100,N_10699,N_10134);
nor U11101 (N_11101,N_10384,N_10020);
nor U11102 (N_11102,N_10777,N_10981);
and U11103 (N_11103,N_10528,N_10478);
xor U11104 (N_11104,N_10335,N_10724);
and U11105 (N_11105,N_10959,N_10437);
or U11106 (N_11106,N_10795,N_10361);
nand U11107 (N_11107,N_10824,N_10964);
nand U11108 (N_11108,N_10053,N_10040);
nor U11109 (N_11109,N_10058,N_10003);
nor U11110 (N_11110,N_10380,N_10879);
xnor U11111 (N_11111,N_10066,N_10105);
xor U11112 (N_11112,N_10449,N_10044);
nor U11113 (N_11113,N_10706,N_10181);
nand U11114 (N_11114,N_10921,N_10573);
nor U11115 (N_11115,N_10738,N_10967);
nand U11116 (N_11116,N_10188,N_10935);
and U11117 (N_11117,N_10589,N_10201);
nand U11118 (N_11118,N_10258,N_10109);
or U11119 (N_11119,N_10231,N_10834);
nand U11120 (N_11120,N_10077,N_10651);
nand U11121 (N_11121,N_10407,N_10262);
or U11122 (N_11122,N_10543,N_10632);
nand U11123 (N_11123,N_10015,N_10198);
or U11124 (N_11124,N_10533,N_10486);
xor U11125 (N_11125,N_10787,N_10334);
nand U11126 (N_11126,N_10799,N_10019);
xnor U11127 (N_11127,N_10197,N_10860);
nor U11128 (N_11128,N_10155,N_10554);
nor U11129 (N_11129,N_10776,N_10298);
and U11130 (N_11130,N_10755,N_10084);
xnor U11131 (N_11131,N_10256,N_10969);
nor U11132 (N_11132,N_10664,N_10368);
xor U11133 (N_11133,N_10418,N_10308);
and U11134 (N_11134,N_10911,N_10500);
or U11135 (N_11135,N_10804,N_10740);
or U11136 (N_11136,N_10000,N_10537);
nand U11137 (N_11137,N_10419,N_10997);
xnor U11138 (N_11138,N_10545,N_10120);
nor U11139 (N_11139,N_10943,N_10213);
nand U11140 (N_11140,N_10615,N_10948);
nand U11141 (N_11141,N_10610,N_10202);
or U11142 (N_11142,N_10616,N_10898);
and U11143 (N_11143,N_10966,N_10639);
and U11144 (N_11144,N_10037,N_10666);
nor U11145 (N_11145,N_10596,N_10900);
or U11146 (N_11146,N_10331,N_10060);
xor U11147 (N_11147,N_10428,N_10585);
and U11148 (N_11148,N_10126,N_10240);
xnor U11149 (N_11149,N_10054,N_10243);
xnor U11150 (N_11150,N_10435,N_10391);
or U11151 (N_11151,N_10863,N_10686);
xnor U11152 (N_11152,N_10854,N_10160);
xnor U11153 (N_11153,N_10174,N_10457);
nor U11154 (N_11154,N_10709,N_10749);
and U11155 (N_11155,N_10351,N_10977);
xor U11156 (N_11156,N_10504,N_10326);
nand U11157 (N_11157,N_10926,N_10381);
or U11158 (N_11158,N_10791,N_10353);
and U11159 (N_11159,N_10846,N_10395);
xnor U11160 (N_11160,N_10936,N_10338);
nor U11161 (N_11161,N_10035,N_10413);
nand U11162 (N_11162,N_10159,N_10339);
xor U11163 (N_11163,N_10729,N_10867);
xnor U11164 (N_11164,N_10992,N_10248);
nor U11165 (N_11165,N_10039,N_10770);
nor U11166 (N_11166,N_10257,N_10125);
or U11167 (N_11167,N_10587,N_10085);
and U11168 (N_11168,N_10057,N_10715);
or U11169 (N_11169,N_10111,N_10195);
nor U11170 (N_11170,N_10779,N_10820);
nand U11171 (N_11171,N_10978,N_10074);
nand U11172 (N_11172,N_10006,N_10771);
nor U11173 (N_11173,N_10087,N_10963);
or U11174 (N_11174,N_10446,N_10440);
xnor U11175 (N_11175,N_10461,N_10767);
and U11176 (N_11176,N_10279,N_10333);
and U11177 (N_11177,N_10136,N_10376);
xor U11178 (N_11178,N_10725,N_10379);
or U11179 (N_11179,N_10439,N_10882);
or U11180 (N_11180,N_10608,N_10780);
and U11181 (N_11181,N_10688,N_10957);
or U11182 (N_11182,N_10051,N_10527);
or U11183 (N_11183,N_10370,N_10875);
xnor U11184 (N_11184,N_10756,N_10460);
nor U11185 (N_11185,N_10481,N_10392);
or U11186 (N_11186,N_10154,N_10473);
nand U11187 (N_11187,N_10572,N_10274);
nand U11188 (N_11188,N_10371,N_10300);
nor U11189 (N_11189,N_10031,N_10430);
nor U11190 (N_11190,N_10821,N_10292);
and U11191 (N_11191,N_10970,N_10176);
or U11192 (N_11192,N_10604,N_10378);
nor U11193 (N_11193,N_10644,N_10151);
and U11194 (N_11194,N_10284,N_10761);
and U11195 (N_11195,N_10913,N_10502);
nor U11196 (N_11196,N_10903,N_10954);
nor U11197 (N_11197,N_10765,N_10036);
or U11198 (N_11198,N_10952,N_10364);
nor U11199 (N_11199,N_10470,N_10547);
nor U11200 (N_11200,N_10847,N_10432);
and U11201 (N_11201,N_10049,N_10757);
nand U11202 (N_11202,N_10802,N_10816);
or U11203 (N_11203,N_10177,N_10012);
nor U11204 (N_11204,N_10549,N_10227);
nor U11205 (N_11205,N_10024,N_10121);
xor U11206 (N_11206,N_10336,N_10497);
xnor U11207 (N_11207,N_10404,N_10467);
nor U11208 (N_11208,N_10079,N_10747);
nand U11209 (N_11209,N_10906,N_10208);
nand U11210 (N_11210,N_10365,N_10447);
and U11211 (N_11211,N_10260,N_10546);
and U11212 (N_11212,N_10752,N_10551);
or U11213 (N_11213,N_10796,N_10112);
nand U11214 (N_11214,N_10577,N_10807);
or U11215 (N_11215,N_10949,N_10113);
nor U11216 (N_11216,N_10045,N_10717);
and U11217 (N_11217,N_10844,N_10582);
or U11218 (N_11218,N_10406,N_10236);
nand U11219 (N_11219,N_10100,N_10316);
xor U11220 (N_11220,N_10341,N_10961);
nand U11221 (N_11221,N_10189,N_10968);
xnor U11222 (N_11222,N_10141,N_10912);
xnor U11223 (N_11223,N_10806,N_10597);
xor U11224 (N_11224,N_10944,N_10520);
xor U11225 (N_11225,N_10890,N_10785);
nor U11226 (N_11226,N_10866,N_10786);
and U11227 (N_11227,N_10482,N_10670);
nand U11228 (N_11228,N_10831,N_10444);
nand U11229 (N_11229,N_10748,N_10750);
xor U11230 (N_11230,N_10073,N_10280);
nand U11231 (N_11231,N_10798,N_10814);
or U11232 (N_11232,N_10209,N_10693);
and U11233 (N_11233,N_10822,N_10251);
nor U11234 (N_11234,N_10255,N_10634);
nor U11235 (N_11235,N_10212,N_10532);
xor U11236 (N_11236,N_10745,N_10010);
and U11237 (N_11237,N_10161,N_10660);
nand U11238 (N_11238,N_10168,N_10133);
or U11239 (N_11239,N_10228,N_10506);
or U11240 (N_11240,N_10367,N_10094);
nand U11241 (N_11241,N_10179,N_10009);
and U11242 (N_11242,N_10163,N_10318);
nor U11243 (N_11243,N_10679,N_10783);
or U11244 (N_11244,N_10678,N_10951);
xor U11245 (N_11245,N_10683,N_10800);
and U11246 (N_11246,N_10222,N_10856);
nand U11247 (N_11247,N_10617,N_10919);
and U11248 (N_11248,N_10781,N_10602);
nand U11249 (N_11249,N_10249,N_10494);
and U11250 (N_11250,N_10873,N_10048);
xnor U11251 (N_11251,N_10237,N_10828);
nand U11252 (N_11252,N_10103,N_10042);
or U11253 (N_11253,N_10838,N_10910);
or U11254 (N_11254,N_10590,N_10238);
xnor U11255 (N_11255,N_10685,N_10322);
xnor U11256 (N_11256,N_10116,N_10217);
nor U11257 (N_11257,N_10669,N_10214);
nand U11258 (N_11258,N_10095,N_10947);
xor U11259 (N_11259,N_10485,N_10059);
and U11260 (N_11260,N_10928,N_10267);
and U11261 (N_11261,N_10123,N_10052);
xnor U11262 (N_11262,N_10984,N_10496);
nand U11263 (N_11263,N_10989,N_10313);
or U11264 (N_11264,N_10534,N_10489);
xnor U11265 (N_11265,N_10886,N_10171);
xor U11266 (N_11266,N_10934,N_10096);
nor U11267 (N_11267,N_10190,N_10330);
or U11268 (N_11268,N_10894,N_10897);
nand U11269 (N_11269,N_10386,N_10398);
and U11270 (N_11270,N_10165,N_10946);
or U11271 (N_11271,N_10974,N_10720);
or U11272 (N_11272,N_10902,N_10028);
and U11273 (N_11273,N_10072,N_10716);
xnor U11274 (N_11274,N_10701,N_10215);
nand U11275 (N_11275,N_10099,N_10071);
xnor U11276 (N_11276,N_10405,N_10146);
xnor U11277 (N_11277,N_10410,N_10578);
nand U11278 (N_11278,N_10076,N_10301);
or U11279 (N_11279,N_10252,N_10266);
or U11280 (N_11280,N_10417,N_10175);
nor U11281 (N_11281,N_10157,N_10086);
nand U11282 (N_11282,N_10224,N_10642);
nor U11283 (N_11283,N_10401,N_10092);
nor U11284 (N_11284,N_10833,N_10332);
or U11285 (N_11285,N_10114,N_10345);
or U11286 (N_11286,N_10988,N_10817);
xor U11287 (N_11287,N_10098,N_10742);
nand U11288 (N_11288,N_10204,N_10891);
xnor U11289 (N_11289,N_10744,N_10102);
nand U11290 (N_11290,N_10431,N_10523);
and U11291 (N_11291,N_10865,N_10859);
or U11292 (N_11292,N_10626,N_10689);
nor U11293 (N_11293,N_10841,N_10924);
xnor U11294 (N_11294,N_10029,N_10922);
or U11295 (N_11295,N_10973,N_10147);
and U11296 (N_11296,N_10403,N_10241);
or U11297 (N_11297,N_10995,N_10294);
xnor U11298 (N_11298,N_10915,N_10463);
xor U11299 (N_11299,N_10695,N_10580);
or U11300 (N_11300,N_10062,N_10453);
nor U11301 (N_11301,N_10396,N_10746);
xnor U11302 (N_11302,N_10047,N_10366);
xnor U11303 (N_11303,N_10186,N_10857);
or U11304 (N_11304,N_10905,N_10811);
or U11305 (N_11305,N_10618,N_10837);
xor U11306 (N_11306,N_10312,N_10574);
and U11307 (N_11307,N_10021,N_10704);
xor U11308 (N_11308,N_10667,N_10139);
and U11309 (N_11309,N_10515,N_10621);
nor U11310 (N_11310,N_10067,N_10375);
xor U11311 (N_11311,N_10107,N_10090);
and U11312 (N_11312,N_10356,N_10309);
nor U11313 (N_11313,N_10288,N_10488);
nor U11314 (N_11314,N_10531,N_10479);
nor U11315 (N_11315,N_10476,N_10722);
nor U11316 (N_11316,N_10263,N_10372);
nand U11317 (N_11317,N_10684,N_10383);
nor U11318 (N_11318,N_10929,N_10357);
or U11319 (N_11319,N_10836,N_10627);
or U11320 (N_11320,N_10895,N_10239);
nor U11321 (N_11321,N_10156,N_10016);
xor U11322 (N_11322,N_10150,N_10319);
and U11323 (N_11323,N_10672,N_10868);
and U11324 (N_11324,N_10920,N_10591);
nand U11325 (N_11325,N_10254,N_10234);
nor U11326 (N_11326,N_10938,N_10736);
or U11327 (N_11327,N_10614,N_10362);
nand U11328 (N_11328,N_10250,N_10612);
and U11329 (N_11329,N_10268,N_10348);
nor U11330 (N_11330,N_10751,N_10408);
or U11331 (N_11331,N_10495,N_10907);
xor U11332 (N_11332,N_10004,N_10472);
and U11333 (N_11333,N_10491,N_10813);
xor U11334 (N_11334,N_10916,N_10877);
nor U11335 (N_11335,N_10571,N_10142);
nand U11336 (N_11336,N_10083,N_10445);
and U11337 (N_11337,N_10719,N_10206);
xnor U11338 (N_11338,N_10662,N_10697);
or U11339 (N_11339,N_10373,N_10210);
and U11340 (N_11340,N_10526,N_10080);
nand U11341 (N_11341,N_10302,N_10412);
or U11342 (N_11342,N_10553,N_10304);
nor U11343 (N_11343,N_10979,N_10593);
nor U11344 (N_11344,N_10281,N_10323);
and U11345 (N_11345,N_10609,N_10409);
xnor U11346 (N_11346,N_10732,N_10994);
nand U11347 (N_11347,N_10089,N_10540);
or U11348 (N_11348,N_10637,N_10987);
or U11349 (N_11349,N_10888,N_10908);
or U11350 (N_11350,N_10676,N_10723);
or U11351 (N_11351,N_10861,N_10493);
xnor U11352 (N_11352,N_10592,N_10173);
or U11353 (N_11353,N_10687,N_10801);
xor U11354 (N_11354,N_10416,N_10883);
and U11355 (N_11355,N_10870,N_10982);
and U11356 (N_11356,N_10007,N_10788);
nand U11357 (N_11357,N_10562,N_10216);
nor U11358 (N_11358,N_10603,N_10359);
or U11359 (N_11359,N_10892,N_10414);
nand U11360 (N_11360,N_10138,N_10584);
and U11361 (N_11361,N_10315,N_10342);
nor U11362 (N_11362,N_10945,N_10731);
and U11363 (N_11363,N_10794,N_10975);
and U11364 (N_11364,N_10536,N_10942);
and U11365 (N_11365,N_10675,N_10862);
nor U11366 (N_11366,N_10424,N_10451);
nand U11367 (N_11367,N_10735,N_10933);
or U11368 (N_11368,N_10483,N_10511);
xor U11369 (N_11369,N_10754,N_10130);
xor U11370 (N_11370,N_10972,N_10586);
and U11371 (N_11371,N_10484,N_10576);
nor U11372 (N_11372,N_10827,N_10852);
and U11373 (N_11373,N_10137,N_10605);
or U11374 (N_11374,N_10475,N_10550);
or U11375 (N_11375,N_10990,N_10681);
and U11376 (N_11376,N_10600,N_10760);
nand U11377 (N_11377,N_10631,N_10097);
xnor U11378 (N_11378,N_10842,N_10018);
nand U11379 (N_11379,N_10329,N_10694);
and U11380 (N_11380,N_10638,N_10282);
or U11381 (N_11381,N_10122,N_10046);
nand U11382 (N_11382,N_10548,N_10700);
xnor U11383 (N_11383,N_10002,N_10043);
nand U11384 (N_11384,N_10855,N_10411);
and U11385 (N_11385,N_10885,N_10106);
nor U11386 (N_11386,N_10393,N_10299);
or U11387 (N_11387,N_10285,N_10194);
or U11388 (N_11388,N_10219,N_10340);
and U11389 (N_11389,N_10950,N_10211);
nor U11390 (N_11390,N_10358,N_10499);
nand U11391 (N_11391,N_10187,N_10235);
xor U11392 (N_11392,N_10454,N_10182);
nand U11393 (N_11393,N_10429,N_10598);
and U11394 (N_11394,N_10881,N_10741);
or U11395 (N_11395,N_10253,N_10369);
or U11396 (N_11396,N_10081,N_10017);
and U11397 (N_11397,N_10682,N_10220);
or U11398 (N_11398,N_10022,N_10918);
or U11399 (N_11399,N_10519,N_10069);
nor U11400 (N_11400,N_10713,N_10148);
nand U11401 (N_11401,N_10128,N_10034);
and U11402 (N_11402,N_10360,N_10487);
or U11403 (N_11403,N_10965,N_10296);
or U11404 (N_11404,N_10117,N_10739);
and U11405 (N_11405,N_10962,N_10880);
nor U11406 (N_11406,N_10026,N_10230);
nor U11407 (N_11407,N_10327,N_10784);
nor U11408 (N_11408,N_10169,N_10185);
nand U11409 (N_11409,N_10710,N_10909);
xor U11410 (N_11410,N_10343,N_10674);
nor U11411 (N_11411,N_10269,N_10061);
nor U11412 (N_11412,N_10809,N_10773);
nand U11413 (N_11413,N_10265,N_10851);
nand U11414 (N_11414,N_10718,N_10876);
nand U11415 (N_11415,N_10063,N_10399);
or U11416 (N_11416,N_10306,N_10797);
nor U11417 (N_11417,N_10759,N_10158);
nor U11418 (N_11418,N_10001,N_10438);
and U11419 (N_11419,N_10887,N_10579);
nand U11420 (N_11420,N_10552,N_10606);
xor U11421 (N_11421,N_10712,N_10272);
nand U11422 (N_11422,N_10643,N_10808);
or U11423 (N_11423,N_10825,N_10661);
nand U11424 (N_11424,N_10023,N_10510);
or U11425 (N_11425,N_10507,N_10355);
or U11426 (N_11426,N_10477,N_10471);
xnor U11427 (N_11427,N_10896,N_10557);
nand U11428 (N_11428,N_10524,N_10124);
nand U11429 (N_11429,N_10884,N_10041);
nand U11430 (N_11430,N_10363,N_10397);
xnor U11431 (N_11431,N_10819,N_10078);
nor U11432 (N_11432,N_10843,N_10180);
nand U11433 (N_11433,N_10762,N_10091);
nor U11434 (N_11434,N_10075,N_10640);
nand U11435 (N_11435,N_10542,N_10101);
nor U11436 (N_11436,N_10730,N_10442);
and U11437 (N_11437,N_10556,N_10377);
and U11438 (N_11438,N_10104,N_10668);
xnor U11439 (N_11439,N_10986,N_10145);
xor U11440 (N_11440,N_10501,N_10203);
xnor U11441 (N_11441,N_10958,N_10233);
or U11442 (N_11442,N_10889,N_10629);
or U11443 (N_11443,N_10649,N_10673);
or U11444 (N_11444,N_10344,N_10633);
or U11445 (N_11445,N_10183,N_10569);
nand U11446 (N_11446,N_10901,N_10655);
nor U11447 (N_11447,N_10196,N_10914);
or U11448 (N_11448,N_10691,N_10503);
and U11449 (N_11449,N_10325,N_10152);
and U11450 (N_11450,N_10772,N_10352);
and U11451 (N_11451,N_10636,N_10619);
xor U11452 (N_11452,N_10792,N_10647);
nor U11453 (N_11453,N_10115,N_10200);
nor U11454 (N_11454,N_10826,N_10570);
or U11455 (N_11455,N_10996,N_10423);
nor U11456 (N_11456,N_10170,N_10624);
and U11457 (N_11457,N_10869,N_10563);
and U11458 (N_11458,N_10993,N_10815);
or U11459 (N_11459,N_10321,N_10131);
xor U11460 (N_11460,N_10941,N_10056);
xor U11461 (N_11461,N_10310,N_10270);
and U11462 (N_11462,N_10420,N_10599);
nor U11463 (N_11463,N_10480,N_10129);
and U11464 (N_11464,N_10468,N_10789);
and U11465 (N_11465,N_10702,N_10374);
nor U11466 (N_11466,N_10132,N_10427);
or U11467 (N_11467,N_10766,N_10764);
and U11468 (N_11468,N_10980,N_10521);
and U11469 (N_11469,N_10927,N_10714);
and U11470 (N_11470,N_10601,N_10245);
nor U11471 (N_11471,N_10782,N_10518);
and U11472 (N_11472,N_10778,N_10065);
and U11473 (N_11473,N_10657,N_10839);
nand U11474 (N_11474,N_10205,N_10595);
or U11475 (N_11475,N_10008,N_10433);
nor U11476 (N_11476,N_10307,N_10999);
xnor U11477 (N_11477,N_10513,N_10874);
or U11478 (N_11478,N_10068,N_10733);
nand U11479 (N_11479,N_10070,N_10734);
or U11480 (N_11480,N_10925,N_10153);
xor U11481 (N_11481,N_10505,N_10753);
and U11482 (N_11482,N_10871,N_10707);
or U11483 (N_11483,N_10728,N_10166);
xnor U11484 (N_11484,N_10853,N_10088);
xnor U11485 (N_11485,N_10849,N_10535);
nor U11486 (N_11486,N_10452,N_10038);
nand U11487 (N_11487,N_10337,N_10830);
and U11488 (N_11488,N_10459,N_10303);
nand U11489 (N_11489,N_10904,N_10421);
or U11490 (N_11490,N_10544,N_10244);
and U11491 (N_11491,N_10394,N_10110);
xor U11492 (N_11492,N_10143,N_10652);
or U11493 (N_11493,N_10349,N_10027);
nor U11494 (N_11494,N_10872,N_10845);
and U11495 (N_11495,N_10711,N_10937);
nand U11496 (N_11496,N_10140,N_10538);
nand U11497 (N_11497,N_10108,N_10848);
nor U11498 (N_11498,N_10259,N_10135);
nand U11499 (N_11499,N_10030,N_10917);
nand U11500 (N_11500,N_10874,N_10379);
nand U11501 (N_11501,N_10085,N_10333);
xor U11502 (N_11502,N_10776,N_10963);
or U11503 (N_11503,N_10655,N_10672);
and U11504 (N_11504,N_10760,N_10064);
nor U11505 (N_11505,N_10692,N_10154);
nor U11506 (N_11506,N_10018,N_10835);
xnor U11507 (N_11507,N_10291,N_10562);
xnor U11508 (N_11508,N_10082,N_10736);
xor U11509 (N_11509,N_10999,N_10029);
nor U11510 (N_11510,N_10951,N_10634);
nor U11511 (N_11511,N_10542,N_10129);
nor U11512 (N_11512,N_10349,N_10845);
and U11513 (N_11513,N_10276,N_10500);
and U11514 (N_11514,N_10943,N_10533);
nor U11515 (N_11515,N_10309,N_10350);
or U11516 (N_11516,N_10166,N_10542);
nor U11517 (N_11517,N_10087,N_10663);
nor U11518 (N_11518,N_10280,N_10015);
and U11519 (N_11519,N_10141,N_10365);
and U11520 (N_11520,N_10353,N_10768);
or U11521 (N_11521,N_10329,N_10292);
nor U11522 (N_11522,N_10366,N_10666);
nand U11523 (N_11523,N_10607,N_10760);
nor U11524 (N_11524,N_10342,N_10054);
xnor U11525 (N_11525,N_10532,N_10602);
nor U11526 (N_11526,N_10741,N_10806);
and U11527 (N_11527,N_10605,N_10785);
xnor U11528 (N_11528,N_10842,N_10203);
nand U11529 (N_11529,N_10439,N_10909);
xnor U11530 (N_11530,N_10292,N_10686);
nand U11531 (N_11531,N_10803,N_10095);
or U11532 (N_11532,N_10713,N_10824);
xor U11533 (N_11533,N_10405,N_10392);
nand U11534 (N_11534,N_10683,N_10467);
nor U11535 (N_11535,N_10839,N_10759);
or U11536 (N_11536,N_10412,N_10172);
and U11537 (N_11537,N_10264,N_10758);
xnor U11538 (N_11538,N_10723,N_10319);
nor U11539 (N_11539,N_10689,N_10782);
xor U11540 (N_11540,N_10306,N_10104);
or U11541 (N_11541,N_10836,N_10426);
nor U11542 (N_11542,N_10903,N_10081);
xnor U11543 (N_11543,N_10728,N_10239);
nand U11544 (N_11544,N_10669,N_10810);
nand U11545 (N_11545,N_10062,N_10963);
xnor U11546 (N_11546,N_10922,N_10378);
or U11547 (N_11547,N_10578,N_10561);
or U11548 (N_11548,N_10312,N_10065);
and U11549 (N_11549,N_10631,N_10316);
and U11550 (N_11550,N_10016,N_10380);
or U11551 (N_11551,N_10529,N_10719);
xnor U11552 (N_11552,N_10441,N_10744);
nor U11553 (N_11553,N_10117,N_10252);
or U11554 (N_11554,N_10872,N_10667);
xor U11555 (N_11555,N_10543,N_10503);
nor U11556 (N_11556,N_10279,N_10746);
nor U11557 (N_11557,N_10316,N_10394);
or U11558 (N_11558,N_10802,N_10969);
xnor U11559 (N_11559,N_10498,N_10919);
nor U11560 (N_11560,N_10199,N_10375);
nor U11561 (N_11561,N_10785,N_10555);
xnor U11562 (N_11562,N_10070,N_10643);
nor U11563 (N_11563,N_10946,N_10076);
xnor U11564 (N_11564,N_10186,N_10574);
xnor U11565 (N_11565,N_10570,N_10262);
nor U11566 (N_11566,N_10931,N_10064);
or U11567 (N_11567,N_10345,N_10927);
nand U11568 (N_11568,N_10564,N_10137);
nor U11569 (N_11569,N_10386,N_10298);
or U11570 (N_11570,N_10100,N_10290);
xnor U11571 (N_11571,N_10521,N_10392);
nand U11572 (N_11572,N_10859,N_10226);
nor U11573 (N_11573,N_10721,N_10500);
xor U11574 (N_11574,N_10034,N_10300);
or U11575 (N_11575,N_10074,N_10053);
nand U11576 (N_11576,N_10553,N_10429);
or U11577 (N_11577,N_10620,N_10921);
and U11578 (N_11578,N_10030,N_10833);
xnor U11579 (N_11579,N_10653,N_10966);
xor U11580 (N_11580,N_10902,N_10484);
xor U11581 (N_11581,N_10965,N_10451);
or U11582 (N_11582,N_10771,N_10566);
nand U11583 (N_11583,N_10690,N_10071);
and U11584 (N_11584,N_10032,N_10831);
xnor U11585 (N_11585,N_10135,N_10710);
or U11586 (N_11586,N_10027,N_10798);
or U11587 (N_11587,N_10269,N_10978);
xnor U11588 (N_11588,N_10296,N_10366);
nand U11589 (N_11589,N_10089,N_10211);
xor U11590 (N_11590,N_10182,N_10743);
xor U11591 (N_11591,N_10958,N_10466);
or U11592 (N_11592,N_10899,N_10164);
nor U11593 (N_11593,N_10180,N_10656);
nand U11594 (N_11594,N_10407,N_10990);
xor U11595 (N_11595,N_10805,N_10712);
xnor U11596 (N_11596,N_10871,N_10599);
nand U11597 (N_11597,N_10473,N_10438);
or U11598 (N_11598,N_10073,N_10572);
nand U11599 (N_11599,N_10392,N_10906);
nand U11600 (N_11600,N_10804,N_10494);
nand U11601 (N_11601,N_10440,N_10866);
and U11602 (N_11602,N_10567,N_10401);
nor U11603 (N_11603,N_10124,N_10207);
nand U11604 (N_11604,N_10430,N_10988);
xnor U11605 (N_11605,N_10345,N_10850);
nor U11606 (N_11606,N_10098,N_10124);
nand U11607 (N_11607,N_10177,N_10778);
nand U11608 (N_11608,N_10679,N_10766);
and U11609 (N_11609,N_10868,N_10242);
and U11610 (N_11610,N_10296,N_10722);
and U11611 (N_11611,N_10131,N_10878);
nor U11612 (N_11612,N_10284,N_10314);
or U11613 (N_11613,N_10484,N_10434);
xor U11614 (N_11614,N_10544,N_10122);
xnor U11615 (N_11615,N_10696,N_10348);
nor U11616 (N_11616,N_10417,N_10982);
and U11617 (N_11617,N_10123,N_10210);
xnor U11618 (N_11618,N_10928,N_10563);
nand U11619 (N_11619,N_10307,N_10819);
nand U11620 (N_11620,N_10047,N_10790);
and U11621 (N_11621,N_10578,N_10952);
nand U11622 (N_11622,N_10908,N_10728);
and U11623 (N_11623,N_10302,N_10166);
xor U11624 (N_11624,N_10888,N_10389);
nor U11625 (N_11625,N_10006,N_10341);
nand U11626 (N_11626,N_10555,N_10384);
or U11627 (N_11627,N_10355,N_10653);
xor U11628 (N_11628,N_10590,N_10265);
nand U11629 (N_11629,N_10219,N_10494);
or U11630 (N_11630,N_10610,N_10131);
nand U11631 (N_11631,N_10526,N_10929);
and U11632 (N_11632,N_10838,N_10466);
or U11633 (N_11633,N_10710,N_10822);
and U11634 (N_11634,N_10994,N_10707);
and U11635 (N_11635,N_10200,N_10970);
xor U11636 (N_11636,N_10859,N_10697);
nor U11637 (N_11637,N_10959,N_10962);
xor U11638 (N_11638,N_10052,N_10621);
and U11639 (N_11639,N_10118,N_10459);
xor U11640 (N_11640,N_10465,N_10289);
or U11641 (N_11641,N_10386,N_10958);
xnor U11642 (N_11642,N_10469,N_10071);
or U11643 (N_11643,N_10929,N_10975);
and U11644 (N_11644,N_10812,N_10767);
xor U11645 (N_11645,N_10200,N_10071);
xor U11646 (N_11646,N_10348,N_10730);
xor U11647 (N_11647,N_10021,N_10659);
xnor U11648 (N_11648,N_10535,N_10370);
or U11649 (N_11649,N_10506,N_10195);
and U11650 (N_11650,N_10604,N_10867);
xor U11651 (N_11651,N_10391,N_10593);
xor U11652 (N_11652,N_10307,N_10682);
or U11653 (N_11653,N_10347,N_10503);
and U11654 (N_11654,N_10111,N_10526);
nand U11655 (N_11655,N_10128,N_10511);
or U11656 (N_11656,N_10329,N_10888);
or U11657 (N_11657,N_10402,N_10850);
or U11658 (N_11658,N_10726,N_10369);
and U11659 (N_11659,N_10996,N_10605);
or U11660 (N_11660,N_10000,N_10297);
and U11661 (N_11661,N_10676,N_10708);
or U11662 (N_11662,N_10765,N_10797);
xnor U11663 (N_11663,N_10277,N_10157);
nor U11664 (N_11664,N_10257,N_10441);
and U11665 (N_11665,N_10682,N_10135);
and U11666 (N_11666,N_10666,N_10649);
or U11667 (N_11667,N_10694,N_10050);
or U11668 (N_11668,N_10584,N_10957);
and U11669 (N_11669,N_10791,N_10046);
xnor U11670 (N_11670,N_10003,N_10278);
nor U11671 (N_11671,N_10161,N_10285);
xnor U11672 (N_11672,N_10933,N_10069);
nor U11673 (N_11673,N_10354,N_10842);
nor U11674 (N_11674,N_10966,N_10671);
xnor U11675 (N_11675,N_10718,N_10716);
xnor U11676 (N_11676,N_10106,N_10055);
nor U11677 (N_11677,N_10102,N_10283);
nand U11678 (N_11678,N_10681,N_10730);
nor U11679 (N_11679,N_10650,N_10997);
nor U11680 (N_11680,N_10889,N_10547);
nor U11681 (N_11681,N_10795,N_10401);
nand U11682 (N_11682,N_10086,N_10383);
xor U11683 (N_11683,N_10411,N_10369);
and U11684 (N_11684,N_10019,N_10304);
and U11685 (N_11685,N_10445,N_10672);
or U11686 (N_11686,N_10952,N_10305);
or U11687 (N_11687,N_10067,N_10261);
or U11688 (N_11688,N_10490,N_10575);
or U11689 (N_11689,N_10925,N_10979);
xnor U11690 (N_11690,N_10104,N_10143);
or U11691 (N_11691,N_10015,N_10335);
nand U11692 (N_11692,N_10757,N_10904);
and U11693 (N_11693,N_10370,N_10734);
nor U11694 (N_11694,N_10811,N_10927);
nand U11695 (N_11695,N_10661,N_10852);
nor U11696 (N_11696,N_10616,N_10768);
nand U11697 (N_11697,N_10620,N_10728);
or U11698 (N_11698,N_10252,N_10247);
nor U11699 (N_11699,N_10472,N_10858);
nor U11700 (N_11700,N_10590,N_10480);
and U11701 (N_11701,N_10295,N_10829);
nand U11702 (N_11702,N_10632,N_10459);
nor U11703 (N_11703,N_10411,N_10846);
nand U11704 (N_11704,N_10629,N_10436);
nor U11705 (N_11705,N_10862,N_10045);
nor U11706 (N_11706,N_10658,N_10810);
xnor U11707 (N_11707,N_10760,N_10498);
or U11708 (N_11708,N_10680,N_10541);
and U11709 (N_11709,N_10953,N_10489);
and U11710 (N_11710,N_10105,N_10060);
or U11711 (N_11711,N_10418,N_10306);
nor U11712 (N_11712,N_10379,N_10481);
and U11713 (N_11713,N_10512,N_10445);
or U11714 (N_11714,N_10207,N_10331);
nor U11715 (N_11715,N_10730,N_10978);
or U11716 (N_11716,N_10600,N_10553);
nand U11717 (N_11717,N_10012,N_10263);
xor U11718 (N_11718,N_10322,N_10751);
or U11719 (N_11719,N_10959,N_10969);
nor U11720 (N_11720,N_10040,N_10961);
nand U11721 (N_11721,N_10103,N_10752);
nor U11722 (N_11722,N_10961,N_10225);
xnor U11723 (N_11723,N_10069,N_10755);
xor U11724 (N_11724,N_10536,N_10847);
nor U11725 (N_11725,N_10078,N_10757);
and U11726 (N_11726,N_10107,N_10730);
and U11727 (N_11727,N_10153,N_10676);
nand U11728 (N_11728,N_10288,N_10217);
and U11729 (N_11729,N_10795,N_10529);
xor U11730 (N_11730,N_10166,N_10026);
nand U11731 (N_11731,N_10765,N_10949);
or U11732 (N_11732,N_10176,N_10777);
nor U11733 (N_11733,N_10720,N_10253);
xnor U11734 (N_11734,N_10226,N_10531);
nand U11735 (N_11735,N_10175,N_10137);
nand U11736 (N_11736,N_10813,N_10063);
nor U11737 (N_11737,N_10564,N_10494);
nand U11738 (N_11738,N_10839,N_10945);
xor U11739 (N_11739,N_10602,N_10396);
or U11740 (N_11740,N_10155,N_10518);
or U11741 (N_11741,N_10563,N_10492);
nor U11742 (N_11742,N_10248,N_10768);
xor U11743 (N_11743,N_10154,N_10319);
nor U11744 (N_11744,N_10901,N_10554);
and U11745 (N_11745,N_10426,N_10629);
nand U11746 (N_11746,N_10740,N_10824);
xor U11747 (N_11747,N_10838,N_10181);
xor U11748 (N_11748,N_10234,N_10441);
nand U11749 (N_11749,N_10394,N_10498);
xnor U11750 (N_11750,N_10516,N_10610);
and U11751 (N_11751,N_10324,N_10868);
and U11752 (N_11752,N_10588,N_10170);
nand U11753 (N_11753,N_10631,N_10741);
nand U11754 (N_11754,N_10147,N_10307);
or U11755 (N_11755,N_10357,N_10856);
xnor U11756 (N_11756,N_10524,N_10648);
nand U11757 (N_11757,N_10141,N_10870);
nor U11758 (N_11758,N_10883,N_10287);
nand U11759 (N_11759,N_10019,N_10731);
nand U11760 (N_11760,N_10709,N_10266);
xnor U11761 (N_11761,N_10861,N_10065);
nand U11762 (N_11762,N_10075,N_10363);
nor U11763 (N_11763,N_10719,N_10754);
nor U11764 (N_11764,N_10198,N_10894);
nand U11765 (N_11765,N_10900,N_10047);
or U11766 (N_11766,N_10377,N_10820);
xnor U11767 (N_11767,N_10459,N_10606);
and U11768 (N_11768,N_10964,N_10087);
nor U11769 (N_11769,N_10248,N_10904);
xor U11770 (N_11770,N_10953,N_10334);
or U11771 (N_11771,N_10453,N_10957);
nand U11772 (N_11772,N_10968,N_10198);
xnor U11773 (N_11773,N_10340,N_10147);
nor U11774 (N_11774,N_10180,N_10339);
or U11775 (N_11775,N_10408,N_10758);
or U11776 (N_11776,N_10426,N_10724);
nor U11777 (N_11777,N_10245,N_10911);
and U11778 (N_11778,N_10167,N_10339);
nand U11779 (N_11779,N_10532,N_10488);
and U11780 (N_11780,N_10970,N_10012);
or U11781 (N_11781,N_10899,N_10194);
or U11782 (N_11782,N_10870,N_10411);
nand U11783 (N_11783,N_10072,N_10297);
xor U11784 (N_11784,N_10498,N_10726);
nand U11785 (N_11785,N_10336,N_10056);
or U11786 (N_11786,N_10682,N_10253);
and U11787 (N_11787,N_10196,N_10863);
or U11788 (N_11788,N_10917,N_10104);
or U11789 (N_11789,N_10422,N_10625);
xor U11790 (N_11790,N_10882,N_10931);
and U11791 (N_11791,N_10340,N_10361);
nor U11792 (N_11792,N_10421,N_10367);
and U11793 (N_11793,N_10418,N_10673);
nand U11794 (N_11794,N_10011,N_10585);
and U11795 (N_11795,N_10537,N_10322);
nand U11796 (N_11796,N_10079,N_10040);
nor U11797 (N_11797,N_10257,N_10755);
and U11798 (N_11798,N_10972,N_10748);
and U11799 (N_11799,N_10696,N_10936);
nor U11800 (N_11800,N_10155,N_10616);
nor U11801 (N_11801,N_10712,N_10810);
or U11802 (N_11802,N_10393,N_10529);
nand U11803 (N_11803,N_10162,N_10894);
nand U11804 (N_11804,N_10468,N_10687);
or U11805 (N_11805,N_10298,N_10388);
xor U11806 (N_11806,N_10930,N_10648);
or U11807 (N_11807,N_10791,N_10299);
and U11808 (N_11808,N_10240,N_10289);
or U11809 (N_11809,N_10907,N_10019);
and U11810 (N_11810,N_10494,N_10892);
nand U11811 (N_11811,N_10626,N_10995);
nor U11812 (N_11812,N_10867,N_10840);
xor U11813 (N_11813,N_10356,N_10018);
nand U11814 (N_11814,N_10616,N_10314);
or U11815 (N_11815,N_10122,N_10373);
nor U11816 (N_11816,N_10183,N_10672);
or U11817 (N_11817,N_10467,N_10325);
and U11818 (N_11818,N_10885,N_10470);
and U11819 (N_11819,N_10418,N_10067);
nand U11820 (N_11820,N_10985,N_10770);
and U11821 (N_11821,N_10773,N_10970);
and U11822 (N_11822,N_10541,N_10566);
and U11823 (N_11823,N_10441,N_10309);
or U11824 (N_11824,N_10924,N_10623);
or U11825 (N_11825,N_10241,N_10323);
and U11826 (N_11826,N_10104,N_10940);
nor U11827 (N_11827,N_10215,N_10838);
nor U11828 (N_11828,N_10822,N_10266);
and U11829 (N_11829,N_10899,N_10724);
nor U11830 (N_11830,N_10021,N_10259);
and U11831 (N_11831,N_10459,N_10841);
or U11832 (N_11832,N_10476,N_10341);
xnor U11833 (N_11833,N_10459,N_10314);
nand U11834 (N_11834,N_10086,N_10682);
and U11835 (N_11835,N_10457,N_10721);
nand U11836 (N_11836,N_10323,N_10360);
nor U11837 (N_11837,N_10430,N_10802);
and U11838 (N_11838,N_10613,N_10097);
nand U11839 (N_11839,N_10400,N_10994);
or U11840 (N_11840,N_10859,N_10557);
nor U11841 (N_11841,N_10985,N_10781);
nand U11842 (N_11842,N_10020,N_10381);
xnor U11843 (N_11843,N_10190,N_10081);
nand U11844 (N_11844,N_10393,N_10255);
nand U11845 (N_11845,N_10764,N_10621);
nand U11846 (N_11846,N_10759,N_10587);
and U11847 (N_11847,N_10842,N_10342);
and U11848 (N_11848,N_10680,N_10677);
nand U11849 (N_11849,N_10476,N_10509);
xor U11850 (N_11850,N_10345,N_10538);
nor U11851 (N_11851,N_10347,N_10626);
nor U11852 (N_11852,N_10453,N_10412);
nand U11853 (N_11853,N_10167,N_10071);
or U11854 (N_11854,N_10257,N_10855);
and U11855 (N_11855,N_10473,N_10268);
and U11856 (N_11856,N_10673,N_10346);
or U11857 (N_11857,N_10822,N_10943);
or U11858 (N_11858,N_10279,N_10732);
xor U11859 (N_11859,N_10514,N_10901);
or U11860 (N_11860,N_10180,N_10142);
and U11861 (N_11861,N_10924,N_10902);
or U11862 (N_11862,N_10963,N_10166);
or U11863 (N_11863,N_10587,N_10641);
nor U11864 (N_11864,N_10032,N_10494);
nor U11865 (N_11865,N_10063,N_10670);
nor U11866 (N_11866,N_10537,N_10438);
nor U11867 (N_11867,N_10919,N_10064);
xnor U11868 (N_11868,N_10547,N_10655);
and U11869 (N_11869,N_10469,N_10204);
nand U11870 (N_11870,N_10689,N_10108);
xnor U11871 (N_11871,N_10546,N_10710);
and U11872 (N_11872,N_10494,N_10738);
nor U11873 (N_11873,N_10768,N_10961);
xnor U11874 (N_11874,N_10689,N_10648);
nand U11875 (N_11875,N_10721,N_10239);
nand U11876 (N_11876,N_10320,N_10997);
nand U11877 (N_11877,N_10761,N_10016);
nor U11878 (N_11878,N_10250,N_10184);
and U11879 (N_11879,N_10643,N_10677);
nor U11880 (N_11880,N_10665,N_10738);
nor U11881 (N_11881,N_10841,N_10040);
nand U11882 (N_11882,N_10653,N_10980);
or U11883 (N_11883,N_10772,N_10456);
and U11884 (N_11884,N_10586,N_10668);
nor U11885 (N_11885,N_10390,N_10890);
and U11886 (N_11886,N_10848,N_10587);
and U11887 (N_11887,N_10024,N_10295);
nor U11888 (N_11888,N_10119,N_10744);
nor U11889 (N_11889,N_10670,N_10384);
xor U11890 (N_11890,N_10000,N_10531);
nand U11891 (N_11891,N_10102,N_10929);
nand U11892 (N_11892,N_10361,N_10294);
and U11893 (N_11893,N_10166,N_10593);
nand U11894 (N_11894,N_10138,N_10612);
or U11895 (N_11895,N_10198,N_10749);
or U11896 (N_11896,N_10665,N_10395);
or U11897 (N_11897,N_10252,N_10721);
nor U11898 (N_11898,N_10431,N_10989);
and U11899 (N_11899,N_10008,N_10149);
nand U11900 (N_11900,N_10853,N_10626);
nor U11901 (N_11901,N_10446,N_10271);
or U11902 (N_11902,N_10816,N_10544);
and U11903 (N_11903,N_10856,N_10965);
and U11904 (N_11904,N_10679,N_10172);
or U11905 (N_11905,N_10818,N_10785);
nand U11906 (N_11906,N_10208,N_10385);
xor U11907 (N_11907,N_10602,N_10597);
nor U11908 (N_11908,N_10876,N_10030);
xnor U11909 (N_11909,N_10971,N_10489);
or U11910 (N_11910,N_10194,N_10002);
and U11911 (N_11911,N_10659,N_10604);
nand U11912 (N_11912,N_10749,N_10041);
nor U11913 (N_11913,N_10455,N_10358);
or U11914 (N_11914,N_10409,N_10921);
nand U11915 (N_11915,N_10838,N_10273);
or U11916 (N_11916,N_10634,N_10694);
xnor U11917 (N_11917,N_10981,N_10856);
and U11918 (N_11918,N_10920,N_10507);
xor U11919 (N_11919,N_10683,N_10240);
nor U11920 (N_11920,N_10608,N_10626);
or U11921 (N_11921,N_10602,N_10239);
or U11922 (N_11922,N_10057,N_10226);
nand U11923 (N_11923,N_10912,N_10669);
nor U11924 (N_11924,N_10847,N_10699);
nor U11925 (N_11925,N_10505,N_10540);
nor U11926 (N_11926,N_10739,N_10175);
xnor U11927 (N_11927,N_10548,N_10868);
and U11928 (N_11928,N_10510,N_10555);
xnor U11929 (N_11929,N_10396,N_10184);
xor U11930 (N_11930,N_10223,N_10204);
xor U11931 (N_11931,N_10062,N_10889);
nand U11932 (N_11932,N_10630,N_10351);
and U11933 (N_11933,N_10512,N_10532);
or U11934 (N_11934,N_10855,N_10623);
nor U11935 (N_11935,N_10455,N_10355);
and U11936 (N_11936,N_10109,N_10140);
nand U11937 (N_11937,N_10114,N_10786);
xnor U11938 (N_11938,N_10823,N_10897);
xor U11939 (N_11939,N_10271,N_10557);
nand U11940 (N_11940,N_10590,N_10091);
nor U11941 (N_11941,N_10837,N_10900);
nand U11942 (N_11942,N_10581,N_10496);
nor U11943 (N_11943,N_10783,N_10341);
nand U11944 (N_11944,N_10559,N_10195);
or U11945 (N_11945,N_10519,N_10800);
or U11946 (N_11946,N_10759,N_10445);
and U11947 (N_11947,N_10783,N_10511);
nand U11948 (N_11948,N_10330,N_10575);
xnor U11949 (N_11949,N_10139,N_10181);
xor U11950 (N_11950,N_10532,N_10004);
nand U11951 (N_11951,N_10859,N_10524);
xor U11952 (N_11952,N_10388,N_10129);
and U11953 (N_11953,N_10053,N_10190);
xnor U11954 (N_11954,N_10354,N_10516);
or U11955 (N_11955,N_10094,N_10760);
xnor U11956 (N_11956,N_10830,N_10924);
or U11957 (N_11957,N_10057,N_10213);
or U11958 (N_11958,N_10367,N_10610);
xnor U11959 (N_11959,N_10311,N_10506);
or U11960 (N_11960,N_10156,N_10004);
nor U11961 (N_11961,N_10818,N_10145);
nand U11962 (N_11962,N_10365,N_10717);
or U11963 (N_11963,N_10976,N_10503);
or U11964 (N_11964,N_10912,N_10751);
and U11965 (N_11965,N_10862,N_10072);
xnor U11966 (N_11966,N_10955,N_10833);
nand U11967 (N_11967,N_10047,N_10427);
or U11968 (N_11968,N_10296,N_10225);
xor U11969 (N_11969,N_10507,N_10209);
xor U11970 (N_11970,N_10226,N_10581);
nor U11971 (N_11971,N_10536,N_10370);
xor U11972 (N_11972,N_10751,N_10458);
nor U11973 (N_11973,N_10601,N_10044);
or U11974 (N_11974,N_10039,N_10235);
xor U11975 (N_11975,N_10717,N_10010);
nor U11976 (N_11976,N_10735,N_10061);
and U11977 (N_11977,N_10266,N_10150);
and U11978 (N_11978,N_10561,N_10369);
xnor U11979 (N_11979,N_10604,N_10022);
or U11980 (N_11980,N_10275,N_10490);
xor U11981 (N_11981,N_10323,N_10320);
nand U11982 (N_11982,N_10110,N_10199);
xnor U11983 (N_11983,N_10359,N_10566);
or U11984 (N_11984,N_10861,N_10833);
xnor U11985 (N_11985,N_10423,N_10578);
nor U11986 (N_11986,N_10006,N_10384);
xnor U11987 (N_11987,N_10724,N_10731);
nand U11988 (N_11988,N_10715,N_10198);
xnor U11989 (N_11989,N_10233,N_10204);
xnor U11990 (N_11990,N_10474,N_10121);
nand U11991 (N_11991,N_10592,N_10738);
nor U11992 (N_11992,N_10886,N_10378);
and U11993 (N_11993,N_10828,N_10111);
nand U11994 (N_11994,N_10630,N_10763);
nand U11995 (N_11995,N_10881,N_10679);
nand U11996 (N_11996,N_10347,N_10981);
and U11997 (N_11997,N_10628,N_10069);
and U11998 (N_11998,N_10510,N_10503);
or U11999 (N_11999,N_10882,N_10936);
and U12000 (N_12000,N_11105,N_11199);
nor U12001 (N_12001,N_11760,N_11115);
and U12002 (N_12002,N_11797,N_11129);
and U12003 (N_12003,N_11877,N_11252);
nand U12004 (N_12004,N_11694,N_11064);
nand U12005 (N_12005,N_11516,N_11088);
nand U12006 (N_12006,N_11791,N_11518);
xnor U12007 (N_12007,N_11764,N_11122);
xor U12008 (N_12008,N_11986,N_11261);
xnor U12009 (N_12009,N_11159,N_11809);
nor U12010 (N_12010,N_11511,N_11755);
or U12011 (N_12011,N_11557,N_11651);
nand U12012 (N_12012,N_11433,N_11234);
nand U12013 (N_12013,N_11905,N_11412);
or U12014 (N_12014,N_11339,N_11533);
or U12015 (N_12015,N_11928,N_11155);
nand U12016 (N_12016,N_11019,N_11883);
nand U12017 (N_12017,N_11524,N_11272);
nor U12018 (N_12018,N_11571,N_11202);
or U12019 (N_12019,N_11145,N_11930);
or U12020 (N_12020,N_11157,N_11648);
nor U12021 (N_12021,N_11285,N_11506);
or U12022 (N_12022,N_11204,N_11615);
xnor U12023 (N_12023,N_11074,N_11871);
or U12024 (N_12024,N_11832,N_11778);
and U12025 (N_12025,N_11484,N_11772);
xnor U12026 (N_12026,N_11513,N_11885);
nor U12027 (N_12027,N_11825,N_11711);
and U12028 (N_12028,N_11971,N_11927);
nand U12029 (N_12029,N_11320,N_11593);
nand U12030 (N_12030,N_11283,N_11109);
or U12031 (N_12031,N_11439,N_11813);
nand U12032 (N_12032,N_11541,N_11025);
nor U12033 (N_12033,N_11034,N_11999);
xnor U12034 (N_12034,N_11340,N_11017);
xor U12035 (N_12035,N_11162,N_11287);
or U12036 (N_12036,N_11539,N_11676);
nor U12037 (N_12037,N_11512,N_11151);
nand U12038 (N_12038,N_11842,N_11410);
nand U12039 (N_12039,N_11085,N_11112);
nor U12040 (N_12040,N_11914,N_11800);
xnor U12041 (N_12041,N_11787,N_11841);
nand U12042 (N_12042,N_11701,N_11814);
nand U12043 (N_12043,N_11087,N_11812);
xnor U12044 (N_12044,N_11881,N_11070);
nand U12045 (N_12045,N_11917,N_11544);
nor U12046 (N_12046,N_11035,N_11817);
xor U12047 (N_12047,N_11644,N_11780);
nand U12048 (N_12048,N_11414,N_11464);
nor U12049 (N_12049,N_11437,N_11231);
or U12050 (N_12050,N_11203,N_11373);
xor U12051 (N_12051,N_11100,N_11956);
xnor U12052 (N_12052,N_11688,N_11063);
and U12053 (N_12053,N_11251,N_11700);
xnor U12054 (N_12054,N_11384,N_11417);
nand U12055 (N_12055,N_11776,N_11564);
or U12056 (N_12056,N_11292,N_11096);
or U12057 (N_12057,N_11654,N_11879);
or U12058 (N_12058,N_11818,N_11808);
xor U12059 (N_12059,N_11200,N_11635);
nand U12060 (N_12060,N_11582,N_11728);
nor U12061 (N_12061,N_11893,N_11827);
nor U12062 (N_12062,N_11041,N_11628);
nand U12063 (N_12063,N_11387,N_11121);
xnor U12064 (N_12064,N_11233,N_11845);
xor U12065 (N_12065,N_11829,N_11055);
xor U12066 (N_12066,N_11084,N_11784);
xnor U12067 (N_12067,N_11349,N_11972);
and U12068 (N_12068,N_11163,N_11957);
nor U12069 (N_12069,N_11048,N_11082);
xnor U12070 (N_12070,N_11196,N_11678);
nand U12071 (N_12071,N_11996,N_11907);
and U12072 (N_12072,N_11699,N_11527);
or U12073 (N_12073,N_11172,N_11781);
nor U12074 (N_12074,N_11810,N_11566);
or U12075 (N_12075,N_11482,N_11355);
and U12076 (N_12076,N_11762,N_11835);
or U12077 (N_12077,N_11455,N_11021);
xor U12078 (N_12078,N_11898,N_11480);
or U12079 (N_12079,N_11449,N_11395);
xnor U12080 (N_12080,N_11529,N_11941);
and U12081 (N_12081,N_11418,N_11993);
or U12082 (N_12082,N_11794,N_11696);
or U12083 (N_12083,N_11577,N_11614);
nand U12084 (N_12084,N_11719,N_11337);
nor U12085 (N_12085,N_11868,N_11773);
xnor U12086 (N_12086,N_11193,N_11637);
xnor U12087 (N_12087,N_11580,N_11168);
or U12088 (N_12088,N_11618,N_11771);
xnor U12089 (N_12089,N_11232,N_11132);
xor U12090 (N_12090,N_11515,N_11954);
or U12091 (N_12091,N_11627,N_11562);
and U12092 (N_12092,N_11182,N_11592);
xnor U12093 (N_12093,N_11181,N_11785);
or U12094 (N_12094,N_11896,N_11820);
nor U12095 (N_12095,N_11046,N_11262);
nand U12096 (N_12096,N_11360,N_11134);
nor U12097 (N_12097,N_11811,N_11698);
xor U12098 (N_12098,N_11052,N_11989);
and U12099 (N_12099,N_11622,N_11640);
and U12100 (N_12100,N_11265,N_11271);
xnor U12101 (N_12101,N_11729,N_11077);
nor U12102 (N_12102,N_11454,N_11201);
nor U12103 (N_12103,N_11805,N_11542);
and U12104 (N_12104,N_11118,N_11740);
nand U12105 (N_12105,N_11016,N_11596);
or U12106 (N_12106,N_11466,N_11291);
nor U12107 (N_12107,N_11472,N_11369);
or U12108 (N_12108,N_11311,N_11921);
nand U12109 (N_12109,N_11278,N_11469);
xnor U12110 (N_12110,N_11220,N_11419);
nand U12111 (N_12111,N_11668,N_11040);
or U12112 (N_12112,N_11816,N_11943);
nand U12113 (N_12113,N_11844,N_11401);
or U12114 (N_12114,N_11804,N_11894);
or U12115 (N_12115,N_11207,N_11004);
or U12116 (N_12116,N_11236,N_11543);
nand U12117 (N_12117,N_11144,N_11248);
nor U12118 (N_12118,N_11028,N_11938);
and U12119 (N_12119,N_11324,N_11937);
nor U12120 (N_12120,N_11214,N_11803);
xnor U12121 (N_12121,N_11366,N_11370);
xnor U12122 (N_12122,N_11655,N_11742);
nand U12123 (N_12123,N_11448,N_11487);
and U12124 (N_12124,N_11570,N_11951);
and U12125 (N_12125,N_11107,N_11260);
nand U12126 (N_12126,N_11873,N_11522);
or U12127 (N_12127,N_11257,N_11583);
nor U12128 (N_12128,N_11974,N_11409);
xnor U12129 (N_12129,N_11421,N_11225);
or U12130 (N_12130,N_11975,N_11763);
xnor U12131 (N_12131,N_11081,N_11191);
nor U12132 (N_12132,N_11589,N_11884);
xnor U12133 (N_12133,N_11836,N_11576);
nand U12134 (N_12134,N_11607,N_11208);
or U12135 (N_12135,N_11294,N_11826);
and U12136 (N_12136,N_11428,N_11631);
nor U12137 (N_12137,N_11362,N_11058);
nand U12138 (N_12138,N_11978,N_11737);
xor U12139 (N_12139,N_11407,N_11056);
nor U12140 (N_12140,N_11333,N_11237);
nor U12141 (N_12141,N_11602,N_11586);
nand U12142 (N_12142,N_11343,N_11356);
and U12143 (N_12143,N_11766,N_11459);
or U12144 (N_12144,N_11666,N_11377);
and U12145 (N_12145,N_11590,N_11530);
or U12146 (N_12146,N_11749,N_11500);
or U12147 (N_12147,N_11429,N_11652);
nand U12148 (N_12148,N_11397,N_11758);
and U12149 (N_12149,N_11920,N_11347);
nor U12150 (N_12150,N_11940,N_11626);
and U12151 (N_12151,N_11024,N_11682);
and U12152 (N_12152,N_11057,N_11612);
or U12153 (N_12153,N_11065,N_11686);
nand U12154 (N_12154,N_11127,N_11741);
and U12155 (N_12155,N_11315,N_11858);
nor U12156 (N_12156,N_11752,N_11479);
xor U12157 (N_12157,N_11359,N_11504);
xor U12158 (N_12158,N_11317,N_11600);
xnor U12159 (N_12159,N_11910,N_11973);
xnor U12160 (N_12160,N_11069,N_11756);
nor U12161 (N_12161,N_11759,N_11226);
nor U12162 (N_12162,N_11197,N_11657);
and U12163 (N_12163,N_11146,N_11244);
nand U12164 (N_12164,N_11638,N_11367);
or U12165 (N_12165,N_11430,N_11497);
nor U12166 (N_12166,N_11636,N_11344);
and U12167 (N_12167,N_11326,N_11446);
nor U12168 (N_12168,N_11661,N_11662);
nor U12169 (N_12169,N_11492,N_11890);
nor U12170 (N_12170,N_11946,N_11030);
xor U12171 (N_12171,N_11212,N_11258);
and U12172 (N_12172,N_11131,N_11018);
nand U12173 (N_12173,N_11241,N_11388);
nand U12174 (N_12174,N_11866,N_11290);
nand U12175 (N_12175,N_11850,N_11076);
nor U12176 (N_12176,N_11150,N_11789);
nand U12177 (N_12177,N_11922,N_11748);
xnor U12178 (N_12178,N_11286,N_11926);
nand U12179 (N_12179,N_11133,N_11486);
xnor U12180 (N_12180,N_11819,N_11843);
nor U12181 (N_12181,N_11451,N_11059);
xor U12182 (N_12182,N_11381,N_11924);
xor U12183 (N_12183,N_11436,N_11601);
nor U12184 (N_12184,N_11372,N_11350);
nand U12185 (N_12185,N_11086,N_11572);
nand U12186 (N_12186,N_11736,N_11135);
nand U12187 (N_12187,N_11153,N_11323);
and U12188 (N_12188,N_11620,N_11619);
nor U12189 (N_12189,N_11724,N_11945);
or U12190 (N_12190,N_11983,N_11665);
and U12191 (N_12191,N_11867,N_11177);
or U12192 (N_12192,N_11992,N_11495);
xor U12193 (N_12193,N_11870,N_11848);
xor U12194 (N_12194,N_11123,N_11432);
nand U12195 (N_12195,N_11965,N_11806);
nand U12196 (N_12196,N_11379,N_11205);
or U12197 (N_12197,N_11005,N_11083);
nand U12198 (N_12198,N_11009,N_11139);
xnor U12199 (N_12199,N_11739,N_11880);
xor U12200 (N_12200,N_11138,N_11091);
nor U12201 (N_12201,N_11693,N_11610);
and U12202 (N_12202,N_11319,N_11649);
nand U12203 (N_12203,N_11673,N_11213);
nor U12204 (N_12204,N_11282,N_11427);
nor U12205 (N_12205,N_11962,N_11793);
and U12206 (N_12206,N_11659,N_11705);
nor U12207 (N_12207,N_11855,N_11033);
nor U12208 (N_12208,N_11561,N_11392);
or U12209 (N_12209,N_11629,N_11186);
xnor U12210 (N_12210,N_11551,N_11568);
nand U12211 (N_12211,N_11585,N_11802);
and U12212 (N_12212,N_11130,N_11958);
nand U12213 (N_12213,N_11857,N_11253);
nand U12214 (N_12214,N_11066,N_11211);
nor U12215 (N_12215,N_11509,N_11779);
and U12216 (N_12216,N_11221,N_11830);
or U12217 (N_12217,N_11000,N_11476);
and U12218 (N_12218,N_11434,N_11591);
or U12219 (N_12219,N_11488,N_11932);
nand U12220 (N_12220,N_11458,N_11523);
xor U12221 (N_12221,N_11578,N_11243);
nor U12222 (N_12222,N_11695,N_11738);
xor U12223 (N_12223,N_11901,N_11909);
nand U12224 (N_12224,N_11995,N_11703);
nor U12225 (N_12225,N_11833,N_11042);
nor U12226 (N_12226,N_11303,N_11185);
nand U12227 (N_12227,N_11113,N_11308);
nor U12228 (N_12228,N_11939,N_11677);
nand U12229 (N_12229,N_11923,N_11950);
and U12230 (N_12230,N_11936,N_11403);
nand U12231 (N_12231,N_11953,N_11230);
nand U12232 (N_12232,N_11704,N_11330);
and U12233 (N_12233,N_11106,N_11156);
or U12234 (N_12234,N_11672,N_11959);
or U12235 (N_12235,N_11918,N_11273);
or U12236 (N_12236,N_11102,N_11603);
or U12237 (N_12237,N_11908,N_11416);
xor U12238 (N_12238,N_11322,N_11111);
nand U12239 (N_12239,N_11613,N_11475);
xor U12240 (N_12240,N_11117,N_11223);
and U12241 (N_12241,N_11643,N_11616);
nand U12242 (N_12242,N_11535,N_11807);
xor U12243 (N_12243,N_11768,N_11089);
nor U12244 (N_12244,N_11716,N_11148);
or U12245 (N_12245,N_11297,N_11404);
or U12246 (N_12246,N_11167,N_11815);
and U12247 (N_12247,N_11567,N_11663);
nand U12248 (N_12248,N_11653,N_11043);
or U12249 (N_12249,N_11777,N_11534);
xnor U12250 (N_12250,N_11228,N_11702);
or U12251 (N_12251,N_11862,N_11691);
and U12252 (N_12252,N_11264,N_11537);
or U12253 (N_12253,N_11210,N_11517);
or U12254 (N_12254,N_11068,N_11003);
nand U12255 (N_12255,N_11708,N_11667);
xnor U12256 (N_12256,N_11722,N_11865);
nand U12257 (N_12257,N_11119,N_11438);
xnor U12258 (N_12258,N_11423,N_11239);
xor U12259 (N_12259,N_11481,N_11269);
and U12260 (N_12260,N_11948,N_11354);
and U12261 (N_12261,N_11714,N_11465);
and U12262 (N_12262,N_11092,N_11398);
xor U12263 (N_12263,N_11002,N_11011);
nor U12264 (N_12264,N_11987,N_11679);
and U12265 (N_12265,N_11605,N_11067);
and U12266 (N_12266,N_11071,N_11967);
nor U12267 (N_12267,N_11980,N_11413);
and U12268 (N_12268,N_11240,N_11745);
nand U12269 (N_12269,N_11735,N_11604);
nor U12270 (N_12270,N_11249,N_11647);
and U12271 (N_12271,N_11710,N_11934);
xor U12272 (N_12272,N_11621,N_11357);
nand U12273 (N_12273,N_11846,N_11912);
xor U12274 (N_12274,N_11502,N_11963);
nand U12275 (N_12275,N_11094,N_11555);
or U12276 (N_12276,N_11669,N_11284);
or U12277 (N_12277,N_11318,N_11027);
and U12278 (N_12278,N_11770,N_11450);
xnor U12279 (N_12279,N_11425,N_11184);
xnor U12280 (N_12280,N_11942,N_11528);
and U12281 (N_12281,N_11329,N_11888);
or U12282 (N_12282,N_11470,N_11546);
or U12283 (N_12283,N_11097,N_11491);
xnor U12284 (N_12284,N_11723,N_11206);
nor U12285 (N_12285,N_11902,N_11863);
or U12286 (N_12286,N_11494,N_11152);
xnor U12287 (N_12287,N_11180,N_11166);
xor U12288 (N_12288,N_11911,N_11897);
nand U12289 (N_12289,N_11852,N_11720);
or U12290 (N_12290,N_11851,N_11140);
and U12291 (N_12291,N_11020,N_11597);
nand U12292 (N_12292,N_11411,N_11899);
and U12293 (N_12293,N_11903,N_11949);
xor U12294 (N_12294,N_11994,N_11358);
nand U12295 (N_12295,N_11985,N_11933);
nor U12296 (N_12296,N_11161,N_11548);
nor U12297 (N_12297,N_11179,N_11685);
and U12298 (N_12298,N_11242,N_11501);
nand U12299 (N_12299,N_11977,N_11442);
and U12300 (N_12300,N_11692,N_11375);
nand U12301 (N_12301,N_11731,N_11889);
nand U12302 (N_12302,N_11222,N_11374);
nor U12303 (N_12303,N_11821,N_11382);
xnor U12304 (N_12304,N_11733,N_11715);
nor U12305 (N_12305,N_11468,N_11037);
or U12306 (N_12306,N_11219,N_11001);
or U12307 (N_12307,N_11099,N_11431);
and U12308 (N_12308,N_11031,N_11312);
and U12309 (N_12309,N_11051,N_11498);
xnor U12310 (N_12310,N_11141,N_11732);
nor U12311 (N_12311,N_11368,N_11854);
and U12312 (N_12312,N_11964,N_11399);
nand U12313 (N_12313,N_11757,N_11120);
nor U12314 (N_12314,N_11215,N_11514);
nand U12315 (N_12315,N_11010,N_11376);
nand U12316 (N_12316,N_11026,N_11380);
and U12317 (N_12317,N_11961,N_11725);
nand U12318 (N_12318,N_11859,N_11298);
nor U12319 (N_12319,N_11396,N_11520);
or U12320 (N_12320,N_11584,N_11970);
nor U12321 (N_12321,N_11485,N_11108);
and U12322 (N_12322,N_11915,N_11681);
nand U12323 (N_12323,N_11408,N_11050);
xnor U12324 (N_12324,N_11190,N_11183);
nor U12325 (N_12325,N_11378,N_11887);
xnor U12326 (N_12326,N_11435,N_11706);
xor U12327 (N_12327,N_11245,N_11675);
or U12328 (N_12328,N_11875,N_11038);
nor U12329 (N_12329,N_11558,N_11164);
nor U12330 (N_12330,N_11301,N_11327);
nand U12331 (N_12331,N_11878,N_11062);
xor U12332 (N_12332,N_11274,N_11697);
nand U12333 (N_12333,N_11295,N_11095);
nand U12334 (N_12334,N_11982,N_11171);
nor U12335 (N_12335,N_11104,N_11746);
xor U12336 (N_12336,N_11137,N_11683);
nor U12337 (N_12337,N_11952,N_11314);
and U12338 (N_12338,N_11124,N_11633);
nand U12339 (N_12339,N_11554,N_11526);
and U12340 (N_12340,N_11743,N_11856);
nor U12341 (N_12341,N_11402,N_11981);
and U12342 (N_12342,N_11521,N_11801);
nand U12343 (N_12343,N_11300,N_11254);
nor U12344 (N_12344,N_11008,N_11839);
xor U12345 (N_12345,N_11581,N_11727);
nor U12346 (N_12346,N_11462,N_11712);
and U12347 (N_12347,N_11632,N_11767);
nand U12348 (N_12348,N_11642,N_11158);
or U12349 (N_12349,N_11473,N_11641);
and U12350 (N_12350,N_11029,N_11178);
nor U12351 (N_12351,N_11721,N_11840);
xor U12352 (N_12352,N_11707,N_11299);
xor U12353 (N_12353,N_11538,N_11338);
and U12354 (N_12354,N_11049,N_11078);
xor U12355 (N_12355,N_11919,N_11796);
nor U12356 (N_12356,N_11363,N_11828);
or U12357 (N_12357,N_11553,N_11611);
nor U12358 (N_12358,N_11393,N_11080);
xor U12359 (N_12359,N_11467,N_11309);
and U12360 (N_12360,N_11490,N_11391);
xor U12361 (N_12361,N_11900,N_11114);
nor U12362 (N_12362,N_11460,N_11969);
or U12363 (N_12363,N_11255,N_11445);
xnor U12364 (N_12364,N_11718,N_11510);
nor U12365 (N_12365,N_11192,N_11098);
and U12366 (N_12366,N_11276,N_11335);
and U12367 (N_12367,N_11575,N_11457);
or U12368 (N_12368,N_11882,N_11966);
or U12369 (N_12369,N_11302,N_11991);
xnor U12370 (N_12370,N_11559,N_11194);
nor U12371 (N_12371,N_11352,N_11799);
nor U12372 (N_12372,N_11864,N_11054);
nor U12373 (N_12373,N_11047,N_11405);
and U12374 (N_12374,N_11573,N_11861);
or U12375 (N_12375,N_11128,N_11471);
nand U12376 (N_12376,N_11444,N_11147);
or U12377 (N_12377,N_11976,N_11838);
nor U12378 (N_12378,N_11422,N_11594);
or U12379 (N_12379,N_11935,N_11606);
nor U12380 (N_12380,N_11660,N_11493);
and U12381 (N_12381,N_11831,N_11508);
and U12382 (N_12382,N_11783,N_11872);
nand U12383 (N_12383,N_11891,N_11609);
or U12384 (N_12384,N_11307,N_11280);
and U12385 (N_12385,N_11136,N_11288);
nand U12386 (N_12386,N_11406,N_11625);
or U12387 (N_12387,N_11023,N_11342);
xnor U12388 (N_12388,N_11321,N_11012);
nand U12389 (N_12389,N_11126,N_11713);
nand U12390 (N_12390,N_11424,N_11664);
and U12391 (N_12391,N_11990,N_11750);
or U12392 (N_12392,N_11545,N_11540);
xnor U12393 (N_12393,N_11906,N_11014);
or U12394 (N_12394,N_11536,N_11684);
or U12395 (N_12395,N_11947,N_11765);
xnor U12396 (N_12396,N_11658,N_11798);
xor U12397 (N_12397,N_11579,N_11630);
xor U12398 (N_12398,N_11217,N_11170);
and U12399 (N_12399,N_11256,N_11656);
and U12400 (N_12400,N_11519,N_11453);
xnor U12401 (N_12401,N_11569,N_11036);
xnor U12402 (N_12402,N_11726,N_11447);
nor U12403 (N_12403,N_11173,N_11013);
nand U12404 (N_12404,N_11267,N_11400);
xor U12405 (N_12405,N_11925,N_11053);
xor U12406 (N_12406,N_11477,N_11198);
and U12407 (N_12407,N_11525,N_11270);
and U12408 (N_12408,N_11674,N_11503);
or U12409 (N_12409,N_11560,N_11671);
xor U12410 (N_12410,N_11348,N_11929);
nand U12411 (N_12411,N_11823,N_11116);
nor U12412 (N_12412,N_11176,N_11824);
nand U12413 (N_12413,N_11496,N_11792);
or U12414 (N_12414,N_11505,N_11175);
nor U12415 (N_12415,N_11761,N_11279);
or U12416 (N_12416,N_11006,N_11385);
or U12417 (N_12417,N_11061,N_11849);
nand U12418 (N_12418,N_11461,N_11931);
or U12419 (N_12419,N_11709,N_11263);
or U12420 (N_12420,N_11336,N_11142);
nand U12421 (N_12421,N_11645,N_11277);
nand U12422 (N_12422,N_11289,N_11623);
nor U12423 (N_12423,N_11390,N_11268);
and U12424 (N_12424,N_11103,N_11690);
xor U12425 (N_12425,N_11531,N_11224);
nor U12426 (N_12426,N_11440,N_11774);
xor U12427 (N_12427,N_11730,N_11227);
and U12428 (N_12428,N_11499,N_11822);
nand U12429 (N_12429,N_11165,N_11689);
nor U12430 (N_12430,N_11913,N_11984);
or U12431 (N_12431,N_11853,N_11478);
xnor U12432 (N_12432,N_11415,N_11332);
or U12433 (N_12433,N_11550,N_11895);
and U12434 (N_12434,N_11598,N_11426);
xor U12435 (N_12435,N_11015,N_11782);
nand U12436 (N_12436,N_11775,N_11364);
nand U12437 (N_12437,N_11997,N_11670);
nor U12438 (N_12438,N_11316,N_11751);
xnor U12439 (N_12439,N_11532,N_11747);
and U12440 (N_12440,N_11552,N_11646);
nand U12441 (N_12441,N_11944,N_11328);
nor U12442 (N_12442,N_11547,N_11754);
xnor U12443 (N_12443,N_11079,N_11574);
xor U12444 (N_12444,N_11275,N_11331);
xnor U12445 (N_12445,N_11687,N_11229);
nand U12446 (N_12446,N_11904,N_11916);
and U12447 (N_12447,N_11310,N_11022);
nand U12448 (N_12448,N_11383,N_11187);
or U12449 (N_12449,N_11365,N_11639);
and U12450 (N_12450,N_11874,N_11565);
xnor U12451 (N_12451,N_11281,N_11195);
nor U12452 (N_12452,N_11045,N_11353);
nor U12453 (N_12453,N_11039,N_11634);
nand U12454 (N_12454,N_11456,N_11624);
xor U12455 (N_12455,N_11563,N_11834);
or U12456 (N_12456,N_11345,N_11998);
nand U12457 (N_12457,N_11093,N_11305);
nand U12458 (N_12458,N_11044,N_11032);
nor U12459 (N_12459,N_11608,N_11617);
xnor U12460 (N_12460,N_11452,N_11717);
or U12461 (N_12461,N_11489,N_11125);
xnor U12462 (N_12462,N_11734,N_11110);
xnor U12463 (N_12463,N_11386,N_11266);
nand U12464 (N_12464,N_11296,N_11968);
or U12465 (N_12465,N_11892,N_11876);
nand U12466 (N_12466,N_11325,N_11143);
or U12467 (N_12467,N_11250,N_11209);
nor U12468 (N_12468,N_11247,N_11744);
nand U12469 (N_12469,N_11007,N_11988);
nand U12470 (N_12470,N_11073,N_11588);
xor U12471 (N_12471,N_11351,N_11860);
nand U12472 (N_12472,N_11101,N_11090);
or U12473 (N_12473,N_11304,N_11218);
xnor U12474 (N_12474,N_11341,N_11389);
and U12475 (N_12475,N_11886,N_11955);
nor U12476 (N_12476,N_11680,N_11869);
and U12477 (N_12477,N_11075,N_11149);
or U12478 (N_12478,N_11753,N_11246);
nand U12479 (N_12479,N_11443,N_11463);
nor U12480 (N_12480,N_11371,N_11060);
nand U12481 (N_12481,N_11313,N_11769);
or U12482 (N_12482,N_11235,N_11587);
nand U12483 (N_12483,N_11788,N_11420);
nand U12484 (N_12484,N_11346,N_11154);
xor U12485 (N_12485,N_11790,N_11441);
and U12486 (N_12486,N_11394,N_11847);
and U12487 (N_12487,N_11188,N_11507);
or U12488 (N_12488,N_11259,N_11293);
or U12489 (N_12489,N_11306,N_11072);
or U12490 (N_12490,N_11556,N_11174);
nand U12491 (N_12491,N_11837,N_11189);
and U12492 (N_12492,N_11334,N_11650);
nor U12493 (N_12493,N_11795,N_11169);
or U12494 (N_12494,N_11595,N_11979);
and U12495 (N_12495,N_11238,N_11786);
nor U12496 (N_12496,N_11599,N_11216);
and U12497 (N_12497,N_11361,N_11160);
xor U12498 (N_12498,N_11483,N_11474);
nand U12499 (N_12499,N_11960,N_11549);
nand U12500 (N_12500,N_11631,N_11408);
and U12501 (N_12501,N_11183,N_11433);
or U12502 (N_12502,N_11089,N_11442);
and U12503 (N_12503,N_11401,N_11653);
or U12504 (N_12504,N_11690,N_11613);
and U12505 (N_12505,N_11250,N_11855);
xnor U12506 (N_12506,N_11678,N_11263);
nand U12507 (N_12507,N_11562,N_11833);
and U12508 (N_12508,N_11632,N_11187);
nor U12509 (N_12509,N_11439,N_11666);
xnor U12510 (N_12510,N_11535,N_11368);
nand U12511 (N_12511,N_11023,N_11668);
or U12512 (N_12512,N_11635,N_11327);
nand U12513 (N_12513,N_11875,N_11416);
and U12514 (N_12514,N_11014,N_11563);
xnor U12515 (N_12515,N_11034,N_11081);
xnor U12516 (N_12516,N_11862,N_11447);
nand U12517 (N_12517,N_11340,N_11591);
or U12518 (N_12518,N_11391,N_11441);
xor U12519 (N_12519,N_11629,N_11761);
nand U12520 (N_12520,N_11636,N_11299);
or U12521 (N_12521,N_11374,N_11862);
xnor U12522 (N_12522,N_11133,N_11848);
nand U12523 (N_12523,N_11247,N_11258);
or U12524 (N_12524,N_11539,N_11345);
or U12525 (N_12525,N_11017,N_11589);
and U12526 (N_12526,N_11343,N_11796);
and U12527 (N_12527,N_11944,N_11166);
xnor U12528 (N_12528,N_11014,N_11373);
nor U12529 (N_12529,N_11888,N_11838);
nand U12530 (N_12530,N_11104,N_11983);
nor U12531 (N_12531,N_11543,N_11453);
nor U12532 (N_12532,N_11330,N_11805);
and U12533 (N_12533,N_11051,N_11774);
and U12534 (N_12534,N_11750,N_11900);
nand U12535 (N_12535,N_11812,N_11673);
nand U12536 (N_12536,N_11568,N_11939);
or U12537 (N_12537,N_11696,N_11214);
or U12538 (N_12538,N_11521,N_11939);
and U12539 (N_12539,N_11671,N_11857);
nand U12540 (N_12540,N_11919,N_11946);
xor U12541 (N_12541,N_11488,N_11650);
nand U12542 (N_12542,N_11363,N_11829);
nand U12543 (N_12543,N_11954,N_11617);
xor U12544 (N_12544,N_11915,N_11325);
or U12545 (N_12545,N_11600,N_11764);
xnor U12546 (N_12546,N_11626,N_11438);
nand U12547 (N_12547,N_11041,N_11899);
nor U12548 (N_12548,N_11192,N_11013);
nand U12549 (N_12549,N_11210,N_11520);
or U12550 (N_12550,N_11553,N_11002);
or U12551 (N_12551,N_11395,N_11028);
or U12552 (N_12552,N_11243,N_11886);
xnor U12553 (N_12553,N_11247,N_11996);
nor U12554 (N_12554,N_11668,N_11821);
xnor U12555 (N_12555,N_11213,N_11871);
xnor U12556 (N_12556,N_11471,N_11714);
nand U12557 (N_12557,N_11058,N_11706);
and U12558 (N_12558,N_11024,N_11945);
nand U12559 (N_12559,N_11049,N_11503);
nor U12560 (N_12560,N_11174,N_11238);
or U12561 (N_12561,N_11643,N_11321);
xor U12562 (N_12562,N_11168,N_11526);
or U12563 (N_12563,N_11023,N_11753);
or U12564 (N_12564,N_11815,N_11921);
or U12565 (N_12565,N_11858,N_11746);
nor U12566 (N_12566,N_11568,N_11567);
xnor U12567 (N_12567,N_11059,N_11254);
xnor U12568 (N_12568,N_11425,N_11502);
xor U12569 (N_12569,N_11144,N_11434);
nor U12570 (N_12570,N_11823,N_11656);
nor U12571 (N_12571,N_11216,N_11684);
and U12572 (N_12572,N_11527,N_11470);
nor U12573 (N_12573,N_11582,N_11493);
and U12574 (N_12574,N_11955,N_11238);
xor U12575 (N_12575,N_11754,N_11282);
xnor U12576 (N_12576,N_11912,N_11739);
and U12577 (N_12577,N_11729,N_11059);
or U12578 (N_12578,N_11193,N_11223);
or U12579 (N_12579,N_11095,N_11113);
nand U12580 (N_12580,N_11064,N_11731);
nand U12581 (N_12581,N_11807,N_11377);
nand U12582 (N_12582,N_11917,N_11168);
or U12583 (N_12583,N_11347,N_11502);
nor U12584 (N_12584,N_11329,N_11139);
and U12585 (N_12585,N_11126,N_11097);
nand U12586 (N_12586,N_11642,N_11740);
and U12587 (N_12587,N_11714,N_11617);
or U12588 (N_12588,N_11991,N_11321);
or U12589 (N_12589,N_11489,N_11351);
or U12590 (N_12590,N_11001,N_11762);
xnor U12591 (N_12591,N_11820,N_11792);
and U12592 (N_12592,N_11620,N_11682);
or U12593 (N_12593,N_11801,N_11137);
nand U12594 (N_12594,N_11550,N_11977);
and U12595 (N_12595,N_11966,N_11449);
nand U12596 (N_12596,N_11777,N_11465);
nand U12597 (N_12597,N_11122,N_11481);
and U12598 (N_12598,N_11780,N_11855);
xor U12599 (N_12599,N_11161,N_11206);
nor U12600 (N_12600,N_11502,N_11316);
xor U12601 (N_12601,N_11593,N_11678);
xnor U12602 (N_12602,N_11038,N_11314);
nor U12603 (N_12603,N_11822,N_11630);
or U12604 (N_12604,N_11193,N_11205);
nand U12605 (N_12605,N_11654,N_11125);
nor U12606 (N_12606,N_11848,N_11840);
xnor U12607 (N_12607,N_11850,N_11563);
nor U12608 (N_12608,N_11454,N_11922);
or U12609 (N_12609,N_11564,N_11500);
and U12610 (N_12610,N_11300,N_11570);
or U12611 (N_12611,N_11194,N_11352);
nand U12612 (N_12612,N_11810,N_11499);
or U12613 (N_12613,N_11523,N_11350);
and U12614 (N_12614,N_11340,N_11795);
and U12615 (N_12615,N_11601,N_11066);
nand U12616 (N_12616,N_11510,N_11733);
xor U12617 (N_12617,N_11638,N_11356);
xnor U12618 (N_12618,N_11222,N_11891);
xor U12619 (N_12619,N_11286,N_11026);
and U12620 (N_12620,N_11390,N_11578);
nand U12621 (N_12621,N_11485,N_11667);
nor U12622 (N_12622,N_11096,N_11429);
or U12623 (N_12623,N_11319,N_11956);
nand U12624 (N_12624,N_11308,N_11479);
nand U12625 (N_12625,N_11250,N_11252);
or U12626 (N_12626,N_11041,N_11024);
nand U12627 (N_12627,N_11220,N_11781);
nor U12628 (N_12628,N_11967,N_11898);
nand U12629 (N_12629,N_11735,N_11594);
xnor U12630 (N_12630,N_11181,N_11095);
nand U12631 (N_12631,N_11271,N_11600);
xor U12632 (N_12632,N_11232,N_11807);
or U12633 (N_12633,N_11300,N_11356);
nor U12634 (N_12634,N_11952,N_11303);
and U12635 (N_12635,N_11123,N_11074);
nand U12636 (N_12636,N_11079,N_11798);
nor U12637 (N_12637,N_11495,N_11878);
and U12638 (N_12638,N_11491,N_11275);
xor U12639 (N_12639,N_11629,N_11656);
xor U12640 (N_12640,N_11127,N_11017);
and U12641 (N_12641,N_11344,N_11843);
or U12642 (N_12642,N_11821,N_11347);
xor U12643 (N_12643,N_11836,N_11804);
xnor U12644 (N_12644,N_11300,N_11887);
xnor U12645 (N_12645,N_11175,N_11544);
or U12646 (N_12646,N_11183,N_11693);
nand U12647 (N_12647,N_11054,N_11846);
xnor U12648 (N_12648,N_11845,N_11314);
nand U12649 (N_12649,N_11362,N_11641);
or U12650 (N_12650,N_11689,N_11445);
and U12651 (N_12651,N_11751,N_11308);
nor U12652 (N_12652,N_11699,N_11203);
or U12653 (N_12653,N_11302,N_11147);
or U12654 (N_12654,N_11813,N_11494);
nand U12655 (N_12655,N_11686,N_11579);
nor U12656 (N_12656,N_11257,N_11320);
nand U12657 (N_12657,N_11639,N_11519);
xnor U12658 (N_12658,N_11030,N_11524);
xnor U12659 (N_12659,N_11618,N_11493);
or U12660 (N_12660,N_11915,N_11698);
nand U12661 (N_12661,N_11321,N_11961);
and U12662 (N_12662,N_11138,N_11552);
and U12663 (N_12663,N_11999,N_11233);
nor U12664 (N_12664,N_11634,N_11340);
and U12665 (N_12665,N_11493,N_11485);
nand U12666 (N_12666,N_11424,N_11222);
nand U12667 (N_12667,N_11829,N_11998);
and U12668 (N_12668,N_11822,N_11784);
or U12669 (N_12669,N_11440,N_11978);
nand U12670 (N_12670,N_11888,N_11532);
nor U12671 (N_12671,N_11657,N_11045);
nor U12672 (N_12672,N_11816,N_11365);
and U12673 (N_12673,N_11480,N_11326);
or U12674 (N_12674,N_11349,N_11963);
or U12675 (N_12675,N_11880,N_11465);
or U12676 (N_12676,N_11741,N_11828);
nor U12677 (N_12677,N_11585,N_11115);
nand U12678 (N_12678,N_11126,N_11572);
or U12679 (N_12679,N_11099,N_11551);
xnor U12680 (N_12680,N_11503,N_11663);
and U12681 (N_12681,N_11588,N_11940);
nand U12682 (N_12682,N_11740,N_11138);
nor U12683 (N_12683,N_11620,N_11149);
and U12684 (N_12684,N_11043,N_11351);
nor U12685 (N_12685,N_11652,N_11347);
xor U12686 (N_12686,N_11562,N_11154);
nor U12687 (N_12687,N_11221,N_11154);
xnor U12688 (N_12688,N_11157,N_11550);
nand U12689 (N_12689,N_11051,N_11483);
and U12690 (N_12690,N_11433,N_11163);
and U12691 (N_12691,N_11082,N_11994);
nand U12692 (N_12692,N_11834,N_11779);
or U12693 (N_12693,N_11688,N_11794);
nor U12694 (N_12694,N_11725,N_11686);
nand U12695 (N_12695,N_11930,N_11264);
xor U12696 (N_12696,N_11639,N_11023);
xor U12697 (N_12697,N_11143,N_11660);
xnor U12698 (N_12698,N_11543,N_11212);
or U12699 (N_12699,N_11630,N_11670);
nand U12700 (N_12700,N_11847,N_11512);
nor U12701 (N_12701,N_11295,N_11373);
or U12702 (N_12702,N_11701,N_11877);
nor U12703 (N_12703,N_11714,N_11387);
or U12704 (N_12704,N_11010,N_11751);
and U12705 (N_12705,N_11198,N_11278);
xnor U12706 (N_12706,N_11260,N_11035);
nand U12707 (N_12707,N_11736,N_11887);
nor U12708 (N_12708,N_11080,N_11938);
xor U12709 (N_12709,N_11970,N_11844);
or U12710 (N_12710,N_11289,N_11740);
nand U12711 (N_12711,N_11036,N_11897);
xor U12712 (N_12712,N_11484,N_11847);
nand U12713 (N_12713,N_11443,N_11427);
nor U12714 (N_12714,N_11752,N_11309);
xor U12715 (N_12715,N_11559,N_11830);
nand U12716 (N_12716,N_11278,N_11201);
xnor U12717 (N_12717,N_11358,N_11196);
nor U12718 (N_12718,N_11558,N_11833);
and U12719 (N_12719,N_11963,N_11051);
nand U12720 (N_12720,N_11412,N_11846);
and U12721 (N_12721,N_11134,N_11425);
nand U12722 (N_12722,N_11412,N_11750);
and U12723 (N_12723,N_11076,N_11434);
nor U12724 (N_12724,N_11733,N_11746);
and U12725 (N_12725,N_11022,N_11923);
nand U12726 (N_12726,N_11925,N_11328);
nand U12727 (N_12727,N_11753,N_11570);
nor U12728 (N_12728,N_11477,N_11311);
xor U12729 (N_12729,N_11527,N_11962);
xor U12730 (N_12730,N_11118,N_11587);
or U12731 (N_12731,N_11073,N_11564);
nor U12732 (N_12732,N_11114,N_11208);
xor U12733 (N_12733,N_11557,N_11348);
nor U12734 (N_12734,N_11480,N_11203);
and U12735 (N_12735,N_11788,N_11663);
nor U12736 (N_12736,N_11606,N_11002);
xor U12737 (N_12737,N_11001,N_11696);
or U12738 (N_12738,N_11936,N_11581);
nor U12739 (N_12739,N_11470,N_11486);
or U12740 (N_12740,N_11564,N_11704);
nand U12741 (N_12741,N_11131,N_11860);
nor U12742 (N_12742,N_11083,N_11037);
xnor U12743 (N_12743,N_11641,N_11274);
nand U12744 (N_12744,N_11689,N_11529);
xnor U12745 (N_12745,N_11092,N_11195);
xnor U12746 (N_12746,N_11621,N_11985);
xor U12747 (N_12747,N_11723,N_11211);
and U12748 (N_12748,N_11321,N_11246);
nand U12749 (N_12749,N_11177,N_11359);
nor U12750 (N_12750,N_11576,N_11969);
nand U12751 (N_12751,N_11271,N_11583);
and U12752 (N_12752,N_11335,N_11325);
or U12753 (N_12753,N_11899,N_11268);
nor U12754 (N_12754,N_11286,N_11176);
xor U12755 (N_12755,N_11209,N_11320);
xor U12756 (N_12756,N_11250,N_11095);
or U12757 (N_12757,N_11444,N_11495);
xor U12758 (N_12758,N_11024,N_11667);
nand U12759 (N_12759,N_11504,N_11426);
nand U12760 (N_12760,N_11199,N_11443);
and U12761 (N_12761,N_11992,N_11920);
xor U12762 (N_12762,N_11416,N_11114);
nor U12763 (N_12763,N_11490,N_11695);
and U12764 (N_12764,N_11960,N_11425);
and U12765 (N_12765,N_11850,N_11321);
or U12766 (N_12766,N_11714,N_11937);
or U12767 (N_12767,N_11084,N_11863);
and U12768 (N_12768,N_11988,N_11129);
xor U12769 (N_12769,N_11747,N_11305);
and U12770 (N_12770,N_11334,N_11321);
xor U12771 (N_12771,N_11322,N_11318);
and U12772 (N_12772,N_11785,N_11551);
xnor U12773 (N_12773,N_11482,N_11010);
and U12774 (N_12774,N_11625,N_11855);
nor U12775 (N_12775,N_11052,N_11367);
or U12776 (N_12776,N_11343,N_11785);
xor U12777 (N_12777,N_11098,N_11158);
and U12778 (N_12778,N_11214,N_11343);
nand U12779 (N_12779,N_11319,N_11900);
nor U12780 (N_12780,N_11764,N_11963);
xnor U12781 (N_12781,N_11709,N_11526);
nand U12782 (N_12782,N_11394,N_11622);
or U12783 (N_12783,N_11470,N_11860);
nand U12784 (N_12784,N_11760,N_11122);
or U12785 (N_12785,N_11048,N_11803);
nor U12786 (N_12786,N_11491,N_11371);
nand U12787 (N_12787,N_11021,N_11473);
or U12788 (N_12788,N_11823,N_11586);
xnor U12789 (N_12789,N_11155,N_11046);
nand U12790 (N_12790,N_11007,N_11257);
nor U12791 (N_12791,N_11637,N_11257);
and U12792 (N_12792,N_11099,N_11448);
or U12793 (N_12793,N_11411,N_11190);
and U12794 (N_12794,N_11375,N_11336);
and U12795 (N_12795,N_11268,N_11296);
xor U12796 (N_12796,N_11053,N_11224);
nand U12797 (N_12797,N_11087,N_11083);
or U12798 (N_12798,N_11941,N_11846);
or U12799 (N_12799,N_11463,N_11459);
or U12800 (N_12800,N_11428,N_11269);
and U12801 (N_12801,N_11212,N_11254);
nor U12802 (N_12802,N_11808,N_11552);
and U12803 (N_12803,N_11024,N_11784);
xnor U12804 (N_12804,N_11008,N_11845);
nand U12805 (N_12805,N_11615,N_11020);
nor U12806 (N_12806,N_11125,N_11114);
xor U12807 (N_12807,N_11064,N_11886);
nand U12808 (N_12808,N_11611,N_11002);
xor U12809 (N_12809,N_11694,N_11470);
and U12810 (N_12810,N_11131,N_11198);
xor U12811 (N_12811,N_11020,N_11702);
nor U12812 (N_12812,N_11290,N_11251);
nor U12813 (N_12813,N_11434,N_11273);
or U12814 (N_12814,N_11483,N_11517);
nand U12815 (N_12815,N_11762,N_11177);
and U12816 (N_12816,N_11087,N_11600);
nor U12817 (N_12817,N_11682,N_11961);
nand U12818 (N_12818,N_11318,N_11232);
nor U12819 (N_12819,N_11637,N_11571);
nand U12820 (N_12820,N_11558,N_11589);
nor U12821 (N_12821,N_11045,N_11855);
or U12822 (N_12822,N_11092,N_11023);
nand U12823 (N_12823,N_11658,N_11502);
and U12824 (N_12824,N_11925,N_11631);
nor U12825 (N_12825,N_11139,N_11933);
nand U12826 (N_12826,N_11707,N_11054);
or U12827 (N_12827,N_11343,N_11435);
nor U12828 (N_12828,N_11896,N_11965);
nand U12829 (N_12829,N_11630,N_11488);
nor U12830 (N_12830,N_11586,N_11345);
nor U12831 (N_12831,N_11559,N_11287);
xnor U12832 (N_12832,N_11536,N_11975);
nand U12833 (N_12833,N_11653,N_11714);
xnor U12834 (N_12834,N_11419,N_11335);
nand U12835 (N_12835,N_11583,N_11865);
nor U12836 (N_12836,N_11199,N_11521);
xnor U12837 (N_12837,N_11371,N_11269);
or U12838 (N_12838,N_11690,N_11014);
and U12839 (N_12839,N_11889,N_11323);
nor U12840 (N_12840,N_11745,N_11128);
and U12841 (N_12841,N_11895,N_11489);
nor U12842 (N_12842,N_11263,N_11233);
nand U12843 (N_12843,N_11035,N_11579);
or U12844 (N_12844,N_11742,N_11575);
and U12845 (N_12845,N_11292,N_11913);
or U12846 (N_12846,N_11451,N_11795);
xor U12847 (N_12847,N_11503,N_11433);
and U12848 (N_12848,N_11345,N_11762);
xor U12849 (N_12849,N_11573,N_11118);
nand U12850 (N_12850,N_11343,N_11622);
and U12851 (N_12851,N_11758,N_11220);
or U12852 (N_12852,N_11275,N_11049);
nand U12853 (N_12853,N_11865,N_11676);
nor U12854 (N_12854,N_11968,N_11509);
nand U12855 (N_12855,N_11026,N_11924);
or U12856 (N_12856,N_11774,N_11900);
or U12857 (N_12857,N_11358,N_11230);
nand U12858 (N_12858,N_11453,N_11462);
nand U12859 (N_12859,N_11389,N_11928);
and U12860 (N_12860,N_11538,N_11806);
nor U12861 (N_12861,N_11718,N_11575);
or U12862 (N_12862,N_11232,N_11075);
nand U12863 (N_12863,N_11041,N_11390);
and U12864 (N_12864,N_11433,N_11216);
nor U12865 (N_12865,N_11295,N_11289);
and U12866 (N_12866,N_11023,N_11843);
nor U12867 (N_12867,N_11556,N_11092);
xnor U12868 (N_12868,N_11126,N_11257);
nand U12869 (N_12869,N_11232,N_11205);
or U12870 (N_12870,N_11252,N_11202);
or U12871 (N_12871,N_11222,N_11184);
nor U12872 (N_12872,N_11392,N_11009);
nand U12873 (N_12873,N_11629,N_11698);
nor U12874 (N_12874,N_11531,N_11565);
xnor U12875 (N_12875,N_11379,N_11349);
or U12876 (N_12876,N_11094,N_11541);
and U12877 (N_12877,N_11413,N_11996);
and U12878 (N_12878,N_11814,N_11310);
xor U12879 (N_12879,N_11778,N_11389);
or U12880 (N_12880,N_11506,N_11642);
and U12881 (N_12881,N_11760,N_11486);
and U12882 (N_12882,N_11273,N_11582);
nand U12883 (N_12883,N_11084,N_11914);
and U12884 (N_12884,N_11849,N_11707);
xnor U12885 (N_12885,N_11423,N_11146);
nand U12886 (N_12886,N_11044,N_11877);
nand U12887 (N_12887,N_11892,N_11891);
or U12888 (N_12888,N_11499,N_11902);
nand U12889 (N_12889,N_11820,N_11723);
nand U12890 (N_12890,N_11533,N_11253);
and U12891 (N_12891,N_11893,N_11164);
xor U12892 (N_12892,N_11811,N_11309);
and U12893 (N_12893,N_11491,N_11283);
xnor U12894 (N_12894,N_11940,N_11110);
nor U12895 (N_12895,N_11099,N_11347);
and U12896 (N_12896,N_11496,N_11394);
and U12897 (N_12897,N_11266,N_11122);
xnor U12898 (N_12898,N_11987,N_11218);
and U12899 (N_12899,N_11527,N_11960);
and U12900 (N_12900,N_11195,N_11536);
nor U12901 (N_12901,N_11521,N_11810);
xnor U12902 (N_12902,N_11972,N_11145);
and U12903 (N_12903,N_11452,N_11767);
or U12904 (N_12904,N_11434,N_11565);
xnor U12905 (N_12905,N_11598,N_11985);
nor U12906 (N_12906,N_11998,N_11426);
nor U12907 (N_12907,N_11509,N_11158);
and U12908 (N_12908,N_11374,N_11112);
xor U12909 (N_12909,N_11425,N_11018);
and U12910 (N_12910,N_11043,N_11434);
xnor U12911 (N_12911,N_11427,N_11675);
nand U12912 (N_12912,N_11494,N_11613);
or U12913 (N_12913,N_11695,N_11227);
xor U12914 (N_12914,N_11156,N_11030);
or U12915 (N_12915,N_11860,N_11058);
and U12916 (N_12916,N_11212,N_11817);
xor U12917 (N_12917,N_11891,N_11906);
nand U12918 (N_12918,N_11127,N_11436);
xor U12919 (N_12919,N_11781,N_11920);
xnor U12920 (N_12920,N_11002,N_11788);
xnor U12921 (N_12921,N_11581,N_11962);
xnor U12922 (N_12922,N_11367,N_11436);
or U12923 (N_12923,N_11637,N_11945);
and U12924 (N_12924,N_11378,N_11185);
nand U12925 (N_12925,N_11456,N_11269);
nor U12926 (N_12926,N_11881,N_11462);
nor U12927 (N_12927,N_11547,N_11427);
and U12928 (N_12928,N_11994,N_11216);
xor U12929 (N_12929,N_11617,N_11425);
nand U12930 (N_12930,N_11967,N_11905);
nand U12931 (N_12931,N_11043,N_11752);
and U12932 (N_12932,N_11976,N_11544);
or U12933 (N_12933,N_11077,N_11836);
and U12934 (N_12934,N_11743,N_11095);
or U12935 (N_12935,N_11891,N_11483);
and U12936 (N_12936,N_11851,N_11890);
nand U12937 (N_12937,N_11135,N_11859);
nand U12938 (N_12938,N_11908,N_11002);
xnor U12939 (N_12939,N_11834,N_11154);
or U12940 (N_12940,N_11766,N_11283);
xor U12941 (N_12941,N_11153,N_11499);
and U12942 (N_12942,N_11035,N_11381);
or U12943 (N_12943,N_11137,N_11824);
and U12944 (N_12944,N_11058,N_11259);
nor U12945 (N_12945,N_11724,N_11457);
and U12946 (N_12946,N_11374,N_11896);
nand U12947 (N_12947,N_11437,N_11033);
and U12948 (N_12948,N_11617,N_11849);
nand U12949 (N_12949,N_11459,N_11333);
and U12950 (N_12950,N_11180,N_11701);
and U12951 (N_12951,N_11088,N_11586);
nand U12952 (N_12952,N_11193,N_11371);
nor U12953 (N_12953,N_11508,N_11652);
nand U12954 (N_12954,N_11640,N_11250);
nor U12955 (N_12955,N_11282,N_11711);
or U12956 (N_12956,N_11839,N_11723);
nor U12957 (N_12957,N_11338,N_11823);
nand U12958 (N_12958,N_11240,N_11039);
xor U12959 (N_12959,N_11381,N_11437);
or U12960 (N_12960,N_11637,N_11011);
nand U12961 (N_12961,N_11444,N_11125);
nand U12962 (N_12962,N_11919,N_11043);
nor U12963 (N_12963,N_11263,N_11335);
nor U12964 (N_12964,N_11803,N_11354);
xor U12965 (N_12965,N_11161,N_11045);
and U12966 (N_12966,N_11210,N_11661);
nand U12967 (N_12967,N_11250,N_11211);
xor U12968 (N_12968,N_11650,N_11915);
or U12969 (N_12969,N_11590,N_11899);
nor U12970 (N_12970,N_11654,N_11222);
xnor U12971 (N_12971,N_11104,N_11850);
nor U12972 (N_12972,N_11248,N_11408);
and U12973 (N_12973,N_11908,N_11305);
and U12974 (N_12974,N_11376,N_11379);
xor U12975 (N_12975,N_11747,N_11547);
or U12976 (N_12976,N_11049,N_11090);
nand U12977 (N_12977,N_11463,N_11569);
or U12978 (N_12978,N_11909,N_11572);
nand U12979 (N_12979,N_11825,N_11291);
xnor U12980 (N_12980,N_11342,N_11545);
xnor U12981 (N_12981,N_11960,N_11765);
or U12982 (N_12982,N_11711,N_11232);
nor U12983 (N_12983,N_11339,N_11198);
or U12984 (N_12984,N_11220,N_11382);
and U12985 (N_12985,N_11982,N_11396);
nor U12986 (N_12986,N_11108,N_11665);
or U12987 (N_12987,N_11336,N_11252);
xnor U12988 (N_12988,N_11463,N_11022);
nor U12989 (N_12989,N_11223,N_11408);
nand U12990 (N_12990,N_11567,N_11254);
or U12991 (N_12991,N_11041,N_11052);
nor U12992 (N_12992,N_11236,N_11457);
or U12993 (N_12993,N_11385,N_11304);
xnor U12994 (N_12994,N_11707,N_11991);
or U12995 (N_12995,N_11866,N_11047);
xnor U12996 (N_12996,N_11138,N_11034);
and U12997 (N_12997,N_11925,N_11906);
nand U12998 (N_12998,N_11804,N_11848);
xnor U12999 (N_12999,N_11399,N_11029);
or U13000 (N_13000,N_12231,N_12983);
or U13001 (N_13001,N_12192,N_12777);
xnor U13002 (N_13002,N_12428,N_12481);
xor U13003 (N_13003,N_12506,N_12013);
and U13004 (N_13004,N_12573,N_12441);
or U13005 (N_13005,N_12408,N_12136);
nand U13006 (N_13006,N_12423,N_12034);
nand U13007 (N_13007,N_12512,N_12942);
nand U13008 (N_13008,N_12724,N_12095);
and U13009 (N_13009,N_12044,N_12529);
and U13010 (N_13010,N_12885,N_12356);
and U13011 (N_13011,N_12761,N_12659);
nor U13012 (N_13012,N_12985,N_12023);
xor U13013 (N_13013,N_12680,N_12910);
nand U13014 (N_13014,N_12490,N_12899);
xnor U13015 (N_13015,N_12503,N_12120);
nor U13016 (N_13016,N_12598,N_12909);
or U13017 (N_13017,N_12113,N_12030);
or U13018 (N_13018,N_12784,N_12210);
or U13019 (N_13019,N_12997,N_12400);
nand U13020 (N_13020,N_12066,N_12736);
nand U13021 (N_13021,N_12774,N_12867);
xor U13022 (N_13022,N_12650,N_12460);
nor U13023 (N_13023,N_12072,N_12035);
xor U13024 (N_13024,N_12263,N_12339);
or U13025 (N_13025,N_12752,N_12473);
xnor U13026 (N_13026,N_12472,N_12211);
nor U13027 (N_13027,N_12522,N_12103);
nand U13028 (N_13028,N_12563,N_12841);
nand U13029 (N_13029,N_12002,N_12275);
xnor U13030 (N_13030,N_12001,N_12438);
xnor U13031 (N_13031,N_12298,N_12897);
nor U13032 (N_13032,N_12766,N_12468);
nand U13033 (N_13033,N_12905,N_12756);
and U13034 (N_13034,N_12809,N_12178);
nor U13035 (N_13035,N_12803,N_12638);
or U13036 (N_13036,N_12243,N_12031);
nor U13037 (N_13037,N_12975,N_12943);
xor U13038 (N_13038,N_12854,N_12163);
and U13039 (N_13039,N_12209,N_12966);
nand U13040 (N_13040,N_12050,N_12973);
or U13041 (N_13041,N_12218,N_12951);
nand U13042 (N_13042,N_12729,N_12139);
nor U13043 (N_13043,N_12620,N_12632);
and U13044 (N_13044,N_12306,N_12362);
nor U13045 (N_13045,N_12168,N_12076);
nor U13046 (N_13046,N_12492,N_12179);
and U13047 (N_13047,N_12737,N_12292);
nand U13048 (N_13048,N_12797,N_12117);
xnor U13049 (N_13049,N_12253,N_12456);
xor U13050 (N_13050,N_12182,N_12334);
and U13051 (N_13051,N_12222,N_12068);
nor U13052 (N_13052,N_12452,N_12319);
or U13053 (N_13053,N_12501,N_12080);
xor U13054 (N_13054,N_12554,N_12486);
or U13055 (N_13055,N_12061,N_12735);
nor U13056 (N_13056,N_12954,N_12961);
or U13057 (N_13057,N_12892,N_12206);
nand U13058 (N_13058,N_12596,N_12556);
nand U13059 (N_13059,N_12886,N_12183);
xor U13060 (N_13060,N_12697,N_12682);
or U13061 (N_13061,N_12717,N_12419);
nand U13062 (N_13062,N_12753,N_12592);
nand U13063 (N_13063,N_12439,N_12232);
and U13064 (N_13064,N_12545,N_12330);
nor U13065 (N_13065,N_12345,N_12581);
nor U13066 (N_13066,N_12491,N_12177);
nand U13067 (N_13067,N_12842,N_12517);
xnor U13068 (N_13068,N_12546,N_12691);
or U13069 (N_13069,N_12935,N_12602);
and U13070 (N_13070,N_12436,N_12042);
and U13071 (N_13071,N_12432,N_12130);
xnor U13072 (N_13072,N_12974,N_12270);
or U13073 (N_13073,N_12744,N_12692);
xnor U13074 (N_13074,N_12149,N_12838);
xor U13075 (N_13075,N_12722,N_12685);
xor U13076 (N_13076,N_12134,N_12584);
xor U13077 (N_13077,N_12824,N_12391);
xnor U13078 (N_13078,N_12091,N_12302);
and U13079 (N_13079,N_12967,N_12863);
and U13080 (N_13080,N_12213,N_12336);
and U13081 (N_13081,N_12241,N_12521);
nor U13082 (N_13082,N_12881,N_12461);
or U13083 (N_13083,N_12763,N_12748);
xor U13084 (N_13084,N_12977,N_12953);
or U13085 (N_13085,N_12105,N_12559);
nor U13086 (N_13086,N_12081,N_12937);
nand U13087 (N_13087,N_12660,N_12200);
nand U13088 (N_13088,N_12971,N_12949);
nor U13089 (N_13089,N_12415,N_12127);
xor U13090 (N_13090,N_12317,N_12033);
nor U13091 (N_13091,N_12564,N_12955);
nand U13092 (N_13092,N_12769,N_12877);
or U13093 (N_13093,N_12626,N_12739);
or U13094 (N_13094,N_12706,N_12801);
nor U13095 (N_13095,N_12026,N_12301);
nand U13096 (N_13096,N_12143,N_12403);
and U13097 (N_13097,N_12643,N_12010);
nand U13098 (N_13098,N_12174,N_12131);
xor U13099 (N_13099,N_12625,N_12508);
and U13100 (N_13100,N_12695,N_12151);
xor U13101 (N_13101,N_12252,N_12984);
nand U13102 (N_13102,N_12202,N_12500);
xor U13103 (N_13103,N_12229,N_12039);
nor U13104 (N_13104,N_12537,N_12772);
and U13105 (N_13105,N_12819,N_12580);
nor U13106 (N_13106,N_12681,N_12274);
and U13107 (N_13107,N_12184,N_12327);
xor U13108 (N_13108,N_12687,N_12276);
nand U13109 (N_13109,N_12762,N_12226);
nand U13110 (N_13110,N_12725,N_12431);
and U13111 (N_13111,N_12324,N_12058);
nand U13112 (N_13112,N_12250,N_12849);
nor U13113 (N_13113,N_12048,N_12121);
and U13114 (N_13114,N_12579,N_12893);
nor U13115 (N_13115,N_12147,N_12440);
or U13116 (N_13116,N_12913,N_12020);
and U13117 (N_13117,N_12212,N_12623);
and U13118 (N_13118,N_12287,N_12426);
and U13119 (N_13119,N_12845,N_12323);
and U13120 (N_13120,N_12145,N_12670);
or U13121 (N_13121,N_12561,N_12982);
nand U13122 (N_13122,N_12173,N_12606);
nor U13123 (N_13123,N_12360,N_12219);
nand U13124 (N_13124,N_12126,N_12227);
xnor U13125 (N_13125,N_12783,N_12217);
nor U13126 (N_13126,N_12349,N_12815);
nand U13127 (N_13127,N_12645,N_12203);
and U13128 (N_13128,N_12237,N_12847);
nand U13129 (N_13129,N_12382,N_12810);
nand U13130 (N_13130,N_12853,N_12363);
nand U13131 (N_13131,N_12560,N_12884);
or U13132 (N_13132,N_12822,N_12085);
and U13133 (N_13133,N_12940,N_12991);
nor U13134 (N_13134,N_12731,N_12914);
xor U13135 (N_13135,N_12751,N_12607);
or U13136 (N_13136,N_12280,N_12032);
xnor U13137 (N_13137,N_12021,N_12873);
or U13138 (N_13138,N_12365,N_12814);
and U13139 (N_13139,N_12547,N_12467);
and U13140 (N_13140,N_12871,N_12194);
and U13141 (N_13141,N_12236,N_12583);
or U13142 (N_13142,N_12102,N_12862);
or U13143 (N_13143,N_12962,N_12075);
or U13144 (N_13144,N_12417,N_12109);
nor U13145 (N_13145,N_12511,N_12829);
nand U13146 (N_13146,N_12480,N_12358);
nand U13147 (N_13147,N_12668,N_12894);
nor U13148 (N_13148,N_12679,N_12310);
and U13149 (N_13149,N_12525,N_12843);
nor U13150 (N_13150,N_12666,N_12006);
xnor U13151 (N_13151,N_12123,N_12390);
xor U13152 (N_13152,N_12097,N_12007);
nor U13153 (N_13153,N_12989,N_12826);
xor U13154 (N_13154,N_12510,N_12443);
xnor U13155 (N_13155,N_12667,N_12247);
xnor U13156 (N_13156,N_12255,N_12883);
nand U13157 (N_13157,N_12749,N_12344);
nand U13158 (N_13158,N_12536,N_12996);
or U13159 (N_13159,N_12703,N_12792);
and U13160 (N_13160,N_12656,N_12214);
nand U13161 (N_13161,N_12577,N_12342);
nor U13162 (N_13162,N_12693,N_12240);
xnor U13163 (N_13163,N_12812,N_12465);
xor U13164 (N_13164,N_12807,N_12868);
or U13165 (N_13165,N_12768,N_12383);
and U13166 (N_13166,N_12187,N_12233);
nor U13167 (N_13167,N_12278,N_12542);
and U13168 (N_13168,N_12716,N_12662);
or U13169 (N_13169,N_12856,N_12267);
or U13170 (N_13170,N_12958,N_12552);
nor U13171 (N_13171,N_12300,N_12321);
and U13172 (N_13172,N_12290,N_12830);
or U13173 (N_13173,N_12470,N_12303);
nand U13174 (N_13174,N_12029,N_12540);
and U13175 (N_13175,N_12462,N_12515);
xor U13176 (N_13176,N_12994,N_12129);
xor U13177 (N_13177,N_12159,N_12538);
xnor U13178 (N_13178,N_12291,N_12543);
and U13179 (N_13179,N_12057,N_12568);
nand U13180 (N_13180,N_12037,N_12857);
xnor U13181 (N_13181,N_12496,N_12702);
and U13182 (N_13182,N_12530,N_12992);
nand U13183 (N_13183,N_12939,N_12256);
and U13184 (N_13184,N_12874,N_12934);
and U13185 (N_13185,N_12089,N_12099);
xor U13186 (N_13186,N_12347,N_12686);
and U13187 (N_13187,N_12981,N_12605);
and U13188 (N_13188,N_12879,N_12947);
nor U13189 (N_13189,N_12759,N_12180);
xor U13190 (N_13190,N_12112,N_12926);
or U13191 (N_13191,N_12396,N_12464);
xor U13192 (N_13192,N_12457,N_12789);
nand U13193 (N_13193,N_12335,N_12088);
nor U13194 (N_13194,N_12155,N_12566);
xnor U13195 (N_13195,N_12442,N_12313);
nor U13196 (N_13196,N_12017,N_12395);
nor U13197 (N_13197,N_12906,N_12189);
or U13198 (N_13198,N_12377,N_12137);
xor U13199 (N_13199,N_12713,N_12993);
nor U13200 (N_13200,N_12435,N_12533);
or U13201 (N_13201,N_12084,N_12312);
or U13202 (N_13202,N_12535,N_12701);
and U13203 (N_13203,N_12271,N_12927);
or U13204 (N_13204,N_12534,N_12786);
and U13205 (N_13205,N_12086,N_12888);
and U13206 (N_13206,N_12328,N_12728);
or U13207 (N_13207,N_12562,N_12098);
nor U13208 (N_13208,N_12146,N_12705);
nand U13209 (N_13209,N_12311,N_12631);
or U13210 (N_13210,N_12889,N_12073);
nor U13211 (N_13211,N_12925,N_12646);
or U13212 (N_13212,N_12876,N_12730);
nor U13213 (N_13213,N_12627,N_12633);
xnor U13214 (N_13214,N_12230,N_12844);
and U13215 (N_13215,N_12498,N_12808);
nor U13216 (N_13216,N_12069,N_12289);
xnor U13217 (N_13217,N_12272,N_12524);
or U13218 (N_13218,N_12639,N_12388);
xor U13219 (N_13219,N_12776,N_12316);
nand U13220 (N_13220,N_12594,N_12615);
nand U13221 (N_13221,N_12455,N_12389);
nor U13222 (N_13222,N_12671,N_12049);
nor U13223 (N_13223,N_12657,N_12418);
and U13224 (N_13224,N_12348,N_12448);
nor U13225 (N_13225,N_12025,N_12340);
xor U13226 (N_13226,N_12652,N_12721);
xor U13227 (N_13227,N_12157,N_12239);
or U13228 (N_13228,N_12489,N_12019);
xnor U13229 (N_13229,N_12795,N_12640);
or U13230 (N_13230,N_12320,N_12374);
or U13231 (N_13231,N_12518,N_12434);
nor U13232 (N_13232,N_12188,N_12065);
nor U13233 (N_13233,N_12082,N_12308);
nor U13234 (N_13234,N_12016,N_12135);
nor U13235 (N_13235,N_12454,N_12848);
or U13236 (N_13236,N_12478,N_12800);
xor U13237 (N_13237,N_12411,N_12921);
nor U13238 (N_13238,N_12223,N_12637);
and U13239 (N_13239,N_12254,N_12970);
nand U13240 (N_13240,N_12846,N_12850);
and U13241 (N_13241,N_12946,N_12917);
and U13242 (N_13242,N_12198,N_12595);
xnor U13243 (N_13243,N_12437,N_12351);
or U13244 (N_13244,N_12047,N_12414);
and U13245 (N_13245,N_12285,N_12726);
nor U13246 (N_13246,N_12858,N_12495);
or U13247 (N_13247,N_12908,N_12235);
or U13248 (N_13248,N_12128,N_12555);
and U13249 (N_13249,N_12618,N_12141);
and U13250 (N_13250,N_12197,N_12684);
or U13251 (N_13251,N_12746,N_12059);
nor U13252 (N_13252,N_12251,N_12354);
and U13253 (N_13253,N_12386,N_12181);
or U13254 (N_13254,N_12372,N_12244);
nor U13255 (N_13255,N_12635,N_12449);
xnor U13256 (N_13256,N_12930,N_12170);
and U13257 (N_13257,N_12046,N_12790);
or U13258 (N_13258,N_12060,N_12787);
nand U13259 (N_13259,N_12932,N_12164);
or U13260 (N_13260,N_12648,N_12928);
xor U13261 (N_13261,N_12882,N_12591);
nand U13262 (N_13262,N_12798,N_12264);
or U13263 (N_13263,N_12972,N_12907);
xor U13264 (N_13264,N_12794,N_12176);
xnor U13265 (N_13265,N_12333,N_12754);
nand U13266 (N_13266,N_12661,N_12331);
and U13267 (N_13267,N_12322,N_12315);
and U13268 (N_13268,N_12720,N_12575);
and U13269 (N_13269,N_12096,N_12523);
xor U13270 (N_13270,N_12453,N_12869);
nor U13271 (N_13271,N_12444,N_12870);
nor U13272 (N_13272,N_12549,N_12696);
and U13273 (N_13273,N_12484,N_12507);
nand U13274 (N_13274,N_12835,N_12420);
nor U13275 (N_13275,N_12804,N_12038);
nand U13276 (N_13276,N_12343,N_12262);
xnor U13277 (N_13277,N_12269,N_12911);
nand U13278 (N_13278,N_12788,N_12249);
and U13279 (N_13279,N_12427,N_12544);
and U13280 (N_13280,N_12663,N_12410);
xnor U13281 (N_13281,N_12369,N_12572);
and U13282 (N_13282,N_12916,N_12630);
xor U13283 (N_13283,N_12248,N_12502);
nor U13284 (N_13284,N_12053,N_12169);
xnor U13285 (N_13285,N_12709,N_12688);
nor U13286 (N_13286,N_12895,N_12375);
xnor U13287 (N_13287,N_12265,N_12837);
and U13288 (N_13288,N_12036,N_12266);
xnor U13289 (N_13289,N_12475,N_12150);
xnor U13290 (N_13290,N_12000,N_12959);
xnor U13291 (N_13291,N_12132,N_12405);
or U13292 (N_13292,N_12152,N_12509);
and U13293 (N_13293,N_12407,N_12541);
nand U13294 (N_13294,N_12381,N_12373);
and U13295 (N_13295,N_12821,N_12074);
xnor U13296 (N_13296,N_12471,N_12352);
xor U13297 (N_13297,N_12379,N_12477);
nor U13298 (N_13298,N_12872,N_12664);
or U13299 (N_13299,N_12919,N_12171);
nor U13300 (N_13300,N_12293,N_12782);
or U13301 (N_13301,N_12234,N_12451);
nand U13302 (N_13302,N_12531,N_12952);
nor U13303 (N_13303,N_12571,N_12487);
nand U13304 (N_13304,N_12430,N_12398);
xor U13305 (N_13305,N_12516,N_12100);
nand U13306 (N_13306,N_12865,N_12111);
and U13307 (N_13307,N_12378,N_12497);
and U13308 (N_13308,N_12887,N_12931);
xor U13309 (N_13309,N_12208,N_12422);
xnor U13310 (N_13310,N_12649,N_12305);
nand U13311 (N_13311,N_12108,N_12778);
nor U13312 (N_13312,N_12576,N_12578);
xnor U13313 (N_13313,N_12175,N_12401);
and U13314 (N_13314,N_12063,N_12834);
or U13315 (N_13315,N_12077,N_12669);
xor U13316 (N_13316,N_12228,N_12677);
or U13317 (N_13317,N_12307,N_12604);
or U13318 (N_13318,N_12104,N_12380);
nand U13319 (N_13319,N_12964,N_12647);
nand U13320 (N_13320,N_12160,N_12505);
nand U13321 (N_13321,N_12738,N_12676);
and U13322 (N_13322,N_12008,N_12817);
and U13323 (N_13323,N_12610,N_12366);
and U13324 (N_13324,N_12732,N_12785);
nor U13325 (N_13325,N_12570,N_12755);
xnor U13326 (N_13326,N_12186,N_12476);
and U13327 (N_13327,N_12963,N_12424);
or U13328 (N_13328,N_12153,N_12624);
or U13329 (N_13329,N_12294,N_12459);
nand U13330 (N_13330,N_12162,N_12041);
xnor U13331 (N_13331,N_12723,N_12585);
xor U13332 (N_13332,N_12929,N_12941);
or U13333 (N_13333,N_12124,N_12586);
or U13334 (N_13334,N_12043,N_12799);
nor U13335 (N_13335,N_12960,N_12698);
and U13336 (N_13336,N_12742,N_12326);
or U13337 (N_13337,N_12384,N_12158);
xor U13338 (N_13338,N_12483,N_12079);
nand U13339 (N_13339,N_12318,N_12770);
and U13340 (N_13340,N_12968,N_12519);
and U13341 (N_13341,N_12548,N_12840);
or U13342 (N_13342,N_12864,N_12654);
nand U13343 (N_13343,N_12779,N_12195);
nor U13344 (N_13344,N_12745,N_12704);
nand U13345 (N_13345,N_12413,N_12499);
nand U13346 (N_13346,N_12904,N_12791);
xnor U13347 (N_13347,N_12012,N_12558);
or U13348 (N_13348,N_12998,N_12027);
nor U13349 (N_13349,N_12614,N_12070);
xor U13350 (N_13350,N_12936,N_12167);
nand U13351 (N_13351,N_12004,N_12283);
nand U13352 (N_13352,N_12781,N_12933);
nor U13353 (N_13353,N_12603,N_12458);
and U13354 (N_13354,N_12593,N_12711);
nor U13355 (N_13355,N_12148,N_12273);
or U13356 (N_13356,N_12675,N_12793);
and U13357 (N_13357,N_12969,N_12092);
nand U13358 (N_13358,N_12304,N_12634);
nand U13359 (N_13359,N_12504,N_12775);
nand U13360 (N_13360,N_12689,N_12071);
nand U13361 (N_13361,N_12172,N_12694);
xnor U13362 (N_13362,N_12474,N_12527);
or U13363 (N_13363,N_12553,N_12446);
nor U13364 (N_13364,N_12945,N_12140);
nor U13365 (N_13365,N_12064,N_12938);
xor U13366 (N_13366,N_12513,N_12062);
nor U13367 (N_13367,N_12851,N_12839);
nand U13368 (N_13368,N_12976,N_12642);
nor U13369 (N_13369,N_12205,N_12221);
or U13370 (N_13370,N_12878,N_12715);
xnor U13371 (N_13371,N_12918,N_12101);
or U13372 (N_13372,N_12118,N_12813);
nor U13373 (N_13373,N_12806,N_12619);
nand U13374 (N_13374,N_12258,N_12052);
xnor U13375 (N_13375,N_12040,N_12286);
nor U13376 (N_13376,N_12616,N_12599);
and U13377 (N_13377,N_12820,N_12245);
nor U13378 (N_13378,N_12611,N_12674);
and U13379 (N_13379,N_12574,N_12028);
and U13380 (N_13380,N_12811,N_12980);
xnor U13381 (N_13381,N_12597,N_12718);
xnor U13382 (N_13382,N_12528,N_12116);
or U13383 (N_13383,N_12196,N_12370);
nor U13384 (N_13384,N_12295,N_12346);
or U13385 (N_13385,N_12710,N_12796);
xnor U13386 (N_13386,N_12609,N_12397);
and U13387 (N_13387,N_12714,N_12394);
nor U13388 (N_13388,N_12412,N_12056);
xnor U13389 (N_13389,N_12087,N_12242);
or U13390 (N_13390,N_12199,N_12995);
nor U13391 (N_13391,N_12780,N_12204);
or U13392 (N_13392,N_12297,N_12246);
or U13393 (N_13393,N_12156,N_12133);
xor U13394 (N_13394,N_12433,N_12896);
and U13395 (N_13395,N_12760,N_12055);
or U13396 (N_13396,N_12683,N_12387);
and U13397 (N_13397,N_12622,N_12402);
nor U13398 (N_13398,N_12831,N_12651);
nor U13399 (N_13399,N_12083,N_12416);
nand U13400 (N_13400,N_12257,N_12225);
nand U13401 (N_13401,N_12757,N_12220);
and U13402 (N_13402,N_12003,N_12207);
and U13403 (N_13403,N_12185,N_12353);
or U13404 (N_13404,N_12015,N_12987);
xnor U13405 (N_13405,N_12641,N_12371);
nor U13406 (N_13406,N_12282,N_12700);
nor U13407 (N_13407,N_12915,N_12224);
xor U13408 (N_13408,N_12268,N_12690);
or U13409 (N_13409,N_12828,N_12665);
nand U13410 (N_13410,N_12277,N_12296);
nor U13411 (N_13411,N_12836,N_12009);
nor U13412 (N_13412,N_12747,N_12341);
nor U13413 (N_13413,N_12469,N_12765);
nand U13414 (N_13414,N_12361,N_12106);
nor U13415 (N_13415,N_12773,N_12364);
nor U13416 (N_13416,N_12161,N_12833);
nand U13417 (N_13417,N_12332,N_12022);
or U13418 (N_13418,N_12166,N_12950);
and U13419 (N_13419,N_12903,N_12750);
nor U13420 (N_13420,N_12466,N_12314);
nand U13421 (N_13421,N_12912,N_12890);
or U13422 (N_13422,N_12485,N_12014);
xor U13423 (N_13423,N_12337,N_12672);
and U13424 (N_13424,N_12891,N_12482);
or U13425 (N_13425,N_12350,N_12238);
nand U13426 (N_13426,N_12190,N_12708);
nor U13427 (N_13427,N_12357,N_12613);
nand U13428 (N_13428,N_12601,N_12367);
nand U13429 (N_13429,N_12557,N_12758);
xnor U13430 (N_13430,N_12409,N_12825);
and U13431 (N_13431,N_12582,N_12565);
nand U13432 (N_13432,N_12924,N_12743);
or U13433 (N_13433,N_12902,N_12107);
nor U13434 (N_13434,N_12406,N_12110);
nor U13435 (N_13435,N_12447,N_12154);
and U13436 (N_13436,N_12191,N_12024);
and U13437 (N_13437,N_12957,N_12018);
and U13438 (N_13438,N_12284,N_12201);
xnor U13439 (N_13439,N_12514,N_12122);
nor U13440 (N_13440,N_12054,N_12653);
xnor U13441 (N_13441,N_12093,N_12532);
or U13442 (N_13442,N_12488,N_12404);
nor U13443 (N_13443,N_12011,N_12922);
and U13444 (N_13444,N_12045,N_12673);
xnor U13445 (N_13445,N_12832,N_12771);
nand U13446 (N_13446,N_12621,N_12355);
nor U13447 (N_13447,N_12429,N_12978);
nand U13448 (N_13448,N_12988,N_12115);
xnor U13449 (N_13449,N_12090,N_12727);
or U13450 (N_13450,N_12986,N_12965);
xor U13451 (N_13451,N_12590,N_12094);
nand U13452 (N_13452,N_12078,N_12551);
xnor U13453 (N_13453,N_12617,N_12425);
xnor U13454 (N_13454,N_12678,N_12259);
nand U13455 (N_13455,N_12067,N_12636);
xnor U13456 (N_13456,N_12299,N_12866);
nor U13457 (N_13457,N_12629,N_12880);
xor U13458 (N_13458,N_12144,N_12260);
and U13459 (N_13459,N_12920,N_12421);
or U13460 (N_13460,N_12125,N_12368);
and U13461 (N_13461,N_12325,N_12338);
nor U13462 (N_13462,N_12861,N_12493);
xnor U13463 (N_13463,N_12138,N_12526);
xor U13464 (N_13464,N_12165,N_12588);
nor U13465 (N_13465,N_12216,N_12463);
xor U13466 (N_13466,N_12733,N_12445);
xnor U13467 (N_13467,N_12818,N_12923);
or U13468 (N_13468,N_12600,N_12567);
nand U13469 (N_13469,N_12005,N_12051);
and U13470 (N_13470,N_12900,N_12309);
nor U13471 (N_13471,N_12802,N_12450);
and U13472 (N_13472,N_12261,N_12589);
xnor U13473 (N_13473,N_12979,N_12644);
or U13474 (N_13474,N_12569,N_12948);
nand U13475 (N_13475,N_12215,N_12628);
and U13476 (N_13476,N_12658,N_12898);
nor U13477 (N_13477,N_12740,N_12279);
xor U13478 (N_13478,N_12699,N_12944);
or U13479 (N_13479,N_12712,N_12393);
and U13480 (N_13480,N_12119,N_12479);
xnor U13481 (N_13481,N_12281,N_12859);
nand U13482 (N_13482,N_12852,N_12608);
xnor U13483 (N_13483,N_12612,N_12359);
and U13484 (N_13484,N_12734,N_12707);
xnor U13485 (N_13485,N_12767,N_12827);
nor U13486 (N_13486,N_12816,N_12142);
and U13487 (N_13487,N_12855,N_12999);
nor U13488 (N_13488,N_12193,N_12587);
or U13489 (N_13489,N_12288,N_12385);
nor U13490 (N_13490,N_12823,N_12764);
xnor U13491 (N_13491,N_12741,N_12392);
xor U13492 (N_13492,N_12376,N_12329);
nand U13493 (N_13493,N_12399,N_12901);
nand U13494 (N_13494,N_12990,N_12550);
or U13495 (N_13495,N_12956,N_12655);
or U13496 (N_13496,N_12494,N_12520);
xnor U13497 (N_13497,N_12860,N_12114);
or U13498 (N_13498,N_12805,N_12875);
nand U13499 (N_13499,N_12719,N_12539);
nand U13500 (N_13500,N_12685,N_12406);
xnor U13501 (N_13501,N_12353,N_12386);
nor U13502 (N_13502,N_12185,N_12925);
or U13503 (N_13503,N_12757,N_12108);
xor U13504 (N_13504,N_12527,N_12362);
nand U13505 (N_13505,N_12586,N_12015);
nand U13506 (N_13506,N_12383,N_12709);
nor U13507 (N_13507,N_12858,N_12927);
nor U13508 (N_13508,N_12303,N_12188);
and U13509 (N_13509,N_12140,N_12381);
xnor U13510 (N_13510,N_12048,N_12251);
and U13511 (N_13511,N_12999,N_12335);
and U13512 (N_13512,N_12365,N_12451);
and U13513 (N_13513,N_12192,N_12128);
nor U13514 (N_13514,N_12526,N_12236);
or U13515 (N_13515,N_12161,N_12752);
xnor U13516 (N_13516,N_12480,N_12963);
and U13517 (N_13517,N_12506,N_12665);
and U13518 (N_13518,N_12566,N_12861);
or U13519 (N_13519,N_12489,N_12482);
nor U13520 (N_13520,N_12190,N_12584);
nand U13521 (N_13521,N_12149,N_12416);
nand U13522 (N_13522,N_12469,N_12964);
or U13523 (N_13523,N_12867,N_12740);
and U13524 (N_13524,N_12088,N_12044);
and U13525 (N_13525,N_12578,N_12900);
xnor U13526 (N_13526,N_12075,N_12239);
and U13527 (N_13527,N_12081,N_12100);
nand U13528 (N_13528,N_12990,N_12892);
xor U13529 (N_13529,N_12000,N_12498);
and U13530 (N_13530,N_12543,N_12742);
nor U13531 (N_13531,N_12285,N_12821);
and U13532 (N_13532,N_12578,N_12868);
nand U13533 (N_13533,N_12441,N_12399);
xor U13534 (N_13534,N_12711,N_12853);
or U13535 (N_13535,N_12544,N_12680);
xnor U13536 (N_13536,N_12893,N_12935);
nand U13537 (N_13537,N_12819,N_12095);
nor U13538 (N_13538,N_12521,N_12923);
nor U13539 (N_13539,N_12064,N_12532);
and U13540 (N_13540,N_12623,N_12700);
xnor U13541 (N_13541,N_12775,N_12413);
nor U13542 (N_13542,N_12330,N_12354);
nand U13543 (N_13543,N_12868,N_12576);
nand U13544 (N_13544,N_12126,N_12489);
nor U13545 (N_13545,N_12737,N_12734);
and U13546 (N_13546,N_12759,N_12608);
xnor U13547 (N_13547,N_12219,N_12913);
xnor U13548 (N_13548,N_12746,N_12013);
nor U13549 (N_13549,N_12850,N_12342);
nand U13550 (N_13550,N_12675,N_12152);
and U13551 (N_13551,N_12929,N_12948);
xor U13552 (N_13552,N_12244,N_12695);
nor U13553 (N_13553,N_12080,N_12957);
nand U13554 (N_13554,N_12371,N_12591);
or U13555 (N_13555,N_12808,N_12153);
nor U13556 (N_13556,N_12508,N_12266);
and U13557 (N_13557,N_12885,N_12041);
or U13558 (N_13558,N_12405,N_12156);
or U13559 (N_13559,N_12580,N_12592);
xnor U13560 (N_13560,N_12653,N_12129);
nor U13561 (N_13561,N_12979,N_12016);
xnor U13562 (N_13562,N_12159,N_12283);
or U13563 (N_13563,N_12968,N_12354);
or U13564 (N_13564,N_12569,N_12729);
xnor U13565 (N_13565,N_12837,N_12922);
or U13566 (N_13566,N_12231,N_12317);
nor U13567 (N_13567,N_12484,N_12433);
or U13568 (N_13568,N_12438,N_12808);
and U13569 (N_13569,N_12386,N_12964);
or U13570 (N_13570,N_12053,N_12635);
and U13571 (N_13571,N_12614,N_12474);
nand U13572 (N_13572,N_12249,N_12907);
nor U13573 (N_13573,N_12699,N_12908);
and U13574 (N_13574,N_12003,N_12755);
xnor U13575 (N_13575,N_12472,N_12946);
and U13576 (N_13576,N_12403,N_12064);
nor U13577 (N_13577,N_12481,N_12651);
and U13578 (N_13578,N_12353,N_12106);
nand U13579 (N_13579,N_12905,N_12440);
nand U13580 (N_13580,N_12311,N_12966);
xnor U13581 (N_13581,N_12960,N_12745);
and U13582 (N_13582,N_12822,N_12926);
and U13583 (N_13583,N_12905,N_12804);
nand U13584 (N_13584,N_12639,N_12201);
and U13585 (N_13585,N_12599,N_12908);
and U13586 (N_13586,N_12560,N_12791);
nand U13587 (N_13587,N_12347,N_12093);
xnor U13588 (N_13588,N_12243,N_12007);
or U13589 (N_13589,N_12196,N_12647);
and U13590 (N_13590,N_12054,N_12131);
nand U13591 (N_13591,N_12545,N_12041);
nand U13592 (N_13592,N_12483,N_12937);
nor U13593 (N_13593,N_12452,N_12504);
or U13594 (N_13594,N_12054,N_12571);
or U13595 (N_13595,N_12653,N_12429);
nor U13596 (N_13596,N_12639,N_12577);
and U13597 (N_13597,N_12636,N_12396);
or U13598 (N_13598,N_12782,N_12938);
nor U13599 (N_13599,N_12372,N_12558);
nand U13600 (N_13600,N_12078,N_12622);
or U13601 (N_13601,N_12279,N_12602);
nand U13602 (N_13602,N_12303,N_12748);
nor U13603 (N_13603,N_12223,N_12050);
or U13604 (N_13604,N_12322,N_12433);
nand U13605 (N_13605,N_12709,N_12489);
and U13606 (N_13606,N_12718,N_12364);
and U13607 (N_13607,N_12358,N_12804);
xor U13608 (N_13608,N_12473,N_12178);
nor U13609 (N_13609,N_12512,N_12882);
nand U13610 (N_13610,N_12095,N_12768);
nor U13611 (N_13611,N_12982,N_12116);
xnor U13612 (N_13612,N_12093,N_12070);
or U13613 (N_13613,N_12486,N_12472);
and U13614 (N_13614,N_12915,N_12568);
nand U13615 (N_13615,N_12526,N_12613);
or U13616 (N_13616,N_12326,N_12170);
and U13617 (N_13617,N_12060,N_12996);
and U13618 (N_13618,N_12226,N_12938);
nand U13619 (N_13619,N_12732,N_12912);
and U13620 (N_13620,N_12158,N_12053);
or U13621 (N_13621,N_12500,N_12220);
nor U13622 (N_13622,N_12736,N_12015);
nor U13623 (N_13623,N_12749,N_12805);
nand U13624 (N_13624,N_12317,N_12278);
xor U13625 (N_13625,N_12015,N_12966);
nor U13626 (N_13626,N_12595,N_12065);
and U13627 (N_13627,N_12607,N_12814);
nand U13628 (N_13628,N_12473,N_12345);
nor U13629 (N_13629,N_12650,N_12349);
nor U13630 (N_13630,N_12623,N_12844);
xor U13631 (N_13631,N_12476,N_12447);
xnor U13632 (N_13632,N_12219,N_12328);
xnor U13633 (N_13633,N_12827,N_12103);
nor U13634 (N_13634,N_12147,N_12453);
nor U13635 (N_13635,N_12491,N_12931);
nor U13636 (N_13636,N_12252,N_12481);
xor U13637 (N_13637,N_12292,N_12221);
nand U13638 (N_13638,N_12001,N_12481);
nor U13639 (N_13639,N_12365,N_12924);
nor U13640 (N_13640,N_12848,N_12182);
or U13641 (N_13641,N_12236,N_12576);
nor U13642 (N_13642,N_12113,N_12990);
nand U13643 (N_13643,N_12235,N_12200);
or U13644 (N_13644,N_12862,N_12034);
nor U13645 (N_13645,N_12460,N_12842);
and U13646 (N_13646,N_12834,N_12923);
or U13647 (N_13647,N_12462,N_12793);
xnor U13648 (N_13648,N_12583,N_12491);
xnor U13649 (N_13649,N_12549,N_12315);
or U13650 (N_13650,N_12171,N_12438);
nand U13651 (N_13651,N_12160,N_12310);
nand U13652 (N_13652,N_12463,N_12237);
and U13653 (N_13653,N_12111,N_12446);
nand U13654 (N_13654,N_12930,N_12276);
and U13655 (N_13655,N_12477,N_12057);
or U13656 (N_13656,N_12215,N_12799);
nand U13657 (N_13657,N_12632,N_12889);
or U13658 (N_13658,N_12281,N_12379);
or U13659 (N_13659,N_12814,N_12841);
nor U13660 (N_13660,N_12323,N_12300);
nor U13661 (N_13661,N_12520,N_12033);
nor U13662 (N_13662,N_12605,N_12880);
xor U13663 (N_13663,N_12766,N_12159);
nor U13664 (N_13664,N_12933,N_12977);
and U13665 (N_13665,N_12843,N_12528);
or U13666 (N_13666,N_12355,N_12931);
or U13667 (N_13667,N_12532,N_12670);
or U13668 (N_13668,N_12931,N_12016);
xor U13669 (N_13669,N_12756,N_12894);
nand U13670 (N_13670,N_12325,N_12598);
xor U13671 (N_13671,N_12400,N_12369);
and U13672 (N_13672,N_12802,N_12348);
and U13673 (N_13673,N_12207,N_12037);
and U13674 (N_13674,N_12853,N_12271);
xor U13675 (N_13675,N_12692,N_12072);
or U13676 (N_13676,N_12507,N_12564);
nor U13677 (N_13677,N_12694,N_12747);
xnor U13678 (N_13678,N_12775,N_12798);
nor U13679 (N_13679,N_12521,N_12821);
or U13680 (N_13680,N_12707,N_12097);
or U13681 (N_13681,N_12322,N_12323);
or U13682 (N_13682,N_12680,N_12746);
nor U13683 (N_13683,N_12796,N_12854);
nor U13684 (N_13684,N_12223,N_12081);
xnor U13685 (N_13685,N_12893,N_12388);
xnor U13686 (N_13686,N_12640,N_12922);
nor U13687 (N_13687,N_12026,N_12630);
and U13688 (N_13688,N_12023,N_12946);
or U13689 (N_13689,N_12404,N_12377);
nor U13690 (N_13690,N_12207,N_12759);
nand U13691 (N_13691,N_12639,N_12517);
xnor U13692 (N_13692,N_12885,N_12008);
and U13693 (N_13693,N_12870,N_12727);
nor U13694 (N_13694,N_12681,N_12981);
or U13695 (N_13695,N_12670,N_12167);
nor U13696 (N_13696,N_12363,N_12328);
xor U13697 (N_13697,N_12348,N_12440);
or U13698 (N_13698,N_12909,N_12117);
nor U13699 (N_13699,N_12733,N_12810);
xnor U13700 (N_13700,N_12390,N_12208);
and U13701 (N_13701,N_12405,N_12546);
nand U13702 (N_13702,N_12854,N_12325);
nand U13703 (N_13703,N_12276,N_12072);
nor U13704 (N_13704,N_12009,N_12809);
xnor U13705 (N_13705,N_12935,N_12547);
xnor U13706 (N_13706,N_12779,N_12317);
nand U13707 (N_13707,N_12798,N_12393);
nor U13708 (N_13708,N_12228,N_12362);
and U13709 (N_13709,N_12915,N_12290);
and U13710 (N_13710,N_12265,N_12078);
or U13711 (N_13711,N_12082,N_12799);
nand U13712 (N_13712,N_12013,N_12596);
or U13713 (N_13713,N_12675,N_12021);
xor U13714 (N_13714,N_12873,N_12053);
xnor U13715 (N_13715,N_12420,N_12714);
nor U13716 (N_13716,N_12665,N_12596);
and U13717 (N_13717,N_12447,N_12264);
nand U13718 (N_13718,N_12546,N_12357);
or U13719 (N_13719,N_12453,N_12267);
xor U13720 (N_13720,N_12804,N_12040);
xor U13721 (N_13721,N_12173,N_12082);
xor U13722 (N_13722,N_12113,N_12373);
xnor U13723 (N_13723,N_12730,N_12903);
or U13724 (N_13724,N_12887,N_12809);
nor U13725 (N_13725,N_12762,N_12541);
nor U13726 (N_13726,N_12093,N_12374);
or U13727 (N_13727,N_12452,N_12823);
or U13728 (N_13728,N_12913,N_12847);
and U13729 (N_13729,N_12455,N_12175);
nor U13730 (N_13730,N_12906,N_12480);
nand U13731 (N_13731,N_12657,N_12119);
nor U13732 (N_13732,N_12093,N_12057);
and U13733 (N_13733,N_12688,N_12406);
or U13734 (N_13734,N_12663,N_12453);
nor U13735 (N_13735,N_12527,N_12571);
or U13736 (N_13736,N_12876,N_12978);
xnor U13737 (N_13737,N_12712,N_12699);
nand U13738 (N_13738,N_12448,N_12946);
and U13739 (N_13739,N_12618,N_12245);
xnor U13740 (N_13740,N_12894,N_12510);
or U13741 (N_13741,N_12460,N_12205);
nand U13742 (N_13742,N_12180,N_12219);
or U13743 (N_13743,N_12635,N_12313);
xor U13744 (N_13744,N_12191,N_12200);
and U13745 (N_13745,N_12064,N_12302);
and U13746 (N_13746,N_12959,N_12318);
or U13747 (N_13747,N_12401,N_12230);
nor U13748 (N_13748,N_12762,N_12507);
or U13749 (N_13749,N_12581,N_12901);
and U13750 (N_13750,N_12442,N_12832);
or U13751 (N_13751,N_12426,N_12695);
and U13752 (N_13752,N_12842,N_12567);
xnor U13753 (N_13753,N_12290,N_12997);
or U13754 (N_13754,N_12789,N_12398);
or U13755 (N_13755,N_12452,N_12812);
xor U13756 (N_13756,N_12431,N_12809);
nand U13757 (N_13757,N_12448,N_12727);
or U13758 (N_13758,N_12843,N_12624);
or U13759 (N_13759,N_12077,N_12323);
or U13760 (N_13760,N_12438,N_12554);
nor U13761 (N_13761,N_12502,N_12424);
nor U13762 (N_13762,N_12677,N_12608);
nor U13763 (N_13763,N_12398,N_12625);
nand U13764 (N_13764,N_12485,N_12043);
and U13765 (N_13765,N_12442,N_12836);
or U13766 (N_13766,N_12617,N_12865);
nor U13767 (N_13767,N_12310,N_12589);
or U13768 (N_13768,N_12972,N_12069);
xnor U13769 (N_13769,N_12608,N_12401);
nor U13770 (N_13770,N_12751,N_12954);
nand U13771 (N_13771,N_12685,N_12094);
nand U13772 (N_13772,N_12724,N_12738);
and U13773 (N_13773,N_12487,N_12567);
or U13774 (N_13774,N_12476,N_12727);
and U13775 (N_13775,N_12130,N_12519);
nor U13776 (N_13776,N_12273,N_12033);
nand U13777 (N_13777,N_12061,N_12762);
xnor U13778 (N_13778,N_12030,N_12681);
xor U13779 (N_13779,N_12702,N_12905);
nor U13780 (N_13780,N_12388,N_12544);
nand U13781 (N_13781,N_12263,N_12374);
or U13782 (N_13782,N_12508,N_12946);
or U13783 (N_13783,N_12768,N_12644);
and U13784 (N_13784,N_12576,N_12465);
xnor U13785 (N_13785,N_12458,N_12957);
nor U13786 (N_13786,N_12466,N_12706);
nor U13787 (N_13787,N_12651,N_12007);
nor U13788 (N_13788,N_12311,N_12516);
or U13789 (N_13789,N_12417,N_12101);
and U13790 (N_13790,N_12340,N_12508);
nor U13791 (N_13791,N_12119,N_12005);
and U13792 (N_13792,N_12172,N_12608);
and U13793 (N_13793,N_12771,N_12712);
nand U13794 (N_13794,N_12848,N_12960);
and U13795 (N_13795,N_12079,N_12143);
nor U13796 (N_13796,N_12368,N_12200);
or U13797 (N_13797,N_12240,N_12470);
or U13798 (N_13798,N_12133,N_12442);
nand U13799 (N_13799,N_12960,N_12409);
and U13800 (N_13800,N_12246,N_12547);
xnor U13801 (N_13801,N_12733,N_12518);
or U13802 (N_13802,N_12635,N_12469);
and U13803 (N_13803,N_12622,N_12924);
nand U13804 (N_13804,N_12980,N_12256);
and U13805 (N_13805,N_12333,N_12039);
xnor U13806 (N_13806,N_12840,N_12610);
and U13807 (N_13807,N_12251,N_12836);
xnor U13808 (N_13808,N_12794,N_12609);
xor U13809 (N_13809,N_12708,N_12104);
nor U13810 (N_13810,N_12921,N_12528);
nor U13811 (N_13811,N_12558,N_12182);
nor U13812 (N_13812,N_12959,N_12385);
or U13813 (N_13813,N_12417,N_12895);
nand U13814 (N_13814,N_12799,N_12000);
nor U13815 (N_13815,N_12246,N_12649);
or U13816 (N_13816,N_12021,N_12063);
and U13817 (N_13817,N_12319,N_12355);
or U13818 (N_13818,N_12800,N_12588);
nor U13819 (N_13819,N_12096,N_12050);
xor U13820 (N_13820,N_12864,N_12095);
and U13821 (N_13821,N_12269,N_12478);
nor U13822 (N_13822,N_12772,N_12785);
and U13823 (N_13823,N_12032,N_12047);
nand U13824 (N_13824,N_12891,N_12642);
nor U13825 (N_13825,N_12551,N_12607);
xor U13826 (N_13826,N_12902,N_12991);
and U13827 (N_13827,N_12325,N_12318);
nand U13828 (N_13828,N_12974,N_12764);
or U13829 (N_13829,N_12852,N_12876);
xnor U13830 (N_13830,N_12039,N_12785);
and U13831 (N_13831,N_12863,N_12026);
and U13832 (N_13832,N_12477,N_12892);
or U13833 (N_13833,N_12984,N_12058);
nor U13834 (N_13834,N_12938,N_12526);
nand U13835 (N_13835,N_12367,N_12804);
nand U13836 (N_13836,N_12265,N_12397);
nor U13837 (N_13837,N_12823,N_12130);
xor U13838 (N_13838,N_12888,N_12812);
nand U13839 (N_13839,N_12721,N_12499);
xor U13840 (N_13840,N_12140,N_12166);
or U13841 (N_13841,N_12128,N_12969);
nand U13842 (N_13842,N_12696,N_12669);
nor U13843 (N_13843,N_12722,N_12457);
nand U13844 (N_13844,N_12965,N_12890);
or U13845 (N_13845,N_12325,N_12385);
nor U13846 (N_13846,N_12156,N_12487);
or U13847 (N_13847,N_12519,N_12620);
nand U13848 (N_13848,N_12347,N_12763);
nor U13849 (N_13849,N_12292,N_12668);
and U13850 (N_13850,N_12082,N_12271);
nor U13851 (N_13851,N_12077,N_12036);
xnor U13852 (N_13852,N_12193,N_12876);
nand U13853 (N_13853,N_12210,N_12024);
nand U13854 (N_13854,N_12376,N_12485);
nand U13855 (N_13855,N_12690,N_12659);
or U13856 (N_13856,N_12738,N_12019);
and U13857 (N_13857,N_12294,N_12049);
xnor U13858 (N_13858,N_12738,N_12451);
nor U13859 (N_13859,N_12255,N_12197);
nor U13860 (N_13860,N_12901,N_12830);
nand U13861 (N_13861,N_12164,N_12476);
xor U13862 (N_13862,N_12925,N_12640);
nand U13863 (N_13863,N_12466,N_12327);
and U13864 (N_13864,N_12564,N_12513);
nand U13865 (N_13865,N_12618,N_12911);
and U13866 (N_13866,N_12554,N_12317);
xor U13867 (N_13867,N_12225,N_12941);
and U13868 (N_13868,N_12857,N_12714);
nor U13869 (N_13869,N_12309,N_12477);
or U13870 (N_13870,N_12093,N_12585);
nand U13871 (N_13871,N_12084,N_12144);
xnor U13872 (N_13872,N_12196,N_12327);
xor U13873 (N_13873,N_12101,N_12074);
and U13874 (N_13874,N_12335,N_12763);
and U13875 (N_13875,N_12723,N_12406);
nor U13876 (N_13876,N_12593,N_12012);
and U13877 (N_13877,N_12334,N_12035);
or U13878 (N_13878,N_12663,N_12614);
nor U13879 (N_13879,N_12478,N_12427);
xor U13880 (N_13880,N_12588,N_12954);
nand U13881 (N_13881,N_12388,N_12916);
xor U13882 (N_13882,N_12028,N_12383);
xnor U13883 (N_13883,N_12186,N_12259);
nor U13884 (N_13884,N_12997,N_12540);
and U13885 (N_13885,N_12044,N_12950);
and U13886 (N_13886,N_12396,N_12833);
nor U13887 (N_13887,N_12435,N_12130);
or U13888 (N_13888,N_12069,N_12909);
xnor U13889 (N_13889,N_12040,N_12180);
nand U13890 (N_13890,N_12161,N_12802);
or U13891 (N_13891,N_12655,N_12405);
or U13892 (N_13892,N_12177,N_12308);
nand U13893 (N_13893,N_12820,N_12864);
nor U13894 (N_13894,N_12844,N_12116);
nor U13895 (N_13895,N_12301,N_12848);
and U13896 (N_13896,N_12604,N_12864);
nand U13897 (N_13897,N_12589,N_12847);
xnor U13898 (N_13898,N_12279,N_12901);
or U13899 (N_13899,N_12785,N_12774);
and U13900 (N_13900,N_12558,N_12408);
nand U13901 (N_13901,N_12263,N_12074);
xnor U13902 (N_13902,N_12408,N_12427);
nand U13903 (N_13903,N_12322,N_12017);
nor U13904 (N_13904,N_12817,N_12314);
nand U13905 (N_13905,N_12677,N_12773);
or U13906 (N_13906,N_12666,N_12864);
nor U13907 (N_13907,N_12526,N_12107);
or U13908 (N_13908,N_12703,N_12840);
nand U13909 (N_13909,N_12353,N_12340);
nor U13910 (N_13910,N_12771,N_12776);
or U13911 (N_13911,N_12126,N_12067);
xnor U13912 (N_13912,N_12009,N_12558);
and U13913 (N_13913,N_12918,N_12097);
and U13914 (N_13914,N_12872,N_12431);
xnor U13915 (N_13915,N_12752,N_12154);
and U13916 (N_13916,N_12847,N_12119);
nor U13917 (N_13917,N_12814,N_12852);
nor U13918 (N_13918,N_12498,N_12469);
or U13919 (N_13919,N_12034,N_12832);
nor U13920 (N_13920,N_12470,N_12839);
nor U13921 (N_13921,N_12497,N_12263);
nand U13922 (N_13922,N_12471,N_12269);
nand U13923 (N_13923,N_12322,N_12215);
nand U13924 (N_13924,N_12825,N_12548);
xor U13925 (N_13925,N_12040,N_12235);
xor U13926 (N_13926,N_12143,N_12711);
nand U13927 (N_13927,N_12777,N_12885);
nand U13928 (N_13928,N_12139,N_12597);
nand U13929 (N_13929,N_12787,N_12405);
nor U13930 (N_13930,N_12176,N_12298);
or U13931 (N_13931,N_12452,N_12038);
xnor U13932 (N_13932,N_12888,N_12818);
nor U13933 (N_13933,N_12605,N_12018);
and U13934 (N_13934,N_12503,N_12886);
nor U13935 (N_13935,N_12872,N_12875);
and U13936 (N_13936,N_12795,N_12569);
nand U13937 (N_13937,N_12941,N_12059);
nand U13938 (N_13938,N_12819,N_12007);
nor U13939 (N_13939,N_12942,N_12039);
nor U13940 (N_13940,N_12999,N_12006);
nor U13941 (N_13941,N_12209,N_12178);
nand U13942 (N_13942,N_12491,N_12593);
or U13943 (N_13943,N_12326,N_12736);
and U13944 (N_13944,N_12468,N_12890);
nor U13945 (N_13945,N_12418,N_12289);
nand U13946 (N_13946,N_12344,N_12871);
and U13947 (N_13947,N_12987,N_12389);
xor U13948 (N_13948,N_12124,N_12676);
and U13949 (N_13949,N_12222,N_12183);
nand U13950 (N_13950,N_12648,N_12496);
or U13951 (N_13951,N_12813,N_12277);
xor U13952 (N_13952,N_12742,N_12876);
nor U13953 (N_13953,N_12143,N_12697);
and U13954 (N_13954,N_12303,N_12317);
or U13955 (N_13955,N_12777,N_12311);
and U13956 (N_13956,N_12510,N_12769);
or U13957 (N_13957,N_12561,N_12254);
nand U13958 (N_13958,N_12312,N_12679);
xor U13959 (N_13959,N_12532,N_12405);
nand U13960 (N_13960,N_12055,N_12933);
or U13961 (N_13961,N_12885,N_12489);
xnor U13962 (N_13962,N_12963,N_12933);
and U13963 (N_13963,N_12477,N_12574);
nand U13964 (N_13964,N_12969,N_12817);
or U13965 (N_13965,N_12902,N_12156);
or U13966 (N_13966,N_12793,N_12118);
or U13967 (N_13967,N_12816,N_12753);
xor U13968 (N_13968,N_12475,N_12109);
nor U13969 (N_13969,N_12163,N_12656);
and U13970 (N_13970,N_12782,N_12985);
and U13971 (N_13971,N_12462,N_12248);
or U13972 (N_13972,N_12545,N_12519);
and U13973 (N_13973,N_12563,N_12248);
xnor U13974 (N_13974,N_12022,N_12211);
nand U13975 (N_13975,N_12715,N_12732);
and U13976 (N_13976,N_12951,N_12394);
xor U13977 (N_13977,N_12251,N_12386);
nand U13978 (N_13978,N_12787,N_12671);
xor U13979 (N_13979,N_12523,N_12159);
nand U13980 (N_13980,N_12675,N_12089);
nand U13981 (N_13981,N_12634,N_12664);
nor U13982 (N_13982,N_12923,N_12202);
and U13983 (N_13983,N_12848,N_12396);
and U13984 (N_13984,N_12374,N_12020);
or U13985 (N_13985,N_12789,N_12216);
nor U13986 (N_13986,N_12992,N_12742);
nor U13987 (N_13987,N_12625,N_12809);
nor U13988 (N_13988,N_12691,N_12374);
nand U13989 (N_13989,N_12843,N_12802);
nand U13990 (N_13990,N_12583,N_12842);
nor U13991 (N_13991,N_12954,N_12770);
xor U13992 (N_13992,N_12251,N_12252);
xnor U13993 (N_13993,N_12755,N_12266);
and U13994 (N_13994,N_12194,N_12372);
and U13995 (N_13995,N_12250,N_12530);
and U13996 (N_13996,N_12113,N_12406);
nand U13997 (N_13997,N_12408,N_12055);
nand U13998 (N_13998,N_12323,N_12204);
or U13999 (N_13999,N_12882,N_12879);
nor U14000 (N_14000,N_13355,N_13064);
nand U14001 (N_14001,N_13550,N_13472);
and U14002 (N_14002,N_13818,N_13216);
nor U14003 (N_14003,N_13959,N_13704);
xnor U14004 (N_14004,N_13688,N_13175);
or U14005 (N_14005,N_13249,N_13880);
xor U14006 (N_14006,N_13419,N_13933);
nor U14007 (N_14007,N_13821,N_13320);
xor U14008 (N_14008,N_13133,N_13727);
nand U14009 (N_14009,N_13324,N_13083);
and U14010 (N_14010,N_13847,N_13383);
nand U14011 (N_14011,N_13609,N_13327);
nand U14012 (N_14012,N_13108,N_13889);
or U14013 (N_14013,N_13358,N_13316);
xnor U14014 (N_14014,N_13598,N_13370);
xnor U14015 (N_14015,N_13604,N_13169);
nand U14016 (N_14016,N_13984,N_13855);
and U14017 (N_14017,N_13339,N_13899);
nor U14018 (N_14018,N_13375,N_13253);
and U14019 (N_14019,N_13707,N_13329);
nand U14020 (N_14020,N_13399,N_13605);
and U14021 (N_14021,N_13271,N_13751);
or U14022 (N_14022,N_13241,N_13754);
xnor U14023 (N_14023,N_13051,N_13693);
and U14024 (N_14024,N_13166,N_13495);
nand U14025 (N_14025,N_13384,N_13745);
nor U14026 (N_14026,N_13022,N_13357);
nand U14027 (N_14027,N_13513,N_13703);
and U14028 (N_14028,N_13917,N_13671);
and U14029 (N_14029,N_13740,N_13217);
xnor U14030 (N_14030,N_13819,N_13619);
and U14031 (N_14031,N_13924,N_13647);
and U14032 (N_14032,N_13877,N_13502);
xnor U14033 (N_14033,N_13045,N_13509);
xor U14034 (N_14034,N_13638,N_13052);
and U14035 (N_14035,N_13909,N_13637);
xor U14036 (N_14036,N_13603,N_13061);
nor U14037 (N_14037,N_13247,N_13120);
nor U14038 (N_14038,N_13866,N_13049);
nor U14039 (N_14039,N_13627,N_13853);
xor U14040 (N_14040,N_13107,N_13258);
nand U14041 (N_14041,N_13835,N_13769);
xor U14042 (N_14042,N_13245,N_13705);
nand U14043 (N_14043,N_13028,N_13572);
and U14044 (N_14044,N_13838,N_13742);
xor U14045 (N_14045,N_13471,N_13006);
nand U14046 (N_14046,N_13568,N_13070);
nor U14047 (N_14047,N_13189,N_13158);
xor U14048 (N_14048,N_13341,N_13687);
or U14049 (N_14049,N_13306,N_13515);
or U14050 (N_14050,N_13228,N_13338);
nor U14051 (N_14051,N_13611,N_13369);
nor U14052 (N_14052,N_13330,N_13012);
nor U14053 (N_14053,N_13165,N_13564);
and U14054 (N_14054,N_13171,N_13451);
nor U14055 (N_14055,N_13673,N_13981);
or U14056 (N_14056,N_13709,N_13719);
nor U14057 (N_14057,N_13825,N_13672);
nand U14058 (N_14058,N_13788,N_13718);
nor U14059 (N_14059,N_13469,N_13063);
and U14060 (N_14060,N_13039,N_13473);
xor U14061 (N_14061,N_13391,N_13987);
nand U14062 (N_14062,N_13440,N_13577);
and U14063 (N_14063,N_13967,N_13467);
nand U14064 (N_14064,N_13438,N_13633);
nand U14065 (N_14065,N_13490,N_13335);
nor U14066 (N_14066,N_13277,N_13177);
and U14067 (N_14067,N_13616,N_13027);
nor U14068 (N_14068,N_13965,N_13411);
nand U14069 (N_14069,N_13274,N_13916);
or U14070 (N_14070,N_13717,N_13910);
and U14071 (N_14071,N_13920,N_13958);
nor U14072 (N_14072,N_13413,N_13793);
xor U14073 (N_14073,N_13592,N_13626);
xnor U14074 (N_14074,N_13903,N_13199);
nor U14075 (N_14075,N_13945,N_13852);
or U14076 (N_14076,N_13173,N_13016);
or U14077 (N_14077,N_13864,N_13677);
xnor U14078 (N_14078,N_13506,N_13313);
and U14079 (N_14079,N_13914,N_13535);
xor U14080 (N_14080,N_13090,N_13284);
nor U14081 (N_14081,N_13919,N_13681);
or U14082 (N_14082,N_13311,N_13906);
nand U14083 (N_14083,N_13779,N_13486);
nand U14084 (N_14084,N_13966,N_13393);
and U14085 (N_14085,N_13174,N_13820);
xnor U14086 (N_14086,N_13887,N_13511);
xor U14087 (N_14087,N_13492,N_13547);
nand U14088 (N_14088,N_13724,N_13214);
xor U14089 (N_14089,N_13305,N_13892);
nand U14090 (N_14090,N_13433,N_13470);
and U14091 (N_14091,N_13043,N_13979);
xnor U14092 (N_14092,N_13430,N_13303);
xnor U14093 (N_14093,N_13566,N_13757);
nor U14094 (N_14094,N_13344,N_13334);
nor U14095 (N_14095,N_13787,N_13901);
nand U14096 (N_14096,N_13215,N_13168);
nand U14097 (N_14097,N_13992,N_13435);
and U14098 (N_14098,N_13222,N_13362);
nor U14099 (N_14099,N_13239,N_13332);
nor U14100 (N_14100,N_13813,N_13553);
xor U14101 (N_14101,N_13921,N_13696);
and U14102 (N_14102,N_13071,N_13744);
xnor U14103 (N_14103,N_13570,N_13285);
or U14104 (N_14104,N_13477,N_13831);
nand U14105 (N_14105,N_13099,N_13695);
and U14106 (N_14106,N_13498,N_13651);
or U14107 (N_14107,N_13101,N_13885);
and U14108 (N_14108,N_13066,N_13573);
nor U14109 (N_14109,N_13985,N_13653);
and U14110 (N_14110,N_13003,N_13333);
nand U14111 (N_14111,N_13770,N_13888);
xor U14112 (N_14112,N_13129,N_13237);
or U14113 (N_14113,N_13663,N_13102);
and U14114 (N_14114,N_13211,N_13118);
nor U14115 (N_14115,N_13698,N_13366);
or U14116 (N_14116,N_13947,N_13230);
or U14117 (N_14117,N_13345,N_13229);
or U14118 (N_14118,N_13977,N_13036);
or U14119 (N_14119,N_13762,N_13008);
and U14120 (N_14120,N_13635,N_13447);
or U14121 (N_14121,N_13731,N_13454);
nand U14122 (N_14122,N_13541,N_13581);
and U14123 (N_14123,N_13319,N_13233);
and U14124 (N_14124,N_13658,N_13849);
nor U14125 (N_14125,N_13312,N_13579);
nor U14126 (N_14126,N_13092,N_13210);
nand U14127 (N_14127,N_13105,N_13364);
or U14128 (N_14128,N_13766,N_13878);
nor U14129 (N_14129,N_13523,N_13014);
or U14130 (N_14130,N_13645,N_13331);
and U14131 (N_14131,N_13997,N_13278);
or U14132 (N_14132,N_13797,N_13396);
nor U14133 (N_14133,N_13857,N_13976);
nand U14134 (N_14134,N_13656,N_13529);
and U14135 (N_14135,N_13531,N_13085);
xor U14136 (N_14136,N_13466,N_13532);
nor U14137 (N_14137,N_13244,N_13336);
or U14138 (N_14138,N_13072,N_13408);
nand U14139 (N_14139,N_13373,N_13374);
or U14140 (N_14140,N_13346,N_13046);
and U14141 (N_14141,N_13275,N_13980);
and U14142 (N_14142,N_13881,N_13743);
or U14143 (N_14143,N_13716,N_13771);
xnor U14144 (N_14144,N_13096,N_13939);
xnor U14145 (N_14145,N_13053,N_13748);
nor U14146 (N_14146,N_13227,N_13879);
nand U14147 (N_14147,N_13426,N_13208);
and U14148 (N_14148,N_13936,N_13248);
nor U14149 (N_14149,N_13512,N_13734);
nor U14150 (N_14150,N_13415,N_13802);
and U14151 (N_14151,N_13224,N_13025);
and U14152 (N_14152,N_13429,N_13600);
xor U14153 (N_14153,N_13584,N_13272);
or U14154 (N_14154,N_13033,N_13670);
and U14155 (N_14155,N_13462,N_13507);
and U14156 (N_14156,N_13388,N_13442);
nor U14157 (N_14157,N_13680,N_13406);
nand U14158 (N_14158,N_13519,N_13389);
xor U14159 (N_14159,N_13928,N_13843);
or U14160 (N_14160,N_13870,N_13679);
xor U14161 (N_14161,N_13824,N_13178);
nor U14162 (N_14162,N_13259,N_13463);
or U14163 (N_14163,N_13407,N_13126);
xor U14164 (N_14164,N_13546,N_13814);
xnor U14165 (N_14165,N_13262,N_13112);
or U14166 (N_14166,N_13994,N_13382);
and U14167 (N_14167,N_13543,N_13202);
nand U14168 (N_14168,N_13733,N_13706);
nor U14169 (N_14169,N_13200,N_13646);
and U14170 (N_14170,N_13701,N_13464);
nor U14171 (N_14171,N_13434,N_13405);
nor U14172 (N_14172,N_13642,N_13869);
xnor U14173 (N_14173,N_13806,N_13154);
nor U14174 (N_14174,N_13489,N_13685);
xnor U14175 (N_14175,N_13895,N_13162);
or U14176 (N_14176,N_13951,N_13386);
or U14177 (N_14177,N_13678,N_13078);
or U14178 (N_14178,N_13268,N_13134);
nor U14179 (N_14179,N_13503,N_13141);
or U14180 (N_14180,N_13574,N_13193);
and U14181 (N_14181,N_13035,N_13161);
xor U14182 (N_14182,N_13093,N_13381);
nand U14183 (N_14183,N_13534,N_13865);
nor U14184 (N_14184,N_13428,N_13636);
xor U14185 (N_14185,N_13796,N_13774);
nand U14186 (N_14186,N_13628,N_13088);
nor U14187 (N_14187,N_13952,N_13504);
nor U14188 (N_14188,N_13385,N_13363);
nand U14189 (N_14189,N_13896,N_13893);
nand U14190 (N_14190,N_13606,N_13905);
nor U14191 (N_14191,N_13423,N_13772);
and U14192 (N_14192,N_13368,N_13516);
xor U14193 (N_14193,N_13739,N_13974);
nor U14194 (N_14194,N_13279,N_13163);
xor U14195 (N_14195,N_13964,N_13076);
or U14196 (N_14196,N_13932,N_13292);
or U14197 (N_14197,N_13474,N_13062);
nor U14198 (N_14198,N_13294,N_13493);
xor U14199 (N_14199,N_13048,N_13069);
nor U14200 (N_14200,N_13295,N_13290);
nor U14201 (N_14201,N_13167,N_13710);
and U14202 (N_14202,N_13218,N_13747);
nand U14203 (N_14203,N_13721,N_13595);
nor U14204 (N_14204,N_13378,N_13569);
and U14205 (N_14205,N_13019,N_13293);
nand U14206 (N_14206,N_13722,N_13439);
or U14207 (N_14207,N_13223,N_13197);
xnor U14208 (N_14208,N_13459,N_13833);
xor U14209 (N_14209,N_13669,N_13587);
nand U14210 (N_14210,N_13115,N_13773);
nor U14211 (N_14211,N_13170,N_13675);
nor U14212 (N_14212,N_13927,N_13962);
nand U14213 (N_14213,N_13191,N_13020);
xor U14214 (N_14214,N_13392,N_13394);
nand U14215 (N_14215,N_13668,N_13851);
nand U14216 (N_14216,N_13926,N_13314);
nand U14217 (N_14217,N_13940,N_13876);
nor U14218 (N_14218,N_13827,N_13556);
nand U14219 (N_14219,N_13360,N_13956);
nand U14220 (N_14220,N_13094,N_13525);
and U14221 (N_14221,N_13084,N_13047);
nand U14222 (N_14222,N_13823,N_13460);
nand U14223 (N_14223,N_13361,N_13077);
or U14224 (N_14224,N_13784,N_13037);
or U14225 (N_14225,N_13270,N_13883);
and U14226 (N_14226,N_13728,N_13978);
and U14227 (N_14227,N_13975,N_13983);
and U14228 (N_14228,N_13255,N_13941);
and U14229 (N_14229,N_13181,N_13242);
or U14230 (N_14230,N_13643,N_13453);
or U14231 (N_14231,N_13436,N_13289);
nand U14232 (N_14232,N_13667,N_13597);
and U14233 (N_14233,N_13935,N_13192);
nand U14234 (N_14234,N_13617,N_13923);
nor U14235 (N_14235,N_13480,N_13220);
nand U14236 (N_14236,N_13449,N_13702);
and U14237 (N_14237,N_13351,N_13195);
nor U14238 (N_14238,N_13252,N_13356);
or U14239 (N_14239,N_13452,N_13723);
or U14240 (N_14240,N_13794,N_13682);
or U14241 (N_14241,N_13184,N_13836);
xor U14242 (N_14242,N_13982,N_13807);
or U14243 (N_14243,N_13136,N_13528);
or U14244 (N_14244,N_13148,N_13376);
and U14245 (N_14245,N_13159,N_13686);
and U14246 (N_14246,N_13652,N_13476);
nor U14247 (N_14247,N_13666,N_13575);
nor U14248 (N_14248,N_13571,N_13768);
or U14249 (N_14249,N_13427,N_13634);
nor U14250 (N_14250,N_13999,N_13082);
xnor U14251 (N_14251,N_13953,N_13055);
nor U14252 (N_14252,N_13790,N_13432);
or U14253 (N_14253,N_13726,N_13585);
nor U14254 (N_14254,N_13894,N_13755);
or U14255 (N_14255,N_13131,N_13044);
and U14256 (N_14256,N_13461,N_13030);
and U14257 (N_14257,N_13315,N_13783);
nand U14258 (N_14258,N_13805,N_13801);
xor U14259 (N_14259,N_13741,N_13100);
and U14260 (N_14260,N_13538,N_13445);
and U14261 (N_14261,N_13955,N_13536);
nand U14262 (N_14262,N_13589,N_13815);
xor U14263 (N_14263,N_13552,N_13132);
nor U14264 (N_14264,N_13545,N_13913);
or U14265 (N_14265,N_13343,N_13380);
xor U14266 (N_14266,N_13563,N_13950);
nand U14267 (N_14267,N_13139,N_13826);
or U14268 (N_14268,N_13699,N_13013);
or U14269 (N_14269,N_13557,N_13152);
xnor U14270 (N_14270,N_13146,N_13468);
nor U14271 (N_14271,N_13455,N_13138);
or U14272 (N_14272,N_13720,N_13684);
nand U14273 (N_14273,N_13127,N_13778);
or U14274 (N_14274,N_13613,N_13310);
or U14275 (N_14275,N_13007,N_13904);
or U14276 (N_14276,N_13714,N_13238);
xor U14277 (N_14277,N_13157,N_13273);
and U14278 (N_14278,N_13004,N_13861);
nand U14279 (N_14279,N_13322,N_13845);
and U14280 (N_14280,N_13488,N_13123);
or U14281 (N_14281,N_13402,N_13232);
nor U14282 (N_14282,N_13288,N_13204);
xor U14283 (N_14283,N_13086,N_13860);
nand U14284 (N_14284,N_13697,N_13122);
nand U14285 (N_14285,N_13444,N_13015);
and U14286 (N_14286,N_13113,N_13095);
and U14287 (N_14287,N_13097,N_13961);
nor U14288 (N_14288,N_13321,N_13811);
nor U14289 (N_14289,N_13863,N_13834);
or U14290 (N_14290,N_13610,N_13588);
nor U14291 (N_14291,N_13567,N_13337);
and U14292 (N_14292,N_13009,N_13297);
xnor U14293 (N_14293,N_13622,N_13871);
or U14294 (N_14294,N_13882,N_13180);
nand U14295 (N_14295,N_13185,N_13624);
and U14296 (N_14296,N_13261,N_13657);
or U14297 (N_14297,N_13998,N_13712);
or U14298 (N_14298,N_13265,N_13856);
and U14299 (N_14299,N_13347,N_13664);
nand U14300 (N_14300,N_13282,N_13257);
nand U14301 (N_14301,N_13114,N_13812);
xnor U14302 (N_14302,N_13993,N_13188);
and U14303 (N_14303,N_13365,N_13140);
and U14304 (N_14304,N_13450,N_13342);
or U14305 (N_14305,N_13164,N_13810);
nor U14306 (N_14306,N_13874,N_13533);
xor U14307 (N_14307,N_13789,N_13260);
nor U14308 (N_14308,N_13011,N_13377);
nor U14309 (N_14309,N_13886,N_13350);
nand U14310 (N_14310,N_13304,N_13640);
nor U14311 (N_14311,N_13608,N_13510);
nor U14312 (N_14312,N_13130,N_13483);
or U14313 (N_14313,N_13649,N_13829);
nand U14314 (N_14314,N_13264,N_13425);
nor U14315 (N_14315,N_13986,N_13946);
xor U14316 (N_14316,N_13963,N_13119);
xor U14317 (N_14317,N_13087,N_13943);
and U14318 (N_14318,N_13352,N_13186);
nor U14319 (N_14319,N_13848,N_13340);
nor U14320 (N_14320,N_13729,N_13816);
xor U14321 (N_14321,N_13944,N_13026);
and U14322 (N_14322,N_13795,N_13738);
xor U14323 (N_14323,N_13465,N_13074);
and U14324 (N_14324,N_13558,N_13073);
and U14325 (N_14325,N_13508,N_13650);
nand U14326 (N_14326,N_13367,N_13151);
nor U14327 (N_14327,N_13854,N_13555);
and U14328 (N_14328,N_13032,N_13050);
nor U14329 (N_14329,N_13590,N_13485);
or U14330 (N_14330,N_13736,N_13593);
and U14331 (N_14331,N_13764,N_13307);
xor U14332 (N_14332,N_13804,N_13867);
nor U14333 (N_14333,N_13424,N_13900);
nor U14334 (N_14334,N_13091,N_13155);
and U14335 (N_14335,N_13746,N_13251);
xnor U14336 (N_14336,N_13024,N_13700);
xor U14337 (N_14337,N_13412,N_13858);
and U14338 (N_14338,N_13187,N_13898);
or U14339 (N_14339,N_13010,N_13286);
or U14340 (N_14340,N_13395,N_13711);
nor U14341 (N_14341,N_13281,N_13017);
or U14342 (N_14342,N_13798,N_13021);
and U14343 (N_14343,N_13110,N_13121);
nor U14344 (N_14344,N_13496,N_13890);
nor U14345 (N_14345,N_13328,N_13891);
and U14346 (N_14346,N_13398,N_13639);
and U14347 (N_14347,N_13591,N_13137);
nor U14348 (N_14348,N_13599,N_13548);
nand U14349 (N_14349,N_13596,N_13296);
nand U14350 (N_14350,N_13578,N_13194);
xnor U14351 (N_14351,N_13840,N_13457);
nand U14352 (N_14352,N_13594,N_13031);
nand U14353 (N_14353,N_13929,N_13499);
or U14354 (N_14354,N_13203,N_13456);
nand U14355 (N_14355,N_13147,N_13676);
xor U14356 (N_14356,N_13309,N_13897);
or U14357 (N_14357,N_13526,N_13149);
nor U14358 (N_14358,N_13996,N_13692);
and U14359 (N_14359,N_13540,N_13614);
xnor U14360 (N_14360,N_13844,N_13287);
nand U14361 (N_14361,N_13206,N_13018);
nor U14362 (N_14362,N_13737,N_13907);
or U14363 (N_14363,N_13875,N_13786);
and U14364 (N_14364,N_13930,N_13859);
and U14365 (N_14365,N_13256,N_13246);
nand U14366 (N_14366,N_13971,N_13562);
nand U14367 (N_14367,N_13799,N_13918);
or U14368 (N_14368,N_13111,N_13198);
nor U14369 (N_14369,N_13756,N_13409);
or U14370 (N_14370,N_13862,N_13625);
xor U14371 (N_14371,N_13458,N_13002);
nand U14372 (N_14372,N_13353,N_13235);
xor U14373 (N_14373,N_13785,N_13058);
nor U14374 (N_14374,N_13583,N_13841);
nand U14375 (N_14375,N_13410,N_13659);
xnor U14376 (N_14376,N_13414,N_13655);
nor U14377 (N_14377,N_13484,N_13038);
xor U14378 (N_14378,N_13942,N_13908);
and U14379 (N_14379,N_13448,N_13128);
xnor U14380 (N_14380,N_13042,N_13694);
nand U14381 (N_14381,N_13995,N_13949);
or U14382 (N_14382,N_13212,N_13902);
nand U14383 (N_14383,N_13505,N_13931);
xnor U14384 (N_14384,N_13234,N_13884);
xnor U14385 (N_14385,N_13623,N_13221);
and U14386 (N_14386,N_13359,N_13660);
and U14387 (N_14387,N_13179,N_13276);
nand U14388 (N_14388,N_13475,N_13830);
xnor U14389 (N_14389,N_13243,N_13832);
nand U14390 (N_14390,N_13551,N_13518);
and U14391 (N_14391,N_13089,N_13060);
and U14392 (N_14392,N_13103,N_13231);
nand U14393 (N_14393,N_13759,N_13539);
nand U14394 (N_14394,N_13420,N_13732);
nor U14395 (N_14395,N_13300,N_13143);
or U14396 (N_14396,N_13615,N_13403);
nor U14397 (N_14397,N_13582,N_13842);
xnor U14398 (N_14398,N_13846,N_13326);
nor U14399 (N_14399,N_13629,N_13182);
nand U14400 (N_14400,N_13837,N_13437);
xnor U14401 (N_14401,N_13960,N_13683);
nor U14402 (N_14402,N_13792,N_13054);
or U14403 (N_14403,N_13354,N_13431);
or U14404 (N_14404,N_13501,N_13318);
and U14405 (N_14405,N_13079,N_13775);
and U14406 (N_14406,N_13478,N_13522);
or U14407 (N_14407,N_13183,N_13780);
nor U14408 (N_14408,N_13446,N_13648);
nand U14409 (N_14409,N_13116,N_13250);
xor U14410 (N_14410,N_13912,N_13665);
nor U14411 (N_14411,N_13266,N_13298);
nor U14412 (N_14412,N_13560,N_13631);
nor U14413 (N_14413,N_13372,N_13517);
xor U14414 (N_14414,N_13416,N_13417);
or U14415 (N_14415,N_13109,N_13632);
nor U14416 (N_14416,N_13145,N_13379);
nor U14417 (N_14417,N_13207,N_13809);
nor U14418 (N_14418,N_13040,N_13443);
and U14419 (N_14419,N_13482,N_13401);
or U14420 (N_14420,N_13991,N_13968);
xor U14421 (N_14421,N_13544,N_13586);
nor U14422 (N_14422,N_13970,N_13990);
and U14423 (N_14423,N_13497,N_13973);
nor U14424 (N_14424,N_13160,N_13301);
nor U14425 (N_14425,N_13299,N_13404);
or U14426 (N_14426,N_13868,N_13576);
and U14427 (N_14427,N_13005,N_13325);
and U14428 (N_14428,N_13621,N_13911);
and U14429 (N_14429,N_13822,N_13514);
xnor U14430 (N_14430,N_13915,N_13752);
xor U14431 (N_14431,N_13873,N_13654);
xor U14432 (N_14432,N_13481,N_13559);
xor U14433 (N_14433,N_13172,N_13034);
or U14434 (N_14434,N_13674,N_13390);
nor U14435 (N_14435,N_13068,N_13422);
and U14436 (N_14436,N_13839,N_13349);
or U14437 (N_14437,N_13972,N_13753);
xor U14438 (N_14438,N_13225,N_13808);
or U14439 (N_14439,N_13758,N_13520);
or U14440 (N_14440,N_13527,N_13782);
or U14441 (N_14441,N_13641,N_13954);
nor U14442 (N_14442,N_13749,N_13291);
xnor U14443 (N_14443,N_13661,N_13267);
xor U14444 (N_14444,N_13713,N_13612);
and U14445 (N_14445,N_13715,N_13620);
xnor U14446 (N_14446,N_13001,N_13630);
or U14447 (N_14447,N_13059,N_13117);
and U14448 (N_14448,N_13075,N_13542);
nand U14449 (N_14449,N_13269,N_13776);
xnor U14450 (N_14450,N_13969,N_13791);
xor U14451 (N_14451,N_13153,N_13190);
xnor U14452 (N_14452,N_13209,N_13421);
and U14453 (N_14453,N_13580,N_13662);
nand U14454 (N_14454,N_13348,N_13205);
nand U14455 (N_14455,N_13565,N_13607);
nand U14456 (N_14456,N_13081,N_13254);
or U14457 (N_14457,N_13150,N_13065);
nand U14458 (N_14458,N_13925,N_13441);
nor U14459 (N_14459,N_13708,N_13125);
nor U14460 (N_14460,N_13317,N_13691);
xnor U14461 (N_14461,N_13280,N_13781);
or U14462 (N_14462,N_13803,N_13524);
or U14463 (N_14463,N_13521,N_13948);
nand U14464 (N_14464,N_13850,N_13500);
nand U14465 (N_14465,N_13029,N_13240);
nor U14466 (N_14466,N_13226,N_13041);
or U14467 (N_14467,N_13323,N_13735);
nor U14468 (N_14468,N_13957,N_13828);
or U14469 (N_14469,N_13989,N_13689);
nor U14470 (N_14470,N_13371,N_13763);
nor U14471 (N_14471,N_13387,N_13080);
nand U14472 (N_14472,N_13602,N_13479);
or U14473 (N_14473,N_13201,N_13000);
nor U14474 (N_14474,N_13537,N_13213);
or U14475 (N_14475,N_13730,N_13283);
and U14476 (N_14476,N_13725,N_13922);
nor U14477 (N_14477,N_13765,N_13530);
or U14478 (N_14478,N_13196,N_13988);
nand U14479 (N_14479,N_13057,N_13494);
nor U14480 (N_14480,N_13176,N_13098);
nor U14481 (N_14481,N_13690,N_13124);
or U14482 (N_14482,N_13236,N_13302);
nor U14483 (N_14483,N_13934,N_13817);
or U14484 (N_14484,N_13400,N_13750);
nor U14485 (N_14485,N_13777,N_13487);
or U14486 (N_14486,N_13491,N_13760);
nand U14487 (N_14487,N_13397,N_13761);
or U14488 (N_14488,N_13554,N_13144);
nand U14489 (N_14489,N_13156,N_13618);
and U14490 (N_14490,N_13023,N_13767);
and U14491 (N_14491,N_13938,N_13800);
and U14492 (N_14492,N_13561,N_13549);
nand U14493 (N_14493,N_13219,N_13056);
nand U14494 (N_14494,N_13067,N_13135);
and U14495 (N_14495,N_13263,N_13601);
or U14496 (N_14496,N_13104,N_13644);
nand U14497 (N_14497,N_13937,N_13308);
and U14498 (N_14498,N_13142,N_13106);
and U14499 (N_14499,N_13872,N_13418);
or U14500 (N_14500,N_13808,N_13376);
or U14501 (N_14501,N_13188,N_13482);
and U14502 (N_14502,N_13166,N_13862);
nand U14503 (N_14503,N_13838,N_13074);
nor U14504 (N_14504,N_13786,N_13069);
and U14505 (N_14505,N_13368,N_13766);
nor U14506 (N_14506,N_13050,N_13659);
and U14507 (N_14507,N_13104,N_13062);
and U14508 (N_14508,N_13077,N_13674);
nand U14509 (N_14509,N_13645,N_13401);
and U14510 (N_14510,N_13634,N_13740);
and U14511 (N_14511,N_13971,N_13484);
or U14512 (N_14512,N_13013,N_13218);
nor U14513 (N_14513,N_13924,N_13460);
nand U14514 (N_14514,N_13576,N_13814);
and U14515 (N_14515,N_13401,N_13648);
nand U14516 (N_14516,N_13518,N_13709);
or U14517 (N_14517,N_13788,N_13231);
xor U14518 (N_14518,N_13535,N_13334);
or U14519 (N_14519,N_13960,N_13010);
nor U14520 (N_14520,N_13951,N_13849);
nand U14521 (N_14521,N_13728,N_13299);
and U14522 (N_14522,N_13459,N_13571);
xor U14523 (N_14523,N_13585,N_13381);
nand U14524 (N_14524,N_13682,N_13608);
or U14525 (N_14525,N_13775,N_13512);
nor U14526 (N_14526,N_13640,N_13879);
nor U14527 (N_14527,N_13273,N_13134);
nand U14528 (N_14528,N_13041,N_13784);
or U14529 (N_14529,N_13246,N_13319);
and U14530 (N_14530,N_13265,N_13589);
nor U14531 (N_14531,N_13393,N_13925);
xnor U14532 (N_14532,N_13004,N_13386);
nor U14533 (N_14533,N_13207,N_13563);
nor U14534 (N_14534,N_13972,N_13604);
or U14535 (N_14535,N_13250,N_13063);
xor U14536 (N_14536,N_13556,N_13228);
and U14537 (N_14537,N_13019,N_13655);
or U14538 (N_14538,N_13051,N_13219);
nand U14539 (N_14539,N_13225,N_13216);
nand U14540 (N_14540,N_13263,N_13156);
nor U14541 (N_14541,N_13384,N_13829);
xnor U14542 (N_14542,N_13213,N_13430);
and U14543 (N_14543,N_13221,N_13580);
nor U14544 (N_14544,N_13952,N_13248);
nor U14545 (N_14545,N_13076,N_13242);
or U14546 (N_14546,N_13749,N_13691);
xnor U14547 (N_14547,N_13288,N_13259);
and U14548 (N_14548,N_13711,N_13773);
and U14549 (N_14549,N_13804,N_13081);
xor U14550 (N_14550,N_13091,N_13526);
xnor U14551 (N_14551,N_13778,N_13986);
and U14552 (N_14552,N_13310,N_13392);
or U14553 (N_14553,N_13554,N_13383);
or U14554 (N_14554,N_13821,N_13398);
or U14555 (N_14555,N_13427,N_13108);
and U14556 (N_14556,N_13781,N_13257);
nand U14557 (N_14557,N_13137,N_13842);
nor U14558 (N_14558,N_13973,N_13273);
and U14559 (N_14559,N_13708,N_13931);
xnor U14560 (N_14560,N_13895,N_13512);
or U14561 (N_14561,N_13883,N_13318);
nor U14562 (N_14562,N_13082,N_13617);
or U14563 (N_14563,N_13548,N_13224);
nor U14564 (N_14564,N_13936,N_13182);
nand U14565 (N_14565,N_13854,N_13804);
nand U14566 (N_14566,N_13478,N_13868);
xnor U14567 (N_14567,N_13230,N_13764);
nor U14568 (N_14568,N_13247,N_13114);
nand U14569 (N_14569,N_13260,N_13925);
and U14570 (N_14570,N_13556,N_13036);
nor U14571 (N_14571,N_13188,N_13533);
or U14572 (N_14572,N_13127,N_13280);
or U14573 (N_14573,N_13816,N_13098);
nand U14574 (N_14574,N_13574,N_13449);
nor U14575 (N_14575,N_13061,N_13572);
or U14576 (N_14576,N_13741,N_13179);
and U14577 (N_14577,N_13111,N_13222);
or U14578 (N_14578,N_13575,N_13238);
nand U14579 (N_14579,N_13104,N_13875);
nand U14580 (N_14580,N_13276,N_13889);
nor U14581 (N_14581,N_13752,N_13157);
xor U14582 (N_14582,N_13332,N_13073);
nor U14583 (N_14583,N_13640,N_13463);
nand U14584 (N_14584,N_13729,N_13748);
and U14585 (N_14585,N_13668,N_13055);
and U14586 (N_14586,N_13768,N_13561);
and U14587 (N_14587,N_13768,N_13365);
nand U14588 (N_14588,N_13548,N_13140);
xnor U14589 (N_14589,N_13012,N_13129);
nor U14590 (N_14590,N_13811,N_13345);
xnor U14591 (N_14591,N_13509,N_13676);
or U14592 (N_14592,N_13531,N_13219);
and U14593 (N_14593,N_13338,N_13621);
and U14594 (N_14594,N_13250,N_13977);
or U14595 (N_14595,N_13565,N_13156);
nand U14596 (N_14596,N_13667,N_13736);
nor U14597 (N_14597,N_13727,N_13158);
xor U14598 (N_14598,N_13810,N_13924);
and U14599 (N_14599,N_13615,N_13159);
nor U14600 (N_14600,N_13705,N_13107);
or U14601 (N_14601,N_13901,N_13296);
and U14602 (N_14602,N_13593,N_13958);
nor U14603 (N_14603,N_13207,N_13744);
nor U14604 (N_14604,N_13419,N_13641);
and U14605 (N_14605,N_13336,N_13253);
or U14606 (N_14606,N_13732,N_13637);
xor U14607 (N_14607,N_13058,N_13338);
nor U14608 (N_14608,N_13561,N_13066);
and U14609 (N_14609,N_13392,N_13124);
nor U14610 (N_14610,N_13025,N_13201);
xnor U14611 (N_14611,N_13018,N_13732);
and U14612 (N_14612,N_13139,N_13539);
xnor U14613 (N_14613,N_13224,N_13327);
or U14614 (N_14614,N_13556,N_13754);
nand U14615 (N_14615,N_13225,N_13499);
nand U14616 (N_14616,N_13345,N_13348);
and U14617 (N_14617,N_13718,N_13941);
or U14618 (N_14618,N_13961,N_13313);
and U14619 (N_14619,N_13750,N_13456);
nor U14620 (N_14620,N_13744,N_13124);
nand U14621 (N_14621,N_13059,N_13326);
nor U14622 (N_14622,N_13190,N_13270);
and U14623 (N_14623,N_13713,N_13567);
nand U14624 (N_14624,N_13770,N_13108);
nor U14625 (N_14625,N_13658,N_13996);
nor U14626 (N_14626,N_13040,N_13557);
or U14627 (N_14627,N_13493,N_13096);
nand U14628 (N_14628,N_13909,N_13133);
nor U14629 (N_14629,N_13648,N_13804);
xnor U14630 (N_14630,N_13293,N_13260);
nand U14631 (N_14631,N_13955,N_13208);
or U14632 (N_14632,N_13439,N_13423);
nor U14633 (N_14633,N_13392,N_13383);
nor U14634 (N_14634,N_13141,N_13829);
xor U14635 (N_14635,N_13528,N_13184);
and U14636 (N_14636,N_13707,N_13958);
and U14637 (N_14637,N_13579,N_13489);
and U14638 (N_14638,N_13218,N_13116);
nor U14639 (N_14639,N_13622,N_13456);
xnor U14640 (N_14640,N_13399,N_13078);
or U14641 (N_14641,N_13724,N_13613);
xnor U14642 (N_14642,N_13831,N_13005);
nor U14643 (N_14643,N_13465,N_13874);
or U14644 (N_14644,N_13608,N_13474);
xnor U14645 (N_14645,N_13348,N_13023);
nand U14646 (N_14646,N_13511,N_13815);
nor U14647 (N_14647,N_13849,N_13997);
nand U14648 (N_14648,N_13981,N_13900);
nor U14649 (N_14649,N_13098,N_13010);
and U14650 (N_14650,N_13389,N_13073);
and U14651 (N_14651,N_13705,N_13696);
nor U14652 (N_14652,N_13350,N_13558);
nand U14653 (N_14653,N_13798,N_13858);
and U14654 (N_14654,N_13202,N_13988);
or U14655 (N_14655,N_13778,N_13059);
or U14656 (N_14656,N_13957,N_13430);
and U14657 (N_14657,N_13591,N_13348);
and U14658 (N_14658,N_13431,N_13525);
nand U14659 (N_14659,N_13040,N_13087);
nor U14660 (N_14660,N_13543,N_13759);
or U14661 (N_14661,N_13597,N_13924);
or U14662 (N_14662,N_13107,N_13812);
xor U14663 (N_14663,N_13801,N_13315);
nor U14664 (N_14664,N_13642,N_13500);
nand U14665 (N_14665,N_13006,N_13386);
nor U14666 (N_14666,N_13254,N_13691);
or U14667 (N_14667,N_13336,N_13525);
xnor U14668 (N_14668,N_13773,N_13107);
nand U14669 (N_14669,N_13060,N_13923);
nor U14670 (N_14670,N_13009,N_13160);
and U14671 (N_14671,N_13700,N_13990);
xor U14672 (N_14672,N_13611,N_13233);
or U14673 (N_14673,N_13171,N_13119);
xnor U14674 (N_14674,N_13194,N_13919);
nor U14675 (N_14675,N_13625,N_13195);
nand U14676 (N_14676,N_13099,N_13861);
nand U14677 (N_14677,N_13187,N_13066);
nand U14678 (N_14678,N_13083,N_13031);
xor U14679 (N_14679,N_13490,N_13917);
and U14680 (N_14680,N_13285,N_13144);
nand U14681 (N_14681,N_13539,N_13800);
xnor U14682 (N_14682,N_13746,N_13210);
nor U14683 (N_14683,N_13069,N_13964);
nand U14684 (N_14684,N_13614,N_13015);
nand U14685 (N_14685,N_13071,N_13669);
and U14686 (N_14686,N_13038,N_13066);
xor U14687 (N_14687,N_13743,N_13268);
nand U14688 (N_14688,N_13544,N_13451);
nand U14689 (N_14689,N_13956,N_13369);
or U14690 (N_14690,N_13054,N_13134);
nand U14691 (N_14691,N_13961,N_13129);
xor U14692 (N_14692,N_13147,N_13253);
or U14693 (N_14693,N_13171,N_13360);
nor U14694 (N_14694,N_13517,N_13812);
and U14695 (N_14695,N_13737,N_13400);
nor U14696 (N_14696,N_13229,N_13744);
or U14697 (N_14697,N_13045,N_13967);
nor U14698 (N_14698,N_13544,N_13766);
xnor U14699 (N_14699,N_13787,N_13196);
nor U14700 (N_14700,N_13482,N_13408);
xnor U14701 (N_14701,N_13909,N_13980);
xor U14702 (N_14702,N_13276,N_13158);
nor U14703 (N_14703,N_13721,N_13125);
and U14704 (N_14704,N_13551,N_13186);
nor U14705 (N_14705,N_13129,N_13030);
and U14706 (N_14706,N_13148,N_13092);
xor U14707 (N_14707,N_13640,N_13053);
xor U14708 (N_14708,N_13472,N_13933);
nand U14709 (N_14709,N_13266,N_13959);
nor U14710 (N_14710,N_13571,N_13606);
xor U14711 (N_14711,N_13909,N_13507);
and U14712 (N_14712,N_13021,N_13684);
xnor U14713 (N_14713,N_13684,N_13468);
xnor U14714 (N_14714,N_13858,N_13906);
nand U14715 (N_14715,N_13315,N_13277);
or U14716 (N_14716,N_13072,N_13414);
nor U14717 (N_14717,N_13822,N_13195);
nand U14718 (N_14718,N_13422,N_13423);
or U14719 (N_14719,N_13965,N_13548);
nor U14720 (N_14720,N_13118,N_13784);
or U14721 (N_14721,N_13870,N_13807);
or U14722 (N_14722,N_13901,N_13645);
nand U14723 (N_14723,N_13619,N_13687);
nor U14724 (N_14724,N_13456,N_13058);
or U14725 (N_14725,N_13017,N_13597);
and U14726 (N_14726,N_13136,N_13228);
nand U14727 (N_14727,N_13041,N_13484);
nand U14728 (N_14728,N_13834,N_13179);
and U14729 (N_14729,N_13768,N_13096);
nand U14730 (N_14730,N_13886,N_13131);
and U14731 (N_14731,N_13223,N_13512);
and U14732 (N_14732,N_13302,N_13411);
and U14733 (N_14733,N_13550,N_13143);
nand U14734 (N_14734,N_13910,N_13840);
nand U14735 (N_14735,N_13930,N_13815);
or U14736 (N_14736,N_13125,N_13439);
xnor U14737 (N_14737,N_13971,N_13708);
and U14738 (N_14738,N_13886,N_13991);
nor U14739 (N_14739,N_13189,N_13526);
nand U14740 (N_14740,N_13325,N_13392);
nor U14741 (N_14741,N_13573,N_13713);
nor U14742 (N_14742,N_13393,N_13684);
xor U14743 (N_14743,N_13550,N_13819);
and U14744 (N_14744,N_13606,N_13082);
xor U14745 (N_14745,N_13906,N_13820);
and U14746 (N_14746,N_13896,N_13582);
and U14747 (N_14747,N_13240,N_13641);
and U14748 (N_14748,N_13543,N_13335);
nor U14749 (N_14749,N_13479,N_13318);
nor U14750 (N_14750,N_13834,N_13255);
and U14751 (N_14751,N_13678,N_13522);
or U14752 (N_14752,N_13446,N_13356);
and U14753 (N_14753,N_13518,N_13968);
xnor U14754 (N_14754,N_13916,N_13313);
nor U14755 (N_14755,N_13089,N_13915);
or U14756 (N_14756,N_13584,N_13897);
nor U14757 (N_14757,N_13773,N_13366);
or U14758 (N_14758,N_13549,N_13138);
or U14759 (N_14759,N_13178,N_13813);
nor U14760 (N_14760,N_13281,N_13922);
nand U14761 (N_14761,N_13206,N_13266);
nor U14762 (N_14762,N_13442,N_13292);
and U14763 (N_14763,N_13161,N_13289);
nor U14764 (N_14764,N_13202,N_13476);
xor U14765 (N_14765,N_13707,N_13253);
xor U14766 (N_14766,N_13321,N_13859);
or U14767 (N_14767,N_13241,N_13835);
and U14768 (N_14768,N_13348,N_13673);
or U14769 (N_14769,N_13410,N_13390);
or U14770 (N_14770,N_13763,N_13656);
xor U14771 (N_14771,N_13183,N_13759);
nor U14772 (N_14772,N_13700,N_13731);
and U14773 (N_14773,N_13022,N_13165);
nor U14774 (N_14774,N_13952,N_13098);
or U14775 (N_14775,N_13451,N_13431);
or U14776 (N_14776,N_13374,N_13149);
xnor U14777 (N_14777,N_13556,N_13971);
nor U14778 (N_14778,N_13370,N_13935);
and U14779 (N_14779,N_13231,N_13095);
nand U14780 (N_14780,N_13919,N_13285);
nand U14781 (N_14781,N_13484,N_13170);
or U14782 (N_14782,N_13484,N_13193);
nand U14783 (N_14783,N_13194,N_13473);
nor U14784 (N_14784,N_13482,N_13034);
nor U14785 (N_14785,N_13210,N_13101);
or U14786 (N_14786,N_13210,N_13274);
nor U14787 (N_14787,N_13340,N_13085);
nor U14788 (N_14788,N_13002,N_13862);
xor U14789 (N_14789,N_13850,N_13497);
or U14790 (N_14790,N_13837,N_13247);
nand U14791 (N_14791,N_13646,N_13262);
and U14792 (N_14792,N_13540,N_13002);
nand U14793 (N_14793,N_13791,N_13039);
and U14794 (N_14794,N_13175,N_13583);
xnor U14795 (N_14795,N_13333,N_13441);
and U14796 (N_14796,N_13403,N_13253);
and U14797 (N_14797,N_13989,N_13834);
xor U14798 (N_14798,N_13040,N_13705);
or U14799 (N_14799,N_13469,N_13665);
nand U14800 (N_14800,N_13358,N_13908);
nand U14801 (N_14801,N_13199,N_13839);
nand U14802 (N_14802,N_13429,N_13848);
nand U14803 (N_14803,N_13022,N_13511);
nand U14804 (N_14804,N_13264,N_13064);
nand U14805 (N_14805,N_13887,N_13982);
and U14806 (N_14806,N_13918,N_13192);
xnor U14807 (N_14807,N_13289,N_13298);
and U14808 (N_14808,N_13428,N_13283);
or U14809 (N_14809,N_13001,N_13971);
xnor U14810 (N_14810,N_13783,N_13206);
xnor U14811 (N_14811,N_13462,N_13435);
or U14812 (N_14812,N_13559,N_13777);
or U14813 (N_14813,N_13125,N_13194);
nand U14814 (N_14814,N_13136,N_13088);
nor U14815 (N_14815,N_13922,N_13129);
or U14816 (N_14816,N_13047,N_13837);
nor U14817 (N_14817,N_13498,N_13945);
or U14818 (N_14818,N_13936,N_13232);
nand U14819 (N_14819,N_13391,N_13137);
nor U14820 (N_14820,N_13115,N_13054);
and U14821 (N_14821,N_13674,N_13591);
and U14822 (N_14822,N_13813,N_13310);
nand U14823 (N_14823,N_13084,N_13217);
and U14824 (N_14824,N_13848,N_13431);
nor U14825 (N_14825,N_13704,N_13589);
or U14826 (N_14826,N_13897,N_13962);
nor U14827 (N_14827,N_13926,N_13498);
or U14828 (N_14828,N_13538,N_13104);
nor U14829 (N_14829,N_13639,N_13694);
or U14830 (N_14830,N_13842,N_13341);
nor U14831 (N_14831,N_13426,N_13955);
and U14832 (N_14832,N_13617,N_13827);
or U14833 (N_14833,N_13192,N_13177);
or U14834 (N_14834,N_13789,N_13170);
xor U14835 (N_14835,N_13542,N_13937);
or U14836 (N_14836,N_13525,N_13919);
nor U14837 (N_14837,N_13884,N_13766);
xnor U14838 (N_14838,N_13213,N_13814);
or U14839 (N_14839,N_13877,N_13144);
nor U14840 (N_14840,N_13065,N_13736);
nand U14841 (N_14841,N_13705,N_13265);
xnor U14842 (N_14842,N_13952,N_13846);
or U14843 (N_14843,N_13737,N_13833);
xnor U14844 (N_14844,N_13117,N_13123);
nand U14845 (N_14845,N_13718,N_13518);
nor U14846 (N_14846,N_13833,N_13217);
xnor U14847 (N_14847,N_13855,N_13360);
nand U14848 (N_14848,N_13702,N_13736);
or U14849 (N_14849,N_13180,N_13001);
nor U14850 (N_14850,N_13528,N_13263);
or U14851 (N_14851,N_13457,N_13712);
nor U14852 (N_14852,N_13302,N_13201);
xor U14853 (N_14853,N_13736,N_13821);
nand U14854 (N_14854,N_13991,N_13327);
xnor U14855 (N_14855,N_13846,N_13453);
and U14856 (N_14856,N_13205,N_13551);
nand U14857 (N_14857,N_13400,N_13827);
nor U14858 (N_14858,N_13734,N_13097);
and U14859 (N_14859,N_13459,N_13517);
nor U14860 (N_14860,N_13863,N_13310);
xor U14861 (N_14861,N_13698,N_13992);
and U14862 (N_14862,N_13266,N_13826);
nor U14863 (N_14863,N_13055,N_13190);
xnor U14864 (N_14864,N_13240,N_13314);
nand U14865 (N_14865,N_13464,N_13756);
nor U14866 (N_14866,N_13316,N_13229);
nor U14867 (N_14867,N_13340,N_13909);
and U14868 (N_14868,N_13407,N_13459);
nand U14869 (N_14869,N_13105,N_13632);
xnor U14870 (N_14870,N_13181,N_13419);
and U14871 (N_14871,N_13265,N_13471);
nand U14872 (N_14872,N_13358,N_13077);
or U14873 (N_14873,N_13448,N_13056);
xnor U14874 (N_14874,N_13294,N_13262);
and U14875 (N_14875,N_13287,N_13086);
or U14876 (N_14876,N_13244,N_13417);
or U14877 (N_14877,N_13148,N_13914);
nor U14878 (N_14878,N_13725,N_13687);
nand U14879 (N_14879,N_13996,N_13827);
nand U14880 (N_14880,N_13772,N_13985);
or U14881 (N_14881,N_13823,N_13143);
and U14882 (N_14882,N_13438,N_13275);
and U14883 (N_14883,N_13345,N_13691);
and U14884 (N_14884,N_13984,N_13646);
xnor U14885 (N_14885,N_13871,N_13169);
xor U14886 (N_14886,N_13507,N_13373);
or U14887 (N_14887,N_13457,N_13290);
nand U14888 (N_14888,N_13203,N_13360);
nor U14889 (N_14889,N_13215,N_13625);
or U14890 (N_14890,N_13301,N_13196);
and U14891 (N_14891,N_13193,N_13874);
nor U14892 (N_14892,N_13074,N_13357);
and U14893 (N_14893,N_13146,N_13996);
xnor U14894 (N_14894,N_13266,N_13488);
and U14895 (N_14895,N_13228,N_13734);
nand U14896 (N_14896,N_13332,N_13001);
xnor U14897 (N_14897,N_13556,N_13309);
xor U14898 (N_14898,N_13835,N_13822);
xnor U14899 (N_14899,N_13191,N_13410);
xnor U14900 (N_14900,N_13027,N_13867);
or U14901 (N_14901,N_13134,N_13628);
and U14902 (N_14902,N_13392,N_13692);
and U14903 (N_14903,N_13213,N_13143);
nand U14904 (N_14904,N_13292,N_13037);
nand U14905 (N_14905,N_13330,N_13714);
nand U14906 (N_14906,N_13996,N_13634);
nor U14907 (N_14907,N_13789,N_13640);
nor U14908 (N_14908,N_13867,N_13514);
nand U14909 (N_14909,N_13786,N_13086);
or U14910 (N_14910,N_13287,N_13146);
xnor U14911 (N_14911,N_13774,N_13572);
xnor U14912 (N_14912,N_13543,N_13887);
xor U14913 (N_14913,N_13118,N_13787);
nor U14914 (N_14914,N_13678,N_13108);
nor U14915 (N_14915,N_13947,N_13565);
and U14916 (N_14916,N_13816,N_13850);
and U14917 (N_14917,N_13072,N_13608);
nor U14918 (N_14918,N_13878,N_13362);
nand U14919 (N_14919,N_13285,N_13728);
xor U14920 (N_14920,N_13173,N_13526);
nor U14921 (N_14921,N_13799,N_13084);
or U14922 (N_14922,N_13652,N_13892);
or U14923 (N_14923,N_13944,N_13752);
nand U14924 (N_14924,N_13049,N_13082);
or U14925 (N_14925,N_13315,N_13518);
and U14926 (N_14926,N_13054,N_13800);
xnor U14927 (N_14927,N_13034,N_13373);
or U14928 (N_14928,N_13715,N_13907);
xor U14929 (N_14929,N_13169,N_13992);
nor U14930 (N_14930,N_13789,N_13243);
and U14931 (N_14931,N_13827,N_13148);
nor U14932 (N_14932,N_13425,N_13671);
nand U14933 (N_14933,N_13388,N_13941);
nor U14934 (N_14934,N_13988,N_13645);
nor U14935 (N_14935,N_13614,N_13891);
nand U14936 (N_14936,N_13747,N_13542);
nand U14937 (N_14937,N_13366,N_13353);
or U14938 (N_14938,N_13759,N_13730);
xor U14939 (N_14939,N_13073,N_13052);
xnor U14940 (N_14940,N_13239,N_13780);
nor U14941 (N_14941,N_13945,N_13074);
xor U14942 (N_14942,N_13198,N_13969);
and U14943 (N_14943,N_13330,N_13377);
or U14944 (N_14944,N_13589,N_13973);
or U14945 (N_14945,N_13572,N_13662);
and U14946 (N_14946,N_13903,N_13591);
nor U14947 (N_14947,N_13249,N_13768);
xnor U14948 (N_14948,N_13963,N_13705);
or U14949 (N_14949,N_13236,N_13422);
and U14950 (N_14950,N_13359,N_13402);
xnor U14951 (N_14951,N_13835,N_13094);
or U14952 (N_14952,N_13779,N_13246);
xor U14953 (N_14953,N_13388,N_13002);
and U14954 (N_14954,N_13960,N_13638);
and U14955 (N_14955,N_13240,N_13977);
or U14956 (N_14956,N_13542,N_13431);
and U14957 (N_14957,N_13268,N_13823);
or U14958 (N_14958,N_13585,N_13700);
or U14959 (N_14959,N_13525,N_13144);
and U14960 (N_14960,N_13113,N_13063);
xnor U14961 (N_14961,N_13159,N_13778);
and U14962 (N_14962,N_13145,N_13692);
xor U14963 (N_14963,N_13209,N_13082);
nand U14964 (N_14964,N_13948,N_13251);
nor U14965 (N_14965,N_13623,N_13220);
and U14966 (N_14966,N_13687,N_13005);
and U14967 (N_14967,N_13578,N_13949);
or U14968 (N_14968,N_13318,N_13406);
or U14969 (N_14969,N_13272,N_13235);
or U14970 (N_14970,N_13579,N_13212);
nor U14971 (N_14971,N_13923,N_13473);
xnor U14972 (N_14972,N_13396,N_13545);
xnor U14973 (N_14973,N_13810,N_13778);
and U14974 (N_14974,N_13120,N_13096);
and U14975 (N_14975,N_13452,N_13899);
nand U14976 (N_14976,N_13187,N_13389);
nand U14977 (N_14977,N_13784,N_13368);
xor U14978 (N_14978,N_13647,N_13592);
nand U14979 (N_14979,N_13254,N_13377);
nand U14980 (N_14980,N_13008,N_13995);
and U14981 (N_14981,N_13219,N_13738);
or U14982 (N_14982,N_13921,N_13277);
or U14983 (N_14983,N_13599,N_13363);
xnor U14984 (N_14984,N_13578,N_13279);
nand U14985 (N_14985,N_13776,N_13573);
nor U14986 (N_14986,N_13619,N_13585);
xor U14987 (N_14987,N_13273,N_13574);
xnor U14988 (N_14988,N_13872,N_13569);
and U14989 (N_14989,N_13867,N_13352);
or U14990 (N_14990,N_13870,N_13552);
nand U14991 (N_14991,N_13027,N_13904);
and U14992 (N_14992,N_13743,N_13361);
nand U14993 (N_14993,N_13391,N_13617);
nand U14994 (N_14994,N_13368,N_13228);
or U14995 (N_14995,N_13889,N_13605);
xor U14996 (N_14996,N_13897,N_13396);
or U14997 (N_14997,N_13833,N_13520);
nor U14998 (N_14998,N_13246,N_13928);
or U14999 (N_14999,N_13476,N_13307);
or U15000 (N_15000,N_14981,N_14423);
nor U15001 (N_15001,N_14693,N_14625);
and U15002 (N_15002,N_14692,N_14300);
nor U15003 (N_15003,N_14001,N_14074);
xnor U15004 (N_15004,N_14867,N_14105);
and U15005 (N_15005,N_14909,N_14958);
or U15006 (N_15006,N_14233,N_14882);
nor U15007 (N_15007,N_14401,N_14457);
and U15008 (N_15008,N_14435,N_14740);
and U15009 (N_15009,N_14648,N_14148);
nor U15010 (N_15010,N_14192,N_14470);
xnor U15011 (N_15011,N_14309,N_14136);
nor U15012 (N_15012,N_14903,N_14044);
nand U15013 (N_15013,N_14913,N_14473);
nand U15014 (N_15014,N_14095,N_14091);
nand U15015 (N_15015,N_14033,N_14516);
nand U15016 (N_15016,N_14606,N_14107);
and U15017 (N_15017,N_14014,N_14721);
xor U15018 (N_15018,N_14902,N_14504);
and U15019 (N_15019,N_14809,N_14102);
nor U15020 (N_15020,N_14156,N_14904);
nor U15021 (N_15021,N_14539,N_14489);
xor U15022 (N_15022,N_14260,N_14694);
and U15023 (N_15023,N_14326,N_14803);
nor U15024 (N_15024,N_14346,N_14293);
and U15025 (N_15025,N_14143,N_14840);
nor U15026 (N_15026,N_14733,N_14822);
or U15027 (N_15027,N_14094,N_14264);
and U15028 (N_15028,N_14591,N_14350);
nand U15029 (N_15029,N_14535,N_14086);
nand U15030 (N_15030,N_14492,N_14420);
and U15031 (N_15031,N_14615,N_14607);
xnor U15032 (N_15032,N_14180,N_14240);
nand U15033 (N_15033,N_14170,N_14378);
nand U15034 (N_15034,N_14668,N_14275);
xor U15035 (N_15035,N_14667,N_14491);
or U15036 (N_15036,N_14093,N_14732);
and U15037 (N_15037,N_14449,N_14421);
or U15038 (N_15038,N_14334,N_14816);
or U15039 (N_15039,N_14511,N_14187);
and U15040 (N_15040,N_14938,N_14076);
nor U15041 (N_15041,N_14598,N_14638);
or U15042 (N_15042,N_14532,N_14720);
xor U15043 (N_15043,N_14222,N_14796);
or U15044 (N_15044,N_14277,N_14128);
nand U15045 (N_15045,N_14994,N_14020);
nor U15046 (N_15046,N_14345,N_14905);
or U15047 (N_15047,N_14000,N_14654);
xor U15048 (N_15048,N_14567,N_14211);
or U15049 (N_15049,N_14786,N_14769);
nand U15050 (N_15050,N_14603,N_14292);
nand U15051 (N_15051,N_14734,N_14032);
or U15052 (N_15052,N_14442,N_14447);
xnor U15053 (N_15053,N_14568,N_14430);
or U15054 (N_15054,N_14810,N_14026);
nor U15055 (N_15055,N_14730,N_14077);
and U15056 (N_15056,N_14827,N_14058);
and U15057 (N_15057,N_14040,N_14670);
nand U15058 (N_15058,N_14820,N_14963);
and U15059 (N_15059,N_14198,N_14324);
or U15060 (N_15060,N_14529,N_14487);
and U15061 (N_15061,N_14967,N_14787);
and U15062 (N_15062,N_14616,N_14499);
xor U15063 (N_15063,N_14906,N_14917);
nor U15064 (N_15064,N_14150,N_14363);
nor U15065 (N_15065,N_14267,N_14377);
and U15066 (N_15066,N_14851,N_14579);
or U15067 (N_15067,N_14046,N_14676);
and U15068 (N_15068,N_14137,N_14593);
and U15069 (N_15069,N_14776,N_14565);
xnor U15070 (N_15070,N_14066,N_14551);
xor U15071 (N_15071,N_14812,N_14237);
nand U15072 (N_15072,N_14775,N_14836);
nor U15073 (N_15073,N_14555,N_14817);
nand U15074 (N_15074,N_14548,N_14484);
nor U15075 (N_15075,N_14242,N_14847);
xnor U15076 (N_15076,N_14117,N_14488);
or U15077 (N_15077,N_14444,N_14992);
nand U15078 (N_15078,N_14856,N_14357);
nor U15079 (N_15079,N_14258,N_14877);
nand U15080 (N_15080,N_14830,N_14496);
nand U15081 (N_15081,N_14713,N_14084);
nand U15082 (N_15082,N_14316,N_14842);
and U15083 (N_15083,N_14062,N_14764);
xor U15084 (N_15084,N_14053,N_14605);
or U15085 (N_15085,N_14415,N_14898);
or U15086 (N_15086,N_14518,N_14110);
nand U15087 (N_15087,N_14250,N_14849);
xor U15088 (N_15088,N_14151,N_14104);
nand U15089 (N_15089,N_14212,N_14149);
xnor U15090 (N_15090,N_14653,N_14660);
nor U15091 (N_15091,N_14715,N_14742);
and U15092 (N_15092,N_14722,N_14129);
xnor U15093 (N_15093,N_14572,N_14343);
xnor U15094 (N_15094,N_14699,N_14171);
nand U15095 (N_15095,N_14411,N_14587);
nand U15096 (N_15096,N_14295,N_14498);
or U15097 (N_15097,N_14834,N_14090);
xor U15098 (N_15098,N_14096,N_14333);
and U15099 (N_15099,N_14768,N_14626);
nor U15100 (N_15100,N_14883,N_14220);
xnor U15101 (N_15101,N_14658,N_14079);
or U15102 (N_15102,N_14244,N_14520);
nand U15103 (N_15103,N_14749,N_14179);
or U15104 (N_15104,N_14761,N_14805);
or U15105 (N_15105,N_14235,N_14880);
or U15106 (N_15106,N_14055,N_14627);
and U15107 (N_15107,N_14164,N_14544);
or U15108 (N_15108,N_14203,N_14331);
and U15109 (N_15109,N_14045,N_14861);
or U15110 (N_15110,N_14866,N_14098);
xnor U15111 (N_15111,N_14312,N_14416);
and U15112 (N_15112,N_14841,N_14405);
nand U15113 (N_15113,N_14330,N_14344);
nand U15114 (N_15114,N_14513,N_14092);
nor U15115 (N_15115,N_14410,N_14234);
nand U15116 (N_15116,N_14177,N_14213);
or U15117 (N_15117,N_14017,N_14640);
and U15118 (N_15118,N_14811,N_14596);
and U15119 (N_15119,N_14945,N_14819);
and U15120 (N_15120,N_14747,N_14426);
xor U15121 (N_15121,N_14123,N_14563);
and U15122 (N_15122,N_14298,N_14229);
or U15123 (N_15123,N_14621,N_14783);
and U15124 (N_15124,N_14160,N_14048);
xor U15125 (N_15125,N_14631,N_14007);
xnor U15126 (N_15126,N_14808,N_14208);
xnor U15127 (N_15127,N_14673,N_14885);
or U15128 (N_15128,N_14113,N_14131);
and U15129 (N_15129,N_14610,N_14839);
or U15130 (N_15130,N_14698,N_14986);
or U15131 (N_15131,N_14506,N_14288);
nor U15132 (N_15132,N_14801,N_14075);
and U15133 (N_15133,N_14038,N_14678);
xnor U15134 (N_15134,N_14845,N_14463);
nand U15135 (N_15135,N_14940,N_14894);
xor U15136 (N_15136,N_14448,N_14739);
nor U15137 (N_15137,N_14680,N_14282);
nor U15138 (N_15138,N_14521,N_14388);
xor U15139 (N_15139,N_14818,N_14085);
or U15140 (N_15140,N_14697,N_14569);
nor U15141 (N_15141,N_14995,N_14087);
nor U15142 (N_15142,N_14051,N_14710);
xnor U15143 (N_15143,N_14735,N_14329);
nand U15144 (N_15144,N_14942,N_14462);
nand U15145 (N_15145,N_14303,N_14646);
nand U15146 (N_15146,N_14273,N_14534);
xnor U15147 (N_15147,N_14554,N_14467);
xnor U15148 (N_15148,N_14056,N_14297);
or U15149 (N_15149,N_14174,N_14952);
nand U15150 (N_15150,N_14912,N_14528);
nand U15151 (N_15151,N_14481,N_14083);
xnor U15152 (N_15152,N_14666,N_14469);
nor U15153 (N_15153,N_14404,N_14766);
and U15154 (N_15154,N_14159,N_14474);
or U15155 (N_15155,N_14990,N_14527);
nand U15156 (N_15156,N_14974,N_14407);
nand U15157 (N_15157,N_14009,N_14620);
nor U15158 (N_15158,N_14550,N_14750);
nor U15159 (N_15159,N_14061,N_14858);
xor U15160 (N_15160,N_14276,N_14207);
nand U15161 (N_15161,N_14310,N_14552);
nor U15162 (N_15162,N_14980,N_14672);
nor U15163 (N_15163,N_14006,N_14386);
nor U15164 (N_15164,N_14547,N_14635);
and U15165 (N_15165,N_14854,N_14762);
nand U15166 (N_15166,N_14478,N_14623);
nor U15167 (N_15167,N_14389,N_14439);
and U15168 (N_15168,N_14935,N_14614);
xnor U15169 (N_15169,N_14997,N_14328);
xor U15170 (N_15170,N_14073,N_14140);
nand U15171 (N_15171,N_14919,N_14976);
nand U15172 (N_15172,N_14645,N_14723);
nand U15173 (N_15173,N_14023,N_14533);
and U15174 (N_15174,N_14600,N_14925);
and U15175 (N_15175,N_14526,N_14376);
or U15176 (N_15176,N_14384,N_14115);
nand U15177 (N_15177,N_14018,N_14857);
nand U15178 (N_15178,N_14443,N_14753);
nand U15179 (N_15179,N_14375,N_14785);
nor U15180 (N_15180,N_14332,N_14826);
nor U15181 (N_15181,N_14949,N_14209);
or U15182 (N_15182,N_14057,N_14978);
and U15183 (N_15183,N_14262,N_14950);
nand U15184 (N_15184,N_14153,N_14173);
or U15185 (N_15185,N_14690,N_14434);
xnor U15186 (N_15186,N_14438,N_14178);
and U15187 (N_15187,N_14687,N_14688);
xnor U15188 (N_15188,N_14936,N_14396);
and U15189 (N_15189,N_14991,N_14167);
nand U15190 (N_15190,N_14285,N_14706);
or U15191 (N_15191,N_14947,N_14500);
xor U15192 (N_15192,N_14025,N_14597);
nor U15193 (N_15193,N_14479,N_14705);
and U15194 (N_15194,N_14590,N_14127);
xnor U15195 (N_15195,N_14955,N_14099);
or U15196 (N_15196,N_14249,N_14800);
nor U15197 (N_15197,N_14542,N_14944);
xnor U15198 (N_15198,N_14793,N_14712);
xor U15199 (N_15199,N_14147,N_14274);
or U15200 (N_15200,N_14510,N_14899);
nor U15201 (N_15201,N_14726,N_14582);
nor U15202 (N_15202,N_14281,N_14195);
nor U15203 (N_15203,N_14973,N_14746);
nand U15204 (N_15204,N_14251,N_14729);
nand U15205 (N_15205,N_14838,N_14985);
or U15206 (N_15206,N_14193,N_14910);
nand U15207 (N_15207,N_14709,N_14964);
or U15208 (N_15208,N_14379,N_14825);
xnor U15209 (N_15209,N_14215,N_14414);
xnor U15210 (N_15210,N_14185,N_14155);
and U15211 (N_15211,N_14770,N_14558);
and U15212 (N_15212,N_14794,N_14029);
or U15213 (N_15213,N_14814,N_14427);
xor U15214 (N_15214,N_14372,N_14031);
xor U15215 (N_15215,N_14662,N_14078);
and U15216 (N_15216,N_14369,N_14966);
nand U15217 (N_15217,N_14704,N_14194);
nand U15218 (N_15218,N_14863,N_14340);
and U15219 (N_15219,N_14731,N_14509);
or U15220 (N_15220,N_14915,N_14987);
nand U15221 (N_15221,N_14920,N_14860);
nor U15222 (N_15222,N_14373,N_14684);
or U15223 (N_15223,N_14921,N_14719);
nor U15224 (N_15224,N_14097,N_14381);
xor U15225 (N_15225,N_14517,N_14119);
xnor U15226 (N_15226,N_14538,N_14868);
and U15227 (N_15227,N_14755,N_14617);
xor U15228 (N_15228,N_14308,N_14772);
xnor U15229 (N_15229,N_14395,N_14422);
or U15230 (N_15230,N_14887,N_14953);
nand U15231 (N_15231,N_14320,N_14541);
or U15232 (N_15232,N_14613,N_14199);
and U15233 (N_15233,N_14961,N_14546);
nand U15234 (N_15234,N_14279,N_14677);
and U15235 (N_15235,N_14190,N_14774);
nand U15236 (N_15236,N_14465,N_14937);
nor U15237 (N_15237,N_14881,N_14486);
and U15238 (N_15238,N_14429,N_14412);
or U15239 (N_15239,N_14652,N_14134);
xor U15240 (N_15240,N_14711,N_14717);
or U15241 (N_15241,N_14959,N_14307);
and U15242 (N_15242,N_14556,N_14927);
nor U15243 (N_15243,N_14485,N_14356);
and U15244 (N_15244,N_14864,N_14599);
nand U15245 (N_15245,N_14304,N_14639);
and U15246 (N_15246,N_14394,N_14252);
and U15247 (N_15247,N_14374,N_14080);
xor U15248 (N_15248,N_14657,N_14475);
xor U15249 (N_15249,N_14176,N_14828);
nand U15250 (N_15250,N_14999,N_14067);
or U15251 (N_15251,N_14790,N_14270);
xnor U15252 (N_15252,N_14525,N_14853);
nor U15253 (N_15253,N_14124,N_14269);
and U15254 (N_15254,N_14446,N_14951);
nand U15255 (N_15255,N_14191,N_14313);
and U15256 (N_15256,N_14675,N_14502);
nor U15257 (N_15257,N_14743,N_14789);
xor U15258 (N_15258,N_14941,N_14184);
nor U15259 (N_15259,N_14060,N_14765);
nor U15260 (N_15260,N_14618,N_14072);
nor U15261 (N_15261,N_14889,N_14779);
or U15262 (N_15262,N_14294,N_14022);
nor U15263 (N_15263,N_14965,N_14897);
nor U15264 (N_15264,N_14760,N_14108);
nor U15265 (N_15265,N_14266,N_14054);
or U15266 (N_15266,N_14960,N_14459);
xor U15267 (N_15267,N_14247,N_14352);
nor U15268 (N_15268,N_14571,N_14358);
or U15269 (N_15269,N_14027,N_14259);
and U15270 (N_15270,N_14089,N_14665);
nand U15271 (N_15271,N_14869,N_14268);
nor U15272 (N_15272,N_14852,N_14561);
and U15273 (N_15273,N_14788,N_14450);
nand U15274 (N_15274,N_14289,N_14763);
nor U15275 (N_15275,N_14196,N_14172);
xnor U15276 (N_15276,N_14829,N_14166);
nor U15277 (N_15277,N_14169,N_14361);
xnor U15278 (N_15278,N_14862,N_14855);
nor U15279 (N_15279,N_14968,N_14633);
and U15280 (N_15280,N_14335,N_14402);
nand U15281 (N_15281,N_14100,N_14983);
or U15282 (N_15282,N_14342,N_14336);
and U15283 (N_15283,N_14773,N_14219);
or U15284 (N_15284,N_14004,N_14907);
or U15285 (N_15285,N_14557,N_14306);
xor U15286 (N_15286,N_14878,N_14918);
and U15287 (N_15287,N_14581,N_14553);
and U15288 (N_15288,N_14042,N_14230);
nor U15289 (N_15289,N_14428,N_14714);
nor U15290 (N_15290,N_14649,N_14321);
nand U15291 (N_15291,N_14183,N_14243);
nand U15292 (N_15292,N_14458,N_14232);
nand U15293 (N_15293,N_14681,N_14664);
or U15294 (N_15294,N_14175,N_14791);
nor U15295 (N_15295,N_14998,N_14716);
nor U15296 (N_15296,N_14609,N_14030);
and U15297 (N_15297,N_14744,N_14146);
xor U15298 (N_15298,N_14708,N_14745);
nand U15299 (N_15299,N_14683,N_14926);
nand U15300 (N_15300,N_14189,N_14201);
and U15301 (N_15301,N_14537,N_14253);
xor U15302 (N_15302,N_14515,N_14707);
nor U15303 (N_15303,N_14122,N_14011);
nand U15304 (N_15304,N_14392,N_14323);
xor U15305 (N_15305,N_14549,N_14695);
nor U15306 (N_15306,N_14126,N_14302);
nand U15307 (N_15307,N_14512,N_14049);
and U15308 (N_15308,N_14691,N_14135);
xor U15309 (N_15309,N_14390,N_14391);
and U15310 (N_15310,N_14290,N_14612);
and U15311 (N_15311,N_14939,N_14585);
or U15312 (N_15312,N_14319,N_14759);
nor U15313 (N_15313,N_14837,N_14069);
nor U15314 (N_15314,N_14387,N_14035);
or U15315 (N_15315,N_14043,N_14874);
or U15316 (N_15316,N_14041,N_14911);
or U15317 (N_15317,N_14573,N_14931);
or U15318 (N_15318,N_14685,N_14341);
xnor U15319 (N_15319,N_14493,N_14641);
nor U15320 (N_15320,N_14299,N_14891);
nor U15321 (N_15321,N_14756,N_14133);
or U15322 (N_15322,N_14154,N_14956);
xnor U15323 (N_15323,N_14659,N_14651);
xor U15324 (N_15324,N_14021,N_14417);
xnor U15325 (N_15325,N_14296,N_14005);
nand U15326 (N_15326,N_14900,N_14236);
xnor U15327 (N_15327,N_14979,N_14574);
nor U15328 (N_15328,N_14844,N_14577);
nand U15329 (N_15329,N_14476,N_14188);
and U15330 (N_15330,N_14116,N_14895);
nand U15331 (N_15331,N_14576,N_14637);
and U15332 (N_15332,N_14255,N_14461);
and U15333 (N_15333,N_14647,N_14975);
or U15334 (N_15334,N_14013,N_14993);
nand U15335 (N_15335,N_14519,N_14608);
nor U15336 (N_15336,N_14239,N_14118);
and U15337 (N_15337,N_14231,N_14368);
xor U15338 (N_15338,N_14928,N_14480);
nand U15339 (N_15339,N_14957,N_14636);
nor U15340 (N_15340,N_14970,N_14466);
and U15341 (N_15341,N_14325,N_14052);
xor U15342 (N_15342,N_14455,N_14367);
and U15343 (N_15343,N_14888,N_14317);
and U15344 (N_15344,N_14162,N_14531);
or U15345 (N_15345,N_14360,N_14318);
nor U15346 (N_15346,N_14514,N_14003);
and U15347 (N_15347,N_14065,N_14972);
xnor U15348 (N_15348,N_14286,N_14752);
xnor U15349 (N_15349,N_14622,N_14010);
xor U15350 (N_15350,N_14454,N_14948);
xor U15351 (N_15351,N_14497,N_14284);
nor U15352 (N_15352,N_14832,N_14624);
nor U15353 (N_15353,N_14923,N_14916);
nor U15354 (N_15354,N_14471,N_14034);
nor U15355 (N_15355,N_14322,N_14703);
nand U15356 (N_15356,N_14217,N_14111);
xor U15357 (N_15357,N_14767,N_14901);
or U15358 (N_15358,N_14425,N_14545);
or U15359 (N_15359,N_14644,N_14634);
nand U15360 (N_15360,N_14835,N_14120);
nand U15361 (N_15361,N_14103,N_14595);
nand U15362 (N_15362,N_14962,N_14327);
xnor U15363 (N_15363,N_14969,N_14380);
nor U15364 (N_15364,N_14807,N_14047);
xor U15365 (N_15365,N_14393,N_14804);
xnor U15366 (N_15366,N_14399,N_14109);
or U15367 (N_15367,N_14523,N_14437);
nor U15368 (N_15368,N_14452,N_14725);
and U15369 (N_15369,N_14748,N_14197);
and U15370 (N_15370,N_14833,N_14798);
and U15371 (N_15371,N_14403,N_14524);
and U15372 (N_15372,N_14382,N_14797);
nand U15373 (N_15373,N_14751,N_14163);
or U15374 (N_15374,N_14943,N_14996);
and U15375 (N_15375,N_14248,N_14204);
or U15376 (N_15376,N_14879,N_14337);
and U15377 (N_15377,N_14737,N_14221);
nor U15378 (N_15378,N_14540,N_14406);
and U15379 (N_15379,N_14460,N_14924);
and U15380 (N_15380,N_14037,N_14601);
xnor U15381 (N_15381,N_14280,N_14141);
xnor U15382 (N_15382,N_14016,N_14566);
or U15383 (N_15383,N_14586,N_14059);
and U15384 (N_15384,N_14784,N_14139);
xor U15385 (N_15385,N_14210,N_14263);
xor U15386 (N_15386,N_14152,N_14946);
nand U15387 (N_15387,N_14815,N_14144);
nand U15388 (N_15388,N_14383,N_14371);
and U15389 (N_15389,N_14101,N_14588);
and U15390 (N_15390,N_14971,N_14806);
nor U15391 (N_15391,N_14872,N_14145);
xnor U15392 (N_15392,N_14589,N_14850);
or U15393 (N_15393,N_14674,N_14158);
and U15394 (N_15394,N_14696,N_14315);
xnor U15395 (N_15395,N_14291,N_14503);
nand U15396 (N_15396,N_14629,N_14702);
and U15397 (N_15397,N_14397,N_14205);
and U15398 (N_15398,N_14663,N_14088);
nor U15399 (N_15399,N_14771,N_14349);
xnor U15400 (N_15400,N_14339,N_14218);
nor U15401 (N_15401,N_14799,N_14934);
nand U15402 (N_15402,N_14200,N_14314);
nand U15403 (N_15403,N_14843,N_14831);
nand U15404 (N_15404,N_14870,N_14224);
or U15405 (N_15405,N_14050,N_14256);
nor U15406 (N_15406,N_14039,N_14802);
and U15407 (N_15407,N_14792,N_14669);
nor U15408 (N_15408,N_14477,N_14884);
nor U15409 (N_15409,N_14977,N_14223);
or U15410 (N_15410,N_14821,N_14875);
nand U15411 (N_15411,N_14578,N_14954);
nand U15412 (N_15412,N_14464,N_14930);
nand U15413 (N_15413,N_14272,N_14494);
and U15414 (N_15414,N_14206,N_14351);
xnor U15415 (N_15415,N_14604,N_14445);
and U15416 (N_15416,N_14728,N_14892);
nand U15417 (N_15417,N_14778,N_14984);
or U15418 (N_15418,N_14536,N_14305);
or U15419 (N_15419,N_14226,N_14679);
xnor U15420 (N_15420,N_14643,N_14575);
xnor U15421 (N_15421,N_14245,N_14758);
nand U15422 (N_15422,N_14451,N_14813);
and U15423 (N_15423,N_14311,N_14355);
nand U15424 (N_15424,N_14246,N_14227);
or U15425 (N_15425,N_14142,N_14370);
and U15426 (N_15426,N_14125,N_14922);
or U15427 (N_15427,N_14441,N_14543);
xnor U15428 (N_15428,N_14165,N_14738);
nor U15429 (N_15429,N_14482,N_14409);
nor U15430 (N_15430,N_14254,N_14873);
and U15431 (N_15431,N_14824,N_14216);
xor U15432 (N_15432,N_14932,N_14718);
and U15433 (N_15433,N_14064,N_14650);
nand U15434 (N_15434,N_14570,N_14366);
or U15435 (N_15435,N_14161,N_14436);
xnor U15436 (N_15436,N_14347,N_14081);
or U15437 (N_15437,N_14238,N_14202);
nor U15438 (N_15438,N_14419,N_14865);
and U15439 (N_15439,N_14661,N_14655);
nand U15440 (N_15440,N_14283,N_14068);
nand U15441 (N_15441,N_14472,N_14780);
and U15442 (N_15442,N_14456,N_14724);
xnor U15443 (N_15443,N_14271,N_14070);
xnor U15444 (N_15444,N_14559,N_14182);
xnor U15445 (N_15445,N_14359,N_14036);
nand U15446 (N_15446,N_14989,N_14602);
and U15447 (N_15447,N_14353,N_14795);
and U15448 (N_15448,N_14008,N_14632);
xor U15449 (N_15449,N_14988,N_14408);
and U15450 (N_15450,N_14241,N_14619);
or U15451 (N_15451,N_14583,N_14157);
nand U15452 (N_15452,N_14781,N_14413);
nor U15453 (N_15453,N_14982,N_14214);
and U15454 (N_15454,N_14741,N_14265);
xor U15455 (N_15455,N_14777,N_14301);
nor U15456 (N_15456,N_14754,N_14893);
and U15457 (N_15457,N_14757,N_14261);
nand U15458 (N_15458,N_14012,N_14896);
and U15459 (N_15459,N_14522,N_14398);
nor U15460 (N_15460,N_14611,N_14656);
and U15461 (N_15461,N_14019,N_14354);
and U15462 (N_15462,N_14121,N_14228);
xor U15463 (N_15463,N_14400,N_14418);
xor U15464 (N_15464,N_14727,N_14348);
and U15465 (N_15465,N_14671,N_14490);
and U15466 (N_15466,N_14562,N_14112);
nor U15467 (N_15467,N_14560,N_14908);
nor U15468 (N_15468,N_14440,N_14138);
nor U15469 (N_15469,N_14929,N_14132);
nand U15470 (N_15470,N_14181,N_14225);
nor U15471 (N_15471,N_14564,N_14468);
and U15472 (N_15472,N_14063,N_14483);
xnor U15473 (N_15473,N_14823,N_14848);
xor U15474 (N_15474,N_14002,N_14364);
nor U15475 (N_15475,N_14106,N_14584);
nor U15476 (N_15476,N_14782,N_14508);
nor U15477 (N_15477,N_14362,N_14365);
and U15478 (N_15478,N_14682,N_14257);
and U15479 (N_15479,N_14028,N_14278);
xnor U15480 (N_15480,N_14338,N_14890);
xnor U15481 (N_15481,N_14431,N_14186);
nor U15482 (N_15482,N_14015,N_14505);
xnor U15483 (N_15483,N_14024,N_14933);
nand U15484 (N_15484,N_14846,N_14071);
and U15485 (N_15485,N_14686,N_14385);
nand U15486 (N_15486,N_14859,N_14082);
or U15487 (N_15487,N_14736,N_14114);
and U15488 (N_15488,N_14501,N_14453);
nor U15489 (N_15489,N_14168,N_14914);
and U15490 (N_15490,N_14594,N_14507);
nor U15491 (N_15491,N_14689,N_14130);
and U15492 (N_15492,N_14424,N_14592);
nor U15493 (N_15493,N_14642,N_14630);
nor U15494 (N_15494,N_14700,N_14886);
xnor U15495 (N_15495,N_14433,N_14628);
nand U15496 (N_15496,N_14287,N_14495);
xnor U15497 (N_15497,N_14432,N_14876);
or U15498 (N_15498,N_14530,N_14701);
or U15499 (N_15499,N_14580,N_14871);
nor U15500 (N_15500,N_14013,N_14209);
and U15501 (N_15501,N_14244,N_14232);
nor U15502 (N_15502,N_14751,N_14496);
nand U15503 (N_15503,N_14491,N_14030);
or U15504 (N_15504,N_14680,N_14257);
xor U15505 (N_15505,N_14467,N_14724);
xnor U15506 (N_15506,N_14270,N_14878);
nor U15507 (N_15507,N_14941,N_14420);
and U15508 (N_15508,N_14535,N_14156);
nor U15509 (N_15509,N_14203,N_14948);
xor U15510 (N_15510,N_14740,N_14185);
nor U15511 (N_15511,N_14585,N_14100);
xnor U15512 (N_15512,N_14234,N_14903);
xor U15513 (N_15513,N_14086,N_14745);
nand U15514 (N_15514,N_14989,N_14798);
or U15515 (N_15515,N_14327,N_14982);
and U15516 (N_15516,N_14438,N_14347);
and U15517 (N_15517,N_14187,N_14891);
nor U15518 (N_15518,N_14564,N_14451);
xnor U15519 (N_15519,N_14300,N_14072);
or U15520 (N_15520,N_14670,N_14930);
nand U15521 (N_15521,N_14027,N_14690);
and U15522 (N_15522,N_14373,N_14936);
nand U15523 (N_15523,N_14418,N_14610);
nor U15524 (N_15524,N_14886,N_14854);
nand U15525 (N_15525,N_14942,N_14926);
xor U15526 (N_15526,N_14678,N_14611);
and U15527 (N_15527,N_14171,N_14308);
nand U15528 (N_15528,N_14547,N_14126);
nand U15529 (N_15529,N_14959,N_14779);
nand U15530 (N_15530,N_14492,N_14098);
xnor U15531 (N_15531,N_14510,N_14373);
nand U15532 (N_15532,N_14870,N_14753);
and U15533 (N_15533,N_14331,N_14946);
and U15534 (N_15534,N_14277,N_14790);
or U15535 (N_15535,N_14940,N_14005);
xor U15536 (N_15536,N_14968,N_14236);
or U15537 (N_15537,N_14339,N_14929);
and U15538 (N_15538,N_14509,N_14538);
nand U15539 (N_15539,N_14965,N_14421);
xnor U15540 (N_15540,N_14062,N_14897);
nand U15541 (N_15541,N_14826,N_14660);
nor U15542 (N_15542,N_14414,N_14732);
or U15543 (N_15543,N_14267,N_14305);
nand U15544 (N_15544,N_14007,N_14917);
xnor U15545 (N_15545,N_14948,N_14342);
nand U15546 (N_15546,N_14166,N_14279);
xnor U15547 (N_15547,N_14407,N_14343);
and U15548 (N_15548,N_14693,N_14179);
nand U15549 (N_15549,N_14878,N_14680);
and U15550 (N_15550,N_14672,N_14058);
xor U15551 (N_15551,N_14867,N_14079);
xor U15552 (N_15552,N_14616,N_14440);
nand U15553 (N_15553,N_14337,N_14757);
and U15554 (N_15554,N_14546,N_14288);
nand U15555 (N_15555,N_14319,N_14979);
or U15556 (N_15556,N_14660,N_14009);
xor U15557 (N_15557,N_14090,N_14489);
xor U15558 (N_15558,N_14610,N_14599);
and U15559 (N_15559,N_14941,N_14521);
and U15560 (N_15560,N_14172,N_14671);
nand U15561 (N_15561,N_14036,N_14450);
and U15562 (N_15562,N_14195,N_14980);
and U15563 (N_15563,N_14601,N_14215);
nor U15564 (N_15564,N_14009,N_14103);
and U15565 (N_15565,N_14977,N_14045);
and U15566 (N_15566,N_14624,N_14456);
xnor U15567 (N_15567,N_14844,N_14345);
nor U15568 (N_15568,N_14294,N_14745);
xnor U15569 (N_15569,N_14330,N_14928);
or U15570 (N_15570,N_14309,N_14743);
nor U15571 (N_15571,N_14821,N_14519);
nand U15572 (N_15572,N_14478,N_14025);
nand U15573 (N_15573,N_14136,N_14023);
nand U15574 (N_15574,N_14761,N_14264);
and U15575 (N_15575,N_14330,N_14202);
and U15576 (N_15576,N_14821,N_14474);
xnor U15577 (N_15577,N_14714,N_14591);
nor U15578 (N_15578,N_14904,N_14533);
nor U15579 (N_15579,N_14978,N_14868);
nor U15580 (N_15580,N_14646,N_14109);
nor U15581 (N_15581,N_14934,N_14341);
nand U15582 (N_15582,N_14877,N_14180);
nor U15583 (N_15583,N_14631,N_14863);
or U15584 (N_15584,N_14710,N_14094);
and U15585 (N_15585,N_14578,N_14827);
xnor U15586 (N_15586,N_14868,N_14688);
or U15587 (N_15587,N_14343,N_14138);
or U15588 (N_15588,N_14598,N_14557);
or U15589 (N_15589,N_14126,N_14466);
or U15590 (N_15590,N_14645,N_14619);
xor U15591 (N_15591,N_14578,N_14411);
nand U15592 (N_15592,N_14286,N_14200);
or U15593 (N_15593,N_14821,N_14156);
or U15594 (N_15594,N_14043,N_14884);
and U15595 (N_15595,N_14314,N_14655);
or U15596 (N_15596,N_14715,N_14723);
or U15597 (N_15597,N_14748,N_14758);
xnor U15598 (N_15598,N_14188,N_14530);
nor U15599 (N_15599,N_14224,N_14433);
and U15600 (N_15600,N_14079,N_14177);
nand U15601 (N_15601,N_14154,N_14405);
xnor U15602 (N_15602,N_14166,N_14858);
and U15603 (N_15603,N_14151,N_14450);
xor U15604 (N_15604,N_14961,N_14005);
or U15605 (N_15605,N_14689,N_14529);
and U15606 (N_15606,N_14365,N_14102);
nand U15607 (N_15607,N_14495,N_14624);
nor U15608 (N_15608,N_14738,N_14823);
xnor U15609 (N_15609,N_14079,N_14542);
and U15610 (N_15610,N_14156,N_14587);
xor U15611 (N_15611,N_14728,N_14309);
and U15612 (N_15612,N_14536,N_14013);
nand U15613 (N_15613,N_14968,N_14332);
nor U15614 (N_15614,N_14562,N_14900);
or U15615 (N_15615,N_14386,N_14294);
xnor U15616 (N_15616,N_14279,N_14230);
or U15617 (N_15617,N_14364,N_14523);
nand U15618 (N_15618,N_14553,N_14198);
xor U15619 (N_15619,N_14909,N_14403);
nand U15620 (N_15620,N_14949,N_14758);
nor U15621 (N_15621,N_14794,N_14180);
nor U15622 (N_15622,N_14149,N_14306);
and U15623 (N_15623,N_14151,N_14688);
xor U15624 (N_15624,N_14694,N_14913);
xnor U15625 (N_15625,N_14775,N_14308);
nand U15626 (N_15626,N_14955,N_14056);
nor U15627 (N_15627,N_14043,N_14734);
or U15628 (N_15628,N_14357,N_14417);
nor U15629 (N_15629,N_14601,N_14305);
and U15630 (N_15630,N_14421,N_14998);
or U15631 (N_15631,N_14131,N_14164);
and U15632 (N_15632,N_14567,N_14779);
or U15633 (N_15633,N_14057,N_14562);
xnor U15634 (N_15634,N_14622,N_14024);
and U15635 (N_15635,N_14327,N_14279);
nand U15636 (N_15636,N_14524,N_14788);
or U15637 (N_15637,N_14292,N_14536);
nand U15638 (N_15638,N_14213,N_14778);
xnor U15639 (N_15639,N_14092,N_14611);
and U15640 (N_15640,N_14356,N_14918);
xnor U15641 (N_15641,N_14868,N_14955);
xor U15642 (N_15642,N_14866,N_14038);
and U15643 (N_15643,N_14704,N_14755);
or U15644 (N_15644,N_14859,N_14623);
or U15645 (N_15645,N_14814,N_14364);
nor U15646 (N_15646,N_14797,N_14036);
nor U15647 (N_15647,N_14032,N_14197);
xor U15648 (N_15648,N_14881,N_14027);
nor U15649 (N_15649,N_14573,N_14957);
nand U15650 (N_15650,N_14134,N_14334);
or U15651 (N_15651,N_14533,N_14179);
nor U15652 (N_15652,N_14633,N_14809);
xnor U15653 (N_15653,N_14934,N_14438);
nor U15654 (N_15654,N_14988,N_14912);
and U15655 (N_15655,N_14762,N_14280);
or U15656 (N_15656,N_14738,N_14017);
nor U15657 (N_15657,N_14084,N_14327);
nand U15658 (N_15658,N_14668,N_14393);
nand U15659 (N_15659,N_14118,N_14990);
nor U15660 (N_15660,N_14591,N_14636);
nor U15661 (N_15661,N_14276,N_14536);
or U15662 (N_15662,N_14934,N_14252);
nand U15663 (N_15663,N_14526,N_14403);
nor U15664 (N_15664,N_14357,N_14393);
or U15665 (N_15665,N_14733,N_14931);
xnor U15666 (N_15666,N_14141,N_14786);
or U15667 (N_15667,N_14736,N_14141);
xnor U15668 (N_15668,N_14318,N_14400);
nand U15669 (N_15669,N_14528,N_14884);
nand U15670 (N_15670,N_14752,N_14991);
and U15671 (N_15671,N_14888,N_14120);
and U15672 (N_15672,N_14787,N_14885);
and U15673 (N_15673,N_14220,N_14445);
nand U15674 (N_15674,N_14245,N_14750);
xnor U15675 (N_15675,N_14955,N_14532);
nor U15676 (N_15676,N_14762,N_14281);
nor U15677 (N_15677,N_14936,N_14360);
or U15678 (N_15678,N_14981,N_14428);
nor U15679 (N_15679,N_14268,N_14592);
and U15680 (N_15680,N_14858,N_14668);
and U15681 (N_15681,N_14426,N_14829);
or U15682 (N_15682,N_14885,N_14660);
xor U15683 (N_15683,N_14790,N_14350);
nand U15684 (N_15684,N_14034,N_14865);
or U15685 (N_15685,N_14516,N_14849);
and U15686 (N_15686,N_14131,N_14953);
or U15687 (N_15687,N_14465,N_14217);
and U15688 (N_15688,N_14602,N_14907);
nand U15689 (N_15689,N_14049,N_14738);
nand U15690 (N_15690,N_14260,N_14043);
or U15691 (N_15691,N_14410,N_14366);
or U15692 (N_15692,N_14389,N_14137);
or U15693 (N_15693,N_14669,N_14492);
xnor U15694 (N_15694,N_14726,N_14157);
nand U15695 (N_15695,N_14648,N_14000);
and U15696 (N_15696,N_14670,N_14113);
nor U15697 (N_15697,N_14404,N_14468);
xor U15698 (N_15698,N_14613,N_14211);
and U15699 (N_15699,N_14812,N_14651);
nand U15700 (N_15700,N_14901,N_14990);
nand U15701 (N_15701,N_14515,N_14686);
nand U15702 (N_15702,N_14615,N_14967);
nand U15703 (N_15703,N_14288,N_14882);
and U15704 (N_15704,N_14207,N_14702);
nor U15705 (N_15705,N_14920,N_14010);
or U15706 (N_15706,N_14178,N_14496);
nor U15707 (N_15707,N_14858,N_14304);
and U15708 (N_15708,N_14588,N_14947);
and U15709 (N_15709,N_14718,N_14745);
nand U15710 (N_15710,N_14321,N_14024);
and U15711 (N_15711,N_14902,N_14071);
nor U15712 (N_15712,N_14423,N_14373);
nand U15713 (N_15713,N_14166,N_14088);
nand U15714 (N_15714,N_14949,N_14600);
nand U15715 (N_15715,N_14499,N_14449);
nand U15716 (N_15716,N_14489,N_14532);
and U15717 (N_15717,N_14529,N_14618);
nand U15718 (N_15718,N_14871,N_14089);
nor U15719 (N_15719,N_14419,N_14578);
or U15720 (N_15720,N_14683,N_14234);
nand U15721 (N_15721,N_14952,N_14388);
and U15722 (N_15722,N_14254,N_14471);
nor U15723 (N_15723,N_14947,N_14034);
or U15724 (N_15724,N_14622,N_14935);
or U15725 (N_15725,N_14554,N_14603);
and U15726 (N_15726,N_14077,N_14896);
xor U15727 (N_15727,N_14754,N_14461);
nor U15728 (N_15728,N_14131,N_14132);
or U15729 (N_15729,N_14158,N_14774);
nand U15730 (N_15730,N_14934,N_14574);
xor U15731 (N_15731,N_14392,N_14621);
xnor U15732 (N_15732,N_14793,N_14942);
nand U15733 (N_15733,N_14917,N_14637);
nor U15734 (N_15734,N_14802,N_14455);
xor U15735 (N_15735,N_14280,N_14094);
xor U15736 (N_15736,N_14150,N_14811);
nor U15737 (N_15737,N_14148,N_14987);
nand U15738 (N_15738,N_14872,N_14564);
nand U15739 (N_15739,N_14039,N_14388);
and U15740 (N_15740,N_14007,N_14621);
nor U15741 (N_15741,N_14780,N_14949);
xor U15742 (N_15742,N_14345,N_14994);
and U15743 (N_15743,N_14754,N_14519);
nand U15744 (N_15744,N_14301,N_14320);
nor U15745 (N_15745,N_14169,N_14389);
or U15746 (N_15746,N_14459,N_14882);
or U15747 (N_15747,N_14461,N_14741);
or U15748 (N_15748,N_14402,N_14897);
or U15749 (N_15749,N_14813,N_14385);
and U15750 (N_15750,N_14100,N_14760);
xnor U15751 (N_15751,N_14588,N_14928);
or U15752 (N_15752,N_14761,N_14414);
or U15753 (N_15753,N_14218,N_14881);
and U15754 (N_15754,N_14749,N_14645);
or U15755 (N_15755,N_14303,N_14074);
xnor U15756 (N_15756,N_14864,N_14174);
nor U15757 (N_15757,N_14010,N_14949);
nor U15758 (N_15758,N_14242,N_14289);
xor U15759 (N_15759,N_14654,N_14988);
nor U15760 (N_15760,N_14186,N_14781);
nand U15761 (N_15761,N_14795,N_14267);
nor U15762 (N_15762,N_14153,N_14550);
nand U15763 (N_15763,N_14176,N_14108);
nand U15764 (N_15764,N_14319,N_14936);
nor U15765 (N_15765,N_14940,N_14970);
or U15766 (N_15766,N_14303,N_14277);
and U15767 (N_15767,N_14069,N_14430);
xor U15768 (N_15768,N_14219,N_14377);
nor U15769 (N_15769,N_14993,N_14024);
nor U15770 (N_15770,N_14781,N_14157);
or U15771 (N_15771,N_14079,N_14855);
xnor U15772 (N_15772,N_14231,N_14163);
nand U15773 (N_15773,N_14789,N_14723);
or U15774 (N_15774,N_14178,N_14415);
nor U15775 (N_15775,N_14178,N_14963);
xor U15776 (N_15776,N_14685,N_14893);
nor U15777 (N_15777,N_14407,N_14706);
and U15778 (N_15778,N_14876,N_14392);
nand U15779 (N_15779,N_14782,N_14003);
nor U15780 (N_15780,N_14806,N_14594);
or U15781 (N_15781,N_14743,N_14389);
or U15782 (N_15782,N_14066,N_14208);
nor U15783 (N_15783,N_14633,N_14408);
xnor U15784 (N_15784,N_14172,N_14555);
and U15785 (N_15785,N_14265,N_14239);
xor U15786 (N_15786,N_14271,N_14359);
and U15787 (N_15787,N_14626,N_14690);
nor U15788 (N_15788,N_14041,N_14113);
nor U15789 (N_15789,N_14832,N_14214);
and U15790 (N_15790,N_14049,N_14892);
nand U15791 (N_15791,N_14977,N_14893);
or U15792 (N_15792,N_14639,N_14373);
xor U15793 (N_15793,N_14307,N_14319);
nor U15794 (N_15794,N_14060,N_14751);
xnor U15795 (N_15795,N_14267,N_14974);
or U15796 (N_15796,N_14788,N_14631);
nand U15797 (N_15797,N_14144,N_14556);
nor U15798 (N_15798,N_14688,N_14741);
and U15799 (N_15799,N_14321,N_14670);
and U15800 (N_15800,N_14194,N_14773);
or U15801 (N_15801,N_14610,N_14884);
and U15802 (N_15802,N_14864,N_14146);
and U15803 (N_15803,N_14326,N_14495);
nor U15804 (N_15804,N_14839,N_14360);
nor U15805 (N_15805,N_14297,N_14518);
and U15806 (N_15806,N_14467,N_14862);
nor U15807 (N_15807,N_14096,N_14425);
or U15808 (N_15808,N_14883,N_14998);
nor U15809 (N_15809,N_14541,N_14146);
or U15810 (N_15810,N_14931,N_14882);
or U15811 (N_15811,N_14433,N_14506);
and U15812 (N_15812,N_14925,N_14362);
nor U15813 (N_15813,N_14889,N_14147);
xor U15814 (N_15814,N_14472,N_14228);
xnor U15815 (N_15815,N_14431,N_14356);
and U15816 (N_15816,N_14910,N_14306);
and U15817 (N_15817,N_14067,N_14580);
nor U15818 (N_15818,N_14810,N_14127);
nor U15819 (N_15819,N_14173,N_14866);
or U15820 (N_15820,N_14817,N_14999);
or U15821 (N_15821,N_14321,N_14495);
nor U15822 (N_15822,N_14767,N_14827);
or U15823 (N_15823,N_14959,N_14028);
nand U15824 (N_15824,N_14323,N_14734);
or U15825 (N_15825,N_14387,N_14113);
nand U15826 (N_15826,N_14210,N_14264);
xor U15827 (N_15827,N_14372,N_14143);
and U15828 (N_15828,N_14359,N_14537);
nand U15829 (N_15829,N_14457,N_14779);
and U15830 (N_15830,N_14916,N_14010);
xor U15831 (N_15831,N_14298,N_14056);
xnor U15832 (N_15832,N_14764,N_14992);
and U15833 (N_15833,N_14705,N_14082);
nand U15834 (N_15834,N_14337,N_14041);
and U15835 (N_15835,N_14472,N_14174);
nor U15836 (N_15836,N_14661,N_14441);
nand U15837 (N_15837,N_14228,N_14018);
xnor U15838 (N_15838,N_14077,N_14158);
nor U15839 (N_15839,N_14791,N_14997);
nor U15840 (N_15840,N_14033,N_14536);
and U15841 (N_15841,N_14959,N_14533);
nor U15842 (N_15842,N_14808,N_14369);
xor U15843 (N_15843,N_14153,N_14927);
and U15844 (N_15844,N_14918,N_14518);
nand U15845 (N_15845,N_14547,N_14534);
nand U15846 (N_15846,N_14510,N_14300);
or U15847 (N_15847,N_14063,N_14924);
xor U15848 (N_15848,N_14561,N_14299);
and U15849 (N_15849,N_14871,N_14378);
nand U15850 (N_15850,N_14518,N_14203);
nand U15851 (N_15851,N_14943,N_14857);
and U15852 (N_15852,N_14621,N_14063);
or U15853 (N_15853,N_14965,N_14143);
nor U15854 (N_15854,N_14235,N_14465);
and U15855 (N_15855,N_14784,N_14914);
and U15856 (N_15856,N_14757,N_14072);
nand U15857 (N_15857,N_14283,N_14644);
and U15858 (N_15858,N_14812,N_14600);
xor U15859 (N_15859,N_14413,N_14616);
and U15860 (N_15860,N_14238,N_14389);
or U15861 (N_15861,N_14000,N_14614);
xor U15862 (N_15862,N_14957,N_14802);
and U15863 (N_15863,N_14850,N_14995);
nor U15864 (N_15864,N_14484,N_14285);
nand U15865 (N_15865,N_14487,N_14660);
and U15866 (N_15866,N_14038,N_14848);
or U15867 (N_15867,N_14916,N_14869);
nor U15868 (N_15868,N_14035,N_14149);
xor U15869 (N_15869,N_14974,N_14521);
and U15870 (N_15870,N_14371,N_14380);
nand U15871 (N_15871,N_14710,N_14225);
or U15872 (N_15872,N_14775,N_14072);
nand U15873 (N_15873,N_14196,N_14318);
nor U15874 (N_15874,N_14918,N_14095);
nor U15875 (N_15875,N_14216,N_14570);
nand U15876 (N_15876,N_14596,N_14967);
nand U15877 (N_15877,N_14565,N_14045);
xnor U15878 (N_15878,N_14046,N_14337);
xnor U15879 (N_15879,N_14072,N_14689);
nor U15880 (N_15880,N_14403,N_14504);
or U15881 (N_15881,N_14318,N_14214);
nand U15882 (N_15882,N_14062,N_14448);
xnor U15883 (N_15883,N_14413,N_14315);
xnor U15884 (N_15884,N_14375,N_14061);
or U15885 (N_15885,N_14078,N_14707);
nand U15886 (N_15886,N_14438,N_14087);
xnor U15887 (N_15887,N_14684,N_14651);
xor U15888 (N_15888,N_14075,N_14761);
nand U15889 (N_15889,N_14109,N_14084);
nor U15890 (N_15890,N_14914,N_14933);
xnor U15891 (N_15891,N_14025,N_14733);
nor U15892 (N_15892,N_14363,N_14336);
nor U15893 (N_15893,N_14228,N_14848);
or U15894 (N_15894,N_14597,N_14914);
or U15895 (N_15895,N_14044,N_14710);
nand U15896 (N_15896,N_14883,N_14968);
or U15897 (N_15897,N_14166,N_14731);
nor U15898 (N_15898,N_14028,N_14211);
nand U15899 (N_15899,N_14777,N_14740);
nor U15900 (N_15900,N_14620,N_14112);
xnor U15901 (N_15901,N_14024,N_14635);
xnor U15902 (N_15902,N_14526,N_14259);
nand U15903 (N_15903,N_14277,N_14756);
xor U15904 (N_15904,N_14378,N_14380);
nor U15905 (N_15905,N_14327,N_14917);
or U15906 (N_15906,N_14689,N_14649);
and U15907 (N_15907,N_14584,N_14249);
and U15908 (N_15908,N_14071,N_14724);
or U15909 (N_15909,N_14162,N_14254);
nand U15910 (N_15910,N_14342,N_14956);
and U15911 (N_15911,N_14796,N_14026);
nand U15912 (N_15912,N_14166,N_14647);
and U15913 (N_15913,N_14576,N_14289);
or U15914 (N_15914,N_14148,N_14008);
nand U15915 (N_15915,N_14808,N_14798);
and U15916 (N_15916,N_14631,N_14300);
and U15917 (N_15917,N_14606,N_14193);
nor U15918 (N_15918,N_14679,N_14681);
nand U15919 (N_15919,N_14875,N_14704);
xor U15920 (N_15920,N_14063,N_14539);
nand U15921 (N_15921,N_14448,N_14144);
xor U15922 (N_15922,N_14333,N_14849);
xnor U15923 (N_15923,N_14617,N_14043);
and U15924 (N_15924,N_14423,N_14600);
xor U15925 (N_15925,N_14115,N_14086);
or U15926 (N_15926,N_14178,N_14382);
nor U15927 (N_15927,N_14840,N_14720);
xor U15928 (N_15928,N_14412,N_14049);
nand U15929 (N_15929,N_14999,N_14720);
xor U15930 (N_15930,N_14528,N_14939);
nand U15931 (N_15931,N_14775,N_14844);
nand U15932 (N_15932,N_14000,N_14465);
and U15933 (N_15933,N_14891,N_14430);
or U15934 (N_15934,N_14511,N_14171);
or U15935 (N_15935,N_14567,N_14087);
and U15936 (N_15936,N_14898,N_14864);
or U15937 (N_15937,N_14031,N_14382);
and U15938 (N_15938,N_14682,N_14098);
or U15939 (N_15939,N_14163,N_14837);
xor U15940 (N_15940,N_14979,N_14377);
and U15941 (N_15941,N_14066,N_14082);
xor U15942 (N_15942,N_14316,N_14680);
nand U15943 (N_15943,N_14311,N_14398);
nand U15944 (N_15944,N_14196,N_14238);
nand U15945 (N_15945,N_14386,N_14399);
xnor U15946 (N_15946,N_14154,N_14324);
nor U15947 (N_15947,N_14319,N_14310);
nand U15948 (N_15948,N_14592,N_14852);
xor U15949 (N_15949,N_14336,N_14985);
or U15950 (N_15950,N_14455,N_14684);
nand U15951 (N_15951,N_14172,N_14989);
nand U15952 (N_15952,N_14695,N_14404);
xor U15953 (N_15953,N_14433,N_14544);
xor U15954 (N_15954,N_14742,N_14109);
nor U15955 (N_15955,N_14287,N_14448);
and U15956 (N_15956,N_14298,N_14647);
nor U15957 (N_15957,N_14047,N_14656);
nand U15958 (N_15958,N_14177,N_14469);
and U15959 (N_15959,N_14681,N_14087);
xor U15960 (N_15960,N_14624,N_14383);
nand U15961 (N_15961,N_14022,N_14887);
nand U15962 (N_15962,N_14774,N_14870);
nor U15963 (N_15963,N_14332,N_14242);
or U15964 (N_15964,N_14308,N_14362);
xnor U15965 (N_15965,N_14951,N_14957);
nand U15966 (N_15966,N_14542,N_14685);
or U15967 (N_15967,N_14990,N_14699);
and U15968 (N_15968,N_14958,N_14657);
nand U15969 (N_15969,N_14271,N_14207);
and U15970 (N_15970,N_14344,N_14782);
and U15971 (N_15971,N_14713,N_14454);
nor U15972 (N_15972,N_14407,N_14587);
xnor U15973 (N_15973,N_14509,N_14799);
nor U15974 (N_15974,N_14853,N_14085);
nand U15975 (N_15975,N_14884,N_14130);
nand U15976 (N_15976,N_14955,N_14315);
nand U15977 (N_15977,N_14717,N_14667);
and U15978 (N_15978,N_14062,N_14893);
and U15979 (N_15979,N_14758,N_14676);
nor U15980 (N_15980,N_14213,N_14555);
nand U15981 (N_15981,N_14425,N_14013);
xor U15982 (N_15982,N_14030,N_14676);
nand U15983 (N_15983,N_14337,N_14935);
and U15984 (N_15984,N_14512,N_14566);
nor U15985 (N_15985,N_14079,N_14581);
xnor U15986 (N_15986,N_14968,N_14374);
nand U15987 (N_15987,N_14747,N_14427);
or U15988 (N_15988,N_14930,N_14860);
or U15989 (N_15989,N_14852,N_14094);
xnor U15990 (N_15990,N_14537,N_14644);
xor U15991 (N_15991,N_14484,N_14826);
nor U15992 (N_15992,N_14529,N_14133);
nand U15993 (N_15993,N_14372,N_14082);
and U15994 (N_15994,N_14096,N_14882);
nand U15995 (N_15995,N_14763,N_14091);
nor U15996 (N_15996,N_14556,N_14781);
and U15997 (N_15997,N_14217,N_14461);
or U15998 (N_15998,N_14508,N_14831);
xor U15999 (N_15999,N_14521,N_14850);
nor U16000 (N_16000,N_15539,N_15490);
and U16001 (N_16001,N_15352,N_15933);
or U16002 (N_16002,N_15750,N_15835);
nor U16003 (N_16003,N_15924,N_15288);
nor U16004 (N_16004,N_15322,N_15422);
or U16005 (N_16005,N_15391,N_15110);
xnor U16006 (N_16006,N_15012,N_15002);
and U16007 (N_16007,N_15788,N_15133);
nand U16008 (N_16008,N_15158,N_15244);
nand U16009 (N_16009,N_15725,N_15084);
and U16010 (N_16010,N_15390,N_15282);
or U16011 (N_16011,N_15602,N_15846);
and U16012 (N_16012,N_15532,N_15299);
nor U16013 (N_16013,N_15603,N_15050);
nand U16014 (N_16014,N_15239,N_15544);
nand U16015 (N_16015,N_15384,N_15693);
nor U16016 (N_16016,N_15307,N_15097);
or U16017 (N_16017,N_15087,N_15464);
xnor U16018 (N_16018,N_15626,N_15219);
or U16019 (N_16019,N_15722,N_15120);
xor U16020 (N_16020,N_15954,N_15781);
nor U16021 (N_16021,N_15971,N_15191);
and U16022 (N_16022,N_15396,N_15445);
nand U16023 (N_16023,N_15981,N_15362);
or U16024 (N_16024,N_15421,N_15301);
nand U16025 (N_16025,N_15053,N_15991);
nand U16026 (N_16026,N_15508,N_15964);
nand U16027 (N_16027,N_15775,N_15952);
xnor U16028 (N_16028,N_15766,N_15751);
nand U16029 (N_16029,N_15435,N_15517);
xor U16030 (N_16030,N_15795,N_15556);
nor U16031 (N_16031,N_15811,N_15724);
or U16032 (N_16032,N_15709,N_15470);
or U16033 (N_16033,N_15814,N_15297);
and U16034 (N_16034,N_15455,N_15542);
xor U16035 (N_16035,N_15618,N_15161);
nand U16036 (N_16036,N_15142,N_15504);
nor U16037 (N_16037,N_15871,N_15430);
nand U16038 (N_16038,N_15173,N_15137);
or U16039 (N_16039,N_15222,N_15912);
xor U16040 (N_16040,N_15653,N_15529);
nor U16041 (N_16041,N_15836,N_15278);
or U16042 (N_16042,N_15999,N_15507);
or U16043 (N_16043,N_15458,N_15369);
nor U16044 (N_16044,N_15957,N_15048);
or U16045 (N_16045,N_15174,N_15342);
nor U16046 (N_16046,N_15355,N_15807);
nor U16047 (N_16047,N_15292,N_15522);
nor U16048 (N_16048,N_15885,N_15404);
or U16049 (N_16049,N_15230,N_15155);
nand U16050 (N_16050,N_15509,N_15568);
nor U16051 (N_16051,N_15613,N_15157);
or U16052 (N_16052,N_15334,N_15953);
nor U16053 (N_16053,N_15250,N_15176);
nor U16054 (N_16054,N_15630,N_15406);
and U16055 (N_16055,N_15393,N_15280);
or U16056 (N_16056,N_15909,N_15545);
nor U16057 (N_16057,N_15148,N_15798);
and U16058 (N_16058,N_15864,N_15837);
nand U16059 (N_16059,N_15546,N_15644);
nand U16060 (N_16060,N_15842,N_15690);
and U16061 (N_16061,N_15293,N_15913);
nand U16062 (N_16062,N_15030,N_15415);
and U16063 (N_16063,N_15571,N_15428);
nand U16064 (N_16064,N_15303,N_15052);
nor U16065 (N_16065,N_15730,N_15866);
and U16066 (N_16066,N_15881,N_15160);
xor U16067 (N_16067,N_15732,N_15294);
nor U16068 (N_16068,N_15236,N_15525);
and U16069 (N_16069,N_15793,N_15605);
xnor U16070 (N_16070,N_15419,N_15289);
xnor U16071 (N_16071,N_15462,N_15001);
or U16072 (N_16072,N_15733,N_15381);
or U16073 (N_16073,N_15092,N_15668);
and U16074 (N_16074,N_15809,N_15667);
nand U16075 (N_16075,N_15505,N_15283);
nand U16076 (N_16076,N_15256,N_15312);
nor U16077 (N_16077,N_15385,N_15448);
nand U16078 (N_16078,N_15474,N_15460);
nand U16079 (N_16079,N_15822,N_15102);
nand U16080 (N_16080,N_15295,N_15581);
or U16081 (N_16081,N_15869,N_15310);
nor U16082 (N_16082,N_15285,N_15785);
xnor U16083 (N_16083,N_15072,N_15434);
and U16084 (N_16084,N_15410,N_15948);
nand U16085 (N_16085,N_15198,N_15677);
nor U16086 (N_16086,N_15749,N_15850);
nor U16087 (N_16087,N_15333,N_15485);
xor U16088 (N_16088,N_15899,N_15253);
nand U16089 (N_16089,N_15812,N_15938);
and U16090 (N_16090,N_15714,N_15591);
and U16091 (N_16091,N_15966,N_15477);
xor U16092 (N_16092,N_15992,N_15827);
xnor U16093 (N_16093,N_15166,N_15248);
nor U16094 (N_16094,N_15513,N_15365);
nand U16095 (N_16095,N_15985,N_15551);
xnor U16096 (N_16096,N_15945,N_15338);
and U16097 (N_16097,N_15403,N_15825);
and U16098 (N_16098,N_15627,N_15765);
nor U16099 (N_16099,N_15743,N_15387);
and U16100 (N_16100,N_15042,N_15080);
xnor U16101 (N_16101,N_15298,N_15329);
nand U16102 (N_16102,N_15443,N_15206);
xnor U16103 (N_16103,N_15487,N_15780);
nand U16104 (N_16104,N_15363,N_15008);
or U16105 (N_16105,N_15853,N_15577);
nor U16106 (N_16106,N_15043,N_15302);
nand U16107 (N_16107,N_15115,N_15475);
and U16108 (N_16108,N_15423,N_15398);
nor U16109 (N_16109,N_15291,N_15537);
and U16110 (N_16110,N_15600,N_15438);
nor U16111 (N_16111,N_15351,N_15129);
nor U16112 (N_16112,N_15059,N_15375);
xnor U16113 (N_16113,N_15520,N_15791);
and U16114 (N_16114,N_15274,N_15819);
nand U16115 (N_16115,N_15854,N_15796);
nand U16116 (N_16116,N_15922,N_15740);
xnor U16117 (N_16117,N_15927,N_15208);
or U16118 (N_16118,N_15773,N_15220);
and U16119 (N_16119,N_15657,N_15243);
xor U16120 (N_16120,N_15456,N_15000);
nor U16121 (N_16121,N_15955,N_15397);
nand U16122 (N_16122,N_15823,N_15891);
nand U16123 (N_16123,N_15538,N_15701);
and U16124 (N_16124,N_15856,N_15995);
or U16125 (N_16125,N_15958,N_15950);
or U16126 (N_16126,N_15016,N_15411);
xnor U16127 (N_16127,N_15119,N_15700);
nor U16128 (N_16128,N_15116,N_15859);
nand U16129 (N_16129,N_15200,N_15987);
nor U16130 (N_16130,N_15235,N_15405);
nand U16131 (N_16131,N_15717,N_15139);
nor U16132 (N_16132,N_15134,N_15466);
or U16133 (N_16133,N_15339,N_15370);
nor U16134 (N_16134,N_15154,N_15232);
nand U16135 (N_16135,N_15764,N_15440);
nand U16136 (N_16136,N_15572,N_15639);
and U16137 (N_16137,N_15550,N_15664);
xor U16138 (N_16138,N_15136,N_15045);
nor U16139 (N_16139,N_15805,N_15654);
or U16140 (N_16140,N_15665,N_15800);
nor U16141 (N_16141,N_15547,N_15893);
xnor U16142 (N_16142,N_15360,N_15442);
nand U16143 (N_16143,N_15185,N_15768);
nand U16144 (N_16144,N_15126,N_15608);
nand U16145 (N_16145,N_15020,N_15527);
nor U16146 (N_16146,N_15085,N_15179);
and U16147 (N_16147,N_15450,N_15524);
nand U16148 (N_16148,N_15757,N_15172);
nor U16149 (N_16149,N_15802,N_15531);
xor U16150 (N_16150,N_15907,N_15194);
nor U16151 (N_16151,N_15025,N_15229);
or U16152 (N_16152,N_15576,N_15357);
nand U16153 (N_16153,N_15923,N_15186);
xor U16154 (N_16154,N_15673,N_15554);
xor U16155 (N_16155,N_15794,N_15801);
nor U16156 (N_16156,N_15346,N_15883);
nor U16157 (N_16157,N_15318,N_15311);
or U16158 (N_16158,N_15004,N_15648);
nor U16159 (N_16159,N_15787,N_15106);
and U16160 (N_16160,N_15977,N_15699);
and U16161 (N_16161,N_15890,N_15469);
or U16162 (N_16162,N_15121,N_15252);
or U16163 (N_16163,N_15723,N_15359);
nand U16164 (N_16164,N_15862,N_15275);
xnor U16165 (N_16165,N_15367,N_15988);
nand U16166 (N_16166,N_15942,N_15067);
nand U16167 (N_16167,N_15223,N_15007);
or U16168 (N_16168,N_15672,N_15921);
nand U16169 (N_16169,N_15327,N_15151);
nand U16170 (N_16170,N_15408,N_15305);
xnor U16171 (N_16171,N_15489,N_15127);
xor U16172 (N_16172,N_15804,N_15040);
or U16173 (N_16173,N_15710,N_15467);
xor U16174 (N_16174,N_15395,N_15495);
nand U16175 (N_16175,N_15506,N_15642);
and U16176 (N_16176,N_15887,N_15254);
nor U16177 (N_16177,N_15290,N_15399);
xnor U16178 (N_16178,N_15965,N_15840);
xor U16179 (N_16179,N_15328,N_15939);
or U16180 (N_16180,N_15718,N_15374);
xnor U16181 (N_16181,N_15900,N_15473);
nand U16182 (N_16182,N_15070,N_15931);
and U16183 (N_16183,N_15371,N_15062);
xnor U16184 (N_16184,N_15675,N_15078);
nor U16185 (N_16185,N_15936,N_15727);
and U16186 (N_16186,N_15518,N_15582);
xor U16187 (N_16187,N_15707,N_15615);
xor U16188 (N_16188,N_15184,N_15389);
or U16189 (N_16189,N_15875,N_15880);
nand U16190 (N_16190,N_15857,N_15637);
or U16191 (N_16191,N_15433,N_15548);
nand U16192 (N_16192,N_15534,N_15851);
and U16193 (N_16193,N_15562,N_15103);
nand U16194 (N_16194,N_15093,N_15082);
xor U16195 (N_16195,N_15039,N_15152);
and U16196 (N_16196,N_15073,N_15358);
nand U16197 (N_16197,N_15671,N_15861);
xnor U16198 (N_16198,N_15978,N_15839);
nand U16199 (N_16199,N_15079,N_15108);
nand U16200 (N_16200,N_15790,N_15196);
and U16201 (N_16201,N_15388,N_15011);
nand U16202 (N_16202,N_15557,N_15870);
and U16203 (N_16203,N_15560,N_15238);
or U16204 (N_16204,N_15575,N_15728);
nor U16205 (N_16205,N_15246,N_15153);
nor U16206 (N_16206,N_15920,N_15377);
nor U16207 (N_16207,N_15739,N_15946);
nand U16208 (N_16208,N_15604,N_15492);
xor U16209 (N_16209,N_15058,N_15175);
nor U16210 (N_16210,N_15919,N_15313);
nor U16211 (N_16211,N_15702,N_15563);
xnor U16212 (N_16212,N_15656,N_15017);
nor U16213 (N_16213,N_15241,N_15584);
or U16214 (N_16214,N_15810,N_15258);
nor U16215 (N_16215,N_15972,N_15047);
or U16216 (N_16216,N_15799,N_15098);
and U16217 (N_16217,N_15268,N_15417);
or U16218 (N_16218,N_15321,N_15128);
and U16219 (N_16219,N_15240,N_15138);
xor U16220 (N_16220,N_15808,N_15003);
nor U16221 (N_16221,N_15916,N_15130);
xnor U16222 (N_16222,N_15259,N_15366);
or U16223 (N_16223,N_15197,N_15782);
and U16224 (N_16224,N_15849,N_15831);
or U16225 (N_16225,N_15598,N_15684);
and U16226 (N_16226,N_15704,N_15482);
or U16227 (N_16227,N_15593,N_15659);
or U16228 (N_16228,N_15736,N_15567);
and U16229 (N_16229,N_15331,N_15553);
nor U16230 (N_16230,N_15345,N_15650);
nor U16231 (N_16231,N_15863,N_15638);
and U16232 (N_16232,N_15373,N_15569);
and U16233 (N_16233,N_15692,N_15696);
and U16234 (N_16234,N_15409,N_15735);
nand U16235 (N_16235,N_15033,N_15019);
nor U16236 (N_16236,N_15091,N_15414);
nand U16237 (N_16237,N_15027,N_15655);
nor U16238 (N_16238,N_15868,N_15461);
nor U16239 (N_16239,N_15737,N_15269);
nor U16240 (N_16240,N_15914,N_15156);
xor U16241 (N_16241,N_15484,N_15711);
nor U16242 (N_16242,N_15476,N_15803);
xnor U16243 (N_16243,N_15975,N_15759);
nand U16244 (N_16244,N_15496,N_15993);
and U16245 (N_16245,N_15564,N_15832);
and U16246 (N_16246,N_15956,N_15071);
or U16247 (N_16247,N_15202,N_15036);
nor U16248 (N_16248,N_15347,N_15526);
nand U16249 (N_16249,N_15625,N_15878);
xnor U16250 (N_16250,N_15731,N_15426);
nor U16251 (N_16251,N_15143,N_15969);
xnor U16252 (N_16252,N_15237,N_15523);
nor U16253 (N_16253,N_15465,N_15451);
xnor U16254 (N_16254,N_15159,N_15940);
xor U16255 (N_16255,N_15177,N_15064);
xor U16256 (N_16256,N_15612,N_15021);
nand U16257 (N_16257,N_15123,N_15213);
nor U16258 (N_16258,N_15122,N_15037);
nor U16259 (N_16259,N_15855,N_15828);
and U16260 (N_16260,N_15777,N_15276);
xnor U16261 (N_16261,N_15902,N_15695);
nor U16262 (N_16262,N_15325,N_15976);
nor U16263 (N_16263,N_15316,N_15502);
and U16264 (N_16264,N_15623,N_15095);
nor U16265 (N_16265,N_15480,N_15776);
and U16266 (N_16266,N_15189,N_15918);
nand U16267 (N_16267,N_15145,N_15925);
or U16268 (N_16268,N_15898,N_15592);
xnor U16269 (N_16269,N_15218,N_15066);
xor U16270 (N_16270,N_15658,N_15182);
nand U16271 (N_16271,N_15231,N_15454);
nor U16272 (N_16272,N_15233,N_15867);
and U16273 (N_16273,N_15437,N_15943);
or U16274 (N_16274,N_15439,N_15272);
or U16275 (N_16275,N_15847,N_15214);
and U16276 (N_16276,N_15744,N_15353);
xor U16277 (N_16277,N_15873,N_15447);
nand U16278 (N_16278,N_15183,N_15181);
xor U16279 (N_16279,N_15224,N_15686);
xnor U16280 (N_16280,N_15712,N_15094);
xnor U16281 (N_16281,N_15135,N_15081);
nor U16282 (N_16282,N_15498,N_15510);
xor U16283 (N_16283,N_15418,N_15207);
xnor U16284 (N_16284,N_15949,N_15678);
or U16285 (N_16285,N_15029,N_15028);
or U16286 (N_16286,N_15424,N_15380);
nor U16287 (N_16287,N_15528,N_15874);
xnor U16288 (N_16288,N_15588,N_15729);
and U16289 (N_16289,N_15944,N_15144);
xnor U16290 (N_16290,N_15963,N_15150);
nand U16291 (N_16291,N_15962,N_15107);
or U16292 (N_16292,N_15543,N_15713);
or U16293 (N_16293,N_15821,N_15190);
or U16294 (N_16294,N_15903,N_15643);
or U16295 (N_16295,N_15663,N_15745);
or U16296 (N_16296,N_15472,N_15763);
xnor U16297 (N_16297,N_15124,N_15915);
nand U16298 (N_16298,N_15247,N_15296);
and U16299 (N_16299,N_15892,N_15076);
or U16300 (N_16300,N_15959,N_15356);
and U16301 (N_16301,N_15010,N_15561);
xor U16302 (N_16302,N_15586,N_15193);
nor U16303 (N_16303,N_15227,N_15332);
xor U16304 (N_16304,N_15060,N_15610);
xnor U16305 (N_16305,N_15830,N_15580);
and U16306 (N_16306,N_15726,N_15579);
or U16307 (N_16307,N_15441,N_15647);
and U16308 (N_16308,N_15689,N_15748);
nor U16309 (N_16309,N_15783,N_15676);
nor U16310 (N_16310,N_15640,N_15006);
and U16311 (N_16311,N_15994,N_15789);
nand U16312 (N_16312,N_15277,N_15982);
or U16313 (N_16313,N_15601,N_15973);
xor U16314 (N_16314,N_15270,N_15843);
xnor U16315 (N_16315,N_15265,N_15552);
nand U16316 (N_16316,N_15820,N_15452);
or U16317 (N_16317,N_15649,N_15026);
nor U16318 (N_16318,N_15559,N_15015);
xor U16319 (N_16319,N_15599,N_15530);
xor U16320 (N_16320,N_15343,N_15906);
or U16321 (N_16321,N_15570,N_15077);
and U16322 (N_16322,N_15772,N_15323);
nand U16323 (N_16323,N_15488,N_15698);
nor U16324 (N_16324,N_15034,N_15242);
nand U16325 (N_16325,N_15669,N_15666);
xnor U16326 (N_16326,N_15680,N_15061);
or U16327 (N_16327,N_15187,N_15486);
xor U16328 (N_16328,N_15685,N_15314);
or U16329 (N_16329,N_15951,N_15928);
nand U16330 (N_16330,N_15720,N_15459);
xnor U16331 (N_16331,N_15335,N_15225);
and U16332 (N_16332,N_15035,N_15420);
or U16333 (N_16333,N_15741,N_15209);
nand U16334 (N_16334,N_15217,N_15501);
xor U16335 (N_16335,N_15300,N_15372);
nor U16336 (N_16336,N_15834,N_15974);
or U16337 (N_16337,N_15264,N_15416);
and U16338 (N_16338,N_15281,N_15427);
nand U16339 (N_16339,N_15996,N_15088);
and U16340 (N_16340,N_15149,N_15889);
nor U16341 (N_16341,N_15979,N_15444);
xor U16342 (N_16342,N_15271,N_15606);
or U16343 (N_16343,N_15930,N_15350);
or U16344 (N_16344,N_15304,N_15815);
nand U16345 (N_16345,N_15960,N_15917);
and U16346 (N_16346,N_15540,N_15670);
nand U16347 (N_16347,N_15055,N_15386);
and U16348 (N_16348,N_15090,N_15056);
and U16349 (N_16349,N_15112,N_15014);
nand U16350 (N_16350,N_15023,N_15747);
or U16351 (N_16351,N_15566,N_15590);
xnor U16352 (N_16352,N_15057,N_15049);
or U16353 (N_16353,N_15620,N_15607);
nand U16354 (N_16354,N_15514,N_15989);
xnor U16355 (N_16355,N_15257,N_15413);
nand U16356 (N_16356,N_15833,N_15279);
and U16357 (N_16357,N_15046,N_15929);
nor U16358 (N_16358,N_15986,N_15336);
or U16359 (N_16359,N_15984,N_15205);
nor U16360 (N_16360,N_15816,N_15326);
nand U16361 (N_16361,N_15516,N_15018);
nor U16362 (N_16362,N_15860,N_15267);
nor U16363 (N_16363,N_15641,N_15826);
and U16364 (N_16364,N_15573,N_15457);
and U16365 (N_16365,N_15706,N_15687);
nand U16366 (N_16366,N_15719,N_15210);
and U16367 (N_16367,N_15378,N_15941);
xor U16368 (N_16368,N_15646,N_15549);
nor U16369 (N_16369,N_15431,N_15895);
and U16370 (N_16370,N_15674,N_15075);
xnor U16371 (N_16371,N_15463,N_15478);
or U16372 (N_16372,N_15886,N_15512);
xor U16373 (N_16373,N_15635,N_15721);
nand U16374 (N_16374,N_15611,N_15752);
and U16375 (N_16375,N_15896,N_15118);
nor U16376 (N_16376,N_15125,N_15519);
xor U16377 (N_16377,N_15761,N_15628);
or U16378 (N_16378,N_15146,N_15691);
and U16379 (N_16379,N_15894,N_15215);
or U16380 (N_16380,N_15211,N_15503);
or U16381 (N_16381,N_15734,N_15753);
xor U16382 (N_16382,N_15169,N_15491);
and U16383 (N_16383,N_15340,N_15162);
nand U16384 (N_16384,N_15679,N_15624);
and U16385 (N_16385,N_15032,N_15908);
nand U16386 (N_16386,N_15063,N_15319);
nor U16387 (N_16387,N_15705,N_15756);
xnor U16388 (N_16388,N_15715,N_15471);
and U16389 (N_16389,N_15497,N_15167);
or U16390 (N_16390,N_15779,N_15594);
nand U16391 (N_16391,N_15662,N_15578);
and U16392 (N_16392,N_15521,N_15432);
and U16393 (N_16393,N_15660,N_15212);
nor U16394 (N_16394,N_15368,N_15614);
xnor U16395 (N_16395,N_15054,N_15500);
nor U16396 (N_16396,N_15483,N_15383);
xnor U16397 (N_16397,N_15872,N_15786);
nand U16398 (N_16398,N_15364,N_15738);
xor U16399 (N_16399,N_15105,N_15511);
nand U16400 (N_16400,N_15446,N_15865);
and U16401 (N_16401,N_15682,N_15337);
nor U16402 (N_16402,N_15587,N_15970);
and U16403 (N_16403,N_15897,N_15284);
or U16404 (N_16404,N_15622,N_15767);
nor U16405 (N_16405,N_15361,N_15769);
nor U16406 (N_16406,N_15178,N_15758);
and U16407 (N_16407,N_15251,N_15038);
and U16408 (N_16408,N_15844,N_15838);
xnor U16409 (N_16409,N_15852,N_15317);
xnor U16410 (N_16410,N_15221,N_15904);
nand U16411 (N_16411,N_15065,N_15818);
nand U16412 (N_16412,N_15884,N_15558);
nand U16413 (N_16413,N_15792,N_15934);
xnor U16414 (N_16414,N_15813,N_15742);
nand U16415 (N_16415,N_15652,N_15044);
nand U16416 (N_16416,N_15392,N_15425);
nor U16417 (N_16417,N_15402,N_15968);
and U16418 (N_16418,N_15515,N_15170);
nor U16419 (N_16419,N_15997,N_15774);
or U16420 (N_16420,N_15771,N_15829);
nor U16421 (N_16421,N_15645,N_15905);
and U16422 (N_16422,N_15226,N_15636);
nor U16423 (N_16423,N_15536,N_15681);
or U16424 (N_16424,N_15101,N_15201);
nor U16425 (N_16425,N_15204,N_15703);
nand U16426 (N_16426,N_15041,N_15140);
nand U16427 (N_16427,N_15574,N_15400);
xor U16428 (N_16428,N_15778,N_15770);
nand U16429 (N_16429,N_15541,N_15806);
or U16430 (N_16430,N_15089,N_15262);
and U16431 (N_16431,N_15104,N_15315);
or U16432 (N_16432,N_15165,N_15876);
xor U16433 (N_16433,N_15845,N_15634);
or U16434 (N_16434,N_15882,N_15086);
or U16435 (N_16435,N_15376,N_15468);
and U16436 (N_16436,N_15533,N_15379);
nor U16437 (N_16437,N_15535,N_15910);
xnor U16438 (N_16438,N_15068,N_15113);
xor U16439 (N_16439,N_15195,N_15980);
xor U16440 (N_16440,N_15109,N_15817);
nand U16441 (N_16441,N_15132,N_15407);
or U16442 (N_16442,N_15263,N_15412);
nand U16443 (N_16443,N_15858,N_15341);
nor U16444 (N_16444,N_15697,N_15349);
nand U16445 (N_16445,N_15583,N_15493);
and U16446 (N_16446,N_15286,N_15879);
or U16447 (N_16447,N_15688,N_15354);
xor U16448 (N_16448,N_15616,N_15746);
nand U16449 (N_16449,N_15171,N_15848);
nand U16450 (N_16450,N_15716,N_15249);
xnor U16451 (N_16451,N_15760,N_15022);
or U16452 (N_16452,N_15266,N_15932);
xnor U16453 (N_16453,N_15099,N_15453);
nor U16454 (N_16454,N_15111,N_15141);
xor U16455 (N_16455,N_15382,N_15499);
nor U16456 (N_16456,N_15708,N_15192);
and U16457 (N_16457,N_15287,N_15555);
xor U16458 (N_16458,N_15147,N_15199);
nor U16459 (N_16459,N_15449,N_15117);
and U16460 (N_16460,N_15260,N_15324);
xor U16461 (N_16461,N_15273,N_15005);
xor U16462 (N_16462,N_15306,N_15216);
and U16463 (N_16463,N_15619,N_15937);
nor U16464 (N_16464,N_15083,N_15394);
or U16465 (N_16465,N_15234,N_15100);
and U16466 (N_16466,N_15784,N_15481);
nor U16467 (N_16467,N_15877,N_15330);
or U16468 (N_16468,N_15245,N_15180);
nand U16469 (N_16469,N_15401,N_15990);
xor U16470 (N_16470,N_15755,N_15188);
and U16471 (N_16471,N_15320,N_15596);
and U16472 (N_16472,N_15131,N_15926);
and U16473 (N_16473,N_15585,N_15494);
nor U16474 (N_16474,N_15051,N_15348);
or U16475 (N_16475,N_15911,N_15841);
nor U16476 (N_16476,N_15164,N_15617);
xor U16477 (N_16477,N_15754,N_15255);
nand U16478 (N_16478,N_15013,N_15983);
nand U16479 (N_16479,N_15261,N_15074);
or U16480 (N_16480,N_15203,N_15344);
and U16481 (N_16481,N_15967,N_15597);
nor U16482 (N_16482,N_15947,N_15694);
and U16483 (N_16483,N_15888,N_15308);
nand U16484 (N_16484,N_15629,N_15031);
and U16485 (N_16485,N_15683,N_15096);
xnor U16486 (N_16486,N_15762,N_15633);
nand U16487 (N_16487,N_15069,N_15632);
and U16488 (N_16488,N_15651,N_15595);
nand U16489 (N_16489,N_15998,N_15479);
xor U16490 (N_16490,N_15589,N_15429);
xor U16491 (N_16491,N_15114,N_15661);
or U16492 (N_16492,N_15935,N_15961);
nor U16493 (N_16493,N_15168,N_15228);
nand U16494 (N_16494,N_15609,N_15009);
xor U16495 (N_16495,N_15631,N_15309);
and U16496 (N_16496,N_15565,N_15824);
and U16497 (N_16497,N_15901,N_15024);
nor U16498 (N_16498,N_15621,N_15797);
nand U16499 (N_16499,N_15163,N_15436);
and U16500 (N_16500,N_15143,N_15039);
and U16501 (N_16501,N_15634,N_15282);
nand U16502 (N_16502,N_15069,N_15687);
or U16503 (N_16503,N_15821,N_15739);
nor U16504 (N_16504,N_15683,N_15997);
and U16505 (N_16505,N_15747,N_15726);
xnor U16506 (N_16506,N_15899,N_15390);
nand U16507 (N_16507,N_15873,N_15738);
nor U16508 (N_16508,N_15884,N_15125);
xnor U16509 (N_16509,N_15701,N_15440);
and U16510 (N_16510,N_15145,N_15916);
nor U16511 (N_16511,N_15994,N_15920);
or U16512 (N_16512,N_15064,N_15632);
xnor U16513 (N_16513,N_15876,N_15875);
xnor U16514 (N_16514,N_15401,N_15427);
or U16515 (N_16515,N_15074,N_15091);
nand U16516 (N_16516,N_15819,N_15894);
nand U16517 (N_16517,N_15811,N_15414);
or U16518 (N_16518,N_15370,N_15320);
and U16519 (N_16519,N_15389,N_15703);
and U16520 (N_16520,N_15912,N_15090);
and U16521 (N_16521,N_15604,N_15166);
nand U16522 (N_16522,N_15207,N_15807);
and U16523 (N_16523,N_15004,N_15370);
xnor U16524 (N_16524,N_15285,N_15552);
nor U16525 (N_16525,N_15213,N_15691);
xor U16526 (N_16526,N_15649,N_15899);
nand U16527 (N_16527,N_15033,N_15485);
xor U16528 (N_16528,N_15294,N_15832);
nand U16529 (N_16529,N_15701,N_15109);
nand U16530 (N_16530,N_15865,N_15409);
and U16531 (N_16531,N_15302,N_15128);
and U16532 (N_16532,N_15963,N_15666);
nand U16533 (N_16533,N_15994,N_15841);
nand U16534 (N_16534,N_15873,N_15323);
or U16535 (N_16535,N_15764,N_15846);
or U16536 (N_16536,N_15370,N_15899);
nand U16537 (N_16537,N_15013,N_15978);
or U16538 (N_16538,N_15732,N_15252);
nand U16539 (N_16539,N_15314,N_15690);
xnor U16540 (N_16540,N_15960,N_15942);
or U16541 (N_16541,N_15259,N_15722);
or U16542 (N_16542,N_15519,N_15865);
or U16543 (N_16543,N_15926,N_15920);
nor U16544 (N_16544,N_15450,N_15745);
xnor U16545 (N_16545,N_15755,N_15274);
or U16546 (N_16546,N_15863,N_15218);
or U16547 (N_16547,N_15847,N_15383);
or U16548 (N_16548,N_15715,N_15629);
nand U16549 (N_16549,N_15255,N_15645);
xor U16550 (N_16550,N_15986,N_15749);
nand U16551 (N_16551,N_15879,N_15587);
nor U16552 (N_16552,N_15362,N_15337);
and U16553 (N_16553,N_15619,N_15858);
or U16554 (N_16554,N_15890,N_15694);
nand U16555 (N_16555,N_15075,N_15062);
xor U16556 (N_16556,N_15370,N_15578);
nand U16557 (N_16557,N_15982,N_15161);
xor U16558 (N_16558,N_15149,N_15712);
and U16559 (N_16559,N_15614,N_15055);
nand U16560 (N_16560,N_15233,N_15515);
xor U16561 (N_16561,N_15347,N_15199);
nor U16562 (N_16562,N_15116,N_15557);
xnor U16563 (N_16563,N_15573,N_15490);
or U16564 (N_16564,N_15792,N_15634);
nand U16565 (N_16565,N_15845,N_15679);
xor U16566 (N_16566,N_15336,N_15878);
nand U16567 (N_16567,N_15130,N_15027);
nand U16568 (N_16568,N_15773,N_15102);
xnor U16569 (N_16569,N_15047,N_15306);
nand U16570 (N_16570,N_15154,N_15373);
and U16571 (N_16571,N_15077,N_15317);
or U16572 (N_16572,N_15561,N_15636);
nor U16573 (N_16573,N_15738,N_15084);
and U16574 (N_16574,N_15276,N_15014);
nand U16575 (N_16575,N_15536,N_15538);
nor U16576 (N_16576,N_15568,N_15485);
or U16577 (N_16577,N_15901,N_15503);
or U16578 (N_16578,N_15463,N_15741);
xor U16579 (N_16579,N_15483,N_15858);
or U16580 (N_16580,N_15484,N_15750);
and U16581 (N_16581,N_15073,N_15178);
nand U16582 (N_16582,N_15123,N_15069);
and U16583 (N_16583,N_15061,N_15693);
nor U16584 (N_16584,N_15944,N_15002);
xor U16585 (N_16585,N_15634,N_15386);
and U16586 (N_16586,N_15189,N_15372);
nand U16587 (N_16587,N_15847,N_15072);
nand U16588 (N_16588,N_15436,N_15023);
nor U16589 (N_16589,N_15260,N_15326);
xnor U16590 (N_16590,N_15425,N_15861);
nand U16591 (N_16591,N_15421,N_15006);
nand U16592 (N_16592,N_15735,N_15379);
nor U16593 (N_16593,N_15683,N_15154);
or U16594 (N_16594,N_15643,N_15287);
xor U16595 (N_16595,N_15360,N_15966);
and U16596 (N_16596,N_15944,N_15537);
xor U16597 (N_16597,N_15662,N_15580);
xor U16598 (N_16598,N_15448,N_15629);
nor U16599 (N_16599,N_15808,N_15356);
or U16600 (N_16600,N_15848,N_15421);
xor U16601 (N_16601,N_15956,N_15757);
xnor U16602 (N_16602,N_15323,N_15002);
and U16603 (N_16603,N_15320,N_15405);
nor U16604 (N_16604,N_15959,N_15779);
nor U16605 (N_16605,N_15648,N_15900);
xor U16606 (N_16606,N_15219,N_15865);
nand U16607 (N_16607,N_15415,N_15777);
nor U16608 (N_16608,N_15477,N_15619);
or U16609 (N_16609,N_15320,N_15372);
or U16610 (N_16610,N_15868,N_15455);
xnor U16611 (N_16611,N_15067,N_15005);
and U16612 (N_16612,N_15699,N_15935);
nand U16613 (N_16613,N_15248,N_15028);
nor U16614 (N_16614,N_15880,N_15030);
nor U16615 (N_16615,N_15531,N_15635);
xor U16616 (N_16616,N_15419,N_15933);
nor U16617 (N_16617,N_15377,N_15092);
nor U16618 (N_16618,N_15605,N_15107);
and U16619 (N_16619,N_15555,N_15537);
or U16620 (N_16620,N_15003,N_15466);
nor U16621 (N_16621,N_15062,N_15467);
xnor U16622 (N_16622,N_15043,N_15877);
and U16623 (N_16623,N_15091,N_15523);
nor U16624 (N_16624,N_15627,N_15662);
nor U16625 (N_16625,N_15806,N_15309);
nand U16626 (N_16626,N_15816,N_15519);
nand U16627 (N_16627,N_15420,N_15910);
and U16628 (N_16628,N_15166,N_15305);
nand U16629 (N_16629,N_15127,N_15746);
or U16630 (N_16630,N_15537,N_15523);
or U16631 (N_16631,N_15219,N_15637);
and U16632 (N_16632,N_15943,N_15693);
nand U16633 (N_16633,N_15258,N_15655);
or U16634 (N_16634,N_15323,N_15416);
nand U16635 (N_16635,N_15223,N_15867);
nand U16636 (N_16636,N_15365,N_15460);
nand U16637 (N_16637,N_15339,N_15816);
xor U16638 (N_16638,N_15601,N_15788);
xor U16639 (N_16639,N_15342,N_15240);
nand U16640 (N_16640,N_15206,N_15388);
xnor U16641 (N_16641,N_15355,N_15865);
and U16642 (N_16642,N_15273,N_15368);
nor U16643 (N_16643,N_15632,N_15884);
or U16644 (N_16644,N_15576,N_15555);
nor U16645 (N_16645,N_15734,N_15471);
xnor U16646 (N_16646,N_15019,N_15467);
and U16647 (N_16647,N_15898,N_15313);
xnor U16648 (N_16648,N_15265,N_15589);
or U16649 (N_16649,N_15006,N_15820);
or U16650 (N_16650,N_15728,N_15930);
nor U16651 (N_16651,N_15541,N_15363);
and U16652 (N_16652,N_15723,N_15742);
and U16653 (N_16653,N_15328,N_15055);
nor U16654 (N_16654,N_15647,N_15042);
or U16655 (N_16655,N_15674,N_15498);
or U16656 (N_16656,N_15345,N_15161);
or U16657 (N_16657,N_15517,N_15758);
and U16658 (N_16658,N_15267,N_15355);
and U16659 (N_16659,N_15380,N_15294);
and U16660 (N_16660,N_15069,N_15247);
or U16661 (N_16661,N_15389,N_15367);
nor U16662 (N_16662,N_15771,N_15947);
and U16663 (N_16663,N_15341,N_15232);
nor U16664 (N_16664,N_15495,N_15665);
or U16665 (N_16665,N_15146,N_15715);
or U16666 (N_16666,N_15585,N_15144);
nor U16667 (N_16667,N_15014,N_15456);
nand U16668 (N_16668,N_15068,N_15214);
or U16669 (N_16669,N_15027,N_15475);
nand U16670 (N_16670,N_15070,N_15054);
xnor U16671 (N_16671,N_15126,N_15427);
or U16672 (N_16672,N_15820,N_15037);
or U16673 (N_16673,N_15084,N_15221);
nand U16674 (N_16674,N_15523,N_15777);
nand U16675 (N_16675,N_15895,N_15405);
nand U16676 (N_16676,N_15400,N_15687);
xnor U16677 (N_16677,N_15420,N_15436);
nor U16678 (N_16678,N_15935,N_15870);
nor U16679 (N_16679,N_15208,N_15039);
nand U16680 (N_16680,N_15898,N_15127);
nand U16681 (N_16681,N_15449,N_15480);
and U16682 (N_16682,N_15570,N_15749);
or U16683 (N_16683,N_15267,N_15100);
or U16684 (N_16684,N_15818,N_15546);
or U16685 (N_16685,N_15387,N_15547);
and U16686 (N_16686,N_15947,N_15683);
nor U16687 (N_16687,N_15543,N_15437);
and U16688 (N_16688,N_15258,N_15403);
nand U16689 (N_16689,N_15958,N_15601);
xnor U16690 (N_16690,N_15567,N_15818);
nor U16691 (N_16691,N_15558,N_15616);
xnor U16692 (N_16692,N_15859,N_15509);
nor U16693 (N_16693,N_15268,N_15637);
xnor U16694 (N_16694,N_15396,N_15491);
xnor U16695 (N_16695,N_15999,N_15751);
xnor U16696 (N_16696,N_15296,N_15341);
nor U16697 (N_16697,N_15746,N_15855);
nand U16698 (N_16698,N_15903,N_15769);
xnor U16699 (N_16699,N_15516,N_15314);
nor U16700 (N_16700,N_15033,N_15333);
and U16701 (N_16701,N_15344,N_15087);
nor U16702 (N_16702,N_15941,N_15147);
or U16703 (N_16703,N_15088,N_15886);
and U16704 (N_16704,N_15982,N_15412);
nor U16705 (N_16705,N_15895,N_15939);
and U16706 (N_16706,N_15465,N_15355);
nor U16707 (N_16707,N_15469,N_15963);
nand U16708 (N_16708,N_15657,N_15011);
xnor U16709 (N_16709,N_15771,N_15933);
or U16710 (N_16710,N_15374,N_15506);
nor U16711 (N_16711,N_15473,N_15817);
nor U16712 (N_16712,N_15543,N_15804);
and U16713 (N_16713,N_15104,N_15945);
nand U16714 (N_16714,N_15719,N_15526);
or U16715 (N_16715,N_15839,N_15647);
or U16716 (N_16716,N_15269,N_15248);
xor U16717 (N_16717,N_15682,N_15417);
xnor U16718 (N_16718,N_15522,N_15089);
or U16719 (N_16719,N_15520,N_15410);
nand U16720 (N_16720,N_15893,N_15717);
or U16721 (N_16721,N_15067,N_15023);
xnor U16722 (N_16722,N_15170,N_15913);
nor U16723 (N_16723,N_15159,N_15721);
nor U16724 (N_16724,N_15673,N_15564);
nor U16725 (N_16725,N_15528,N_15936);
xor U16726 (N_16726,N_15474,N_15362);
nand U16727 (N_16727,N_15145,N_15353);
nand U16728 (N_16728,N_15541,N_15356);
and U16729 (N_16729,N_15555,N_15029);
nor U16730 (N_16730,N_15075,N_15833);
nand U16731 (N_16731,N_15196,N_15366);
or U16732 (N_16732,N_15398,N_15318);
nor U16733 (N_16733,N_15926,N_15315);
and U16734 (N_16734,N_15187,N_15976);
or U16735 (N_16735,N_15145,N_15151);
nor U16736 (N_16736,N_15687,N_15218);
nand U16737 (N_16737,N_15953,N_15722);
or U16738 (N_16738,N_15808,N_15918);
and U16739 (N_16739,N_15931,N_15027);
xor U16740 (N_16740,N_15974,N_15153);
and U16741 (N_16741,N_15974,N_15370);
nand U16742 (N_16742,N_15231,N_15899);
xor U16743 (N_16743,N_15084,N_15657);
and U16744 (N_16744,N_15999,N_15001);
xor U16745 (N_16745,N_15844,N_15786);
nor U16746 (N_16746,N_15014,N_15798);
nor U16747 (N_16747,N_15846,N_15683);
or U16748 (N_16748,N_15761,N_15137);
or U16749 (N_16749,N_15882,N_15476);
xnor U16750 (N_16750,N_15061,N_15181);
xor U16751 (N_16751,N_15279,N_15432);
or U16752 (N_16752,N_15334,N_15274);
nor U16753 (N_16753,N_15200,N_15880);
nor U16754 (N_16754,N_15727,N_15065);
xor U16755 (N_16755,N_15853,N_15325);
and U16756 (N_16756,N_15678,N_15815);
or U16757 (N_16757,N_15365,N_15473);
nand U16758 (N_16758,N_15864,N_15873);
xnor U16759 (N_16759,N_15761,N_15842);
nand U16760 (N_16760,N_15446,N_15470);
nor U16761 (N_16761,N_15489,N_15417);
and U16762 (N_16762,N_15525,N_15110);
or U16763 (N_16763,N_15321,N_15030);
xor U16764 (N_16764,N_15194,N_15586);
and U16765 (N_16765,N_15892,N_15878);
nor U16766 (N_16766,N_15146,N_15421);
nand U16767 (N_16767,N_15020,N_15472);
xor U16768 (N_16768,N_15934,N_15878);
nor U16769 (N_16769,N_15750,N_15139);
or U16770 (N_16770,N_15393,N_15495);
nand U16771 (N_16771,N_15684,N_15214);
xnor U16772 (N_16772,N_15108,N_15759);
xor U16773 (N_16773,N_15022,N_15051);
nor U16774 (N_16774,N_15879,N_15557);
nand U16775 (N_16775,N_15653,N_15329);
nor U16776 (N_16776,N_15470,N_15204);
nand U16777 (N_16777,N_15810,N_15457);
or U16778 (N_16778,N_15408,N_15160);
nand U16779 (N_16779,N_15382,N_15432);
nor U16780 (N_16780,N_15778,N_15769);
xor U16781 (N_16781,N_15292,N_15779);
nand U16782 (N_16782,N_15427,N_15963);
xnor U16783 (N_16783,N_15513,N_15113);
xor U16784 (N_16784,N_15101,N_15707);
nor U16785 (N_16785,N_15578,N_15311);
xnor U16786 (N_16786,N_15172,N_15687);
or U16787 (N_16787,N_15556,N_15659);
xnor U16788 (N_16788,N_15801,N_15760);
nor U16789 (N_16789,N_15084,N_15369);
nand U16790 (N_16790,N_15306,N_15415);
nor U16791 (N_16791,N_15448,N_15790);
nand U16792 (N_16792,N_15044,N_15346);
nand U16793 (N_16793,N_15371,N_15807);
and U16794 (N_16794,N_15039,N_15696);
and U16795 (N_16795,N_15998,N_15262);
nand U16796 (N_16796,N_15616,N_15045);
or U16797 (N_16797,N_15866,N_15207);
nor U16798 (N_16798,N_15158,N_15528);
and U16799 (N_16799,N_15412,N_15543);
xnor U16800 (N_16800,N_15737,N_15218);
nor U16801 (N_16801,N_15214,N_15626);
and U16802 (N_16802,N_15601,N_15725);
or U16803 (N_16803,N_15200,N_15211);
or U16804 (N_16804,N_15741,N_15516);
and U16805 (N_16805,N_15052,N_15057);
xor U16806 (N_16806,N_15746,N_15729);
and U16807 (N_16807,N_15665,N_15473);
and U16808 (N_16808,N_15538,N_15731);
or U16809 (N_16809,N_15496,N_15670);
and U16810 (N_16810,N_15474,N_15136);
or U16811 (N_16811,N_15294,N_15938);
nand U16812 (N_16812,N_15827,N_15181);
nor U16813 (N_16813,N_15537,N_15481);
and U16814 (N_16814,N_15099,N_15444);
xnor U16815 (N_16815,N_15535,N_15197);
nand U16816 (N_16816,N_15733,N_15345);
or U16817 (N_16817,N_15823,N_15454);
nand U16818 (N_16818,N_15797,N_15617);
and U16819 (N_16819,N_15256,N_15461);
nor U16820 (N_16820,N_15155,N_15705);
or U16821 (N_16821,N_15659,N_15714);
or U16822 (N_16822,N_15903,N_15263);
nand U16823 (N_16823,N_15559,N_15487);
xor U16824 (N_16824,N_15623,N_15965);
and U16825 (N_16825,N_15720,N_15328);
or U16826 (N_16826,N_15739,N_15830);
nand U16827 (N_16827,N_15465,N_15854);
and U16828 (N_16828,N_15268,N_15271);
nor U16829 (N_16829,N_15797,N_15721);
nand U16830 (N_16830,N_15138,N_15137);
or U16831 (N_16831,N_15791,N_15589);
or U16832 (N_16832,N_15455,N_15508);
and U16833 (N_16833,N_15720,N_15994);
and U16834 (N_16834,N_15233,N_15502);
nand U16835 (N_16835,N_15133,N_15684);
nand U16836 (N_16836,N_15389,N_15602);
nand U16837 (N_16837,N_15992,N_15777);
nand U16838 (N_16838,N_15392,N_15072);
and U16839 (N_16839,N_15213,N_15161);
or U16840 (N_16840,N_15950,N_15754);
xor U16841 (N_16841,N_15047,N_15950);
nand U16842 (N_16842,N_15941,N_15140);
nor U16843 (N_16843,N_15415,N_15311);
xor U16844 (N_16844,N_15938,N_15132);
nor U16845 (N_16845,N_15823,N_15540);
nor U16846 (N_16846,N_15402,N_15759);
or U16847 (N_16847,N_15324,N_15115);
or U16848 (N_16848,N_15353,N_15520);
nand U16849 (N_16849,N_15840,N_15530);
nand U16850 (N_16850,N_15704,N_15823);
or U16851 (N_16851,N_15556,N_15840);
and U16852 (N_16852,N_15477,N_15351);
xor U16853 (N_16853,N_15988,N_15173);
or U16854 (N_16854,N_15190,N_15913);
nor U16855 (N_16855,N_15306,N_15282);
and U16856 (N_16856,N_15333,N_15794);
nor U16857 (N_16857,N_15864,N_15340);
or U16858 (N_16858,N_15143,N_15434);
xor U16859 (N_16859,N_15431,N_15706);
nor U16860 (N_16860,N_15954,N_15629);
and U16861 (N_16861,N_15603,N_15735);
nor U16862 (N_16862,N_15848,N_15096);
nor U16863 (N_16863,N_15034,N_15562);
nor U16864 (N_16864,N_15635,N_15361);
and U16865 (N_16865,N_15317,N_15430);
nor U16866 (N_16866,N_15523,N_15283);
nor U16867 (N_16867,N_15731,N_15383);
and U16868 (N_16868,N_15379,N_15275);
nor U16869 (N_16869,N_15121,N_15669);
nand U16870 (N_16870,N_15981,N_15820);
and U16871 (N_16871,N_15528,N_15018);
nor U16872 (N_16872,N_15292,N_15529);
nor U16873 (N_16873,N_15521,N_15355);
or U16874 (N_16874,N_15797,N_15033);
or U16875 (N_16875,N_15543,N_15333);
and U16876 (N_16876,N_15818,N_15109);
nor U16877 (N_16877,N_15475,N_15584);
nand U16878 (N_16878,N_15946,N_15799);
nand U16879 (N_16879,N_15869,N_15345);
and U16880 (N_16880,N_15879,N_15505);
nand U16881 (N_16881,N_15975,N_15971);
nor U16882 (N_16882,N_15952,N_15850);
nand U16883 (N_16883,N_15382,N_15937);
or U16884 (N_16884,N_15625,N_15419);
nor U16885 (N_16885,N_15189,N_15766);
nor U16886 (N_16886,N_15774,N_15190);
and U16887 (N_16887,N_15630,N_15466);
and U16888 (N_16888,N_15263,N_15855);
and U16889 (N_16889,N_15289,N_15532);
nand U16890 (N_16890,N_15381,N_15268);
nand U16891 (N_16891,N_15233,N_15588);
and U16892 (N_16892,N_15740,N_15421);
xnor U16893 (N_16893,N_15135,N_15491);
nand U16894 (N_16894,N_15962,N_15900);
nand U16895 (N_16895,N_15349,N_15617);
xor U16896 (N_16896,N_15015,N_15436);
nand U16897 (N_16897,N_15320,N_15285);
and U16898 (N_16898,N_15120,N_15190);
nor U16899 (N_16899,N_15125,N_15411);
xnor U16900 (N_16900,N_15336,N_15531);
xnor U16901 (N_16901,N_15780,N_15889);
or U16902 (N_16902,N_15139,N_15989);
xor U16903 (N_16903,N_15685,N_15013);
and U16904 (N_16904,N_15765,N_15205);
xnor U16905 (N_16905,N_15100,N_15068);
xnor U16906 (N_16906,N_15890,N_15415);
nand U16907 (N_16907,N_15956,N_15931);
nor U16908 (N_16908,N_15728,N_15276);
and U16909 (N_16909,N_15070,N_15902);
and U16910 (N_16910,N_15406,N_15056);
xnor U16911 (N_16911,N_15383,N_15764);
nand U16912 (N_16912,N_15765,N_15385);
and U16913 (N_16913,N_15528,N_15952);
and U16914 (N_16914,N_15621,N_15184);
or U16915 (N_16915,N_15244,N_15303);
and U16916 (N_16916,N_15966,N_15733);
nand U16917 (N_16917,N_15577,N_15786);
and U16918 (N_16918,N_15861,N_15980);
nand U16919 (N_16919,N_15838,N_15736);
or U16920 (N_16920,N_15835,N_15211);
and U16921 (N_16921,N_15601,N_15520);
nand U16922 (N_16922,N_15647,N_15421);
and U16923 (N_16923,N_15861,N_15385);
or U16924 (N_16924,N_15251,N_15704);
xnor U16925 (N_16925,N_15503,N_15181);
nand U16926 (N_16926,N_15120,N_15313);
nor U16927 (N_16927,N_15993,N_15336);
nor U16928 (N_16928,N_15797,N_15436);
xnor U16929 (N_16929,N_15479,N_15748);
and U16930 (N_16930,N_15930,N_15909);
xnor U16931 (N_16931,N_15522,N_15392);
and U16932 (N_16932,N_15667,N_15959);
xnor U16933 (N_16933,N_15413,N_15554);
nand U16934 (N_16934,N_15346,N_15791);
nand U16935 (N_16935,N_15781,N_15283);
and U16936 (N_16936,N_15583,N_15582);
nand U16937 (N_16937,N_15875,N_15897);
and U16938 (N_16938,N_15222,N_15434);
nand U16939 (N_16939,N_15469,N_15312);
or U16940 (N_16940,N_15019,N_15330);
nand U16941 (N_16941,N_15416,N_15063);
nand U16942 (N_16942,N_15092,N_15541);
and U16943 (N_16943,N_15550,N_15843);
nand U16944 (N_16944,N_15665,N_15515);
and U16945 (N_16945,N_15889,N_15221);
and U16946 (N_16946,N_15029,N_15653);
nor U16947 (N_16947,N_15125,N_15346);
nor U16948 (N_16948,N_15102,N_15728);
and U16949 (N_16949,N_15794,N_15444);
nor U16950 (N_16950,N_15457,N_15536);
and U16951 (N_16951,N_15977,N_15043);
xor U16952 (N_16952,N_15925,N_15399);
and U16953 (N_16953,N_15473,N_15899);
or U16954 (N_16954,N_15554,N_15119);
and U16955 (N_16955,N_15991,N_15584);
xnor U16956 (N_16956,N_15267,N_15081);
nand U16957 (N_16957,N_15551,N_15308);
xnor U16958 (N_16958,N_15233,N_15582);
nor U16959 (N_16959,N_15110,N_15505);
and U16960 (N_16960,N_15613,N_15438);
nor U16961 (N_16961,N_15700,N_15972);
nand U16962 (N_16962,N_15206,N_15151);
nor U16963 (N_16963,N_15212,N_15735);
nand U16964 (N_16964,N_15936,N_15345);
xor U16965 (N_16965,N_15011,N_15709);
xor U16966 (N_16966,N_15925,N_15559);
nor U16967 (N_16967,N_15614,N_15680);
nand U16968 (N_16968,N_15155,N_15709);
nand U16969 (N_16969,N_15282,N_15663);
and U16970 (N_16970,N_15143,N_15758);
nand U16971 (N_16971,N_15421,N_15794);
xor U16972 (N_16972,N_15652,N_15386);
and U16973 (N_16973,N_15683,N_15640);
xor U16974 (N_16974,N_15698,N_15665);
nor U16975 (N_16975,N_15239,N_15382);
nor U16976 (N_16976,N_15036,N_15421);
or U16977 (N_16977,N_15345,N_15105);
nand U16978 (N_16978,N_15954,N_15912);
nand U16979 (N_16979,N_15038,N_15758);
and U16980 (N_16980,N_15017,N_15039);
xnor U16981 (N_16981,N_15370,N_15880);
or U16982 (N_16982,N_15638,N_15201);
or U16983 (N_16983,N_15664,N_15975);
or U16984 (N_16984,N_15322,N_15456);
nor U16985 (N_16985,N_15610,N_15178);
nor U16986 (N_16986,N_15931,N_15013);
and U16987 (N_16987,N_15930,N_15221);
or U16988 (N_16988,N_15292,N_15830);
and U16989 (N_16989,N_15237,N_15419);
nor U16990 (N_16990,N_15160,N_15936);
or U16991 (N_16991,N_15439,N_15840);
nor U16992 (N_16992,N_15826,N_15136);
and U16993 (N_16993,N_15429,N_15293);
nor U16994 (N_16994,N_15020,N_15321);
and U16995 (N_16995,N_15708,N_15089);
or U16996 (N_16996,N_15002,N_15893);
nor U16997 (N_16997,N_15294,N_15217);
and U16998 (N_16998,N_15094,N_15102);
nand U16999 (N_16999,N_15750,N_15978);
nand U17000 (N_17000,N_16231,N_16248);
xor U17001 (N_17001,N_16925,N_16139);
and U17002 (N_17002,N_16195,N_16209);
xnor U17003 (N_17003,N_16520,N_16972);
or U17004 (N_17004,N_16136,N_16971);
nor U17005 (N_17005,N_16626,N_16164);
xor U17006 (N_17006,N_16372,N_16780);
and U17007 (N_17007,N_16947,N_16535);
nand U17008 (N_17008,N_16783,N_16640);
nand U17009 (N_17009,N_16381,N_16038);
or U17010 (N_17010,N_16361,N_16552);
nand U17011 (N_17011,N_16108,N_16496);
nand U17012 (N_17012,N_16879,N_16923);
xor U17013 (N_17013,N_16308,N_16194);
xor U17014 (N_17014,N_16881,N_16781);
xor U17015 (N_17015,N_16866,N_16823);
xor U17016 (N_17016,N_16675,N_16031);
or U17017 (N_17017,N_16206,N_16886);
and U17018 (N_17018,N_16294,N_16803);
xnor U17019 (N_17019,N_16794,N_16912);
nand U17020 (N_17020,N_16313,N_16908);
or U17021 (N_17021,N_16926,N_16698);
xor U17022 (N_17022,N_16754,N_16157);
xor U17023 (N_17023,N_16325,N_16272);
nand U17024 (N_17024,N_16216,N_16589);
nand U17025 (N_17025,N_16184,N_16207);
xor U17026 (N_17026,N_16402,N_16688);
and U17027 (N_17027,N_16077,N_16270);
or U17028 (N_17028,N_16760,N_16735);
xnor U17029 (N_17029,N_16861,N_16653);
xor U17030 (N_17030,N_16828,N_16942);
and U17031 (N_17031,N_16582,N_16906);
or U17032 (N_17032,N_16138,N_16648);
and U17033 (N_17033,N_16793,N_16562);
nand U17034 (N_17034,N_16696,N_16091);
xnor U17035 (N_17035,N_16235,N_16302);
and U17036 (N_17036,N_16468,N_16197);
and U17037 (N_17037,N_16320,N_16305);
xnor U17038 (N_17038,N_16901,N_16475);
xor U17039 (N_17039,N_16343,N_16175);
and U17040 (N_17040,N_16799,N_16674);
or U17041 (N_17041,N_16182,N_16769);
xnor U17042 (N_17042,N_16763,N_16960);
xnor U17043 (N_17043,N_16580,N_16782);
or U17044 (N_17044,N_16183,N_16765);
xnor U17045 (N_17045,N_16287,N_16795);
xor U17046 (N_17046,N_16465,N_16717);
nor U17047 (N_17047,N_16524,N_16009);
or U17048 (N_17048,N_16187,N_16286);
or U17049 (N_17049,N_16643,N_16303);
or U17050 (N_17050,N_16497,N_16340);
nor U17051 (N_17051,N_16113,N_16899);
xor U17052 (N_17052,N_16099,N_16507);
xor U17053 (N_17053,N_16579,N_16721);
or U17054 (N_17054,N_16893,N_16008);
xor U17055 (N_17055,N_16957,N_16629);
nor U17056 (N_17056,N_16444,N_16853);
xor U17057 (N_17057,N_16602,N_16642);
and U17058 (N_17058,N_16217,N_16658);
nor U17059 (N_17059,N_16169,N_16262);
or U17060 (N_17060,N_16620,N_16723);
nor U17061 (N_17061,N_16924,N_16992);
or U17062 (N_17062,N_16558,N_16669);
or U17063 (N_17063,N_16436,N_16953);
nor U17064 (N_17064,N_16985,N_16454);
nand U17065 (N_17065,N_16508,N_16610);
nand U17066 (N_17066,N_16239,N_16132);
xor U17067 (N_17067,N_16536,N_16479);
and U17068 (N_17068,N_16291,N_16137);
nand U17069 (N_17069,N_16776,N_16938);
or U17070 (N_17070,N_16153,N_16577);
nand U17071 (N_17071,N_16115,N_16488);
nand U17072 (N_17072,N_16683,N_16612);
nand U17073 (N_17073,N_16718,N_16598);
xnor U17074 (N_17074,N_16800,N_16847);
nand U17075 (N_17075,N_16198,N_16822);
and U17076 (N_17076,N_16680,N_16775);
and U17077 (N_17077,N_16254,N_16814);
or U17078 (N_17078,N_16788,N_16097);
nand U17079 (N_17079,N_16990,N_16421);
nand U17080 (N_17080,N_16652,N_16709);
and U17081 (N_17081,N_16314,N_16878);
nor U17082 (N_17082,N_16135,N_16029);
nand U17083 (N_17083,N_16103,N_16647);
or U17084 (N_17084,N_16043,N_16007);
or U17085 (N_17085,N_16489,N_16345);
nor U17086 (N_17086,N_16427,N_16979);
nor U17087 (N_17087,N_16720,N_16913);
or U17088 (N_17088,N_16109,N_16351);
nor U17089 (N_17089,N_16613,N_16080);
and U17090 (N_17090,N_16839,N_16362);
nand U17091 (N_17091,N_16311,N_16166);
and U17092 (N_17092,N_16958,N_16155);
or U17093 (N_17093,N_16202,N_16831);
and U17094 (N_17094,N_16257,N_16641);
or U17095 (N_17095,N_16731,N_16020);
nor U17096 (N_17096,N_16252,N_16162);
nand U17097 (N_17097,N_16596,N_16423);
xnor U17098 (N_17098,N_16172,N_16672);
and U17099 (N_17099,N_16935,N_16900);
and U17100 (N_17100,N_16862,N_16838);
nand U17101 (N_17101,N_16621,N_16040);
and U17102 (N_17102,N_16693,N_16310);
nor U17103 (N_17103,N_16846,N_16048);
or U17104 (N_17104,N_16517,N_16944);
or U17105 (N_17105,N_16107,N_16370);
or U17106 (N_17106,N_16770,N_16758);
nor U17107 (N_17107,N_16282,N_16650);
or U17108 (N_17108,N_16296,N_16028);
xor U17109 (N_17109,N_16073,N_16392);
and U17110 (N_17110,N_16140,N_16388);
xor U17111 (N_17111,N_16976,N_16707);
nand U17112 (N_17112,N_16821,N_16512);
or U17113 (N_17113,N_16564,N_16358);
and U17114 (N_17114,N_16975,N_16263);
nor U17115 (N_17115,N_16882,N_16895);
nand U17116 (N_17116,N_16826,N_16404);
or U17117 (N_17117,N_16159,N_16845);
nor U17118 (N_17118,N_16591,N_16323);
xor U17119 (N_17119,N_16446,N_16335);
and U17120 (N_17120,N_16870,N_16661);
xor U17121 (N_17121,N_16978,N_16954);
nand U17122 (N_17122,N_16529,N_16459);
or U17123 (N_17123,N_16412,N_16685);
xnor U17124 (N_17124,N_16074,N_16911);
nor U17125 (N_17125,N_16749,N_16490);
or U17126 (N_17126,N_16950,N_16111);
and U17127 (N_17127,N_16784,N_16887);
nand U17128 (N_17128,N_16060,N_16728);
xnor U17129 (N_17129,N_16003,N_16330);
or U17130 (N_17130,N_16785,N_16738);
and U17131 (N_17131,N_16393,N_16018);
xor U17132 (N_17132,N_16716,N_16830);
xnor U17133 (N_17133,N_16319,N_16247);
nor U17134 (N_17134,N_16275,N_16176);
xor U17135 (N_17135,N_16486,N_16934);
xor U17136 (N_17136,N_16762,N_16443);
xor U17137 (N_17137,N_16811,N_16245);
nand U17138 (N_17138,N_16120,N_16767);
nand U17139 (N_17139,N_16185,N_16131);
xnor U17140 (N_17140,N_16530,N_16289);
or U17141 (N_17141,N_16416,N_16122);
nor U17142 (N_17142,N_16356,N_16952);
or U17143 (N_17143,N_16228,N_16857);
or U17144 (N_17144,N_16092,N_16143);
nor U17145 (N_17145,N_16342,N_16125);
nor U17146 (N_17146,N_16051,N_16012);
or U17147 (N_17147,N_16449,N_16067);
xor U17148 (N_17148,N_16951,N_16898);
and U17149 (N_17149,N_16116,N_16736);
xor U17150 (N_17150,N_16128,N_16970);
xor U17151 (N_17151,N_16929,N_16548);
nor U17152 (N_17152,N_16883,N_16428);
or U17153 (N_17153,N_16452,N_16057);
nor U17154 (N_17154,N_16922,N_16079);
xor U17155 (N_17155,N_16405,N_16902);
nor U17156 (N_17156,N_16329,N_16001);
nand U17157 (N_17157,N_16331,N_16075);
or U17158 (N_17158,N_16606,N_16982);
and U17159 (N_17159,N_16400,N_16130);
and U17160 (N_17160,N_16438,N_16044);
nor U17161 (N_17161,N_16391,N_16690);
nand U17162 (N_17162,N_16165,N_16715);
nor U17163 (N_17163,N_16743,N_16750);
xor U17164 (N_17164,N_16730,N_16588);
or U17165 (N_17165,N_16142,N_16694);
nor U17166 (N_17166,N_16434,N_16484);
nor U17167 (N_17167,N_16849,N_16890);
or U17168 (N_17168,N_16095,N_16081);
and U17169 (N_17169,N_16387,N_16016);
and U17170 (N_17170,N_16431,N_16493);
or U17171 (N_17171,N_16868,N_16915);
xor U17172 (N_17172,N_16295,N_16625);
nand U17173 (N_17173,N_16203,N_16819);
xor U17174 (N_17174,N_16677,N_16071);
xor U17175 (N_17175,N_16753,N_16632);
nor U17176 (N_17176,N_16991,N_16789);
nand U17177 (N_17177,N_16355,N_16191);
xnor U17178 (N_17178,N_16920,N_16981);
or U17179 (N_17179,N_16733,N_16267);
or U17180 (N_17180,N_16027,N_16312);
nand U17181 (N_17181,N_16943,N_16396);
nor U17182 (N_17182,N_16554,N_16858);
xnor U17183 (N_17183,N_16301,N_16875);
nor U17184 (N_17184,N_16534,N_16059);
or U17185 (N_17185,N_16751,N_16907);
and U17186 (N_17186,N_16583,N_16537);
xor U17187 (N_17187,N_16021,N_16367);
or U17188 (N_17188,N_16514,N_16492);
nand U17189 (N_17189,N_16528,N_16840);
or U17190 (N_17190,N_16742,N_16386);
or U17191 (N_17191,N_16983,N_16773);
or U17192 (N_17192,N_16959,N_16557);
nor U17193 (N_17193,N_16725,N_16719);
xor U17194 (N_17194,N_16212,N_16590);
and U17195 (N_17195,N_16076,N_16933);
nor U17196 (N_17196,N_16581,N_16098);
nand U17197 (N_17197,N_16965,N_16987);
nand U17198 (N_17198,N_16570,N_16699);
and U17199 (N_17199,N_16605,N_16631);
xnor U17200 (N_17200,N_16413,N_16124);
nor U17201 (N_17201,N_16424,N_16279);
and U17202 (N_17202,N_16984,N_16339);
and U17203 (N_17203,N_16186,N_16377);
and U17204 (N_17204,N_16792,N_16595);
nor U17205 (N_17205,N_16039,N_16461);
nand U17206 (N_17206,N_16764,N_16365);
and U17207 (N_17207,N_16927,N_16518);
xnor U17208 (N_17208,N_16790,N_16394);
and U17209 (N_17209,N_16101,N_16315);
nand U17210 (N_17210,N_16084,N_16961);
and U17211 (N_17211,N_16201,N_16168);
nand U17212 (N_17212,N_16258,N_16255);
nand U17213 (N_17213,N_16288,N_16772);
nor U17214 (N_17214,N_16498,N_16119);
or U17215 (N_17215,N_16178,N_16664);
or U17216 (N_17216,N_16714,N_16442);
nand U17217 (N_17217,N_16264,N_16072);
nor U17218 (N_17218,N_16324,N_16474);
nand U17219 (N_17219,N_16285,N_16036);
nand U17220 (N_17220,N_16170,N_16724);
xor U17221 (N_17221,N_16877,N_16188);
and U17222 (N_17222,N_16024,N_16274);
and U17223 (N_17223,N_16336,N_16668);
and U17224 (N_17224,N_16466,N_16807);
xnor U17225 (N_17225,N_16271,N_16005);
nand U17226 (N_17226,N_16854,N_16622);
and U17227 (N_17227,N_16578,N_16656);
nor U17228 (N_17228,N_16487,N_16608);
nor U17229 (N_17229,N_16410,N_16181);
nor U17230 (N_17230,N_16786,N_16069);
or U17231 (N_17231,N_16993,N_16727);
or U17232 (N_17232,N_16567,N_16568);
nor U17233 (N_17233,N_16236,N_16757);
or U17234 (N_17234,N_16834,N_16112);
or U17235 (N_17235,N_16682,N_16418);
nor U17236 (N_17236,N_16321,N_16994);
nor U17237 (N_17237,N_16050,N_16237);
xnor U17238 (N_17238,N_16322,N_16090);
nor U17239 (N_17239,N_16948,N_16349);
nand U17240 (N_17240,N_16617,N_16798);
xor U17241 (N_17241,N_16277,N_16777);
and U17242 (N_17242,N_16284,N_16937);
or U17243 (N_17243,N_16056,N_16888);
nand U17244 (N_17244,N_16663,N_16333);
or U17245 (N_17245,N_16916,N_16070);
nor U17246 (N_17246,N_16941,N_16290);
xor U17247 (N_17247,N_16032,N_16177);
or U17248 (N_17248,N_16499,N_16238);
xnor U17249 (N_17249,N_16085,N_16566);
nor U17250 (N_17250,N_16472,N_16670);
xor U17251 (N_17251,N_16654,N_16977);
nor U17252 (N_17252,N_16549,N_16249);
nor U17253 (N_17253,N_16110,N_16932);
nor U17254 (N_17254,N_16746,N_16855);
nor U17255 (N_17255,N_16378,N_16986);
nor U17256 (N_17256,N_16561,N_16768);
nor U17257 (N_17257,N_16919,N_16966);
nand U17258 (N_17258,N_16017,N_16711);
and U17259 (N_17259,N_16004,N_16480);
nor U17260 (N_17260,N_16041,N_16037);
or U17261 (N_17261,N_16945,N_16604);
xnor U17262 (N_17262,N_16766,N_16167);
nand U17263 (N_17263,N_16797,N_16317);
and U17264 (N_17264,N_16455,N_16283);
nand U17265 (N_17265,N_16628,N_16246);
xnor U17266 (N_17266,N_16384,N_16094);
nand U17267 (N_17267,N_16306,N_16515);
nand U17268 (N_17268,N_16417,N_16597);
and U17269 (N_17269,N_16456,N_16500);
nand U17270 (N_17270,N_16379,N_16657);
or U17271 (N_17271,N_16841,N_16281);
nor U17272 (N_17272,N_16667,N_16093);
and U17273 (N_17273,N_16265,N_16892);
or U17274 (N_17274,N_16261,N_16513);
and U17275 (N_17275,N_16745,N_16747);
nand U17276 (N_17276,N_16635,N_16504);
xnor U17277 (N_17277,N_16510,N_16541);
nor U17278 (N_17278,N_16376,N_16706);
nand U17279 (N_17279,N_16220,N_16755);
nor U17280 (N_17280,N_16481,N_16451);
xnor U17281 (N_17281,N_16891,N_16627);
and U17282 (N_17282,N_16569,N_16353);
nand U17283 (N_17283,N_16052,N_16914);
nor U17284 (N_17284,N_16430,N_16199);
and U17285 (N_17285,N_16519,N_16433);
nor U17286 (N_17286,N_16885,N_16815);
nor U17287 (N_17287,N_16824,N_16068);
and U17288 (N_17288,N_16033,N_16382);
nor U17289 (N_17289,N_16221,N_16872);
nand U17290 (N_17290,N_16133,N_16390);
or U17291 (N_17291,N_16563,N_16019);
and U17292 (N_17292,N_16752,N_16023);
and U17293 (N_17293,N_16399,N_16470);
nand U17294 (N_17294,N_16904,N_16936);
nand U17295 (N_17295,N_16350,N_16623);
and U17296 (N_17296,N_16173,N_16158);
nor U17297 (N_17297,N_16676,N_16665);
or U17298 (N_17298,N_16226,N_16930);
and U17299 (N_17299,N_16467,N_16369);
and U17300 (N_17300,N_16211,N_16850);
nor U17301 (N_17301,N_16998,N_16867);
nand U17302 (N_17302,N_16684,N_16161);
xor U17303 (N_17303,N_16100,N_16619);
nor U17304 (N_17304,N_16089,N_16114);
nand U17305 (N_17305,N_16251,N_16955);
or U17306 (N_17306,N_16420,N_16796);
nor U17307 (N_17307,N_16527,N_16827);
nand U17308 (N_17308,N_16852,N_16545);
nor U17309 (N_17309,N_16860,N_16058);
xor U17310 (N_17310,N_16681,N_16835);
nor U17311 (N_17311,N_16575,N_16364);
or U17312 (N_17312,N_16156,N_16859);
nor U17313 (N_17313,N_16047,N_16522);
or U17314 (N_17314,N_16088,N_16842);
and U17315 (N_17315,N_16874,N_16903);
nor U17316 (N_17316,N_16204,N_16660);
or U17317 (N_17317,N_16460,N_16639);
nand U17318 (N_17318,N_16734,N_16425);
xor U17319 (N_17319,N_16448,N_16546);
nand U17320 (N_17320,N_16832,N_16638);
xnor U17321 (N_17321,N_16999,N_16398);
xor U17322 (N_17322,N_16214,N_16704);
and U17323 (N_17323,N_16939,N_16607);
xnor U17324 (N_17324,N_16121,N_16962);
and U17325 (N_17325,N_16973,N_16844);
nand U17326 (N_17326,N_16179,N_16594);
nand U17327 (N_17327,N_16278,N_16791);
or U17328 (N_17328,N_16910,N_16458);
and U17329 (N_17329,N_16509,N_16837);
xor U17330 (N_17330,N_16624,N_16414);
or U17331 (N_17331,N_16587,N_16437);
and U17332 (N_17332,N_16547,N_16483);
xnor U17333 (N_17333,N_16087,N_16326);
and U17334 (N_17334,N_16374,N_16147);
nand U17335 (N_17335,N_16851,N_16145);
nand U17336 (N_17336,N_16599,N_16066);
nand U17337 (N_17337,N_16909,N_16055);
xnor U17338 (N_17338,N_16700,N_16316);
xor U17339 (N_17339,N_16415,N_16980);
xor U17340 (N_17340,N_16737,N_16559);
nand U17341 (N_17341,N_16542,N_16778);
or U17342 (N_17342,N_16229,N_16045);
nand U17343 (N_17343,N_16897,N_16880);
or U17344 (N_17344,N_16232,N_16836);
and U17345 (N_17345,N_16478,N_16250);
xnor U17346 (N_17346,N_16969,N_16601);
nand U17347 (N_17347,N_16560,N_16543);
nand U17348 (N_17348,N_16011,N_16432);
or U17349 (N_17349,N_16726,N_16544);
xor U17350 (N_17350,N_16025,N_16967);
or U17351 (N_17351,N_16586,N_16219);
or U17352 (N_17352,N_16555,N_16825);
xor U17353 (N_17353,N_16256,N_16227);
xnor U17354 (N_17354,N_16964,N_16096);
xor U17355 (N_17355,N_16689,N_16222);
xor U17356 (N_17356,N_16525,N_16856);
nor U17357 (N_17357,N_16869,N_16634);
nor U17358 (N_17358,N_16553,N_16401);
xnor U17359 (N_17359,N_16026,N_16804);
nor U17360 (N_17360,N_16334,N_16889);
or U17361 (N_17361,N_16729,N_16104);
or U17362 (N_17362,N_16297,N_16395);
nor U17363 (N_17363,N_16896,N_16651);
nor U17364 (N_17364,N_16348,N_16495);
nor U17365 (N_17365,N_16533,N_16917);
nor U17366 (N_17366,N_16759,N_16300);
and U17367 (N_17367,N_16538,N_16328);
xnor U17368 (N_17368,N_16779,N_16485);
xor U17369 (N_17369,N_16710,N_16118);
nand U17370 (N_17370,N_16469,N_16189);
or U17371 (N_17371,N_16141,N_16637);
and U17372 (N_17372,N_16603,N_16053);
xnor U17373 (N_17373,N_16233,N_16154);
xor U17374 (N_17374,N_16686,N_16304);
or U17375 (N_17375,N_16453,N_16210);
xnor U17376 (N_17376,N_16833,N_16064);
nand U17377 (N_17377,N_16813,N_16440);
xnor U17378 (N_17378,N_16439,N_16963);
xnor U17379 (N_17379,N_16659,N_16574);
nor U17380 (N_17380,N_16692,N_16268);
xnor U17381 (N_17381,N_16464,N_16450);
nand U17382 (N_17382,N_16732,N_16307);
nand U17383 (N_17383,N_16192,N_16573);
nand U17384 (N_17384,N_16344,N_16332);
nand U17385 (N_17385,N_16082,N_16352);
and U17386 (N_17386,N_16593,N_16148);
and U17387 (N_17387,N_16298,N_16863);
nand U17388 (N_17388,N_16809,N_16988);
nand U17389 (N_17389,N_16380,N_16995);
nand U17390 (N_17390,N_16429,N_16441);
or U17391 (N_17391,N_16949,N_16940);
or U17392 (N_17392,N_16666,N_16697);
nand U17393 (N_17393,N_16225,N_16477);
xor U17394 (N_17394,N_16054,N_16805);
xnor U17395 (N_17395,N_16447,N_16242);
or U17396 (N_17396,N_16234,N_16609);
xnor U17397 (N_17397,N_16494,N_16360);
nor U17398 (N_17398,N_16293,N_16174);
xnor U17399 (N_17399,N_16426,N_16357);
or U17400 (N_17400,N_16389,N_16010);
or U17401 (N_17401,N_16102,N_16708);
nand U17402 (N_17402,N_16463,N_16403);
nor U17403 (N_17403,N_16213,N_16280);
nor U17404 (N_17404,N_16701,N_16457);
or U17405 (N_17405,N_16523,N_16230);
nand U17406 (N_17406,N_16633,N_16042);
or U17407 (N_17407,N_16373,N_16756);
xor U17408 (N_17408,N_16063,N_16347);
or U17409 (N_17409,N_16002,N_16884);
or U17410 (N_17410,N_16383,N_16190);
nand U17411 (N_17411,N_16471,N_16572);
xor U17412 (N_17412,N_16894,N_16030);
nor U17413 (N_17413,N_16034,N_16144);
or U17414 (N_17414,N_16806,N_16152);
and U17415 (N_17415,N_16539,N_16208);
nand U17416 (N_17416,N_16218,N_16163);
and U17417 (N_17417,N_16327,N_16259);
xnor U17418 (N_17418,N_16801,N_16946);
xor U17419 (N_17419,N_16864,N_16371);
nand U17420 (N_17420,N_16614,N_16200);
xor U17421 (N_17421,N_16820,N_16502);
and U17422 (N_17422,N_16550,N_16106);
xor U17423 (N_17423,N_16501,N_16818);
and U17424 (N_17424,N_16810,N_16771);
and U17425 (N_17425,N_16241,N_16748);
or U17426 (N_17426,N_16687,N_16997);
nand U17427 (N_17427,N_16921,N_16151);
nor U17428 (N_17428,N_16761,N_16375);
and U17429 (N_17429,N_16812,N_16385);
and U17430 (N_17430,N_16215,N_16615);
xor U17431 (N_17431,N_16407,N_16014);
or U17432 (N_17432,N_16611,N_16253);
xnor U17433 (N_17433,N_16592,N_16363);
xnor U17434 (N_17434,N_16292,N_16816);
nand U17435 (N_17435,N_16540,N_16243);
or U17436 (N_17436,N_16865,N_16526);
nand U17437 (N_17437,N_16240,N_16630);
and U17438 (N_17438,N_16505,N_16411);
and U17439 (N_17439,N_16829,N_16408);
xor U17440 (N_17440,N_16744,N_16532);
nor U17441 (N_17441,N_16171,N_16565);
xnor U17442 (N_17442,N_16713,N_16655);
nor U17443 (N_17443,N_16989,N_16366);
and U17444 (N_17444,N_16649,N_16266);
xor U17445 (N_17445,N_16022,N_16061);
xor U17446 (N_17446,N_16150,N_16035);
nor U17447 (N_17447,N_16695,N_16065);
nor U17448 (N_17448,N_16705,N_16722);
xnor U17449 (N_17449,N_16931,N_16808);
xnor U17450 (N_17450,N_16521,N_16013);
nand U17451 (N_17451,N_16585,N_16046);
and U17452 (N_17452,N_16260,N_16397);
nand U17453 (N_17453,N_16905,N_16015);
xnor U17454 (N_17454,N_16006,N_16273);
and U17455 (N_17455,N_16506,N_16873);
or U17456 (N_17456,N_16337,N_16741);
nand U17457 (N_17457,N_16636,N_16703);
and U17458 (N_17458,N_16740,N_16445);
nand U17459 (N_17459,N_16968,N_16774);
or U17460 (N_17460,N_16871,N_16476);
nor U17461 (N_17461,N_16802,N_16584);
xor U17462 (N_17462,N_16149,N_16180);
nand U17463 (N_17463,N_16224,N_16531);
nor U17464 (N_17464,N_16646,N_16422);
and U17465 (N_17465,N_16341,N_16691);
xor U17466 (N_17466,N_16576,N_16000);
and U17467 (N_17467,N_16739,N_16419);
xnor U17468 (N_17468,N_16702,N_16346);
xnor U17469 (N_17469,N_16134,N_16196);
and U17470 (N_17470,N_16516,N_16338);
xnor U17471 (N_17471,N_16406,N_16644);
or U17472 (N_17472,N_16556,N_16511);
nand U17473 (N_17473,N_16359,N_16473);
nand U17474 (N_17474,N_16996,N_16503);
or U17475 (N_17475,N_16928,N_16318);
nand U17476 (N_17476,N_16299,N_16276);
or U17477 (N_17477,N_16600,N_16083);
xnor U17478 (N_17478,N_16129,N_16551);
nand U17479 (N_17479,N_16616,N_16462);
and U17480 (N_17480,N_16049,N_16491);
xor U17481 (N_17481,N_16117,N_16817);
nor U17482 (N_17482,N_16673,N_16244);
nor U17483 (N_17483,N_16787,N_16482);
and U17484 (N_17484,N_16435,N_16223);
xor U17485 (N_17485,N_16848,N_16146);
and U17486 (N_17486,N_16712,N_16843);
and U17487 (N_17487,N_16645,N_16123);
nor U17488 (N_17488,N_16918,N_16126);
nor U17489 (N_17489,N_16309,N_16269);
and U17490 (N_17490,N_16974,N_16671);
nor U17491 (N_17491,N_16571,N_16678);
or U17492 (N_17492,N_16105,N_16160);
and U17493 (N_17493,N_16086,N_16193);
nor U17494 (N_17494,N_16876,N_16368);
or U17495 (N_17495,N_16062,N_16409);
nor U17496 (N_17496,N_16679,N_16205);
and U17497 (N_17497,N_16662,N_16078);
and U17498 (N_17498,N_16618,N_16354);
nand U17499 (N_17499,N_16956,N_16127);
nor U17500 (N_17500,N_16154,N_16005);
and U17501 (N_17501,N_16730,N_16473);
and U17502 (N_17502,N_16269,N_16933);
or U17503 (N_17503,N_16713,N_16756);
nor U17504 (N_17504,N_16209,N_16725);
xor U17505 (N_17505,N_16423,N_16469);
nand U17506 (N_17506,N_16775,N_16749);
and U17507 (N_17507,N_16281,N_16162);
nand U17508 (N_17508,N_16905,N_16497);
and U17509 (N_17509,N_16213,N_16037);
and U17510 (N_17510,N_16790,N_16025);
or U17511 (N_17511,N_16687,N_16557);
or U17512 (N_17512,N_16421,N_16740);
nand U17513 (N_17513,N_16607,N_16257);
or U17514 (N_17514,N_16514,N_16749);
or U17515 (N_17515,N_16649,N_16505);
or U17516 (N_17516,N_16949,N_16337);
nor U17517 (N_17517,N_16840,N_16126);
or U17518 (N_17518,N_16240,N_16263);
or U17519 (N_17519,N_16453,N_16343);
xor U17520 (N_17520,N_16547,N_16035);
nor U17521 (N_17521,N_16152,N_16275);
nor U17522 (N_17522,N_16361,N_16528);
nor U17523 (N_17523,N_16719,N_16041);
nand U17524 (N_17524,N_16594,N_16209);
and U17525 (N_17525,N_16454,N_16281);
or U17526 (N_17526,N_16813,N_16084);
and U17527 (N_17527,N_16605,N_16421);
or U17528 (N_17528,N_16630,N_16191);
or U17529 (N_17529,N_16298,N_16902);
and U17530 (N_17530,N_16103,N_16415);
and U17531 (N_17531,N_16758,N_16589);
and U17532 (N_17532,N_16372,N_16846);
nor U17533 (N_17533,N_16323,N_16935);
or U17534 (N_17534,N_16652,N_16874);
xor U17535 (N_17535,N_16410,N_16886);
nand U17536 (N_17536,N_16209,N_16502);
xnor U17537 (N_17537,N_16161,N_16730);
nand U17538 (N_17538,N_16072,N_16005);
nand U17539 (N_17539,N_16216,N_16991);
nor U17540 (N_17540,N_16053,N_16270);
and U17541 (N_17541,N_16604,N_16789);
nor U17542 (N_17542,N_16112,N_16863);
nand U17543 (N_17543,N_16321,N_16626);
nand U17544 (N_17544,N_16175,N_16786);
nor U17545 (N_17545,N_16722,N_16021);
nand U17546 (N_17546,N_16249,N_16923);
nand U17547 (N_17547,N_16040,N_16359);
nor U17548 (N_17548,N_16397,N_16673);
nand U17549 (N_17549,N_16903,N_16049);
or U17550 (N_17550,N_16900,N_16978);
nand U17551 (N_17551,N_16688,N_16368);
and U17552 (N_17552,N_16039,N_16406);
nand U17553 (N_17553,N_16617,N_16162);
nor U17554 (N_17554,N_16934,N_16720);
or U17555 (N_17555,N_16955,N_16836);
and U17556 (N_17556,N_16204,N_16800);
nor U17557 (N_17557,N_16307,N_16075);
nand U17558 (N_17558,N_16339,N_16192);
xor U17559 (N_17559,N_16719,N_16325);
nor U17560 (N_17560,N_16048,N_16637);
or U17561 (N_17561,N_16517,N_16244);
or U17562 (N_17562,N_16792,N_16352);
nand U17563 (N_17563,N_16295,N_16539);
nand U17564 (N_17564,N_16323,N_16481);
nor U17565 (N_17565,N_16401,N_16508);
or U17566 (N_17566,N_16453,N_16944);
or U17567 (N_17567,N_16480,N_16614);
nand U17568 (N_17568,N_16639,N_16139);
xnor U17569 (N_17569,N_16992,N_16065);
and U17570 (N_17570,N_16355,N_16421);
xnor U17571 (N_17571,N_16211,N_16922);
xor U17572 (N_17572,N_16408,N_16411);
nand U17573 (N_17573,N_16164,N_16249);
nor U17574 (N_17574,N_16783,N_16774);
nand U17575 (N_17575,N_16910,N_16465);
and U17576 (N_17576,N_16241,N_16822);
and U17577 (N_17577,N_16554,N_16888);
nand U17578 (N_17578,N_16078,N_16808);
and U17579 (N_17579,N_16687,N_16818);
nor U17580 (N_17580,N_16044,N_16291);
or U17581 (N_17581,N_16101,N_16757);
nand U17582 (N_17582,N_16072,N_16396);
xnor U17583 (N_17583,N_16049,N_16697);
nor U17584 (N_17584,N_16551,N_16684);
nor U17585 (N_17585,N_16997,N_16410);
or U17586 (N_17586,N_16631,N_16238);
nor U17587 (N_17587,N_16419,N_16467);
nand U17588 (N_17588,N_16363,N_16352);
xnor U17589 (N_17589,N_16471,N_16939);
nor U17590 (N_17590,N_16544,N_16393);
or U17591 (N_17591,N_16597,N_16326);
or U17592 (N_17592,N_16288,N_16063);
nand U17593 (N_17593,N_16756,N_16238);
nand U17594 (N_17594,N_16550,N_16175);
xor U17595 (N_17595,N_16453,N_16536);
and U17596 (N_17596,N_16972,N_16030);
nand U17597 (N_17597,N_16296,N_16791);
nand U17598 (N_17598,N_16233,N_16990);
and U17599 (N_17599,N_16719,N_16350);
nor U17600 (N_17600,N_16797,N_16976);
nand U17601 (N_17601,N_16328,N_16011);
and U17602 (N_17602,N_16488,N_16612);
nand U17603 (N_17603,N_16254,N_16243);
and U17604 (N_17604,N_16557,N_16103);
xor U17605 (N_17605,N_16279,N_16516);
and U17606 (N_17606,N_16457,N_16988);
nand U17607 (N_17607,N_16935,N_16420);
and U17608 (N_17608,N_16269,N_16184);
nor U17609 (N_17609,N_16612,N_16751);
and U17610 (N_17610,N_16730,N_16497);
and U17611 (N_17611,N_16175,N_16837);
or U17612 (N_17612,N_16552,N_16953);
xnor U17613 (N_17613,N_16174,N_16578);
nor U17614 (N_17614,N_16560,N_16339);
nor U17615 (N_17615,N_16849,N_16602);
and U17616 (N_17616,N_16711,N_16475);
nand U17617 (N_17617,N_16885,N_16991);
and U17618 (N_17618,N_16973,N_16993);
nor U17619 (N_17619,N_16926,N_16591);
nor U17620 (N_17620,N_16943,N_16492);
xnor U17621 (N_17621,N_16264,N_16095);
nand U17622 (N_17622,N_16891,N_16207);
nor U17623 (N_17623,N_16734,N_16644);
nor U17624 (N_17624,N_16879,N_16269);
xnor U17625 (N_17625,N_16804,N_16730);
nor U17626 (N_17626,N_16768,N_16492);
or U17627 (N_17627,N_16637,N_16547);
or U17628 (N_17628,N_16073,N_16875);
xor U17629 (N_17629,N_16246,N_16525);
xnor U17630 (N_17630,N_16774,N_16977);
or U17631 (N_17631,N_16203,N_16183);
or U17632 (N_17632,N_16134,N_16706);
nor U17633 (N_17633,N_16131,N_16018);
and U17634 (N_17634,N_16620,N_16539);
nor U17635 (N_17635,N_16260,N_16219);
or U17636 (N_17636,N_16357,N_16893);
nand U17637 (N_17637,N_16350,N_16886);
and U17638 (N_17638,N_16770,N_16319);
xnor U17639 (N_17639,N_16612,N_16860);
xnor U17640 (N_17640,N_16232,N_16100);
nand U17641 (N_17641,N_16693,N_16533);
or U17642 (N_17642,N_16580,N_16239);
nor U17643 (N_17643,N_16678,N_16886);
and U17644 (N_17644,N_16943,N_16895);
or U17645 (N_17645,N_16643,N_16148);
nor U17646 (N_17646,N_16388,N_16268);
or U17647 (N_17647,N_16943,N_16940);
xnor U17648 (N_17648,N_16992,N_16073);
and U17649 (N_17649,N_16418,N_16580);
xor U17650 (N_17650,N_16674,N_16254);
and U17651 (N_17651,N_16444,N_16775);
and U17652 (N_17652,N_16745,N_16090);
nor U17653 (N_17653,N_16762,N_16167);
nor U17654 (N_17654,N_16474,N_16389);
xor U17655 (N_17655,N_16929,N_16061);
xor U17656 (N_17656,N_16706,N_16972);
xor U17657 (N_17657,N_16026,N_16279);
or U17658 (N_17658,N_16155,N_16166);
xnor U17659 (N_17659,N_16697,N_16665);
nor U17660 (N_17660,N_16412,N_16327);
xor U17661 (N_17661,N_16287,N_16000);
xor U17662 (N_17662,N_16225,N_16035);
nor U17663 (N_17663,N_16193,N_16146);
or U17664 (N_17664,N_16799,N_16780);
xor U17665 (N_17665,N_16384,N_16012);
xor U17666 (N_17666,N_16029,N_16052);
nand U17667 (N_17667,N_16270,N_16378);
or U17668 (N_17668,N_16702,N_16341);
or U17669 (N_17669,N_16378,N_16212);
nand U17670 (N_17670,N_16584,N_16075);
nand U17671 (N_17671,N_16142,N_16003);
xnor U17672 (N_17672,N_16706,N_16726);
nor U17673 (N_17673,N_16184,N_16717);
or U17674 (N_17674,N_16687,N_16881);
nand U17675 (N_17675,N_16262,N_16405);
nand U17676 (N_17676,N_16736,N_16806);
nand U17677 (N_17677,N_16002,N_16479);
xnor U17678 (N_17678,N_16050,N_16125);
or U17679 (N_17679,N_16920,N_16613);
nor U17680 (N_17680,N_16529,N_16385);
and U17681 (N_17681,N_16974,N_16006);
nor U17682 (N_17682,N_16756,N_16312);
nand U17683 (N_17683,N_16365,N_16111);
and U17684 (N_17684,N_16423,N_16942);
nand U17685 (N_17685,N_16611,N_16636);
nor U17686 (N_17686,N_16007,N_16675);
nor U17687 (N_17687,N_16977,N_16130);
and U17688 (N_17688,N_16354,N_16897);
xnor U17689 (N_17689,N_16919,N_16640);
and U17690 (N_17690,N_16181,N_16493);
nand U17691 (N_17691,N_16323,N_16579);
nor U17692 (N_17692,N_16451,N_16072);
or U17693 (N_17693,N_16726,N_16955);
xnor U17694 (N_17694,N_16166,N_16532);
and U17695 (N_17695,N_16586,N_16635);
and U17696 (N_17696,N_16482,N_16353);
nor U17697 (N_17697,N_16232,N_16910);
or U17698 (N_17698,N_16649,N_16318);
and U17699 (N_17699,N_16951,N_16502);
or U17700 (N_17700,N_16641,N_16502);
nand U17701 (N_17701,N_16170,N_16235);
or U17702 (N_17702,N_16686,N_16363);
or U17703 (N_17703,N_16317,N_16882);
nor U17704 (N_17704,N_16220,N_16365);
or U17705 (N_17705,N_16894,N_16684);
or U17706 (N_17706,N_16680,N_16049);
and U17707 (N_17707,N_16852,N_16674);
and U17708 (N_17708,N_16357,N_16388);
xnor U17709 (N_17709,N_16354,N_16571);
xnor U17710 (N_17710,N_16390,N_16908);
nand U17711 (N_17711,N_16452,N_16481);
or U17712 (N_17712,N_16352,N_16584);
nor U17713 (N_17713,N_16613,N_16133);
and U17714 (N_17714,N_16415,N_16693);
or U17715 (N_17715,N_16294,N_16769);
nand U17716 (N_17716,N_16035,N_16520);
nand U17717 (N_17717,N_16107,N_16977);
nand U17718 (N_17718,N_16938,N_16734);
or U17719 (N_17719,N_16539,N_16435);
nand U17720 (N_17720,N_16087,N_16956);
nand U17721 (N_17721,N_16150,N_16562);
nor U17722 (N_17722,N_16372,N_16988);
and U17723 (N_17723,N_16724,N_16775);
and U17724 (N_17724,N_16191,N_16331);
nor U17725 (N_17725,N_16827,N_16432);
or U17726 (N_17726,N_16822,N_16063);
and U17727 (N_17727,N_16110,N_16658);
or U17728 (N_17728,N_16450,N_16609);
and U17729 (N_17729,N_16261,N_16976);
nor U17730 (N_17730,N_16329,N_16158);
xnor U17731 (N_17731,N_16076,N_16005);
and U17732 (N_17732,N_16680,N_16356);
nand U17733 (N_17733,N_16034,N_16478);
and U17734 (N_17734,N_16958,N_16272);
and U17735 (N_17735,N_16634,N_16485);
or U17736 (N_17736,N_16594,N_16024);
xor U17737 (N_17737,N_16652,N_16513);
nand U17738 (N_17738,N_16146,N_16044);
nand U17739 (N_17739,N_16506,N_16007);
nor U17740 (N_17740,N_16880,N_16928);
nand U17741 (N_17741,N_16708,N_16074);
or U17742 (N_17742,N_16509,N_16295);
nand U17743 (N_17743,N_16812,N_16529);
or U17744 (N_17744,N_16578,N_16096);
or U17745 (N_17745,N_16447,N_16317);
xnor U17746 (N_17746,N_16195,N_16800);
nor U17747 (N_17747,N_16151,N_16558);
or U17748 (N_17748,N_16661,N_16044);
nor U17749 (N_17749,N_16064,N_16257);
or U17750 (N_17750,N_16808,N_16322);
and U17751 (N_17751,N_16186,N_16242);
or U17752 (N_17752,N_16968,N_16769);
nand U17753 (N_17753,N_16067,N_16966);
xor U17754 (N_17754,N_16519,N_16128);
and U17755 (N_17755,N_16443,N_16471);
nand U17756 (N_17756,N_16964,N_16342);
nor U17757 (N_17757,N_16780,N_16509);
nor U17758 (N_17758,N_16432,N_16479);
xor U17759 (N_17759,N_16289,N_16483);
nor U17760 (N_17760,N_16367,N_16995);
or U17761 (N_17761,N_16559,N_16906);
or U17762 (N_17762,N_16923,N_16133);
nor U17763 (N_17763,N_16651,N_16041);
or U17764 (N_17764,N_16870,N_16694);
xor U17765 (N_17765,N_16728,N_16671);
xor U17766 (N_17766,N_16081,N_16663);
nand U17767 (N_17767,N_16112,N_16397);
or U17768 (N_17768,N_16349,N_16085);
nor U17769 (N_17769,N_16478,N_16025);
nand U17770 (N_17770,N_16226,N_16248);
nor U17771 (N_17771,N_16139,N_16200);
and U17772 (N_17772,N_16726,N_16112);
nand U17773 (N_17773,N_16205,N_16500);
or U17774 (N_17774,N_16476,N_16891);
nand U17775 (N_17775,N_16286,N_16301);
and U17776 (N_17776,N_16557,N_16784);
nand U17777 (N_17777,N_16081,N_16727);
and U17778 (N_17778,N_16082,N_16947);
or U17779 (N_17779,N_16742,N_16889);
and U17780 (N_17780,N_16310,N_16001);
nor U17781 (N_17781,N_16780,N_16796);
nand U17782 (N_17782,N_16548,N_16277);
nand U17783 (N_17783,N_16554,N_16506);
or U17784 (N_17784,N_16242,N_16256);
nor U17785 (N_17785,N_16947,N_16981);
xor U17786 (N_17786,N_16963,N_16526);
or U17787 (N_17787,N_16549,N_16961);
or U17788 (N_17788,N_16857,N_16818);
nand U17789 (N_17789,N_16210,N_16720);
nor U17790 (N_17790,N_16650,N_16088);
xor U17791 (N_17791,N_16618,N_16565);
nor U17792 (N_17792,N_16905,N_16179);
nor U17793 (N_17793,N_16626,N_16635);
xor U17794 (N_17794,N_16353,N_16288);
or U17795 (N_17795,N_16905,N_16156);
or U17796 (N_17796,N_16673,N_16478);
nand U17797 (N_17797,N_16836,N_16567);
or U17798 (N_17798,N_16670,N_16906);
or U17799 (N_17799,N_16237,N_16662);
nand U17800 (N_17800,N_16058,N_16730);
and U17801 (N_17801,N_16575,N_16244);
or U17802 (N_17802,N_16538,N_16913);
or U17803 (N_17803,N_16146,N_16419);
nor U17804 (N_17804,N_16727,N_16448);
nor U17805 (N_17805,N_16108,N_16983);
and U17806 (N_17806,N_16525,N_16548);
and U17807 (N_17807,N_16172,N_16082);
xnor U17808 (N_17808,N_16573,N_16696);
or U17809 (N_17809,N_16743,N_16330);
or U17810 (N_17810,N_16280,N_16283);
nor U17811 (N_17811,N_16856,N_16395);
xor U17812 (N_17812,N_16439,N_16066);
xor U17813 (N_17813,N_16513,N_16027);
or U17814 (N_17814,N_16844,N_16628);
nor U17815 (N_17815,N_16573,N_16727);
and U17816 (N_17816,N_16067,N_16518);
xnor U17817 (N_17817,N_16527,N_16253);
nand U17818 (N_17818,N_16888,N_16739);
nor U17819 (N_17819,N_16727,N_16652);
nor U17820 (N_17820,N_16085,N_16093);
or U17821 (N_17821,N_16502,N_16701);
nand U17822 (N_17822,N_16557,N_16345);
or U17823 (N_17823,N_16171,N_16229);
xnor U17824 (N_17824,N_16323,N_16745);
or U17825 (N_17825,N_16057,N_16427);
and U17826 (N_17826,N_16134,N_16141);
nor U17827 (N_17827,N_16049,N_16155);
xor U17828 (N_17828,N_16495,N_16401);
and U17829 (N_17829,N_16075,N_16646);
xor U17830 (N_17830,N_16836,N_16574);
nand U17831 (N_17831,N_16683,N_16834);
nand U17832 (N_17832,N_16270,N_16781);
nor U17833 (N_17833,N_16619,N_16796);
nand U17834 (N_17834,N_16852,N_16412);
xnor U17835 (N_17835,N_16386,N_16869);
and U17836 (N_17836,N_16137,N_16213);
nor U17837 (N_17837,N_16432,N_16007);
or U17838 (N_17838,N_16315,N_16560);
and U17839 (N_17839,N_16922,N_16235);
and U17840 (N_17840,N_16756,N_16129);
or U17841 (N_17841,N_16071,N_16898);
and U17842 (N_17842,N_16097,N_16583);
nand U17843 (N_17843,N_16586,N_16814);
nand U17844 (N_17844,N_16834,N_16864);
or U17845 (N_17845,N_16077,N_16997);
nor U17846 (N_17846,N_16410,N_16562);
xor U17847 (N_17847,N_16042,N_16119);
or U17848 (N_17848,N_16818,N_16755);
nand U17849 (N_17849,N_16898,N_16698);
xor U17850 (N_17850,N_16377,N_16235);
nor U17851 (N_17851,N_16459,N_16552);
nor U17852 (N_17852,N_16272,N_16177);
nor U17853 (N_17853,N_16271,N_16182);
nand U17854 (N_17854,N_16107,N_16638);
nand U17855 (N_17855,N_16767,N_16902);
nor U17856 (N_17856,N_16897,N_16133);
and U17857 (N_17857,N_16928,N_16953);
and U17858 (N_17858,N_16929,N_16382);
nand U17859 (N_17859,N_16982,N_16172);
xor U17860 (N_17860,N_16897,N_16728);
or U17861 (N_17861,N_16015,N_16613);
or U17862 (N_17862,N_16581,N_16867);
and U17863 (N_17863,N_16108,N_16145);
nand U17864 (N_17864,N_16703,N_16789);
or U17865 (N_17865,N_16484,N_16361);
nor U17866 (N_17866,N_16941,N_16495);
and U17867 (N_17867,N_16436,N_16434);
nand U17868 (N_17868,N_16587,N_16200);
and U17869 (N_17869,N_16699,N_16277);
nor U17870 (N_17870,N_16564,N_16809);
nand U17871 (N_17871,N_16489,N_16382);
and U17872 (N_17872,N_16326,N_16497);
xor U17873 (N_17873,N_16458,N_16621);
xnor U17874 (N_17874,N_16521,N_16112);
nand U17875 (N_17875,N_16547,N_16554);
and U17876 (N_17876,N_16400,N_16026);
nor U17877 (N_17877,N_16694,N_16322);
and U17878 (N_17878,N_16812,N_16314);
and U17879 (N_17879,N_16452,N_16887);
xnor U17880 (N_17880,N_16139,N_16699);
or U17881 (N_17881,N_16131,N_16144);
nor U17882 (N_17882,N_16784,N_16279);
xnor U17883 (N_17883,N_16035,N_16176);
and U17884 (N_17884,N_16203,N_16571);
or U17885 (N_17885,N_16345,N_16615);
nor U17886 (N_17886,N_16223,N_16551);
nor U17887 (N_17887,N_16499,N_16725);
nor U17888 (N_17888,N_16338,N_16442);
and U17889 (N_17889,N_16963,N_16342);
xor U17890 (N_17890,N_16872,N_16671);
nand U17891 (N_17891,N_16927,N_16410);
xnor U17892 (N_17892,N_16367,N_16959);
nor U17893 (N_17893,N_16510,N_16662);
nand U17894 (N_17894,N_16399,N_16652);
nor U17895 (N_17895,N_16363,N_16413);
and U17896 (N_17896,N_16156,N_16682);
xnor U17897 (N_17897,N_16885,N_16186);
nand U17898 (N_17898,N_16850,N_16100);
or U17899 (N_17899,N_16751,N_16282);
and U17900 (N_17900,N_16873,N_16373);
nor U17901 (N_17901,N_16899,N_16361);
nand U17902 (N_17902,N_16762,N_16973);
and U17903 (N_17903,N_16095,N_16675);
nand U17904 (N_17904,N_16558,N_16259);
xor U17905 (N_17905,N_16259,N_16248);
or U17906 (N_17906,N_16755,N_16837);
or U17907 (N_17907,N_16127,N_16033);
nor U17908 (N_17908,N_16231,N_16581);
nor U17909 (N_17909,N_16647,N_16044);
nor U17910 (N_17910,N_16996,N_16768);
nor U17911 (N_17911,N_16662,N_16074);
or U17912 (N_17912,N_16165,N_16946);
xnor U17913 (N_17913,N_16985,N_16726);
xor U17914 (N_17914,N_16088,N_16743);
and U17915 (N_17915,N_16842,N_16060);
nor U17916 (N_17916,N_16120,N_16295);
or U17917 (N_17917,N_16223,N_16198);
xnor U17918 (N_17918,N_16532,N_16547);
or U17919 (N_17919,N_16772,N_16575);
nor U17920 (N_17920,N_16050,N_16750);
or U17921 (N_17921,N_16055,N_16514);
xnor U17922 (N_17922,N_16666,N_16761);
xnor U17923 (N_17923,N_16353,N_16195);
nand U17924 (N_17924,N_16026,N_16479);
nand U17925 (N_17925,N_16939,N_16750);
nor U17926 (N_17926,N_16021,N_16316);
nand U17927 (N_17927,N_16351,N_16430);
nor U17928 (N_17928,N_16048,N_16273);
xor U17929 (N_17929,N_16820,N_16747);
or U17930 (N_17930,N_16273,N_16417);
or U17931 (N_17931,N_16888,N_16799);
and U17932 (N_17932,N_16009,N_16719);
or U17933 (N_17933,N_16520,N_16904);
nand U17934 (N_17934,N_16715,N_16527);
or U17935 (N_17935,N_16528,N_16166);
nand U17936 (N_17936,N_16106,N_16115);
nand U17937 (N_17937,N_16930,N_16880);
nand U17938 (N_17938,N_16145,N_16656);
nand U17939 (N_17939,N_16634,N_16217);
nand U17940 (N_17940,N_16320,N_16389);
nor U17941 (N_17941,N_16120,N_16401);
nor U17942 (N_17942,N_16971,N_16319);
or U17943 (N_17943,N_16841,N_16482);
xnor U17944 (N_17944,N_16895,N_16696);
and U17945 (N_17945,N_16563,N_16711);
nand U17946 (N_17946,N_16847,N_16041);
xnor U17947 (N_17947,N_16983,N_16588);
or U17948 (N_17948,N_16022,N_16384);
nand U17949 (N_17949,N_16150,N_16164);
xor U17950 (N_17950,N_16409,N_16046);
and U17951 (N_17951,N_16500,N_16574);
nor U17952 (N_17952,N_16100,N_16710);
and U17953 (N_17953,N_16288,N_16054);
nand U17954 (N_17954,N_16523,N_16136);
and U17955 (N_17955,N_16998,N_16514);
or U17956 (N_17956,N_16489,N_16998);
and U17957 (N_17957,N_16644,N_16421);
and U17958 (N_17958,N_16380,N_16014);
and U17959 (N_17959,N_16944,N_16581);
or U17960 (N_17960,N_16503,N_16129);
xnor U17961 (N_17961,N_16906,N_16289);
xnor U17962 (N_17962,N_16556,N_16799);
and U17963 (N_17963,N_16159,N_16694);
or U17964 (N_17964,N_16103,N_16169);
xor U17965 (N_17965,N_16464,N_16808);
xnor U17966 (N_17966,N_16212,N_16990);
nand U17967 (N_17967,N_16572,N_16906);
and U17968 (N_17968,N_16660,N_16654);
xor U17969 (N_17969,N_16191,N_16555);
and U17970 (N_17970,N_16163,N_16663);
nand U17971 (N_17971,N_16084,N_16860);
nor U17972 (N_17972,N_16407,N_16949);
xnor U17973 (N_17973,N_16415,N_16701);
or U17974 (N_17974,N_16372,N_16155);
nand U17975 (N_17975,N_16535,N_16714);
or U17976 (N_17976,N_16965,N_16090);
xor U17977 (N_17977,N_16255,N_16271);
and U17978 (N_17978,N_16346,N_16442);
nor U17979 (N_17979,N_16978,N_16726);
and U17980 (N_17980,N_16291,N_16185);
and U17981 (N_17981,N_16710,N_16190);
nor U17982 (N_17982,N_16556,N_16984);
xor U17983 (N_17983,N_16451,N_16812);
or U17984 (N_17984,N_16677,N_16022);
xnor U17985 (N_17985,N_16849,N_16442);
nand U17986 (N_17986,N_16245,N_16150);
nand U17987 (N_17987,N_16456,N_16678);
xor U17988 (N_17988,N_16670,N_16753);
and U17989 (N_17989,N_16322,N_16096);
nand U17990 (N_17990,N_16296,N_16587);
and U17991 (N_17991,N_16524,N_16788);
nor U17992 (N_17992,N_16834,N_16616);
or U17993 (N_17993,N_16526,N_16284);
nor U17994 (N_17994,N_16952,N_16164);
nand U17995 (N_17995,N_16794,N_16845);
and U17996 (N_17996,N_16381,N_16311);
and U17997 (N_17997,N_16628,N_16165);
xor U17998 (N_17998,N_16959,N_16364);
or U17999 (N_17999,N_16748,N_16267);
and U18000 (N_18000,N_17960,N_17931);
xnor U18001 (N_18001,N_17118,N_17881);
and U18002 (N_18002,N_17900,N_17448);
nor U18003 (N_18003,N_17023,N_17499);
or U18004 (N_18004,N_17876,N_17884);
and U18005 (N_18005,N_17864,N_17858);
and U18006 (N_18006,N_17068,N_17832);
or U18007 (N_18007,N_17522,N_17665);
nor U18008 (N_18008,N_17319,N_17403);
nor U18009 (N_18009,N_17315,N_17365);
xnor U18010 (N_18010,N_17214,N_17254);
nand U18011 (N_18011,N_17204,N_17057);
nand U18012 (N_18012,N_17503,N_17898);
xor U18013 (N_18013,N_17276,N_17744);
or U18014 (N_18014,N_17153,N_17021);
nor U18015 (N_18015,N_17887,N_17821);
nor U18016 (N_18016,N_17544,N_17263);
or U18017 (N_18017,N_17280,N_17590);
and U18018 (N_18018,N_17004,N_17194);
nand U18019 (N_18019,N_17048,N_17981);
nand U18020 (N_18020,N_17622,N_17104);
and U18021 (N_18021,N_17570,N_17686);
nand U18022 (N_18022,N_17218,N_17636);
or U18023 (N_18023,N_17650,N_17516);
nand U18024 (N_18024,N_17201,N_17607);
nor U18025 (N_18025,N_17086,N_17666);
nand U18026 (N_18026,N_17661,N_17331);
nand U18027 (N_18027,N_17386,N_17219);
and U18028 (N_18028,N_17682,N_17890);
nand U18029 (N_18029,N_17547,N_17766);
nor U18030 (N_18030,N_17482,N_17537);
and U18031 (N_18031,N_17690,N_17593);
nand U18032 (N_18032,N_17364,N_17402);
nand U18033 (N_18033,N_17565,N_17756);
xor U18034 (N_18034,N_17813,N_17579);
and U18035 (N_18035,N_17974,N_17770);
or U18036 (N_18036,N_17101,N_17188);
or U18037 (N_18037,N_17055,N_17606);
nor U18038 (N_18038,N_17663,N_17352);
or U18039 (N_18039,N_17645,N_17297);
or U18040 (N_18040,N_17562,N_17444);
nor U18041 (N_18041,N_17311,N_17888);
and U18042 (N_18042,N_17385,N_17563);
nor U18043 (N_18043,N_17839,N_17809);
nor U18044 (N_18044,N_17914,N_17873);
xnor U18045 (N_18045,N_17451,N_17082);
and U18046 (N_18046,N_17878,N_17706);
or U18047 (N_18047,N_17715,N_17853);
or U18048 (N_18048,N_17559,N_17374);
xor U18049 (N_18049,N_17735,N_17709);
xnor U18050 (N_18050,N_17024,N_17327);
and U18051 (N_18051,N_17711,N_17928);
nand U18052 (N_18052,N_17626,N_17775);
nand U18053 (N_18053,N_17932,N_17309);
and U18054 (N_18054,N_17748,N_17944);
or U18055 (N_18055,N_17520,N_17697);
and U18056 (N_18056,N_17467,N_17705);
nor U18057 (N_18057,N_17976,N_17029);
and U18058 (N_18058,N_17003,N_17133);
xor U18059 (N_18059,N_17526,N_17824);
and U18060 (N_18060,N_17927,N_17993);
or U18061 (N_18061,N_17883,N_17147);
nor U18062 (N_18062,N_17483,N_17321);
or U18063 (N_18063,N_17217,N_17267);
nand U18064 (N_18064,N_17816,N_17435);
xnor U18065 (N_18065,N_17480,N_17026);
nand U18066 (N_18066,N_17595,N_17288);
nor U18067 (N_18067,N_17936,N_17432);
or U18068 (N_18068,N_17059,N_17320);
nand U18069 (N_18069,N_17774,N_17156);
and U18070 (N_18070,N_17145,N_17238);
and U18071 (N_18071,N_17810,N_17140);
xor U18072 (N_18072,N_17100,N_17693);
xnor U18073 (N_18073,N_17269,N_17558);
nor U18074 (N_18074,N_17621,N_17628);
nand U18075 (N_18075,N_17287,N_17310);
nand U18076 (N_18076,N_17488,N_17151);
or U18077 (N_18077,N_17506,N_17185);
or U18078 (N_18078,N_17507,N_17747);
or U18079 (N_18079,N_17815,N_17787);
and U18080 (N_18080,N_17250,N_17519);
xnor U18081 (N_18081,N_17995,N_17769);
nor U18082 (N_18082,N_17644,N_17283);
nand U18083 (N_18083,N_17417,N_17964);
nor U18084 (N_18084,N_17889,N_17925);
and U18085 (N_18085,N_17175,N_17729);
or U18086 (N_18086,N_17160,N_17253);
and U18087 (N_18087,N_17084,N_17648);
nand U18088 (N_18088,N_17397,N_17973);
xnor U18089 (N_18089,N_17676,N_17657);
and U18090 (N_18090,N_17235,N_17578);
nand U18091 (N_18091,N_17117,N_17349);
nor U18092 (N_18092,N_17796,N_17335);
or U18093 (N_18093,N_17683,N_17861);
and U18094 (N_18094,N_17481,N_17285);
xnor U18095 (N_18095,N_17954,N_17672);
or U18096 (N_18096,N_17505,N_17389);
or U18097 (N_18097,N_17033,N_17486);
or U18098 (N_18098,N_17080,N_17767);
nor U18099 (N_18099,N_17604,N_17571);
xor U18100 (N_18100,N_17660,N_17687);
and U18101 (N_18101,N_17893,N_17536);
and U18102 (N_18102,N_17162,N_17124);
and U18103 (N_18103,N_17865,N_17216);
or U18104 (N_18104,N_17127,N_17679);
or U18105 (N_18105,N_17196,N_17724);
xor U18106 (N_18106,N_17044,N_17172);
xnor U18107 (N_18107,N_17684,N_17500);
and U18108 (N_18108,N_17783,N_17001);
xnor U18109 (N_18109,N_17336,N_17180);
xor U18110 (N_18110,N_17840,N_17996);
and U18111 (N_18111,N_17485,N_17475);
nand U18112 (N_18112,N_17785,N_17983);
or U18113 (N_18113,N_17056,N_17857);
nand U18114 (N_18114,N_17939,N_17305);
nand U18115 (N_18115,N_17940,N_17535);
or U18116 (N_18116,N_17081,N_17961);
nand U18117 (N_18117,N_17491,N_17183);
nor U18118 (N_18118,N_17209,N_17806);
and U18119 (N_18119,N_17047,N_17798);
or U18120 (N_18120,N_17376,N_17064);
and U18121 (N_18121,N_17600,N_17812);
nor U18122 (N_18122,N_17054,N_17521);
nor U18123 (N_18123,N_17306,N_17041);
and U18124 (N_18124,N_17119,N_17399);
nand U18125 (N_18125,N_17843,N_17510);
xnor U18126 (N_18126,N_17249,N_17173);
and U18127 (N_18127,N_17027,N_17191);
nand U18128 (N_18128,N_17777,N_17354);
nor U18129 (N_18129,N_17791,N_17513);
and U18130 (N_18130,N_17831,N_17692);
nor U18131 (N_18131,N_17919,N_17942);
xnor U18132 (N_18132,N_17548,N_17149);
xnor U18133 (N_18133,N_17624,N_17242);
xor U18134 (N_18134,N_17493,N_17805);
nor U18135 (N_18135,N_17459,N_17362);
and U18136 (N_18136,N_17006,N_17233);
nor U18137 (N_18137,N_17159,N_17032);
or U18138 (N_18138,N_17419,N_17130);
and U18139 (N_18139,N_17933,N_17912);
nand U18140 (N_18140,N_17643,N_17018);
and U18141 (N_18141,N_17637,N_17257);
and U18142 (N_18142,N_17552,N_17969);
xnor U18143 (N_18143,N_17065,N_17302);
nor U18144 (N_18144,N_17340,N_17157);
nand U18145 (N_18145,N_17366,N_17759);
nand U18146 (N_18146,N_17398,N_17922);
and U18147 (N_18147,N_17010,N_17886);
xnor U18148 (N_18148,N_17022,N_17241);
nand U18149 (N_18149,N_17923,N_17512);
and U18150 (N_18150,N_17811,N_17163);
and U18151 (N_18151,N_17025,N_17146);
xnor U18152 (N_18152,N_17955,N_17168);
nand U18153 (N_18153,N_17076,N_17358);
and U18154 (N_18154,N_17437,N_17950);
xor U18155 (N_18155,N_17273,N_17430);
and U18156 (N_18156,N_17958,N_17980);
and U18157 (N_18157,N_17746,N_17443);
or U18158 (N_18158,N_17458,N_17685);
xnor U18159 (N_18159,N_17087,N_17719);
or U18160 (N_18160,N_17844,N_17596);
nand U18161 (N_18161,N_17568,N_17763);
or U18162 (N_18162,N_17487,N_17930);
nand U18163 (N_18163,N_17123,N_17136);
xnor U18164 (N_18164,N_17880,N_17765);
nor U18165 (N_18165,N_17538,N_17296);
and U18166 (N_18166,N_17879,N_17557);
nand U18167 (N_18167,N_17126,N_17688);
and U18168 (N_18168,N_17202,N_17268);
and U18169 (N_18169,N_17782,N_17412);
and U18170 (N_18170,N_17633,N_17074);
nand U18171 (N_18171,N_17523,N_17077);
nor U18172 (N_18172,N_17978,N_17083);
xor U18173 (N_18173,N_17051,N_17000);
nand U18174 (N_18174,N_17852,N_17453);
xnor U18175 (N_18175,N_17116,N_17371);
and U18176 (N_18176,N_17792,N_17418);
and U18177 (N_18177,N_17728,N_17921);
nand U18178 (N_18178,N_17885,N_17847);
nor U18179 (N_18179,N_17461,N_17438);
xnor U18180 (N_18180,N_17205,N_17971);
or U18181 (N_18181,N_17870,N_17742);
or U18182 (N_18182,N_17704,N_17441);
xnor U18183 (N_18183,N_17723,N_17727);
xor U18184 (N_18184,N_17028,N_17178);
xnor U18185 (N_18185,N_17042,N_17749);
xnor U18186 (N_18186,N_17429,N_17977);
nand U18187 (N_18187,N_17261,N_17494);
and U18188 (N_18188,N_17129,N_17255);
and U18189 (N_18189,N_17143,N_17407);
nand U18190 (N_18190,N_17308,N_17786);
nor U18191 (N_18191,N_17543,N_17067);
nor U18192 (N_18192,N_17752,N_17150);
nand U18193 (N_18193,N_17471,N_17702);
xnor U18194 (N_18194,N_17089,N_17542);
xor U18195 (N_18195,N_17569,N_17212);
nand U18196 (N_18196,N_17618,N_17328);
or U18197 (N_18197,N_17532,N_17337);
nor U18198 (N_18198,N_17095,N_17525);
nor U18199 (N_18199,N_17445,N_17918);
or U18200 (N_18200,N_17186,N_17620);
nand U18201 (N_18201,N_17612,N_17381);
nor U18202 (N_18202,N_17988,N_17353);
and U18203 (N_18203,N_17017,N_17979);
xnor U18204 (N_18204,N_17841,N_17224);
or U18205 (N_18205,N_17799,N_17192);
nor U18206 (N_18206,N_17608,N_17093);
xor U18207 (N_18207,N_17300,N_17514);
and U18208 (N_18208,N_17098,N_17091);
nand U18209 (N_18209,N_17414,N_17694);
nor U18210 (N_18210,N_17587,N_17479);
xor U18211 (N_18211,N_17793,N_17274);
xor U18212 (N_18212,N_17573,N_17511);
or U18213 (N_18213,N_17314,N_17278);
and U18214 (N_18214,N_17994,N_17073);
nor U18215 (N_18215,N_17710,N_17771);
nor U18216 (N_18216,N_17915,N_17415);
nand U18217 (N_18217,N_17627,N_17154);
nor U18218 (N_18218,N_17721,N_17240);
nor U18219 (N_18219,N_17855,N_17111);
nand U18220 (N_18220,N_17105,N_17322);
or U18221 (N_18221,N_17541,N_17373);
and U18222 (N_18222,N_17016,N_17210);
xor U18223 (N_18223,N_17819,N_17997);
nand U18224 (N_18224,N_17225,N_17518);
xor U18225 (N_18225,N_17141,N_17937);
nand U18226 (N_18226,N_17462,N_17298);
nor U18227 (N_18227,N_17295,N_17052);
and U18228 (N_18228,N_17651,N_17517);
nand U18229 (N_18229,N_17708,N_17303);
and U18230 (N_18230,N_17592,N_17677);
or U18231 (N_18231,N_17442,N_17031);
and U18232 (N_18232,N_17096,N_17072);
nand U18233 (N_18233,N_17422,N_17588);
xor U18234 (N_18234,N_17948,N_17874);
or U18235 (N_18235,N_17013,N_17170);
and U18236 (N_18236,N_17454,N_17700);
or U18237 (N_18237,N_17952,N_17860);
and U18238 (N_18238,N_17470,N_17795);
nand U18239 (N_18239,N_17668,N_17489);
nand U18240 (N_18240,N_17907,N_17316);
nand U18241 (N_18241,N_17058,N_17986);
or U18242 (N_18242,N_17002,N_17972);
xor U18243 (N_18243,N_17911,N_17745);
xor U18244 (N_18244,N_17891,N_17585);
nor U18245 (N_18245,N_17803,N_17991);
nand U18246 (N_18246,N_17797,N_17778);
and U18247 (N_18247,N_17895,N_17780);
xor U18248 (N_18248,N_17121,N_17359);
xor U18249 (N_18249,N_17220,N_17594);
nor U18250 (N_18250,N_17040,N_17099);
or U18251 (N_18251,N_17404,N_17102);
nand U18252 (N_18252,N_17339,N_17773);
nand U18253 (N_18253,N_17670,N_17179);
nand U18254 (N_18254,N_17674,N_17968);
xnor U18255 (N_18255,N_17882,N_17826);
nor U18256 (N_18256,N_17591,N_17369);
xnor U18257 (N_18257,N_17122,N_17182);
and U18258 (N_18258,N_17176,N_17938);
nor U18259 (N_18259,N_17346,N_17158);
and U18260 (N_18260,N_17695,N_17726);
or U18261 (N_18261,N_17265,N_17598);
xnor U18262 (N_18262,N_17602,N_17734);
nor U18263 (N_18263,N_17609,N_17649);
nor U18264 (N_18264,N_17189,N_17334);
nand U18265 (N_18265,N_17085,N_17232);
and U18266 (N_18266,N_17449,N_17851);
xor U18267 (N_18267,N_17312,N_17758);
and U18268 (N_18268,N_17347,N_17393);
xor U18269 (N_18269,N_17820,N_17455);
or U18270 (N_18270,N_17707,N_17601);
and U18271 (N_18271,N_17920,N_17446);
or U18272 (N_18272,N_17534,N_17061);
nor U18273 (N_18273,N_17464,N_17379);
and U18274 (N_18274,N_17575,N_17106);
and U18275 (N_18275,N_17800,N_17753);
or U18276 (N_18276,N_17924,N_17062);
and U18277 (N_18277,N_17460,N_17850);
nand U18278 (N_18278,N_17060,N_17239);
nand U18279 (N_18279,N_17531,N_17007);
or U18280 (N_18280,N_17410,N_17329);
or U18281 (N_18281,N_17050,N_17551);
xnor U18282 (N_18282,N_17867,N_17560);
or U18283 (N_18283,N_17152,N_17277);
nand U18284 (N_18284,N_17063,N_17272);
xor U18285 (N_18285,N_17134,N_17014);
and U18286 (N_18286,N_17229,N_17206);
or U18287 (N_18287,N_17208,N_17474);
and U18288 (N_18288,N_17230,N_17553);
xor U18289 (N_18289,N_17361,N_17236);
and U18290 (N_18290,N_17248,N_17110);
nor U18291 (N_18291,N_17641,N_17228);
nand U18292 (N_18292,N_17681,N_17680);
xor U18293 (N_18293,N_17492,N_17034);
and U18294 (N_18294,N_17664,N_17713);
and U18295 (N_18295,N_17078,N_17463);
xnor U18296 (N_18296,N_17282,N_17781);
nor U18297 (N_18297,N_17762,N_17155);
or U18298 (N_18298,N_17655,N_17258);
and U18299 (N_18299,N_17625,N_17203);
or U18300 (N_18300,N_17975,N_17868);
nand U18301 (N_18301,N_17545,N_17367);
nand U18302 (N_18302,N_17869,N_17350);
nand U18303 (N_18303,N_17355,N_17733);
or U18304 (N_18304,N_17572,N_17112);
nor U18305 (N_18305,N_17425,N_17807);
xnor U18306 (N_18306,N_17356,N_17529);
xnor U18307 (N_18307,N_17689,N_17788);
or U18308 (N_18308,N_17848,N_17019);
xor U18309 (N_18309,N_17577,N_17424);
nor U18310 (N_18310,N_17142,N_17963);
or U18311 (N_18311,N_17834,N_17951);
nor U18312 (N_18312,N_17989,N_17631);
and U18313 (N_18313,N_17131,N_17223);
xor U18314 (N_18314,N_17539,N_17739);
or U18315 (N_18315,N_17408,N_17009);
or U18316 (N_18316,N_17549,N_17862);
nand U18317 (N_18317,N_17957,N_17264);
nand U18318 (N_18318,N_17290,N_17043);
and U18319 (N_18319,N_17830,N_17108);
or U18320 (N_18320,N_17428,N_17910);
xnor U18321 (N_18321,N_17439,N_17431);
nand U18322 (N_18322,N_17699,N_17284);
nor U18323 (N_18323,N_17999,N_17849);
nand U18324 (N_18324,N_17908,N_17671);
xor U18325 (N_18325,N_17956,N_17226);
or U18326 (N_18326,N_17630,N_17751);
or U18327 (N_18327,N_17262,N_17802);
xnor U18328 (N_18328,N_17383,N_17966);
or U18329 (N_18329,N_17351,N_17259);
xnor U18330 (N_18330,N_17754,N_17892);
or U18331 (N_18331,N_17103,N_17243);
or U18332 (N_18332,N_17421,N_17332);
xor U18333 (N_18333,N_17712,N_17164);
xnor U18334 (N_18334,N_17617,N_17294);
nor U18335 (N_18335,N_17396,N_17501);
nor U18336 (N_18336,N_17732,N_17490);
nand U18337 (N_18337,N_17171,N_17270);
nor U18338 (N_18338,N_17360,N_17465);
nand U18339 (N_18339,N_17252,N_17616);
xor U18340 (N_18340,N_17629,N_17846);
nand U18341 (N_18341,N_17401,N_17395);
xor U18342 (N_18342,N_17139,N_17370);
and U18343 (N_18343,N_17597,N_17498);
and U18344 (N_18344,N_17527,N_17835);
nor U18345 (N_18345,N_17720,N_17193);
xor U18346 (N_18346,N_17198,N_17941);
xnor U18347 (N_18347,N_17279,N_17015);
xor U18348 (N_18348,N_17905,N_17825);
or U18349 (N_18349,N_17037,N_17039);
and U18350 (N_18350,N_17266,N_17292);
and U18351 (N_18351,N_17447,N_17906);
xnor U18352 (N_18352,N_17776,N_17213);
and U18353 (N_18353,N_17466,N_17094);
nand U18354 (N_18354,N_17632,N_17184);
nand U18355 (N_18355,N_17662,N_17949);
nor U18356 (N_18356,N_17372,N_17012);
xnor U18357 (N_18357,N_17934,N_17169);
and U18358 (N_18358,N_17363,N_17947);
nor U18359 (N_18359,N_17614,N_17515);
or U18360 (N_18360,N_17231,N_17814);
xor U18361 (N_18361,N_17245,N_17234);
xor U18362 (N_18362,N_17634,N_17605);
xor U18363 (N_18363,N_17829,N_17165);
and U18364 (N_18364,N_17842,N_17987);
and U18365 (N_18365,N_17546,N_17768);
nor U18366 (N_18366,N_17313,N_17789);
xnor U18367 (N_18367,N_17005,N_17066);
xor U18368 (N_18368,N_17181,N_17413);
or U18369 (N_18369,N_17380,N_17992);
nor U18370 (N_18370,N_17528,N_17200);
xor U18371 (N_18371,N_17148,N_17502);
nand U18372 (N_18372,N_17045,N_17187);
or U18373 (N_18373,N_17092,N_17652);
or U18374 (N_18374,N_17576,N_17866);
or U18375 (N_18375,N_17472,N_17678);
and U18376 (N_18376,N_17237,N_17333);
nand U18377 (N_18377,N_17275,N_17701);
or U18378 (N_18378,N_17916,N_17613);
xor U18379 (N_18379,N_17901,N_17642);
nor U18380 (N_18380,N_17097,N_17473);
or U18381 (N_18381,N_17808,N_17669);
and U18382 (N_18382,N_17877,N_17190);
and U18383 (N_18383,N_17260,N_17195);
nor U18384 (N_18384,N_17790,N_17725);
xor U18385 (N_18385,N_17343,N_17524);
nand U18386 (N_18386,N_17875,N_17090);
or U18387 (N_18387,N_17113,N_17132);
nor U18388 (N_18388,N_17138,N_17691);
nand U18389 (N_18389,N_17304,N_17659);
and U18390 (N_18390,N_17069,N_17567);
or U18391 (N_18391,N_17564,N_17833);
nand U18392 (N_18392,N_17495,N_17137);
and U18393 (N_18393,N_17476,N_17456);
nand U18394 (N_18394,N_17375,N_17623);
nand U18395 (N_18395,N_17967,N_17896);
nor U18396 (N_18396,N_17286,N_17998);
and U18397 (N_18397,N_17440,N_17504);
xor U18398 (N_18398,N_17804,N_17740);
and U18399 (N_18399,N_17222,N_17741);
nand U18400 (N_18400,N_17982,N_17426);
xnor U18401 (N_18401,N_17990,N_17391);
nand U18402 (N_18402,N_17049,N_17411);
or U18403 (N_18403,N_17120,N_17390);
xor U18404 (N_18404,N_17902,N_17330);
nand U18405 (N_18405,N_17161,N_17484);
and U18406 (N_18406,N_17619,N_17125);
and U18407 (N_18407,N_17909,N_17817);
nand U18408 (N_18408,N_17075,N_17863);
and U18409 (N_18409,N_17583,N_17897);
nor U18410 (N_18410,N_17667,N_17323);
xor U18411 (N_18411,N_17696,N_17828);
nand U18412 (N_18412,N_17384,N_17008);
or U18413 (N_18413,N_17871,N_17639);
and U18414 (N_18414,N_17859,N_17509);
and U18415 (N_18415,N_17953,N_17342);
and U18416 (N_18416,N_17344,N_17675);
xnor U18417 (N_18417,N_17291,N_17935);
or U18418 (N_18418,N_17635,N_17166);
or U18419 (N_18419,N_17845,N_17736);
nor U18420 (N_18420,N_17345,N_17530);
or U18421 (N_18421,N_17574,N_17409);
xor U18422 (N_18422,N_17088,N_17584);
and U18423 (N_18423,N_17555,N_17221);
nor U18424 (N_18424,N_17293,N_17107);
or U18425 (N_18425,N_17899,N_17450);
and U18426 (N_18426,N_17640,N_17307);
nor U18427 (N_18427,N_17984,N_17038);
xnor U18428 (N_18428,N_17207,N_17838);
or U18429 (N_18429,N_17550,N_17540);
and U18430 (N_18430,N_17737,N_17755);
nand U18431 (N_18431,N_17556,N_17943);
and U18432 (N_18432,N_17357,N_17856);
xor U18433 (N_18433,N_17533,N_17423);
and U18434 (N_18434,N_17581,N_17801);
or U18435 (N_18435,N_17434,N_17582);
nor U18436 (N_18436,N_17392,N_17962);
and U18437 (N_18437,N_17477,N_17247);
nor U18438 (N_18438,N_17603,N_17251);
nor U18439 (N_18439,N_17256,N_17271);
nor U18440 (N_18440,N_17433,N_17109);
or U18441 (N_18441,N_17406,N_17917);
or U18442 (N_18442,N_17654,N_17731);
or U18443 (N_18443,N_17227,N_17128);
nand U18444 (N_18444,N_17611,N_17794);
nor U18445 (N_18445,N_17854,N_17599);
xnor U18446 (N_18446,N_17508,N_17750);
nor U18447 (N_18447,N_17496,N_17325);
and U18448 (N_18448,N_17469,N_17646);
nand U18449 (N_18449,N_17326,N_17743);
and U18450 (N_18450,N_17317,N_17244);
xnor U18451 (N_18451,N_17035,N_17405);
nand U18452 (N_18452,N_17946,N_17554);
and U18453 (N_18453,N_17197,N_17761);
nand U18454 (N_18454,N_17673,N_17904);
and U18455 (N_18455,N_17717,N_17716);
nand U18456 (N_18456,N_17388,N_17289);
nand U18457 (N_18457,N_17427,N_17144);
or U18458 (N_18458,N_17738,N_17382);
nor U18459 (N_18459,N_17341,N_17070);
nand U18460 (N_18460,N_17301,N_17822);
or U18461 (N_18461,N_17653,N_17586);
nand U18462 (N_18462,N_17647,N_17837);
xor U18463 (N_18463,N_17324,N_17730);
xnor U18464 (N_18464,N_17764,N_17478);
nor U18465 (N_18465,N_17615,N_17913);
and U18466 (N_18466,N_17046,N_17377);
or U18467 (N_18467,N_17416,N_17772);
nand U18468 (N_18468,N_17760,N_17656);
nand U18469 (N_18469,N_17215,N_17779);
or U18470 (N_18470,N_17011,N_17945);
nor U18471 (N_18471,N_17965,N_17368);
nor U18472 (N_18472,N_17959,N_17784);
or U18473 (N_18473,N_17020,N_17638);
xor U18474 (N_18474,N_17135,N_17053);
and U18475 (N_18475,N_17114,N_17827);
xnor U18476 (N_18476,N_17348,N_17436);
nor U18477 (N_18477,N_17497,N_17703);
nor U18478 (N_18478,N_17036,N_17589);
or U18479 (N_18479,N_17394,N_17610);
or U18480 (N_18480,N_17929,N_17457);
and U18481 (N_18481,N_17722,N_17823);
xnor U18482 (N_18482,N_17757,N_17658);
xnor U18483 (N_18483,N_17985,N_17970);
or U18484 (N_18484,N_17281,N_17211);
nor U18485 (N_18485,N_17580,N_17338);
nor U18486 (N_18486,N_17836,N_17926);
or U18487 (N_18487,N_17452,N_17872);
nor U18488 (N_18488,N_17566,N_17079);
or U18489 (N_18489,N_17299,N_17468);
nand U18490 (N_18490,N_17115,N_17199);
nand U18491 (N_18491,N_17174,N_17246);
xnor U18492 (N_18492,N_17400,N_17561);
nor U18493 (N_18493,N_17818,N_17420);
and U18494 (N_18494,N_17167,N_17071);
and U18495 (N_18495,N_17177,N_17030);
and U18496 (N_18496,N_17714,N_17718);
or U18497 (N_18497,N_17318,N_17378);
xor U18498 (N_18498,N_17894,N_17698);
and U18499 (N_18499,N_17903,N_17387);
xor U18500 (N_18500,N_17136,N_17138);
xnor U18501 (N_18501,N_17704,N_17970);
nor U18502 (N_18502,N_17642,N_17355);
and U18503 (N_18503,N_17006,N_17617);
and U18504 (N_18504,N_17433,N_17560);
nor U18505 (N_18505,N_17446,N_17988);
and U18506 (N_18506,N_17657,N_17130);
nand U18507 (N_18507,N_17157,N_17124);
nor U18508 (N_18508,N_17403,N_17120);
nand U18509 (N_18509,N_17025,N_17845);
and U18510 (N_18510,N_17113,N_17786);
nand U18511 (N_18511,N_17406,N_17977);
nor U18512 (N_18512,N_17700,N_17467);
or U18513 (N_18513,N_17978,N_17171);
and U18514 (N_18514,N_17336,N_17847);
and U18515 (N_18515,N_17775,N_17127);
or U18516 (N_18516,N_17235,N_17038);
xor U18517 (N_18517,N_17893,N_17486);
xnor U18518 (N_18518,N_17773,N_17018);
nand U18519 (N_18519,N_17362,N_17792);
xnor U18520 (N_18520,N_17858,N_17377);
xnor U18521 (N_18521,N_17430,N_17902);
and U18522 (N_18522,N_17155,N_17981);
nand U18523 (N_18523,N_17543,N_17511);
nor U18524 (N_18524,N_17666,N_17928);
xnor U18525 (N_18525,N_17583,N_17372);
or U18526 (N_18526,N_17358,N_17112);
and U18527 (N_18527,N_17047,N_17821);
nor U18528 (N_18528,N_17998,N_17266);
and U18529 (N_18529,N_17331,N_17607);
xnor U18530 (N_18530,N_17964,N_17897);
nor U18531 (N_18531,N_17912,N_17777);
nand U18532 (N_18532,N_17566,N_17859);
nand U18533 (N_18533,N_17931,N_17647);
nor U18534 (N_18534,N_17918,N_17120);
nand U18535 (N_18535,N_17212,N_17824);
and U18536 (N_18536,N_17863,N_17175);
nand U18537 (N_18537,N_17963,N_17250);
nand U18538 (N_18538,N_17666,N_17497);
nand U18539 (N_18539,N_17326,N_17901);
and U18540 (N_18540,N_17329,N_17721);
or U18541 (N_18541,N_17109,N_17691);
nand U18542 (N_18542,N_17406,N_17696);
and U18543 (N_18543,N_17973,N_17530);
or U18544 (N_18544,N_17100,N_17580);
nor U18545 (N_18545,N_17934,N_17767);
or U18546 (N_18546,N_17134,N_17428);
nor U18547 (N_18547,N_17619,N_17269);
xnor U18548 (N_18548,N_17643,N_17883);
nand U18549 (N_18549,N_17412,N_17308);
xor U18550 (N_18550,N_17039,N_17429);
nand U18551 (N_18551,N_17655,N_17376);
nand U18552 (N_18552,N_17311,N_17426);
xnor U18553 (N_18553,N_17545,N_17109);
xnor U18554 (N_18554,N_17562,N_17677);
nand U18555 (N_18555,N_17608,N_17998);
or U18556 (N_18556,N_17749,N_17887);
and U18557 (N_18557,N_17483,N_17209);
xnor U18558 (N_18558,N_17551,N_17450);
and U18559 (N_18559,N_17694,N_17114);
nor U18560 (N_18560,N_17285,N_17517);
nand U18561 (N_18561,N_17409,N_17367);
xor U18562 (N_18562,N_17651,N_17635);
or U18563 (N_18563,N_17513,N_17066);
nand U18564 (N_18564,N_17378,N_17687);
or U18565 (N_18565,N_17684,N_17120);
or U18566 (N_18566,N_17345,N_17009);
and U18567 (N_18567,N_17213,N_17704);
xnor U18568 (N_18568,N_17900,N_17411);
and U18569 (N_18569,N_17713,N_17995);
or U18570 (N_18570,N_17040,N_17935);
nand U18571 (N_18571,N_17518,N_17399);
nor U18572 (N_18572,N_17096,N_17714);
nand U18573 (N_18573,N_17908,N_17412);
and U18574 (N_18574,N_17785,N_17392);
and U18575 (N_18575,N_17877,N_17028);
nand U18576 (N_18576,N_17003,N_17685);
or U18577 (N_18577,N_17035,N_17285);
nand U18578 (N_18578,N_17802,N_17077);
nand U18579 (N_18579,N_17280,N_17993);
or U18580 (N_18580,N_17065,N_17011);
xor U18581 (N_18581,N_17052,N_17098);
xnor U18582 (N_18582,N_17195,N_17679);
nor U18583 (N_18583,N_17709,N_17414);
and U18584 (N_18584,N_17461,N_17940);
xor U18585 (N_18585,N_17219,N_17143);
or U18586 (N_18586,N_17791,N_17956);
or U18587 (N_18587,N_17785,N_17291);
nor U18588 (N_18588,N_17690,N_17645);
nand U18589 (N_18589,N_17556,N_17134);
or U18590 (N_18590,N_17232,N_17884);
nor U18591 (N_18591,N_17584,N_17650);
and U18592 (N_18592,N_17589,N_17248);
xnor U18593 (N_18593,N_17714,N_17227);
nand U18594 (N_18594,N_17680,N_17634);
nand U18595 (N_18595,N_17693,N_17181);
or U18596 (N_18596,N_17065,N_17569);
xor U18597 (N_18597,N_17992,N_17676);
nor U18598 (N_18598,N_17108,N_17619);
and U18599 (N_18599,N_17304,N_17703);
and U18600 (N_18600,N_17474,N_17595);
and U18601 (N_18601,N_17585,N_17943);
nor U18602 (N_18602,N_17840,N_17720);
nor U18603 (N_18603,N_17308,N_17153);
xor U18604 (N_18604,N_17877,N_17409);
xnor U18605 (N_18605,N_17779,N_17332);
and U18606 (N_18606,N_17141,N_17345);
nor U18607 (N_18607,N_17930,N_17827);
and U18608 (N_18608,N_17264,N_17902);
nor U18609 (N_18609,N_17964,N_17838);
or U18610 (N_18610,N_17074,N_17662);
xnor U18611 (N_18611,N_17154,N_17728);
or U18612 (N_18612,N_17657,N_17009);
and U18613 (N_18613,N_17054,N_17679);
nor U18614 (N_18614,N_17287,N_17261);
and U18615 (N_18615,N_17725,N_17955);
xor U18616 (N_18616,N_17860,N_17732);
nand U18617 (N_18617,N_17406,N_17171);
and U18618 (N_18618,N_17561,N_17560);
and U18619 (N_18619,N_17375,N_17606);
nand U18620 (N_18620,N_17096,N_17549);
nor U18621 (N_18621,N_17804,N_17528);
or U18622 (N_18622,N_17494,N_17121);
and U18623 (N_18623,N_17249,N_17191);
or U18624 (N_18624,N_17283,N_17049);
nand U18625 (N_18625,N_17564,N_17881);
xnor U18626 (N_18626,N_17525,N_17887);
or U18627 (N_18627,N_17834,N_17446);
xnor U18628 (N_18628,N_17566,N_17866);
nor U18629 (N_18629,N_17093,N_17424);
xor U18630 (N_18630,N_17626,N_17049);
xnor U18631 (N_18631,N_17003,N_17311);
and U18632 (N_18632,N_17392,N_17996);
xor U18633 (N_18633,N_17251,N_17142);
nor U18634 (N_18634,N_17070,N_17381);
and U18635 (N_18635,N_17341,N_17606);
and U18636 (N_18636,N_17736,N_17654);
and U18637 (N_18637,N_17852,N_17304);
nand U18638 (N_18638,N_17685,N_17956);
nor U18639 (N_18639,N_17528,N_17964);
and U18640 (N_18640,N_17981,N_17128);
and U18641 (N_18641,N_17588,N_17916);
and U18642 (N_18642,N_17242,N_17619);
and U18643 (N_18643,N_17279,N_17461);
nor U18644 (N_18644,N_17524,N_17047);
and U18645 (N_18645,N_17500,N_17738);
nor U18646 (N_18646,N_17085,N_17997);
nor U18647 (N_18647,N_17048,N_17418);
nand U18648 (N_18648,N_17192,N_17963);
and U18649 (N_18649,N_17453,N_17229);
xor U18650 (N_18650,N_17370,N_17989);
and U18651 (N_18651,N_17319,N_17844);
nand U18652 (N_18652,N_17440,N_17200);
or U18653 (N_18653,N_17165,N_17366);
nand U18654 (N_18654,N_17899,N_17011);
nor U18655 (N_18655,N_17678,N_17634);
and U18656 (N_18656,N_17293,N_17302);
and U18657 (N_18657,N_17177,N_17610);
nand U18658 (N_18658,N_17028,N_17422);
nand U18659 (N_18659,N_17272,N_17905);
nor U18660 (N_18660,N_17638,N_17517);
xnor U18661 (N_18661,N_17890,N_17192);
nor U18662 (N_18662,N_17112,N_17769);
or U18663 (N_18663,N_17904,N_17170);
and U18664 (N_18664,N_17507,N_17375);
nor U18665 (N_18665,N_17155,N_17431);
xor U18666 (N_18666,N_17654,N_17146);
or U18667 (N_18667,N_17618,N_17779);
and U18668 (N_18668,N_17272,N_17575);
nand U18669 (N_18669,N_17716,N_17682);
or U18670 (N_18670,N_17002,N_17862);
xor U18671 (N_18671,N_17852,N_17844);
nor U18672 (N_18672,N_17539,N_17068);
xor U18673 (N_18673,N_17308,N_17073);
xor U18674 (N_18674,N_17384,N_17172);
xnor U18675 (N_18675,N_17659,N_17722);
nor U18676 (N_18676,N_17990,N_17498);
xnor U18677 (N_18677,N_17109,N_17681);
nand U18678 (N_18678,N_17188,N_17408);
nand U18679 (N_18679,N_17700,N_17955);
nand U18680 (N_18680,N_17549,N_17394);
and U18681 (N_18681,N_17028,N_17793);
nor U18682 (N_18682,N_17928,N_17463);
xnor U18683 (N_18683,N_17710,N_17691);
xnor U18684 (N_18684,N_17144,N_17445);
nor U18685 (N_18685,N_17206,N_17866);
and U18686 (N_18686,N_17170,N_17844);
and U18687 (N_18687,N_17885,N_17496);
and U18688 (N_18688,N_17177,N_17855);
nor U18689 (N_18689,N_17422,N_17201);
nor U18690 (N_18690,N_17563,N_17831);
nor U18691 (N_18691,N_17777,N_17679);
nor U18692 (N_18692,N_17358,N_17694);
or U18693 (N_18693,N_17153,N_17993);
nor U18694 (N_18694,N_17422,N_17716);
nor U18695 (N_18695,N_17282,N_17220);
nand U18696 (N_18696,N_17158,N_17376);
or U18697 (N_18697,N_17449,N_17712);
and U18698 (N_18698,N_17448,N_17938);
xor U18699 (N_18699,N_17263,N_17809);
xnor U18700 (N_18700,N_17923,N_17759);
and U18701 (N_18701,N_17725,N_17941);
nand U18702 (N_18702,N_17509,N_17052);
nand U18703 (N_18703,N_17102,N_17214);
nand U18704 (N_18704,N_17017,N_17494);
nand U18705 (N_18705,N_17166,N_17763);
xnor U18706 (N_18706,N_17586,N_17456);
nand U18707 (N_18707,N_17757,N_17730);
or U18708 (N_18708,N_17582,N_17285);
nand U18709 (N_18709,N_17738,N_17209);
nor U18710 (N_18710,N_17264,N_17978);
nor U18711 (N_18711,N_17569,N_17535);
or U18712 (N_18712,N_17507,N_17024);
xnor U18713 (N_18713,N_17685,N_17410);
or U18714 (N_18714,N_17339,N_17417);
nand U18715 (N_18715,N_17910,N_17474);
xor U18716 (N_18716,N_17775,N_17719);
xor U18717 (N_18717,N_17000,N_17642);
or U18718 (N_18718,N_17632,N_17905);
nor U18719 (N_18719,N_17532,N_17369);
and U18720 (N_18720,N_17704,N_17632);
and U18721 (N_18721,N_17984,N_17378);
or U18722 (N_18722,N_17910,N_17093);
and U18723 (N_18723,N_17844,N_17959);
nor U18724 (N_18724,N_17163,N_17128);
and U18725 (N_18725,N_17040,N_17940);
xor U18726 (N_18726,N_17994,N_17804);
nand U18727 (N_18727,N_17257,N_17460);
nor U18728 (N_18728,N_17818,N_17717);
nor U18729 (N_18729,N_17231,N_17717);
or U18730 (N_18730,N_17688,N_17562);
nand U18731 (N_18731,N_17707,N_17577);
and U18732 (N_18732,N_17518,N_17921);
nand U18733 (N_18733,N_17623,N_17084);
nand U18734 (N_18734,N_17127,N_17629);
or U18735 (N_18735,N_17573,N_17701);
nand U18736 (N_18736,N_17838,N_17589);
xor U18737 (N_18737,N_17976,N_17714);
and U18738 (N_18738,N_17953,N_17329);
and U18739 (N_18739,N_17172,N_17947);
nor U18740 (N_18740,N_17262,N_17935);
nor U18741 (N_18741,N_17532,N_17160);
nor U18742 (N_18742,N_17255,N_17865);
nand U18743 (N_18743,N_17560,N_17040);
nor U18744 (N_18744,N_17537,N_17181);
nand U18745 (N_18745,N_17242,N_17700);
and U18746 (N_18746,N_17189,N_17036);
or U18747 (N_18747,N_17658,N_17623);
nor U18748 (N_18748,N_17485,N_17690);
xor U18749 (N_18749,N_17108,N_17820);
nor U18750 (N_18750,N_17753,N_17472);
xnor U18751 (N_18751,N_17259,N_17502);
and U18752 (N_18752,N_17657,N_17397);
nand U18753 (N_18753,N_17637,N_17007);
or U18754 (N_18754,N_17404,N_17743);
nand U18755 (N_18755,N_17433,N_17866);
nor U18756 (N_18756,N_17093,N_17389);
or U18757 (N_18757,N_17289,N_17990);
and U18758 (N_18758,N_17441,N_17955);
nand U18759 (N_18759,N_17848,N_17772);
or U18760 (N_18760,N_17240,N_17261);
or U18761 (N_18761,N_17693,N_17575);
nor U18762 (N_18762,N_17553,N_17397);
or U18763 (N_18763,N_17545,N_17643);
nor U18764 (N_18764,N_17416,N_17326);
and U18765 (N_18765,N_17794,N_17074);
or U18766 (N_18766,N_17301,N_17650);
nor U18767 (N_18767,N_17850,N_17494);
or U18768 (N_18768,N_17546,N_17734);
or U18769 (N_18769,N_17668,N_17473);
nor U18770 (N_18770,N_17325,N_17715);
nand U18771 (N_18771,N_17626,N_17101);
xnor U18772 (N_18772,N_17556,N_17298);
and U18773 (N_18773,N_17034,N_17508);
nor U18774 (N_18774,N_17265,N_17993);
nand U18775 (N_18775,N_17693,N_17468);
nor U18776 (N_18776,N_17365,N_17520);
or U18777 (N_18777,N_17043,N_17514);
or U18778 (N_18778,N_17479,N_17318);
nand U18779 (N_18779,N_17221,N_17917);
xnor U18780 (N_18780,N_17074,N_17496);
nor U18781 (N_18781,N_17705,N_17365);
xor U18782 (N_18782,N_17484,N_17292);
xor U18783 (N_18783,N_17691,N_17830);
and U18784 (N_18784,N_17553,N_17543);
and U18785 (N_18785,N_17367,N_17426);
or U18786 (N_18786,N_17473,N_17861);
and U18787 (N_18787,N_17219,N_17435);
nor U18788 (N_18788,N_17376,N_17281);
xnor U18789 (N_18789,N_17853,N_17119);
nand U18790 (N_18790,N_17212,N_17716);
xnor U18791 (N_18791,N_17587,N_17053);
nand U18792 (N_18792,N_17307,N_17355);
or U18793 (N_18793,N_17704,N_17344);
xnor U18794 (N_18794,N_17358,N_17869);
nand U18795 (N_18795,N_17855,N_17383);
nand U18796 (N_18796,N_17528,N_17944);
nor U18797 (N_18797,N_17116,N_17844);
xnor U18798 (N_18798,N_17956,N_17697);
xor U18799 (N_18799,N_17971,N_17187);
xor U18800 (N_18800,N_17287,N_17132);
nand U18801 (N_18801,N_17493,N_17444);
nand U18802 (N_18802,N_17510,N_17322);
nor U18803 (N_18803,N_17213,N_17022);
or U18804 (N_18804,N_17005,N_17095);
nand U18805 (N_18805,N_17324,N_17033);
nor U18806 (N_18806,N_17723,N_17724);
nor U18807 (N_18807,N_17664,N_17858);
nor U18808 (N_18808,N_17553,N_17237);
and U18809 (N_18809,N_17365,N_17727);
and U18810 (N_18810,N_17401,N_17806);
nand U18811 (N_18811,N_17022,N_17424);
xnor U18812 (N_18812,N_17052,N_17657);
and U18813 (N_18813,N_17703,N_17519);
nand U18814 (N_18814,N_17127,N_17846);
nand U18815 (N_18815,N_17193,N_17004);
nor U18816 (N_18816,N_17362,N_17842);
and U18817 (N_18817,N_17807,N_17293);
nand U18818 (N_18818,N_17820,N_17802);
nand U18819 (N_18819,N_17027,N_17306);
nor U18820 (N_18820,N_17300,N_17417);
xnor U18821 (N_18821,N_17624,N_17511);
and U18822 (N_18822,N_17720,N_17427);
nor U18823 (N_18823,N_17077,N_17071);
nor U18824 (N_18824,N_17379,N_17752);
nor U18825 (N_18825,N_17540,N_17816);
nor U18826 (N_18826,N_17074,N_17250);
xnor U18827 (N_18827,N_17059,N_17640);
and U18828 (N_18828,N_17135,N_17721);
or U18829 (N_18829,N_17456,N_17812);
or U18830 (N_18830,N_17529,N_17536);
or U18831 (N_18831,N_17401,N_17351);
or U18832 (N_18832,N_17202,N_17421);
nand U18833 (N_18833,N_17284,N_17996);
and U18834 (N_18834,N_17799,N_17954);
xnor U18835 (N_18835,N_17741,N_17761);
nand U18836 (N_18836,N_17774,N_17599);
or U18837 (N_18837,N_17107,N_17978);
nand U18838 (N_18838,N_17258,N_17155);
and U18839 (N_18839,N_17834,N_17959);
or U18840 (N_18840,N_17148,N_17875);
or U18841 (N_18841,N_17525,N_17260);
nand U18842 (N_18842,N_17419,N_17581);
xnor U18843 (N_18843,N_17702,N_17300);
nor U18844 (N_18844,N_17499,N_17072);
xnor U18845 (N_18845,N_17923,N_17137);
or U18846 (N_18846,N_17850,N_17068);
nand U18847 (N_18847,N_17194,N_17376);
nor U18848 (N_18848,N_17611,N_17642);
nor U18849 (N_18849,N_17349,N_17299);
or U18850 (N_18850,N_17641,N_17832);
xnor U18851 (N_18851,N_17439,N_17299);
xnor U18852 (N_18852,N_17455,N_17926);
or U18853 (N_18853,N_17933,N_17824);
nand U18854 (N_18854,N_17168,N_17835);
nor U18855 (N_18855,N_17099,N_17180);
xnor U18856 (N_18856,N_17630,N_17300);
nor U18857 (N_18857,N_17520,N_17861);
nor U18858 (N_18858,N_17541,N_17951);
xnor U18859 (N_18859,N_17839,N_17325);
nand U18860 (N_18860,N_17848,N_17872);
nor U18861 (N_18861,N_17835,N_17428);
and U18862 (N_18862,N_17376,N_17675);
nand U18863 (N_18863,N_17180,N_17038);
nand U18864 (N_18864,N_17991,N_17734);
nor U18865 (N_18865,N_17812,N_17502);
xnor U18866 (N_18866,N_17065,N_17593);
nor U18867 (N_18867,N_17878,N_17448);
nand U18868 (N_18868,N_17533,N_17472);
xor U18869 (N_18869,N_17548,N_17575);
xnor U18870 (N_18870,N_17436,N_17082);
xor U18871 (N_18871,N_17926,N_17046);
and U18872 (N_18872,N_17137,N_17239);
nor U18873 (N_18873,N_17454,N_17077);
nor U18874 (N_18874,N_17931,N_17980);
and U18875 (N_18875,N_17115,N_17425);
and U18876 (N_18876,N_17887,N_17505);
nor U18877 (N_18877,N_17144,N_17046);
nand U18878 (N_18878,N_17627,N_17730);
or U18879 (N_18879,N_17926,N_17325);
xnor U18880 (N_18880,N_17106,N_17758);
nor U18881 (N_18881,N_17885,N_17291);
or U18882 (N_18882,N_17919,N_17734);
and U18883 (N_18883,N_17249,N_17669);
or U18884 (N_18884,N_17379,N_17013);
nor U18885 (N_18885,N_17932,N_17420);
nand U18886 (N_18886,N_17359,N_17213);
and U18887 (N_18887,N_17033,N_17540);
nor U18888 (N_18888,N_17931,N_17741);
and U18889 (N_18889,N_17817,N_17142);
and U18890 (N_18890,N_17461,N_17417);
nor U18891 (N_18891,N_17656,N_17651);
nor U18892 (N_18892,N_17609,N_17832);
nand U18893 (N_18893,N_17742,N_17524);
nand U18894 (N_18894,N_17216,N_17301);
nand U18895 (N_18895,N_17259,N_17446);
and U18896 (N_18896,N_17412,N_17334);
xor U18897 (N_18897,N_17217,N_17654);
or U18898 (N_18898,N_17680,N_17684);
or U18899 (N_18899,N_17557,N_17791);
or U18900 (N_18900,N_17061,N_17143);
or U18901 (N_18901,N_17489,N_17047);
and U18902 (N_18902,N_17876,N_17482);
nor U18903 (N_18903,N_17410,N_17074);
or U18904 (N_18904,N_17600,N_17280);
nor U18905 (N_18905,N_17212,N_17837);
xor U18906 (N_18906,N_17550,N_17669);
nand U18907 (N_18907,N_17872,N_17112);
and U18908 (N_18908,N_17161,N_17515);
xnor U18909 (N_18909,N_17698,N_17649);
or U18910 (N_18910,N_17382,N_17300);
or U18911 (N_18911,N_17394,N_17913);
nor U18912 (N_18912,N_17709,N_17820);
nand U18913 (N_18913,N_17486,N_17242);
or U18914 (N_18914,N_17076,N_17042);
xnor U18915 (N_18915,N_17157,N_17554);
and U18916 (N_18916,N_17414,N_17473);
xor U18917 (N_18917,N_17453,N_17157);
nand U18918 (N_18918,N_17966,N_17275);
and U18919 (N_18919,N_17425,N_17592);
xor U18920 (N_18920,N_17107,N_17843);
nor U18921 (N_18921,N_17201,N_17968);
and U18922 (N_18922,N_17512,N_17037);
nor U18923 (N_18923,N_17658,N_17033);
and U18924 (N_18924,N_17783,N_17635);
nand U18925 (N_18925,N_17413,N_17690);
and U18926 (N_18926,N_17068,N_17801);
or U18927 (N_18927,N_17059,N_17602);
or U18928 (N_18928,N_17890,N_17440);
and U18929 (N_18929,N_17969,N_17583);
nand U18930 (N_18930,N_17535,N_17987);
and U18931 (N_18931,N_17148,N_17522);
or U18932 (N_18932,N_17139,N_17978);
nor U18933 (N_18933,N_17359,N_17411);
or U18934 (N_18934,N_17889,N_17423);
and U18935 (N_18935,N_17916,N_17493);
xor U18936 (N_18936,N_17004,N_17689);
or U18937 (N_18937,N_17601,N_17993);
nand U18938 (N_18938,N_17634,N_17048);
nand U18939 (N_18939,N_17502,N_17469);
nand U18940 (N_18940,N_17661,N_17430);
or U18941 (N_18941,N_17984,N_17773);
and U18942 (N_18942,N_17632,N_17886);
and U18943 (N_18943,N_17414,N_17085);
or U18944 (N_18944,N_17993,N_17564);
and U18945 (N_18945,N_17629,N_17490);
nand U18946 (N_18946,N_17084,N_17762);
nand U18947 (N_18947,N_17893,N_17842);
nand U18948 (N_18948,N_17685,N_17261);
or U18949 (N_18949,N_17291,N_17355);
nor U18950 (N_18950,N_17236,N_17272);
xor U18951 (N_18951,N_17224,N_17931);
and U18952 (N_18952,N_17727,N_17176);
nand U18953 (N_18953,N_17929,N_17736);
nor U18954 (N_18954,N_17375,N_17248);
or U18955 (N_18955,N_17593,N_17596);
xor U18956 (N_18956,N_17455,N_17360);
xnor U18957 (N_18957,N_17842,N_17397);
and U18958 (N_18958,N_17174,N_17922);
nor U18959 (N_18959,N_17108,N_17283);
nand U18960 (N_18960,N_17803,N_17378);
and U18961 (N_18961,N_17432,N_17465);
xor U18962 (N_18962,N_17089,N_17945);
or U18963 (N_18963,N_17344,N_17240);
and U18964 (N_18964,N_17770,N_17866);
xnor U18965 (N_18965,N_17567,N_17426);
nor U18966 (N_18966,N_17451,N_17986);
xnor U18967 (N_18967,N_17226,N_17687);
nor U18968 (N_18968,N_17011,N_17312);
xnor U18969 (N_18969,N_17144,N_17434);
nor U18970 (N_18970,N_17836,N_17666);
xnor U18971 (N_18971,N_17896,N_17400);
xnor U18972 (N_18972,N_17033,N_17876);
xor U18973 (N_18973,N_17478,N_17753);
or U18974 (N_18974,N_17228,N_17159);
nand U18975 (N_18975,N_17099,N_17284);
nand U18976 (N_18976,N_17970,N_17742);
xor U18977 (N_18977,N_17757,N_17173);
nor U18978 (N_18978,N_17927,N_17678);
xor U18979 (N_18979,N_17860,N_17238);
and U18980 (N_18980,N_17356,N_17964);
xor U18981 (N_18981,N_17868,N_17751);
or U18982 (N_18982,N_17953,N_17410);
and U18983 (N_18983,N_17631,N_17688);
and U18984 (N_18984,N_17004,N_17988);
nor U18985 (N_18985,N_17734,N_17105);
xnor U18986 (N_18986,N_17995,N_17721);
and U18987 (N_18987,N_17846,N_17072);
xor U18988 (N_18988,N_17186,N_17169);
and U18989 (N_18989,N_17165,N_17820);
nor U18990 (N_18990,N_17168,N_17358);
nor U18991 (N_18991,N_17144,N_17278);
and U18992 (N_18992,N_17047,N_17851);
nand U18993 (N_18993,N_17216,N_17569);
or U18994 (N_18994,N_17818,N_17289);
and U18995 (N_18995,N_17904,N_17431);
nor U18996 (N_18996,N_17989,N_17980);
nor U18997 (N_18997,N_17915,N_17585);
or U18998 (N_18998,N_17561,N_17004);
xnor U18999 (N_18999,N_17030,N_17792);
nor U19000 (N_19000,N_18689,N_18860);
nor U19001 (N_19001,N_18935,N_18126);
nor U19002 (N_19002,N_18966,N_18088);
and U19003 (N_19003,N_18127,N_18299);
or U19004 (N_19004,N_18749,N_18787);
nand U19005 (N_19005,N_18596,N_18652);
xor U19006 (N_19006,N_18928,N_18727);
xor U19007 (N_19007,N_18188,N_18271);
nand U19008 (N_19008,N_18733,N_18506);
xnor U19009 (N_19009,N_18607,N_18021);
and U19010 (N_19010,N_18960,N_18905);
or U19011 (N_19011,N_18736,N_18943);
xor U19012 (N_19012,N_18405,N_18753);
or U19013 (N_19013,N_18063,N_18359);
or U19014 (N_19014,N_18957,N_18911);
nand U19015 (N_19015,N_18648,N_18149);
nand U19016 (N_19016,N_18082,N_18035);
xnor U19017 (N_19017,N_18544,N_18540);
nor U19018 (N_19018,N_18184,N_18942);
xnor U19019 (N_19019,N_18266,N_18570);
or U19020 (N_19020,N_18442,N_18769);
nor U19021 (N_19021,N_18555,N_18818);
xnor U19022 (N_19022,N_18092,N_18304);
nor U19023 (N_19023,N_18402,N_18142);
xnor U19024 (N_19024,N_18851,N_18739);
nor U19025 (N_19025,N_18763,N_18585);
and U19026 (N_19026,N_18455,N_18183);
and U19027 (N_19027,N_18516,N_18283);
or U19028 (N_19028,N_18210,N_18383);
or U19029 (N_19029,N_18480,N_18887);
nor U19030 (N_19030,N_18899,N_18337);
xor U19031 (N_19031,N_18658,N_18123);
or U19032 (N_19032,N_18421,N_18493);
nand U19033 (N_19033,N_18221,N_18466);
nor U19034 (N_19034,N_18656,N_18364);
or U19035 (N_19035,N_18655,N_18186);
or U19036 (N_19036,N_18545,N_18866);
xor U19037 (N_19037,N_18573,N_18986);
xor U19038 (N_19038,N_18125,N_18370);
nor U19039 (N_19039,N_18216,N_18237);
nand U19040 (N_19040,N_18892,N_18253);
or U19041 (N_19041,N_18504,N_18889);
nor U19042 (N_19042,N_18252,N_18649);
or U19043 (N_19043,N_18885,N_18766);
nor U19044 (N_19044,N_18408,N_18486);
xor U19045 (N_19045,N_18117,N_18489);
nand U19046 (N_19046,N_18050,N_18211);
and U19047 (N_19047,N_18691,N_18446);
and U19048 (N_19048,N_18949,N_18635);
or U19049 (N_19049,N_18313,N_18552);
and U19050 (N_19050,N_18686,N_18803);
xor U19051 (N_19051,N_18098,N_18692);
nand U19052 (N_19052,N_18776,N_18549);
nand U19053 (N_19053,N_18135,N_18386);
or U19054 (N_19054,N_18812,N_18533);
nor U19055 (N_19055,N_18610,N_18565);
nor U19056 (N_19056,N_18815,N_18303);
or U19057 (N_19057,N_18706,N_18109);
nand U19058 (N_19058,N_18679,N_18443);
nor U19059 (N_19059,N_18171,N_18830);
nand U19060 (N_19060,N_18485,N_18512);
or U19061 (N_19061,N_18091,N_18701);
xor U19062 (N_19062,N_18112,N_18064);
and U19063 (N_19063,N_18362,N_18426);
and U19064 (N_19064,N_18180,N_18713);
xnor U19065 (N_19065,N_18385,N_18732);
or U19066 (N_19066,N_18011,N_18754);
or U19067 (N_19067,N_18838,N_18326);
or U19068 (N_19068,N_18714,N_18977);
nand U19069 (N_19069,N_18682,N_18490);
nand U19070 (N_19070,N_18626,N_18620);
or U19071 (N_19071,N_18173,N_18642);
or U19072 (N_19072,N_18995,N_18017);
and U19073 (N_19073,N_18828,N_18287);
and U19074 (N_19074,N_18052,N_18666);
and U19075 (N_19075,N_18105,N_18616);
nand U19076 (N_19076,N_18331,N_18548);
or U19077 (N_19077,N_18841,N_18068);
or U19078 (N_19078,N_18280,N_18735);
nand U19079 (N_19079,N_18872,N_18353);
or U19080 (N_19080,N_18031,N_18244);
xor U19081 (N_19081,N_18576,N_18668);
nor U19082 (N_19082,N_18457,N_18718);
or U19083 (N_19083,N_18118,N_18883);
or U19084 (N_19084,N_18392,N_18030);
xor U19085 (N_19085,N_18414,N_18936);
nor U19086 (N_19086,N_18579,N_18639);
or U19087 (N_19087,N_18508,N_18521);
and U19088 (N_19088,N_18672,N_18792);
nand U19089 (N_19089,N_18859,N_18217);
nand U19090 (N_19090,N_18827,N_18006);
nor U19091 (N_19091,N_18282,N_18798);
xor U19092 (N_19092,N_18605,N_18700);
nor U19093 (N_19093,N_18685,N_18542);
or U19094 (N_19094,N_18973,N_18877);
and U19095 (N_19095,N_18247,N_18268);
nand U19096 (N_19096,N_18144,N_18001);
xnor U19097 (N_19097,N_18155,N_18427);
nor U19098 (N_19098,N_18317,N_18674);
and U19099 (N_19099,N_18444,N_18191);
nor U19100 (N_19100,N_18873,N_18153);
nor U19101 (N_19101,N_18786,N_18846);
or U19102 (N_19102,N_18354,N_18908);
nor U19103 (N_19103,N_18275,N_18474);
nand U19104 (N_19104,N_18238,N_18005);
and U19105 (N_19105,N_18397,N_18433);
and U19106 (N_19106,N_18262,N_18454);
or U19107 (N_19107,N_18192,N_18850);
nor U19108 (N_19108,N_18018,N_18844);
and U19109 (N_19109,N_18968,N_18760);
xor U19110 (N_19110,N_18759,N_18762);
nand U19111 (N_19111,N_18875,N_18650);
or U19112 (N_19112,N_18168,N_18559);
nor U19113 (N_19113,N_18752,N_18723);
nand U19114 (N_19114,N_18496,N_18530);
and U19115 (N_19115,N_18143,N_18581);
xnor U19116 (N_19116,N_18481,N_18611);
or U19117 (N_19117,N_18621,N_18081);
xnor U19118 (N_19118,N_18945,N_18561);
and U19119 (N_19119,N_18265,N_18175);
nor U19120 (N_19120,N_18378,N_18156);
xnor U19121 (N_19121,N_18790,N_18219);
or U19122 (N_19122,N_18865,N_18744);
or U19123 (N_19123,N_18166,N_18694);
or U19124 (N_19124,N_18636,N_18254);
nand U19125 (N_19125,N_18609,N_18748);
nor U19126 (N_19126,N_18467,N_18263);
nor U19127 (N_19127,N_18090,N_18437);
and U19128 (N_19128,N_18348,N_18286);
and U19129 (N_19129,N_18350,N_18106);
nand U19130 (N_19130,N_18222,N_18969);
xnor U19131 (N_19131,N_18661,N_18374);
or U19132 (N_19132,N_18964,N_18808);
nand U19133 (N_19133,N_18071,N_18057);
xnor U19134 (N_19134,N_18821,N_18894);
and U19135 (N_19135,N_18336,N_18886);
nor U19136 (N_19136,N_18400,N_18214);
nand U19137 (N_19137,N_18890,N_18203);
xnor U19138 (N_19138,N_18113,N_18878);
or U19139 (N_19139,N_18854,N_18108);
nand U19140 (N_19140,N_18814,N_18740);
xor U19141 (N_19141,N_18334,N_18205);
nand U19142 (N_19142,N_18750,N_18909);
xor U19143 (N_19143,N_18788,N_18780);
nand U19144 (N_19144,N_18065,N_18462);
nor U19145 (N_19145,N_18432,N_18614);
and U19146 (N_19146,N_18472,N_18600);
xor U19147 (N_19147,N_18435,N_18080);
or U19148 (N_19148,N_18996,N_18807);
xnor U19149 (N_19149,N_18743,N_18460);
and U19150 (N_19150,N_18318,N_18721);
xnor U19151 (N_19151,N_18624,N_18152);
nand U19152 (N_19152,N_18419,N_18925);
or U19153 (N_19153,N_18365,N_18116);
xor U19154 (N_19154,N_18978,N_18665);
nor U19155 (N_19155,N_18917,N_18355);
nor U19156 (N_19156,N_18606,N_18963);
nand U19157 (N_19157,N_18308,N_18861);
or U19158 (N_19158,N_18612,N_18629);
nor U19159 (N_19159,N_18534,N_18796);
nor U19160 (N_19160,N_18046,N_18725);
xnor U19161 (N_19161,N_18536,N_18014);
nand U19162 (N_19162,N_18023,N_18837);
nand U19163 (N_19163,N_18097,N_18741);
nor U19164 (N_19164,N_18670,N_18296);
xor U19165 (N_19165,N_18638,N_18187);
nor U19166 (N_19166,N_18985,N_18589);
xor U19167 (N_19167,N_18857,N_18418);
xor U19168 (N_19168,N_18778,N_18320);
xor U19169 (N_19169,N_18864,N_18915);
and U19170 (N_19170,N_18820,N_18562);
xor U19171 (N_19171,N_18133,N_18458);
nor U19172 (N_19172,N_18468,N_18601);
nor U19173 (N_19173,N_18276,N_18518);
xor U19174 (N_19174,N_18411,N_18901);
nor U19175 (N_19175,N_18715,N_18393);
or U19176 (N_19176,N_18231,N_18045);
nand U19177 (N_19177,N_18382,N_18659);
or U19178 (N_19178,N_18755,N_18728);
and U19179 (N_19179,N_18141,N_18495);
nor U19180 (N_19180,N_18038,N_18479);
and U19181 (N_19181,N_18918,N_18025);
nand U19182 (N_19182,N_18608,N_18880);
or U19183 (N_19183,N_18502,N_18070);
xnor U19184 (N_19184,N_18592,N_18122);
or U19185 (N_19185,N_18974,N_18738);
xnor U19186 (N_19186,N_18944,N_18130);
or U19187 (N_19187,N_18779,N_18197);
and U19188 (N_19188,N_18409,N_18301);
or U19189 (N_19189,N_18557,N_18251);
or U19190 (N_19190,N_18121,N_18722);
or U19191 (N_19191,N_18086,N_18465);
xor U19192 (N_19192,N_18781,N_18055);
xnor U19193 (N_19193,N_18288,N_18363);
xor U19194 (N_19194,N_18644,N_18952);
nor U19195 (N_19195,N_18329,N_18920);
or U19196 (N_19196,N_18871,N_18289);
or U19197 (N_19197,N_18012,N_18069);
nor U19198 (N_19198,N_18954,N_18598);
and U19199 (N_19199,N_18697,N_18200);
nor U19200 (N_19200,N_18501,N_18256);
or U19201 (N_19201,N_18212,N_18574);
nand U19202 (N_19202,N_18994,N_18040);
or U19203 (N_19203,N_18136,N_18563);
or U19204 (N_19204,N_18147,N_18084);
xor U19205 (N_19205,N_18929,N_18583);
or U19206 (N_19206,N_18239,N_18225);
nor U19207 (N_19207,N_18235,N_18770);
nand U19208 (N_19208,N_18855,N_18298);
or U19209 (N_19209,N_18321,N_18119);
nor U19210 (N_19210,N_18330,N_18423);
nand U19211 (N_19211,N_18195,N_18907);
nor U19212 (N_19212,N_18096,N_18167);
and U19213 (N_19213,N_18368,N_18595);
xnor U19214 (N_19214,N_18450,N_18078);
nor U19215 (N_19215,N_18311,N_18525);
nand U19216 (N_19216,N_18164,N_18003);
nand U19217 (N_19217,N_18630,N_18927);
nor U19218 (N_19218,N_18604,N_18281);
xnor U19219 (N_19219,N_18671,N_18028);
nor U19220 (N_19220,N_18083,N_18461);
and U19221 (N_19221,N_18751,N_18295);
or U19222 (N_19222,N_18858,N_18795);
or U19223 (N_19223,N_18930,N_18471);
or U19224 (N_19224,N_18228,N_18441);
nand U19225 (N_19225,N_18588,N_18524);
or U19226 (N_19226,N_18747,N_18341);
xor U19227 (N_19227,N_18874,N_18110);
nand U19228 (N_19228,N_18352,N_18989);
nand U19229 (N_19229,N_18094,N_18292);
or U19230 (N_19230,N_18267,N_18193);
xnor U19231 (N_19231,N_18537,N_18048);
nor U19232 (N_19232,N_18953,N_18734);
xnor U19233 (N_19233,N_18967,N_18279);
and U19234 (N_19234,N_18372,N_18477);
nor U19235 (N_19235,N_18793,N_18440);
and U19236 (N_19236,N_18888,N_18801);
xor U19237 (N_19237,N_18811,N_18004);
nand U19238 (N_19238,N_18500,N_18449);
nand U19239 (N_19239,N_18257,N_18416);
xnor U19240 (N_19240,N_18002,N_18036);
nor U19241 (N_19241,N_18972,N_18297);
xor U19242 (N_19242,N_18229,N_18491);
and U19243 (N_19243,N_18946,N_18622);
nand U19244 (N_19244,N_18120,N_18834);
nor U19245 (N_19245,N_18577,N_18475);
and U19246 (N_19246,N_18509,N_18594);
nand U19247 (N_19247,N_18543,N_18514);
or U19248 (N_19248,N_18213,N_18087);
and U19249 (N_19249,N_18654,N_18438);
nor U19250 (N_19250,N_18428,N_18618);
and U19251 (N_19251,N_18615,N_18805);
nand U19252 (N_19252,N_18241,N_18675);
xnor U19253 (N_19253,N_18938,N_18553);
and U19254 (N_19254,N_18019,N_18358);
and U19255 (N_19255,N_18494,N_18054);
and U19256 (N_19256,N_18148,N_18863);
nand U19257 (N_19257,N_18347,N_18882);
or U19258 (N_19258,N_18342,N_18439);
or U19259 (N_19259,N_18020,N_18146);
xnor U19260 (N_19260,N_18862,N_18037);
nor U19261 (N_19261,N_18349,N_18131);
nor U19262 (N_19262,N_18230,N_18934);
and U19263 (N_19263,N_18218,N_18492);
nor U19264 (N_19264,N_18463,N_18488);
xnor U19265 (N_19265,N_18737,N_18705);
nor U19266 (N_19266,N_18274,N_18729);
and U19267 (N_19267,N_18783,N_18169);
nand U19268 (N_19268,N_18902,N_18129);
nand U19269 (N_19269,N_18599,N_18429);
xnor U19270 (N_19270,N_18224,N_18832);
nand U19271 (N_19271,N_18172,N_18360);
and U19272 (N_19272,N_18631,N_18898);
and U19273 (N_19273,N_18566,N_18822);
nand U19274 (N_19274,N_18584,N_18260);
nand U19275 (N_19275,N_18667,N_18306);
xor U19276 (N_19276,N_18140,N_18401);
nand U19277 (N_19277,N_18922,N_18316);
and U19278 (N_19278,N_18556,N_18663);
xor U19279 (N_19279,N_18993,N_18190);
or U19280 (N_19280,N_18245,N_18194);
or U19281 (N_19281,N_18955,N_18842);
xnor U19282 (N_19282,N_18398,N_18422);
and U19283 (N_19283,N_18357,N_18089);
nor U19284 (N_19284,N_18380,N_18528);
xor U19285 (N_19285,N_18285,N_18939);
and U19286 (N_19286,N_18916,N_18568);
nand U19287 (N_19287,N_18538,N_18387);
nand U19288 (N_19288,N_18951,N_18111);
and U19289 (N_19289,N_18074,N_18132);
or U19290 (N_19290,N_18806,N_18487);
xor U19291 (N_19291,N_18531,N_18325);
and U19292 (N_19292,N_18077,N_18976);
and U19293 (N_19293,N_18425,N_18836);
nor U19294 (N_19294,N_18226,N_18983);
and U19295 (N_19295,N_18731,N_18711);
or U19296 (N_19296,N_18453,N_18043);
and U19297 (N_19297,N_18243,N_18093);
nor U19298 (N_19298,N_18424,N_18702);
or U19299 (N_19299,N_18852,N_18338);
nor U19300 (N_19300,N_18079,N_18719);
or U19301 (N_19301,N_18569,N_18699);
and U19302 (N_19302,N_18114,N_18128);
nand U19303 (N_19303,N_18824,N_18690);
xnor U19304 (N_19304,N_18802,N_18520);
xnor U19305 (N_19305,N_18042,N_18240);
nor U19306 (N_19306,N_18204,N_18376);
nor U19307 (N_19307,N_18027,N_18339);
nand U19308 (N_19308,N_18162,N_18910);
xnor U19309 (N_19309,N_18881,N_18066);
and U19310 (N_19310,N_18513,N_18673);
xor U19311 (N_19311,N_18817,N_18277);
nor U19312 (N_19312,N_18617,N_18154);
or U19313 (N_19313,N_18956,N_18484);
and U19314 (N_19314,N_18948,N_18351);
and U19315 (N_19315,N_18984,N_18469);
nand U19316 (N_19316,N_18703,N_18619);
nand U19317 (N_19317,N_18999,N_18765);
xnor U19318 (N_19318,N_18884,N_18590);
nor U19319 (N_19319,N_18041,N_18305);
nor U19320 (N_19320,N_18101,N_18284);
nor U19321 (N_19321,N_18742,N_18933);
nand U19322 (N_19322,N_18526,N_18293);
or U19323 (N_19323,N_18991,N_18307);
and U19324 (N_19324,N_18451,N_18653);
and U19325 (N_19325,N_18693,N_18373);
and U19326 (N_19326,N_18291,N_18498);
xor U19327 (N_19327,N_18998,N_18896);
or U19328 (N_19328,N_18529,N_18470);
nor U19329 (N_19329,N_18868,N_18067);
or U19330 (N_19330,N_18124,N_18634);
and U19331 (N_19331,N_18764,N_18056);
nand U19332 (N_19332,N_18344,N_18161);
nand U19333 (N_19333,N_18771,N_18895);
nand U19334 (N_19334,N_18234,N_18095);
xor U19335 (N_19335,N_18517,N_18100);
nor U19336 (N_19336,N_18523,N_18051);
xnor U19337 (N_19337,N_18511,N_18452);
nor U19338 (N_19338,N_18535,N_18177);
xnor U19339 (N_19339,N_18085,N_18912);
and U19340 (N_19340,N_18150,N_18328);
and U19341 (N_19341,N_18248,N_18013);
nand U19342 (N_19342,N_18924,N_18677);
nor U19343 (N_19343,N_18761,N_18958);
or U19344 (N_19344,N_18008,N_18179);
and U19345 (N_19345,N_18550,N_18772);
or U19346 (N_19346,N_18399,N_18558);
nor U19347 (N_19347,N_18389,N_18931);
nand U19348 (N_19348,N_18395,N_18637);
and U19349 (N_19349,N_18519,N_18613);
or U19350 (N_19350,N_18499,N_18979);
nor U19351 (N_19351,N_18138,N_18163);
and U19352 (N_19352,N_18029,N_18059);
nand U19353 (N_19353,N_18185,N_18151);
and U19354 (N_19354,N_18597,N_18845);
nand U19355 (N_19355,N_18997,N_18436);
and U19356 (N_19356,N_18209,N_18346);
and U19357 (N_19357,N_18708,N_18914);
nand U19358 (N_19358,N_18273,N_18980);
xor U19359 (N_19359,N_18033,N_18923);
and U19360 (N_19360,N_18073,N_18361);
nor U19361 (N_19361,N_18507,N_18698);
nor U19362 (N_19362,N_18580,N_18810);
nor U19363 (N_19363,N_18809,N_18061);
nand U19364 (N_19364,N_18633,N_18407);
and U19365 (N_19365,N_18024,N_18505);
and U19366 (N_19366,N_18825,N_18181);
or U19367 (N_19367,N_18981,N_18940);
or U19368 (N_19368,N_18319,N_18567);
or U19369 (N_19369,N_18582,N_18391);
nor U19370 (N_19370,N_18522,N_18159);
nor U19371 (N_19371,N_18242,N_18961);
nor U19372 (N_19372,N_18941,N_18593);
nand U19373 (N_19373,N_18249,N_18683);
or U19374 (N_19374,N_18932,N_18641);
or U19375 (N_19375,N_18367,N_18390);
nor U19376 (N_19376,N_18848,N_18062);
nand U19377 (N_19377,N_18867,N_18269);
xor U19378 (N_19378,N_18371,N_18053);
nand U19379 (N_19379,N_18165,N_18756);
xnor U19380 (N_19380,N_18270,N_18145);
nand U19381 (N_19381,N_18410,N_18532);
xnor U19382 (N_19382,N_18332,N_18797);
and U19383 (N_19383,N_18826,N_18049);
nand U19384 (N_19384,N_18227,N_18356);
nor U19385 (N_19385,N_18560,N_18403);
xor U19386 (N_19386,N_18345,N_18785);
or U19387 (N_19387,N_18547,N_18799);
xor U19388 (N_19388,N_18034,N_18704);
nand U19389 (N_19389,N_18831,N_18833);
nor U19390 (N_19390,N_18684,N_18646);
or U19391 (N_19391,N_18250,N_18007);
xor U19392 (N_19392,N_18903,N_18182);
nand U19393 (N_19393,N_18921,N_18724);
and U19394 (N_19394,N_18926,N_18343);
or U19395 (N_19395,N_18775,N_18312);
xnor U19396 (N_19396,N_18541,N_18869);
xnor U19397 (N_19397,N_18379,N_18819);
and U19398 (N_19398,N_18645,N_18076);
or U19399 (N_19399,N_18010,N_18632);
and U19400 (N_19400,N_18746,N_18115);
nor U19401 (N_19401,N_18554,N_18139);
and U19402 (N_19402,N_18420,N_18975);
and U19403 (N_19403,N_18075,N_18678);
nand U19404 (N_19404,N_18134,N_18876);
xnor U19405 (N_19405,N_18539,N_18327);
nand U19406 (N_19406,N_18623,N_18396);
nand U19407 (N_19407,N_18160,N_18625);
or U19408 (N_19408,N_18982,N_18310);
xor U19409 (N_19409,N_18476,N_18794);
or U19410 (N_19410,N_18784,N_18236);
xor U19411 (N_19411,N_18856,N_18664);
nand U19412 (N_19412,N_18816,N_18870);
xor U19413 (N_19413,N_18000,N_18527);
nand U19414 (N_19414,N_18300,N_18891);
xnor U19415 (N_19415,N_18309,N_18434);
xor U19416 (N_19416,N_18431,N_18448);
and U19417 (N_19417,N_18196,N_18107);
and U19418 (N_19418,N_18366,N_18777);
and U19419 (N_19419,N_18515,N_18726);
or U19420 (N_19420,N_18791,N_18680);
nand U19421 (N_19421,N_18510,N_18937);
nor U19422 (N_19422,N_18497,N_18009);
or U19423 (N_19423,N_18959,N_18628);
nor U19424 (N_19424,N_18757,N_18278);
nand U19425 (N_19425,N_18189,N_18322);
or U19426 (N_19426,N_18840,N_18294);
or U19427 (N_19427,N_18464,N_18259);
nor U19428 (N_19428,N_18712,N_18207);
and U19429 (N_19429,N_18551,N_18206);
or U19430 (N_19430,N_18767,N_18710);
and U19431 (N_19431,N_18473,N_18717);
xor U19432 (N_19432,N_18377,N_18290);
xor U19433 (N_19433,N_18962,N_18660);
nor U19434 (N_19434,N_18688,N_18335);
and U19435 (N_19435,N_18662,N_18849);
nand U19436 (N_19436,N_18696,N_18201);
or U19437 (N_19437,N_18415,N_18835);
or U19438 (N_19438,N_18823,N_18789);
xnor U19439 (N_19439,N_18323,N_18044);
nor U19440 (N_19440,N_18261,N_18774);
nor U19441 (N_19441,N_18970,N_18990);
or U19442 (N_19442,N_18178,N_18158);
nor U19443 (N_19443,N_18745,N_18099);
nand U19444 (N_19444,N_18853,N_18022);
nor U19445 (N_19445,N_18170,N_18847);
xor U19446 (N_19446,N_18591,N_18987);
nor U19447 (N_19447,N_18264,N_18215);
and U19448 (N_19448,N_18384,N_18375);
nor U19449 (N_19449,N_18627,N_18758);
and U19450 (N_19450,N_18255,N_18406);
nand U19451 (N_19451,N_18947,N_18208);
nand U19452 (N_19452,N_18103,N_18015);
xor U19453 (N_19453,N_18202,N_18919);
nor U19454 (N_19454,N_18800,N_18950);
and U19455 (N_19455,N_18333,N_18829);
and U19456 (N_19456,N_18369,N_18430);
and U19457 (N_19457,N_18879,N_18174);
nand U19458 (N_19458,N_18246,N_18302);
or U19459 (N_19459,N_18233,N_18546);
and U19460 (N_19460,N_18340,N_18971);
and U19461 (N_19461,N_18483,N_18657);
or U19462 (N_19462,N_18404,N_18564);
nor U19463 (N_19463,N_18478,N_18413);
or U19464 (N_19464,N_18965,N_18768);
and U19465 (N_19465,N_18137,N_18016);
nor U19466 (N_19466,N_18047,N_18388);
xnor U19467 (N_19467,N_18503,N_18104);
or U19468 (N_19468,N_18720,N_18906);
and U19469 (N_19469,N_18893,N_18651);
or U19470 (N_19470,N_18687,N_18447);
nand U19471 (N_19471,N_18586,N_18060);
nor U19472 (N_19472,N_18707,N_18176);
xnor U19473 (N_19473,N_18839,N_18199);
nand U19474 (N_19474,N_18102,N_18032);
nand U19475 (N_19475,N_18904,N_18459);
and U19476 (N_19476,N_18843,N_18602);
and U19477 (N_19477,N_18988,N_18913);
xnor U19478 (N_19478,N_18575,N_18232);
xnor U19479 (N_19479,N_18220,N_18571);
nand U19480 (N_19480,N_18603,N_18804);
and U19481 (N_19481,N_18324,N_18482);
nor U19482 (N_19482,N_18897,N_18394);
or U19483 (N_19483,N_18026,N_18587);
and U19484 (N_19484,N_18315,N_18445);
nand U19485 (N_19485,N_18681,N_18730);
xnor U19486 (N_19486,N_18716,N_18773);
or U19487 (N_19487,N_18412,N_18272);
or U19488 (N_19488,N_18900,N_18417);
and U19489 (N_19489,N_18813,N_18381);
or U19490 (N_19490,N_18157,N_18072);
nand U19491 (N_19491,N_18782,N_18456);
xnor U19492 (N_19492,N_18578,N_18198);
nor U19493 (N_19493,N_18695,N_18643);
or U19494 (N_19494,N_18258,N_18640);
nand U19495 (N_19495,N_18223,N_18314);
or U19496 (N_19496,N_18647,N_18992);
xnor U19497 (N_19497,N_18572,N_18709);
xor U19498 (N_19498,N_18058,N_18669);
nand U19499 (N_19499,N_18676,N_18039);
and U19500 (N_19500,N_18121,N_18400);
xnor U19501 (N_19501,N_18938,N_18732);
or U19502 (N_19502,N_18851,N_18202);
nand U19503 (N_19503,N_18488,N_18979);
or U19504 (N_19504,N_18091,N_18497);
nand U19505 (N_19505,N_18780,N_18108);
or U19506 (N_19506,N_18947,N_18074);
xor U19507 (N_19507,N_18996,N_18773);
and U19508 (N_19508,N_18366,N_18285);
nor U19509 (N_19509,N_18177,N_18615);
and U19510 (N_19510,N_18294,N_18036);
or U19511 (N_19511,N_18616,N_18023);
nand U19512 (N_19512,N_18259,N_18256);
or U19513 (N_19513,N_18409,N_18953);
and U19514 (N_19514,N_18400,N_18958);
nand U19515 (N_19515,N_18611,N_18695);
or U19516 (N_19516,N_18555,N_18705);
xnor U19517 (N_19517,N_18461,N_18493);
nor U19518 (N_19518,N_18076,N_18845);
and U19519 (N_19519,N_18835,N_18474);
nand U19520 (N_19520,N_18273,N_18353);
nor U19521 (N_19521,N_18289,N_18797);
xnor U19522 (N_19522,N_18078,N_18589);
nand U19523 (N_19523,N_18149,N_18696);
nand U19524 (N_19524,N_18494,N_18247);
nand U19525 (N_19525,N_18149,N_18284);
nor U19526 (N_19526,N_18294,N_18206);
nand U19527 (N_19527,N_18382,N_18958);
nor U19528 (N_19528,N_18125,N_18656);
nor U19529 (N_19529,N_18112,N_18926);
or U19530 (N_19530,N_18428,N_18699);
nor U19531 (N_19531,N_18990,N_18317);
nor U19532 (N_19532,N_18774,N_18370);
xnor U19533 (N_19533,N_18651,N_18750);
nor U19534 (N_19534,N_18640,N_18599);
xor U19535 (N_19535,N_18201,N_18874);
or U19536 (N_19536,N_18022,N_18001);
xnor U19537 (N_19537,N_18160,N_18222);
or U19538 (N_19538,N_18470,N_18834);
xnor U19539 (N_19539,N_18412,N_18719);
and U19540 (N_19540,N_18144,N_18825);
nand U19541 (N_19541,N_18146,N_18755);
xor U19542 (N_19542,N_18620,N_18795);
or U19543 (N_19543,N_18173,N_18363);
or U19544 (N_19544,N_18185,N_18600);
nor U19545 (N_19545,N_18640,N_18321);
nor U19546 (N_19546,N_18310,N_18085);
nand U19547 (N_19547,N_18269,N_18109);
or U19548 (N_19548,N_18810,N_18602);
nand U19549 (N_19549,N_18298,N_18997);
and U19550 (N_19550,N_18824,N_18705);
nor U19551 (N_19551,N_18562,N_18389);
nor U19552 (N_19552,N_18958,N_18458);
xnor U19553 (N_19553,N_18912,N_18061);
nor U19554 (N_19554,N_18694,N_18956);
or U19555 (N_19555,N_18125,N_18961);
and U19556 (N_19556,N_18176,N_18265);
or U19557 (N_19557,N_18904,N_18456);
xor U19558 (N_19558,N_18731,N_18957);
xor U19559 (N_19559,N_18695,N_18880);
nor U19560 (N_19560,N_18491,N_18760);
nand U19561 (N_19561,N_18054,N_18097);
nor U19562 (N_19562,N_18201,N_18248);
xor U19563 (N_19563,N_18004,N_18835);
xor U19564 (N_19564,N_18962,N_18768);
nand U19565 (N_19565,N_18568,N_18686);
and U19566 (N_19566,N_18215,N_18565);
nor U19567 (N_19567,N_18675,N_18195);
xnor U19568 (N_19568,N_18514,N_18552);
or U19569 (N_19569,N_18223,N_18953);
and U19570 (N_19570,N_18713,N_18678);
nor U19571 (N_19571,N_18939,N_18240);
nand U19572 (N_19572,N_18135,N_18005);
xnor U19573 (N_19573,N_18698,N_18977);
xor U19574 (N_19574,N_18959,N_18533);
nor U19575 (N_19575,N_18695,N_18520);
xor U19576 (N_19576,N_18974,N_18581);
xnor U19577 (N_19577,N_18906,N_18843);
nand U19578 (N_19578,N_18175,N_18595);
nand U19579 (N_19579,N_18823,N_18230);
nand U19580 (N_19580,N_18947,N_18176);
nand U19581 (N_19581,N_18258,N_18458);
or U19582 (N_19582,N_18943,N_18348);
xnor U19583 (N_19583,N_18276,N_18054);
nand U19584 (N_19584,N_18678,N_18053);
and U19585 (N_19585,N_18432,N_18815);
xor U19586 (N_19586,N_18938,N_18144);
nor U19587 (N_19587,N_18864,N_18459);
or U19588 (N_19588,N_18898,N_18718);
or U19589 (N_19589,N_18949,N_18645);
or U19590 (N_19590,N_18207,N_18862);
nand U19591 (N_19591,N_18363,N_18503);
nand U19592 (N_19592,N_18474,N_18993);
or U19593 (N_19593,N_18261,N_18389);
and U19594 (N_19594,N_18573,N_18397);
nand U19595 (N_19595,N_18727,N_18434);
or U19596 (N_19596,N_18550,N_18382);
or U19597 (N_19597,N_18394,N_18022);
nand U19598 (N_19598,N_18339,N_18560);
and U19599 (N_19599,N_18747,N_18142);
nand U19600 (N_19600,N_18548,N_18629);
and U19601 (N_19601,N_18175,N_18681);
nor U19602 (N_19602,N_18046,N_18224);
xnor U19603 (N_19603,N_18606,N_18172);
nand U19604 (N_19604,N_18229,N_18427);
nor U19605 (N_19605,N_18057,N_18325);
nor U19606 (N_19606,N_18747,N_18538);
xor U19607 (N_19607,N_18625,N_18525);
xnor U19608 (N_19608,N_18983,N_18071);
or U19609 (N_19609,N_18701,N_18410);
and U19610 (N_19610,N_18066,N_18799);
nand U19611 (N_19611,N_18262,N_18567);
nand U19612 (N_19612,N_18550,N_18196);
nand U19613 (N_19613,N_18495,N_18091);
nand U19614 (N_19614,N_18964,N_18302);
nor U19615 (N_19615,N_18681,N_18011);
or U19616 (N_19616,N_18324,N_18149);
and U19617 (N_19617,N_18298,N_18822);
xor U19618 (N_19618,N_18901,N_18401);
xor U19619 (N_19619,N_18056,N_18148);
or U19620 (N_19620,N_18525,N_18100);
xnor U19621 (N_19621,N_18205,N_18949);
xor U19622 (N_19622,N_18427,N_18416);
xnor U19623 (N_19623,N_18259,N_18045);
xor U19624 (N_19624,N_18361,N_18422);
xnor U19625 (N_19625,N_18129,N_18222);
and U19626 (N_19626,N_18590,N_18695);
and U19627 (N_19627,N_18848,N_18891);
or U19628 (N_19628,N_18612,N_18876);
nand U19629 (N_19629,N_18494,N_18051);
nand U19630 (N_19630,N_18965,N_18533);
or U19631 (N_19631,N_18334,N_18617);
nor U19632 (N_19632,N_18986,N_18439);
and U19633 (N_19633,N_18644,N_18020);
xor U19634 (N_19634,N_18824,N_18861);
nor U19635 (N_19635,N_18137,N_18472);
xor U19636 (N_19636,N_18973,N_18017);
nand U19637 (N_19637,N_18115,N_18993);
xor U19638 (N_19638,N_18886,N_18344);
xnor U19639 (N_19639,N_18898,N_18228);
or U19640 (N_19640,N_18598,N_18416);
and U19641 (N_19641,N_18717,N_18805);
and U19642 (N_19642,N_18909,N_18664);
or U19643 (N_19643,N_18550,N_18261);
nor U19644 (N_19644,N_18866,N_18290);
xor U19645 (N_19645,N_18160,N_18390);
and U19646 (N_19646,N_18294,N_18990);
or U19647 (N_19647,N_18821,N_18402);
nor U19648 (N_19648,N_18330,N_18227);
and U19649 (N_19649,N_18741,N_18028);
xnor U19650 (N_19650,N_18060,N_18472);
or U19651 (N_19651,N_18871,N_18998);
nor U19652 (N_19652,N_18291,N_18221);
nand U19653 (N_19653,N_18389,N_18779);
xnor U19654 (N_19654,N_18849,N_18191);
xor U19655 (N_19655,N_18017,N_18621);
and U19656 (N_19656,N_18851,N_18985);
or U19657 (N_19657,N_18981,N_18263);
nand U19658 (N_19658,N_18861,N_18620);
nor U19659 (N_19659,N_18380,N_18634);
xor U19660 (N_19660,N_18889,N_18690);
xnor U19661 (N_19661,N_18200,N_18491);
nor U19662 (N_19662,N_18934,N_18023);
nor U19663 (N_19663,N_18134,N_18522);
nand U19664 (N_19664,N_18137,N_18390);
and U19665 (N_19665,N_18567,N_18161);
xnor U19666 (N_19666,N_18531,N_18608);
xnor U19667 (N_19667,N_18922,N_18089);
xnor U19668 (N_19668,N_18558,N_18724);
nand U19669 (N_19669,N_18646,N_18323);
xnor U19670 (N_19670,N_18739,N_18057);
and U19671 (N_19671,N_18409,N_18507);
nand U19672 (N_19672,N_18358,N_18338);
or U19673 (N_19673,N_18391,N_18979);
nor U19674 (N_19674,N_18819,N_18752);
nand U19675 (N_19675,N_18420,N_18724);
nor U19676 (N_19676,N_18548,N_18562);
or U19677 (N_19677,N_18295,N_18071);
and U19678 (N_19678,N_18588,N_18565);
nand U19679 (N_19679,N_18702,N_18335);
xnor U19680 (N_19680,N_18527,N_18041);
nand U19681 (N_19681,N_18760,N_18101);
and U19682 (N_19682,N_18367,N_18145);
nand U19683 (N_19683,N_18603,N_18370);
nor U19684 (N_19684,N_18501,N_18252);
or U19685 (N_19685,N_18514,N_18364);
nand U19686 (N_19686,N_18898,N_18485);
nand U19687 (N_19687,N_18893,N_18660);
xor U19688 (N_19688,N_18915,N_18682);
and U19689 (N_19689,N_18283,N_18022);
nand U19690 (N_19690,N_18748,N_18494);
and U19691 (N_19691,N_18047,N_18245);
and U19692 (N_19692,N_18354,N_18293);
nand U19693 (N_19693,N_18014,N_18436);
nor U19694 (N_19694,N_18636,N_18213);
nor U19695 (N_19695,N_18469,N_18118);
and U19696 (N_19696,N_18302,N_18452);
xnor U19697 (N_19697,N_18623,N_18233);
xor U19698 (N_19698,N_18154,N_18266);
nor U19699 (N_19699,N_18817,N_18628);
and U19700 (N_19700,N_18378,N_18452);
nand U19701 (N_19701,N_18191,N_18353);
and U19702 (N_19702,N_18335,N_18893);
or U19703 (N_19703,N_18704,N_18631);
xnor U19704 (N_19704,N_18679,N_18406);
nand U19705 (N_19705,N_18343,N_18755);
nor U19706 (N_19706,N_18396,N_18148);
and U19707 (N_19707,N_18295,N_18709);
nand U19708 (N_19708,N_18453,N_18800);
nor U19709 (N_19709,N_18374,N_18965);
xor U19710 (N_19710,N_18562,N_18529);
and U19711 (N_19711,N_18446,N_18049);
nand U19712 (N_19712,N_18659,N_18705);
and U19713 (N_19713,N_18113,N_18634);
or U19714 (N_19714,N_18805,N_18813);
nand U19715 (N_19715,N_18776,N_18662);
nor U19716 (N_19716,N_18228,N_18272);
nand U19717 (N_19717,N_18068,N_18333);
nor U19718 (N_19718,N_18945,N_18997);
nor U19719 (N_19719,N_18837,N_18049);
nand U19720 (N_19720,N_18773,N_18630);
xor U19721 (N_19721,N_18349,N_18996);
or U19722 (N_19722,N_18892,N_18165);
xor U19723 (N_19723,N_18896,N_18852);
or U19724 (N_19724,N_18189,N_18832);
xnor U19725 (N_19725,N_18655,N_18215);
xnor U19726 (N_19726,N_18032,N_18221);
xnor U19727 (N_19727,N_18013,N_18879);
nand U19728 (N_19728,N_18179,N_18122);
xnor U19729 (N_19729,N_18482,N_18288);
nand U19730 (N_19730,N_18779,N_18110);
nand U19731 (N_19731,N_18506,N_18948);
and U19732 (N_19732,N_18523,N_18003);
xnor U19733 (N_19733,N_18623,N_18171);
or U19734 (N_19734,N_18264,N_18424);
and U19735 (N_19735,N_18522,N_18489);
nor U19736 (N_19736,N_18360,N_18422);
nor U19737 (N_19737,N_18219,N_18652);
nor U19738 (N_19738,N_18952,N_18148);
and U19739 (N_19739,N_18425,N_18379);
nand U19740 (N_19740,N_18076,N_18684);
or U19741 (N_19741,N_18089,N_18836);
nand U19742 (N_19742,N_18178,N_18655);
or U19743 (N_19743,N_18532,N_18722);
xor U19744 (N_19744,N_18465,N_18578);
nor U19745 (N_19745,N_18211,N_18951);
nor U19746 (N_19746,N_18129,N_18694);
xor U19747 (N_19747,N_18282,N_18610);
xnor U19748 (N_19748,N_18680,N_18319);
or U19749 (N_19749,N_18451,N_18141);
or U19750 (N_19750,N_18370,N_18555);
nand U19751 (N_19751,N_18503,N_18507);
and U19752 (N_19752,N_18254,N_18701);
nand U19753 (N_19753,N_18532,N_18820);
or U19754 (N_19754,N_18068,N_18310);
xnor U19755 (N_19755,N_18964,N_18166);
nor U19756 (N_19756,N_18067,N_18268);
and U19757 (N_19757,N_18611,N_18265);
xor U19758 (N_19758,N_18309,N_18817);
or U19759 (N_19759,N_18784,N_18147);
nor U19760 (N_19760,N_18036,N_18211);
and U19761 (N_19761,N_18052,N_18990);
nor U19762 (N_19762,N_18796,N_18600);
xor U19763 (N_19763,N_18118,N_18308);
or U19764 (N_19764,N_18815,N_18236);
and U19765 (N_19765,N_18307,N_18410);
nor U19766 (N_19766,N_18095,N_18805);
or U19767 (N_19767,N_18167,N_18499);
nand U19768 (N_19768,N_18131,N_18482);
and U19769 (N_19769,N_18681,N_18127);
xor U19770 (N_19770,N_18854,N_18439);
nor U19771 (N_19771,N_18381,N_18991);
nand U19772 (N_19772,N_18415,N_18619);
or U19773 (N_19773,N_18885,N_18910);
nor U19774 (N_19774,N_18785,N_18683);
nand U19775 (N_19775,N_18537,N_18591);
nand U19776 (N_19776,N_18665,N_18171);
or U19777 (N_19777,N_18337,N_18819);
nor U19778 (N_19778,N_18907,N_18955);
or U19779 (N_19779,N_18099,N_18446);
nand U19780 (N_19780,N_18872,N_18156);
or U19781 (N_19781,N_18556,N_18899);
nor U19782 (N_19782,N_18101,N_18412);
nand U19783 (N_19783,N_18655,N_18258);
nand U19784 (N_19784,N_18172,N_18877);
nor U19785 (N_19785,N_18501,N_18789);
nand U19786 (N_19786,N_18828,N_18203);
xor U19787 (N_19787,N_18990,N_18345);
or U19788 (N_19788,N_18465,N_18610);
xor U19789 (N_19789,N_18983,N_18255);
nor U19790 (N_19790,N_18125,N_18533);
nand U19791 (N_19791,N_18168,N_18353);
and U19792 (N_19792,N_18584,N_18652);
xnor U19793 (N_19793,N_18189,N_18586);
or U19794 (N_19794,N_18015,N_18611);
nor U19795 (N_19795,N_18592,N_18733);
xor U19796 (N_19796,N_18058,N_18610);
nand U19797 (N_19797,N_18883,N_18892);
or U19798 (N_19798,N_18921,N_18352);
xnor U19799 (N_19799,N_18014,N_18049);
and U19800 (N_19800,N_18073,N_18997);
and U19801 (N_19801,N_18665,N_18235);
nor U19802 (N_19802,N_18338,N_18133);
nor U19803 (N_19803,N_18203,N_18957);
and U19804 (N_19804,N_18715,N_18572);
or U19805 (N_19805,N_18961,N_18609);
nand U19806 (N_19806,N_18688,N_18798);
or U19807 (N_19807,N_18985,N_18844);
nand U19808 (N_19808,N_18667,N_18550);
nand U19809 (N_19809,N_18510,N_18224);
nand U19810 (N_19810,N_18634,N_18591);
nand U19811 (N_19811,N_18115,N_18596);
and U19812 (N_19812,N_18482,N_18188);
nand U19813 (N_19813,N_18897,N_18767);
or U19814 (N_19814,N_18000,N_18718);
and U19815 (N_19815,N_18885,N_18268);
nor U19816 (N_19816,N_18467,N_18813);
nor U19817 (N_19817,N_18524,N_18964);
and U19818 (N_19818,N_18482,N_18132);
xnor U19819 (N_19819,N_18302,N_18443);
and U19820 (N_19820,N_18181,N_18602);
nand U19821 (N_19821,N_18257,N_18577);
nand U19822 (N_19822,N_18075,N_18712);
nand U19823 (N_19823,N_18359,N_18973);
or U19824 (N_19824,N_18438,N_18091);
nand U19825 (N_19825,N_18511,N_18192);
or U19826 (N_19826,N_18703,N_18949);
or U19827 (N_19827,N_18039,N_18009);
nand U19828 (N_19828,N_18394,N_18645);
or U19829 (N_19829,N_18339,N_18880);
or U19830 (N_19830,N_18548,N_18056);
or U19831 (N_19831,N_18622,N_18911);
or U19832 (N_19832,N_18091,N_18204);
and U19833 (N_19833,N_18769,N_18398);
xor U19834 (N_19834,N_18885,N_18044);
xnor U19835 (N_19835,N_18299,N_18753);
nand U19836 (N_19836,N_18517,N_18313);
and U19837 (N_19837,N_18106,N_18831);
nand U19838 (N_19838,N_18061,N_18998);
xnor U19839 (N_19839,N_18000,N_18887);
or U19840 (N_19840,N_18841,N_18365);
nor U19841 (N_19841,N_18437,N_18034);
nand U19842 (N_19842,N_18903,N_18682);
or U19843 (N_19843,N_18113,N_18950);
or U19844 (N_19844,N_18592,N_18785);
nand U19845 (N_19845,N_18486,N_18591);
nor U19846 (N_19846,N_18130,N_18807);
nor U19847 (N_19847,N_18716,N_18109);
nor U19848 (N_19848,N_18027,N_18874);
or U19849 (N_19849,N_18578,N_18508);
xnor U19850 (N_19850,N_18104,N_18326);
or U19851 (N_19851,N_18558,N_18436);
or U19852 (N_19852,N_18543,N_18377);
nand U19853 (N_19853,N_18522,N_18414);
or U19854 (N_19854,N_18061,N_18895);
or U19855 (N_19855,N_18966,N_18429);
nand U19856 (N_19856,N_18864,N_18545);
or U19857 (N_19857,N_18888,N_18058);
nand U19858 (N_19858,N_18184,N_18638);
nor U19859 (N_19859,N_18141,N_18013);
or U19860 (N_19860,N_18467,N_18326);
and U19861 (N_19861,N_18280,N_18855);
nand U19862 (N_19862,N_18681,N_18766);
or U19863 (N_19863,N_18842,N_18919);
or U19864 (N_19864,N_18819,N_18062);
xor U19865 (N_19865,N_18320,N_18309);
or U19866 (N_19866,N_18151,N_18429);
and U19867 (N_19867,N_18471,N_18574);
or U19868 (N_19868,N_18289,N_18052);
and U19869 (N_19869,N_18267,N_18479);
nor U19870 (N_19870,N_18916,N_18131);
nand U19871 (N_19871,N_18585,N_18407);
or U19872 (N_19872,N_18874,N_18999);
nand U19873 (N_19873,N_18776,N_18728);
nor U19874 (N_19874,N_18751,N_18216);
nand U19875 (N_19875,N_18002,N_18678);
and U19876 (N_19876,N_18493,N_18641);
nand U19877 (N_19877,N_18836,N_18062);
or U19878 (N_19878,N_18773,N_18588);
nor U19879 (N_19879,N_18168,N_18635);
nand U19880 (N_19880,N_18672,N_18830);
xor U19881 (N_19881,N_18587,N_18644);
nor U19882 (N_19882,N_18781,N_18657);
and U19883 (N_19883,N_18743,N_18172);
or U19884 (N_19884,N_18604,N_18968);
nand U19885 (N_19885,N_18851,N_18735);
and U19886 (N_19886,N_18084,N_18232);
nor U19887 (N_19887,N_18358,N_18139);
and U19888 (N_19888,N_18866,N_18420);
xor U19889 (N_19889,N_18618,N_18256);
and U19890 (N_19890,N_18928,N_18968);
xnor U19891 (N_19891,N_18569,N_18106);
or U19892 (N_19892,N_18533,N_18160);
xor U19893 (N_19893,N_18304,N_18976);
nor U19894 (N_19894,N_18728,N_18071);
xnor U19895 (N_19895,N_18689,N_18815);
or U19896 (N_19896,N_18850,N_18289);
xnor U19897 (N_19897,N_18139,N_18840);
xor U19898 (N_19898,N_18499,N_18592);
xnor U19899 (N_19899,N_18296,N_18399);
and U19900 (N_19900,N_18264,N_18181);
nand U19901 (N_19901,N_18262,N_18696);
nand U19902 (N_19902,N_18622,N_18825);
and U19903 (N_19903,N_18022,N_18280);
xor U19904 (N_19904,N_18893,N_18940);
or U19905 (N_19905,N_18867,N_18514);
nor U19906 (N_19906,N_18893,N_18188);
or U19907 (N_19907,N_18194,N_18022);
xnor U19908 (N_19908,N_18782,N_18945);
xnor U19909 (N_19909,N_18828,N_18930);
and U19910 (N_19910,N_18063,N_18289);
xor U19911 (N_19911,N_18194,N_18344);
nor U19912 (N_19912,N_18611,N_18067);
nor U19913 (N_19913,N_18529,N_18668);
xnor U19914 (N_19914,N_18702,N_18376);
and U19915 (N_19915,N_18817,N_18127);
xor U19916 (N_19916,N_18318,N_18929);
or U19917 (N_19917,N_18587,N_18501);
xor U19918 (N_19918,N_18755,N_18659);
xnor U19919 (N_19919,N_18310,N_18882);
nor U19920 (N_19920,N_18332,N_18778);
xnor U19921 (N_19921,N_18650,N_18579);
or U19922 (N_19922,N_18687,N_18054);
xnor U19923 (N_19923,N_18602,N_18575);
xor U19924 (N_19924,N_18987,N_18897);
nor U19925 (N_19925,N_18662,N_18956);
and U19926 (N_19926,N_18426,N_18249);
and U19927 (N_19927,N_18186,N_18766);
nand U19928 (N_19928,N_18676,N_18012);
nand U19929 (N_19929,N_18321,N_18438);
nor U19930 (N_19930,N_18695,N_18639);
nand U19931 (N_19931,N_18193,N_18793);
or U19932 (N_19932,N_18320,N_18659);
nor U19933 (N_19933,N_18624,N_18506);
and U19934 (N_19934,N_18180,N_18423);
xnor U19935 (N_19935,N_18993,N_18138);
nand U19936 (N_19936,N_18325,N_18552);
nand U19937 (N_19937,N_18502,N_18819);
nand U19938 (N_19938,N_18773,N_18012);
xnor U19939 (N_19939,N_18476,N_18439);
or U19940 (N_19940,N_18492,N_18538);
nor U19941 (N_19941,N_18577,N_18889);
xor U19942 (N_19942,N_18819,N_18498);
and U19943 (N_19943,N_18149,N_18116);
xnor U19944 (N_19944,N_18221,N_18583);
and U19945 (N_19945,N_18736,N_18162);
xnor U19946 (N_19946,N_18130,N_18340);
xor U19947 (N_19947,N_18936,N_18954);
and U19948 (N_19948,N_18141,N_18835);
or U19949 (N_19949,N_18723,N_18011);
nand U19950 (N_19950,N_18355,N_18414);
nand U19951 (N_19951,N_18981,N_18044);
nor U19952 (N_19952,N_18872,N_18779);
or U19953 (N_19953,N_18210,N_18889);
nand U19954 (N_19954,N_18480,N_18116);
nand U19955 (N_19955,N_18599,N_18991);
nor U19956 (N_19956,N_18526,N_18587);
nor U19957 (N_19957,N_18124,N_18457);
nor U19958 (N_19958,N_18900,N_18111);
nor U19959 (N_19959,N_18831,N_18111);
or U19960 (N_19960,N_18943,N_18992);
and U19961 (N_19961,N_18595,N_18051);
or U19962 (N_19962,N_18029,N_18300);
and U19963 (N_19963,N_18260,N_18010);
nand U19964 (N_19964,N_18316,N_18796);
nand U19965 (N_19965,N_18700,N_18637);
xnor U19966 (N_19966,N_18718,N_18986);
nand U19967 (N_19967,N_18595,N_18952);
nand U19968 (N_19968,N_18659,N_18467);
and U19969 (N_19969,N_18237,N_18752);
xor U19970 (N_19970,N_18548,N_18115);
and U19971 (N_19971,N_18484,N_18740);
xnor U19972 (N_19972,N_18958,N_18159);
nand U19973 (N_19973,N_18657,N_18013);
xor U19974 (N_19974,N_18575,N_18936);
nand U19975 (N_19975,N_18938,N_18930);
and U19976 (N_19976,N_18874,N_18162);
nor U19977 (N_19977,N_18940,N_18692);
nor U19978 (N_19978,N_18311,N_18140);
xnor U19979 (N_19979,N_18319,N_18167);
and U19980 (N_19980,N_18992,N_18619);
xnor U19981 (N_19981,N_18933,N_18787);
nand U19982 (N_19982,N_18514,N_18229);
or U19983 (N_19983,N_18075,N_18668);
or U19984 (N_19984,N_18182,N_18303);
xnor U19985 (N_19985,N_18607,N_18957);
and U19986 (N_19986,N_18687,N_18876);
xnor U19987 (N_19987,N_18334,N_18170);
nor U19988 (N_19988,N_18488,N_18969);
nand U19989 (N_19989,N_18609,N_18885);
and U19990 (N_19990,N_18884,N_18700);
nand U19991 (N_19991,N_18163,N_18924);
or U19992 (N_19992,N_18771,N_18266);
xor U19993 (N_19993,N_18210,N_18140);
or U19994 (N_19994,N_18676,N_18892);
xnor U19995 (N_19995,N_18427,N_18619);
nor U19996 (N_19996,N_18081,N_18281);
or U19997 (N_19997,N_18135,N_18263);
nand U19998 (N_19998,N_18832,N_18214);
or U19999 (N_19999,N_18091,N_18601);
or U20000 (N_20000,N_19116,N_19041);
xor U20001 (N_20001,N_19557,N_19595);
and U20002 (N_20002,N_19330,N_19596);
nand U20003 (N_20003,N_19804,N_19807);
xor U20004 (N_20004,N_19609,N_19624);
and U20005 (N_20005,N_19376,N_19813);
nor U20006 (N_20006,N_19738,N_19126);
nor U20007 (N_20007,N_19146,N_19363);
and U20008 (N_20008,N_19823,N_19833);
nor U20009 (N_20009,N_19753,N_19350);
or U20010 (N_20010,N_19638,N_19963);
nor U20011 (N_20011,N_19160,N_19802);
or U20012 (N_20012,N_19108,N_19263);
nor U20013 (N_20013,N_19635,N_19282);
xor U20014 (N_20014,N_19888,N_19106);
nor U20015 (N_20015,N_19852,N_19284);
or U20016 (N_20016,N_19790,N_19630);
and U20017 (N_20017,N_19599,N_19406);
or U20018 (N_20018,N_19837,N_19361);
nand U20019 (N_20019,N_19656,N_19188);
xnor U20020 (N_20020,N_19567,N_19791);
xnor U20021 (N_20021,N_19362,N_19469);
nor U20022 (N_20022,N_19522,N_19054);
and U20023 (N_20023,N_19558,N_19201);
xnor U20024 (N_20024,N_19264,N_19682);
nand U20025 (N_20025,N_19096,N_19409);
or U20026 (N_20026,N_19497,N_19795);
nand U20027 (N_20027,N_19576,N_19371);
xor U20028 (N_20028,N_19826,N_19112);
nor U20029 (N_20029,N_19550,N_19746);
xor U20030 (N_20030,N_19899,N_19944);
nand U20031 (N_20031,N_19989,N_19966);
xor U20032 (N_20032,N_19506,N_19243);
nor U20033 (N_20033,N_19772,N_19326);
xnor U20034 (N_20034,N_19980,N_19815);
or U20035 (N_20035,N_19655,N_19098);
nor U20036 (N_20036,N_19820,N_19461);
or U20037 (N_20037,N_19505,N_19246);
nand U20038 (N_20038,N_19622,N_19265);
nor U20039 (N_20039,N_19117,N_19847);
nand U20040 (N_20040,N_19299,N_19631);
nor U20041 (N_20041,N_19415,N_19431);
or U20042 (N_20042,N_19030,N_19043);
nand U20043 (N_20043,N_19907,N_19977);
nor U20044 (N_20044,N_19306,N_19140);
xnor U20045 (N_20045,N_19370,N_19389);
and U20046 (N_20046,N_19339,N_19173);
nor U20047 (N_20047,N_19968,N_19958);
and U20048 (N_20048,N_19278,N_19249);
xnor U20049 (N_20049,N_19590,N_19592);
xnor U20050 (N_20050,N_19085,N_19903);
and U20051 (N_20051,N_19713,N_19464);
nor U20052 (N_20052,N_19355,N_19620);
xnor U20053 (N_20053,N_19209,N_19070);
and U20054 (N_20054,N_19718,N_19083);
nor U20055 (N_20055,N_19894,N_19741);
xnor U20056 (N_20056,N_19854,N_19318);
or U20057 (N_20057,N_19358,N_19094);
nor U20058 (N_20058,N_19541,N_19955);
nand U20059 (N_20059,N_19102,N_19189);
or U20060 (N_20060,N_19751,N_19923);
nand U20061 (N_20061,N_19392,N_19679);
nand U20062 (N_20062,N_19764,N_19716);
nor U20063 (N_20063,N_19485,N_19100);
nor U20064 (N_20064,N_19953,N_19933);
or U20065 (N_20065,N_19918,N_19077);
xor U20066 (N_20066,N_19231,N_19238);
or U20067 (N_20067,N_19879,N_19237);
or U20068 (N_20068,N_19002,N_19623);
and U20069 (N_20069,N_19875,N_19049);
and U20070 (N_20070,N_19143,N_19474);
and U20071 (N_20071,N_19244,N_19686);
xor U20072 (N_20072,N_19683,N_19781);
or U20073 (N_20073,N_19042,N_19202);
nand U20074 (N_20074,N_19915,N_19033);
nand U20075 (N_20075,N_19147,N_19297);
or U20076 (N_20076,N_19736,N_19827);
xnor U20077 (N_20077,N_19164,N_19908);
or U20078 (N_20078,N_19583,N_19549);
nor U20079 (N_20079,N_19479,N_19774);
nor U20080 (N_20080,N_19521,N_19304);
nor U20081 (N_20081,N_19004,N_19385);
xor U20082 (N_20082,N_19843,N_19695);
xor U20083 (N_20083,N_19706,N_19008);
and U20084 (N_20084,N_19568,N_19593);
nor U20085 (N_20085,N_19196,N_19690);
xor U20086 (N_20086,N_19972,N_19144);
nand U20087 (N_20087,N_19436,N_19612);
nor U20088 (N_20088,N_19769,N_19709);
nand U20089 (N_20089,N_19353,N_19768);
xnor U20090 (N_20090,N_19692,N_19611);
and U20091 (N_20091,N_19867,N_19491);
and U20092 (N_20092,N_19673,N_19207);
or U20093 (N_20093,N_19229,N_19993);
nand U20094 (N_20094,N_19941,N_19783);
xor U20095 (N_20095,N_19806,N_19555);
nand U20096 (N_20096,N_19312,N_19642);
nor U20097 (N_20097,N_19171,N_19562);
nor U20098 (N_20098,N_19494,N_19489);
nor U20099 (N_20099,N_19271,N_19313);
nand U20100 (N_20100,N_19281,N_19535);
nor U20101 (N_20101,N_19051,N_19156);
nor U20102 (N_20102,N_19315,N_19296);
and U20103 (N_20103,N_19165,N_19660);
nor U20104 (N_20104,N_19463,N_19473);
and U20105 (N_20105,N_19861,N_19668);
xnor U20106 (N_20106,N_19180,N_19458);
xor U20107 (N_20107,N_19342,N_19341);
xnor U20108 (N_20108,N_19982,N_19740);
or U20109 (N_20109,N_19708,N_19259);
xor U20110 (N_20110,N_19195,N_19619);
and U20111 (N_20111,N_19857,N_19747);
nor U20112 (N_20112,N_19884,N_19369);
or U20113 (N_20113,N_19752,N_19825);
nor U20114 (N_20114,N_19035,N_19641);
nor U20115 (N_20115,N_19063,N_19031);
xor U20116 (N_20116,N_19137,N_19671);
xor U20117 (N_20117,N_19836,N_19976);
and U20118 (N_20118,N_19771,N_19808);
and U20119 (N_20119,N_19302,N_19443);
nand U20120 (N_20120,N_19516,N_19684);
or U20121 (N_20121,N_19215,N_19074);
nor U20122 (N_20122,N_19667,N_19203);
nor U20123 (N_20123,N_19509,N_19184);
nand U20124 (N_20124,N_19314,N_19733);
xor U20125 (N_20125,N_19168,N_19954);
and U20126 (N_20126,N_19058,N_19013);
and U20127 (N_20127,N_19084,N_19681);
and U20128 (N_20128,N_19710,N_19336);
and U20129 (N_20129,N_19224,N_19761);
nor U20130 (N_20130,N_19909,N_19255);
xor U20131 (N_20131,N_19756,N_19883);
and U20132 (N_20132,N_19187,N_19577);
nand U20133 (N_20133,N_19145,N_19528);
nor U20134 (N_20134,N_19161,N_19998);
xor U20135 (N_20135,N_19556,N_19992);
nand U20136 (N_20136,N_19329,N_19386);
or U20137 (N_20137,N_19366,N_19492);
nand U20138 (N_20138,N_19563,N_19719);
and U20139 (N_20139,N_19864,N_19711);
or U20140 (N_20140,N_19210,N_19166);
nand U20141 (N_20141,N_19014,N_19703);
nor U20142 (N_20142,N_19242,N_19453);
and U20143 (N_20143,N_19354,N_19571);
nand U20144 (N_20144,N_19732,N_19250);
nand U20145 (N_20145,N_19896,N_19338);
or U20146 (N_20146,N_19845,N_19142);
nand U20147 (N_20147,N_19331,N_19649);
or U20148 (N_20148,N_19546,N_19024);
xnor U20149 (N_20149,N_19348,N_19935);
nand U20150 (N_20150,N_19975,N_19637);
or U20151 (N_20151,N_19604,N_19372);
nand U20152 (N_20152,N_19378,N_19865);
nor U20153 (N_20153,N_19948,N_19482);
nand U20154 (N_20154,N_19914,N_19036);
xnor U20155 (N_20155,N_19937,N_19507);
nor U20156 (N_20156,N_19005,N_19529);
nor U20157 (N_20157,N_19470,N_19818);
and U20158 (N_20158,N_19893,N_19261);
and U20159 (N_20159,N_19554,N_19828);
nand U20160 (N_20160,N_19393,N_19892);
and U20161 (N_20161,N_19434,N_19869);
nand U20162 (N_20162,N_19324,N_19456);
xor U20163 (N_20163,N_19407,N_19887);
or U20164 (N_20164,N_19566,N_19585);
and U20165 (N_20165,N_19375,N_19748);
xnor U20166 (N_20166,N_19007,N_19862);
nand U20167 (N_20167,N_19351,N_19524);
nor U20168 (N_20168,N_19979,N_19704);
nor U20169 (N_20169,N_19579,N_19245);
nand U20170 (N_20170,N_19057,N_19841);
and U20171 (N_20171,N_19225,N_19334);
or U20172 (N_20172,N_19107,N_19978);
nand U20173 (N_20173,N_19552,N_19547);
and U20174 (N_20174,N_19186,N_19927);
xor U20175 (N_20175,N_19515,N_19323);
nand U20176 (N_20176,N_19784,N_19427);
or U20177 (N_20177,N_19119,N_19158);
nand U20178 (N_20178,N_19830,N_19122);
nand U20179 (N_20179,N_19542,N_19775);
nand U20180 (N_20180,N_19858,N_19572);
or U20181 (N_20181,N_19512,N_19228);
or U20182 (N_20182,N_19999,N_19866);
nor U20183 (N_20183,N_19066,N_19067);
or U20184 (N_20184,N_19408,N_19253);
nor U20185 (N_20185,N_19471,N_19019);
and U20186 (N_20186,N_19356,N_19367);
nand U20187 (N_20187,N_19834,N_19983);
nand U20188 (N_20188,N_19154,N_19850);
and U20189 (N_20189,N_19310,N_19422);
nor U20190 (N_20190,N_19991,N_19446);
and U20191 (N_20191,N_19454,N_19659);
nand U20192 (N_20192,N_19573,N_19676);
nor U20193 (N_20193,N_19885,N_19621);
xnor U20194 (N_20194,N_19481,N_19969);
nor U20195 (N_20195,N_19678,N_19193);
and U20196 (N_20196,N_19091,N_19429);
xor U20197 (N_20197,N_19928,N_19816);
nor U20198 (N_20198,N_19924,N_19625);
or U20199 (N_20199,N_19000,N_19105);
or U20200 (N_20200,N_19728,N_19787);
or U20201 (N_20201,N_19500,N_19055);
xnor U20202 (N_20202,N_19050,N_19420);
or U20203 (N_20203,N_19234,N_19699);
nand U20204 (N_20204,N_19499,N_19097);
nand U20205 (N_20205,N_19477,N_19696);
and U20206 (N_20206,N_19988,N_19905);
and U20207 (N_20207,N_19486,N_19672);
nand U20208 (N_20208,N_19868,N_19423);
nor U20209 (N_20209,N_19113,N_19459);
or U20210 (N_20210,N_19487,N_19587);
or U20211 (N_20211,N_19260,N_19086);
nand U20212 (N_20212,N_19048,N_19729);
nand U20213 (N_20213,N_19026,N_19110);
and U20214 (N_20214,N_19551,N_19332);
and U20215 (N_20215,N_19922,N_19629);
or U20216 (N_20216,N_19929,N_19380);
nand U20217 (N_20217,N_19151,N_19071);
nand U20218 (N_20218,N_19230,N_19269);
or U20219 (N_20219,N_19859,N_19646);
xor U20220 (N_20220,N_19871,N_19088);
or U20221 (N_20221,N_19608,N_19352);
or U20222 (N_20222,N_19010,N_19029);
xor U20223 (N_20223,N_19449,N_19947);
xnor U20224 (N_20224,N_19942,N_19061);
nand U20225 (N_20225,N_19693,N_19817);
nand U20226 (N_20226,N_19089,N_19803);
nand U20227 (N_20227,N_19020,N_19930);
xnor U20228 (N_20228,N_19603,N_19731);
xnor U20229 (N_20229,N_19200,N_19744);
nor U20230 (N_20230,N_19939,N_19211);
or U20231 (N_20231,N_19799,N_19523);
nand U20232 (N_20232,N_19198,N_19517);
and U20233 (N_20233,N_19068,N_19997);
nand U20234 (N_20234,N_19325,N_19543);
or U20235 (N_20235,N_19131,N_19400);
and U20236 (N_20236,N_19967,N_19322);
or U20237 (N_20237,N_19786,N_19056);
and U20238 (N_20238,N_19971,N_19360);
nor U20239 (N_20239,N_19412,N_19416);
xor U20240 (N_20240,N_19346,N_19654);
nand U20241 (N_20241,N_19586,N_19092);
nor U20242 (N_20242,N_19410,N_19379);
nand U20243 (N_20243,N_19270,N_19123);
xnor U20244 (N_20244,N_19457,N_19961);
and U20245 (N_20245,N_19636,N_19782);
xor U20246 (N_20246,N_19065,N_19616);
or U20247 (N_20247,N_19028,N_19996);
nand U20248 (N_20248,N_19374,N_19870);
or U20249 (N_20249,N_19127,N_19633);
and U20250 (N_20250,N_19974,N_19952);
nand U20251 (N_20251,N_19132,N_19418);
and U20252 (N_20252,N_19093,N_19544);
xnor U20253 (N_20253,N_19344,N_19832);
xor U20254 (N_20254,N_19150,N_19645);
or U20255 (N_20255,N_19037,N_19388);
and U20256 (N_20256,N_19257,N_19938);
nand U20257 (N_20257,N_19789,N_19478);
nor U20258 (N_20258,N_19565,N_19290);
nor U20259 (N_20259,N_19419,N_19588);
and U20260 (N_20260,N_19973,N_19442);
and U20261 (N_20261,N_19570,N_19536);
nor U20262 (N_20262,N_19995,N_19805);
nor U20263 (N_20263,N_19880,N_19949);
or U20264 (N_20264,N_19797,N_19900);
or U20265 (N_20265,N_19185,N_19001);
nand U20266 (N_20266,N_19448,N_19809);
or U20267 (N_20267,N_19222,N_19714);
nor U20268 (N_20268,N_19465,N_19598);
nor U20269 (N_20269,N_19990,N_19793);
nand U20270 (N_20270,N_19040,N_19317);
and U20271 (N_20271,N_19316,N_19812);
nor U20272 (N_20272,N_19428,N_19767);
nand U20273 (N_20273,N_19950,N_19663);
xor U20274 (N_20274,N_19021,N_19440);
or U20275 (N_20275,N_19652,N_19985);
or U20276 (N_20276,N_19776,N_19758);
xnor U20277 (N_20277,N_19569,N_19090);
nor U20278 (N_20278,N_19027,N_19800);
nor U20279 (N_20279,N_19627,N_19666);
or U20280 (N_20280,N_19589,N_19095);
nor U20281 (N_20281,N_19307,N_19513);
nor U20282 (N_20282,N_19175,N_19876);
or U20283 (N_20283,N_19488,N_19006);
xnor U20284 (N_20284,N_19438,N_19578);
and U20285 (N_20285,N_19421,N_19581);
and U20286 (N_20286,N_19911,N_19430);
nand U20287 (N_20287,N_19717,N_19680);
or U20288 (N_20288,N_19722,N_19981);
and U20289 (N_20289,N_19901,N_19136);
xnor U20290 (N_20290,N_19159,N_19677);
and U20291 (N_20291,N_19349,N_19890);
xnor U20292 (N_20292,N_19664,N_19219);
nand U20293 (N_20293,N_19532,N_19226);
xnor U20294 (N_20294,N_19221,N_19182);
nor U20295 (N_20295,N_19130,N_19204);
or U20296 (N_20296,N_19044,N_19912);
or U20297 (N_20297,N_19720,N_19287);
and U20298 (N_20298,N_19294,N_19755);
xor U20299 (N_20299,N_19432,N_19082);
nor U20300 (N_20300,N_19046,N_19076);
and U20301 (N_20301,N_19450,N_19582);
nor U20302 (N_20302,N_19397,N_19594);
or U20303 (N_20303,N_19530,N_19697);
nand U20304 (N_20304,N_19561,N_19754);
nor U20305 (N_20305,N_19032,N_19886);
and U20306 (N_20306,N_19447,N_19519);
xnor U20307 (N_20307,N_19333,N_19653);
or U20308 (N_20308,N_19757,N_19670);
and U20309 (N_20309,N_19648,N_19610);
nor U20310 (N_20310,N_19384,N_19829);
and U20311 (N_20311,N_19181,N_19291);
and U20312 (N_20312,N_19694,N_19335);
nand U20313 (N_20313,N_19468,N_19626);
nor U20314 (N_20314,N_19176,N_19398);
and U20315 (N_20315,N_19538,N_19560);
nor U20316 (N_20316,N_19606,N_19214);
and U20317 (N_20317,N_19936,N_19514);
or U20318 (N_20318,N_19881,N_19233);
xnor U20319 (N_20319,N_19405,N_19467);
and U20320 (N_20320,N_19839,N_19128);
xnor U20321 (N_20321,N_19760,N_19762);
nand U20322 (N_20322,N_19657,N_19658);
xnor U20323 (N_20323,N_19232,N_19258);
and U20324 (N_20324,N_19700,N_19220);
xnor U20325 (N_20325,N_19618,N_19383);
nand U20326 (N_20326,N_19962,N_19526);
and U20327 (N_20327,N_19012,N_19838);
xnor U20328 (N_20328,N_19252,N_19882);
xor U20329 (N_20329,N_19749,N_19502);
nor U20330 (N_20330,N_19853,N_19614);
xnor U20331 (N_20331,N_19039,N_19819);
nor U20332 (N_20332,N_19194,N_19280);
nand U20333 (N_20333,N_19247,N_19466);
and U20334 (N_20334,N_19452,N_19701);
xor U20335 (N_20335,N_19121,N_19129);
nand U20336 (N_20336,N_19511,N_19404);
xor U20337 (N_20337,N_19288,N_19381);
and U20338 (N_20338,N_19064,N_19273);
and U20339 (N_20339,N_19311,N_19080);
xor U20340 (N_20340,N_19213,N_19275);
nor U20341 (N_20341,N_19022,N_19399);
nand U20342 (N_20342,N_19498,N_19135);
xnor U20343 (N_20343,N_19617,N_19347);
nand U20344 (N_20344,N_19277,N_19268);
or U20345 (N_20345,N_19235,N_19591);
and U20346 (N_20346,N_19739,N_19527);
xor U20347 (N_20347,N_19946,N_19015);
nand U20348 (N_20348,N_19889,N_19742);
nand U20349 (N_20349,N_19301,N_19860);
nor U20350 (N_20350,N_19956,N_19357);
or U20351 (N_20351,N_19283,N_19337);
or U20352 (N_20352,N_19345,N_19223);
and U20353 (N_20353,N_19831,N_19778);
and U20354 (N_20354,N_19730,N_19373);
xnor U20355 (N_20355,N_19099,N_19072);
or U20356 (N_20356,N_19639,N_19917);
xnor U20357 (N_20357,N_19038,N_19218);
nor U20358 (N_20358,N_19279,N_19691);
nor U20359 (N_20359,N_19665,N_19661);
xnor U20360 (N_20360,N_19504,N_19208);
and U20361 (N_20361,N_19179,N_19897);
nor U20362 (N_20362,N_19723,N_19874);
nand U20363 (N_20363,N_19824,N_19846);
or U20364 (N_20364,N_19745,N_19003);
and U20365 (N_20365,N_19079,N_19904);
xnor U20366 (N_20366,N_19674,N_19017);
xnor U20367 (N_20367,N_19320,N_19285);
xor U20368 (N_20368,N_19267,N_19062);
nand U20369 (N_20369,N_19548,N_19177);
and U20370 (N_20370,N_19863,N_19564);
and U20371 (N_20371,N_19932,N_19777);
nor U20372 (N_20372,N_19239,N_19364);
and U20373 (N_20373,N_19726,N_19798);
or U20374 (N_20374,N_19075,N_19855);
nor U20375 (N_20375,N_19559,N_19248);
nand U20376 (N_20376,N_19734,N_19125);
and U20377 (N_20377,N_19023,N_19785);
and U20378 (N_20378,N_19715,N_19945);
and U20379 (N_20379,N_19060,N_19687);
xnor U20380 (N_20380,N_19721,N_19272);
and U20381 (N_20381,N_19878,N_19501);
or U20382 (N_20382,N_19286,N_19920);
nand U20383 (N_20383,N_19898,N_19169);
nand U20384 (N_20384,N_19844,N_19327);
or U20385 (N_20385,N_19309,N_19451);
or U20386 (N_20386,N_19134,N_19574);
or U20387 (N_20387,N_19340,N_19835);
or U20388 (N_20388,N_19640,N_19293);
nand U20389 (N_20389,N_19387,N_19120);
and U20390 (N_20390,N_19647,N_19437);
nor U20391 (N_20391,N_19087,N_19750);
and U20392 (N_20392,N_19508,N_19395);
nand U20393 (N_20393,N_19779,N_19197);
nor U20394 (N_20394,N_19227,N_19111);
nor U20395 (N_20395,N_19433,N_19822);
nand U20396 (N_20396,N_19045,N_19382);
or U20397 (N_20397,N_19913,N_19849);
and U20398 (N_20398,N_19476,N_19444);
nor U20399 (N_20399,N_19851,N_19368);
xor U20400 (N_20400,N_19689,N_19483);
nor U20401 (N_20401,N_19462,N_19289);
or U20402 (N_20402,N_19155,N_19240);
and U20403 (N_20403,N_19484,N_19580);
xor U20404 (N_20404,N_19455,N_19951);
or U20405 (N_20405,N_19411,N_19540);
nor U20406 (N_20406,N_19759,N_19401);
nand U20407 (N_20407,N_19216,N_19199);
and U20408 (N_20408,N_19727,N_19052);
or U20409 (N_20409,N_19891,N_19359);
xnor U20410 (N_20410,N_19537,N_19601);
nor U20411 (N_20411,N_19765,N_19178);
and U20412 (N_20412,N_19274,N_19439);
nand U20413 (N_20413,N_19480,N_19531);
xor U20414 (N_20414,N_19262,N_19424);
and U20415 (N_20415,N_19895,N_19931);
xor U20416 (N_20416,N_19906,N_19441);
and U20417 (N_20417,N_19205,N_19069);
nor U20418 (N_20418,N_19669,N_19810);
nand U20419 (N_20419,N_19047,N_19192);
nand U20420 (N_20420,N_19133,N_19959);
nor U20421 (N_20421,N_19493,N_19236);
nor U20422 (N_20422,N_19735,N_19520);
or U20423 (N_20423,N_19725,N_19533);
or U20424 (N_20424,N_19081,N_19644);
and U20425 (N_20425,N_19662,N_19174);
nor U20426 (N_20426,N_19321,N_19943);
xnor U20427 (N_20427,N_19104,N_19510);
nand U20428 (N_20428,N_19413,N_19534);
or U20429 (N_20429,N_19114,N_19600);
and U20430 (N_20430,N_19545,N_19190);
and U20431 (N_20431,N_19821,N_19766);
and U20432 (N_20432,N_19607,N_19584);
nor U20433 (N_20433,N_19016,N_19926);
nand U20434 (N_20434,N_19217,N_19792);
nor U20435 (N_20435,N_19475,N_19149);
xnor U20436 (N_20436,N_19685,N_19212);
and U20437 (N_20437,N_19602,N_19138);
nand U20438 (N_20438,N_19152,N_19934);
or U20439 (N_20439,N_19919,N_19305);
nand U20440 (N_20440,N_19109,N_19018);
or U20441 (N_20441,N_19814,N_19328);
or U20442 (N_20442,N_19796,N_19773);
xnor U20443 (N_20443,N_19396,N_19183);
nand U20444 (N_20444,N_19256,N_19472);
nand U20445 (N_20445,N_19403,N_19402);
and U20446 (N_20446,N_19298,N_19503);
nor U20447 (N_20447,N_19872,N_19254);
nand U20448 (N_20448,N_19994,N_19206);
and U20449 (N_20449,N_19877,N_19780);
nand U20450 (N_20450,N_19241,N_19856);
xnor U20451 (N_20451,N_19251,N_19763);
nand U20452 (N_20452,N_19575,N_19840);
xnor U20453 (N_20453,N_19115,N_19987);
nor U20454 (N_20454,N_19650,N_19634);
or U20455 (N_20455,N_19632,N_19425);
nor U20456 (N_20456,N_19009,N_19391);
or U20457 (N_20457,N_19518,N_19167);
and U20458 (N_20458,N_19414,N_19163);
nor U20459 (N_20459,N_19921,N_19688);
and U20460 (N_20460,N_19794,N_19842);
xnor U20461 (N_20461,N_19539,N_19490);
or U20462 (N_20462,N_19984,N_19525);
xnor U20463 (N_20463,N_19737,N_19319);
xnor U20464 (N_20464,N_19073,N_19011);
nand U20465 (N_20465,N_19675,N_19162);
nor U20466 (N_20466,N_19698,N_19148);
nand U20467 (N_20467,N_19495,N_19276);
and U20468 (N_20468,N_19295,N_19365);
xnor U20469 (N_20469,N_19910,N_19153);
or U20470 (N_20470,N_19377,N_19613);
or U20471 (N_20471,N_19101,N_19390);
and U20472 (N_20472,N_19124,N_19025);
nand U20473 (N_20473,N_19925,N_19615);
nor U20474 (N_20474,N_19902,N_19873);
nand U20475 (N_20475,N_19916,N_19705);
or U20476 (N_20476,N_19770,N_19643);
and U20477 (N_20477,N_19170,N_19426);
nor U20478 (N_20478,N_19605,N_19788);
and U20479 (N_20479,N_19957,N_19811);
and U20480 (N_20480,N_19417,N_19964);
and U20481 (N_20481,N_19435,N_19986);
or U20482 (N_20482,N_19965,N_19724);
or U20483 (N_20483,N_19141,N_19460);
and U20484 (N_20484,N_19053,N_19292);
xnor U20485 (N_20485,N_19103,N_19848);
xor U20486 (N_20486,N_19743,N_19707);
xor U20487 (N_20487,N_19034,N_19300);
or U20488 (N_20488,N_19303,N_19628);
and U20489 (N_20489,N_19308,N_19553);
or U20490 (N_20490,N_19597,N_19651);
and U20491 (N_20491,N_19118,N_19960);
xor U20492 (N_20492,N_19702,N_19078);
nor U20493 (N_20493,N_19496,N_19343);
nor U20494 (N_20494,N_19157,N_19801);
nand U20495 (N_20495,N_19445,N_19940);
or U20496 (N_20496,N_19394,N_19191);
or U20497 (N_20497,N_19139,N_19172);
xnor U20498 (N_20498,N_19059,N_19970);
xnor U20499 (N_20499,N_19266,N_19712);
and U20500 (N_20500,N_19983,N_19756);
and U20501 (N_20501,N_19959,N_19626);
and U20502 (N_20502,N_19852,N_19890);
and U20503 (N_20503,N_19496,N_19461);
or U20504 (N_20504,N_19062,N_19066);
xnor U20505 (N_20505,N_19528,N_19269);
nor U20506 (N_20506,N_19301,N_19700);
nand U20507 (N_20507,N_19686,N_19773);
nand U20508 (N_20508,N_19090,N_19930);
xor U20509 (N_20509,N_19939,N_19840);
nor U20510 (N_20510,N_19440,N_19494);
nor U20511 (N_20511,N_19726,N_19514);
nand U20512 (N_20512,N_19225,N_19589);
xnor U20513 (N_20513,N_19783,N_19949);
or U20514 (N_20514,N_19015,N_19417);
and U20515 (N_20515,N_19618,N_19439);
or U20516 (N_20516,N_19795,N_19024);
xor U20517 (N_20517,N_19690,N_19193);
and U20518 (N_20518,N_19606,N_19771);
or U20519 (N_20519,N_19478,N_19710);
and U20520 (N_20520,N_19032,N_19429);
xor U20521 (N_20521,N_19211,N_19926);
nand U20522 (N_20522,N_19589,N_19662);
xor U20523 (N_20523,N_19133,N_19678);
nor U20524 (N_20524,N_19045,N_19364);
xnor U20525 (N_20525,N_19140,N_19577);
xor U20526 (N_20526,N_19773,N_19555);
and U20527 (N_20527,N_19979,N_19269);
or U20528 (N_20528,N_19668,N_19630);
and U20529 (N_20529,N_19868,N_19320);
nand U20530 (N_20530,N_19350,N_19401);
nor U20531 (N_20531,N_19817,N_19315);
xnor U20532 (N_20532,N_19297,N_19652);
or U20533 (N_20533,N_19625,N_19864);
or U20534 (N_20534,N_19325,N_19697);
nand U20535 (N_20535,N_19175,N_19924);
nand U20536 (N_20536,N_19013,N_19338);
nor U20537 (N_20537,N_19977,N_19311);
or U20538 (N_20538,N_19979,N_19031);
nand U20539 (N_20539,N_19941,N_19287);
nor U20540 (N_20540,N_19242,N_19611);
or U20541 (N_20541,N_19267,N_19598);
nand U20542 (N_20542,N_19142,N_19289);
or U20543 (N_20543,N_19802,N_19603);
xor U20544 (N_20544,N_19305,N_19945);
and U20545 (N_20545,N_19892,N_19460);
and U20546 (N_20546,N_19029,N_19995);
nor U20547 (N_20547,N_19583,N_19332);
nor U20548 (N_20548,N_19620,N_19802);
xor U20549 (N_20549,N_19919,N_19710);
and U20550 (N_20550,N_19980,N_19707);
or U20551 (N_20551,N_19068,N_19866);
or U20552 (N_20552,N_19845,N_19668);
nand U20553 (N_20553,N_19759,N_19854);
or U20554 (N_20554,N_19465,N_19258);
nor U20555 (N_20555,N_19763,N_19962);
xnor U20556 (N_20556,N_19350,N_19442);
xnor U20557 (N_20557,N_19066,N_19519);
nand U20558 (N_20558,N_19794,N_19223);
nor U20559 (N_20559,N_19096,N_19796);
nor U20560 (N_20560,N_19634,N_19312);
and U20561 (N_20561,N_19893,N_19783);
nand U20562 (N_20562,N_19854,N_19324);
or U20563 (N_20563,N_19402,N_19220);
nand U20564 (N_20564,N_19631,N_19900);
or U20565 (N_20565,N_19530,N_19466);
and U20566 (N_20566,N_19352,N_19714);
nand U20567 (N_20567,N_19045,N_19661);
or U20568 (N_20568,N_19516,N_19720);
xor U20569 (N_20569,N_19000,N_19202);
and U20570 (N_20570,N_19794,N_19578);
nor U20571 (N_20571,N_19865,N_19987);
nor U20572 (N_20572,N_19232,N_19299);
nand U20573 (N_20573,N_19054,N_19744);
nor U20574 (N_20574,N_19671,N_19585);
xor U20575 (N_20575,N_19378,N_19392);
or U20576 (N_20576,N_19583,N_19764);
xnor U20577 (N_20577,N_19595,N_19672);
or U20578 (N_20578,N_19656,N_19088);
nor U20579 (N_20579,N_19166,N_19470);
nand U20580 (N_20580,N_19620,N_19680);
xnor U20581 (N_20581,N_19317,N_19580);
nand U20582 (N_20582,N_19495,N_19804);
nand U20583 (N_20583,N_19518,N_19338);
xor U20584 (N_20584,N_19561,N_19372);
nor U20585 (N_20585,N_19333,N_19607);
nor U20586 (N_20586,N_19264,N_19987);
nand U20587 (N_20587,N_19171,N_19415);
nor U20588 (N_20588,N_19773,N_19177);
xnor U20589 (N_20589,N_19936,N_19232);
xnor U20590 (N_20590,N_19271,N_19072);
and U20591 (N_20591,N_19500,N_19639);
or U20592 (N_20592,N_19229,N_19061);
and U20593 (N_20593,N_19937,N_19002);
or U20594 (N_20594,N_19098,N_19504);
nor U20595 (N_20595,N_19199,N_19256);
or U20596 (N_20596,N_19417,N_19384);
xor U20597 (N_20597,N_19379,N_19005);
xnor U20598 (N_20598,N_19668,N_19921);
nor U20599 (N_20599,N_19282,N_19746);
nor U20600 (N_20600,N_19959,N_19058);
nand U20601 (N_20601,N_19390,N_19475);
xnor U20602 (N_20602,N_19316,N_19532);
and U20603 (N_20603,N_19950,N_19737);
or U20604 (N_20604,N_19601,N_19541);
xnor U20605 (N_20605,N_19304,N_19563);
and U20606 (N_20606,N_19649,N_19080);
xor U20607 (N_20607,N_19858,N_19381);
or U20608 (N_20608,N_19262,N_19490);
nor U20609 (N_20609,N_19686,N_19375);
and U20610 (N_20610,N_19019,N_19849);
nand U20611 (N_20611,N_19302,N_19062);
and U20612 (N_20612,N_19502,N_19565);
xnor U20613 (N_20613,N_19245,N_19260);
nand U20614 (N_20614,N_19846,N_19216);
xnor U20615 (N_20615,N_19269,N_19045);
nor U20616 (N_20616,N_19458,N_19966);
nor U20617 (N_20617,N_19331,N_19360);
nand U20618 (N_20618,N_19624,N_19979);
or U20619 (N_20619,N_19058,N_19389);
or U20620 (N_20620,N_19351,N_19633);
nor U20621 (N_20621,N_19499,N_19010);
and U20622 (N_20622,N_19147,N_19153);
and U20623 (N_20623,N_19846,N_19879);
xnor U20624 (N_20624,N_19070,N_19464);
xnor U20625 (N_20625,N_19868,N_19401);
xor U20626 (N_20626,N_19152,N_19445);
and U20627 (N_20627,N_19001,N_19682);
xnor U20628 (N_20628,N_19039,N_19687);
nor U20629 (N_20629,N_19604,N_19686);
xnor U20630 (N_20630,N_19765,N_19188);
nor U20631 (N_20631,N_19941,N_19102);
nand U20632 (N_20632,N_19648,N_19173);
xnor U20633 (N_20633,N_19381,N_19166);
nor U20634 (N_20634,N_19026,N_19903);
nand U20635 (N_20635,N_19401,N_19703);
nand U20636 (N_20636,N_19500,N_19797);
nor U20637 (N_20637,N_19075,N_19377);
or U20638 (N_20638,N_19029,N_19701);
xnor U20639 (N_20639,N_19300,N_19503);
xor U20640 (N_20640,N_19163,N_19055);
nor U20641 (N_20641,N_19533,N_19510);
and U20642 (N_20642,N_19553,N_19671);
nand U20643 (N_20643,N_19966,N_19532);
xnor U20644 (N_20644,N_19478,N_19694);
nand U20645 (N_20645,N_19872,N_19708);
nor U20646 (N_20646,N_19655,N_19506);
xnor U20647 (N_20647,N_19332,N_19220);
xnor U20648 (N_20648,N_19478,N_19470);
xor U20649 (N_20649,N_19421,N_19535);
or U20650 (N_20650,N_19143,N_19101);
nor U20651 (N_20651,N_19134,N_19584);
xnor U20652 (N_20652,N_19512,N_19959);
xor U20653 (N_20653,N_19560,N_19124);
nand U20654 (N_20654,N_19362,N_19254);
nand U20655 (N_20655,N_19939,N_19065);
and U20656 (N_20656,N_19939,N_19476);
xnor U20657 (N_20657,N_19763,N_19916);
nand U20658 (N_20658,N_19821,N_19184);
xnor U20659 (N_20659,N_19716,N_19794);
or U20660 (N_20660,N_19460,N_19555);
nor U20661 (N_20661,N_19787,N_19183);
nand U20662 (N_20662,N_19019,N_19630);
or U20663 (N_20663,N_19035,N_19011);
nand U20664 (N_20664,N_19810,N_19554);
nor U20665 (N_20665,N_19547,N_19335);
nor U20666 (N_20666,N_19882,N_19092);
and U20667 (N_20667,N_19145,N_19069);
or U20668 (N_20668,N_19098,N_19044);
nand U20669 (N_20669,N_19151,N_19492);
nor U20670 (N_20670,N_19093,N_19864);
xnor U20671 (N_20671,N_19902,N_19714);
or U20672 (N_20672,N_19399,N_19665);
nor U20673 (N_20673,N_19101,N_19342);
nor U20674 (N_20674,N_19168,N_19213);
or U20675 (N_20675,N_19207,N_19559);
and U20676 (N_20676,N_19051,N_19549);
xnor U20677 (N_20677,N_19691,N_19962);
and U20678 (N_20678,N_19846,N_19369);
nor U20679 (N_20679,N_19584,N_19284);
xor U20680 (N_20680,N_19779,N_19042);
xnor U20681 (N_20681,N_19221,N_19268);
xor U20682 (N_20682,N_19146,N_19257);
nor U20683 (N_20683,N_19183,N_19158);
and U20684 (N_20684,N_19871,N_19912);
nor U20685 (N_20685,N_19952,N_19116);
xnor U20686 (N_20686,N_19645,N_19744);
nand U20687 (N_20687,N_19982,N_19881);
xor U20688 (N_20688,N_19531,N_19333);
xnor U20689 (N_20689,N_19404,N_19262);
or U20690 (N_20690,N_19933,N_19204);
xnor U20691 (N_20691,N_19845,N_19416);
nor U20692 (N_20692,N_19723,N_19936);
or U20693 (N_20693,N_19300,N_19484);
nand U20694 (N_20694,N_19865,N_19724);
and U20695 (N_20695,N_19878,N_19769);
or U20696 (N_20696,N_19078,N_19805);
nand U20697 (N_20697,N_19851,N_19816);
and U20698 (N_20698,N_19350,N_19334);
xor U20699 (N_20699,N_19125,N_19394);
or U20700 (N_20700,N_19944,N_19951);
nand U20701 (N_20701,N_19969,N_19483);
nor U20702 (N_20702,N_19289,N_19556);
or U20703 (N_20703,N_19225,N_19027);
nand U20704 (N_20704,N_19181,N_19149);
and U20705 (N_20705,N_19335,N_19032);
xnor U20706 (N_20706,N_19330,N_19022);
nand U20707 (N_20707,N_19036,N_19750);
nor U20708 (N_20708,N_19569,N_19330);
or U20709 (N_20709,N_19595,N_19090);
or U20710 (N_20710,N_19323,N_19611);
nor U20711 (N_20711,N_19371,N_19578);
nand U20712 (N_20712,N_19805,N_19923);
or U20713 (N_20713,N_19060,N_19051);
nand U20714 (N_20714,N_19397,N_19207);
nand U20715 (N_20715,N_19483,N_19376);
or U20716 (N_20716,N_19120,N_19719);
or U20717 (N_20717,N_19241,N_19498);
and U20718 (N_20718,N_19948,N_19983);
nand U20719 (N_20719,N_19646,N_19475);
and U20720 (N_20720,N_19533,N_19322);
xor U20721 (N_20721,N_19291,N_19629);
xnor U20722 (N_20722,N_19660,N_19424);
or U20723 (N_20723,N_19619,N_19469);
and U20724 (N_20724,N_19891,N_19190);
xor U20725 (N_20725,N_19283,N_19743);
or U20726 (N_20726,N_19738,N_19220);
and U20727 (N_20727,N_19892,N_19845);
and U20728 (N_20728,N_19311,N_19736);
and U20729 (N_20729,N_19823,N_19456);
nand U20730 (N_20730,N_19549,N_19799);
or U20731 (N_20731,N_19571,N_19504);
xor U20732 (N_20732,N_19476,N_19511);
or U20733 (N_20733,N_19457,N_19175);
nor U20734 (N_20734,N_19664,N_19549);
xnor U20735 (N_20735,N_19763,N_19690);
nand U20736 (N_20736,N_19700,N_19809);
nand U20737 (N_20737,N_19914,N_19864);
and U20738 (N_20738,N_19692,N_19282);
nand U20739 (N_20739,N_19354,N_19277);
nand U20740 (N_20740,N_19237,N_19263);
and U20741 (N_20741,N_19576,N_19461);
and U20742 (N_20742,N_19417,N_19171);
xnor U20743 (N_20743,N_19518,N_19535);
nand U20744 (N_20744,N_19388,N_19918);
nor U20745 (N_20745,N_19071,N_19410);
and U20746 (N_20746,N_19188,N_19732);
nor U20747 (N_20747,N_19514,N_19637);
and U20748 (N_20748,N_19082,N_19503);
nor U20749 (N_20749,N_19138,N_19236);
xor U20750 (N_20750,N_19994,N_19821);
and U20751 (N_20751,N_19360,N_19733);
and U20752 (N_20752,N_19177,N_19551);
or U20753 (N_20753,N_19343,N_19483);
nand U20754 (N_20754,N_19427,N_19435);
xnor U20755 (N_20755,N_19922,N_19059);
xnor U20756 (N_20756,N_19381,N_19074);
xor U20757 (N_20757,N_19462,N_19713);
nor U20758 (N_20758,N_19283,N_19805);
nand U20759 (N_20759,N_19640,N_19236);
nor U20760 (N_20760,N_19624,N_19711);
and U20761 (N_20761,N_19850,N_19322);
nand U20762 (N_20762,N_19602,N_19298);
and U20763 (N_20763,N_19125,N_19872);
nand U20764 (N_20764,N_19336,N_19535);
xnor U20765 (N_20765,N_19902,N_19705);
and U20766 (N_20766,N_19401,N_19887);
xor U20767 (N_20767,N_19934,N_19144);
xor U20768 (N_20768,N_19506,N_19522);
nand U20769 (N_20769,N_19199,N_19858);
nand U20770 (N_20770,N_19073,N_19417);
xor U20771 (N_20771,N_19848,N_19879);
nor U20772 (N_20772,N_19535,N_19841);
nand U20773 (N_20773,N_19318,N_19762);
nor U20774 (N_20774,N_19176,N_19024);
and U20775 (N_20775,N_19194,N_19155);
nor U20776 (N_20776,N_19467,N_19153);
xor U20777 (N_20777,N_19170,N_19858);
and U20778 (N_20778,N_19656,N_19290);
xor U20779 (N_20779,N_19851,N_19211);
nand U20780 (N_20780,N_19378,N_19175);
or U20781 (N_20781,N_19379,N_19404);
and U20782 (N_20782,N_19021,N_19597);
and U20783 (N_20783,N_19938,N_19955);
nand U20784 (N_20784,N_19916,N_19231);
xnor U20785 (N_20785,N_19965,N_19417);
or U20786 (N_20786,N_19867,N_19618);
nand U20787 (N_20787,N_19601,N_19121);
or U20788 (N_20788,N_19097,N_19359);
nand U20789 (N_20789,N_19317,N_19994);
nor U20790 (N_20790,N_19846,N_19828);
and U20791 (N_20791,N_19991,N_19097);
and U20792 (N_20792,N_19162,N_19122);
nor U20793 (N_20793,N_19531,N_19516);
or U20794 (N_20794,N_19642,N_19165);
nor U20795 (N_20795,N_19950,N_19648);
xor U20796 (N_20796,N_19949,N_19523);
xnor U20797 (N_20797,N_19518,N_19962);
xnor U20798 (N_20798,N_19785,N_19090);
or U20799 (N_20799,N_19987,N_19272);
nand U20800 (N_20800,N_19195,N_19684);
or U20801 (N_20801,N_19547,N_19084);
or U20802 (N_20802,N_19534,N_19275);
nor U20803 (N_20803,N_19465,N_19958);
xor U20804 (N_20804,N_19443,N_19409);
and U20805 (N_20805,N_19813,N_19509);
xor U20806 (N_20806,N_19823,N_19596);
nand U20807 (N_20807,N_19749,N_19674);
nand U20808 (N_20808,N_19665,N_19035);
and U20809 (N_20809,N_19691,N_19731);
or U20810 (N_20810,N_19268,N_19753);
or U20811 (N_20811,N_19245,N_19802);
and U20812 (N_20812,N_19313,N_19937);
nor U20813 (N_20813,N_19653,N_19026);
nor U20814 (N_20814,N_19325,N_19127);
xor U20815 (N_20815,N_19187,N_19911);
nand U20816 (N_20816,N_19716,N_19959);
xnor U20817 (N_20817,N_19505,N_19108);
xor U20818 (N_20818,N_19489,N_19528);
or U20819 (N_20819,N_19090,N_19561);
and U20820 (N_20820,N_19016,N_19058);
and U20821 (N_20821,N_19248,N_19427);
nor U20822 (N_20822,N_19948,N_19571);
and U20823 (N_20823,N_19921,N_19776);
nand U20824 (N_20824,N_19967,N_19957);
nor U20825 (N_20825,N_19589,N_19999);
nor U20826 (N_20826,N_19760,N_19829);
and U20827 (N_20827,N_19782,N_19339);
and U20828 (N_20828,N_19819,N_19420);
xor U20829 (N_20829,N_19042,N_19808);
xor U20830 (N_20830,N_19063,N_19159);
nor U20831 (N_20831,N_19137,N_19546);
nor U20832 (N_20832,N_19460,N_19152);
or U20833 (N_20833,N_19782,N_19058);
nor U20834 (N_20834,N_19161,N_19773);
and U20835 (N_20835,N_19642,N_19521);
or U20836 (N_20836,N_19250,N_19728);
xor U20837 (N_20837,N_19706,N_19329);
xor U20838 (N_20838,N_19232,N_19862);
xor U20839 (N_20839,N_19783,N_19573);
nor U20840 (N_20840,N_19784,N_19321);
nand U20841 (N_20841,N_19924,N_19181);
or U20842 (N_20842,N_19989,N_19317);
nor U20843 (N_20843,N_19547,N_19504);
xnor U20844 (N_20844,N_19655,N_19652);
xnor U20845 (N_20845,N_19874,N_19627);
nor U20846 (N_20846,N_19301,N_19432);
xnor U20847 (N_20847,N_19008,N_19444);
or U20848 (N_20848,N_19714,N_19757);
xor U20849 (N_20849,N_19430,N_19719);
and U20850 (N_20850,N_19139,N_19464);
nor U20851 (N_20851,N_19074,N_19646);
xnor U20852 (N_20852,N_19700,N_19433);
xor U20853 (N_20853,N_19260,N_19407);
nor U20854 (N_20854,N_19419,N_19469);
or U20855 (N_20855,N_19720,N_19817);
and U20856 (N_20856,N_19483,N_19965);
xnor U20857 (N_20857,N_19655,N_19046);
xnor U20858 (N_20858,N_19631,N_19858);
or U20859 (N_20859,N_19563,N_19785);
xor U20860 (N_20860,N_19041,N_19776);
or U20861 (N_20861,N_19989,N_19849);
nor U20862 (N_20862,N_19573,N_19543);
xnor U20863 (N_20863,N_19404,N_19324);
nand U20864 (N_20864,N_19159,N_19138);
nand U20865 (N_20865,N_19118,N_19040);
nand U20866 (N_20866,N_19501,N_19516);
nand U20867 (N_20867,N_19807,N_19376);
nor U20868 (N_20868,N_19056,N_19290);
nand U20869 (N_20869,N_19164,N_19489);
nor U20870 (N_20870,N_19508,N_19424);
xor U20871 (N_20871,N_19087,N_19373);
or U20872 (N_20872,N_19406,N_19867);
nor U20873 (N_20873,N_19201,N_19741);
xnor U20874 (N_20874,N_19011,N_19369);
nor U20875 (N_20875,N_19261,N_19565);
xnor U20876 (N_20876,N_19054,N_19917);
and U20877 (N_20877,N_19551,N_19126);
nor U20878 (N_20878,N_19299,N_19015);
xor U20879 (N_20879,N_19458,N_19244);
nor U20880 (N_20880,N_19281,N_19774);
or U20881 (N_20881,N_19894,N_19505);
nand U20882 (N_20882,N_19445,N_19809);
or U20883 (N_20883,N_19328,N_19638);
and U20884 (N_20884,N_19921,N_19605);
and U20885 (N_20885,N_19673,N_19920);
xnor U20886 (N_20886,N_19778,N_19374);
xnor U20887 (N_20887,N_19536,N_19008);
nand U20888 (N_20888,N_19114,N_19206);
and U20889 (N_20889,N_19888,N_19059);
nand U20890 (N_20890,N_19467,N_19245);
or U20891 (N_20891,N_19722,N_19711);
nor U20892 (N_20892,N_19670,N_19198);
or U20893 (N_20893,N_19204,N_19824);
nor U20894 (N_20894,N_19644,N_19306);
xor U20895 (N_20895,N_19318,N_19588);
xor U20896 (N_20896,N_19423,N_19056);
nor U20897 (N_20897,N_19700,N_19936);
or U20898 (N_20898,N_19687,N_19724);
nor U20899 (N_20899,N_19860,N_19552);
nor U20900 (N_20900,N_19132,N_19852);
nor U20901 (N_20901,N_19418,N_19850);
xor U20902 (N_20902,N_19998,N_19061);
nor U20903 (N_20903,N_19831,N_19100);
and U20904 (N_20904,N_19268,N_19925);
nor U20905 (N_20905,N_19743,N_19461);
nand U20906 (N_20906,N_19400,N_19518);
nor U20907 (N_20907,N_19632,N_19232);
or U20908 (N_20908,N_19013,N_19389);
nor U20909 (N_20909,N_19255,N_19405);
nand U20910 (N_20910,N_19036,N_19423);
nand U20911 (N_20911,N_19674,N_19931);
nor U20912 (N_20912,N_19317,N_19351);
or U20913 (N_20913,N_19089,N_19885);
nor U20914 (N_20914,N_19536,N_19537);
nor U20915 (N_20915,N_19134,N_19483);
or U20916 (N_20916,N_19456,N_19758);
xor U20917 (N_20917,N_19307,N_19404);
and U20918 (N_20918,N_19200,N_19905);
nor U20919 (N_20919,N_19263,N_19140);
nand U20920 (N_20920,N_19184,N_19128);
or U20921 (N_20921,N_19097,N_19841);
xor U20922 (N_20922,N_19305,N_19718);
or U20923 (N_20923,N_19473,N_19793);
or U20924 (N_20924,N_19546,N_19365);
and U20925 (N_20925,N_19961,N_19449);
nand U20926 (N_20926,N_19831,N_19575);
xnor U20927 (N_20927,N_19606,N_19391);
nand U20928 (N_20928,N_19619,N_19986);
xor U20929 (N_20929,N_19998,N_19650);
or U20930 (N_20930,N_19612,N_19764);
or U20931 (N_20931,N_19161,N_19618);
nor U20932 (N_20932,N_19932,N_19315);
and U20933 (N_20933,N_19297,N_19063);
xnor U20934 (N_20934,N_19524,N_19451);
and U20935 (N_20935,N_19134,N_19510);
xor U20936 (N_20936,N_19764,N_19711);
xor U20937 (N_20937,N_19333,N_19131);
xnor U20938 (N_20938,N_19888,N_19840);
nor U20939 (N_20939,N_19307,N_19659);
nor U20940 (N_20940,N_19333,N_19829);
nand U20941 (N_20941,N_19883,N_19643);
or U20942 (N_20942,N_19083,N_19189);
nand U20943 (N_20943,N_19001,N_19276);
xnor U20944 (N_20944,N_19046,N_19166);
and U20945 (N_20945,N_19864,N_19373);
and U20946 (N_20946,N_19352,N_19382);
or U20947 (N_20947,N_19789,N_19262);
nor U20948 (N_20948,N_19156,N_19188);
nand U20949 (N_20949,N_19949,N_19823);
xor U20950 (N_20950,N_19804,N_19126);
nor U20951 (N_20951,N_19264,N_19581);
xnor U20952 (N_20952,N_19953,N_19471);
and U20953 (N_20953,N_19420,N_19787);
and U20954 (N_20954,N_19960,N_19827);
xnor U20955 (N_20955,N_19611,N_19249);
nor U20956 (N_20956,N_19774,N_19731);
nor U20957 (N_20957,N_19243,N_19630);
nor U20958 (N_20958,N_19269,N_19518);
and U20959 (N_20959,N_19190,N_19492);
nand U20960 (N_20960,N_19692,N_19064);
nand U20961 (N_20961,N_19962,N_19608);
and U20962 (N_20962,N_19220,N_19749);
and U20963 (N_20963,N_19759,N_19837);
and U20964 (N_20964,N_19414,N_19475);
nor U20965 (N_20965,N_19283,N_19546);
xor U20966 (N_20966,N_19404,N_19574);
nand U20967 (N_20967,N_19786,N_19266);
or U20968 (N_20968,N_19695,N_19234);
xnor U20969 (N_20969,N_19954,N_19299);
nor U20970 (N_20970,N_19039,N_19861);
xor U20971 (N_20971,N_19640,N_19679);
and U20972 (N_20972,N_19051,N_19777);
xor U20973 (N_20973,N_19402,N_19781);
nor U20974 (N_20974,N_19051,N_19920);
and U20975 (N_20975,N_19974,N_19552);
or U20976 (N_20976,N_19872,N_19082);
and U20977 (N_20977,N_19035,N_19784);
nor U20978 (N_20978,N_19248,N_19201);
xnor U20979 (N_20979,N_19850,N_19589);
xor U20980 (N_20980,N_19445,N_19286);
nand U20981 (N_20981,N_19044,N_19376);
nor U20982 (N_20982,N_19079,N_19696);
nand U20983 (N_20983,N_19418,N_19991);
nor U20984 (N_20984,N_19512,N_19053);
and U20985 (N_20985,N_19742,N_19225);
and U20986 (N_20986,N_19499,N_19983);
xnor U20987 (N_20987,N_19357,N_19948);
or U20988 (N_20988,N_19724,N_19722);
nand U20989 (N_20989,N_19636,N_19709);
nand U20990 (N_20990,N_19347,N_19802);
xnor U20991 (N_20991,N_19351,N_19543);
or U20992 (N_20992,N_19578,N_19240);
nand U20993 (N_20993,N_19244,N_19834);
or U20994 (N_20994,N_19343,N_19166);
nor U20995 (N_20995,N_19273,N_19523);
or U20996 (N_20996,N_19909,N_19935);
or U20997 (N_20997,N_19250,N_19622);
or U20998 (N_20998,N_19428,N_19476);
xor U20999 (N_20999,N_19274,N_19099);
nand U21000 (N_21000,N_20036,N_20968);
or U21001 (N_21001,N_20848,N_20502);
nand U21002 (N_21002,N_20196,N_20141);
or U21003 (N_21003,N_20399,N_20137);
xor U21004 (N_21004,N_20165,N_20274);
nor U21005 (N_21005,N_20197,N_20259);
or U21006 (N_21006,N_20297,N_20143);
nor U21007 (N_21007,N_20433,N_20486);
and U21008 (N_21008,N_20641,N_20246);
xor U21009 (N_21009,N_20917,N_20015);
xnor U21010 (N_21010,N_20513,N_20214);
nor U21011 (N_21011,N_20842,N_20612);
xor U21012 (N_21012,N_20822,N_20591);
xor U21013 (N_21013,N_20555,N_20028);
xor U21014 (N_21014,N_20097,N_20409);
nand U21015 (N_21015,N_20900,N_20172);
or U21016 (N_21016,N_20262,N_20990);
and U21017 (N_21017,N_20147,N_20057);
or U21018 (N_21018,N_20098,N_20017);
and U21019 (N_21019,N_20955,N_20412);
xor U21020 (N_21020,N_20898,N_20133);
and U21021 (N_21021,N_20031,N_20293);
nor U21022 (N_21022,N_20897,N_20609);
and U21023 (N_21023,N_20339,N_20943);
xnor U21024 (N_21024,N_20876,N_20084);
xor U21025 (N_21025,N_20786,N_20923);
nand U21026 (N_21026,N_20813,N_20243);
nor U21027 (N_21027,N_20765,N_20635);
xnor U21028 (N_21028,N_20276,N_20422);
nand U21029 (N_21029,N_20066,N_20270);
or U21030 (N_21030,N_20739,N_20527);
and U21031 (N_21031,N_20628,N_20020);
xnor U21032 (N_21032,N_20070,N_20731);
and U21033 (N_21033,N_20021,N_20489);
nor U21034 (N_21034,N_20154,N_20504);
nand U21035 (N_21035,N_20414,N_20785);
nand U21036 (N_21036,N_20878,N_20524);
or U21037 (N_21037,N_20784,N_20920);
or U21038 (N_21038,N_20152,N_20815);
nand U21039 (N_21039,N_20494,N_20799);
or U21040 (N_21040,N_20948,N_20092);
xor U21041 (N_21041,N_20940,N_20523);
nor U21042 (N_21042,N_20417,N_20039);
nor U21043 (N_21043,N_20597,N_20983);
and U21044 (N_21044,N_20620,N_20073);
and U21045 (N_21045,N_20460,N_20462);
nand U21046 (N_21046,N_20931,N_20171);
or U21047 (N_21047,N_20024,N_20327);
xnor U21048 (N_21048,N_20134,N_20730);
xnor U21049 (N_21049,N_20729,N_20715);
xnor U21050 (N_21050,N_20738,N_20312);
and U21051 (N_21051,N_20338,N_20218);
xor U21052 (N_21052,N_20025,N_20836);
nand U21053 (N_21053,N_20491,N_20603);
or U21054 (N_21054,N_20888,N_20874);
or U21055 (N_21055,N_20488,N_20007);
and U21056 (N_21056,N_20574,N_20265);
and U21057 (N_21057,N_20384,N_20185);
nand U21058 (N_21058,N_20778,N_20182);
and U21059 (N_21059,N_20446,N_20862);
and U21060 (N_21060,N_20249,N_20717);
nor U21061 (N_21061,N_20631,N_20072);
xor U21062 (N_21062,N_20088,N_20803);
nor U21063 (N_21063,N_20860,N_20238);
or U21064 (N_21064,N_20775,N_20354);
or U21065 (N_21065,N_20104,N_20754);
nand U21066 (N_21066,N_20053,N_20205);
xor U21067 (N_21067,N_20429,N_20038);
or U21068 (N_21068,N_20300,N_20012);
xnor U21069 (N_21069,N_20546,N_20379);
nand U21070 (N_21070,N_20101,N_20664);
xor U21071 (N_21071,N_20938,N_20065);
nand U21072 (N_21072,N_20936,N_20544);
and U21073 (N_21073,N_20183,N_20180);
nor U21074 (N_21074,N_20734,N_20564);
and U21075 (N_21075,N_20304,N_20884);
and U21076 (N_21076,N_20869,N_20213);
or U21077 (N_21077,N_20699,N_20311);
nand U21078 (N_21078,N_20618,N_20081);
and U21079 (N_21079,N_20964,N_20117);
nand U21080 (N_21080,N_20385,N_20161);
and U21081 (N_21081,N_20688,N_20740);
nand U21082 (N_21082,N_20541,N_20672);
nand U21083 (N_21083,N_20903,N_20946);
nand U21084 (N_21084,N_20347,N_20288);
and U21085 (N_21085,N_20201,N_20014);
xnor U21086 (N_21086,N_20334,N_20498);
xor U21087 (N_21087,N_20830,N_20211);
and U21088 (N_21088,N_20518,N_20472);
nand U21089 (N_21089,N_20596,N_20475);
xnor U21090 (N_21090,N_20168,N_20932);
xor U21091 (N_21091,N_20144,N_20291);
and U21092 (N_21092,N_20616,N_20637);
xnor U21093 (N_21093,N_20941,N_20724);
nor U21094 (N_21094,N_20352,N_20742);
and U21095 (N_21095,N_20549,N_20642);
and U21096 (N_21096,N_20411,N_20459);
or U21097 (N_21097,N_20284,N_20970);
xnor U21098 (N_21098,N_20625,N_20646);
and U21099 (N_21099,N_20834,N_20400);
xor U21100 (N_21100,N_20711,N_20187);
xor U21101 (N_21101,N_20426,N_20126);
or U21102 (N_21102,N_20059,N_20050);
or U21103 (N_21103,N_20610,N_20617);
nor U21104 (N_21104,N_20112,N_20669);
xor U21105 (N_21105,N_20146,N_20330);
xor U21106 (N_21106,N_20272,N_20814);
nand U21107 (N_21107,N_20841,N_20985);
and U21108 (N_21108,N_20561,N_20107);
and U21109 (N_21109,N_20175,N_20962);
and U21110 (N_21110,N_20481,N_20006);
and U21111 (N_21111,N_20566,N_20080);
or U21112 (N_21112,N_20883,N_20391);
nor U21113 (N_21113,N_20812,N_20468);
and U21114 (N_21114,N_20294,N_20174);
xor U21115 (N_21115,N_20124,N_20782);
and U21116 (N_21116,N_20693,N_20000);
nand U21117 (N_21117,N_20844,N_20105);
nor U21118 (N_21118,N_20747,N_20956);
nor U21119 (N_21119,N_20856,N_20506);
or U21120 (N_21120,N_20068,N_20278);
nand U21121 (N_21121,N_20167,N_20766);
or U21122 (N_21122,N_20027,N_20316);
or U21123 (N_21123,N_20054,N_20444);
xor U21124 (N_21124,N_20593,N_20443);
or U21125 (N_21125,N_20753,N_20662);
nand U21126 (N_21126,N_20223,N_20333);
and U21127 (N_21127,N_20470,N_20816);
or U21128 (N_21128,N_20567,N_20415);
nor U21129 (N_21129,N_20684,N_20335);
and U21130 (N_21130,N_20599,N_20727);
nand U21131 (N_21131,N_20780,N_20957);
and U21132 (N_21132,N_20085,N_20111);
nor U21133 (N_21133,N_20380,N_20351);
nand U21134 (N_21134,N_20592,N_20255);
or U21135 (N_21135,N_20198,N_20933);
xor U21136 (N_21136,N_20536,N_20037);
nand U21137 (N_21137,N_20353,N_20975);
nand U21138 (N_21138,N_20003,N_20594);
nor U21139 (N_21139,N_20302,N_20530);
xor U21140 (N_21140,N_20403,N_20295);
xor U21141 (N_21141,N_20543,N_20418);
or U21142 (N_21142,N_20222,N_20774);
and U21143 (N_21143,N_20621,N_20716);
nand U21144 (N_21144,N_20115,N_20756);
xor U21145 (N_21145,N_20389,N_20652);
or U21146 (N_21146,N_20170,N_20763);
nor U21147 (N_21147,N_20689,N_20306);
xor U21148 (N_21148,N_20551,N_20078);
or U21149 (N_21149,N_20916,N_20921);
or U21150 (N_21150,N_20273,N_20156);
nand U21151 (N_21151,N_20926,N_20209);
and U21152 (N_21152,N_20582,N_20746);
nand U21153 (N_21153,N_20407,N_20367);
nor U21154 (N_21154,N_20863,N_20533);
nand U21155 (N_21155,N_20480,N_20509);
nor U21156 (N_21156,N_20553,N_20539);
nor U21157 (N_21157,N_20336,N_20852);
or U21158 (N_21158,N_20918,N_20733);
xnor U21159 (N_21159,N_20030,N_20363);
or U21160 (N_21160,N_20944,N_20953);
xor U21161 (N_21161,N_20675,N_20911);
and U21162 (N_21162,N_20366,N_20627);
nor U21163 (N_21163,N_20548,N_20645);
nor U21164 (N_21164,N_20705,N_20034);
and U21165 (N_21165,N_20531,N_20887);
nor U21166 (N_21166,N_20889,N_20991);
xnor U21167 (N_21167,N_20685,N_20683);
xor U21168 (N_21168,N_20934,N_20718);
nor U21169 (N_21169,N_20648,N_20679);
or U21170 (N_21170,N_20189,N_20503);
nor U21171 (N_21171,N_20476,N_20035);
and U21172 (N_21172,N_20356,N_20710);
nor U21173 (N_21173,N_20419,N_20239);
nor U21174 (N_21174,N_20307,N_20033);
and U21175 (N_21175,N_20914,N_20691);
nor U21176 (N_21176,N_20195,N_20508);
and U21177 (N_21177,N_20629,N_20492);
or U21178 (N_21178,N_20535,N_20952);
xnor U21179 (N_21179,N_20893,N_20708);
nand U21180 (N_21180,N_20163,N_20723);
nand U21181 (N_21181,N_20505,N_20136);
and U21182 (N_21182,N_20455,N_20589);
or U21183 (N_21183,N_20919,N_20169);
or U21184 (N_21184,N_20817,N_20925);
nand U21185 (N_21185,N_20374,N_20581);
xor U21186 (N_21186,N_20980,N_20299);
xnor U21187 (N_21187,N_20252,N_20714);
nand U21188 (N_21188,N_20695,N_20974);
nand U21189 (N_21189,N_20483,N_20935);
nor U21190 (N_21190,N_20788,N_20118);
nor U21191 (N_21191,N_20741,N_20216);
and U21192 (N_21192,N_20212,N_20381);
nor U21193 (N_21193,N_20737,N_20789);
or U21194 (N_21194,N_20478,N_20682);
and U21195 (N_21195,N_20881,N_20280);
xor U21196 (N_21196,N_20692,N_20364);
nor U21197 (N_21197,N_20110,N_20927);
xor U21198 (N_21198,N_20305,N_20560);
nand U21199 (N_21199,N_20668,N_20382);
xor U21200 (N_21200,N_20989,N_20891);
nor U21201 (N_21201,N_20202,N_20702);
or U21202 (N_21202,N_20752,N_20082);
and U21203 (N_21203,N_20721,N_20512);
nor U21204 (N_21204,N_20430,N_20296);
or U21205 (N_21205,N_20556,N_20559);
nor U21206 (N_21206,N_20401,N_20833);
nor U21207 (N_21207,N_20630,N_20859);
or U21208 (N_21208,N_20829,N_20767);
or U21209 (N_21209,N_20632,N_20557);
nand U21210 (N_21210,N_20639,N_20359);
or U21211 (N_21211,N_20448,N_20537);
nand U21212 (N_21212,N_20160,N_20231);
and U21213 (N_21213,N_20271,N_20150);
nor U21214 (N_21214,N_20976,N_20602);
xor U21215 (N_21215,N_20485,N_20371);
or U21216 (N_21216,N_20571,N_20377);
and U21217 (N_21217,N_20845,N_20849);
and U21218 (N_21218,N_20395,N_20796);
or U21219 (N_21219,N_20640,N_20200);
or U21220 (N_21220,N_20586,N_20580);
xor U21221 (N_21221,N_20453,N_20858);
xnor U21222 (N_21222,N_20011,N_20886);
or U21223 (N_21223,N_20166,N_20406);
xor U21224 (N_21224,N_20568,N_20540);
xnor U21225 (N_21225,N_20096,N_20447);
xor U21226 (N_21226,N_20744,N_20676);
nor U21227 (N_21227,N_20009,N_20431);
nand U21228 (N_21228,N_20994,N_20001);
nand U21229 (N_21229,N_20607,N_20947);
xor U21230 (N_21230,N_20386,N_20469);
nor U21231 (N_21231,N_20519,N_20130);
nand U21232 (N_21232,N_20230,N_20058);
nand U21233 (N_21233,N_20119,N_20832);
xnor U21234 (N_21234,N_20987,N_20142);
nor U21235 (N_21235,N_20315,N_20824);
and U21236 (N_21236,N_20658,N_20062);
and U21237 (N_21237,N_20343,N_20713);
xor U21238 (N_21238,N_20825,N_20821);
nor U21239 (N_21239,N_20242,N_20611);
and U21240 (N_21240,N_20457,N_20759);
nor U21241 (N_21241,N_20572,N_20465);
nor U21242 (N_21242,N_20387,N_20704);
xnor U21243 (N_21243,N_20529,N_20452);
nor U21244 (N_21244,N_20971,N_20383);
xnor U21245 (N_21245,N_20314,N_20114);
or U21246 (N_21246,N_20499,N_20838);
nand U21247 (N_21247,N_20719,N_20982);
xnor U21248 (N_21248,N_20690,N_20321);
xnor U21249 (N_21249,N_20584,N_20232);
and U21250 (N_21250,N_20922,N_20538);
xor U21251 (N_21251,N_20224,N_20360);
nand U21252 (N_21252,N_20048,N_20550);
and U21253 (N_21253,N_20240,N_20608);
and U21254 (N_21254,N_20521,N_20855);
or U21255 (N_21255,N_20945,N_20042);
nand U21256 (N_21256,N_20969,N_20258);
nor U21257 (N_21257,N_20570,N_20928);
and U21258 (N_21258,N_20471,N_20768);
xor U21259 (N_21259,N_20257,N_20965);
nor U21260 (N_21260,N_20177,N_20372);
or U21261 (N_21261,N_20349,N_20215);
xor U21262 (N_21262,N_20002,N_20850);
and U21263 (N_21263,N_20425,N_20787);
nor U21264 (N_21264,N_20826,N_20275);
nor U21265 (N_21265,N_20287,N_20781);
or U21266 (N_21266,N_20325,N_20576);
nor U21267 (N_21267,N_20861,N_20261);
and U21268 (N_21268,N_20507,N_20398);
and U21269 (N_21269,N_20251,N_20913);
or U21270 (N_21270,N_20558,N_20600);
xnor U21271 (N_21271,N_20751,N_20879);
nand U21272 (N_21272,N_20516,N_20866);
xnor U21273 (N_21273,N_20487,N_20819);
and U21274 (N_21274,N_20896,N_20905);
or U21275 (N_21275,N_20776,N_20199);
nand U21276 (N_21276,N_20966,N_20253);
or U21277 (N_21277,N_20977,N_20100);
xnor U21278 (N_21278,N_20678,N_20902);
nor U21279 (N_21279,N_20466,N_20633);
nand U21280 (N_21280,N_20432,N_20158);
or U21281 (N_21281,N_20667,N_20378);
nor U21282 (N_21282,N_20707,N_20442);
nor U21283 (N_21283,N_20127,N_20697);
and U21284 (N_21284,N_20086,N_20565);
and U21285 (N_21285,N_20904,N_20102);
xnor U21286 (N_21286,N_20004,N_20424);
and U21287 (N_21287,N_20461,N_20496);
and U21288 (N_21288,N_20484,N_20959);
or U21289 (N_21289,N_20263,N_20585);
xor U21290 (N_21290,N_20563,N_20319);
nand U21291 (N_21291,N_20661,N_20873);
or U21292 (N_21292,N_20915,N_20256);
nor U21293 (N_21293,N_20772,N_20846);
and U21294 (N_21294,N_20277,N_20140);
xor U21295 (N_21295,N_20317,N_20208);
or U21296 (N_21296,N_20342,N_20290);
nor U21297 (N_21297,N_20234,N_20203);
nand U21298 (N_21298,N_20798,N_20190);
xnor U21299 (N_21299,N_20909,N_20770);
nor U21300 (N_21300,N_20043,N_20217);
or U21301 (N_21301,N_20666,N_20064);
xor U21302 (N_21302,N_20748,N_20026);
nand U21303 (N_21303,N_20388,N_20912);
and U21304 (N_21304,N_20283,N_20008);
xnor U21305 (N_21305,N_20247,N_20906);
nand U21306 (N_21306,N_20885,N_20963);
and U21307 (N_21307,N_20298,N_20619);
nor U21308 (N_21308,N_20226,N_20547);
or U21309 (N_21309,N_20245,N_20532);
or U21310 (N_21310,N_20427,N_20369);
xor U21311 (N_21311,N_20791,N_20286);
nand U21312 (N_21312,N_20857,N_20355);
or U21313 (N_21313,N_20099,N_20606);
xnor U21314 (N_21314,N_20810,N_20601);
xor U21315 (N_21315,N_20542,N_20434);
nor U21316 (N_21316,N_20949,N_20060);
or U21317 (N_21317,N_20501,N_20981);
nor U21318 (N_21318,N_20820,N_20954);
nor U21319 (N_21319,N_20750,N_20960);
and U21320 (N_21320,N_20663,N_20194);
and U21321 (N_21321,N_20522,N_20178);
nor U21322 (N_21322,N_20103,N_20157);
or U21323 (N_21323,N_20520,N_20041);
nand U21324 (N_21324,N_20871,N_20698);
xor U21325 (N_21325,N_20010,N_20394);
and U21326 (N_21326,N_20318,N_20076);
nand U21327 (N_21327,N_20901,N_20650);
or U21328 (N_21328,N_20292,N_20063);
xor U21329 (N_21329,N_20598,N_20326);
or U21330 (N_21330,N_20595,N_20743);
and U21331 (N_21331,N_20895,N_20908);
xor U21332 (N_21332,N_20375,N_20647);
or U21333 (N_21333,N_20077,N_20095);
nand U21334 (N_21334,N_20764,N_20517);
and U21335 (N_21335,N_20404,N_20924);
nor U21336 (N_21336,N_20075,N_20303);
xnor U21337 (N_21337,N_20069,N_20390);
or U21338 (N_21338,N_20206,N_20473);
nor U21339 (N_21339,N_20324,N_20942);
or U21340 (N_21340,N_20309,N_20313);
xnor U21341 (N_21341,N_20227,N_20090);
or U21342 (N_21342,N_20345,N_20526);
nor U21343 (N_21343,N_20769,N_20653);
and U21344 (N_21344,N_20464,N_20583);
or U21345 (N_21345,N_20792,N_20638);
nor U21346 (N_21346,N_20587,N_20843);
xnor U21347 (N_21347,N_20951,N_20220);
nor U21348 (N_21348,N_20332,N_20757);
or U21349 (N_21349,N_20973,N_20622);
xor U21350 (N_21350,N_20801,N_20545);
and U21351 (N_21351,N_20986,N_20049);
nand U21352 (N_21352,N_20978,N_20145);
nor U21353 (N_21353,N_20282,N_20651);
nor U21354 (N_21354,N_20660,N_20510);
nor U21355 (N_21355,N_20839,N_20569);
nand U21356 (N_21356,N_20013,N_20123);
nor U21357 (N_21357,N_20827,N_20458);
nand U21358 (N_21358,N_20939,N_20435);
or U21359 (N_21359,N_20368,N_20758);
and U21360 (N_21360,N_20807,N_20410);
nor U21361 (N_21361,N_20396,N_20525);
nor U21362 (N_21362,N_20162,N_20323);
or U21363 (N_21363,N_20773,N_20674);
and U21364 (N_21364,N_20248,N_20877);
and U21365 (N_21365,N_20700,N_20837);
or U21366 (N_21366,N_20310,N_20191);
or U21367 (N_21367,N_20121,N_20806);
xor U21368 (N_21368,N_20018,N_20413);
and U21369 (N_21369,N_20735,N_20937);
nor U21370 (N_21370,N_20999,N_20657);
and U21371 (N_21371,N_20184,N_20929);
nor U21372 (N_21372,N_20655,N_20087);
nor U21373 (N_21373,N_20495,N_20445);
xor U21374 (N_21374,N_20864,N_20930);
nand U21375 (N_21375,N_20726,N_20677);
xor U21376 (N_21376,N_20882,N_20696);
nand U21377 (N_21377,N_20490,N_20229);
nand U21378 (N_21378,N_20135,N_20865);
nand U21379 (N_21379,N_20493,N_20228);
nand U21380 (N_21380,N_20654,N_20588);
nand U21381 (N_21381,N_20055,N_20818);
xor U21382 (N_21382,N_20755,N_20659);
nand U21383 (N_21383,N_20720,N_20762);
and U21384 (N_21384,N_20260,N_20793);
and U21385 (N_21385,N_20370,N_20420);
nand U21386 (N_21386,N_20267,N_20188);
nor U21387 (N_21387,N_20680,N_20344);
or U21388 (N_21388,N_20346,N_20109);
nand U21389 (N_21389,N_20173,N_20337);
nor U21390 (N_21390,N_20301,N_20040);
nand U21391 (N_21391,N_20210,N_20463);
xor U21392 (N_21392,N_20736,N_20996);
nor U21393 (N_21393,N_20106,N_20131);
xnor U21394 (N_21394,N_20416,N_20074);
or U21395 (N_21395,N_20428,N_20071);
or U21396 (N_21396,N_20761,N_20079);
nor U21397 (N_21397,N_20835,N_20760);
nand U21398 (N_21398,N_20264,N_20155);
xnor U21399 (N_21399,N_20623,N_20797);
nor U21400 (N_21400,N_20061,N_20089);
nor U21401 (N_21401,N_20393,N_20179);
nor U21402 (N_21402,N_20643,N_20113);
or U21403 (N_21403,N_20235,N_20083);
xnor U21404 (N_21404,N_20056,N_20808);
or U21405 (N_21405,N_20441,N_20809);
xor U21406 (N_21406,N_20497,N_20578);
xnor U21407 (N_21407,N_20779,N_20467);
nand U21408 (N_21408,N_20790,N_20029);
xnor U21409 (N_21409,N_20528,N_20802);
nor U21410 (N_21410,N_20149,N_20614);
and U21411 (N_21411,N_20439,N_20500);
and U21412 (N_21412,N_20362,N_20725);
nor U21413 (N_21413,N_20482,N_20450);
nand U21414 (N_21414,N_20328,N_20984);
nand U21415 (N_21415,N_20613,N_20233);
xor U21416 (N_21416,N_20853,N_20219);
or U21417 (N_21417,N_20093,N_20051);
and U21418 (N_21418,N_20128,N_20783);
nor U21419 (N_21419,N_20350,N_20281);
xnor U21420 (N_21420,N_20044,N_20046);
nand U21421 (N_21421,N_20122,N_20132);
nor U21422 (N_21422,N_20722,N_20047);
xnor U21423 (N_21423,N_20045,N_20870);
or U21424 (N_21424,N_20795,N_20108);
nor U21425 (N_21425,N_20022,N_20285);
xnor U21426 (N_21426,N_20438,N_20266);
nor U21427 (N_21427,N_20005,N_20204);
nand U21428 (N_21428,N_20604,N_20289);
xnor U21429 (N_21429,N_20579,N_20225);
or U21430 (N_21430,N_20732,N_20749);
nor U21431 (N_21431,N_20615,N_20254);
nand U21432 (N_21432,N_20479,N_20811);
or U21433 (N_21433,N_20237,N_20148);
nand U21434 (N_21434,N_20880,N_20153);
or U21435 (N_21435,N_20348,N_20624);
nand U21436 (N_21436,N_20340,N_20554);
nor U21437 (N_21437,N_20192,N_20997);
and U21438 (N_21438,N_20397,N_20995);
or U21439 (N_21439,N_20176,N_20241);
or U21440 (N_21440,N_20405,N_20244);
and U21441 (N_21441,N_20577,N_20474);
and U21442 (N_21442,N_20186,N_20320);
xor U21443 (N_21443,N_20910,N_20032);
and U21444 (N_21444,N_20421,N_20534);
and U21445 (N_21445,N_20575,N_20402);
xor U21446 (N_21446,N_20828,N_20671);
xnor U21447 (N_21447,N_20673,N_20894);
and U21448 (N_21448,N_20139,N_20120);
nand U21449 (N_21449,N_20193,N_20890);
and U21450 (N_21450,N_20331,N_20023);
and U21451 (N_21451,N_20605,N_20573);
and U21452 (N_21452,N_20590,N_20998);
xnor U21453 (N_21453,N_20847,N_20052);
nand U21454 (N_21454,N_20125,N_20644);
nor U21455 (N_21455,N_20341,N_20562);
and U21456 (N_21456,N_20514,N_20670);
nor U21457 (N_21457,N_20703,N_20656);
and U21458 (N_21458,N_20322,N_20992);
xor U21459 (N_21459,N_20357,N_20159);
xor U21460 (N_21460,N_20972,N_20840);
nor U21461 (N_21461,N_20777,N_20687);
nand U21462 (N_21462,N_20511,N_20709);
xor U21463 (N_21463,N_20423,N_20408);
and U21464 (N_21464,N_20449,N_20268);
or U21465 (N_21465,N_20854,N_20164);
xnor U21466 (N_21466,N_20950,N_20181);
xor U21467 (N_21467,N_20805,N_20993);
or U21468 (N_21468,N_20823,N_20067);
and U21469 (N_21469,N_20712,N_20831);
nand U21470 (N_21470,N_20988,N_20376);
nor U21471 (N_21471,N_20236,N_20094);
nand U21472 (N_21472,N_20686,N_20701);
xor U21473 (N_21473,N_20358,N_20800);
or U21474 (N_21474,N_20269,N_20892);
xnor U21475 (N_21475,N_20091,N_20019);
or U21476 (N_21476,N_20308,N_20329);
nand U21477 (N_21477,N_20899,N_20867);
and U21478 (N_21478,N_20907,N_20016);
xor U21479 (N_21479,N_20361,N_20151);
nor U21480 (N_21480,N_20967,N_20552);
nand U21481 (N_21481,N_20868,N_20745);
or U21482 (N_21482,N_20851,N_20116);
xor U21483 (N_21483,N_20279,N_20771);
and U21484 (N_21484,N_20694,N_20436);
or U21485 (N_21485,N_20451,N_20681);
xor U21486 (N_21486,N_20392,N_20440);
xor U21487 (N_21487,N_20207,N_20477);
nand U21488 (N_21488,N_20875,N_20250);
nor U21489 (N_21489,N_20129,N_20515);
and U21490 (N_21490,N_20649,N_20636);
and U21491 (N_21491,N_20979,N_20634);
xnor U21492 (N_21492,N_20872,N_20221);
xor U21493 (N_21493,N_20961,N_20626);
and U21494 (N_21494,N_20373,N_20456);
nor U21495 (N_21495,N_20437,N_20804);
nand U21496 (N_21496,N_20138,N_20794);
or U21497 (N_21497,N_20665,N_20958);
xnor U21498 (N_21498,N_20365,N_20454);
xnor U21499 (N_21499,N_20706,N_20728);
xor U21500 (N_21500,N_20895,N_20139);
nand U21501 (N_21501,N_20366,N_20522);
nand U21502 (N_21502,N_20394,N_20196);
nor U21503 (N_21503,N_20316,N_20067);
or U21504 (N_21504,N_20748,N_20638);
xor U21505 (N_21505,N_20128,N_20589);
nor U21506 (N_21506,N_20573,N_20990);
nand U21507 (N_21507,N_20077,N_20187);
nand U21508 (N_21508,N_20908,N_20410);
nand U21509 (N_21509,N_20158,N_20973);
and U21510 (N_21510,N_20888,N_20223);
xor U21511 (N_21511,N_20523,N_20007);
xor U21512 (N_21512,N_20394,N_20121);
xor U21513 (N_21513,N_20845,N_20212);
or U21514 (N_21514,N_20518,N_20231);
nand U21515 (N_21515,N_20833,N_20903);
and U21516 (N_21516,N_20869,N_20723);
or U21517 (N_21517,N_20629,N_20898);
xor U21518 (N_21518,N_20959,N_20828);
and U21519 (N_21519,N_20515,N_20759);
or U21520 (N_21520,N_20654,N_20949);
xnor U21521 (N_21521,N_20300,N_20200);
and U21522 (N_21522,N_20401,N_20810);
and U21523 (N_21523,N_20656,N_20411);
or U21524 (N_21524,N_20636,N_20278);
and U21525 (N_21525,N_20357,N_20023);
xnor U21526 (N_21526,N_20169,N_20980);
or U21527 (N_21527,N_20698,N_20717);
nand U21528 (N_21528,N_20322,N_20970);
nand U21529 (N_21529,N_20433,N_20025);
nand U21530 (N_21530,N_20031,N_20760);
nand U21531 (N_21531,N_20901,N_20930);
nor U21532 (N_21532,N_20792,N_20465);
or U21533 (N_21533,N_20998,N_20288);
nand U21534 (N_21534,N_20816,N_20102);
nand U21535 (N_21535,N_20165,N_20401);
xnor U21536 (N_21536,N_20784,N_20987);
nand U21537 (N_21537,N_20968,N_20431);
xor U21538 (N_21538,N_20817,N_20281);
nand U21539 (N_21539,N_20874,N_20875);
nand U21540 (N_21540,N_20769,N_20339);
or U21541 (N_21541,N_20994,N_20402);
nor U21542 (N_21542,N_20685,N_20152);
xor U21543 (N_21543,N_20558,N_20172);
nand U21544 (N_21544,N_20850,N_20393);
xor U21545 (N_21545,N_20130,N_20393);
or U21546 (N_21546,N_20283,N_20496);
or U21547 (N_21547,N_20422,N_20087);
nor U21548 (N_21548,N_20476,N_20795);
nand U21549 (N_21549,N_20351,N_20363);
xor U21550 (N_21550,N_20562,N_20285);
and U21551 (N_21551,N_20547,N_20669);
and U21552 (N_21552,N_20024,N_20442);
xor U21553 (N_21553,N_20350,N_20505);
or U21554 (N_21554,N_20855,N_20176);
and U21555 (N_21555,N_20148,N_20833);
or U21556 (N_21556,N_20269,N_20899);
and U21557 (N_21557,N_20382,N_20789);
nor U21558 (N_21558,N_20682,N_20588);
and U21559 (N_21559,N_20041,N_20479);
nand U21560 (N_21560,N_20597,N_20406);
nor U21561 (N_21561,N_20036,N_20158);
xor U21562 (N_21562,N_20426,N_20560);
or U21563 (N_21563,N_20456,N_20223);
and U21564 (N_21564,N_20712,N_20457);
nor U21565 (N_21565,N_20038,N_20161);
xnor U21566 (N_21566,N_20177,N_20029);
nor U21567 (N_21567,N_20748,N_20484);
nor U21568 (N_21568,N_20771,N_20650);
and U21569 (N_21569,N_20483,N_20407);
nand U21570 (N_21570,N_20351,N_20279);
or U21571 (N_21571,N_20909,N_20176);
or U21572 (N_21572,N_20920,N_20425);
nand U21573 (N_21573,N_20372,N_20149);
and U21574 (N_21574,N_20041,N_20204);
and U21575 (N_21575,N_20614,N_20479);
nor U21576 (N_21576,N_20399,N_20568);
and U21577 (N_21577,N_20318,N_20003);
nor U21578 (N_21578,N_20868,N_20074);
nand U21579 (N_21579,N_20448,N_20735);
and U21580 (N_21580,N_20939,N_20078);
or U21581 (N_21581,N_20438,N_20236);
nor U21582 (N_21582,N_20011,N_20985);
xor U21583 (N_21583,N_20722,N_20433);
and U21584 (N_21584,N_20129,N_20680);
nand U21585 (N_21585,N_20004,N_20571);
nor U21586 (N_21586,N_20896,N_20109);
and U21587 (N_21587,N_20699,N_20168);
nand U21588 (N_21588,N_20951,N_20558);
or U21589 (N_21589,N_20199,N_20971);
nor U21590 (N_21590,N_20526,N_20176);
xnor U21591 (N_21591,N_20996,N_20127);
nor U21592 (N_21592,N_20801,N_20307);
and U21593 (N_21593,N_20974,N_20746);
xnor U21594 (N_21594,N_20022,N_20766);
and U21595 (N_21595,N_20688,N_20786);
or U21596 (N_21596,N_20133,N_20094);
nor U21597 (N_21597,N_20955,N_20388);
nor U21598 (N_21598,N_20786,N_20145);
xor U21599 (N_21599,N_20381,N_20830);
nand U21600 (N_21600,N_20514,N_20846);
or U21601 (N_21601,N_20861,N_20398);
xor U21602 (N_21602,N_20616,N_20087);
or U21603 (N_21603,N_20998,N_20514);
xor U21604 (N_21604,N_20354,N_20649);
nor U21605 (N_21605,N_20032,N_20583);
or U21606 (N_21606,N_20725,N_20486);
nand U21607 (N_21607,N_20315,N_20697);
or U21608 (N_21608,N_20939,N_20070);
nor U21609 (N_21609,N_20688,N_20677);
and U21610 (N_21610,N_20074,N_20400);
xor U21611 (N_21611,N_20976,N_20177);
nand U21612 (N_21612,N_20785,N_20195);
xnor U21613 (N_21613,N_20981,N_20594);
and U21614 (N_21614,N_20301,N_20015);
or U21615 (N_21615,N_20224,N_20310);
nand U21616 (N_21616,N_20194,N_20583);
or U21617 (N_21617,N_20467,N_20237);
or U21618 (N_21618,N_20562,N_20773);
nand U21619 (N_21619,N_20299,N_20178);
nor U21620 (N_21620,N_20070,N_20325);
nand U21621 (N_21621,N_20781,N_20279);
xor U21622 (N_21622,N_20354,N_20469);
or U21623 (N_21623,N_20240,N_20189);
xnor U21624 (N_21624,N_20717,N_20764);
or U21625 (N_21625,N_20759,N_20656);
xnor U21626 (N_21626,N_20221,N_20206);
and U21627 (N_21627,N_20830,N_20905);
and U21628 (N_21628,N_20726,N_20800);
or U21629 (N_21629,N_20083,N_20566);
or U21630 (N_21630,N_20635,N_20026);
nand U21631 (N_21631,N_20510,N_20135);
nand U21632 (N_21632,N_20925,N_20326);
or U21633 (N_21633,N_20072,N_20487);
and U21634 (N_21634,N_20009,N_20779);
xnor U21635 (N_21635,N_20016,N_20038);
xnor U21636 (N_21636,N_20952,N_20264);
xor U21637 (N_21637,N_20448,N_20818);
nand U21638 (N_21638,N_20673,N_20921);
nor U21639 (N_21639,N_20577,N_20250);
xnor U21640 (N_21640,N_20413,N_20456);
nand U21641 (N_21641,N_20174,N_20746);
xnor U21642 (N_21642,N_20897,N_20520);
and U21643 (N_21643,N_20151,N_20051);
and U21644 (N_21644,N_20244,N_20868);
and U21645 (N_21645,N_20203,N_20131);
or U21646 (N_21646,N_20948,N_20147);
nor U21647 (N_21647,N_20575,N_20370);
and U21648 (N_21648,N_20726,N_20308);
or U21649 (N_21649,N_20227,N_20936);
nor U21650 (N_21650,N_20660,N_20545);
nand U21651 (N_21651,N_20865,N_20530);
nand U21652 (N_21652,N_20382,N_20295);
or U21653 (N_21653,N_20421,N_20982);
xnor U21654 (N_21654,N_20139,N_20223);
xor U21655 (N_21655,N_20242,N_20638);
nand U21656 (N_21656,N_20764,N_20899);
and U21657 (N_21657,N_20523,N_20366);
or U21658 (N_21658,N_20081,N_20817);
and U21659 (N_21659,N_20231,N_20146);
and U21660 (N_21660,N_20054,N_20811);
or U21661 (N_21661,N_20391,N_20469);
or U21662 (N_21662,N_20262,N_20716);
and U21663 (N_21663,N_20117,N_20698);
and U21664 (N_21664,N_20523,N_20888);
or U21665 (N_21665,N_20727,N_20129);
nor U21666 (N_21666,N_20921,N_20999);
xor U21667 (N_21667,N_20000,N_20575);
nor U21668 (N_21668,N_20513,N_20652);
nor U21669 (N_21669,N_20162,N_20534);
nor U21670 (N_21670,N_20636,N_20339);
nand U21671 (N_21671,N_20261,N_20901);
nand U21672 (N_21672,N_20435,N_20060);
xnor U21673 (N_21673,N_20933,N_20764);
xnor U21674 (N_21674,N_20982,N_20015);
or U21675 (N_21675,N_20919,N_20944);
or U21676 (N_21676,N_20493,N_20678);
xnor U21677 (N_21677,N_20693,N_20631);
or U21678 (N_21678,N_20053,N_20294);
xor U21679 (N_21679,N_20211,N_20523);
or U21680 (N_21680,N_20977,N_20539);
xor U21681 (N_21681,N_20783,N_20801);
and U21682 (N_21682,N_20905,N_20179);
nand U21683 (N_21683,N_20087,N_20726);
nor U21684 (N_21684,N_20771,N_20950);
or U21685 (N_21685,N_20552,N_20503);
and U21686 (N_21686,N_20510,N_20234);
and U21687 (N_21687,N_20292,N_20744);
or U21688 (N_21688,N_20287,N_20539);
xnor U21689 (N_21689,N_20219,N_20629);
xnor U21690 (N_21690,N_20167,N_20004);
or U21691 (N_21691,N_20678,N_20275);
or U21692 (N_21692,N_20108,N_20859);
and U21693 (N_21693,N_20215,N_20574);
nor U21694 (N_21694,N_20487,N_20942);
or U21695 (N_21695,N_20469,N_20578);
nor U21696 (N_21696,N_20332,N_20705);
xor U21697 (N_21697,N_20387,N_20439);
nand U21698 (N_21698,N_20599,N_20832);
or U21699 (N_21699,N_20848,N_20675);
xor U21700 (N_21700,N_20728,N_20509);
nand U21701 (N_21701,N_20480,N_20318);
nand U21702 (N_21702,N_20988,N_20372);
xnor U21703 (N_21703,N_20404,N_20224);
xnor U21704 (N_21704,N_20496,N_20929);
nand U21705 (N_21705,N_20933,N_20356);
nor U21706 (N_21706,N_20844,N_20367);
and U21707 (N_21707,N_20332,N_20477);
and U21708 (N_21708,N_20491,N_20808);
nand U21709 (N_21709,N_20538,N_20357);
and U21710 (N_21710,N_20455,N_20820);
and U21711 (N_21711,N_20842,N_20013);
or U21712 (N_21712,N_20060,N_20798);
nand U21713 (N_21713,N_20272,N_20740);
or U21714 (N_21714,N_20697,N_20586);
nor U21715 (N_21715,N_20091,N_20242);
and U21716 (N_21716,N_20985,N_20311);
nand U21717 (N_21717,N_20592,N_20179);
nand U21718 (N_21718,N_20190,N_20314);
nand U21719 (N_21719,N_20356,N_20689);
xnor U21720 (N_21720,N_20661,N_20325);
nand U21721 (N_21721,N_20213,N_20850);
nand U21722 (N_21722,N_20759,N_20903);
and U21723 (N_21723,N_20883,N_20979);
xor U21724 (N_21724,N_20533,N_20626);
or U21725 (N_21725,N_20321,N_20043);
xnor U21726 (N_21726,N_20359,N_20754);
nand U21727 (N_21727,N_20975,N_20994);
xnor U21728 (N_21728,N_20052,N_20935);
xor U21729 (N_21729,N_20649,N_20722);
xor U21730 (N_21730,N_20109,N_20741);
or U21731 (N_21731,N_20554,N_20465);
nor U21732 (N_21732,N_20437,N_20825);
xnor U21733 (N_21733,N_20448,N_20831);
nor U21734 (N_21734,N_20593,N_20027);
xor U21735 (N_21735,N_20221,N_20257);
or U21736 (N_21736,N_20827,N_20978);
nor U21737 (N_21737,N_20903,N_20353);
xnor U21738 (N_21738,N_20512,N_20358);
or U21739 (N_21739,N_20521,N_20975);
and U21740 (N_21740,N_20281,N_20566);
or U21741 (N_21741,N_20975,N_20392);
or U21742 (N_21742,N_20273,N_20383);
xnor U21743 (N_21743,N_20995,N_20648);
or U21744 (N_21744,N_20066,N_20382);
nor U21745 (N_21745,N_20204,N_20349);
nand U21746 (N_21746,N_20268,N_20109);
nand U21747 (N_21747,N_20625,N_20000);
nand U21748 (N_21748,N_20132,N_20139);
and U21749 (N_21749,N_20692,N_20216);
xnor U21750 (N_21750,N_20109,N_20778);
or U21751 (N_21751,N_20459,N_20865);
and U21752 (N_21752,N_20318,N_20711);
nor U21753 (N_21753,N_20557,N_20434);
nor U21754 (N_21754,N_20559,N_20704);
nor U21755 (N_21755,N_20562,N_20044);
xor U21756 (N_21756,N_20025,N_20911);
nor U21757 (N_21757,N_20701,N_20639);
and U21758 (N_21758,N_20121,N_20447);
or U21759 (N_21759,N_20451,N_20558);
xor U21760 (N_21760,N_20707,N_20893);
or U21761 (N_21761,N_20028,N_20775);
nand U21762 (N_21762,N_20622,N_20220);
or U21763 (N_21763,N_20751,N_20990);
nand U21764 (N_21764,N_20569,N_20950);
nand U21765 (N_21765,N_20210,N_20879);
nor U21766 (N_21766,N_20068,N_20513);
or U21767 (N_21767,N_20902,N_20812);
and U21768 (N_21768,N_20028,N_20615);
and U21769 (N_21769,N_20514,N_20199);
or U21770 (N_21770,N_20030,N_20888);
nand U21771 (N_21771,N_20959,N_20685);
and U21772 (N_21772,N_20273,N_20748);
nor U21773 (N_21773,N_20612,N_20247);
or U21774 (N_21774,N_20344,N_20369);
nand U21775 (N_21775,N_20830,N_20328);
and U21776 (N_21776,N_20638,N_20889);
xor U21777 (N_21777,N_20645,N_20978);
xor U21778 (N_21778,N_20819,N_20812);
nand U21779 (N_21779,N_20617,N_20277);
and U21780 (N_21780,N_20795,N_20314);
and U21781 (N_21781,N_20103,N_20018);
nand U21782 (N_21782,N_20559,N_20206);
xnor U21783 (N_21783,N_20375,N_20868);
nor U21784 (N_21784,N_20758,N_20831);
or U21785 (N_21785,N_20174,N_20718);
nand U21786 (N_21786,N_20308,N_20866);
xor U21787 (N_21787,N_20784,N_20527);
xnor U21788 (N_21788,N_20921,N_20701);
nand U21789 (N_21789,N_20293,N_20445);
nor U21790 (N_21790,N_20374,N_20776);
or U21791 (N_21791,N_20826,N_20091);
and U21792 (N_21792,N_20004,N_20350);
nor U21793 (N_21793,N_20654,N_20885);
nor U21794 (N_21794,N_20813,N_20425);
xor U21795 (N_21795,N_20384,N_20355);
and U21796 (N_21796,N_20767,N_20780);
or U21797 (N_21797,N_20209,N_20976);
xnor U21798 (N_21798,N_20163,N_20677);
nand U21799 (N_21799,N_20343,N_20476);
nand U21800 (N_21800,N_20794,N_20230);
and U21801 (N_21801,N_20948,N_20716);
xor U21802 (N_21802,N_20878,N_20412);
nand U21803 (N_21803,N_20454,N_20407);
xor U21804 (N_21804,N_20186,N_20081);
nand U21805 (N_21805,N_20401,N_20902);
nor U21806 (N_21806,N_20037,N_20238);
nor U21807 (N_21807,N_20045,N_20349);
xor U21808 (N_21808,N_20367,N_20324);
nor U21809 (N_21809,N_20492,N_20075);
or U21810 (N_21810,N_20695,N_20749);
nor U21811 (N_21811,N_20909,N_20520);
or U21812 (N_21812,N_20197,N_20948);
xnor U21813 (N_21813,N_20228,N_20384);
nand U21814 (N_21814,N_20955,N_20790);
or U21815 (N_21815,N_20031,N_20892);
xor U21816 (N_21816,N_20539,N_20422);
nand U21817 (N_21817,N_20415,N_20228);
or U21818 (N_21818,N_20952,N_20690);
xor U21819 (N_21819,N_20113,N_20508);
xor U21820 (N_21820,N_20052,N_20702);
and U21821 (N_21821,N_20090,N_20707);
nor U21822 (N_21822,N_20921,N_20317);
nand U21823 (N_21823,N_20620,N_20350);
and U21824 (N_21824,N_20573,N_20229);
nor U21825 (N_21825,N_20391,N_20884);
or U21826 (N_21826,N_20596,N_20038);
and U21827 (N_21827,N_20949,N_20981);
xor U21828 (N_21828,N_20226,N_20283);
or U21829 (N_21829,N_20459,N_20985);
or U21830 (N_21830,N_20003,N_20214);
nor U21831 (N_21831,N_20690,N_20367);
nand U21832 (N_21832,N_20404,N_20478);
nor U21833 (N_21833,N_20713,N_20308);
or U21834 (N_21834,N_20591,N_20922);
xnor U21835 (N_21835,N_20300,N_20325);
xnor U21836 (N_21836,N_20311,N_20903);
nor U21837 (N_21837,N_20408,N_20098);
or U21838 (N_21838,N_20602,N_20651);
xor U21839 (N_21839,N_20671,N_20628);
or U21840 (N_21840,N_20835,N_20602);
nor U21841 (N_21841,N_20159,N_20806);
nand U21842 (N_21842,N_20366,N_20986);
nand U21843 (N_21843,N_20904,N_20812);
or U21844 (N_21844,N_20562,N_20296);
or U21845 (N_21845,N_20954,N_20262);
or U21846 (N_21846,N_20412,N_20923);
xor U21847 (N_21847,N_20923,N_20972);
nor U21848 (N_21848,N_20752,N_20411);
or U21849 (N_21849,N_20783,N_20075);
and U21850 (N_21850,N_20723,N_20680);
nor U21851 (N_21851,N_20674,N_20324);
nand U21852 (N_21852,N_20689,N_20425);
xnor U21853 (N_21853,N_20585,N_20656);
xnor U21854 (N_21854,N_20016,N_20589);
and U21855 (N_21855,N_20227,N_20763);
nand U21856 (N_21856,N_20873,N_20274);
and U21857 (N_21857,N_20575,N_20091);
or U21858 (N_21858,N_20649,N_20745);
nor U21859 (N_21859,N_20090,N_20506);
nor U21860 (N_21860,N_20368,N_20619);
nand U21861 (N_21861,N_20784,N_20519);
nand U21862 (N_21862,N_20856,N_20603);
and U21863 (N_21863,N_20258,N_20293);
nand U21864 (N_21864,N_20799,N_20511);
xnor U21865 (N_21865,N_20511,N_20470);
nand U21866 (N_21866,N_20038,N_20776);
or U21867 (N_21867,N_20564,N_20964);
or U21868 (N_21868,N_20085,N_20195);
nand U21869 (N_21869,N_20634,N_20450);
nor U21870 (N_21870,N_20168,N_20436);
xor U21871 (N_21871,N_20915,N_20293);
or U21872 (N_21872,N_20572,N_20070);
or U21873 (N_21873,N_20620,N_20843);
nor U21874 (N_21874,N_20786,N_20886);
nor U21875 (N_21875,N_20625,N_20806);
nor U21876 (N_21876,N_20636,N_20053);
nand U21877 (N_21877,N_20161,N_20349);
nand U21878 (N_21878,N_20621,N_20527);
nand U21879 (N_21879,N_20956,N_20263);
nand U21880 (N_21880,N_20239,N_20316);
xnor U21881 (N_21881,N_20464,N_20007);
and U21882 (N_21882,N_20947,N_20877);
or U21883 (N_21883,N_20983,N_20326);
and U21884 (N_21884,N_20567,N_20804);
nand U21885 (N_21885,N_20463,N_20274);
or U21886 (N_21886,N_20865,N_20870);
or U21887 (N_21887,N_20773,N_20469);
xnor U21888 (N_21888,N_20005,N_20052);
or U21889 (N_21889,N_20429,N_20565);
nand U21890 (N_21890,N_20232,N_20347);
nand U21891 (N_21891,N_20784,N_20566);
nor U21892 (N_21892,N_20925,N_20378);
or U21893 (N_21893,N_20225,N_20272);
nand U21894 (N_21894,N_20404,N_20491);
nor U21895 (N_21895,N_20461,N_20381);
nand U21896 (N_21896,N_20816,N_20746);
nor U21897 (N_21897,N_20550,N_20218);
nor U21898 (N_21898,N_20704,N_20057);
or U21899 (N_21899,N_20332,N_20664);
nand U21900 (N_21900,N_20450,N_20144);
or U21901 (N_21901,N_20080,N_20614);
and U21902 (N_21902,N_20605,N_20497);
nor U21903 (N_21903,N_20479,N_20594);
nand U21904 (N_21904,N_20607,N_20972);
and U21905 (N_21905,N_20948,N_20715);
nor U21906 (N_21906,N_20586,N_20996);
nor U21907 (N_21907,N_20205,N_20871);
nand U21908 (N_21908,N_20327,N_20622);
or U21909 (N_21909,N_20662,N_20882);
or U21910 (N_21910,N_20346,N_20648);
xnor U21911 (N_21911,N_20460,N_20996);
and U21912 (N_21912,N_20879,N_20733);
nand U21913 (N_21913,N_20408,N_20835);
xnor U21914 (N_21914,N_20648,N_20563);
or U21915 (N_21915,N_20212,N_20549);
nand U21916 (N_21916,N_20585,N_20607);
and U21917 (N_21917,N_20157,N_20248);
or U21918 (N_21918,N_20595,N_20264);
xor U21919 (N_21919,N_20436,N_20214);
nand U21920 (N_21920,N_20930,N_20376);
or U21921 (N_21921,N_20483,N_20091);
nand U21922 (N_21922,N_20630,N_20931);
nor U21923 (N_21923,N_20860,N_20883);
nor U21924 (N_21924,N_20771,N_20978);
and U21925 (N_21925,N_20797,N_20120);
or U21926 (N_21926,N_20174,N_20722);
nand U21927 (N_21927,N_20855,N_20252);
nor U21928 (N_21928,N_20042,N_20644);
nor U21929 (N_21929,N_20568,N_20311);
nor U21930 (N_21930,N_20630,N_20071);
xor U21931 (N_21931,N_20860,N_20794);
nand U21932 (N_21932,N_20655,N_20992);
and U21933 (N_21933,N_20148,N_20034);
and U21934 (N_21934,N_20793,N_20980);
or U21935 (N_21935,N_20421,N_20723);
xnor U21936 (N_21936,N_20291,N_20288);
nand U21937 (N_21937,N_20433,N_20412);
or U21938 (N_21938,N_20045,N_20115);
and U21939 (N_21939,N_20255,N_20494);
and U21940 (N_21940,N_20654,N_20236);
nor U21941 (N_21941,N_20362,N_20789);
nor U21942 (N_21942,N_20079,N_20686);
nor U21943 (N_21943,N_20260,N_20263);
and U21944 (N_21944,N_20216,N_20269);
nor U21945 (N_21945,N_20957,N_20383);
xnor U21946 (N_21946,N_20634,N_20639);
or U21947 (N_21947,N_20967,N_20271);
or U21948 (N_21948,N_20866,N_20806);
nand U21949 (N_21949,N_20434,N_20752);
or U21950 (N_21950,N_20284,N_20146);
nand U21951 (N_21951,N_20735,N_20474);
xnor U21952 (N_21952,N_20637,N_20785);
nor U21953 (N_21953,N_20266,N_20381);
xnor U21954 (N_21954,N_20247,N_20729);
xnor U21955 (N_21955,N_20789,N_20741);
xnor U21956 (N_21956,N_20736,N_20285);
and U21957 (N_21957,N_20581,N_20840);
nor U21958 (N_21958,N_20837,N_20422);
xor U21959 (N_21959,N_20602,N_20805);
and U21960 (N_21960,N_20114,N_20575);
and U21961 (N_21961,N_20272,N_20149);
nand U21962 (N_21962,N_20595,N_20814);
or U21963 (N_21963,N_20880,N_20174);
and U21964 (N_21964,N_20238,N_20280);
and U21965 (N_21965,N_20804,N_20140);
xnor U21966 (N_21966,N_20864,N_20163);
and U21967 (N_21967,N_20094,N_20017);
nor U21968 (N_21968,N_20939,N_20940);
or U21969 (N_21969,N_20179,N_20378);
and U21970 (N_21970,N_20880,N_20453);
nand U21971 (N_21971,N_20021,N_20127);
or U21972 (N_21972,N_20276,N_20947);
nor U21973 (N_21973,N_20431,N_20486);
nor U21974 (N_21974,N_20754,N_20778);
or U21975 (N_21975,N_20670,N_20949);
xor U21976 (N_21976,N_20185,N_20651);
xnor U21977 (N_21977,N_20507,N_20448);
nand U21978 (N_21978,N_20853,N_20124);
nand U21979 (N_21979,N_20405,N_20241);
nand U21980 (N_21980,N_20448,N_20707);
nor U21981 (N_21981,N_20023,N_20502);
or U21982 (N_21982,N_20062,N_20392);
and U21983 (N_21983,N_20607,N_20822);
or U21984 (N_21984,N_20341,N_20941);
nand U21985 (N_21985,N_20916,N_20751);
or U21986 (N_21986,N_20641,N_20423);
or U21987 (N_21987,N_20189,N_20302);
nand U21988 (N_21988,N_20719,N_20327);
xnor U21989 (N_21989,N_20630,N_20755);
or U21990 (N_21990,N_20287,N_20048);
xnor U21991 (N_21991,N_20342,N_20809);
xor U21992 (N_21992,N_20956,N_20707);
and U21993 (N_21993,N_20536,N_20495);
and U21994 (N_21994,N_20165,N_20570);
nor U21995 (N_21995,N_20838,N_20482);
or U21996 (N_21996,N_20447,N_20535);
nand U21997 (N_21997,N_20317,N_20363);
nor U21998 (N_21998,N_20746,N_20117);
nor U21999 (N_21999,N_20695,N_20162);
or U22000 (N_22000,N_21684,N_21339);
nor U22001 (N_22001,N_21292,N_21063);
xnor U22002 (N_22002,N_21344,N_21807);
nor U22003 (N_22003,N_21636,N_21989);
nand U22004 (N_22004,N_21088,N_21779);
and U22005 (N_22005,N_21407,N_21284);
or U22006 (N_22006,N_21534,N_21094);
xnor U22007 (N_22007,N_21512,N_21409);
and U22008 (N_22008,N_21624,N_21111);
nor U22009 (N_22009,N_21789,N_21499);
and U22010 (N_22010,N_21559,N_21629);
nand U22011 (N_22011,N_21658,N_21209);
or U22012 (N_22012,N_21225,N_21932);
or U22013 (N_22013,N_21328,N_21297);
and U22014 (N_22014,N_21736,N_21296);
nand U22015 (N_22015,N_21238,N_21047);
or U22016 (N_22016,N_21659,N_21640);
nand U22017 (N_22017,N_21199,N_21536);
nor U22018 (N_22018,N_21928,N_21473);
nand U22019 (N_22019,N_21436,N_21605);
nor U22020 (N_22020,N_21431,N_21160);
and U22021 (N_22021,N_21946,N_21362);
or U22022 (N_22022,N_21885,N_21260);
nor U22023 (N_22023,N_21745,N_21654);
nand U22024 (N_22024,N_21738,N_21428);
or U22025 (N_22025,N_21938,N_21445);
nand U22026 (N_22026,N_21870,N_21994);
nor U22027 (N_22027,N_21136,N_21583);
nand U22028 (N_22028,N_21894,N_21934);
nor U22029 (N_22029,N_21718,N_21776);
or U22030 (N_22030,N_21053,N_21993);
xnor U22031 (N_22031,N_21236,N_21579);
and U22032 (N_22032,N_21118,N_21501);
or U22033 (N_22033,N_21137,N_21502);
or U22034 (N_22034,N_21358,N_21283);
xor U22035 (N_22035,N_21714,N_21844);
xor U22036 (N_22036,N_21641,N_21150);
or U22037 (N_22037,N_21850,N_21661);
xnor U22038 (N_22038,N_21530,N_21325);
and U22039 (N_22039,N_21140,N_21333);
nand U22040 (N_22040,N_21315,N_21656);
xor U22041 (N_22041,N_21628,N_21016);
and U22042 (N_22042,N_21911,N_21737);
and U22043 (N_22043,N_21625,N_21207);
and U22044 (N_22044,N_21538,N_21183);
nand U22045 (N_22045,N_21816,N_21293);
xor U22046 (N_22046,N_21769,N_21637);
nor U22047 (N_22047,N_21185,N_21206);
nor U22048 (N_22048,N_21398,N_21275);
or U22049 (N_22049,N_21319,N_21954);
xnor U22050 (N_22050,N_21890,N_21569);
xor U22051 (N_22051,N_21271,N_21177);
or U22052 (N_22052,N_21146,N_21895);
and U22053 (N_22053,N_21696,N_21755);
xnor U22054 (N_22054,N_21316,N_21467);
xor U22055 (N_22055,N_21197,N_21313);
and U22056 (N_22056,N_21359,N_21215);
nor U22057 (N_22057,N_21517,N_21848);
or U22058 (N_22058,N_21253,N_21231);
nand U22059 (N_22059,N_21670,N_21560);
nand U22060 (N_22060,N_21123,N_21263);
and U22061 (N_22061,N_21212,N_21607);
nand U22062 (N_22062,N_21385,N_21280);
and U22063 (N_22063,N_21775,N_21320);
or U22064 (N_22064,N_21087,N_21335);
or U22065 (N_22065,N_21672,N_21771);
xnor U22066 (N_22066,N_21376,N_21978);
xnor U22067 (N_22067,N_21960,N_21809);
and U22068 (N_22068,N_21105,N_21674);
or U22069 (N_22069,N_21759,N_21852);
xnor U22070 (N_22070,N_21104,N_21553);
or U22071 (N_22071,N_21195,N_21575);
xor U22072 (N_22072,N_21290,N_21015);
or U22073 (N_22073,N_21233,N_21814);
xnor U22074 (N_22074,N_21478,N_21375);
nor U22075 (N_22075,N_21457,N_21777);
nor U22076 (N_22076,N_21999,N_21794);
nor U22077 (N_22077,N_21336,N_21214);
xnor U22078 (N_22078,N_21144,N_21109);
xnor U22079 (N_22079,N_21049,N_21797);
nor U22080 (N_22080,N_21285,N_21429);
xor U22081 (N_22081,N_21472,N_21089);
or U22082 (N_22082,N_21190,N_21606);
and U22083 (N_22083,N_21617,N_21305);
nor U22084 (N_22084,N_21166,N_21947);
nor U22085 (N_22085,N_21391,N_21623);
nor U22086 (N_22086,N_21036,N_21544);
or U22087 (N_22087,N_21026,N_21237);
nand U22088 (N_22088,N_21121,N_21338);
and U22089 (N_22089,N_21519,N_21732);
and U22090 (N_22090,N_21592,N_21399);
and U22091 (N_22091,N_21829,N_21787);
nand U22092 (N_22092,N_21318,N_21649);
xor U22093 (N_22093,N_21835,N_21308);
xor U22094 (N_22094,N_21991,N_21688);
nor U22095 (N_22095,N_21493,N_21154);
xor U22096 (N_22096,N_21984,N_21168);
or U22097 (N_22097,N_21303,N_21784);
nand U22098 (N_22098,N_21124,N_21521);
xnor U22099 (N_22099,N_21572,N_21581);
xor U22100 (N_22100,N_21926,N_21093);
nand U22101 (N_22101,N_21471,N_21372);
nor U22102 (N_22102,N_21642,N_21173);
or U22103 (N_22103,N_21956,N_21044);
nand U22104 (N_22104,N_21007,N_21891);
and U22105 (N_22105,N_21716,N_21011);
nor U22106 (N_22106,N_21985,N_21614);
and U22107 (N_22107,N_21198,N_21252);
xnor U22108 (N_22108,N_21447,N_21347);
or U22109 (N_22109,N_21145,N_21180);
and U22110 (N_22110,N_21005,N_21753);
nor U22111 (N_22111,N_21261,N_21806);
nor U22112 (N_22112,N_21576,N_21241);
xor U22113 (N_22113,N_21821,N_21465);
or U22114 (N_22114,N_21090,N_21153);
and U22115 (N_22115,N_21662,N_21570);
nor U22116 (N_22116,N_21176,N_21772);
nor U22117 (N_22117,N_21849,N_21324);
nand U22118 (N_22118,N_21446,N_21799);
or U22119 (N_22119,N_21065,N_21029);
xnor U22120 (N_22120,N_21915,N_21227);
and U22121 (N_22121,N_21615,N_21485);
and U22122 (N_22122,N_21676,N_21919);
nor U22123 (N_22123,N_21550,N_21585);
nor U22124 (N_22124,N_21685,N_21076);
nand U22125 (N_22125,N_21669,N_21880);
nand U22126 (N_22126,N_21059,N_21980);
xor U22127 (N_22127,N_21998,N_21413);
xnor U22128 (N_22128,N_21546,N_21596);
or U22129 (N_22129,N_21773,N_21851);
nand U22130 (N_22130,N_21506,N_21223);
nor U22131 (N_22131,N_21108,N_21700);
nor U22132 (N_22132,N_21668,N_21069);
nor U22133 (N_22133,N_21634,N_21652);
and U22134 (N_22134,N_21189,N_21792);
xnor U22135 (N_22135,N_21057,N_21403);
or U22136 (N_22136,N_21229,N_21356);
xnor U22137 (N_22137,N_21143,N_21631);
xor U22138 (N_22138,N_21205,N_21497);
nand U22139 (N_22139,N_21783,N_21027);
xor U22140 (N_22140,N_21416,N_21766);
xnor U22141 (N_22141,N_21510,N_21874);
and U22142 (N_22142,N_21620,N_21922);
nand U22143 (N_22143,N_21235,N_21132);
nand U22144 (N_22144,N_21962,N_21255);
nand U22145 (N_22145,N_21170,N_21957);
nand U22146 (N_22146,N_21925,N_21474);
xor U22147 (N_22147,N_21883,N_21547);
nand U22148 (N_22148,N_21393,N_21839);
nor U22149 (N_22149,N_21125,N_21704);
nor U22150 (N_22150,N_21479,N_21912);
nand U22151 (N_22151,N_21520,N_21077);
nor U22152 (N_22152,N_21566,N_21348);
nand U22153 (N_22153,N_21720,N_21217);
or U22154 (N_22154,N_21580,N_21887);
and U22155 (N_22155,N_21020,N_21360);
nand U22156 (N_22156,N_21451,N_21908);
or U22157 (N_22157,N_21749,N_21882);
and U22158 (N_22158,N_21635,N_21188);
nand U22159 (N_22159,N_21258,N_21099);
nor U22160 (N_22160,N_21349,N_21167);
nor U22161 (N_22161,N_21781,N_21708);
nand U22162 (N_22162,N_21054,N_21495);
and U22163 (N_22163,N_21010,N_21172);
xor U22164 (N_22164,N_21441,N_21815);
xor U22165 (N_22165,N_21147,N_21646);
nand U22166 (N_22166,N_21001,N_21793);
and U22167 (N_22167,N_21687,N_21317);
and U22168 (N_22168,N_21128,N_21936);
nand U22169 (N_22169,N_21548,N_21698);
or U22170 (N_22170,N_21159,N_21556);
nand U22171 (N_22171,N_21706,N_21003);
xnor U22172 (N_22172,N_21950,N_21847);
nand U22173 (N_22173,N_21910,N_21463);
and U22174 (N_22174,N_21804,N_21216);
and U22175 (N_22175,N_21500,N_21552);
nand U22176 (N_22176,N_21655,N_21056);
nand U22177 (N_22177,N_21110,N_21892);
nor U22178 (N_22178,N_21958,N_21224);
nor U22179 (N_22179,N_21918,N_21062);
nor U22180 (N_22180,N_21332,N_21876);
or U22181 (N_22181,N_21509,N_21304);
and U22182 (N_22182,N_21148,N_21249);
and U22183 (N_22183,N_21419,N_21481);
nand U22184 (N_22184,N_21751,N_21830);
nor U22185 (N_22185,N_21211,N_21130);
xor U22186 (N_22186,N_21435,N_21055);
nor U22187 (N_22187,N_21460,N_21394);
nor U22188 (N_22188,N_21450,N_21306);
nand U22189 (N_22189,N_21854,N_21459);
and U22190 (N_22190,N_21196,N_21012);
xor U22191 (N_22191,N_21555,N_21837);
xnor U22192 (N_22192,N_21272,N_21256);
xnor U22193 (N_22193,N_21037,N_21959);
or U22194 (N_22194,N_21721,N_21486);
nor U22195 (N_22195,N_21423,N_21082);
or U22196 (N_22196,N_21786,N_21941);
or U22197 (N_22197,N_21013,N_21232);
or U22198 (N_22198,N_21432,N_21475);
xnor U22199 (N_22199,N_21587,N_21192);
or U22200 (N_22200,N_21097,N_21187);
xnor U22201 (N_22201,N_21265,N_21469);
or U22202 (N_22202,N_21021,N_21905);
or U22203 (N_22203,N_21071,N_21856);
and U22204 (N_22204,N_21357,N_21643);
or U22205 (N_22205,N_21009,N_21599);
nand U22206 (N_22206,N_21503,N_21203);
nor U22207 (N_22207,N_21135,N_21677);
nand U22208 (N_22208,N_21571,N_21330);
or U22209 (N_22209,N_21299,N_21302);
or U22210 (N_22210,N_21683,N_21909);
nor U22211 (N_22211,N_21609,N_21392);
and U22212 (N_22212,N_21412,N_21279);
nand U22213 (N_22213,N_21343,N_21632);
or U22214 (N_22214,N_21161,N_21788);
or U22215 (N_22215,N_21162,N_21767);
xnor U22216 (N_22216,N_21014,N_21595);
nor U22217 (N_22217,N_21757,N_21386);
nor U22218 (N_22218,N_21041,N_21120);
nor U22219 (N_22219,N_21411,N_21884);
or U22220 (N_22220,N_21370,N_21401);
nand U22221 (N_22221,N_21484,N_21597);
xnor U22222 (N_22222,N_21095,N_21404);
nand U22223 (N_22223,N_21591,N_21080);
xor U22224 (N_22224,N_21052,N_21417);
xnor U22225 (N_22225,N_21100,N_21836);
nand U22226 (N_22226,N_21384,N_21897);
and U22227 (N_22227,N_21711,N_21184);
xnor U22228 (N_22228,N_21964,N_21365);
nor U22229 (N_22229,N_21245,N_21528);
nand U22230 (N_22230,N_21537,N_21803);
and U22231 (N_22231,N_21045,N_21762);
nand U22232 (N_22232,N_21701,N_21179);
nor U22233 (N_22233,N_21174,N_21778);
and U22234 (N_22234,N_21420,N_21115);
or U22235 (N_22235,N_21156,N_21462);
nor U22236 (N_22236,N_21675,N_21443);
nand U22237 (N_22237,N_21035,N_21933);
nand U22238 (N_22238,N_21453,N_21322);
nand U22239 (N_22239,N_21931,N_21254);
and U22240 (N_22240,N_21877,N_21327);
nor U22241 (N_22241,N_21748,N_21096);
or U22242 (N_22242,N_21639,N_21812);
nor U22243 (N_22243,N_21865,N_21171);
xor U22244 (N_22244,N_21752,N_21702);
and U22245 (N_22245,N_21942,N_21692);
and U22246 (N_22246,N_21564,N_21660);
xor U22247 (N_22247,N_21667,N_21981);
nor U22248 (N_22248,N_21782,N_21378);
nor U22249 (N_22249,N_21487,N_21855);
and U22250 (N_22250,N_21801,N_21201);
and U22251 (N_22251,N_21665,N_21971);
nor U22252 (N_22252,N_21951,N_21619);
and U22253 (N_22253,N_21006,N_21785);
or U22254 (N_22254,N_21899,N_21200);
nand U22255 (N_22255,N_21276,N_21651);
xor U22256 (N_22256,N_21274,N_21158);
and U22257 (N_22257,N_21731,N_21827);
nand U22258 (N_22258,N_21067,N_21246);
or U22259 (N_22259,N_21907,N_21425);
xnor U22260 (N_22260,N_21540,N_21562);
and U22261 (N_22261,N_21030,N_21050);
and U22262 (N_22262,N_21191,N_21524);
xor U22263 (N_22263,N_21741,N_21878);
and U22264 (N_22264,N_21278,N_21664);
nor U22265 (N_22265,N_21833,N_21813);
or U22266 (N_22266,N_21454,N_21647);
nand U22267 (N_22267,N_21390,N_21522);
and U22268 (N_22268,N_21103,N_21477);
and U22269 (N_22269,N_21987,N_21355);
nand U22270 (N_22270,N_21397,N_21970);
and U22271 (N_22271,N_21992,N_21131);
nand U22272 (N_22272,N_21307,N_21722);
nor U22273 (N_22273,N_21439,N_21542);
xnor U22274 (N_22274,N_21842,N_21935);
and U22275 (N_22275,N_21515,N_21712);
nor U22276 (N_22276,N_21221,N_21818);
and U22277 (N_22277,N_21997,N_21367);
nor U22278 (N_22278,N_21734,N_21653);
or U22279 (N_22279,N_21598,N_21588);
nand U22280 (N_22280,N_21374,N_21742);
xnor U22281 (N_22281,N_21577,N_21976);
xnor U22282 (N_22282,N_21511,N_21418);
xnor U22283 (N_22283,N_21289,N_21139);
or U22284 (N_22284,N_21526,N_21427);
nand U22285 (N_22285,N_21387,N_21220);
or U22286 (N_22286,N_21996,N_21081);
or U22287 (N_22287,N_21808,N_21600);
nand U22288 (N_22288,N_21025,N_21551);
xor U22289 (N_22289,N_21549,N_21323);
xnor U22290 (N_22290,N_21682,N_21995);
or U22291 (N_22291,N_21841,N_21068);
nand U22292 (N_22292,N_21155,N_21175);
xor U22293 (N_22293,N_21298,N_21230);
or U22294 (N_22294,N_21226,N_21079);
nand U22295 (N_22295,N_21165,N_21686);
and U22296 (N_22296,N_21151,N_21843);
or U22297 (N_22297,N_21483,N_21612);
xor U22298 (N_22298,N_21904,N_21066);
and U22299 (N_22299,N_21291,N_21824);
or U22300 (N_22300,N_21380,N_21898);
or U22301 (N_22301,N_21930,N_21273);
or U22302 (N_22302,N_21990,N_21955);
xor U22303 (N_22303,N_21248,N_21482);
xor U22304 (N_22304,N_21354,N_21948);
xnor U22305 (N_22305,N_21092,N_21680);
and U22306 (N_22306,N_21149,N_21456);
nor U22307 (N_22307,N_21314,N_21868);
nor U22308 (N_22308,N_21084,N_21590);
nand U22309 (N_22309,N_21532,N_21896);
nand U22310 (N_22310,N_21507,N_21917);
and U22311 (N_22311,N_21480,N_21589);
or U22312 (N_22312,N_21601,N_21886);
and U22313 (N_22313,N_21949,N_21138);
and U22314 (N_22314,N_21798,N_21494);
xor U22315 (N_22315,N_21790,N_21965);
nor U22316 (N_22316,N_21492,N_21690);
xor U22317 (N_22317,N_21114,N_21944);
nand U22318 (N_22318,N_21703,N_21630);
nand U22319 (N_22319,N_21421,N_21262);
or U22320 (N_22320,N_21287,N_21901);
and U22321 (N_22321,N_21468,N_21545);
nor U22322 (N_22322,N_21846,N_21710);
nand U22323 (N_22323,N_21913,N_21604);
or U22324 (N_22324,N_21234,N_21764);
or U22325 (N_22325,N_21414,N_21770);
nand U22326 (N_22326,N_21717,N_21040);
xnor U22327 (N_22327,N_21337,N_21920);
and U22328 (N_22328,N_21043,N_21210);
or U22329 (N_22329,N_21295,N_21361);
or U22330 (N_22330,N_21018,N_21881);
or U22331 (N_22331,N_21780,N_21527);
or U22332 (N_22332,N_21430,N_21747);
nand U22333 (N_22333,N_21986,N_21709);
and U22334 (N_22334,N_21645,N_21134);
and U22335 (N_22335,N_21610,N_21193);
nor U22336 (N_22336,N_21750,N_21893);
nand U22337 (N_22337,N_21679,N_21098);
nor U22338 (N_22338,N_21763,N_21405);
nand U22339 (N_22339,N_21754,N_21961);
and U22340 (N_22340,N_21730,N_21832);
and U22341 (N_22341,N_21496,N_21019);
nand U22342 (N_22342,N_21142,N_21657);
nand U22343 (N_22343,N_21004,N_21903);
nor U22344 (N_22344,N_21074,N_21705);
xor U22345 (N_22345,N_21437,N_21440);
xnor U22346 (N_22346,N_21022,N_21963);
and U22347 (N_22347,N_21578,N_21264);
xnor U22348 (N_22348,N_21085,N_21523);
and U22349 (N_22349,N_21396,N_21294);
nand U22350 (N_22350,N_21728,N_21715);
nor U22351 (N_22351,N_21678,N_21765);
nand U22352 (N_22352,N_21796,N_21239);
or U22353 (N_22353,N_21584,N_21694);
or U22354 (N_22354,N_21389,N_21426);
or U22355 (N_22355,N_21565,N_21377);
and U22356 (N_22356,N_21247,N_21558);
nor U22357 (N_22357,N_21689,N_21573);
xor U22358 (N_22358,N_21194,N_21823);
or U22359 (N_22359,N_21663,N_21000);
or U22360 (N_22360,N_21864,N_21321);
xnor U22361 (N_22361,N_21611,N_21567);
nor U22362 (N_22362,N_21438,N_21363);
xnor U22363 (N_22363,N_21017,N_21400);
xor U22364 (N_22364,N_21034,N_21086);
or U22365 (N_22365,N_21863,N_21574);
nor U22366 (N_22366,N_21444,N_21743);
or U22367 (N_22367,N_21383,N_21373);
xor U22368 (N_22368,N_21906,N_21972);
and U22369 (N_22369,N_21541,N_21860);
nand U22370 (N_22370,N_21967,N_21859);
and U22371 (N_22371,N_21916,N_21593);
nor U22372 (N_22372,N_21504,N_21433);
xnor U22373 (N_22373,N_21603,N_21760);
or U22374 (N_22374,N_21464,N_21023);
nor U22375 (N_22375,N_21008,N_21288);
or U22376 (N_22376,N_21382,N_21204);
nand U22377 (N_22377,N_21648,N_21352);
and U22378 (N_22378,N_21845,N_21379);
xor U22379 (N_22379,N_21873,N_21529);
xnor U22380 (N_22380,N_21982,N_21921);
xnor U22381 (N_22381,N_21697,N_21539);
nand U22382 (N_22382,N_21758,N_21724);
and U22383 (N_22383,N_21442,N_21070);
and U22384 (N_22384,N_21244,N_21133);
or U22385 (N_22385,N_21113,N_21723);
or U22386 (N_22386,N_21927,N_21518);
or U22387 (N_22387,N_21448,N_21825);
nor U22388 (N_22388,N_21046,N_21939);
nand U22389 (N_22389,N_21719,N_21761);
and U22390 (N_22390,N_21726,N_21351);
nand U22391 (N_22391,N_21106,N_21811);
nor U22392 (N_22392,N_21902,N_21740);
nand U22393 (N_22393,N_21002,N_21800);
or U22394 (N_22394,N_21735,N_21557);
and U22395 (N_22395,N_21681,N_21461);
nand U22396 (N_22396,N_21282,N_21458);
nand U22397 (N_22397,N_21650,N_21107);
or U22398 (N_22398,N_21119,N_21988);
and U22399 (N_22399,N_21673,N_21817);
and U22400 (N_22400,N_21281,N_21466);
and U22401 (N_22401,N_21300,N_21822);
and U22402 (N_22402,N_21819,N_21310);
xnor U22403 (N_22403,N_21756,N_21953);
nor U22404 (N_22404,N_21102,N_21112);
xor U22405 (N_22405,N_21943,N_21693);
and U22406 (N_22406,N_21060,N_21408);
xnor U22407 (N_22407,N_21270,N_21739);
nor U22408 (N_22408,N_21627,N_21117);
and U22409 (N_22409,N_21489,N_21434);
and U22410 (N_22410,N_21422,N_21979);
nor U22411 (N_22411,N_21410,N_21340);
or U22412 (N_22412,N_21038,N_21369);
xor U22413 (N_22413,N_21586,N_21031);
xor U22414 (N_22414,N_21810,N_21508);
nor U22415 (N_22415,N_21582,N_21805);
and U22416 (N_22416,N_21622,N_21350);
xnor U22417 (N_22417,N_21346,N_21309);
and U22418 (N_22418,N_21101,N_21608);
or U22419 (N_22419,N_21768,N_21415);
nand U22420 (N_22420,N_21455,N_21301);
xnor U22421 (N_22421,N_21072,N_21498);
and U22422 (N_22422,N_21061,N_21618);
or U22423 (N_22423,N_21857,N_21866);
and U22424 (N_22424,N_21032,N_21802);
and U22425 (N_22425,N_21152,N_21388);
and U22426 (N_22426,N_21516,N_21476);
nor U22427 (N_22427,N_21312,N_21078);
and U22428 (N_22428,N_21795,N_21831);
xor U22429 (N_22429,N_21406,N_21733);
and U22430 (N_22430,N_21621,N_21725);
xor U22431 (N_22431,N_21838,N_21381);
or U22432 (N_22432,N_21364,N_21286);
nor U22433 (N_22433,N_21186,N_21341);
nand U22434 (N_22434,N_21969,N_21353);
and U22435 (N_22435,N_21983,N_21858);
nor U22436 (N_22436,N_21525,N_21940);
or U22437 (N_22437,N_21277,N_21242);
and U22438 (N_22438,N_21028,N_21695);
nor U22439 (N_22439,N_21181,N_21975);
nor U22440 (N_22440,N_21218,N_21488);
nand U22441 (N_22441,N_21867,N_21977);
nor U22442 (N_22442,N_21853,N_21974);
and U22443 (N_22443,N_21116,N_21157);
xor U22444 (N_22444,N_21729,N_21083);
nor U22445 (N_22445,N_21543,N_21869);
nor U22446 (N_22446,N_21671,N_21644);
and U22447 (N_22447,N_21240,N_21937);
or U22448 (N_22448,N_21929,N_21505);
nand U22449 (N_22449,N_21535,N_21638);
xor U22450 (N_22450,N_21250,N_21042);
nand U22451 (N_22451,N_21871,N_21875);
and U22452 (N_22452,N_21329,N_21311);
nor U22453 (N_22453,N_21127,N_21924);
nor U22454 (N_22454,N_21952,N_21923);
xnor U22455 (N_22455,N_21602,N_21470);
nor U22456 (N_22456,N_21395,N_21533);
and U22457 (N_22457,N_21744,N_21208);
xor U22458 (N_22458,N_21269,N_21727);
and U22459 (N_22459,N_21945,N_21219);
nand U22460 (N_22460,N_21973,N_21213);
and U22461 (N_22461,N_21129,N_21914);
and U22462 (N_22462,N_21064,N_21122);
xor U22463 (N_22463,N_21126,N_21251);
nor U22464 (N_22464,N_21490,N_21164);
nor U22465 (N_22465,N_21024,N_21345);
and U22466 (N_22466,N_21368,N_21699);
xor U22467 (N_22467,N_21202,N_21563);
nor U22468 (N_22468,N_21326,N_21058);
nand U22469 (N_22469,N_21222,N_21691);
and U22470 (N_22470,N_21073,N_21834);
xor U22471 (N_22471,N_21568,N_21826);
and U22472 (N_22472,N_21091,N_21257);
nor U22473 (N_22473,N_21554,N_21514);
and U22474 (N_22474,N_21594,N_21424);
or U22475 (N_22475,N_21840,N_21228);
xnor U22476 (N_22476,N_21182,N_21774);
or U22477 (N_22477,N_21334,N_21561);
and U22478 (N_22478,N_21075,N_21666);
nand U22479 (N_22479,N_21889,N_21371);
and U22480 (N_22480,N_21169,N_21513);
xor U22481 (N_22481,N_21266,N_21968);
nor U22482 (N_22482,N_21900,N_21616);
nor U22483 (N_22483,N_21626,N_21243);
or U22484 (N_22484,N_21791,N_21707);
and U22485 (N_22485,N_21178,N_21342);
or U22486 (N_22486,N_21452,N_21888);
nor U22487 (N_22487,N_21613,N_21449);
nand U22488 (N_22488,N_21862,N_21331);
or U22489 (N_22489,N_21141,N_21966);
xnor U22490 (N_22490,N_21048,N_21268);
nand U22491 (N_22491,N_21828,N_21872);
nand U22492 (N_22492,N_21879,N_21861);
nor U22493 (N_22493,N_21713,N_21491);
nor U22494 (N_22494,N_21531,N_21366);
or U22495 (N_22495,N_21039,N_21051);
nand U22496 (N_22496,N_21259,N_21163);
and U22497 (N_22497,N_21746,N_21402);
or U22498 (N_22498,N_21267,N_21820);
and U22499 (N_22499,N_21633,N_21033);
or U22500 (N_22500,N_21337,N_21288);
or U22501 (N_22501,N_21587,N_21109);
nor U22502 (N_22502,N_21079,N_21164);
and U22503 (N_22503,N_21804,N_21970);
nand U22504 (N_22504,N_21662,N_21526);
or U22505 (N_22505,N_21667,N_21616);
or U22506 (N_22506,N_21088,N_21368);
and U22507 (N_22507,N_21207,N_21361);
nand U22508 (N_22508,N_21008,N_21885);
nand U22509 (N_22509,N_21508,N_21363);
nand U22510 (N_22510,N_21190,N_21174);
xor U22511 (N_22511,N_21316,N_21201);
xnor U22512 (N_22512,N_21621,N_21790);
nor U22513 (N_22513,N_21167,N_21335);
or U22514 (N_22514,N_21566,N_21284);
xor U22515 (N_22515,N_21052,N_21091);
and U22516 (N_22516,N_21469,N_21305);
xor U22517 (N_22517,N_21139,N_21281);
or U22518 (N_22518,N_21862,N_21020);
or U22519 (N_22519,N_21270,N_21121);
nor U22520 (N_22520,N_21421,N_21928);
nor U22521 (N_22521,N_21772,N_21166);
nor U22522 (N_22522,N_21756,N_21673);
nand U22523 (N_22523,N_21649,N_21612);
or U22524 (N_22524,N_21584,N_21391);
nand U22525 (N_22525,N_21129,N_21241);
nand U22526 (N_22526,N_21332,N_21217);
xor U22527 (N_22527,N_21251,N_21821);
or U22528 (N_22528,N_21759,N_21684);
nor U22529 (N_22529,N_21407,N_21317);
xor U22530 (N_22530,N_21647,N_21064);
xnor U22531 (N_22531,N_21792,N_21753);
or U22532 (N_22532,N_21386,N_21082);
or U22533 (N_22533,N_21473,N_21536);
nand U22534 (N_22534,N_21158,N_21478);
xnor U22535 (N_22535,N_21463,N_21172);
and U22536 (N_22536,N_21162,N_21865);
and U22537 (N_22537,N_21400,N_21959);
nand U22538 (N_22538,N_21306,N_21202);
nand U22539 (N_22539,N_21715,N_21123);
nand U22540 (N_22540,N_21465,N_21615);
or U22541 (N_22541,N_21049,N_21682);
and U22542 (N_22542,N_21580,N_21308);
and U22543 (N_22543,N_21372,N_21302);
and U22544 (N_22544,N_21207,N_21757);
nand U22545 (N_22545,N_21421,N_21548);
nand U22546 (N_22546,N_21816,N_21587);
nor U22547 (N_22547,N_21904,N_21418);
and U22548 (N_22548,N_21787,N_21228);
nor U22549 (N_22549,N_21979,N_21831);
or U22550 (N_22550,N_21307,N_21503);
nand U22551 (N_22551,N_21135,N_21434);
xor U22552 (N_22552,N_21951,N_21849);
and U22553 (N_22553,N_21021,N_21611);
or U22554 (N_22554,N_21058,N_21853);
nor U22555 (N_22555,N_21138,N_21631);
xor U22556 (N_22556,N_21359,N_21795);
and U22557 (N_22557,N_21374,N_21208);
and U22558 (N_22558,N_21821,N_21235);
nor U22559 (N_22559,N_21783,N_21572);
nand U22560 (N_22560,N_21467,N_21242);
nand U22561 (N_22561,N_21738,N_21524);
nand U22562 (N_22562,N_21283,N_21625);
nor U22563 (N_22563,N_21380,N_21823);
nand U22564 (N_22564,N_21008,N_21018);
nor U22565 (N_22565,N_21904,N_21023);
nand U22566 (N_22566,N_21657,N_21312);
and U22567 (N_22567,N_21786,N_21419);
nor U22568 (N_22568,N_21206,N_21690);
xnor U22569 (N_22569,N_21139,N_21699);
or U22570 (N_22570,N_21152,N_21804);
nand U22571 (N_22571,N_21790,N_21019);
nor U22572 (N_22572,N_21209,N_21076);
and U22573 (N_22573,N_21901,N_21130);
and U22574 (N_22574,N_21287,N_21165);
nand U22575 (N_22575,N_21314,N_21216);
and U22576 (N_22576,N_21589,N_21970);
xnor U22577 (N_22577,N_21108,N_21134);
or U22578 (N_22578,N_21271,N_21437);
and U22579 (N_22579,N_21436,N_21468);
xnor U22580 (N_22580,N_21699,N_21761);
and U22581 (N_22581,N_21788,N_21230);
nand U22582 (N_22582,N_21469,N_21890);
or U22583 (N_22583,N_21215,N_21009);
xor U22584 (N_22584,N_21046,N_21959);
xor U22585 (N_22585,N_21314,N_21929);
nand U22586 (N_22586,N_21058,N_21821);
xor U22587 (N_22587,N_21790,N_21509);
nand U22588 (N_22588,N_21883,N_21675);
xor U22589 (N_22589,N_21910,N_21140);
and U22590 (N_22590,N_21834,N_21134);
or U22591 (N_22591,N_21519,N_21403);
xnor U22592 (N_22592,N_21372,N_21227);
nand U22593 (N_22593,N_21712,N_21870);
nand U22594 (N_22594,N_21147,N_21184);
nand U22595 (N_22595,N_21439,N_21494);
nor U22596 (N_22596,N_21365,N_21962);
nand U22597 (N_22597,N_21078,N_21636);
xor U22598 (N_22598,N_21007,N_21316);
xor U22599 (N_22599,N_21359,N_21123);
and U22600 (N_22600,N_21831,N_21964);
nor U22601 (N_22601,N_21972,N_21619);
nand U22602 (N_22602,N_21630,N_21753);
nand U22603 (N_22603,N_21191,N_21567);
and U22604 (N_22604,N_21700,N_21253);
or U22605 (N_22605,N_21194,N_21156);
nor U22606 (N_22606,N_21871,N_21495);
xnor U22607 (N_22607,N_21343,N_21450);
nand U22608 (N_22608,N_21940,N_21315);
nor U22609 (N_22609,N_21725,N_21359);
xnor U22610 (N_22610,N_21051,N_21717);
nor U22611 (N_22611,N_21486,N_21039);
nand U22612 (N_22612,N_21158,N_21229);
and U22613 (N_22613,N_21557,N_21085);
xnor U22614 (N_22614,N_21187,N_21656);
nand U22615 (N_22615,N_21607,N_21207);
xor U22616 (N_22616,N_21770,N_21837);
and U22617 (N_22617,N_21653,N_21932);
or U22618 (N_22618,N_21839,N_21065);
nand U22619 (N_22619,N_21407,N_21040);
xor U22620 (N_22620,N_21961,N_21016);
or U22621 (N_22621,N_21828,N_21928);
and U22622 (N_22622,N_21122,N_21243);
nor U22623 (N_22623,N_21323,N_21377);
nand U22624 (N_22624,N_21772,N_21813);
nand U22625 (N_22625,N_21926,N_21200);
nand U22626 (N_22626,N_21839,N_21696);
nand U22627 (N_22627,N_21261,N_21705);
nand U22628 (N_22628,N_21531,N_21787);
xor U22629 (N_22629,N_21176,N_21634);
nand U22630 (N_22630,N_21633,N_21592);
and U22631 (N_22631,N_21575,N_21250);
xor U22632 (N_22632,N_21629,N_21493);
nand U22633 (N_22633,N_21294,N_21158);
xor U22634 (N_22634,N_21219,N_21193);
or U22635 (N_22635,N_21273,N_21076);
nor U22636 (N_22636,N_21654,N_21116);
or U22637 (N_22637,N_21478,N_21781);
or U22638 (N_22638,N_21240,N_21473);
nor U22639 (N_22639,N_21974,N_21562);
nand U22640 (N_22640,N_21278,N_21025);
or U22641 (N_22641,N_21768,N_21522);
nor U22642 (N_22642,N_21363,N_21091);
and U22643 (N_22643,N_21439,N_21577);
nor U22644 (N_22644,N_21509,N_21838);
xor U22645 (N_22645,N_21258,N_21926);
or U22646 (N_22646,N_21029,N_21318);
or U22647 (N_22647,N_21524,N_21872);
and U22648 (N_22648,N_21740,N_21369);
and U22649 (N_22649,N_21970,N_21368);
and U22650 (N_22650,N_21535,N_21421);
xor U22651 (N_22651,N_21498,N_21730);
nor U22652 (N_22652,N_21243,N_21154);
nand U22653 (N_22653,N_21012,N_21973);
xor U22654 (N_22654,N_21646,N_21322);
nor U22655 (N_22655,N_21268,N_21018);
and U22656 (N_22656,N_21628,N_21106);
nor U22657 (N_22657,N_21057,N_21068);
xor U22658 (N_22658,N_21755,N_21409);
and U22659 (N_22659,N_21888,N_21857);
and U22660 (N_22660,N_21443,N_21247);
nor U22661 (N_22661,N_21354,N_21761);
or U22662 (N_22662,N_21918,N_21747);
xnor U22663 (N_22663,N_21504,N_21472);
xor U22664 (N_22664,N_21579,N_21588);
or U22665 (N_22665,N_21717,N_21888);
xor U22666 (N_22666,N_21793,N_21091);
and U22667 (N_22667,N_21184,N_21329);
or U22668 (N_22668,N_21607,N_21149);
nand U22669 (N_22669,N_21085,N_21397);
and U22670 (N_22670,N_21902,N_21758);
nand U22671 (N_22671,N_21826,N_21381);
nor U22672 (N_22672,N_21459,N_21343);
nand U22673 (N_22673,N_21011,N_21707);
nand U22674 (N_22674,N_21835,N_21675);
xor U22675 (N_22675,N_21218,N_21940);
nor U22676 (N_22676,N_21081,N_21810);
or U22677 (N_22677,N_21180,N_21510);
or U22678 (N_22678,N_21638,N_21785);
xor U22679 (N_22679,N_21695,N_21762);
xor U22680 (N_22680,N_21472,N_21044);
nor U22681 (N_22681,N_21530,N_21631);
or U22682 (N_22682,N_21435,N_21268);
xor U22683 (N_22683,N_21970,N_21042);
nor U22684 (N_22684,N_21832,N_21641);
nand U22685 (N_22685,N_21358,N_21823);
xor U22686 (N_22686,N_21891,N_21509);
and U22687 (N_22687,N_21762,N_21714);
nand U22688 (N_22688,N_21507,N_21582);
nand U22689 (N_22689,N_21232,N_21494);
or U22690 (N_22690,N_21231,N_21611);
nand U22691 (N_22691,N_21498,N_21077);
or U22692 (N_22692,N_21892,N_21421);
and U22693 (N_22693,N_21751,N_21640);
xnor U22694 (N_22694,N_21616,N_21906);
nor U22695 (N_22695,N_21473,N_21026);
xor U22696 (N_22696,N_21638,N_21572);
xnor U22697 (N_22697,N_21669,N_21924);
xnor U22698 (N_22698,N_21621,N_21505);
nand U22699 (N_22699,N_21638,N_21683);
nand U22700 (N_22700,N_21657,N_21796);
xor U22701 (N_22701,N_21431,N_21402);
nor U22702 (N_22702,N_21154,N_21854);
nand U22703 (N_22703,N_21896,N_21623);
nor U22704 (N_22704,N_21001,N_21155);
xor U22705 (N_22705,N_21418,N_21114);
xor U22706 (N_22706,N_21344,N_21862);
nand U22707 (N_22707,N_21899,N_21897);
nor U22708 (N_22708,N_21149,N_21682);
nand U22709 (N_22709,N_21772,N_21899);
xnor U22710 (N_22710,N_21332,N_21412);
xnor U22711 (N_22711,N_21759,N_21732);
and U22712 (N_22712,N_21605,N_21572);
and U22713 (N_22713,N_21528,N_21369);
nor U22714 (N_22714,N_21661,N_21674);
or U22715 (N_22715,N_21338,N_21997);
nand U22716 (N_22716,N_21423,N_21547);
and U22717 (N_22717,N_21400,N_21853);
and U22718 (N_22718,N_21737,N_21219);
and U22719 (N_22719,N_21564,N_21504);
or U22720 (N_22720,N_21347,N_21619);
nor U22721 (N_22721,N_21462,N_21912);
and U22722 (N_22722,N_21788,N_21157);
and U22723 (N_22723,N_21452,N_21724);
and U22724 (N_22724,N_21317,N_21691);
xor U22725 (N_22725,N_21015,N_21973);
nand U22726 (N_22726,N_21937,N_21188);
xnor U22727 (N_22727,N_21846,N_21815);
nor U22728 (N_22728,N_21761,N_21038);
or U22729 (N_22729,N_21671,N_21180);
nand U22730 (N_22730,N_21055,N_21667);
nor U22731 (N_22731,N_21545,N_21891);
and U22732 (N_22732,N_21805,N_21060);
or U22733 (N_22733,N_21677,N_21997);
or U22734 (N_22734,N_21305,N_21284);
and U22735 (N_22735,N_21409,N_21471);
nor U22736 (N_22736,N_21659,N_21808);
or U22737 (N_22737,N_21309,N_21329);
and U22738 (N_22738,N_21361,N_21754);
nand U22739 (N_22739,N_21226,N_21717);
nor U22740 (N_22740,N_21983,N_21687);
or U22741 (N_22741,N_21507,N_21356);
and U22742 (N_22742,N_21240,N_21972);
nor U22743 (N_22743,N_21749,N_21599);
xnor U22744 (N_22744,N_21411,N_21156);
nor U22745 (N_22745,N_21355,N_21939);
and U22746 (N_22746,N_21236,N_21446);
or U22747 (N_22747,N_21249,N_21317);
nor U22748 (N_22748,N_21664,N_21644);
nor U22749 (N_22749,N_21147,N_21846);
xor U22750 (N_22750,N_21594,N_21821);
nand U22751 (N_22751,N_21713,N_21846);
nor U22752 (N_22752,N_21021,N_21999);
nor U22753 (N_22753,N_21060,N_21441);
xnor U22754 (N_22754,N_21202,N_21236);
nor U22755 (N_22755,N_21000,N_21835);
nor U22756 (N_22756,N_21845,N_21856);
and U22757 (N_22757,N_21689,N_21642);
nand U22758 (N_22758,N_21238,N_21120);
xnor U22759 (N_22759,N_21854,N_21534);
or U22760 (N_22760,N_21931,N_21890);
nand U22761 (N_22761,N_21174,N_21941);
and U22762 (N_22762,N_21649,N_21045);
or U22763 (N_22763,N_21985,N_21480);
xor U22764 (N_22764,N_21373,N_21998);
nor U22765 (N_22765,N_21255,N_21123);
or U22766 (N_22766,N_21825,N_21373);
and U22767 (N_22767,N_21843,N_21497);
and U22768 (N_22768,N_21125,N_21251);
xor U22769 (N_22769,N_21833,N_21247);
or U22770 (N_22770,N_21672,N_21209);
nand U22771 (N_22771,N_21471,N_21779);
and U22772 (N_22772,N_21351,N_21872);
or U22773 (N_22773,N_21110,N_21216);
xnor U22774 (N_22774,N_21886,N_21905);
xnor U22775 (N_22775,N_21397,N_21178);
and U22776 (N_22776,N_21054,N_21090);
or U22777 (N_22777,N_21972,N_21316);
xor U22778 (N_22778,N_21414,N_21313);
nand U22779 (N_22779,N_21193,N_21113);
and U22780 (N_22780,N_21196,N_21592);
nand U22781 (N_22781,N_21522,N_21385);
or U22782 (N_22782,N_21110,N_21475);
or U22783 (N_22783,N_21071,N_21148);
nand U22784 (N_22784,N_21312,N_21836);
nor U22785 (N_22785,N_21673,N_21232);
nor U22786 (N_22786,N_21639,N_21333);
xor U22787 (N_22787,N_21595,N_21289);
or U22788 (N_22788,N_21385,N_21921);
nor U22789 (N_22789,N_21126,N_21366);
and U22790 (N_22790,N_21338,N_21360);
nand U22791 (N_22791,N_21608,N_21590);
or U22792 (N_22792,N_21572,N_21805);
and U22793 (N_22793,N_21852,N_21033);
nand U22794 (N_22794,N_21089,N_21644);
nand U22795 (N_22795,N_21274,N_21987);
nor U22796 (N_22796,N_21508,N_21381);
or U22797 (N_22797,N_21844,N_21255);
and U22798 (N_22798,N_21092,N_21870);
or U22799 (N_22799,N_21948,N_21171);
xor U22800 (N_22800,N_21004,N_21459);
xnor U22801 (N_22801,N_21455,N_21865);
nor U22802 (N_22802,N_21055,N_21160);
or U22803 (N_22803,N_21845,N_21761);
or U22804 (N_22804,N_21192,N_21176);
and U22805 (N_22805,N_21593,N_21461);
and U22806 (N_22806,N_21688,N_21161);
or U22807 (N_22807,N_21520,N_21348);
or U22808 (N_22808,N_21284,N_21120);
xor U22809 (N_22809,N_21881,N_21754);
or U22810 (N_22810,N_21766,N_21065);
nor U22811 (N_22811,N_21261,N_21646);
and U22812 (N_22812,N_21778,N_21518);
xnor U22813 (N_22813,N_21494,N_21199);
and U22814 (N_22814,N_21547,N_21216);
nor U22815 (N_22815,N_21885,N_21317);
nand U22816 (N_22816,N_21535,N_21775);
nand U22817 (N_22817,N_21005,N_21543);
and U22818 (N_22818,N_21967,N_21962);
and U22819 (N_22819,N_21679,N_21226);
xnor U22820 (N_22820,N_21485,N_21256);
or U22821 (N_22821,N_21115,N_21555);
nor U22822 (N_22822,N_21226,N_21071);
nand U22823 (N_22823,N_21453,N_21065);
nor U22824 (N_22824,N_21157,N_21709);
or U22825 (N_22825,N_21842,N_21397);
nand U22826 (N_22826,N_21080,N_21173);
nor U22827 (N_22827,N_21127,N_21052);
and U22828 (N_22828,N_21475,N_21757);
xor U22829 (N_22829,N_21620,N_21848);
xor U22830 (N_22830,N_21920,N_21937);
nor U22831 (N_22831,N_21397,N_21045);
and U22832 (N_22832,N_21462,N_21053);
nand U22833 (N_22833,N_21942,N_21509);
and U22834 (N_22834,N_21471,N_21012);
xnor U22835 (N_22835,N_21873,N_21231);
and U22836 (N_22836,N_21046,N_21369);
and U22837 (N_22837,N_21217,N_21983);
xor U22838 (N_22838,N_21517,N_21960);
xnor U22839 (N_22839,N_21227,N_21494);
and U22840 (N_22840,N_21649,N_21408);
nor U22841 (N_22841,N_21760,N_21144);
and U22842 (N_22842,N_21015,N_21489);
nor U22843 (N_22843,N_21349,N_21232);
or U22844 (N_22844,N_21047,N_21457);
and U22845 (N_22845,N_21647,N_21858);
nand U22846 (N_22846,N_21728,N_21717);
xor U22847 (N_22847,N_21047,N_21057);
nand U22848 (N_22848,N_21115,N_21297);
xor U22849 (N_22849,N_21957,N_21190);
nor U22850 (N_22850,N_21260,N_21464);
and U22851 (N_22851,N_21904,N_21475);
xnor U22852 (N_22852,N_21417,N_21259);
nand U22853 (N_22853,N_21834,N_21655);
nand U22854 (N_22854,N_21279,N_21738);
or U22855 (N_22855,N_21907,N_21581);
nor U22856 (N_22856,N_21951,N_21953);
nand U22857 (N_22857,N_21519,N_21915);
nand U22858 (N_22858,N_21051,N_21269);
xor U22859 (N_22859,N_21757,N_21392);
and U22860 (N_22860,N_21231,N_21493);
or U22861 (N_22861,N_21433,N_21474);
nor U22862 (N_22862,N_21522,N_21815);
and U22863 (N_22863,N_21046,N_21271);
and U22864 (N_22864,N_21945,N_21847);
nand U22865 (N_22865,N_21863,N_21409);
nor U22866 (N_22866,N_21712,N_21378);
and U22867 (N_22867,N_21698,N_21915);
or U22868 (N_22868,N_21031,N_21160);
nor U22869 (N_22869,N_21068,N_21088);
or U22870 (N_22870,N_21431,N_21944);
xor U22871 (N_22871,N_21376,N_21450);
xnor U22872 (N_22872,N_21767,N_21098);
nand U22873 (N_22873,N_21896,N_21979);
xnor U22874 (N_22874,N_21277,N_21612);
nor U22875 (N_22875,N_21799,N_21585);
and U22876 (N_22876,N_21991,N_21341);
and U22877 (N_22877,N_21233,N_21328);
and U22878 (N_22878,N_21876,N_21886);
nor U22879 (N_22879,N_21629,N_21182);
nor U22880 (N_22880,N_21252,N_21221);
xnor U22881 (N_22881,N_21753,N_21795);
xor U22882 (N_22882,N_21421,N_21776);
and U22883 (N_22883,N_21854,N_21937);
xor U22884 (N_22884,N_21842,N_21408);
nand U22885 (N_22885,N_21088,N_21377);
nor U22886 (N_22886,N_21677,N_21487);
nand U22887 (N_22887,N_21972,N_21253);
xor U22888 (N_22888,N_21174,N_21390);
and U22889 (N_22889,N_21394,N_21783);
or U22890 (N_22890,N_21570,N_21167);
and U22891 (N_22891,N_21302,N_21939);
nand U22892 (N_22892,N_21117,N_21175);
xnor U22893 (N_22893,N_21513,N_21063);
or U22894 (N_22894,N_21435,N_21440);
or U22895 (N_22895,N_21876,N_21563);
and U22896 (N_22896,N_21441,N_21785);
xor U22897 (N_22897,N_21167,N_21340);
nor U22898 (N_22898,N_21228,N_21591);
or U22899 (N_22899,N_21774,N_21692);
nand U22900 (N_22900,N_21044,N_21370);
nand U22901 (N_22901,N_21520,N_21217);
and U22902 (N_22902,N_21834,N_21439);
xnor U22903 (N_22903,N_21162,N_21098);
nand U22904 (N_22904,N_21300,N_21228);
xor U22905 (N_22905,N_21115,N_21049);
nor U22906 (N_22906,N_21813,N_21290);
and U22907 (N_22907,N_21152,N_21320);
or U22908 (N_22908,N_21034,N_21254);
nand U22909 (N_22909,N_21150,N_21408);
and U22910 (N_22910,N_21666,N_21655);
and U22911 (N_22911,N_21081,N_21135);
xnor U22912 (N_22912,N_21602,N_21721);
and U22913 (N_22913,N_21180,N_21093);
or U22914 (N_22914,N_21054,N_21468);
nand U22915 (N_22915,N_21290,N_21986);
xor U22916 (N_22916,N_21971,N_21101);
and U22917 (N_22917,N_21515,N_21209);
nor U22918 (N_22918,N_21458,N_21349);
or U22919 (N_22919,N_21396,N_21104);
and U22920 (N_22920,N_21722,N_21694);
or U22921 (N_22921,N_21235,N_21381);
nor U22922 (N_22922,N_21002,N_21116);
xor U22923 (N_22923,N_21999,N_21329);
xnor U22924 (N_22924,N_21615,N_21845);
nand U22925 (N_22925,N_21522,N_21342);
xor U22926 (N_22926,N_21362,N_21320);
nand U22927 (N_22927,N_21073,N_21000);
xor U22928 (N_22928,N_21304,N_21353);
nor U22929 (N_22929,N_21811,N_21555);
nor U22930 (N_22930,N_21089,N_21408);
nand U22931 (N_22931,N_21986,N_21649);
xor U22932 (N_22932,N_21765,N_21065);
or U22933 (N_22933,N_21255,N_21870);
nor U22934 (N_22934,N_21173,N_21381);
xnor U22935 (N_22935,N_21249,N_21931);
or U22936 (N_22936,N_21562,N_21250);
xnor U22937 (N_22937,N_21836,N_21765);
or U22938 (N_22938,N_21971,N_21386);
nor U22939 (N_22939,N_21158,N_21943);
nand U22940 (N_22940,N_21720,N_21429);
and U22941 (N_22941,N_21963,N_21253);
nor U22942 (N_22942,N_21829,N_21597);
or U22943 (N_22943,N_21121,N_21681);
nand U22944 (N_22944,N_21546,N_21761);
xor U22945 (N_22945,N_21153,N_21274);
nor U22946 (N_22946,N_21356,N_21915);
xnor U22947 (N_22947,N_21482,N_21253);
xor U22948 (N_22948,N_21810,N_21449);
xor U22949 (N_22949,N_21379,N_21953);
or U22950 (N_22950,N_21006,N_21559);
nor U22951 (N_22951,N_21288,N_21053);
nor U22952 (N_22952,N_21255,N_21017);
nor U22953 (N_22953,N_21459,N_21958);
or U22954 (N_22954,N_21260,N_21653);
or U22955 (N_22955,N_21568,N_21940);
or U22956 (N_22956,N_21213,N_21383);
or U22957 (N_22957,N_21975,N_21954);
or U22958 (N_22958,N_21836,N_21496);
nor U22959 (N_22959,N_21529,N_21724);
nor U22960 (N_22960,N_21863,N_21085);
nor U22961 (N_22961,N_21895,N_21841);
xor U22962 (N_22962,N_21211,N_21242);
nor U22963 (N_22963,N_21402,N_21215);
xnor U22964 (N_22964,N_21557,N_21511);
and U22965 (N_22965,N_21927,N_21854);
nor U22966 (N_22966,N_21326,N_21378);
nand U22967 (N_22967,N_21143,N_21570);
nand U22968 (N_22968,N_21114,N_21642);
or U22969 (N_22969,N_21900,N_21494);
or U22970 (N_22970,N_21699,N_21374);
and U22971 (N_22971,N_21355,N_21354);
xor U22972 (N_22972,N_21320,N_21959);
or U22973 (N_22973,N_21691,N_21931);
or U22974 (N_22974,N_21043,N_21084);
nor U22975 (N_22975,N_21505,N_21467);
or U22976 (N_22976,N_21355,N_21491);
nand U22977 (N_22977,N_21450,N_21400);
nand U22978 (N_22978,N_21477,N_21425);
nand U22979 (N_22979,N_21451,N_21642);
xor U22980 (N_22980,N_21075,N_21781);
xnor U22981 (N_22981,N_21277,N_21530);
xnor U22982 (N_22982,N_21625,N_21285);
nor U22983 (N_22983,N_21818,N_21910);
nand U22984 (N_22984,N_21854,N_21548);
nand U22985 (N_22985,N_21740,N_21998);
xnor U22986 (N_22986,N_21983,N_21287);
xor U22987 (N_22987,N_21465,N_21089);
nor U22988 (N_22988,N_21370,N_21813);
or U22989 (N_22989,N_21402,N_21908);
and U22990 (N_22990,N_21999,N_21342);
nor U22991 (N_22991,N_21401,N_21411);
nor U22992 (N_22992,N_21320,N_21018);
and U22993 (N_22993,N_21384,N_21474);
or U22994 (N_22994,N_21692,N_21812);
and U22995 (N_22995,N_21726,N_21621);
xor U22996 (N_22996,N_21116,N_21535);
or U22997 (N_22997,N_21045,N_21654);
nor U22998 (N_22998,N_21538,N_21410);
and U22999 (N_22999,N_21971,N_21856);
nor U23000 (N_23000,N_22674,N_22041);
or U23001 (N_23001,N_22425,N_22679);
and U23002 (N_23002,N_22358,N_22624);
or U23003 (N_23003,N_22652,N_22946);
or U23004 (N_23004,N_22701,N_22743);
nor U23005 (N_23005,N_22825,N_22289);
nand U23006 (N_23006,N_22308,N_22860);
nand U23007 (N_23007,N_22572,N_22996);
xnor U23008 (N_23008,N_22299,N_22565);
or U23009 (N_23009,N_22536,N_22325);
and U23010 (N_23010,N_22011,N_22907);
nand U23011 (N_23011,N_22801,N_22886);
xor U23012 (N_23012,N_22528,N_22714);
nor U23013 (N_23013,N_22274,N_22884);
nor U23014 (N_23014,N_22779,N_22715);
nand U23015 (N_23015,N_22310,N_22874);
or U23016 (N_23016,N_22066,N_22157);
nor U23017 (N_23017,N_22344,N_22955);
xnor U23018 (N_23018,N_22669,N_22204);
xor U23019 (N_23019,N_22768,N_22290);
and U23020 (N_23020,N_22340,N_22795);
nand U23021 (N_23021,N_22793,N_22196);
xor U23022 (N_23022,N_22977,N_22003);
or U23023 (N_23023,N_22038,N_22058);
nor U23024 (N_23024,N_22747,N_22691);
or U23025 (N_23025,N_22685,N_22297);
nand U23026 (N_23026,N_22769,N_22116);
nand U23027 (N_23027,N_22931,N_22987);
and U23028 (N_23028,N_22170,N_22859);
nor U23029 (N_23029,N_22489,N_22929);
nand U23030 (N_23030,N_22141,N_22903);
nand U23031 (N_23031,N_22756,N_22577);
xor U23032 (N_23032,N_22850,N_22269);
xnor U23033 (N_23033,N_22229,N_22730);
nand U23034 (N_23034,N_22953,N_22608);
nand U23035 (N_23035,N_22702,N_22542);
and U23036 (N_23036,N_22605,N_22316);
and U23037 (N_23037,N_22879,N_22478);
or U23038 (N_23038,N_22321,N_22905);
nand U23039 (N_23039,N_22045,N_22128);
nor U23040 (N_23040,N_22546,N_22544);
nor U23041 (N_23041,N_22262,N_22418);
nor U23042 (N_23042,N_22979,N_22354);
nand U23043 (N_23043,N_22563,N_22307);
or U23044 (N_23044,N_22463,N_22593);
or U23045 (N_23045,N_22926,N_22798);
xor U23046 (N_23046,N_22503,N_22488);
nand U23047 (N_23047,N_22723,N_22149);
nand U23048 (N_23048,N_22568,N_22194);
and U23049 (N_23049,N_22688,N_22604);
xor U23050 (N_23050,N_22981,N_22915);
nor U23051 (N_23051,N_22689,N_22687);
xor U23052 (N_23052,N_22295,N_22312);
or U23053 (N_23053,N_22439,N_22826);
or U23054 (N_23054,N_22921,N_22322);
xnor U23055 (N_23055,N_22384,N_22147);
or U23056 (N_23056,N_22390,N_22518);
nand U23057 (N_23057,N_22595,N_22772);
or U23058 (N_23058,N_22615,N_22783);
nor U23059 (N_23059,N_22517,N_22805);
xor U23060 (N_23060,N_22190,N_22240);
and U23061 (N_23061,N_22751,N_22569);
nor U23062 (N_23062,N_22121,N_22006);
xor U23063 (N_23063,N_22893,N_22001);
or U23064 (N_23064,N_22386,N_22252);
nor U23065 (N_23065,N_22725,N_22978);
xor U23066 (N_23066,N_22416,N_22298);
nand U23067 (N_23067,N_22245,N_22070);
xor U23068 (N_23068,N_22823,N_22509);
nor U23069 (N_23069,N_22830,N_22985);
and U23070 (N_23070,N_22056,N_22704);
and U23071 (N_23071,N_22403,N_22226);
nand U23072 (N_23072,N_22242,N_22109);
xnor U23073 (N_23073,N_22369,N_22382);
nor U23074 (N_23074,N_22952,N_22136);
nor U23075 (N_23075,N_22510,N_22100);
nand U23076 (N_23076,N_22502,N_22639);
or U23077 (N_23077,N_22039,N_22426);
nand U23078 (N_23078,N_22071,N_22318);
nor U23079 (N_23079,N_22500,N_22827);
and U23080 (N_23080,N_22256,N_22734);
nand U23081 (N_23081,N_22838,N_22590);
xor U23082 (N_23082,N_22917,N_22219);
and U23083 (N_23083,N_22789,N_22048);
and U23084 (N_23084,N_22806,N_22005);
xor U23085 (N_23085,N_22753,N_22947);
and U23086 (N_23086,N_22068,N_22847);
nand U23087 (N_23087,N_22394,N_22641);
nor U23088 (N_23088,N_22144,N_22995);
or U23089 (N_23089,N_22705,N_22437);
or U23090 (N_23090,N_22207,N_22677);
or U23091 (N_23091,N_22026,N_22537);
nand U23092 (N_23092,N_22267,N_22078);
nand U23093 (N_23093,N_22336,N_22868);
nor U23094 (N_23094,N_22765,N_22417);
nor U23095 (N_23095,N_22086,N_22460);
and U23096 (N_23096,N_22928,N_22800);
nor U23097 (N_23097,N_22130,N_22694);
or U23098 (N_23098,N_22529,N_22139);
and U23099 (N_23099,N_22986,N_22348);
nor U23100 (N_23100,N_22212,N_22659);
nand U23101 (N_23101,N_22012,N_22650);
nor U23102 (N_23102,N_22712,N_22771);
and U23103 (N_23103,N_22970,N_22623);
or U23104 (N_23104,N_22328,N_22232);
nand U23105 (N_23105,N_22958,N_22525);
and U23106 (N_23106,N_22966,N_22738);
xor U23107 (N_23107,N_22633,N_22904);
nor U23108 (N_23108,N_22832,N_22241);
nand U23109 (N_23109,N_22627,N_22167);
or U23110 (N_23110,N_22023,N_22551);
xor U23111 (N_23111,N_22151,N_22531);
or U23112 (N_23112,N_22468,N_22575);
and U23113 (N_23113,N_22837,N_22341);
and U23114 (N_23114,N_22203,N_22483);
nand U23115 (N_23115,N_22560,N_22492);
xnor U23116 (N_23116,N_22137,N_22927);
and U23117 (N_23117,N_22337,N_22871);
or U23118 (N_23118,N_22494,N_22506);
or U23119 (N_23119,N_22469,N_22745);
nand U23120 (N_23120,N_22866,N_22960);
or U23121 (N_23121,N_22522,N_22213);
xnor U23122 (N_23122,N_22018,N_22201);
nor U23123 (N_23123,N_22813,N_22414);
nand U23124 (N_23124,N_22407,N_22710);
nor U23125 (N_23125,N_22236,N_22657);
nand U23126 (N_23126,N_22067,N_22278);
nand U23127 (N_23127,N_22935,N_22719);
nor U23128 (N_23128,N_22357,N_22102);
and U23129 (N_23129,N_22916,N_22740);
nand U23130 (N_23130,N_22622,N_22788);
nor U23131 (N_23131,N_22748,N_22746);
nand U23132 (N_23132,N_22853,N_22690);
nand U23133 (N_23133,N_22974,N_22431);
or U23134 (N_23134,N_22762,N_22470);
and U23135 (N_23135,N_22754,N_22975);
xor U23136 (N_23136,N_22291,N_22261);
or U23137 (N_23137,N_22392,N_22535);
nor U23138 (N_23138,N_22628,N_22890);
and U23139 (N_23139,N_22471,N_22131);
or U23140 (N_23140,N_22811,N_22758);
and U23141 (N_23141,N_22703,N_22835);
nor U23142 (N_23142,N_22984,N_22814);
nor U23143 (N_23143,N_22095,N_22294);
or U23144 (N_23144,N_22653,N_22330);
or U23145 (N_23145,N_22467,N_22664);
or U23146 (N_23146,N_22558,N_22363);
or U23147 (N_23147,N_22968,N_22179);
and U23148 (N_23148,N_22332,N_22271);
nand U23149 (N_23149,N_22776,N_22976);
xor U23150 (N_23150,N_22351,N_22303);
or U23151 (N_23151,N_22275,N_22101);
and U23152 (N_23152,N_22475,N_22942);
and U23153 (N_23153,N_22739,N_22474);
nor U23154 (N_23154,N_22352,N_22711);
or U23155 (N_23155,N_22932,N_22780);
nor U23156 (N_23156,N_22964,N_22027);
or U23157 (N_23157,N_22661,N_22925);
xnor U23158 (N_23158,N_22864,N_22146);
nand U23159 (N_23159,N_22513,N_22231);
or U23160 (N_23160,N_22698,N_22224);
xnor U23161 (N_23161,N_22446,N_22395);
and U23162 (N_23162,N_22085,N_22962);
and U23163 (N_23163,N_22276,N_22367);
and U23164 (N_23164,N_22693,N_22658);
or U23165 (N_23165,N_22611,N_22106);
and U23166 (N_23166,N_22186,N_22684);
and U23167 (N_23167,N_22616,N_22549);
and U23168 (N_23168,N_22896,N_22557);
and U23169 (N_23169,N_22949,N_22098);
nand U23170 (N_23170,N_22851,N_22237);
or U23171 (N_23171,N_22377,N_22075);
nor U23172 (N_23172,N_22279,N_22620);
nor U23173 (N_23173,N_22234,N_22586);
xor U23174 (N_23174,N_22302,N_22594);
nor U23175 (N_23175,N_22355,N_22857);
nor U23176 (N_23176,N_22314,N_22938);
or U23177 (N_23177,N_22877,N_22726);
and U23178 (N_23178,N_22087,N_22065);
or U23179 (N_23179,N_22326,N_22644);
nand U23180 (N_23180,N_22706,N_22514);
nor U23181 (N_23181,N_22613,N_22309);
nand U23182 (N_23182,N_22582,N_22777);
nand U23183 (N_23183,N_22254,N_22399);
nand U23184 (N_23184,N_22749,N_22466);
nand U23185 (N_23185,N_22580,N_22539);
nor U23186 (N_23186,N_22948,N_22496);
xor U23187 (N_23187,N_22831,N_22389);
nand U23188 (N_23188,N_22554,N_22767);
and U23189 (N_23189,N_22858,N_22887);
nor U23190 (N_23190,N_22797,N_22020);
or U23191 (N_23191,N_22869,N_22413);
nand U23192 (N_23192,N_22610,N_22374);
nand U23193 (N_23193,N_22770,N_22108);
xor U23194 (N_23194,N_22600,N_22404);
nor U23195 (N_23195,N_22211,N_22848);
nor U23196 (N_23196,N_22183,N_22052);
xor U23197 (N_23197,N_22880,N_22816);
nand U23198 (N_23198,N_22264,N_22516);
or U23199 (N_23199,N_22487,N_22799);
nand U23200 (N_23200,N_22526,N_22989);
xnor U23201 (N_23201,N_22579,N_22944);
xnor U23202 (N_23202,N_22251,N_22965);
nand U23203 (N_23203,N_22030,N_22368);
nand U23204 (N_23204,N_22922,N_22988);
and U23205 (N_23205,N_22364,N_22888);
nor U23206 (N_23206,N_22258,N_22126);
or U23207 (N_23207,N_22453,N_22646);
and U23208 (N_23208,N_22961,N_22440);
and U23209 (N_23209,N_22617,N_22206);
and U23210 (N_23210,N_22587,N_22187);
and U23211 (N_23211,N_22632,N_22540);
nor U23212 (N_23212,N_22521,N_22150);
or U23213 (N_23213,N_22461,N_22373);
or U23214 (N_23214,N_22457,N_22497);
xor U23215 (N_23215,N_22032,N_22643);
nor U23216 (N_23216,N_22548,N_22043);
nand U23217 (N_23217,N_22089,N_22077);
or U23218 (N_23218,N_22225,N_22459);
or U23219 (N_23219,N_22519,N_22875);
or U23220 (N_23220,N_22381,N_22550);
nor U23221 (N_23221,N_22244,N_22950);
nand U23222 (N_23222,N_22682,N_22490);
nand U23223 (N_23223,N_22235,N_22809);
nand U23224 (N_23224,N_22485,N_22385);
nand U23225 (N_23225,N_22794,N_22662);
or U23226 (N_23226,N_22882,N_22993);
nand U23227 (N_23227,N_22178,N_22499);
nor U23228 (N_23228,N_22564,N_22840);
xnor U23229 (N_23229,N_22420,N_22200);
or U23230 (N_23230,N_22443,N_22555);
nor U23231 (N_23231,N_22724,N_22156);
nor U23232 (N_23232,N_22222,N_22317);
xor U23233 (N_23233,N_22193,N_22619);
xnor U23234 (N_23234,N_22504,N_22218);
xnor U23235 (N_23235,N_22454,N_22338);
xor U23236 (N_23236,N_22073,N_22117);
nor U23237 (N_23237,N_22670,N_22473);
nand U23238 (N_23238,N_22401,N_22113);
xor U23239 (N_23239,N_22603,N_22000);
or U23240 (N_23240,N_22422,N_22982);
and U23241 (N_23241,N_22455,N_22969);
or U23242 (N_23242,N_22843,N_22940);
xnor U23243 (N_23243,N_22421,N_22876);
xnor U23244 (N_23244,N_22400,N_22596);
nand U23245 (N_23245,N_22164,N_22649);
nand U23246 (N_23246,N_22372,N_22821);
nor U23247 (N_23247,N_22849,N_22050);
xnor U23248 (N_23248,N_22356,N_22296);
nor U23249 (N_23249,N_22683,N_22119);
or U23250 (N_23250,N_22614,N_22967);
xor U23251 (N_23251,N_22054,N_22597);
nand U23252 (N_23252,N_22347,N_22692);
and U23253 (N_23253,N_22956,N_22865);
and U23254 (N_23254,N_22733,N_22450);
and U23255 (N_23255,N_22900,N_22094);
nand U23256 (N_23256,N_22076,N_22834);
nand U23257 (N_23257,N_22057,N_22323);
xor U23258 (N_23258,N_22999,N_22523);
or U23259 (N_23259,N_22124,N_22462);
and U23260 (N_23260,N_22578,N_22177);
or U23261 (N_23261,N_22430,N_22263);
nand U23262 (N_23262,N_22284,N_22479);
xnor U23263 (N_23263,N_22335,N_22943);
xnor U23264 (N_23264,N_22963,N_22663);
xnor U23265 (N_23265,N_22238,N_22375);
nand U23266 (N_23266,N_22040,N_22629);
and U23267 (N_23267,N_22447,N_22361);
and U23268 (N_23268,N_22173,N_22304);
nand U23269 (N_23269,N_22735,N_22079);
nand U23270 (N_23270,N_22423,N_22083);
nand U23271 (N_23271,N_22718,N_22306);
nand U23272 (N_23272,N_22415,N_22112);
xor U23273 (N_23273,N_22655,N_22573);
xor U23274 (N_23274,N_22675,N_22686);
and U23275 (N_23275,N_22477,N_22648);
and U23276 (N_23276,N_22438,N_22990);
nand U23277 (N_23277,N_22744,N_22665);
xor U23278 (N_23278,N_22429,N_22584);
and U23279 (N_23279,N_22750,N_22448);
or U23280 (N_23280,N_22697,N_22198);
or U23281 (N_23281,N_22366,N_22331);
or U23282 (N_23282,N_22630,N_22349);
and U23283 (N_23283,N_22640,N_22992);
and U23284 (N_23284,N_22161,N_22345);
nor U23285 (N_23285,N_22668,N_22371);
or U23286 (N_23286,N_22379,N_22634);
nor U23287 (N_23287,N_22191,N_22647);
nor U23288 (N_23288,N_22508,N_22168);
nand U23289 (N_23289,N_22773,N_22607);
nor U23290 (N_23290,N_22804,N_22120);
xnor U23291 (N_23291,N_22017,N_22515);
nand U23292 (N_23292,N_22110,N_22074);
nor U23293 (N_23293,N_22036,N_22524);
xor U23294 (N_23294,N_22288,N_22883);
nor U23295 (N_23295,N_22031,N_22913);
xor U23296 (N_23296,N_22132,N_22171);
nor U23297 (N_23297,N_22424,N_22885);
nor U23298 (N_23298,N_22599,N_22376);
xnor U23299 (N_23299,N_22727,N_22872);
nand U23300 (N_23300,N_22637,N_22656);
or U23301 (N_23301,N_22125,N_22741);
xor U23302 (N_23302,N_22181,N_22445);
xor U23303 (N_23303,N_22409,N_22383);
and U23304 (N_23304,N_22861,N_22021);
or U23305 (N_23305,N_22016,N_22362);
and U23306 (N_23306,N_22360,N_22791);
and U23307 (N_23307,N_22937,N_22760);
or U23308 (N_23308,N_22195,N_22971);
and U23309 (N_23309,N_22481,N_22035);
nand U23310 (N_23310,N_22081,N_22997);
nand U23311 (N_23311,N_22855,N_22228);
nor U23312 (N_23312,N_22166,N_22924);
nor U23313 (N_23313,N_22626,N_22681);
and U23314 (N_23314,N_22280,N_22700);
nand U23315 (N_23315,N_22583,N_22666);
nor U23316 (N_23316,N_22538,N_22396);
nand U23317 (N_23317,N_22651,N_22642);
or U23318 (N_23318,N_22895,N_22053);
nand U23319 (N_23319,N_22411,N_22327);
and U23320 (N_23320,N_22829,N_22854);
xor U23321 (N_23321,N_22220,N_22159);
nor U23322 (N_23322,N_22024,N_22778);
and U23323 (N_23323,N_22678,N_22581);
xnor U23324 (N_23324,N_22458,N_22930);
nand U23325 (N_23325,N_22870,N_22398);
nand U23326 (N_23326,N_22359,N_22350);
nor U23327 (N_23327,N_22836,N_22097);
and U23328 (N_23328,N_22918,N_22301);
xor U23329 (N_23329,N_22589,N_22602);
xor U23330 (N_23330,N_22556,N_22621);
or U23331 (N_23331,N_22285,N_22716);
nand U23332 (N_23332,N_22210,N_22954);
nor U23333 (N_23333,N_22833,N_22878);
nor U23334 (N_23334,N_22123,N_22774);
or U23335 (N_23335,N_22093,N_22239);
xor U23336 (N_23336,N_22759,N_22936);
nand U23337 (N_23337,N_22033,N_22188);
nor U23338 (N_23338,N_22208,N_22272);
nand U23339 (N_23339,N_22576,N_22215);
and U23340 (N_23340,N_22182,N_22807);
nand U23341 (N_23341,N_22742,N_22051);
nand U23342 (N_23342,N_22785,N_22585);
nor U23343 (N_23343,N_22873,N_22266);
and U23344 (N_23344,N_22015,N_22342);
and U23345 (N_23345,N_22552,N_22660);
nor U23346 (N_23346,N_22107,N_22781);
nand U23347 (N_23347,N_22625,N_22061);
or U23348 (N_23348,N_22442,N_22612);
and U23349 (N_23349,N_22636,N_22428);
xnor U23350 (N_23350,N_22209,N_22260);
and U23351 (N_23351,N_22197,N_22533);
xor U23352 (N_23352,N_22566,N_22983);
nor U23353 (N_23353,N_22072,N_22175);
xor U23354 (N_23354,N_22324,N_22911);
and U23355 (N_23355,N_22898,N_22410);
nand U23356 (N_23356,N_22062,N_22792);
and U23357 (N_23357,N_22273,N_22154);
nand U23358 (N_23358,N_22270,N_22764);
nor U23359 (N_23359,N_22717,N_22365);
nor U23360 (N_23360,N_22214,N_22129);
or U23361 (N_23361,N_22391,N_22845);
xnor U23362 (N_23362,N_22047,N_22134);
and U23363 (N_23363,N_22096,N_22484);
nor U23364 (N_23364,N_22545,N_22919);
nor U23365 (N_23365,N_22008,N_22019);
xnor U23366 (N_23366,N_22782,N_22370);
nor U23367 (N_23367,N_22894,N_22380);
nand U23368 (N_23368,N_22255,N_22311);
or U23369 (N_23369,N_22227,N_22881);
xnor U23370 (N_23370,N_22160,N_22567);
nor U23371 (N_23371,N_22223,N_22007);
or U23372 (N_23372,N_22037,N_22221);
nand U23373 (N_23373,N_22169,N_22172);
nand U23374 (N_23374,N_22755,N_22547);
nand U23375 (N_23375,N_22939,N_22432);
nor U23376 (N_23376,N_22787,N_22319);
nor U23377 (N_23377,N_22265,N_22553);
nor U23378 (N_23378,N_22064,N_22654);
or U23379 (N_23379,N_22511,N_22444);
nand U23380 (N_23380,N_22722,N_22456);
xor U23381 (N_23381,N_22165,N_22202);
or U23382 (N_23382,N_22713,N_22028);
xor U23383 (N_23383,N_22472,N_22591);
nand U23384 (N_23384,N_22757,N_22217);
nand U23385 (N_23385,N_22482,N_22574);
xnor U23386 (N_23386,N_22998,N_22084);
nand U23387 (N_23387,N_22143,N_22010);
xnor U23388 (N_23388,N_22192,N_22709);
nand U23389 (N_23389,N_22004,N_22824);
and U23390 (N_23390,N_22945,N_22029);
nand U23391 (N_23391,N_22959,N_22063);
xnor U23392 (N_23392,N_22104,N_22732);
or U23393 (N_23393,N_22696,N_22387);
nor U23394 (N_23394,N_22464,N_22699);
or U23395 (N_23395,N_22505,N_22737);
nand U23396 (N_23396,N_22598,N_22820);
nor U23397 (N_23397,N_22507,N_22320);
nand U23398 (N_23398,N_22163,N_22189);
nor U23399 (N_23399,N_22667,N_22520);
and U23400 (N_23400,N_22268,N_22761);
xnor U23401 (N_23401,N_22480,N_22818);
nand U23402 (N_23402,N_22645,N_22846);
nand U23403 (N_23403,N_22092,N_22609);
or U23404 (N_23404,N_22449,N_22088);
and U23405 (N_23405,N_22180,N_22934);
and U23406 (N_23406,N_22080,N_22991);
nor U23407 (N_23407,N_22412,N_22133);
nor U23408 (N_23408,N_22530,N_22817);
xor U23409 (N_23409,N_22819,N_22022);
nor U23410 (N_23410,N_22862,N_22592);
xnor U23411 (N_23411,N_22973,N_22333);
or U23412 (N_23412,N_22631,N_22909);
nand U23413 (N_23413,N_22436,N_22728);
nand U23414 (N_23414,N_22863,N_22434);
and U23415 (N_23415,N_22543,N_22707);
and U23416 (N_23416,N_22287,N_22844);
and U23417 (N_23417,N_22841,N_22099);
or U23418 (N_23418,N_22090,N_22891);
nand U23419 (N_23419,N_22148,N_22752);
xnor U23420 (N_23420,N_22406,N_22281);
and U23421 (N_23421,N_22378,N_22082);
nand U23422 (N_23422,N_22638,N_22671);
and U23423 (N_23423,N_22114,N_22541);
nand U23424 (N_23424,N_22796,N_22812);
and U23425 (N_23425,N_22142,N_22618);
or U23426 (N_23426,N_22115,N_22532);
and U23427 (N_23427,N_22118,N_22127);
or U23428 (N_23428,N_22914,N_22230);
xnor U23429 (N_23429,N_22736,N_22512);
xnor U23430 (N_23430,N_22339,N_22185);
nor U23431 (N_23431,N_22721,N_22353);
xnor U23432 (N_23432,N_22920,N_22451);
nand U23433 (N_23433,N_22111,N_22606);
and U23434 (N_23434,N_22695,N_22912);
xor U23435 (N_23435,N_22486,N_22889);
xor U23436 (N_23436,N_22972,N_22559);
nor U23437 (N_23437,N_22784,N_22676);
and U23438 (N_23438,N_22534,N_22562);
nand U23439 (N_23439,N_22014,N_22763);
and U23440 (N_23440,N_22002,N_22828);
nand U23441 (N_23441,N_22305,N_22892);
or U23442 (N_23442,N_22122,N_22049);
nor U23443 (N_23443,N_22465,N_22923);
nor U23444 (N_23444,N_22034,N_22205);
xor U23445 (N_23445,N_22672,N_22315);
or U23446 (N_23446,N_22902,N_22055);
and U23447 (N_23447,N_22174,N_22046);
xnor U23448 (N_23448,N_22527,N_22493);
xnor U23449 (N_23449,N_22729,N_22571);
xnor U23450 (N_23450,N_22588,N_22060);
or U23451 (N_23451,N_22491,N_22293);
xor U23452 (N_23452,N_22334,N_22994);
and U23453 (N_23453,N_22158,N_22561);
nor U23454 (N_23454,N_22257,N_22808);
nor U23455 (N_23455,N_22856,N_22906);
nor U23456 (N_23456,N_22250,N_22405);
and U23457 (N_23457,N_22495,N_22790);
and U23458 (N_23458,N_22408,N_22140);
xnor U23459 (N_23459,N_22815,N_22277);
and U23460 (N_23460,N_22822,N_22803);
nor U23461 (N_23461,N_22397,N_22313);
xor U23462 (N_23462,N_22680,N_22708);
nor U23463 (N_23463,N_22957,N_22498);
nor U23464 (N_23464,N_22908,N_22091);
nand U23465 (N_23465,N_22282,N_22259);
and U23466 (N_23466,N_22145,N_22673);
xor U23467 (N_23467,N_22388,N_22009);
and U23468 (N_23468,N_22199,N_22899);
or U23469 (N_23469,N_22980,N_22842);
xnor U23470 (N_23470,N_22138,N_22135);
nor U23471 (N_23471,N_22419,N_22720);
nor U23472 (N_23472,N_22393,N_22802);
and U23473 (N_23473,N_22103,N_22184);
nand U23474 (N_23474,N_22852,N_22402);
nand U23475 (N_23475,N_22300,N_22233);
xnor U23476 (N_23476,N_22933,N_22283);
nand U23477 (N_23477,N_22044,N_22501);
xor U23478 (N_23478,N_22247,N_22941);
xnor U23479 (N_23479,N_22476,N_22152);
nand U23480 (N_23480,N_22570,N_22059);
nor U23481 (N_23481,N_22013,N_22153);
xor U23482 (N_23482,N_22427,N_22775);
or U23483 (N_23483,N_22246,N_22329);
and U23484 (N_23484,N_22910,N_22731);
xor U23485 (N_23485,N_22105,N_22601);
nor U23486 (N_23486,N_22216,N_22786);
and U23487 (N_23487,N_22635,N_22249);
nor U23488 (N_23488,N_22243,N_22839);
and U23489 (N_23489,N_22286,N_22176);
xnor U23490 (N_23490,N_22441,N_22025);
and U23491 (N_23491,N_22901,N_22042);
or U23492 (N_23492,N_22897,N_22766);
or U23493 (N_23493,N_22951,N_22433);
and U23494 (N_23494,N_22253,N_22346);
nor U23495 (N_23495,N_22867,N_22069);
nor U23496 (N_23496,N_22248,N_22452);
nor U23497 (N_23497,N_22292,N_22343);
and U23498 (N_23498,N_22155,N_22162);
xor U23499 (N_23499,N_22810,N_22435);
and U23500 (N_23500,N_22722,N_22162);
or U23501 (N_23501,N_22047,N_22419);
xnor U23502 (N_23502,N_22090,N_22359);
and U23503 (N_23503,N_22303,N_22685);
nand U23504 (N_23504,N_22566,N_22329);
xnor U23505 (N_23505,N_22941,N_22848);
or U23506 (N_23506,N_22410,N_22738);
nor U23507 (N_23507,N_22909,N_22551);
nor U23508 (N_23508,N_22879,N_22083);
nor U23509 (N_23509,N_22438,N_22627);
xor U23510 (N_23510,N_22072,N_22972);
xor U23511 (N_23511,N_22299,N_22989);
and U23512 (N_23512,N_22084,N_22578);
or U23513 (N_23513,N_22157,N_22445);
nor U23514 (N_23514,N_22232,N_22819);
or U23515 (N_23515,N_22180,N_22048);
and U23516 (N_23516,N_22677,N_22342);
or U23517 (N_23517,N_22108,N_22045);
or U23518 (N_23518,N_22415,N_22695);
xor U23519 (N_23519,N_22965,N_22264);
or U23520 (N_23520,N_22991,N_22153);
and U23521 (N_23521,N_22802,N_22618);
nor U23522 (N_23522,N_22114,N_22425);
nor U23523 (N_23523,N_22678,N_22224);
nor U23524 (N_23524,N_22668,N_22742);
or U23525 (N_23525,N_22085,N_22345);
nand U23526 (N_23526,N_22740,N_22601);
xor U23527 (N_23527,N_22417,N_22116);
and U23528 (N_23528,N_22548,N_22579);
and U23529 (N_23529,N_22682,N_22888);
nor U23530 (N_23530,N_22095,N_22549);
nand U23531 (N_23531,N_22720,N_22754);
xor U23532 (N_23532,N_22591,N_22509);
nand U23533 (N_23533,N_22440,N_22937);
nor U23534 (N_23534,N_22426,N_22055);
and U23535 (N_23535,N_22439,N_22847);
nor U23536 (N_23536,N_22033,N_22517);
nor U23537 (N_23537,N_22378,N_22633);
nand U23538 (N_23538,N_22355,N_22739);
nor U23539 (N_23539,N_22140,N_22775);
and U23540 (N_23540,N_22374,N_22289);
nor U23541 (N_23541,N_22099,N_22641);
and U23542 (N_23542,N_22315,N_22701);
or U23543 (N_23543,N_22425,N_22948);
xor U23544 (N_23544,N_22593,N_22263);
xor U23545 (N_23545,N_22421,N_22962);
xnor U23546 (N_23546,N_22833,N_22971);
and U23547 (N_23547,N_22924,N_22100);
nand U23548 (N_23548,N_22303,N_22175);
and U23549 (N_23549,N_22459,N_22920);
or U23550 (N_23550,N_22157,N_22404);
and U23551 (N_23551,N_22023,N_22894);
nor U23552 (N_23552,N_22606,N_22555);
and U23553 (N_23553,N_22739,N_22361);
and U23554 (N_23554,N_22435,N_22212);
and U23555 (N_23555,N_22140,N_22161);
and U23556 (N_23556,N_22565,N_22869);
and U23557 (N_23557,N_22368,N_22076);
or U23558 (N_23558,N_22541,N_22276);
and U23559 (N_23559,N_22126,N_22792);
nor U23560 (N_23560,N_22653,N_22981);
nor U23561 (N_23561,N_22641,N_22537);
or U23562 (N_23562,N_22354,N_22850);
nor U23563 (N_23563,N_22225,N_22594);
nor U23564 (N_23564,N_22596,N_22869);
or U23565 (N_23565,N_22098,N_22863);
nor U23566 (N_23566,N_22004,N_22877);
nand U23567 (N_23567,N_22684,N_22487);
nand U23568 (N_23568,N_22959,N_22096);
or U23569 (N_23569,N_22064,N_22358);
xor U23570 (N_23570,N_22456,N_22715);
nor U23571 (N_23571,N_22749,N_22722);
nor U23572 (N_23572,N_22273,N_22576);
or U23573 (N_23573,N_22624,N_22265);
xnor U23574 (N_23574,N_22781,N_22833);
nor U23575 (N_23575,N_22297,N_22436);
nand U23576 (N_23576,N_22155,N_22779);
or U23577 (N_23577,N_22987,N_22528);
nand U23578 (N_23578,N_22162,N_22387);
nand U23579 (N_23579,N_22901,N_22096);
and U23580 (N_23580,N_22917,N_22587);
xor U23581 (N_23581,N_22944,N_22094);
nand U23582 (N_23582,N_22009,N_22521);
xnor U23583 (N_23583,N_22228,N_22420);
nand U23584 (N_23584,N_22889,N_22652);
or U23585 (N_23585,N_22152,N_22023);
nor U23586 (N_23586,N_22439,N_22823);
nor U23587 (N_23587,N_22153,N_22516);
xnor U23588 (N_23588,N_22885,N_22507);
nand U23589 (N_23589,N_22980,N_22540);
and U23590 (N_23590,N_22485,N_22805);
nand U23591 (N_23591,N_22169,N_22640);
nor U23592 (N_23592,N_22076,N_22475);
nand U23593 (N_23593,N_22422,N_22374);
xor U23594 (N_23594,N_22099,N_22680);
or U23595 (N_23595,N_22808,N_22977);
or U23596 (N_23596,N_22738,N_22661);
nand U23597 (N_23597,N_22069,N_22182);
nor U23598 (N_23598,N_22130,N_22380);
or U23599 (N_23599,N_22251,N_22178);
xnor U23600 (N_23600,N_22390,N_22735);
xnor U23601 (N_23601,N_22543,N_22257);
nor U23602 (N_23602,N_22965,N_22154);
xor U23603 (N_23603,N_22304,N_22777);
or U23604 (N_23604,N_22073,N_22891);
xor U23605 (N_23605,N_22955,N_22100);
or U23606 (N_23606,N_22641,N_22521);
nand U23607 (N_23607,N_22569,N_22132);
xor U23608 (N_23608,N_22444,N_22571);
nand U23609 (N_23609,N_22428,N_22322);
nand U23610 (N_23610,N_22216,N_22793);
or U23611 (N_23611,N_22192,N_22861);
or U23612 (N_23612,N_22779,N_22922);
xor U23613 (N_23613,N_22600,N_22082);
or U23614 (N_23614,N_22850,N_22648);
nor U23615 (N_23615,N_22541,N_22291);
and U23616 (N_23616,N_22147,N_22576);
nor U23617 (N_23617,N_22285,N_22181);
xnor U23618 (N_23618,N_22190,N_22153);
and U23619 (N_23619,N_22921,N_22205);
and U23620 (N_23620,N_22232,N_22073);
and U23621 (N_23621,N_22948,N_22063);
nand U23622 (N_23622,N_22478,N_22883);
nand U23623 (N_23623,N_22787,N_22867);
and U23624 (N_23624,N_22386,N_22097);
or U23625 (N_23625,N_22827,N_22840);
and U23626 (N_23626,N_22560,N_22536);
xnor U23627 (N_23627,N_22355,N_22114);
or U23628 (N_23628,N_22754,N_22426);
and U23629 (N_23629,N_22312,N_22888);
and U23630 (N_23630,N_22756,N_22113);
or U23631 (N_23631,N_22745,N_22162);
and U23632 (N_23632,N_22241,N_22819);
or U23633 (N_23633,N_22889,N_22820);
or U23634 (N_23634,N_22580,N_22815);
nor U23635 (N_23635,N_22103,N_22484);
and U23636 (N_23636,N_22246,N_22765);
xnor U23637 (N_23637,N_22924,N_22071);
and U23638 (N_23638,N_22257,N_22422);
or U23639 (N_23639,N_22167,N_22030);
nand U23640 (N_23640,N_22801,N_22288);
or U23641 (N_23641,N_22006,N_22744);
and U23642 (N_23642,N_22533,N_22510);
xor U23643 (N_23643,N_22511,N_22202);
and U23644 (N_23644,N_22902,N_22754);
and U23645 (N_23645,N_22616,N_22460);
xnor U23646 (N_23646,N_22802,N_22037);
nor U23647 (N_23647,N_22932,N_22018);
nor U23648 (N_23648,N_22469,N_22292);
nor U23649 (N_23649,N_22973,N_22078);
nand U23650 (N_23650,N_22371,N_22248);
nor U23651 (N_23651,N_22611,N_22830);
xor U23652 (N_23652,N_22393,N_22981);
nand U23653 (N_23653,N_22702,N_22739);
and U23654 (N_23654,N_22031,N_22666);
nand U23655 (N_23655,N_22834,N_22289);
or U23656 (N_23656,N_22243,N_22933);
and U23657 (N_23657,N_22199,N_22555);
nor U23658 (N_23658,N_22689,N_22505);
nand U23659 (N_23659,N_22561,N_22284);
and U23660 (N_23660,N_22652,N_22410);
or U23661 (N_23661,N_22798,N_22529);
xor U23662 (N_23662,N_22653,N_22234);
xor U23663 (N_23663,N_22192,N_22505);
xnor U23664 (N_23664,N_22757,N_22516);
and U23665 (N_23665,N_22452,N_22250);
xor U23666 (N_23666,N_22629,N_22105);
or U23667 (N_23667,N_22155,N_22114);
and U23668 (N_23668,N_22200,N_22982);
and U23669 (N_23669,N_22528,N_22518);
or U23670 (N_23670,N_22304,N_22685);
nand U23671 (N_23671,N_22191,N_22139);
nand U23672 (N_23672,N_22111,N_22712);
nand U23673 (N_23673,N_22881,N_22713);
nor U23674 (N_23674,N_22195,N_22457);
and U23675 (N_23675,N_22792,N_22509);
and U23676 (N_23676,N_22892,N_22537);
or U23677 (N_23677,N_22973,N_22958);
or U23678 (N_23678,N_22494,N_22558);
or U23679 (N_23679,N_22947,N_22857);
or U23680 (N_23680,N_22777,N_22071);
nand U23681 (N_23681,N_22537,N_22886);
nand U23682 (N_23682,N_22367,N_22376);
nor U23683 (N_23683,N_22747,N_22251);
or U23684 (N_23684,N_22376,N_22440);
or U23685 (N_23685,N_22535,N_22506);
and U23686 (N_23686,N_22654,N_22311);
or U23687 (N_23687,N_22123,N_22026);
and U23688 (N_23688,N_22238,N_22630);
and U23689 (N_23689,N_22433,N_22321);
xnor U23690 (N_23690,N_22341,N_22186);
nand U23691 (N_23691,N_22824,N_22244);
xnor U23692 (N_23692,N_22354,N_22144);
xor U23693 (N_23693,N_22530,N_22556);
or U23694 (N_23694,N_22326,N_22181);
nand U23695 (N_23695,N_22739,N_22208);
and U23696 (N_23696,N_22061,N_22122);
or U23697 (N_23697,N_22417,N_22925);
nand U23698 (N_23698,N_22896,N_22444);
or U23699 (N_23699,N_22027,N_22903);
and U23700 (N_23700,N_22571,N_22824);
nand U23701 (N_23701,N_22420,N_22773);
nand U23702 (N_23702,N_22054,N_22551);
and U23703 (N_23703,N_22134,N_22319);
or U23704 (N_23704,N_22787,N_22003);
and U23705 (N_23705,N_22071,N_22314);
xnor U23706 (N_23706,N_22148,N_22322);
or U23707 (N_23707,N_22548,N_22697);
nor U23708 (N_23708,N_22091,N_22475);
nand U23709 (N_23709,N_22859,N_22689);
nand U23710 (N_23710,N_22260,N_22003);
and U23711 (N_23711,N_22223,N_22623);
nand U23712 (N_23712,N_22308,N_22414);
nand U23713 (N_23713,N_22457,N_22537);
nor U23714 (N_23714,N_22141,N_22463);
nand U23715 (N_23715,N_22678,N_22687);
or U23716 (N_23716,N_22381,N_22432);
nor U23717 (N_23717,N_22573,N_22306);
nor U23718 (N_23718,N_22162,N_22380);
xnor U23719 (N_23719,N_22270,N_22211);
and U23720 (N_23720,N_22070,N_22600);
nor U23721 (N_23721,N_22750,N_22216);
and U23722 (N_23722,N_22793,N_22052);
nor U23723 (N_23723,N_22147,N_22786);
nor U23724 (N_23724,N_22971,N_22291);
or U23725 (N_23725,N_22010,N_22051);
nand U23726 (N_23726,N_22842,N_22936);
xnor U23727 (N_23727,N_22628,N_22419);
xnor U23728 (N_23728,N_22825,N_22709);
nor U23729 (N_23729,N_22027,N_22665);
and U23730 (N_23730,N_22530,N_22486);
and U23731 (N_23731,N_22940,N_22120);
nor U23732 (N_23732,N_22954,N_22246);
nand U23733 (N_23733,N_22031,N_22068);
and U23734 (N_23734,N_22772,N_22062);
xnor U23735 (N_23735,N_22465,N_22064);
xor U23736 (N_23736,N_22473,N_22257);
nor U23737 (N_23737,N_22199,N_22961);
and U23738 (N_23738,N_22388,N_22536);
or U23739 (N_23739,N_22765,N_22378);
nand U23740 (N_23740,N_22900,N_22041);
or U23741 (N_23741,N_22966,N_22464);
nor U23742 (N_23742,N_22545,N_22666);
nor U23743 (N_23743,N_22217,N_22593);
nor U23744 (N_23744,N_22645,N_22609);
nand U23745 (N_23745,N_22107,N_22815);
nand U23746 (N_23746,N_22608,N_22191);
nor U23747 (N_23747,N_22497,N_22618);
nor U23748 (N_23748,N_22548,N_22375);
and U23749 (N_23749,N_22611,N_22175);
or U23750 (N_23750,N_22199,N_22978);
and U23751 (N_23751,N_22950,N_22079);
or U23752 (N_23752,N_22839,N_22214);
nand U23753 (N_23753,N_22290,N_22750);
and U23754 (N_23754,N_22127,N_22329);
and U23755 (N_23755,N_22162,N_22358);
nand U23756 (N_23756,N_22201,N_22959);
nand U23757 (N_23757,N_22711,N_22846);
or U23758 (N_23758,N_22625,N_22710);
xor U23759 (N_23759,N_22133,N_22145);
nor U23760 (N_23760,N_22536,N_22906);
xnor U23761 (N_23761,N_22323,N_22105);
nand U23762 (N_23762,N_22811,N_22603);
or U23763 (N_23763,N_22421,N_22160);
or U23764 (N_23764,N_22898,N_22444);
nand U23765 (N_23765,N_22386,N_22873);
or U23766 (N_23766,N_22644,N_22474);
nor U23767 (N_23767,N_22420,N_22294);
xor U23768 (N_23768,N_22667,N_22323);
or U23769 (N_23769,N_22266,N_22168);
nor U23770 (N_23770,N_22071,N_22151);
xor U23771 (N_23771,N_22852,N_22981);
xor U23772 (N_23772,N_22560,N_22741);
xnor U23773 (N_23773,N_22702,N_22071);
nor U23774 (N_23774,N_22902,N_22174);
xor U23775 (N_23775,N_22437,N_22641);
nand U23776 (N_23776,N_22654,N_22238);
nor U23777 (N_23777,N_22299,N_22504);
nand U23778 (N_23778,N_22995,N_22228);
nand U23779 (N_23779,N_22008,N_22370);
or U23780 (N_23780,N_22905,N_22151);
nor U23781 (N_23781,N_22393,N_22759);
nor U23782 (N_23782,N_22495,N_22868);
xor U23783 (N_23783,N_22481,N_22879);
or U23784 (N_23784,N_22982,N_22726);
or U23785 (N_23785,N_22168,N_22237);
nand U23786 (N_23786,N_22063,N_22376);
nand U23787 (N_23787,N_22306,N_22585);
nand U23788 (N_23788,N_22191,N_22410);
and U23789 (N_23789,N_22387,N_22491);
nor U23790 (N_23790,N_22828,N_22012);
or U23791 (N_23791,N_22906,N_22292);
xor U23792 (N_23792,N_22850,N_22108);
nor U23793 (N_23793,N_22699,N_22608);
and U23794 (N_23794,N_22944,N_22004);
nor U23795 (N_23795,N_22219,N_22102);
xnor U23796 (N_23796,N_22120,N_22515);
or U23797 (N_23797,N_22471,N_22854);
nor U23798 (N_23798,N_22704,N_22771);
and U23799 (N_23799,N_22570,N_22037);
nor U23800 (N_23800,N_22060,N_22028);
xnor U23801 (N_23801,N_22470,N_22682);
xor U23802 (N_23802,N_22631,N_22072);
xor U23803 (N_23803,N_22012,N_22961);
nor U23804 (N_23804,N_22024,N_22774);
nor U23805 (N_23805,N_22571,N_22456);
and U23806 (N_23806,N_22313,N_22322);
nor U23807 (N_23807,N_22520,N_22644);
or U23808 (N_23808,N_22425,N_22433);
xnor U23809 (N_23809,N_22420,N_22902);
nand U23810 (N_23810,N_22819,N_22124);
nand U23811 (N_23811,N_22582,N_22304);
and U23812 (N_23812,N_22800,N_22158);
or U23813 (N_23813,N_22255,N_22918);
xnor U23814 (N_23814,N_22248,N_22408);
xnor U23815 (N_23815,N_22491,N_22959);
xor U23816 (N_23816,N_22836,N_22609);
xor U23817 (N_23817,N_22791,N_22906);
and U23818 (N_23818,N_22796,N_22860);
xnor U23819 (N_23819,N_22729,N_22956);
nand U23820 (N_23820,N_22029,N_22969);
and U23821 (N_23821,N_22282,N_22054);
nor U23822 (N_23822,N_22939,N_22407);
and U23823 (N_23823,N_22572,N_22253);
or U23824 (N_23824,N_22936,N_22176);
nor U23825 (N_23825,N_22354,N_22635);
nor U23826 (N_23826,N_22154,N_22084);
xor U23827 (N_23827,N_22639,N_22158);
nand U23828 (N_23828,N_22890,N_22167);
or U23829 (N_23829,N_22394,N_22009);
xor U23830 (N_23830,N_22972,N_22459);
or U23831 (N_23831,N_22282,N_22482);
nand U23832 (N_23832,N_22300,N_22929);
nand U23833 (N_23833,N_22218,N_22920);
and U23834 (N_23834,N_22626,N_22662);
nand U23835 (N_23835,N_22746,N_22809);
and U23836 (N_23836,N_22872,N_22543);
nor U23837 (N_23837,N_22587,N_22708);
xor U23838 (N_23838,N_22281,N_22593);
nor U23839 (N_23839,N_22562,N_22866);
xor U23840 (N_23840,N_22432,N_22270);
nor U23841 (N_23841,N_22278,N_22095);
and U23842 (N_23842,N_22388,N_22561);
and U23843 (N_23843,N_22837,N_22081);
nor U23844 (N_23844,N_22394,N_22550);
nor U23845 (N_23845,N_22190,N_22244);
xor U23846 (N_23846,N_22156,N_22445);
and U23847 (N_23847,N_22852,N_22242);
nor U23848 (N_23848,N_22461,N_22376);
xor U23849 (N_23849,N_22945,N_22117);
or U23850 (N_23850,N_22648,N_22202);
nand U23851 (N_23851,N_22516,N_22219);
nor U23852 (N_23852,N_22032,N_22422);
xor U23853 (N_23853,N_22273,N_22797);
nand U23854 (N_23854,N_22599,N_22090);
and U23855 (N_23855,N_22517,N_22325);
xor U23856 (N_23856,N_22198,N_22674);
nor U23857 (N_23857,N_22544,N_22714);
and U23858 (N_23858,N_22600,N_22958);
nand U23859 (N_23859,N_22123,N_22028);
xor U23860 (N_23860,N_22613,N_22577);
and U23861 (N_23861,N_22203,N_22418);
nor U23862 (N_23862,N_22503,N_22713);
nand U23863 (N_23863,N_22855,N_22562);
or U23864 (N_23864,N_22192,N_22610);
nor U23865 (N_23865,N_22762,N_22719);
xnor U23866 (N_23866,N_22912,N_22270);
xor U23867 (N_23867,N_22214,N_22900);
and U23868 (N_23868,N_22745,N_22658);
nor U23869 (N_23869,N_22052,N_22114);
nor U23870 (N_23870,N_22057,N_22898);
nand U23871 (N_23871,N_22800,N_22867);
nor U23872 (N_23872,N_22905,N_22420);
or U23873 (N_23873,N_22665,N_22225);
nand U23874 (N_23874,N_22831,N_22193);
or U23875 (N_23875,N_22128,N_22510);
or U23876 (N_23876,N_22416,N_22934);
nand U23877 (N_23877,N_22055,N_22789);
or U23878 (N_23878,N_22708,N_22614);
nand U23879 (N_23879,N_22692,N_22531);
xnor U23880 (N_23880,N_22301,N_22498);
xnor U23881 (N_23881,N_22087,N_22758);
or U23882 (N_23882,N_22991,N_22152);
or U23883 (N_23883,N_22466,N_22236);
nor U23884 (N_23884,N_22807,N_22940);
or U23885 (N_23885,N_22443,N_22981);
xnor U23886 (N_23886,N_22285,N_22349);
or U23887 (N_23887,N_22662,N_22964);
and U23888 (N_23888,N_22849,N_22161);
nand U23889 (N_23889,N_22907,N_22978);
and U23890 (N_23890,N_22214,N_22256);
nor U23891 (N_23891,N_22396,N_22077);
and U23892 (N_23892,N_22255,N_22830);
nor U23893 (N_23893,N_22233,N_22780);
and U23894 (N_23894,N_22809,N_22487);
and U23895 (N_23895,N_22556,N_22877);
nand U23896 (N_23896,N_22708,N_22792);
xor U23897 (N_23897,N_22228,N_22865);
xor U23898 (N_23898,N_22557,N_22109);
or U23899 (N_23899,N_22929,N_22147);
nand U23900 (N_23900,N_22169,N_22231);
xnor U23901 (N_23901,N_22434,N_22419);
nor U23902 (N_23902,N_22307,N_22622);
and U23903 (N_23903,N_22337,N_22487);
or U23904 (N_23904,N_22915,N_22705);
nor U23905 (N_23905,N_22719,N_22869);
nor U23906 (N_23906,N_22549,N_22225);
nand U23907 (N_23907,N_22817,N_22291);
and U23908 (N_23908,N_22734,N_22649);
xor U23909 (N_23909,N_22315,N_22130);
and U23910 (N_23910,N_22692,N_22005);
nand U23911 (N_23911,N_22921,N_22381);
and U23912 (N_23912,N_22931,N_22984);
nor U23913 (N_23913,N_22736,N_22680);
or U23914 (N_23914,N_22261,N_22827);
xnor U23915 (N_23915,N_22680,N_22365);
and U23916 (N_23916,N_22367,N_22148);
nor U23917 (N_23917,N_22447,N_22116);
nand U23918 (N_23918,N_22399,N_22287);
nand U23919 (N_23919,N_22036,N_22481);
nand U23920 (N_23920,N_22529,N_22864);
nand U23921 (N_23921,N_22124,N_22220);
nor U23922 (N_23922,N_22235,N_22920);
or U23923 (N_23923,N_22796,N_22043);
and U23924 (N_23924,N_22316,N_22615);
nor U23925 (N_23925,N_22888,N_22059);
nand U23926 (N_23926,N_22274,N_22017);
and U23927 (N_23927,N_22050,N_22028);
nand U23928 (N_23928,N_22185,N_22746);
nor U23929 (N_23929,N_22568,N_22769);
xnor U23930 (N_23930,N_22934,N_22500);
nor U23931 (N_23931,N_22679,N_22604);
nor U23932 (N_23932,N_22025,N_22457);
and U23933 (N_23933,N_22697,N_22344);
nand U23934 (N_23934,N_22428,N_22485);
and U23935 (N_23935,N_22432,N_22134);
nor U23936 (N_23936,N_22740,N_22904);
and U23937 (N_23937,N_22478,N_22230);
and U23938 (N_23938,N_22963,N_22240);
xor U23939 (N_23939,N_22636,N_22018);
nor U23940 (N_23940,N_22091,N_22291);
or U23941 (N_23941,N_22046,N_22829);
or U23942 (N_23942,N_22879,N_22290);
nor U23943 (N_23943,N_22118,N_22066);
or U23944 (N_23944,N_22579,N_22889);
nor U23945 (N_23945,N_22928,N_22528);
or U23946 (N_23946,N_22712,N_22990);
nand U23947 (N_23947,N_22944,N_22018);
or U23948 (N_23948,N_22864,N_22786);
and U23949 (N_23949,N_22406,N_22156);
xnor U23950 (N_23950,N_22276,N_22819);
nor U23951 (N_23951,N_22900,N_22501);
and U23952 (N_23952,N_22269,N_22281);
and U23953 (N_23953,N_22733,N_22680);
and U23954 (N_23954,N_22199,N_22233);
xor U23955 (N_23955,N_22667,N_22943);
nor U23956 (N_23956,N_22863,N_22315);
and U23957 (N_23957,N_22785,N_22366);
nand U23958 (N_23958,N_22120,N_22433);
xnor U23959 (N_23959,N_22349,N_22033);
nor U23960 (N_23960,N_22772,N_22934);
or U23961 (N_23961,N_22154,N_22161);
or U23962 (N_23962,N_22603,N_22533);
nor U23963 (N_23963,N_22947,N_22201);
nor U23964 (N_23964,N_22342,N_22982);
nand U23965 (N_23965,N_22902,N_22217);
or U23966 (N_23966,N_22714,N_22534);
nand U23967 (N_23967,N_22797,N_22063);
and U23968 (N_23968,N_22248,N_22292);
nand U23969 (N_23969,N_22943,N_22577);
nor U23970 (N_23970,N_22787,N_22146);
nand U23971 (N_23971,N_22868,N_22748);
nand U23972 (N_23972,N_22038,N_22105);
xor U23973 (N_23973,N_22256,N_22688);
and U23974 (N_23974,N_22841,N_22136);
nand U23975 (N_23975,N_22963,N_22229);
or U23976 (N_23976,N_22136,N_22116);
xor U23977 (N_23977,N_22294,N_22837);
or U23978 (N_23978,N_22228,N_22408);
xor U23979 (N_23979,N_22039,N_22613);
xnor U23980 (N_23980,N_22439,N_22899);
nor U23981 (N_23981,N_22765,N_22664);
or U23982 (N_23982,N_22377,N_22693);
and U23983 (N_23983,N_22358,N_22243);
nand U23984 (N_23984,N_22645,N_22722);
nand U23985 (N_23985,N_22523,N_22765);
xor U23986 (N_23986,N_22786,N_22716);
and U23987 (N_23987,N_22003,N_22235);
nor U23988 (N_23988,N_22890,N_22258);
and U23989 (N_23989,N_22430,N_22910);
and U23990 (N_23990,N_22213,N_22054);
xnor U23991 (N_23991,N_22147,N_22300);
xnor U23992 (N_23992,N_22662,N_22576);
or U23993 (N_23993,N_22708,N_22297);
xor U23994 (N_23994,N_22482,N_22619);
nor U23995 (N_23995,N_22256,N_22149);
xnor U23996 (N_23996,N_22591,N_22191);
and U23997 (N_23997,N_22329,N_22123);
nand U23998 (N_23998,N_22743,N_22791);
xnor U23999 (N_23999,N_22156,N_22964);
nand U24000 (N_24000,N_23323,N_23753);
nor U24001 (N_24001,N_23372,N_23455);
and U24002 (N_24002,N_23214,N_23571);
nor U24003 (N_24003,N_23120,N_23164);
xor U24004 (N_24004,N_23770,N_23781);
xor U24005 (N_24005,N_23004,N_23773);
and U24006 (N_24006,N_23168,N_23337);
xor U24007 (N_24007,N_23996,N_23142);
or U24008 (N_24008,N_23071,N_23900);
xnor U24009 (N_24009,N_23161,N_23495);
nor U24010 (N_24010,N_23944,N_23356);
or U24011 (N_24011,N_23492,N_23371);
nand U24012 (N_24012,N_23688,N_23799);
nand U24013 (N_24013,N_23267,N_23244);
and U24014 (N_24014,N_23025,N_23233);
xor U24015 (N_24015,N_23437,N_23442);
xor U24016 (N_24016,N_23384,N_23870);
nand U24017 (N_24017,N_23335,N_23529);
or U24018 (N_24018,N_23293,N_23227);
nand U24019 (N_24019,N_23292,N_23978);
nor U24020 (N_24020,N_23763,N_23821);
xor U24021 (N_24021,N_23157,N_23835);
xnor U24022 (N_24022,N_23787,N_23617);
nand U24023 (N_24023,N_23136,N_23092);
or U24024 (N_24024,N_23045,N_23199);
and U24025 (N_24025,N_23922,N_23370);
xnor U24026 (N_24026,N_23429,N_23677);
xor U24027 (N_24027,N_23351,N_23880);
xnor U24028 (N_24028,N_23287,N_23568);
and U24029 (N_24029,N_23731,N_23990);
or U24030 (N_24030,N_23908,N_23038);
nor U24031 (N_24031,N_23683,N_23423);
nor U24032 (N_24032,N_23203,N_23863);
and U24033 (N_24033,N_23628,N_23816);
xor U24034 (N_24034,N_23374,N_23473);
xor U24035 (N_24035,N_23091,N_23618);
nand U24036 (N_24036,N_23424,N_23848);
nor U24037 (N_24037,N_23265,N_23663);
xor U24038 (N_24038,N_23786,N_23151);
nor U24039 (N_24039,N_23130,N_23604);
or U24040 (N_24040,N_23512,N_23145);
nor U24041 (N_24041,N_23614,N_23684);
nor U24042 (N_24042,N_23928,N_23768);
xnor U24043 (N_24043,N_23884,N_23923);
and U24044 (N_24044,N_23599,N_23084);
and U24045 (N_24045,N_23710,N_23407);
and U24046 (N_24046,N_23002,N_23017);
and U24047 (N_24047,N_23317,N_23564);
and U24048 (N_24048,N_23232,N_23468);
or U24049 (N_24049,N_23822,N_23301);
or U24050 (N_24050,N_23426,N_23919);
or U24051 (N_24051,N_23373,N_23324);
xor U24052 (N_24052,N_23672,N_23970);
nand U24053 (N_24053,N_23388,N_23439);
nand U24054 (N_24054,N_23463,N_23026);
xor U24055 (N_24055,N_23148,N_23534);
nor U24056 (N_24056,N_23242,N_23619);
and U24057 (N_24057,N_23237,N_23976);
nand U24058 (N_24058,N_23701,N_23270);
nand U24059 (N_24059,N_23254,N_23703);
or U24060 (N_24060,N_23825,N_23462);
nand U24061 (N_24061,N_23447,N_23917);
nor U24062 (N_24062,N_23706,N_23275);
or U24063 (N_24063,N_23807,N_23221);
and U24064 (N_24064,N_23813,N_23645);
or U24065 (N_24065,N_23088,N_23031);
nand U24066 (N_24066,N_23850,N_23561);
xor U24067 (N_24067,N_23842,N_23048);
nor U24068 (N_24068,N_23115,N_23399);
xor U24069 (N_24069,N_23208,N_23500);
or U24070 (N_24070,N_23624,N_23118);
nor U24071 (N_24071,N_23566,N_23217);
xor U24072 (N_24072,N_23841,N_23650);
nand U24073 (N_24073,N_23176,N_23404);
or U24074 (N_24074,N_23887,N_23538);
or U24075 (N_24075,N_23975,N_23319);
nand U24076 (N_24076,N_23491,N_23847);
nor U24077 (N_24077,N_23304,N_23828);
and U24078 (N_24078,N_23470,N_23393);
xor U24079 (N_24079,N_23222,N_23851);
xor U24080 (N_24080,N_23702,N_23480);
xor U24081 (N_24081,N_23751,N_23644);
and U24082 (N_24082,N_23076,N_23300);
nor U24083 (N_24083,N_23250,N_23985);
nor U24084 (N_24084,N_23349,N_23111);
nand U24085 (N_24085,N_23581,N_23955);
xnor U24086 (N_24086,N_23195,N_23119);
xor U24087 (N_24087,N_23339,N_23152);
nand U24088 (N_24088,N_23137,N_23268);
nand U24089 (N_24089,N_23022,N_23478);
or U24090 (N_24090,N_23269,N_23635);
and U24091 (N_24091,N_23637,N_23907);
nor U24092 (N_24092,N_23752,N_23094);
nor U24093 (N_24093,N_23428,N_23431);
or U24094 (N_24094,N_23105,N_23519);
and U24095 (N_24095,N_23550,N_23971);
nand U24096 (N_24096,N_23836,N_23942);
nor U24097 (N_24097,N_23090,N_23732);
xnor U24098 (N_24098,N_23679,N_23612);
or U24099 (N_24099,N_23893,N_23106);
xor U24100 (N_24100,N_23032,N_23059);
or U24101 (N_24101,N_23591,N_23926);
nor U24102 (N_24102,N_23068,N_23359);
nand U24103 (N_24103,N_23814,N_23072);
or U24104 (N_24104,N_23569,N_23406);
nand U24105 (N_24105,N_23046,N_23416);
or U24106 (N_24106,N_23585,N_23818);
nor U24107 (N_24107,N_23494,N_23875);
or U24108 (N_24108,N_23030,N_23162);
xor U24109 (N_24109,N_23991,N_23108);
nand U24110 (N_24110,N_23365,N_23555);
nor U24111 (N_24111,N_23466,N_23170);
and U24112 (N_24112,N_23586,N_23865);
and U24113 (N_24113,N_23066,N_23750);
or U24114 (N_24114,N_23128,N_23541);
nand U24115 (N_24115,N_23338,N_23789);
nand U24116 (N_24116,N_23409,N_23489);
or U24117 (N_24117,N_23280,N_23283);
and U24118 (N_24118,N_23129,N_23475);
xor U24119 (N_24119,N_23326,N_23100);
nor U24120 (N_24120,N_23685,N_23943);
and U24121 (N_24121,N_23602,N_23929);
nand U24122 (N_24122,N_23224,N_23951);
nor U24123 (N_24123,N_23941,N_23657);
xor U24124 (N_24124,N_23749,N_23518);
or U24125 (N_24125,N_23008,N_23110);
or U24126 (N_24126,N_23190,N_23389);
and U24127 (N_24127,N_23024,N_23725);
nand U24128 (N_24128,N_23421,N_23109);
nand U24129 (N_24129,N_23296,N_23047);
and U24130 (N_24130,N_23903,N_23554);
or U24131 (N_24131,N_23631,N_23675);
or U24132 (N_24132,N_23665,N_23213);
or U24133 (N_24133,N_23918,N_23140);
nand U24134 (N_24134,N_23273,N_23352);
nor U24135 (N_24135,N_23589,N_23327);
and U24136 (N_24136,N_23403,N_23674);
nor U24137 (N_24137,N_23889,N_23775);
or U24138 (N_24138,N_23150,N_23952);
xor U24139 (N_24139,N_23185,N_23009);
nand U24140 (N_24140,N_23358,N_23112);
nand U24141 (N_24141,N_23769,N_23797);
xor U24142 (N_24142,N_23594,N_23994);
nand U24143 (N_24143,N_23459,N_23720);
xnor U24144 (N_24144,N_23973,N_23180);
or U24145 (N_24145,N_23476,N_23306);
and U24146 (N_24146,N_23791,N_23510);
nor U24147 (N_24147,N_23843,N_23745);
nand U24148 (N_24148,N_23123,N_23829);
nor U24149 (N_24149,N_23949,N_23827);
or U24150 (N_24150,N_23866,N_23549);
xor U24151 (N_24151,N_23877,N_23697);
and U24152 (N_24152,N_23515,N_23400);
nand U24153 (N_24153,N_23995,N_23694);
and U24154 (N_24154,N_23632,N_23098);
and U24155 (N_24155,N_23114,N_23307);
or U24156 (N_24156,N_23715,N_23433);
xor U24157 (N_24157,N_23014,N_23113);
and U24158 (N_24158,N_23499,N_23159);
and U24159 (N_24159,N_23837,N_23945);
xnor U24160 (N_24160,N_23346,N_23838);
xor U24161 (N_24161,N_23450,N_23989);
and U24162 (N_24162,N_23528,N_23933);
nor U24163 (N_24163,N_23334,N_23616);
nand U24164 (N_24164,N_23078,N_23754);
and U24165 (N_24165,N_23959,N_23210);
xnor U24166 (N_24166,N_23178,N_23065);
and U24167 (N_24167,N_23678,N_23039);
nand U24168 (N_24168,N_23761,N_23805);
xor U24169 (N_24169,N_23704,N_23759);
and U24170 (N_24170,N_23931,N_23241);
nand U24171 (N_24171,N_23856,N_23737);
nand U24172 (N_24172,N_23667,N_23689);
nand U24173 (N_24173,N_23264,N_23597);
nand U24174 (N_24174,N_23297,N_23007);
and U24175 (N_24175,N_23531,N_23392);
xor U24176 (N_24176,N_23206,N_23215);
nand U24177 (N_24177,N_23288,N_23023);
nor U24178 (N_24178,N_23496,N_23143);
or U24179 (N_24179,N_23800,N_23193);
and U24180 (N_24180,N_23207,N_23006);
or U24181 (N_24181,N_23498,N_23965);
or U24182 (N_24182,N_23879,N_23036);
nand U24183 (N_24183,N_23840,N_23124);
and U24184 (N_24184,N_23896,N_23713);
nor U24185 (N_24185,N_23557,N_23913);
xnor U24186 (N_24186,N_23417,N_23432);
and U24187 (N_24187,N_23669,N_23386);
xnor U24188 (N_24188,N_23643,N_23765);
xnor U24189 (N_24189,N_23303,N_23011);
or U24190 (N_24190,N_23547,N_23497);
xnor U24191 (N_24191,N_23321,N_23378);
xor U24192 (N_24192,N_23397,N_23792);
nor U24193 (N_24193,N_23460,N_23535);
and U24194 (N_24194,N_23956,N_23248);
and U24195 (N_24195,N_23967,N_23261);
and U24196 (N_24196,N_23696,N_23852);
xor U24197 (N_24197,N_23532,N_23166);
xor U24198 (N_24198,N_23660,N_23892);
nand U24199 (N_24199,N_23601,N_23874);
xor U24200 (N_24200,N_23488,N_23575);
or U24201 (N_24201,N_23298,N_23316);
and U24202 (N_24202,N_23544,N_23369);
nor U24203 (N_24203,N_23079,N_23172);
xor U24204 (N_24204,N_23379,N_23181);
nand U24205 (N_24205,N_23451,N_23043);
and U24206 (N_24206,N_23471,N_23686);
nand U24207 (N_24207,N_23340,N_23259);
xor U24208 (N_24208,N_23202,N_23121);
xnor U24209 (N_24209,N_23551,N_23153);
nor U24210 (N_24210,N_23226,N_23061);
nand U24211 (N_24211,N_23655,N_23003);
or U24212 (N_24212,N_23553,N_23739);
xor U24213 (N_24213,N_23653,N_23899);
xor U24214 (N_24214,N_23401,N_23681);
and U24215 (N_24215,N_23169,N_23398);
nand U24216 (N_24216,N_23735,N_23290);
nand U24217 (N_24217,N_23832,N_23289);
nor U24218 (N_24218,N_23698,N_23782);
and U24219 (N_24219,N_23073,N_23276);
xnor U24220 (N_24220,N_23383,N_23074);
or U24221 (N_24221,N_23435,N_23205);
or U24222 (N_24222,N_23320,N_23521);
or U24223 (N_24223,N_23311,N_23051);
nand U24224 (N_24224,N_23778,N_23760);
and U24225 (N_24225,N_23235,N_23132);
nand U24226 (N_24226,N_23651,N_23104);
or U24227 (N_24227,N_23156,N_23484);
and U24228 (N_24228,N_23993,N_23201);
or U24229 (N_24229,N_23277,N_23200);
nor U24230 (N_24230,N_23687,N_23060);
nand U24231 (N_24231,N_23709,N_23891);
nand U24232 (N_24232,N_23777,N_23033);
nand U24233 (N_24233,N_23620,N_23695);
xnor U24234 (N_24234,N_23138,N_23101);
nand U24235 (N_24235,N_23390,N_23723);
nand U24236 (N_24236,N_23229,N_23394);
or U24237 (N_24237,N_23804,N_23490);
nand U24238 (N_24238,N_23191,N_23331);
xnor U24239 (N_24239,N_23219,N_23794);
or U24240 (N_24240,N_23075,N_23888);
xor U24241 (N_24241,N_23000,N_23988);
xnor U24242 (N_24242,N_23155,N_23458);
and U24243 (N_24243,N_23504,N_23691);
xnor U24244 (N_24244,N_23741,N_23730);
nor U24245 (N_24245,N_23693,N_23443);
nor U24246 (N_24246,N_23050,N_23448);
nand U24247 (N_24247,N_23901,N_23165);
xor U24248 (N_24248,N_23175,N_23666);
nand U24249 (N_24249,N_23948,N_23251);
and U24250 (N_24250,N_23905,N_23436);
and U24251 (N_24251,N_23354,N_23318);
nor U24252 (N_24252,N_23826,N_23312);
nor U24253 (N_24253,N_23279,N_23328);
nand U24254 (N_24254,N_23188,N_23187);
xnor U24255 (N_24255,N_23097,N_23353);
nand U24256 (N_24256,N_23795,N_23493);
and U24257 (N_24257,N_23211,N_23154);
nand U24258 (N_24258,N_23367,N_23131);
nand U24259 (N_24259,N_23027,N_23615);
and U24260 (N_24260,N_23536,N_23779);
nand U24261 (N_24261,N_23692,N_23867);
nor U24262 (N_24262,N_23332,N_23295);
or U24263 (N_24263,N_23064,N_23081);
or U24264 (N_24264,N_23921,N_23964);
or U24265 (N_24265,N_23984,N_23158);
nor U24266 (N_24266,N_23871,N_23330);
xor U24267 (N_24267,N_23056,N_23972);
nand U24268 (N_24268,N_23182,N_23600);
nand U24269 (N_24269,N_23209,N_23830);
and U24270 (N_24270,N_23380,N_23664);
xor U24271 (N_24271,N_23579,N_23095);
or U24272 (N_24272,N_23603,N_23034);
or U24273 (N_24273,N_23231,N_23469);
xnor U24274 (N_24274,N_23438,N_23630);
nor U24275 (N_24275,N_23934,N_23873);
and U24276 (N_24276,N_23748,N_23413);
nor U24277 (N_24277,N_23937,N_23236);
nand U24278 (N_24278,N_23141,N_23461);
xnor U24279 (N_24279,N_23588,N_23507);
and U24280 (N_24280,N_23481,N_23015);
nand U24281 (N_24281,N_23345,N_23756);
nand U24282 (N_24282,N_23147,N_23486);
xor U24283 (N_24283,N_23058,N_23271);
or U24284 (N_24284,N_23590,N_23572);
xor U24285 (N_24285,N_23107,N_23482);
and U24286 (N_24286,N_23020,N_23418);
and U24287 (N_24287,N_23285,N_23508);
xnor U24288 (N_24288,N_23347,N_23982);
and U24289 (N_24289,N_23610,N_23505);
or U24290 (N_24290,N_23573,N_23652);
or U24291 (N_24291,N_23134,N_23662);
or U24292 (N_24292,N_23368,N_23823);
nand U24293 (N_24293,N_23998,N_23634);
and U24294 (N_24294,N_23649,N_23912);
nor U24295 (N_24295,N_23344,N_23796);
nor U24296 (N_24296,N_23744,N_23186);
xnor U24297 (N_24297,N_23171,N_23096);
and U24298 (N_24298,N_23381,N_23018);
or U24299 (N_24299,N_23846,N_23758);
nand U24300 (N_24300,N_23950,N_23981);
nor U24301 (N_24301,N_23824,N_23817);
or U24302 (N_24302,N_23196,N_23184);
xor U24303 (N_24303,N_23391,N_23514);
and U24304 (N_24304,N_23559,N_23733);
nand U24305 (N_24305,N_23523,N_23785);
nor U24306 (N_24306,N_23772,N_23886);
or U24307 (N_24307,N_23427,N_23253);
and U24308 (N_24308,N_23743,N_23342);
nor U24309 (N_24309,N_23894,N_23258);
and U24310 (N_24310,N_23979,N_23560);
xnor U24311 (N_24311,N_23216,N_23668);
nor U24312 (N_24312,N_23282,N_23053);
nand U24313 (N_24313,N_23454,N_23013);
and U24314 (N_24314,N_23305,N_23960);
and U24315 (N_24315,N_23444,N_23537);
or U24316 (N_24316,N_23883,N_23966);
and U24317 (N_24317,N_23054,N_23361);
or U24318 (N_24318,N_23576,N_23935);
xnor U24319 (N_24319,N_23636,N_23953);
xor U24320 (N_24320,N_23815,N_23712);
or U24321 (N_24321,N_23160,N_23986);
or U24322 (N_24322,N_23661,N_23911);
nor U24323 (N_24323,N_23801,N_23308);
nor U24324 (N_24324,N_23527,N_23286);
xnor U24325 (N_24325,N_23646,N_23876);
xnor U24326 (N_24326,N_23658,N_23626);
nand U24327 (N_24327,N_23783,N_23997);
or U24328 (N_24328,N_23596,N_23049);
nor U24329 (N_24329,N_23452,N_23167);
nor U24330 (N_24330,N_23525,N_23906);
or U24331 (N_24331,N_23810,N_23310);
nor U24332 (N_24332,N_23360,N_23629);
and U24333 (N_24333,N_23117,N_23639);
nor U24334 (N_24334,N_23093,N_23410);
nor U24335 (N_24335,N_23563,N_23577);
xnor U24336 (N_24336,N_23387,N_23910);
xnor U24337 (N_24337,N_23329,N_23595);
xor U24338 (N_24338,N_23592,N_23747);
and U24339 (N_24339,N_23272,N_23915);
or U24340 (N_24340,N_23256,N_23021);
nand U24341 (N_24341,N_23080,N_23502);
nor U24342 (N_24342,N_23414,N_23240);
nor U24343 (N_24343,N_23540,N_23315);
xor U24344 (N_24344,N_23700,N_23764);
nand U24345 (N_24345,N_23927,N_23642);
or U24346 (N_24346,N_23611,N_23127);
and U24347 (N_24347,N_23052,N_23477);
xor U24348 (N_24348,N_23548,N_23247);
and U24349 (N_24349,N_23946,N_23808);
nor U24350 (N_24350,N_23234,N_23844);
xor U24351 (N_24351,N_23281,N_23890);
and U24352 (N_24352,N_23366,N_23987);
nand U24353 (N_24353,N_23774,N_23126);
nor U24354 (N_24354,N_23062,N_23453);
nand U24355 (N_24355,N_23262,N_23350);
nor U24356 (N_24356,N_23957,N_23278);
xor U24357 (N_24357,N_23472,N_23336);
nor U24358 (N_24358,N_23574,N_23930);
nand U24359 (N_24359,N_23809,N_23968);
or U24360 (N_24360,N_23983,N_23456);
or U24361 (N_24361,N_23717,N_23341);
nor U24362 (N_24362,N_23562,N_23087);
xor U24363 (N_24363,N_23567,N_23977);
and U24364 (N_24364,N_23333,N_23375);
nand U24365 (N_24365,N_23220,N_23430);
nand U24366 (N_24366,N_23582,N_23771);
and U24367 (N_24367,N_23654,N_23909);
and U24368 (N_24368,N_23063,N_23252);
and U24369 (N_24369,N_23294,N_23396);
and U24370 (N_24370,N_23086,N_23938);
nand U24371 (N_24371,N_23446,N_23633);
nor U24372 (N_24372,N_23445,N_23419);
and U24373 (N_24373,N_23144,N_23299);
nand U24374 (N_24374,N_23864,N_23882);
nand U24375 (N_24375,N_23057,N_23405);
and U24376 (N_24376,N_23793,N_23627);
nor U24377 (N_24377,N_23881,N_23558);
nand U24378 (N_24378,N_23606,N_23385);
nor U24379 (N_24379,N_23859,N_23501);
and U24380 (N_24380,N_23539,N_23831);
or U24381 (N_24381,N_23146,N_23246);
xor U24382 (N_24382,N_23895,N_23249);
nand U24383 (N_24383,N_23855,N_23609);
and U24384 (N_24384,N_23016,N_23040);
or U24385 (N_24385,N_23309,N_23395);
nor U24386 (N_24386,N_23578,N_23511);
and U24387 (N_24387,N_23920,N_23343);
and U24388 (N_24388,N_23716,N_23640);
nand U24389 (N_24389,N_23357,N_23099);
nor U24390 (N_24390,N_23449,N_23412);
nand U24391 (N_24391,N_23364,N_23382);
or U24392 (N_24392,N_23806,N_23077);
nor U24393 (N_24393,N_23740,N_23082);
nand U24394 (N_24394,N_23992,N_23411);
xor U24395 (N_24395,N_23868,N_23055);
nor U24396 (N_24396,N_23070,N_23718);
and U24397 (N_24397,N_23485,N_23212);
nand U24398 (N_24398,N_23570,N_23999);
and U24399 (N_24399,N_23853,N_23820);
nand U24400 (N_24400,N_23916,N_23238);
nand U24401 (N_24401,N_23291,N_23483);
and U24402 (N_24402,N_23862,N_23322);
or U24403 (N_24403,N_23947,N_23355);
xnor U24404 (N_24404,N_23656,N_23543);
nand U24405 (N_24405,N_23858,N_23707);
and U24406 (N_24406,N_23545,N_23001);
nor U24407 (N_24407,N_23197,N_23961);
nor U24408 (N_24408,N_23263,N_23598);
xnor U24409 (N_24409,N_23724,N_23625);
nand U24410 (N_24410,N_23776,N_23010);
or U24411 (N_24411,N_23425,N_23362);
nand U24412 (N_24412,N_23122,N_23194);
nor U24413 (N_24413,N_23402,N_23727);
and U24414 (N_24414,N_23530,N_23708);
nand U24415 (N_24415,N_23699,N_23513);
and U24416 (N_24416,N_23936,N_23464);
or U24417 (N_24417,N_23533,N_23638);
nor U24418 (N_24418,N_23622,N_23089);
and U24419 (N_24419,N_23742,N_23019);
or U24420 (N_24420,N_23608,N_23245);
nor U24421 (N_24421,N_23924,N_23854);
nor U24422 (N_24422,N_23621,N_23734);
nor U24423 (N_24423,N_23974,N_23587);
xor U24424 (N_24424,N_23802,N_23125);
or U24425 (N_24425,N_23467,N_23849);
and U24426 (N_24426,N_23257,N_23902);
xnor U24427 (N_24427,N_23542,N_23798);
nand U24428 (N_24428,N_23962,N_23705);
and U24429 (N_24429,N_23659,N_23012);
nand U24430 (N_24430,N_23204,N_23861);
and U24431 (N_24431,N_23613,N_23812);
nand U24432 (N_24432,N_23474,N_23746);
xor U24433 (N_24433,N_23503,N_23834);
nand U24434 (N_24434,N_23174,N_23565);
nor U24435 (N_24435,N_23721,N_23682);
or U24436 (N_24436,N_23198,N_23552);
xnor U24437 (N_24437,N_23035,N_23860);
and U24438 (N_24438,N_23255,N_23584);
nor U24439 (N_24439,N_23083,N_23239);
or U24440 (N_24440,N_23963,N_23302);
or U24441 (N_24441,N_23230,N_23738);
and U24442 (N_24442,N_23788,N_23784);
xnor U24443 (N_24443,N_23583,N_23904);
xnor U24444 (N_24444,N_23487,N_23641);
nor U24445 (N_24445,N_23218,N_23872);
and U24446 (N_24446,N_23593,N_23363);
nand U24447 (N_24447,N_23671,N_23189);
or U24448 (N_24448,N_23376,N_23736);
nor U24449 (N_24449,N_23673,N_23029);
xnor U24450 (N_24450,N_23348,N_23192);
xnor U24451 (N_24451,N_23526,N_23037);
nand U24452 (N_24452,N_23897,N_23878);
nor U24453 (N_24453,N_23434,N_23811);
xor U24454 (N_24454,N_23103,N_23728);
nor U24455 (N_24455,N_23313,N_23914);
xnor U24456 (N_24456,N_23314,N_23516);
xor U24457 (N_24457,N_23260,N_23139);
nand U24458 (N_24458,N_23005,N_23648);
or U24459 (N_24459,N_23898,N_23819);
xor U24460 (N_24460,N_23790,N_23149);
nor U24461 (N_24461,N_23722,N_23266);
xnor U24462 (N_24462,N_23177,N_23607);
xor U24463 (N_24463,N_23958,N_23885);
or U24464 (N_24464,N_23225,N_23325);
nand U24465 (N_24465,N_23780,N_23408);
xnor U24466 (N_24466,N_23845,N_23670);
or U24467 (N_24467,N_23803,N_23932);
xnor U24468 (N_24468,N_23729,N_23546);
or U24469 (N_24469,N_23869,N_23605);
and U24470 (N_24470,N_23680,N_23274);
xor U24471 (N_24471,N_23767,N_23925);
xor U24472 (N_24472,N_23711,N_23517);
or U24473 (N_24473,N_23623,N_23228);
nand U24474 (N_24474,N_23441,N_23839);
nor U24475 (N_24475,N_23954,N_23415);
xor U24476 (N_24476,N_23719,N_23857);
nor U24477 (N_24477,N_23085,N_23243);
xnor U24478 (N_24478,N_23044,N_23457);
nor U24479 (N_24479,N_23556,N_23377);
nand U24480 (N_24480,N_23284,N_23479);
and U24481 (N_24481,N_23420,N_23173);
xnor U24482 (N_24482,N_23223,N_23755);
or U24483 (N_24483,N_23676,N_23939);
nor U24484 (N_24484,N_23440,N_23506);
or U24485 (N_24485,N_23179,N_23757);
nand U24486 (N_24486,N_23042,N_23647);
nand U24487 (N_24487,N_23102,N_23028);
and U24488 (N_24488,N_23133,N_23714);
nor U24489 (N_24489,N_23524,N_23422);
nand U24490 (N_24490,N_23163,N_23762);
and U24491 (N_24491,N_23940,N_23766);
and U24492 (N_24492,N_23465,N_23520);
or U24493 (N_24493,N_23980,N_23522);
nand U24494 (N_24494,N_23183,N_23580);
xor U24495 (N_24495,N_23067,N_23135);
or U24496 (N_24496,N_23833,N_23726);
nor U24497 (N_24497,N_23116,N_23041);
or U24498 (N_24498,N_23069,N_23969);
or U24499 (N_24499,N_23509,N_23690);
and U24500 (N_24500,N_23557,N_23213);
or U24501 (N_24501,N_23556,N_23601);
xnor U24502 (N_24502,N_23604,N_23992);
nand U24503 (N_24503,N_23282,N_23795);
nor U24504 (N_24504,N_23102,N_23011);
or U24505 (N_24505,N_23835,N_23038);
nand U24506 (N_24506,N_23607,N_23204);
nor U24507 (N_24507,N_23009,N_23657);
and U24508 (N_24508,N_23663,N_23248);
nor U24509 (N_24509,N_23756,N_23975);
or U24510 (N_24510,N_23627,N_23149);
nand U24511 (N_24511,N_23151,N_23703);
nor U24512 (N_24512,N_23194,N_23298);
and U24513 (N_24513,N_23377,N_23728);
xor U24514 (N_24514,N_23616,N_23537);
nand U24515 (N_24515,N_23041,N_23505);
xor U24516 (N_24516,N_23247,N_23251);
xor U24517 (N_24517,N_23927,N_23871);
nor U24518 (N_24518,N_23707,N_23552);
xnor U24519 (N_24519,N_23410,N_23203);
or U24520 (N_24520,N_23475,N_23041);
xnor U24521 (N_24521,N_23734,N_23989);
nand U24522 (N_24522,N_23413,N_23708);
nor U24523 (N_24523,N_23281,N_23762);
nor U24524 (N_24524,N_23802,N_23641);
or U24525 (N_24525,N_23065,N_23079);
nor U24526 (N_24526,N_23063,N_23675);
xnor U24527 (N_24527,N_23818,N_23702);
xor U24528 (N_24528,N_23161,N_23584);
and U24529 (N_24529,N_23330,N_23191);
nor U24530 (N_24530,N_23344,N_23231);
nor U24531 (N_24531,N_23449,N_23877);
xor U24532 (N_24532,N_23953,N_23759);
or U24533 (N_24533,N_23180,N_23054);
nor U24534 (N_24534,N_23200,N_23925);
and U24535 (N_24535,N_23970,N_23953);
and U24536 (N_24536,N_23647,N_23657);
and U24537 (N_24537,N_23519,N_23829);
nand U24538 (N_24538,N_23198,N_23805);
or U24539 (N_24539,N_23853,N_23464);
xnor U24540 (N_24540,N_23903,N_23018);
nand U24541 (N_24541,N_23095,N_23572);
nand U24542 (N_24542,N_23079,N_23342);
nor U24543 (N_24543,N_23033,N_23861);
nor U24544 (N_24544,N_23193,N_23151);
and U24545 (N_24545,N_23984,N_23579);
xnor U24546 (N_24546,N_23478,N_23789);
xnor U24547 (N_24547,N_23390,N_23777);
or U24548 (N_24548,N_23345,N_23786);
nand U24549 (N_24549,N_23684,N_23088);
nor U24550 (N_24550,N_23176,N_23670);
xor U24551 (N_24551,N_23853,N_23573);
and U24552 (N_24552,N_23885,N_23956);
or U24553 (N_24553,N_23689,N_23009);
nor U24554 (N_24554,N_23519,N_23093);
or U24555 (N_24555,N_23482,N_23671);
or U24556 (N_24556,N_23097,N_23792);
xnor U24557 (N_24557,N_23179,N_23816);
or U24558 (N_24558,N_23766,N_23176);
and U24559 (N_24559,N_23426,N_23111);
and U24560 (N_24560,N_23139,N_23622);
xnor U24561 (N_24561,N_23986,N_23047);
xor U24562 (N_24562,N_23909,N_23852);
and U24563 (N_24563,N_23336,N_23251);
and U24564 (N_24564,N_23892,N_23861);
xnor U24565 (N_24565,N_23013,N_23786);
nor U24566 (N_24566,N_23915,N_23860);
and U24567 (N_24567,N_23208,N_23254);
nand U24568 (N_24568,N_23700,N_23186);
nand U24569 (N_24569,N_23991,N_23123);
xor U24570 (N_24570,N_23988,N_23375);
nand U24571 (N_24571,N_23092,N_23268);
nor U24572 (N_24572,N_23051,N_23219);
and U24573 (N_24573,N_23136,N_23642);
xor U24574 (N_24574,N_23358,N_23164);
or U24575 (N_24575,N_23025,N_23502);
xnor U24576 (N_24576,N_23266,N_23455);
xor U24577 (N_24577,N_23111,N_23365);
nand U24578 (N_24578,N_23791,N_23888);
nand U24579 (N_24579,N_23107,N_23487);
or U24580 (N_24580,N_23257,N_23935);
or U24581 (N_24581,N_23334,N_23454);
xnor U24582 (N_24582,N_23842,N_23986);
nor U24583 (N_24583,N_23650,N_23621);
xnor U24584 (N_24584,N_23880,N_23391);
xnor U24585 (N_24585,N_23500,N_23345);
xnor U24586 (N_24586,N_23539,N_23153);
and U24587 (N_24587,N_23715,N_23596);
nor U24588 (N_24588,N_23926,N_23597);
and U24589 (N_24589,N_23181,N_23530);
xnor U24590 (N_24590,N_23446,N_23124);
nand U24591 (N_24591,N_23811,N_23306);
xor U24592 (N_24592,N_23732,N_23967);
nor U24593 (N_24593,N_23063,N_23439);
or U24594 (N_24594,N_23671,N_23751);
nand U24595 (N_24595,N_23117,N_23603);
nand U24596 (N_24596,N_23385,N_23526);
nor U24597 (N_24597,N_23959,N_23991);
nor U24598 (N_24598,N_23587,N_23153);
xor U24599 (N_24599,N_23887,N_23945);
xor U24600 (N_24600,N_23311,N_23751);
xor U24601 (N_24601,N_23663,N_23925);
and U24602 (N_24602,N_23612,N_23080);
nor U24603 (N_24603,N_23313,N_23234);
nand U24604 (N_24604,N_23909,N_23931);
nand U24605 (N_24605,N_23674,N_23923);
xnor U24606 (N_24606,N_23643,N_23373);
nand U24607 (N_24607,N_23966,N_23001);
xnor U24608 (N_24608,N_23373,N_23941);
xnor U24609 (N_24609,N_23553,N_23078);
or U24610 (N_24610,N_23365,N_23979);
nand U24611 (N_24611,N_23116,N_23142);
and U24612 (N_24612,N_23982,N_23801);
nand U24613 (N_24613,N_23149,N_23226);
xnor U24614 (N_24614,N_23307,N_23264);
nand U24615 (N_24615,N_23582,N_23335);
xor U24616 (N_24616,N_23329,N_23255);
or U24617 (N_24617,N_23419,N_23441);
xnor U24618 (N_24618,N_23093,N_23556);
nand U24619 (N_24619,N_23239,N_23413);
xor U24620 (N_24620,N_23403,N_23054);
or U24621 (N_24621,N_23956,N_23024);
and U24622 (N_24622,N_23695,N_23113);
or U24623 (N_24623,N_23325,N_23036);
nor U24624 (N_24624,N_23363,N_23159);
or U24625 (N_24625,N_23273,N_23741);
nor U24626 (N_24626,N_23744,N_23266);
xor U24627 (N_24627,N_23834,N_23320);
nor U24628 (N_24628,N_23743,N_23421);
and U24629 (N_24629,N_23188,N_23805);
nor U24630 (N_24630,N_23934,N_23790);
nor U24631 (N_24631,N_23006,N_23915);
nor U24632 (N_24632,N_23000,N_23214);
or U24633 (N_24633,N_23632,N_23974);
nand U24634 (N_24634,N_23051,N_23506);
nor U24635 (N_24635,N_23134,N_23195);
or U24636 (N_24636,N_23840,N_23497);
or U24637 (N_24637,N_23145,N_23505);
xnor U24638 (N_24638,N_23222,N_23035);
and U24639 (N_24639,N_23230,N_23024);
and U24640 (N_24640,N_23686,N_23091);
xnor U24641 (N_24641,N_23482,N_23286);
nor U24642 (N_24642,N_23263,N_23721);
nor U24643 (N_24643,N_23025,N_23967);
nand U24644 (N_24644,N_23456,N_23903);
and U24645 (N_24645,N_23630,N_23144);
and U24646 (N_24646,N_23445,N_23728);
xnor U24647 (N_24647,N_23461,N_23865);
and U24648 (N_24648,N_23708,N_23511);
xnor U24649 (N_24649,N_23951,N_23206);
or U24650 (N_24650,N_23767,N_23219);
nor U24651 (N_24651,N_23391,N_23465);
nand U24652 (N_24652,N_23068,N_23674);
and U24653 (N_24653,N_23155,N_23726);
nor U24654 (N_24654,N_23226,N_23831);
or U24655 (N_24655,N_23299,N_23347);
or U24656 (N_24656,N_23975,N_23760);
xor U24657 (N_24657,N_23916,N_23851);
nor U24658 (N_24658,N_23832,N_23013);
nor U24659 (N_24659,N_23021,N_23539);
nor U24660 (N_24660,N_23089,N_23727);
xor U24661 (N_24661,N_23035,N_23849);
and U24662 (N_24662,N_23181,N_23187);
xor U24663 (N_24663,N_23465,N_23583);
and U24664 (N_24664,N_23332,N_23821);
and U24665 (N_24665,N_23746,N_23840);
or U24666 (N_24666,N_23580,N_23641);
and U24667 (N_24667,N_23489,N_23984);
xor U24668 (N_24668,N_23862,N_23605);
nand U24669 (N_24669,N_23789,N_23254);
and U24670 (N_24670,N_23881,N_23851);
nand U24671 (N_24671,N_23158,N_23370);
nor U24672 (N_24672,N_23010,N_23850);
nor U24673 (N_24673,N_23057,N_23327);
nand U24674 (N_24674,N_23256,N_23839);
nand U24675 (N_24675,N_23067,N_23012);
nand U24676 (N_24676,N_23218,N_23065);
or U24677 (N_24677,N_23178,N_23545);
and U24678 (N_24678,N_23281,N_23291);
and U24679 (N_24679,N_23030,N_23118);
nor U24680 (N_24680,N_23749,N_23651);
nand U24681 (N_24681,N_23764,N_23734);
xor U24682 (N_24682,N_23937,N_23652);
nor U24683 (N_24683,N_23110,N_23866);
and U24684 (N_24684,N_23091,N_23728);
nand U24685 (N_24685,N_23364,N_23673);
nor U24686 (N_24686,N_23559,N_23862);
nor U24687 (N_24687,N_23913,N_23985);
xor U24688 (N_24688,N_23451,N_23872);
nand U24689 (N_24689,N_23894,N_23297);
xor U24690 (N_24690,N_23981,N_23347);
or U24691 (N_24691,N_23675,N_23746);
nand U24692 (N_24692,N_23682,N_23336);
or U24693 (N_24693,N_23805,N_23002);
or U24694 (N_24694,N_23861,N_23148);
and U24695 (N_24695,N_23754,N_23552);
nand U24696 (N_24696,N_23247,N_23560);
and U24697 (N_24697,N_23989,N_23687);
nand U24698 (N_24698,N_23205,N_23905);
or U24699 (N_24699,N_23861,N_23909);
or U24700 (N_24700,N_23547,N_23863);
or U24701 (N_24701,N_23253,N_23251);
and U24702 (N_24702,N_23330,N_23651);
or U24703 (N_24703,N_23935,N_23177);
nand U24704 (N_24704,N_23898,N_23980);
nor U24705 (N_24705,N_23620,N_23014);
nand U24706 (N_24706,N_23342,N_23622);
or U24707 (N_24707,N_23196,N_23821);
xor U24708 (N_24708,N_23655,N_23891);
nand U24709 (N_24709,N_23897,N_23640);
nor U24710 (N_24710,N_23093,N_23499);
and U24711 (N_24711,N_23728,N_23312);
or U24712 (N_24712,N_23491,N_23805);
or U24713 (N_24713,N_23447,N_23596);
or U24714 (N_24714,N_23146,N_23539);
xnor U24715 (N_24715,N_23792,N_23379);
xnor U24716 (N_24716,N_23374,N_23821);
xor U24717 (N_24717,N_23367,N_23789);
or U24718 (N_24718,N_23846,N_23470);
nand U24719 (N_24719,N_23218,N_23605);
nor U24720 (N_24720,N_23568,N_23483);
or U24721 (N_24721,N_23742,N_23018);
or U24722 (N_24722,N_23848,N_23820);
xnor U24723 (N_24723,N_23032,N_23298);
xnor U24724 (N_24724,N_23146,N_23989);
or U24725 (N_24725,N_23359,N_23888);
and U24726 (N_24726,N_23601,N_23824);
nand U24727 (N_24727,N_23956,N_23878);
or U24728 (N_24728,N_23701,N_23844);
and U24729 (N_24729,N_23555,N_23493);
nand U24730 (N_24730,N_23338,N_23955);
and U24731 (N_24731,N_23422,N_23268);
or U24732 (N_24732,N_23425,N_23746);
and U24733 (N_24733,N_23847,N_23985);
and U24734 (N_24734,N_23016,N_23960);
and U24735 (N_24735,N_23640,N_23279);
xnor U24736 (N_24736,N_23015,N_23679);
xnor U24737 (N_24737,N_23941,N_23033);
and U24738 (N_24738,N_23704,N_23644);
nand U24739 (N_24739,N_23367,N_23499);
or U24740 (N_24740,N_23124,N_23021);
or U24741 (N_24741,N_23912,N_23599);
xor U24742 (N_24742,N_23215,N_23372);
or U24743 (N_24743,N_23791,N_23294);
xnor U24744 (N_24744,N_23267,N_23879);
and U24745 (N_24745,N_23439,N_23115);
xor U24746 (N_24746,N_23331,N_23218);
or U24747 (N_24747,N_23944,N_23417);
xor U24748 (N_24748,N_23233,N_23406);
nand U24749 (N_24749,N_23226,N_23394);
xnor U24750 (N_24750,N_23285,N_23359);
nor U24751 (N_24751,N_23738,N_23871);
nand U24752 (N_24752,N_23160,N_23987);
nor U24753 (N_24753,N_23905,N_23906);
xor U24754 (N_24754,N_23498,N_23859);
and U24755 (N_24755,N_23590,N_23724);
nand U24756 (N_24756,N_23245,N_23629);
xnor U24757 (N_24757,N_23966,N_23101);
nand U24758 (N_24758,N_23024,N_23158);
and U24759 (N_24759,N_23420,N_23765);
xor U24760 (N_24760,N_23454,N_23603);
nor U24761 (N_24761,N_23049,N_23668);
and U24762 (N_24762,N_23997,N_23038);
and U24763 (N_24763,N_23362,N_23771);
xnor U24764 (N_24764,N_23899,N_23703);
or U24765 (N_24765,N_23873,N_23421);
or U24766 (N_24766,N_23165,N_23652);
nor U24767 (N_24767,N_23191,N_23717);
nor U24768 (N_24768,N_23605,N_23846);
nor U24769 (N_24769,N_23070,N_23314);
nand U24770 (N_24770,N_23422,N_23312);
xnor U24771 (N_24771,N_23332,N_23662);
and U24772 (N_24772,N_23971,N_23551);
xnor U24773 (N_24773,N_23710,N_23453);
nor U24774 (N_24774,N_23704,N_23426);
nand U24775 (N_24775,N_23003,N_23957);
or U24776 (N_24776,N_23886,N_23133);
and U24777 (N_24777,N_23523,N_23718);
xnor U24778 (N_24778,N_23492,N_23356);
or U24779 (N_24779,N_23750,N_23712);
xor U24780 (N_24780,N_23361,N_23206);
nor U24781 (N_24781,N_23616,N_23696);
and U24782 (N_24782,N_23891,N_23790);
nor U24783 (N_24783,N_23207,N_23507);
nor U24784 (N_24784,N_23642,N_23540);
nand U24785 (N_24785,N_23456,N_23025);
and U24786 (N_24786,N_23410,N_23023);
or U24787 (N_24787,N_23485,N_23831);
xnor U24788 (N_24788,N_23785,N_23266);
or U24789 (N_24789,N_23872,N_23610);
nand U24790 (N_24790,N_23271,N_23446);
xor U24791 (N_24791,N_23070,N_23836);
xnor U24792 (N_24792,N_23686,N_23271);
nor U24793 (N_24793,N_23257,N_23303);
nand U24794 (N_24794,N_23588,N_23258);
xor U24795 (N_24795,N_23482,N_23906);
nor U24796 (N_24796,N_23737,N_23172);
nand U24797 (N_24797,N_23526,N_23118);
nor U24798 (N_24798,N_23200,N_23301);
or U24799 (N_24799,N_23500,N_23742);
nand U24800 (N_24800,N_23098,N_23479);
nor U24801 (N_24801,N_23383,N_23501);
nand U24802 (N_24802,N_23810,N_23806);
xor U24803 (N_24803,N_23582,N_23579);
or U24804 (N_24804,N_23695,N_23400);
and U24805 (N_24805,N_23401,N_23341);
nand U24806 (N_24806,N_23562,N_23334);
nor U24807 (N_24807,N_23802,N_23859);
and U24808 (N_24808,N_23350,N_23224);
nor U24809 (N_24809,N_23191,N_23593);
xnor U24810 (N_24810,N_23198,N_23978);
nor U24811 (N_24811,N_23382,N_23089);
nor U24812 (N_24812,N_23409,N_23567);
or U24813 (N_24813,N_23911,N_23195);
or U24814 (N_24814,N_23151,N_23960);
xnor U24815 (N_24815,N_23067,N_23122);
or U24816 (N_24816,N_23503,N_23458);
nand U24817 (N_24817,N_23770,N_23500);
or U24818 (N_24818,N_23919,N_23018);
nor U24819 (N_24819,N_23676,N_23259);
or U24820 (N_24820,N_23945,N_23415);
xor U24821 (N_24821,N_23463,N_23212);
nand U24822 (N_24822,N_23692,N_23324);
or U24823 (N_24823,N_23490,N_23988);
nand U24824 (N_24824,N_23767,N_23721);
nor U24825 (N_24825,N_23018,N_23516);
nor U24826 (N_24826,N_23952,N_23100);
or U24827 (N_24827,N_23116,N_23567);
nand U24828 (N_24828,N_23466,N_23312);
xnor U24829 (N_24829,N_23425,N_23436);
nand U24830 (N_24830,N_23883,N_23732);
and U24831 (N_24831,N_23336,N_23834);
nand U24832 (N_24832,N_23824,N_23446);
nand U24833 (N_24833,N_23179,N_23045);
and U24834 (N_24834,N_23595,N_23438);
nor U24835 (N_24835,N_23675,N_23917);
or U24836 (N_24836,N_23926,N_23855);
nor U24837 (N_24837,N_23506,N_23048);
nand U24838 (N_24838,N_23310,N_23667);
nor U24839 (N_24839,N_23957,N_23475);
nor U24840 (N_24840,N_23476,N_23905);
and U24841 (N_24841,N_23608,N_23773);
nor U24842 (N_24842,N_23768,N_23314);
and U24843 (N_24843,N_23274,N_23068);
nand U24844 (N_24844,N_23715,N_23360);
xor U24845 (N_24845,N_23884,N_23396);
or U24846 (N_24846,N_23395,N_23136);
xor U24847 (N_24847,N_23630,N_23046);
nand U24848 (N_24848,N_23095,N_23553);
nor U24849 (N_24849,N_23856,N_23708);
nor U24850 (N_24850,N_23320,N_23757);
or U24851 (N_24851,N_23897,N_23099);
xnor U24852 (N_24852,N_23574,N_23554);
or U24853 (N_24853,N_23617,N_23665);
and U24854 (N_24854,N_23223,N_23298);
or U24855 (N_24855,N_23917,N_23358);
nand U24856 (N_24856,N_23904,N_23903);
nor U24857 (N_24857,N_23471,N_23387);
nand U24858 (N_24858,N_23380,N_23909);
and U24859 (N_24859,N_23966,N_23306);
and U24860 (N_24860,N_23777,N_23116);
and U24861 (N_24861,N_23858,N_23171);
nand U24862 (N_24862,N_23332,N_23183);
xor U24863 (N_24863,N_23876,N_23229);
xor U24864 (N_24864,N_23234,N_23500);
or U24865 (N_24865,N_23014,N_23341);
xnor U24866 (N_24866,N_23253,N_23079);
or U24867 (N_24867,N_23749,N_23102);
xor U24868 (N_24868,N_23741,N_23185);
xnor U24869 (N_24869,N_23845,N_23561);
and U24870 (N_24870,N_23022,N_23076);
xnor U24871 (N_24871,N_23789,N_23935);
or U24872 (N_24872,N_23729,N_23785);
nor U24873 (N_24873,N_23911,N_23380);
or U24874 (N_24874,N_23643,N_23898);
or U24875 (N_24875,N_23628,N_23423);
nor U24876 (N_24876,N_23771,N_23316);
nor U24877 (N_24877,N_23058,N_23758);
xnor U24878 (N_24878,N_23588,N_23956);
nand U24879 (N_24879,N_23092,N_23467);
or U24880 (N_24880,N_23409,N_23180);
nand U24881 (N_24881,N_23995,N_23222);
nor U24882 (N_24882,N_23183,N_23966);
xnor U24883 (N_24883,N_23672,N_23076);
xor U24884 (N_24884,N_23797,N_23807);
and U24885 (N_24885,N_23901,N_23334);
and U24886 (N_24886,N_23120,N_23726);
nor U24887 (N_24887,N_23535,N_23894);
nor U24888 (N_24888,N_23406,N_23391);
and U24889 (N_24889,N_23481,N_23271);
and U24890 (N_24890,N_23826,N_23369);
nand U24891 (N_24891,N_23389,N_23322);
and U24892 (N_24892,N_23136,N_23628);
and U24893 (N_24893,N_23546,N_23538);
nand U24894 (N_24894,N_23894,N_23027);
nor U24895 (N_24895,N_23566,N_23798);
nor U24896 (N_24896,N_23027,N_23188);
xor U24897 (N_24897,N_23350,N_23691);
or U24898 (N_24898,N_23413,N_23604);
or U24899 (N_24899,N_23726,N_23012);
or U24900 (N_24900,N_23149,N_23615);
or U24901 (N_24901,N_23066,N_23129);
nor U24902 (N_24902,N_23754,N_23521);
and U24903 (N_24903,N_23301,N_23175);
and U24904 (N_24904,N_23288,N_23615);
and U24905 (N_24905,N_23131,N_23727);
or U24906 (N_24906,N_23962,N_23136);
and U24907 (N_24907,N_23348,N_23267);
nand U24908 (N_24908,N_23830,N_23248);
xor U24909 (N_24909,N_23345,N_23109);
or U24910 (N_24910,N_23453,N_23945);
or U24911 (N_24911,N_23929,N_23205);
nand U24912 (N_24912,N_23308,N_23451);
xnor U24913 (N_24913,N_23351,N_23265);
and U24914 (N_24914,N_23733,N_23859);
or U24915 (N_24915,N_23986,N_23154);
or U24916 (N_24916,N_23821,N_23781);
xor U24917 (N_24917,N_23773,N_23587);
or U24918 (N_24918,N_23877,N_23721);
nor U24919 (N_24919,N_23218,N_23910);
nand U24920 (N_24920,N_23884,N_23569);
xnor U24921 (N_24921,N_23008,N_23577);
xnor U24922 (N_24922,N_23861,N_23859);
nand U24923 (N_24923,N_23308,N_23494);
and U24924 (N_24924,N_23730,N_23058);
nand U24925 (N_24925,N_23820,N_23625);
nor U24926 (N_24926,N_23445,N_23695);
and U24927 (N_24927,N_23234,N_23648);
nand U24928 (N_24928,N_23975,N_23217);
nand U24929 (N_24929,N_23621,N_23416);
or U24930 (N_24930,N_23160,N_23884);
or U24931 (N_24931,N_23157,N_23999);
xnor U24932 (N_24932,N_23517,N_23130);
xor U24933 (N_24933,N_23905,N_23627);
and U24934 (N_24934,N_23258,N_23934);
nor U24935 (N_24935,N_23459,N_23277);
nor U24936 (N_24936,N_23002,N_23550);
or U24937 (N_24937,N_23061,N_23469);
nor U24938 (N_24938,N_23369,N_23020);
nor U24939 (N_24939,N_23748,N_23561);
and U24940 (N_24940,N_23668,N_23290);
and U24941 (N_24941,N_23625,N_23898);
xor U24942 (N_24942,N_23467,N_23473);
xnor U24943 (N_24943,N_23652,N_23952);
nand U24944 (N_24944,N_23568,N_23694);
or U24945 (N_24945,N_23883,N_23022);
xnor U24946 (N_24946,N_23248,N_23558);
nand U24947 (N_24947,N_23290,N_23530);
and U24948 (N_24948,N_23010,N_23303);
nand U24949 (N_24949,N_23523,N_23031);
or U24950 (N_24950,N_23103,N_23820);
xor U24951 (N_24951,N_23758,N_23316);
nor U24952 (N_24952,N_23127,N_23573);
nand U24953 (N_24953,N_23247,N_23465);
nand U24954 (N_24954,N_23386,N_23712);
xor U24955 (N_24955,N_23596,N_23942);
xnor U24956 (N_24956,N_23548,N_23447);
and U24957 (N_24957,N_23238,N_23009);
nand U24958 (N_24958,N_23271,N_23048);
or U24959 (N_24959,N_23316,N_23448);
nand U24960 (N_24960,N_23300,N_23356);
or U24961 (N_24961,N_23405,N_23579);
xnor U24962 (N_24962,N_23003,N_23862);
xor U24963 (N_24963,N_23678,N_23768);
or U24964 (N_24964,N_23784,N_23395);
or U24965 (N_24965,N_23883,N_23494);
nor U24966 (N_24966,N_23857,N_23642);
xnor U24967 (N_24967,N_23873,N_23103);
or U24968 (N_24968,N_23316,N_23546);
or U24969 (N_24969,N_23601,N_23690);
nand U24970 (N_24970,N_23516,N_23096);
nor U24971 (N_24971,N_23780,N_23475);
or U24972 (N_24972,N_23610,N_23217);
nand U24973 (N_24973,N_23141,N_23040);
nor U24974 (N_24974,N_23993,N_23655);
and U24975 (N_24975,N_23884,N_23982);
xnor U24976 (N_24976,N_23976,N_23023);
or U24977 (N_24977,N_23808,N_23257);
and U24978 (N_24978,N_23177,N_23443);
nor U24979 (N_24979,N_23381,N_23114);
or U24980 (N_24980,N_23304,N_23104);
or U24981 (N_24981,N_23502,N_23039);
xor U24982 (N_24982,N_23096,N_23002);
and U24983 (N_24983,N_23688,N_23989);
nand U24984 (N_24984,N_23139,N_23501);
nor U24985 (N_24985,N_23357,N_23782);
and U24986 (N_24986,N_23985,N_23277);
nand U24987 (N_24987,N_23942,N_23913);
and U24988 (N_24988,N_23647,N_23154);
and U24989 (N_24989,N_23394,N_23104);
nor U24990 (N_24990,N_23347,N_23205);
or U24991 (N_24991,N_23689,N_23320);
nor U24992 (N_24992,N_23604,N_23572);
xnor U24993 (N_24993,N_23964,N_23534);
xnor U24994 (N_24994,N_23729,N_23283);
or U24995 (N_24995,N_23248,N_23492);
and U24996 (N_24996,N_23645,N_23156);
nand U24997 (N_24997,N_23921,N_23724);
nand U24998 (N_24998,N_23220,N_23847);
or U24999 (N_24999,N_23695,N_23100);
nor UO_0 (O_0,N_24560,N_24825);
nor UO_1 (O_1,N_24058,N_24201);
and UO_2 (O_2,N_24281,N_24898);
xnor UO_3 (O_3,N_24154,N_24065);
or UO_4 (O_4,N_24419,N_24139);
nand UO_5 (O_5,N_24975,N_24771);
nand UO_6 (O_6,N_24259,N_24725);
or UO_7 (O_7,N_24330,N_24890);
and UO_8 (O_8,N_24857,N_24881);
or UO_9 (O_9,N_24450,N_24336);
or UO_10 (O_10,N_24569,N_24548);
and UO_11 (O_11,N_24213,N_24850);
and UO_12 (O_12,N_24389,N_24808);
xnor UO_13 (O_13,N_24662,N_24634);
nand UO_14 (O_14,N_24282,N_24769);
nand UO_15 (O_15,N_24035,N_24004);
xnor UO_16 (O_16,N_24918,N_24737);
nand UO_17 (O_17,N_24360,N_24165);
and UO_18 (O_18,N_24566,N_24285);
xnor UO_19 (O_19,N_24145,N_24388);
nor UO_20 (O_20,N_24392,N_24511);
and UO_21 (O_21,N_24528,N_24742);
nor UO_22 (O_22,N_24985,N_24351);
nor UO_23 (O_23,N_24135,N_24254);
xor UO_24 (O_24,N_24971,N_24236);
nand UO_25 (O_25,N_24172,N_24822);
nand UO_26 (O_26,N_24289,N_24532);
nand UO_27 (O_27,N_24328,N_24224);
or UO_28 (O_28,N_24432,N_24972);
or UO_29 (O_29,N_24758,N_24365);
xor UO_30 (O_30,N_24160,N_24386);
or UO_31 (O_31,N_24544,N_24372);
or UO_32 (O_32,N_24200,N_24264);
xnor UO_33 (O_33,N_24955,N_24744);
nor UO_34 (O_34,N_24809,N_24494);
xnor UO_35 (O_35,N_24105,N_24377);
and UO_36 (O_36,N_24182,N_24605);
and UO_37 (O_37,N_24618,N_24128);
nor UO_38 (O_38,N_24446,N_24221);
and UO_39 (O_39,N_24789,N_24295);
and UO_40 (O_40,N_24038,N_24722);
nor UO_41 (O_41,N_24531,N_24510);
xor UO_42 (O_42,N_24483,N_24411);
nand UO_43 (O_43,N_24824,N_24148);
xnor UO_44 (O_44,N_24598,N_24417);
and UO_45 (O_45,N_24888,N_24288);
xor UO_46 (O_46,N_24197,N_24029);
or UO_47 (O_47,N_24640,N_24265);
and UO_48 (O_48,N_24358,N_24471);
nor UO_49 (O_49,N_24921,N_24706);
nand UO_50 (O_50,N_24556,N_24699);
or UO_51 (O_51,N_24923,N_24959);
nor UO_52 (O_52,N_24911,N_24858);
nand UO_53 (O_53,N_24420,N_24207);
and UO_54 (O_54,N_24387,N_24986);
or UO_55 (O_55,N_24130,N_24137);
and UO_56 (O_56,N_24472,N_24144);
and UO_57 (O_57,N_24287,N_24781);
nand UO_58 (O_58,N_24501,N_24623);
xnor UO_59 (O_59,N_24841,N_24908);
and UO_60 (O_60,N_24322,N_24700);
nor UO_61 (O_61,N_24210,N_24932);
xnor UO_62 (O_62,N_24622,N_24708);
xnor UO_63 (O_63,N_24924,N_24514);
nand UO_64 (O_64,N_24869,N_24083);
nor UO_65 (O_65,N_24845,N_24516);
xor UO_66 (O_66,N_24997,N_24752);
xor UO_67 (O_67,N_24587,N_24729);
xnor UO_68 (O_68,N_24895,N_24016);
or UO_69 (O_69,N_24939,N_24637);
nor UO_70 (O_70,N_24804,N_24376);
xor UO_71 (O_71,N_24206,N_24068);
nand UO_72 (O_72,N_24436,N_24831);
and UO_73 (O_73,N_24306,N_24175);
and UO_74 (O_74,N_24547,N_24082);
nand UO_75 (O_75,N_24632,N_24780);
nor UO_76 (O_76,N_24627,N_24775);
nand UO_77 (O_77,N_24801,N_24602);
and UO_78 (O_78,N_24813,N_24806);
and UO_79 (O_79,N_24592,N_24084);
or UO_80 (O_80,N_24025,N_24843);
and UO_81 (O_81,N_24063,N_24136);
nand UO_82 (O_82,N_24350,N_24324);
nand UO_83 (O_83,N_24342,N_24162);
nand UO_84 (O_84,N_24127,N_24138);
and UO_85 (O_85,N_24820,N_24188);
and UO_86 (O_86,N_24524,N_24949);
and UO_87 (O_87,N_24694,N_24502);
and UO_88 (O_88,N_24900,N_24507);
nor UO_89 (O_89,N_24456,N_24401);
nand UO_90 (O_90,N_24000,N_24594);
or UO_91 (O_91,N_24051,N_24366);
nor UO_92 (O_92,N_24732,N_24246);
nand UO_93 (O_93,N_24120,N_24668);
nor UO_94 (O_94,N_24909,N_24777);
or UO_95 (O_95,N_24906,N_24710);
xor UO_96 (O_96,N_24107,N_24119);
or UO_97 (O_97,N_24862,N_24665);
nor UO_98 (O_98,N_24071,N_24028);
nand UO_99 (O_99,N_24779,N_24217);
or UO_100 (O_100,N_24014,N_24123);
nand UO_101 (O_101,N_24856,N_24099);
nand UO_102 (O_102,N_24842,N_24400);
xnor UO_103 (O_103,N_24243,N_24458);
or UO_104 (O_104,N_24327,N_24227);
or UO_105 (O_105,N_24826,N_24993);
and UO_106 (O_106,N_24707,N_24043);
and UO_107 (O_107,N_24437,N_24792);
nand UO_108 (O_108,N_24944,N_24457);
nor UO_109 (O_109,N_24301,N_24855);
or UO_110 (O_110,N_24367,N_24509);
and UO_111 (O_111,N_24183,N_24216);
xor UO_112 (O_112,N_24284,N_24428);
or UO_113 (O_113,N_24177,N_24500);
and UO_114 (O_114,N_24169,N_24879);
xnor UO_115 (O_115,N_24108,N_24616);
or UO_116 (O_116,N_24967,N_24423);
and UO_117 (O_117,N_24094,N_24651);
and UO_118 (O_118,N_24149,N_24788);
or UO_119 (O_119,N_24100,N_24290);
nor UO_120 (O_120,N_24689,N_24492);
nand UO_121 (O_121,N_24104,N_24907);
xor UO_122 (O_122,N_24701,N_24125);
and UO_123 (O_123,N_24688,N_24603);
and UO_124 (O_124,N_24333,N_24228);
and UO_125 (O_125,N_24596,N_24931);
and UO_126 (O_126,N_24614,N_24008);
xor UO_127 (O_127,N_24334,N_24656);
xnor UO_128 (O_128,N_24496,N_24899);
or UO_129 (O_129,N_24418,N_24542);
nor UO_130 (O_130,N_24341,N_24678);
or UO_131 (O_131,N_24343,N_24329);
nor UO_132 (O_132,N_24462,N_24155);
or UO_133 (O_133,N_24956,N_24469);
nor UO_134 (O_134,N_24187,N_24089);
and UO_135 (O_135,N_24199,N_24316);
or UO_136 (O_136,N_24272,N_24222);
nand UO_137 (O_137,N_24464,N_24558);
and UO_138 (O_138,N_24961,N_24938);
and UO_139 (O_139,N_24802,N_24247);
nand UO_140 (O_140,N_24146,N_24812);
xor UO_141 (O_141,N_24504,N_24966);
and UO_142 (O_142,N_24168,N_24803);
xor UO_143 (O_143,N_24406,N_24090);
and UO_144 (O_144,N_24977,N_24947);
nand UO_145 (O_145,N_24447,N_24525);
or UO_146 (O_146,N_24021,N_24724);
xor UO_147 (O_147,N_24687,N_24231);
xor UO_148 (O_148,N_24098,N_24134);
xnor UO_149 (O_149,N_24096,N_24913);
or UO_150 (O_150,N_24970,N_24078);
and UO_151 (O_151,N_24589,N_24011);
nor UO_152 (O_152,N_24101,N_24652);
and UO_153 (O_153,N_24092,N_24463);
or UO_154 (O_154,N_24552,N_24362);
nor UO_155 (O_155,N_24621,N_24431);
nand UO_156 (O_156,N_24497,N_24693);
or UO_157 (O_157,N_24703,N_24536);
or UO_158 (O_158,N_24574,N_24421);
and UO_159 (O_159,N_24331,N_24195);
xor UO_160 (O_160,N_24075,N_24866);
and UO_161 (O_161,N_24680,N_24027);
nand UO_162 (O_162,N_24153,N_24761);
and UO_163 (O_163,N_24639,N_24121);
nor UO_164 (O_164,N_24690,N_24452);
nor UO_165 (O_165,N_24278,N_24572);
or UO_166 (O_166,N_24943,N_24647);
nand UO_167 (O_167,N_24522,N_24600);
nor UO_168 (O_168,N_24588,N_24482);
or UO_169 (O_169,N_24359,N_24396);
nand UO_170 (O_170,N_24032,N_24666);
nand UO_171 (O_171,N_24354,N_24299);
or UO_172 (O_172,N_24676,N_24296);
xnor UO_173 (O_173,N_24868,N_24568);
or UO_174 (O_174,N_24193,N_24575);
or UO_175 (O_175,N_24260,N_24076);
nor UO_176 (O_176,N_24764,N_24584);
or UO_177 (O_177,N_24728,N_24529);
or UO_178 (O_178,N_24054,N_24727);
nor UO_179 (O_179,N_24563,N_24205);
nor UO_180 (O_180,N_24186,N_24505);
nor UO_181 (O_181,N_24715,N_24922);
xnor UO_182 (O_182,N_24404,N_24571);
or UO_183 (O_183,N_24756,N_24357);
and UO_184 (O_184,N_24698,N_24981);
and UO_185 (O_185,N_24118,N_24607);
nor UO_186 (O_186,N_24248,N_24747);
or UO_187 (O_187,N_24275,N_24097);
nor UO_188 (O_188,N_24305,N_24905);
nand UO_189 (O_189,N_24633,N_24848);
and UO_190 (O_190,N_24786,N_24992);
nor UO_191 (O_191,N_24562,N_24111);
nand UO_192 (O_192,N_24962,N_24256);
nor UO_193 (O_193,N_24384,N_24237);
nand UO_194 (O_194,N_24355,N_24917);
and UO_195 (O_195,N_24036,N_24682);
xnor UO_196 (O_196,N_24692,N_24671);
or UO_197 (O_197,N_24439,N_24466);
nor UO_198 (O_198,N_24298,N_24581);
and UO_199 (O_199,N_24766,N_24901);
and UO_200 (O_200,N_24585,N_24768);
xnor UO_201 (O_201,N_24540,N_24646);
nand UO_202 (O_202,N_24892,N_24220);
xnor UO_203 (O_203,N_24745,N_24984);
and UO_204 (O_204,N_24723,N_24669);
and UO_205 (O_205,N_24005,N_24846);
and UO_206 (O_206,N_24695,N_24763);
and UO_207 (O_207,N_24987,N_24912);
and UO_208 (O_208,N_24270,N_24867);
and UO_209 (O_209,N_24870,N_24045);
and UO_210 (O_210,N_24915,N_24371);
xnor UO_211 (O_211,N_24499,N_24894);
or UO_212 (O_212,N_24697,N_24515);
and UO_213 (O_213,N_24713,N_24508);
nor UO_214 (O_214,N_24854,N_24310);
and UO_215 (O_215,N_24751,N_24679);
xor UO_216 (O_216,N_24232,N_24626);
and UO_217 (O_217,N_24979,N_24307);
nor UO_218 (O_218,N_24930,N_24555);
nand UO_219 (O_219,N_24748,N_24527);
and UO_220 (O_220,N_24835,N_24258);
nand UO_221 (O_221,N_24079,N_24696);
nand UO_222 (O_222,N_24062,N_24266);
nand UO_223 (O_223,N_24795,N_24648);
and UO_224 (O_224,N_24593,N_24048);
nor UO_225 (O_225,N_24441,N_24942);
or UO_226 (O_226,N_24356,N_24060);
nor UO_227 (O_227,N_24714,N_24778);
nor UO_228 (O_228,N_24185,N_24438);
or UO_229 (O_229,N_24827,N_24022);
and UO_230 (O_230,N_24629,N_24297);
and UO_231 (O_231,N_24670,N_24451);
and UO_232 (O_232,N_24239,N_24218);
xor UO_233 (O_233,N_24664,N_24399);
and UO_234 (O_234,N_24425,N_24044);
nor UO_235 (O_235,N_24049,N_24208);
xor UO_236 (O_236,N_24738,N_24851);
nand UO_237 (O_237,N_24821,N_24176);
or UO_238 (O_238,N_24459,N_24064);
nor UO_239 (O_239,N_24807,N_24958);
and UO_240 (O_240,N_24315,N_24280);
or UO_241 (O_241,N_24945,N_24964);
nor UO_242 (O_242,N_24684,N_24325);
nand UO_243 (O_243,N_24677,N_24631);
or UO_244 (O_244,N_24583,N_24268);
nand UO_245 (O_245,N_24951,N_24353);
nor UO_246 (O_246,N_24833,N_24904);
nand UO_247 (O_247,N_24202,N_24219);
nand UO_248 (O_248,N_24375,N_24013);
nor UO_249 (O_249,N_24152,N_24948);
and UO_250 (O_250,N_24965,N_24567);
xor UO_251 (O_251,N_24624,N_24031);
xor UO_252 (O_252,N_24591,N_24050);
nor UO_253 (O_253,N_24554,N_24262);
nor UO_254 (O_254,N_24817,N_24793);
and UO_255 (O_255,N_24001,N_24364);
and UO_256 (O_256,N_24557,N_24673);
and UO_257 (O_257,N_24481,N_24488);
and UO_258 (O_258,N_24590,N_24348);
xnor UO_259 (O_259,N_24773,N_24171);
and UO_260 (O_260,N_24649,N_24124);
or UO_261 (O_261,N_24929,N_24880);
or UO_262 (O_262,N_24468,N_24211);
or UO_263 (O_263,N_24088,N_24518);
and UO_264 (O_264,N_24642,N_24250);
or UO_265 (O_265,N_24608,N_24704);
or UO_266 (O_266,N_24072,N_24934);
or UO_267 (O_267,N_24147,N_24660);
nor UO_268 (O_268,N_24009,N_24772);
and UO_269 (O_269,N_24445,N_24920);
xnor UO_270 (O_270,N_24429,N_24883);
nand UO_271 (O_271,N_24189,N_24273);
or UO_272 (O_272,N_24040,N_24320);
or UO_273 (O_273,N_24839,N_24974);
nand UO_274 (O_274,N_24887,N_24323);
nor UO_275 (O_275,N_24613,N_24791);
or UO_276 (O_276,N_24115,N_24559);
nand UO_277 (O_277,N_24736,N_24257);
xor UO_278 (O_278,N_24628,N_24319);
nand UO_279 (O_279,N_24369,N_24326);
nor UO_280 (O_280,N_24741,N_24212);
nor UO_281 (O_281,N_24378,N_24828);
xnor UO_282 (O_282,N_24717,N_24102);
nor UO_283 (O_283,N_24655,N_24380);
or UO_284 (O_284,N_24198,N_24361);
nor UO_285 (O_285,N_24398,N_24416);
or UO_286 (O_286,N_24244,N_24784);
and UO_287 (O_287,N_24427,N_24067);
and UO_288 (O_288,N_24312,N_24382);
nand UO_289 (O_289,N_24240,N_24636);
nor UO_290 (O_290,N_24030,N_24910);
and UO_291 (O_291,N_24037,N_24294);
nand UO_292 (O_292,N_24718,N_24338);
or UO_293 (O_293,N_24733,N_24479);
and UO_294 (O_294,N_24283,N_24385);
or UO_295 (O_295,N_24476,N_24782);
nand UO_296 (O_296,N_24345,N_24085);
nand UO_297 (O_297,N_24061,N_24810);
nand UO_298 (O_298,N_24042,N_24512);
xor UO_299 (O_299,N_24767,N_24374);
and UO_300 (O_300,N_24520,N_24988);
and UO_301 (O_301,N_24625,N_24173);
nor UO_302 (O_302,N_24889,N_24156);
nor UO_303 (O_303,N_24167,N_24024);
or UO_304 (O_304,N_24936,N_24233);
or UO_305 (O_305,N_24397,N_24644);
xnor UO_306 (O_306,N_24225,N_24657);
or UO_307 (O_307,N_24480,N_24950);
and UO_308 (O_308,N_24087,N_24755);
and UO_309 (O_309,N_24994,N_24170);
xnor UO_310 (O_310,N_24980,N_24095);
or UO_311 (O_311,N_24012,N_24818);
or UO_312 (O_312,N_24926,N_24976);
nand UO_313 (O_313,N_24790,N_24346);
and UO_314 (O_314,N_24426,N_24599);
or UO_315 (O_315,N_24538,N_24832);
nand UO_316 (O_316,N_24007,N_24586);
nand UO_317 (O_317,N_24263,N_24840);
and UO_318 (O_318,N_24836,N_24370);
nor UO_319 (O_319,N_24150,N_24658);
and UO_320 (O_320,N_24163,N_24513);
nor UO_321 (O_321,N_24081,N_24453);
and UO_322 (O_322,N_24158,N_24271);
nand UO_323 (O_323,N_24034,N_24579);
xnor UO_324 (O_324,N_24897,N_24317);
and UO_325 (O_325,N_24433,N_24352);
and UO_326 (O_326,N_24963,N_24606);
nor UO_327 (O_327,N_24654,N_24597);
and UO_328 (O_328,N_24161,N_24157);
nand UO_329 (O_329,N_24523,N_24953);
or UO_330 (O_330,N_24164,N_24990);
nor UO_331 (O_331,N_24796,N_24521);
and UO_332 (O_332,N_24609,N_24455);
xnor UO_333 (O_333,N_24039,N_24180);
nor UO_334 (O_334,N_24313,N_24863);
or UO_335 (O_335,N_24339,N_24800);
xor UO_336 (O_336,N_24730,N_24490);
and UO_337 (O_337,N_24238,N_24477);
nand UO_338 (O_338,N_24363,N_24543);
or UO_339 (O_339,N_24794,N_24546);
or UO_340 (O_340,N_24335,N_24498);
and UO_341 (O_341,N_24408,N_24675);
nor UO_342 (O_342,N_24415,N_24046);
and UO_343 (O_343,N_24337,N_24739);
or UO_344 (O_344,N_24116,N_24844);
or UO_345 (O_345,N_24533,N_24413);
and UO_346 (O_346,N_24344,N_24873);
xor UO_347 (O_347,N_24847,N_24576);
and UO_348 (O_348,N_24991,N_24267);
xnor UO_349 (O_349,N_24797,N_24059);
and UO_350 (O_350,N_24086,N_24914);
nand UO_351 (O_351,N_24381,N_24823);
or UO_352 (O_352,N_24838,N_24174);
nand UO_353 (O_353,N_24998,N_24578);
and UO_354 (O_354,N_24712,N_24151);
xnor UO_355 (O_355,N_24303,N_24731);
and UO_356 (O_356,N_24077,N_24368);
xor UO_357 (O_357,N_24903,N_24109);
xnor UO_358 (O_358,N_24941,N_24475);
nor UO_359 (O_359,N_24110,N_24989);
or UO_360 (O_360,N_24070,N_24829);
and UO_361 (O_361,N_24875,N_24545);
nand UO_362 (O_362,N_24129,N_24241);
xor UO_363 (O_363,N_24493,N_24018);
nand UO_364 (O_364,N_24709,N_24209);
or UO_365 (O_365,N_24537,N_24349);
and UO_366 (O_366,N_24885,N_24191);
xnor UO_367 (O_367,N_24249,N_24859);
nor UO_368 (O_368,N_24017,N_24734);
nand UO_369 (O_369,N_24896,N_24610);
nor UO_370 (O_370,N_24549,N_24925);
xor UO_371 (O_371,N_24203,N_24830);
and UO_372 (O_372,N_24430,N_24983);
xnor UO_373 (O_373,N_24878,N_24849);
xor UO_374 (O_374,N_24204,N_24661);
xnor UO_375 (O_375,N_24141,N_24969);
xor UO_376 (O_376,N_24300,N_24269);
nor UO_377 (O_377,N_24391,N_24461);
nand UO_378 (O_378,N_24681,N_24442);
nand UO_379 (O_379,N_24865,N_24667);
xnor UO_380 (O_380,N_24982,N_24181);
or UO_381 (O_381,N_24470,N_24686);
and UO_382 (O_382,N_24968,N_24954);
nand UO_383 (O_383,N_24117,N_24530);
xnor UO_384 (O_384,N_24113,N_24519);
xnor UO_385 (O_385,N_24277,N_24776);
and UO_386 (O_386,N_24877,N_24143);
or UO_387 (O_387,N_24837,N_24595);
and UO_388 (O_388,N_24302,N_24960);
nand UO_389 (O_389,N_24122,N_24291);
xor UO_390 (O_390,N_24645,N_24242);
nor UO_391 (O_391,N_24638,N_24672);
xor UO_392 (O_392,N_24485,N_24448);
and UO_393 (O_393,N_24798,N_24819);
and UO_394 (O_394,N_24630,N_24860);
or UO_395 (O_395,N_24814,N_24999);
xnor UO_396 (O_396,N_24659,N_24503);
xor UO_397 (O_397,N_24570,N_24582);
xor UO_398 (O_398,N_24023,N_24226);
xor UO_399 (O_399,N_24190,N_24253);
or UO_400 (O_400,N_24973,N_24757);
nand UO_401 (O_401,N_24192,N_24619);
and UO_402 (O_402,N_24765,N_24019);
xnor UO_403 (O_403,N_24884,N_24716);
nor UO_404 (O_404,N_24166,N_24460);
and UO_405 (O_405,N_24473,N_24978);
xnor UO_406 (O_406,N_24601,N_24314);
nand UO_407 (O_407,N_24422,N_24020);
and UO_408 (O_408,N_24754,N_24215);
xnor UO_409 (O_409,N_24864,N_24783);
or UO_410 (O_410,N_24292,N_24080);
nor UO_411 (O_411,N_24114,N_24952);
xnor UO_412 (O_412,N_24495,N_24279);
nor UO_413 (O_413,N_24726,N_24916);
nor UO_414 (O_414,N_24683,N_24735);
or UO_415 (O_415,N_24946,N_24467);
or UO_416 (O_416,N_24685,N_24465);
and UO_417 (O_417,N_24230,N_24293);
nand UO_418 (O_418,N_24674,N_24304);
and UO_419 (O_419,N_24615,N_24047);
and UO_420 (O_420,N_24142,N_24785);
or UO_421 (O_421,N_24383,N_24140);
nor UO_422 (O_422,N_24106,N_24834);
or UO_423 (O_423,N_24935,N_24740);
nand UO_424 (O_424,N_24551,N_24056);
nand UO_425 (O_425,N_24434,N_24711);
and UO_426 (O_426,N_24274,N_24340);
nor UO_427 (O_427,N_24390,N_24928);
or UO_428 (O_428,N_24573,N_24308);
nand UO_429 (O_429,N_24753,N_24871);
nor UO_430 (O_430,N_24743,N_24235);
or UO_431 (O_431,N_24721,N_24996);
xnor UO_432 (O_432,N_24489,N_24811);
or UO_433 (O_433,N_24405,N_24245);
or UO_434 (O_434,N_24184,N_24759);
and UO_435 (O_435,N_24010,N_24478);
nand UO_436 (O_436,N_24940,N_24379);
nor UO_437 (O_437,N_24760,N_24933);
or UO_438 (O_438,N_24852,N_24332);
nor UO_439 (O_439,N_24815,N_24750);
nor UO_440 (O_440,N_24091,N_24506);
xnor UO_441 (O_441,N_24653,N_24746);
and UO_442 (O_442,N_24650,N_24872);
nor UO_443 (O_443,N_24002,N_24937);
nand UO_444 (O_444,N_24309,N_24234);
xnor UO_445 (O_445,N_24414,N_24286);
nor UO_446 (O_446,N_24057,N_24491);
xor UO_447 (O_447,N_24617,N_24553);
nor UO_448 (O_448,N_24444,N_24749);
and UO_449 (O_449,N_24435,N_24719);
and UO_450 (O_450,N_24440,N_24093);
nor UO_451 (O_451,N_24131,N_24770);
xnor UO_452 (O_452,N_24886,N_24069);
nor UO_453 (O_453,N_24561,N_24604);
xnor UO_454 (O_454,N_24033,N_24026);
and UO_455 (O_455,N_24133,N_24373);
xnor UO_456 (O_456,N_24055,N_24410);
and UO_457 (O_457,N_24774,N_24311);
or UO_458 (O_458,N_24103,N_24159);
xnor UO_459 (O_459,N_24449,N_24691);
or UO_460 (O_460,N_24454,N_24995);
and UO_461 (O_461,N_24517,N_24015);
or UO_462 (O_462,N_24635,N_24564);
or UO_463 (O_463,N_24565,N_24251);
or UO_464 (O_464,N_24705,N_24223);
and UO_465 (O_465,N_24321,N_24347);
nor UO_466 (O_466,N_24893,N_24620);
nand UO_467 (O_467,N_24214,N_24902);
nand UO_468 (O_468,N_24876,N_24066);
or UO_469 (O_469,N_24535,N_24318);
nand UO_470 (O_470,N_24003,N_24957);
and UO_471 (O_471,N_24787,N_24074);
xnor UO_472 (O_472,N_24541,N_24132);
xnor UO_473 (O_473,N_24539,N_24229);
and UO_474 (O_474,N_24805,N_24641);
or UO_475 (O_475,N_24577,N_24276);
xnor UO_476 (O_476,N_24853,N_24412);
nor UO_477 (O_477,N_24874,N_24112);
or UO_478 (O_478,N_24194,N_24550);
nand UO_479 (O_479,N_24474,N_24580);
nor UO_480 (O_480,N_24255,N_24816);
or UO_481 (O_481,N_24927,N_24409);
nand UO_482 (O_482,N_24526,N_24484);
and UO_483 (O_483,N_24402,N_24407);
nor UO_484 (O_484,N_24487,N_24861);
xnor UO_485 (O_485,N_24663,N_24611);
nor UO_486 (O_486,N_24799,N_24261);
nand UO_487 (O_487,N_24702,N_24126);
nand UO_488 (O_488,N_24643,N_24196);
and UO_489 (O_489,N_24053,N_24178);
nand UO_490 (O_490,N_24534,N_24443);
xor UO_491 (O_491,N_24919,N_24424);
nand UO_492 (O_492,N_24179,N_24486);
nor UO_493 (O_493,N_24041,N_24073);
xor UO_494 (O_494,N_24394,N_24052);
or UO_495 (O_495,N_24393,N_24762);
xnor UO_496 (O_496,N_24612,N_24720);
or UO_497 (O_497,N_24403,N_24891);
and UO_498 (O_498,N_24252,N_24006);
xor UO_499 (O_499,N_24395,N_24882);
or UO_500 (O_500,N_24885,N_24650);
or UO_501 (O_501,N_24052,N_24479);
or UO_502 (O_502,N_24161,N_24020);
or UO_503 (O_503,N_24341,N_24444);
nand UO_504 (O_504,N_24453,N_24019);
or UO_505 (O_505,N_24319,N_24167);
nand UO_506 (O_506,N_24555,N_24660);
or UO_507 (O_507,N_24161,N_24840);
and UO_508 (O_508,N_24537,N_24289);
xnor UO_509 (O_509,N_24001,N_24372);
xnor UO_510 (O_510,N_24253,N_24682);
and UO_511 (O_511,N_24771,N_24505);
nand UO_512 (O_512,N_24902,N_24853);
and UO_513 (O_513,N_24060,N_24443);
or UO_514 (O_514,N_24748,N_24978);
nor UO_515 (O_515,N_24901,N_24162);
nand UO_516 (O_516,N_24631,N_24786);
nand UO_517 (O_517,N_24058,N_24031);
xnor UO_518 (O_518,N_24247,N_24971);
nor UO_519 (O_519,N_24975,N_24799);
or UO_520 (O_520,N_24159,N_24132);
nor UO_521 (O_521,N_24493,N_24502);
and UO_522 (O_522,N_24478,N_24312);
or UO_523 (O_523,N_24278,N_24146);
xnor UO_524 (O_524,N_24159,N_24422);
and UO_525 (O_525,N_24187,N_24918);
and UO_526 (O_526,N_24175,N_24072);
nand UO_527 (O_527,N_24994,N_24316);
or UO_528 (O_528,N_24293,N_24254);
and UO_529 (O_529,N_24981,N_24170);
nand UO_530 (O_530,N_24274,N_24208);
and UO_531 (O_531,N_24194,N_24829);
and UO_532 (O_532,N_24871,N_24239);
and UO_533 (O_533,N_24793,N_24781);
nor UO_534 (O_534,N_24094,N_24819);
xnor UO_535 (O_535,N_24529,N_24934);
nor UO_536 (O_536,N_24350,N_24470);
or UO_537 (O_537,N_24977,N_24069);
and UO_538 (O_538,N_24993,N_24084);
nand UO_539 (O_539,N_24067,N_24613);
and UO_540 (O_540,N_24562,N_24532);
xnor UO_541 (O_541,N_24506,N_24327);
nor UO_542 (O_542,N_24667,N_24266);
nand UO_543 (O_543,N_24490,N_24669);
xnor UO_544 (O_544,N_24716,N_24683);
nand UO_545 (O_545,N_24259,N_24446);
and UO_546 (O_546,N_24873,N_24143);
nand UO_547 (O_547,N_24640,N_24132);
xnor UO_548 (O_548,N_24203,N_24769);
nor UO_549 (O_549,N_24577,N_24729);
or UO_550 (O_550,N_24400,N_24000);
xnor UO_551 (O_551,N_24823,N_24163);
nand UO_552 (O_552,N_24820,N_24256);
or UO_553 (O_553,N_24221,N_24742);
nand UO_554 (O_554,N_24136,N_24672);
nand UO_555 (O_555,N_24449,N_24922);
and UO_556 (O_556,N_24233,N_24396);
or UO_557 (O_557,N_24929,N_24699);
nor UO_558 (O_558,N_24359,N_24526);
or UO_559 (O_559,N_24243,N_24619);
nor UO_560 (O_560,N_24887,N_24387);
nor UO_561 (O_561,N_24432,N_24590);
and UO_562 (O_562,N_24983,N_24818);
nor UO_563 (O_563,N_24993,N_24450);
nor UO_564 (O_564,N_24667,N_24705);
or UO_565 (O_565,N_24030,N_24472);
and UO_566 (O_566,N_24415,N_24809);
and UO_567 (O_567,N_24251,N_24199);
nor UO_568 (O_568,N_24224,N_24047);
and UO_569 (O_569,N_24369,N_24301);
nand UO_570 (O_570,N_24051,N_24859);
nor UO_571 (O_571,N_24351,N_24176);
nand UO_572 (O_572,N_24568,N_24573);
xor UO_573 (O_573,N_24400,N_24015);
nor UO_574 (O_574,N_24789,N_24603);
nand UO_575 (O_575,N_24326,N_24010);
xor UO_576 (O_576,N_24465,N_24573);
xor UO_577 (O_577,N_24010,N_24251);
nand UO_578 (O_578,N_24469,N_24370);
or UO_579 (O_579,N_24105,N_24755);
and UO_580 (O_580,N_24361,N_24439);
or UO_581 (O_581,N_24338,N_24384);
xor UO_582 (O_582,N_24207,N_24430);
or UO_583 (O_583,N_24653,N_24606);
nor UO_584 (O_584,N_24861,N_24747);
or UO_585 (O_585,N_24893,N_24446);
nor UO_586 (O_586,N_24845,N_24807);
nand UO_587 (O_587,N_24981,N_24365);
or UO_588 (O_588,N_24530,N_24355);
and UO_589 (O_589,N_24197,N_24977);
and UO_590 (O_590,N_24990,N_24476);
nand UO_591 (O_591,N_24804,N_24892);
nand UO_592 (O_592,N_24297,N_24002);
nand UO_593 (O_593,N_24196,N_24015);
nor UO_594 (O_594,N_24451,N_24604);
nand UO_595 (O_595,N_24023,N_24847);
nor UO_596 (O_596,N_24613,N_24135);
xor UO_597 (O_597,N_24342,N_24115);
nor UO_598 (O_598,N_24843,N_24424);
xnor UO_599 (O_599,N_24878,N_24403);
nand UO_600 (O_600,N_24403,N_24838);
xor UO_601 (O_601,N_24882,N_24298);
and UO_602 (O_602,N_24846,N_24766);
or UO_603 (O_603,N_24809,N_24569);
and UO_604 (O_604,N_24930,N_24415);
nand UO_605 (O_605,N_24852,N_24059);
xor UO_606 (O_606,N_24652,N_24437);
xnor UO_607 (O_607,N_24211,N_24461);
or UO_608 (O_608,N_24171,N_24809);
or UO_609 (O_609,N_24897,N_24339);
xnor UO_610 (O_610,N_24855,N_24782);
nand UO_611 (O_611,N_24606,N_24638);
xnor UO_612 (O_612,N_24223,N_24347);
or UO_613 (O_613,N_24939,N_24034);
nand UO_614 (O_614,N_24034,N_24612);
nor UO_615 (O_615,N_24886,N_24120);
or UO_616 (O_616,N_24696,N_24874);
or UO_617 (O_617,N_24586,N_24026);
nor UO_618 (O_618,N_24960,N_24354);
nor UO_619 (O_619,N_24415,N_24405);
nand UO_620 (O_620,N_24508,N_24054);
or UO_621 (O_621,N_24533,N_24231);
and UO_622 (O_622,N_24862,N_24380);
or UO_623 (O_623,N_24192,N_24103);
nand UO_624 (O_624,N_24748,N_24129);
and UO_625 (O_625,N_24252,N_24268);
nor UO_626 (O_626,N_24575,N_24951);
and UO_627 (O_627,N_24834,N_24183);
or UO_628 (O_628,N_24785,N_24237);
nor UO_629 (O_629,N_24319,N_24633);
nor UO_630 (O_630,N_24396,N_24481);
or UO_631 (O_631,N_24773,N_24453);
nand UO_632 (O_632,N_24860,N_24500);
and UO_633 (O_633,N_24183,N_24773);
or UO_634 (O_634,N_24436,N_24229);
xnor UO_635 (O_635,N_24603,N_24843);
and UO_636 (O_636,N_24603,N_24620);
nand UO_637 (O_637,N_24985,N_24755);
xor UO_638 (O_638,N_24016,N_24515);
or UO_639 (O_639,N_24271,N_24662);
nor UO_640 (O_640,N_24281,N_24276);
and UO_641 (O_641,N_24764,N_24009);
or UO_642 (O_642,N_24348,N_24646);
or UO_643 (O_643,N_24444,N_24276);
nor UO_644 (O_644,N_24314,N_24919);
xnor UO_645 (O_645,N_24961,N_24784);
or UO_646 (O_646,N_24426,N_24111);
nor UO_647 (O_647,N_24424,N_24559);
or UO_648 (O_648,N_24326,N_24461);
or UO_649 (O_649,N_24019,N_24995);
or UO_650 (O_650,N_24317,N_24981);
and UO_651 (O_651,N_24717,N_24043);
nand UO_652 (O_652,N_24798,N_24905);
xnor UO_653 (O_653,N_24050,N_24335);
and UO_654 (O_654,N_24568,N_24284);
xor UO_655 (O_655,N_24178,N_24764);
and UO_656 (O_656,N_24879,N_24453);
and UO_657 (O_657,N_24677,N_24039);
or UO_658 (O_658,N_24876,N_24921);
nand UO_659 (O_659,N_24301,N_24857);
nor UO_660 (O_660,N_24685,N_24381);
nor UO_661 (O_661,N_24299,N_24881);
or UO_662 (O_662,N_24249,N_24332);
and UO_663 (O_663,N_24736,N_24839);
nand UO_664 (O_664,N_24689,N_24596);
nor UO_665 (O_665,N_24166,N_24013);
or UO_666 (O_666,N_24451,N_24030);
nor UO_667 (O_667,N_24442,N_24561);
and UO_668 (O_668,N_24329,N_24993);
or UO_669 (O_669,N_24104,N_24990);
and UO_670 (O_670,N_24489,N_24365);
nand UO_671 (O_671,N_24090,N_24845);
nand UO_672 (O_672,N_24626,N_24102);
or UO_673 (O_673,N_24565,N_24574);
xnor UO_674 (O_674,N_24953,N_24720);
or UO_675 (O_675,N_24969,N_24786);
or UO_676 (O_676,N_24945,N_24654);
nand UO_677 (O_677,N_24775,N_24940);
nor UO_678 (O_678,N_24634,N_24925);
nor UO_679 (O_679,N_24074,N_24013);
and UO_680 (O_680,N_24745,N_24634);
nand UO_681 (O_681,N_24905,N_24561);
xor UO_682 (O_682,N_24874,N_24672);
nor UO_683 (O_683,N_24559,N_24085);
nor UO_684 (O_684,N_24873,N_24501);
or UO_685 (O_685,N_24420,N_24360);
or UO_686 (O_686,N_24174,N_24877);
nor UO_687 (O_687,N_24185,N_24519);
or UO_688 (O_688,N_24348,N_24233);
nor UO_689 (O_689,N_24833,N_24699);
nor UO_690 (O_690,N_24196,N_24684);
and UO_691 (O_691,N_24915,N_24648);
and UO_692 (O_692,N_24960,N_24197);
nand UO_693 (O_693,N_24855,N_24305);
nor UO_694 (O_694,N_24177,N_24311);
nor UO_695 (O_695,N_24308,N_24604);
nor UO_696 (O_696,N_24392,N_24942);
xnor UO_697 (O_697,N_24027,N_24582);
nand UO_698 (O_698,N_24273,N_24697);
and UO_699 (O_699,N_24039,N_24456);
nand UO_700 (O_700,N_24072,N_24865);
nor UO_701 (O_701,N_24779,N_24353);
and UO_702 (O_702,N_24030,N_24855);
or UO_703 (O_703,N_24541,N_24632);
or UO_704 (O_704,N_24732,N_24345);
and UO_705 (O_705,N_24953,N_24753);
xnor UO_706 (O_706,N_24974,N_24453);
xor UO_707 (O_707,N_24358,N_24859);
xnor UO_708 (O_708,N_24923,N_24784);
xnor UO_709 (O_709,N_24552,N_24264);
xor UO_710 (O_710,N_24686,N_24072);
nand UO_711 (O_711,N_24220,N_24994);
xnor UO_712 (O_712,N_24436,N_24446);
and UO_713 (O_713,N_24343,N_24639);
xnor UO_714 (O_714,N_24178,N_24882);
nor UO_715 (O_715,N_24868,N_24702);
or UO_716 (O_716,N_24486,N_24654);
nor UO_717 (O_717,N_24587,N_24474);
xnor UO_718 (O_718,N_24097,N_24994);
and UO_719 (O_719,N_24931,N_24349);
nor UO_720 (O_720,N_24057,N_24271);
nor UO_721 (O_721,N_24944,N_24354);
or UO_722 (O_722,N_24144,N_24781);
or UO_723 (O_723,N_24071,N_24216);
nand UO_724 (O_724,N_24054,N_24000);
and UO_725 (O_725,N_24086,N_24445);
nand UO_726 (O_726,N_24989,N_24491);
or UO_727 (O_727,N_24104,N_24773);
nor UO_728 (O_728,N_24100,N_24696);
or UO_729 (O_729,N_24582,N_24798);
and UO_730 (O_730,N_24454,N_24226);
nand UO_731 (O_731,N_24020,N_24300);
or UO_732 (O_732,N_24452,N_24877);
nor UO_733 (O_733,N_24086,N_24807);
nand UO_734 (O_734,N_24850,N_24630);
xor UO_735 (O_735,N_24150,N_24754);
nor UO_736 (O_736,N_24610,N_24980);
nand UO_737 (O_737,N_24292,N_24828);
or UO_738 (O_738,N_24186,N_24148);
and UO_739 (O_739,N_24866,N_24250);
xor UO_740 (O_740,N_24599,N_24090);
or UO_741 (O_741,N_24579,N_24517);
nor UO_742 (O_742,N_24099,N_24715);
or UO_743 (O_743,N_24103,N_24832);
and UO_744 (O_744,N_24944,N_24112);
and UO_745 (O_745,N_24279,N_24461);
xor UO_746 (O_746,N_24771,N_24132);
nand UO_747 (O_747,N_24498,N_24665);
and UO_748 (O_748,N_24169,N_24998);
or UO_749 (O_749,N_24911,N_24516);
or UO_750 (O_750,N_24776,N_24868);
or UO_751 (O_751,N_24204,N_24035);
and UO_752 (O_752,N_24895,N_24111);
xnor UO_753 (O_753,N_24936,N_24853);
or UO_754 (O_754,N_24300,N_24254);
xnor UO_755 (O_755,N_24335,N_24979);
xnor UO_756 (O_756,N_24030,N_24461);
nor UO_757 (O_757,N_24433,N_24841);
nand UO_758 (O_758,N_24311,N_24185);
nor UO_759 (O_759,N_24780,N_24271);
or UO_760 (O_760,N_24501,N_24263);
nor UO_761 (O_761,N_24474,N_24550);
xnor UO_762 (O_762,N_24868,N_24300);
nand UO_763 (O_763,N_24634,N_24455);
or UO_764 (O_764,N_24737,N_24334);
nor UO_765 (O_765,N_24737,N_24677);
xnor UO_766 (O_766,N_24798,N_24395);
nor UO_767 (O_767,N_24373,N_24309);
nor UO_768 (O_768,N_24386,N_24078);
nor UO_769 (O_769,N_24692,N_24772);
or UO_770 (O_770,N_24682,N_24650);
or UO_771 (O_771,N_24699,N_24052);
nand UO_772 (O_772,N_24301,N_24771);
or UO_773 (O_773,N_24816,N_24397);
and UO_774 (O_774,N_24333,N_24184);
nand UO_775 (O_775,N_24654,N_24968);
and UO_776 (O_776,N_24863,N_24675);
nor UO_777 (O_777,N_24145,N_24324);
or UO_778 (O_778,N_24638,N_24843);
and UO_779 (O_779,N_24446,N_24769);
xnor UO_780 (O_780,N_24064,N_24313);
xor UO_781 (O_781,N_24084,N_24371);
nor UO_782 (O_782,N_24712,N_24074);
xnor UO_783 (O_783,N_24925,N_24240);
nand UO_784 (O_784,N_24405,N_24705);
and UO_785 (O_785,N_24590,N_24135);
or UO_786 (O_786,N_24862,N_24682);
or UO_787 (O_787,N_24276,N_24956);
and UO_788 (O_788,N_24013,N_24734);
nor UO_789 (O_789,N_24813,N_24382);
xor UO_790 (O_790,N_24037,N_24132);
xnor UO_791 (O_791,N_24078,N_24148);
nor UO_792 (O_792,N_24215,N_24252);
and UO_793 (O_793,N_24556,N_24836);
xnor UO_794 (O_794,N_24075,N_24241);
or UO_795 (O_795,N_24043,N_24706);
nand UO_796 (O_796,N_24157,N_24845);
xor UO_797 (O_797,N_24866,N_24919);
and UO_798 (O_798,N_24385,N_24678);
nor UO_799 (O_799,N_24934,N_24338);
and UO_800 (O_800,N_24217,N_24273);
and UO_801 (O_801,N_24460,N_24972);
and UO_802 (O_802,N_24641,N_24911);
and UO_803 (O_803,N_24889,N_24035);
xnor UO_804 (O_804,N_24292,N_24025);
or UO_805 (O_805,N_24849,N_24043);
nand UO_806 (O_806,N_24756,N_24854);
nand UO_807 (O_807,N_24472,N_24127);
and UO_808 (O_808,N_24898,N_24055);
nor UO_809 (O_809,N_24020,N_24961);
and UO_810 (O_810,N_24554,N_24953);
nand UO_811 (O_811,N_24350,N_24337);
nor UO_812 (O_812,N_24946,N_24511);
and UO_813 (O_813,N_24392,N_24823);
nor UO_814 (O_814,N_24193,N_24112);
and UO_815 (O_815,N_24594,N_24801);
nand UO_816 (O_816,N_24821,N_24447);
nand UO_817 (O_817,N_24893,N_24907);
nor UO_818 (O_818,N_24786,N_24732);
nand UO_819 (O_819,N_24923,N_24929);
and UO_820 (O_820,N_24098,N_24506);
xnor UO_821 (O_821,N_24389,N_24074);
and UO_822 (O_822,N_24096,N_24901);
xor UO_823 (O_823,N_24366,N_24879);
nor UO_824 (O_824,N_24581,N_24540);
and UO_825 (O_825,N_24331,N_24964);
xnor UO_826 (O_826,N_24013,N_24237);
xor UO_827 (O_827,N_24050,N_24081);
and UO_828 (O_828,N_24205,N_24809);
nor UO_829 (O_829,N_24691,N_24350);
xor UO_830 (O_830,N_24265,N_24587);
nor UO_831 (O_831,N_24539,N_24112);
or UO_832 (O_832,N_24544,N_24143);
xnor UO_833 (O_833,N_24538,N_24550);
xnor UO_834 (O_834,N_24885,N_24704);
xnor UO_835 (O_835,N_24834,N_24904);
nor UO_836 (O_836,N_24152,N_24885);
nor UO_837 (O_837,N_24833,N_24838);
or UO_838 (O_838,N_24676,N_24769);
xnor UO_839 (O_839,N_24131,N_24399);
xor UO_840 (O_840,N_24246,N_24029);
nand UO_841 (O_841,N_24450,N_24077);
or UO_842 (O_842,N_24022,N_24714);
and UO_843 (O_843,N_24560,N_24593);
and UO_844 (O_844,N_24275,N_24089);
xnor UO_845 (O_845,N_24018,N_24983);
and UO_846 (O_846,N_24273,N_24080);
or UO_847 (O_847,N_24377,N_24047);
nor UO_848 (O_848,N_24193,N_24026);
or UO_849 (O_849,N_24983,N_24687);
nand UO_850 (O_850,N_24034,N_24205);
or UO_851 (O_851,N_24279,N_24969);
nor UO_852 (O_852,N_24747,N_24755);
nand UO_853 (O_853,N_24641,N_24088);
xor UO_854 (O_854,N_24707,N_24066);
or UO_855 (O_855,N_24694,N_24308);
and UO_856 (O_856,N_24472,N_24650);
nor UO_857 (O_857,N_24273,N_24727);
and UO_858 (O_858,N_24744,N_24762);
nand UO_859 (O_859,N_24836,N_24632);
xor UO_860 (O_860,N_24972,N_24683);
and UO_861 (O_861,N_24520,N_24604);
and UO_862 (O_862,N_24804,N_24602);
nor UO_863 (O_863,N_24782,N_24841);
xor UO_864 (O_864,N_24272,N_24813);
xnor UO_865 (O_865,N_24839,N_24301);
nor UO_866 (O_866,N_24115,N_24336);
nor UO_867 (O_867,N_24571,N_24530);
or UO_868 (O_868,N_24328,N_24975);
or UO_869 (O_869,N_24358,N_24014);
nand UO_870 (O_870,N_24497,N_24922);
nor UO_871 (O_871,N_24784,N_24878);
xnor UO_872 (O_872,N_24524,N_24297);
nor UO_873 (O_873,N_24725,N_24108);
nand UO_874 (O_874,N_24560,N_24262);
xor UO_875 (O_875,N_24326,N_24372);
xor UO_876 (O_876,N_24308,N_24699);
and UO_877 (O_877,N_24045,N_24331);
nor UO_878 (O_878,N_24878,N_24710);
nand UO_879 (O_879,N_24498,N_24397);
nor UO_880 (O_880,N_24874,N_24784);
xor UO_881 (O_881,N_24978,N_24737);
xor UO_882 (O_882,N_24441,N_24952);
or UO_883 (O_883,N_24613,N_24533);
and UO_884 (O_884,N_24402,N_24309);
and UO_885 (O_885,N_24287,N_24895);
or UO_886 (O_886,N_24685,N_24590);
nor UO_887 (O_887,N_24570,N_24872);
xnor UO_888 (O_888,N_24626,N_24089);
nand UO_889 (O_889,N_24702,N_24309);
and UO_890 (O_890,N_24326,N_24137);
or UO_891 (O_891,N_24222,N_24070);
nand UO_892 (O_892,N_24256,N_24554);
nand UO_893 (O_893,N_24255,N_24375);
and UO_894 (O_894,N_24702,N_24802);
and UO_895 (O_895,N_24762,N_24757);
nand UO_896 (O_896,N_24821,N_24056);
and UO_897 (O_897,N_24579,N_24713);
xor UO_898 (O_898,N_24502,N_24191);
and UO_899 (O_899,N_24151,N_24609);
or UO_900 (O_900,N_24300,N_24304);
nor UO_901 (O_901,N_24830,N_24001);
nor UO_902 (O_902,N_24430,N_24379);
or UO_903 (O_903,N_24192,N_24667);
or UO_904 (O_904,N_24907,N_24476);
xnor UO_905 (O_905,N_24540,N_24430);
nor UO_906 (O_906,N_24761,N_24164);
xor UO_907 (O_907,N_24382,N_24642);
xor UO_908 (O_908,N_24872,N_24639);
nand UO_909 (O_909,N_24629,N_24449);
nand UO_910 (O_910,N_24453,N_24214);
or UO_911 (O_911,N_24238,N_24574);
nor UO_912 (O_912,N_24189,N_24483);
nand UO_913 (O_913,N_24909,N_24313);
and UO_914 (O_914,N_24752,N_24193);
and UO_915 (O_915,N_24659,N_24056);
nor UO_916 (O_916,N_24350,N_24358);
nor UO_917 (O_917,N_24294,N_24365);
and UO_918 (O_918,N_24265,N_24361);
and UO_919 (O_919,N_24467,N_24742);
nor UO_920 (O_920,N_24941,N_24982);
nand UO_921 (O_921,N_24736,N_24441);
nand UO_922 (O_922,N_24978,N_24639);
nor UO_923 (O_923,N_24540,N_24683);
nand UO_924 (O_924,N_24365,N_24096);
xor UO_925 (O_925,N_24344,N_24257);
xnor UO_926 (O_926,N_24245,N_24287);
xnor UO_927 (O_927,N_24225,N_24151);
nor UO_928 (O_928,N_24872,N_24042);
nor UO_929 (O_929,N_24590,N_24678);
or UO_930 (O_930,N_24048,N_24552);
and UO_931 (O_931,N_24567,N_24856);
nor UO_932 (O_932,N_24295,N_24672);
nor UO_933 (O_933,N_24472,N_24605);
nand UO_934 (O_934,N_24281,N_24807);
xor UO_935 (O_935,N_24064,N_24473);
nor UO_936 (O_936,N_24744,N_24336);
or UO_937 (O_937,N_24405,N_24604);
xnor UO_938 (O_938,N_24997,N_24092);
xor UO_939 (O_939,N_24334,N_24317);
nor UO_940 (O_940,N_24772,N_24122);
xor UO_941 (O_941,N_24169,N_24144);
xor UO_942 (O_942,N_24031,N_24815);
xor UO_943 (O_943,N_24616,N_24986);
nor UO_944 (O_944,N_24321,N_24023);
nor UO_945 (O_945,N_24099,N_24535);
or UO_946 (O_946,N_24500,N_24785);
xor UO_947 (O_947,N_24807,N_24242);
or UO_948 (O_948,N_24667,N_24491);
xnor UO_949 (O_949,N_24230,N_24355);
xnor UO_950 (O_950,N_24195,N_24413);
and UO_951 (O_951,N_24865,N_24642);
and UO_952 (O_952,N_24369,N_24108);
xor UO_953 (O_953,N_24442,N_24458);
xnor UO_954 (O_954,N_24355,N_24328);
and UO_955 (O_955,N_24975,N_24790);
and UO_956 (O_956,N_24283,N_24524);
xor UO_957 (O_957,N_24960,N_24006);
or UO_958 (O_958,N_24543,N_24258);
or UO_959 (O_959,N_24164,N_24444);
or UO_960 (O_960,N_24023,N_24814);
nor UO_961 (O_961,N_24628,N_24100);
or UO_962 (O_962,N_24501,N_24620);
nor UO_963 (O_963,N_24625,N_24192);
nor UO_964 (O_964,N_24601,N_24100);
xor UO_965 (O_965,N_24197,N_24521);
nor UO_966 (O_966,N_24375,N_24639);
nor UO_967 (O_967,N_24841,N_24344);
and UO_968 (O_968,N_24828,N_24398);
and UO_969 (O_969,N_24718,N_24236);
and UO_970 (O_970,N_24662,N_24555);
or UO_971 (O_971,N_24899,N_24823);
and UO_972 (O_972,N_24115,N_24932);
nand UO_973 (O_973,N_24827,N_24499);
nor UO_974 (O_974,N_24637,N_24670);
xnor UO_975 (O_975,N_24116,N_24068);
and UO_976 (O_976,N_24651,N_24870);
nand UO_977 (O_977,N_24933,N_24184);
xor UO_978 (O_978,N_24337,N_24032);
xor UO_979 (O_979,N_24119,N_24749);
or UO_980 (O_980,N_24184,N_24584);
nor UO_981 (O_981,N_24719,N_24103);
nand UO_982 (O_982,N_24190,N_24819);
or UO_983 (O_983,N_24893,N_24042);
and UO_984 (O_984,N_24115,N_24204);
xor UO_985 (O_985,N_24247,N_24214);
nor UO_986 (O_986,N_24955,N_24881);
xor UO_987 (O_987,N_24091,N_24267);
nand UO_988 (O_988,N_24076,N_24030);
xor UO_989 (O_989,N_24408,N_24825);
and UO_990 (O_990,N_24507,N_24398);
nand UO_991 (O_991,N_24247,N_24647);
and UO_992 (O_992,N_24976,N_24284);
nand UO_993 (O_993,N_24571,N_24657);
xnor UO_994 (O_994,N_24905,N_24419);
and UO_995 (O_995,N_24992,N_24743);
or UO_996 (O_996,N_24333,N_24928);
nor UO_997 (O_997,N_24349,N_24377);
and UO_998 (O_998,N_24805,N_24685);
or UO_999 (O_999,N_24596,N_24307);
or UO_1000 (O_1000,N_24042,N_24719);
nor UO_1001 (O_1001,N_24110,N_24365);
and UO_1002 (O_1002,N_24790,N_24015);
nor UO_1003 (O_1003,N_24410,N_24216);
xor UO_1004 (O_1004,N_24137,N_24728);
nor UO_1005 (O_1005,N_24381,N_24873);
nand UO_1006 (O_1006,N_24581,N_24620);
nand UO_1007 (O_1007,N_24948,N_24732);
or UO_1008 (O_1008,N_24732,N_24520);
or UO_1009 (O_1009,N_24306,N_24521);
and UO_1010 (O_1010,N_24108,N_24047);
and UO_1011 (O_1011,N_24254,N_24140);
xor UO_1012 (O_1012,N_24937,N_24205);
nor UO_1013 (O_1013,N_24085,N_24188);
nor UO_1014 (O_1014,N_24506,N_24427);
xnor UO_1015 (O_1015,N_24676,N_24235);
xnor UO_1016 (O_1016,N_24718,N_24995);
nor UO_1017 (O_1017,N_24257,N_24137);
nand UO_1018 (O_1018,N_24116,N_24584);
nor UO_1019 (O_1019,N_24700,N_24433);
nor UO_1020 (O_1020,N_24886,N_24373);
xnor UO_1021 (O_1021,N_24501,N_24474);
xnor UO_1022 (O_1022,N_24146,N_24592);
and UO_1023 (O_1023,N_24069,N_24083);
and UO_1024 (O_1024,N_24794,N_24402);
nor UO_1025 (O_1025,N_24620,N_24793);
nand UO_1026 (O_1026,N_24600,N_24943);
or UO_1027 (O_1027,N_24412,N_24564);
nor UO_1028 (O_1028,N_24158,N_24931);
or UO_1029 (O_1029,N_24834,N_24677);
nand UO_1030 (O_1030,N_24244,N_24112);
xor UO_1031 (O_1031,N_24100,N_24799);
nand UO_1032 (O_1032,N_24990,N_24947);
and UO_1033 (O_1033,N_24812,N_24370);
nor UO_1034 (O_1034,N_24365,N_24684);
xor UO_1035 (O_1035,N_24195,N_24344);
xnor UO_1036 (O_1036,N_24234,N_24436);
xnor UO_1037 (O_1037,N_24983,N_24514);
nor UO_1038 (O_1038,N_24841,N_24051);
nand UO_1039 (O_1039,N_24258,N_24977);
xor UO_1040 (O_1040,N_24001,N_24750);
and UO_1041 (O_1041,N_24308,N_24316);
or UO_1042 (O_1042,N_24200,N_24284);
and UO_1043 (O_1043,N_24315,N_24567);
xor UO_1044 (O_1044,N_24556,N_24423);
or UO_1045 (O_1045,N_24743,N_24873);
nor UO_1046 (O_1046,N_24134,N_24861);
and UO_1047 (O_1047,N_24285,N_24549);
nor UO_1048 (O_1048,N_24281,N_24614);
or UO_1049 (O_1049,N_24574,N_24075);
nand UO_1050 (O_1050,N_24002,N_24284);
xnor UO_1051 (O_1051,N_24271,N_24290);
and UO_1052 (O_1052,N_24175,N_24411);
nor UO_1053 (O_1053,N_24323,N_24769);
xnor UO_1054 (O_1054,N_24066,N_24648);
nand UO_1055 (O_1055,N_24982,N_24469);
and UO_1056 (O_1056,N_24578,N_24287);
or UO_1057 (O_1057,N_24080,N_24985);
nand UO_1058 (O_1058,N_24780,N_24161);
nor UO_1059 (O_1059,N_24577,N_24460);
or UO_1060 (O_1060,N_24207,N_24149);
xor UO_1061 (O_1061,N_24561,N_24010);
nor UO_1062 (O_1062,N_24574,N_24389);
and UO_1063 (O_1063,N_24439,N_24562);
nor UO_1064 (O_1064,N_24655,N_24619);
xor UO_1065 (O_1065,N_24277,N_24992);
and UO_1066 (O_1066,N_24115,N_24176);
nand UO_1067 (O_1067,N_24301,N_24319);
or UO_1068 (O_1068,N_24918,N_24212);
and UO_1069 (O_1069,N_24620,N_24610);
nor UO_1070 (O_1070,N_24296,N_24917);
or UO_1071 (O_1071,N_24765,N_24302);
nor UO_1072 (O_1072,N_24207,N_24028);
and UO_1073 (O_1073,N_24778,N_24338);
nor UO_1074 (O_1074,N_24250,N_24576);
and UO_1075 (O_1075,N_24499,N_24114);
nand UO_1076 (O_1076,N_24490,N_24849);
and UO_1077 (O_1077,N_24641,N_24696);
xnor UO_1078 (O_1078,N_24726,N_24586);
nand UO_1079 (O_1079,N_24203,N_24125);
nor UO_1080 (O_1080,N_24352,N_24384);
nand UO_1081 (O_1081,N_24935,N_24992);
xnor UO_1082 (O_1082,N_24337,N_24081);
or UO_1083 (O_1083,N_24589,N_24685);
nand UO_1084 (O_1084,N_24467,N_24120);
and UO_1085 (O_1085,N_24475,N_24007);
nor UO_1086 (O_1086,N_24507,N_24524);
xor UO_1087 (O_1087,N_24119,N_24177);
or UO_1088 (O_1088,N_24960,N_24553);
nor UO_1089 (O_1089,N_24732,N_24132);
nor UO_1090 (O_1090,N_24159,N_24341);
or UO_1091 (O_1091,N_24366,N_24785);
or UO_1092 (O_1092,N_24509,N_24106);
nand UO_1093 (O_1093,N_24278,N_24283);
and UO_1094 (O_1094,N_24761,N_24699);
or UO_1095 (O_1095,N_24124,N_24667);
nand UO_1096 (O_1096,N_24694,N_24592);
or UO_1097 (O_1097,N_24427,N_24971);
or UO_1098 (O_1098,N_24192,N_24811);
nand UO_1099 (O_1099,N_24529,N_24675);
or UO_1100 (O_1100,N_24289,N_24691);
and UO_1101 (O_1101,N_24417,N_24928);
and UO_1102 (O_1102,N_24640,N_24018);
xnor UO_1103 (O_1103,N_24319,N_24074);
xor UO_1104 (O_1104,N_24780,N_24226);
nand UO_1105 (O_1105,N_24268,N_24700);
nand UO_1106 (O_1106,N_24136,N_24500);
nand UO_1107 (O_1107,N_24539,N_24598);
or UO_1108 (O_1108,N_24641,N_24693);
and UO_1109 (O_1109,N_24287,N_24361);
and UO_1110 (O_1110,N_24902,N_24763);
xnor UO_1111 (O_1111,N_24170,N_24445);
or UO_1112 (O_1112,N_24130,N_24143);
and UO_1113 (O_1113,N_24592,N_24885);
xnor UO_1114 (O_1114,N_24030,N_24337);
and UO_1115 (O_1115,N_24236,N_24695);
nand UO_1116 (O_1116,N_24593,N_24982);
nand UO_1117 (O_1117,N_24945,N_24776);
xor UO_1118 (O_1118,N_24914,N_24473);
xor UO_1119 (O_1119,N_24000,N_24686);
and UO_1120 (O_1120,N_24406,N_24133);
or UO_1121 (O_1121,N_24826,N_24576);
xor UO_1122 (O_1122,N_24422,N_24919);
nand UO_1123 (O_1123,N_24120,N_24266);
nand UO_1124 (O_1124,N_24779,N_24078);
or UO_1125 (O_1125,N_24952,N_24732);
and UO_1126 (O_1126,N_24786,N_24064);
nand UO_1127 (O_1127,N_24250,N_24681);
nand UO_1128 (O_1128,N_24676,N_24955);
or UO_1129 (O_1129,N_24602,N_24065);
xnor UO_1130 (O_1130,N_24012,N_24517);
nor UO_1131 (O_1131,N_24272,N_24902);
or UO_1132 (O_1132,N_24341,N_24535);
xnor UO_1133 (O_1133,N_24642,N_24146);
xnor UO_1134 (O_1134,N_24446,N_24632);
or UO_1135 (O_1135,N_24485,N_24904);
nor UO_1136 (O_1136,N_24566,N_24290);
nand UO_1137 (O_1137,N_24833,N_24511);
nand UO_1138 (O_1138,N_24047,N_24408);
and UO_1139 (O_1139,N_24199,N_24426);
nand UO_1140 (O_1140,N_24444,N_24981);
and UO_1141 (O_1141,N_24469,N_24466);
or UO_1142 (O_1142,N_24373,N_24968);
xor UO_1143 (O_1143,N_24694,N_24902);
and UO_1144 (O_1144,N_24978,N_24478);
nor UO_1145 (O_1145,N_24477,N_24006);
xor UO_1146 (O_1146,N_24613,N_24217);
nand UO_1147 (O_1147,N_24879,N_24581);
and UO_1148 (O_1148,N_24859,N_24157);
xor UO_1149 (O_1149,N_24551,N_24256);
nand UO_1150 (O_1150,N_24170,N_24442);
xnor UO_1151 (O_1151,N_24260,N_24277);
xnor UO_1152 (O_1152,N_24444,N_24372);
nor UO_1153 (O_1153,N_24704,N_24921);
xor UO_1154 (O_1154,N_24294,N_24315);
nand UO_1155 (O_1155,N_24653,N_24398);
xnor UO_1156 (O_1156,N_24824,N_24884);
nand UO_1157 (O_1157,N_24839,N_24368);
nand UO_1158 (O_1158,N_24443,N_24888);
and UO_1159 (O_1159,N_24864,N_24902);
nor UO_1160 (O_1160,N_24411,N_24904);
or UO_1161 (O_1161,N_24540,N_24389);
xor UO_1162 (O_1162,N_24672,N_24257);
xor UO_1163 (O_1163,N_24247,N_24645);
xnor UO_1164 (O_1164,N_24886,N_24268);
nand UO_1165 (O_1165,N_24305,N_24090);
xor UO_1166 (O_1166,N_24218,N_24113);
nand UO_1167 (O_1167,N_24036,N_24432);
nor UO_1168 (O_1168,N_24987,N_24572);
or UO_1169 (O_1169,N_24187,N_24632);
nor UO_1170 (O_1170,N_24507,N_24034);
or UO_1171 (O_1171,N_24266,N_24962);
nor UO_1172 (O_1172,N_24116,N_24679);
nand UO_1173 (O_1173,N_24446,N_24541);
xnor UO_1174 (O_1174,N_24004,N_24876);
nand UO_1175 (O_1175,N_24820,N_24709);
or UO_1176 (O_1176,N_24863,N_24631);
or UO_1177 (O_1177,N_24529,N_24120);
or UO_1178 (O_1178,N_24971,N_24319);
nor UO_1179 (O_1179,N_24280,N_24508);
or UO_1180 (O_1180,N_24198,N_24156);
nand UO_1181 (O_1181,N_24457,N_24523);
or UO_1182 (O_1182,N_24269,N_24918);
nor UO_1183 (O_1183,N_24682,N_24720);
or UO_1184 (O_1184,N_24177,N_24364);
and UO_1185 (O_1185,N_24905,N_24216);
and UO_1186 (O_1186,N_24702,N_24854);
and UO_1187 (O_1187,N_24119,N_24432);
or UO_1188 (O_1188,N_24360,N_24693);
and UO_1189 (O_1189,N_24474,N_24258);
xnor UO_1190 (O_1190,N_24168,N_24454);
xor UO_1191 (O_1191,N_24415,N_24447);
nor UO_1192 (O_1192,N_24116,N_24151);
or UO_1193 (O_1193,N_24084,N_24556);
xor UO_1194 (O_1194,N_24306,N_24118);
nor UO_1195 (O_1195,N_24682,N_24614);
or UO_1196 (O_1196,N_24781,N_24010);
and UO_1197 (O_1197,N_24861,N_24072);
or UO_1198 (O_1198,N_24260,N_24110);
nor UO_1199 (O_1199,N_24681,N_24842);
nor UO_1200 (O_1200,N_24932,N_24841);
xnor UO_1201 (O_1201,N_24704,N_24853);
xnor UO_1202 (O_1202,N_24183,N_24162);
xor UO_1203 (O_1203,N_24623,N_24603);
or UO_1204 (O_1204,N_24144,N_24847);
nand UO_1205 (O_1205,N_24618,N_24978);
and UO_1206 (O_1206,N_24279,N_24105);
or UO_1207 (O_1207,N_24568,N_24111);
xor UO_1208 (O_1208,N_24280,N_24741);
or UO_1209 (O_1209,N_24920,N_24834);
and UO_1210 (O_1210,N_24022,N_24883);
nor UO_1211 (O_1211,N_24296,N_24279);
nand UO_1212 (O_1212,N_24792,N_24123);
and UO_1213 (O_1213,N_24675,N_24345);
nand UO_1214 (O_1214,N_24121,N_24033);
or UO_1215 (O_1215,N_24633,N_24925);
and UO_1216 (O_1216,N_24759,N_24701);
and UO_1217 (O_1217,N_24271,N_24933);
xnor UO_1218 (O_1218,N_24184,N_24537);
nor UO_1219 (O_1219,N_24144,N_24178);
or UO_1220 (O_1220,N_24656,N_24864);
nor UO_1221 (O_1221,N_24817,N_24122);
or UO_1222 (O_1222,N_24551,N_24287);
or UO_1223 (O_1223,N_24977,N_24268);
and UO_1224 (O_1224,N_24704,N_24258);
and UO_1225 (O_1225,N_24005,N_24521);
nor UO_1226 (O_1226,N_24724,N_24471);
nor UO_1227 (O_1227,N_24898,N_24519);
or UO_1228 (O_1228,N_24410,N_24475);
xor UO_1229 (O_1229,N_24996,N_24695);
xnor UO_1230 (O_1230,N_24602,N_24508);
nor UO_1231 (O_1231,N_24320,N_24229);
xnor UO_1232 (O_1232,N_24578,N_24128);
or UO_1233 (O_1233,N_24910,N_24410);
nand UO_1234 (O_1234,N_24193,N_24807);
nor UO_1235 (O_1235,N_24241,N_24193);
xor UO_1236 (O_1236,N_24695,N_24704);
or UO_1237 (O_1237,N_24047,N_24881);
nor UO_1238 (O_1238,N_24617,N_24159);
or UO_1239 (O_1239,N_24307,N_24078);
or UO_1240 (O_1240,N_24048,N_24557);
or UO_1241 (O_1241,N_24108,N_24717);
and UO_1242 (O_1242,N_24743,N_24180);
and UO_1243 (O_1243,N_24747,N_24090);
xor UO_1244 (O_1244,N_24225,N_24614);
nand UO_1245 (O_1245,N_24432,N_24570);
and UO_1246 (O_1246,N_24781,N_24002);
xor UO_1247 (O_1247,N_24326,N_24913);
xor UO_1248 (O_1248,N_24542,N_24169);
or UO_1249 (O_1249,N_24599,N_24508);
nand UO_1250 (O_1250,N_24761,N_24417);
or UO_1251 (O_1251,N_24935,N_24845);
xnor UO_1252 (O_1252,N_24134,N_24791);
and UO_1253 (O_1253,N_24680,N_24988);
or UO_1254 (O_1254,N_24950,N_24898);
and UO_1255 (O_1255,N_24074,N_24780);
nand UO_1256 (O_1256,N_24274,N_24938);
xor UO_1257 (O_1257,N_24764,N_24102);
xnor UO_1258 (O_1258,N_24422,N_24069);
nand UO_1259 (O_1259,N_24408,N_24352);
nor UO_1260 (O_1260,N_24017,N_24179);
nand UO_1261 (O_1261,N_24870,N_24157);
nand UO_1262 (O_1262,N_24663,N_24882);
xor UO_1263 (O_1263,N_24980,N_24746);
and UO_1264 (O_1264,N_24318,N_24170);
nand UO_1265 (O_1265,N_24373,N_24742);
and UO_1266 (O_1266,N_24228,N_24367);
nor UO_1267 (O_1267,N_24854,N_24069);
or UO_1268 (O_1268,N_24165,N_24775);
or UO_1269 (O_1269,N_24082,N_24127);
nor UO_1270 (O_1270,N_24489,N_24298);
nor UO_1271 (O_1271,N_24607,N_24345);
and UO_1272 (O_1272,N_24557,N_24968);
or UO_1273 (O_1273,N_24993,N_24011);
and UO_1274 (O_1274,N_24914,N_24669);
nor UO_1275 (O_1275,N_24484,N_24848);
or UO_1276 (O_1276,N_24998,N_24054);
nand UO_1277 (O_1277,N_24733,N_24216);
nor UO_1278 (O_1278,N_24699,N_24217);
and UO_1279 (O_1279,N_24104,N_24958);
or UO_1280 (O_1280,N_24332,N_24814);
or UO_1281 (O_1281,N_24293,N_24448);
nor UO_1282 (O_1282,N_24773,N_24156);
nand UO_1283 (O_1283,N_24685,N_24484);
xor UO_1284 (O_1284,N_24582,N_24817);
or UO_1285 (O_1285,N_24234,N_24067);
nand UO_1286 (O_1286,N_24144,N_24175);
nand UO_1287 (O_1287,N_24900,N_24783);
or UO_1288 (O_1288,N_24801,N_24522);
xor UO_1289 (O_1289,N_24107,N_24480);
nand UO_1290 (O_1290,N_24788,N_24688);
or UO_1291 (O_1291,N_24608,N_24560);
nand UO_1292 (O_1292,N_24922,N_24978);
and UO_1293 (O_1293,N_24738,N_24177);
and UO_1294 (O_1294,N_24849,N_24163);
nor UO_1295 (O_1295,N_24722,N_24651);
or UO_1296 (O_1296,N_24569,N_24982);
nand UO_1297 (O_1297,N_24076,N_24408);
nand UO_1298 (O_1298,N_24036,N_24316);
nand UO_1299 (O_1299,N_24059,N_24571);
xnor UO_1300 (O_1300,N_24878,N_24893);
or UO_1301 (O_1301,N_24792,N_24045);
or UO_1302 (O_1302,N_24048,N_24974);
xor UO_1303 (O_1303,N_24580,N_24812);
nor UO_1304 (O_1304,N_24249,N_24894);
and UO_1305 (O_1305,N_24216,N_24677);
or UO_1306 (O_1306,N_24746,N_24302);
nor UO_1307 (O_1307,N_24018,N_24578);
nand UO_1308 (O_1308,N_24111,N_24622);
xnor UO_1309 (O_1309,N_24167,N_24291);
nor UO_1310 (O_1310,N_24179,N_24061);
or UO_1311 (O_1311,N_24324,N_24960);
and UO_1312 (O_1312,N_24866,N_24067);
nor UO_1313 (O_1313,N_24719,N_24519);
nand UO_1314 (O_1314,N_24153,N_24920);
xnor UO_1315 (O_1315,N_24883,N_24780);
and UO_1316 (O_1316,N_24842,N_24090);
or UO_1317 (O_1317,N_24767,N_24043);
xnor UO_1318 (O_1318,N_24084,N_24362);
and UO_1319 (O_1319,N_24411,N_24625);
xnor UO_1320 (O_1320,N_24347,N_24441);
nand UO_1321 (O_1321,N_24716,N_24946);
nand UO_1322 (O_1322,N_24965,N_24919);
or UO_1323 (O_1323,N_24707,N_24906);
xor UO_1324 (O_1324,N_24342,N_24868);
xor UO_1325 (O_1325,N_24731,N_24773);
and UO_1326 (O_1326,N_24683,N_24588);
xnor UO_1327 (O_1327,N_24190,N_24683);
or UO_1328 (O_1328,N_24515,N_24213);
nand UO_1329 (O_1329,N_24041,N_24621);
xor UO_1330 (O_1330,N_24036,N_24002);
xnor UO_1331 (O_1331,N_24230,N_24872);
or UO_1332 (O_1332,N_24413,N_24750);
xnor UO_1333 (O_1333,N_24867,N_24919);
nand UO_1334 (O_1334,N_24034,N_24849);
nor UO_1335 (O_1335,N_24815,N_24657);
xor UO_1336 (O_1336,N_24948,N_24911);
nor UO_1337 (O_1337,N_24273,N_24558);
or UO_1338 (O_1338,N_24151,N_24493);
or UO_1339 (O_1339,N_24172,N_24206);
and UO_1340 (O_1340,N_24394,N_24315);
nand UO_1341 (O_1341,N_24844,N_24306);
nand UO_1342 (O_1342,N_24357,N_24486);
nor UO_1343 (O_1343,N_24925,N_24209);
and UO_1344 (O_1344,N_24412,N_24844);
xor UO_1345 (O_1345,N_24594,N_24282);
or UO_1346 (O_1346,N_24384,N_24118);
and UO_1347 (O_1347,N_24591,N_24454);
nand UO_1348 (O_1348,N_24781,N_24114);
or UO_1349 (O_1349,N_24398,N_24516);
xnor UO_1350 (O_1350,N_24944,N_24441);
and UO_1351 (O_1351,N_24593,N_24609);
xnor UO_1352 (O_1352,N_24093,N_24293);
and UO_1353 (O_1353,N_24049,N_24307);
and UO_1354 (O_1354,N_24986,N_24038);
nand UO_1355 (O_1355,N_24662,N_24035);
xor UO_1356 (O_1356,N_24500,N_24573);
or UO_1357 (O_1357,N_24188,N_24523);
and UO_1358 (O_1358,N_24511,N_24037);
and UO_1359 (O_1359,N_24656,N_24216);
or UO_1360 (O_1360,N_24202,N_24275);
xnor UO_1361 (O_1361,N_24560,N_24177);
nand UO_1362 (O_1362,N_24731,N_24566);
xor UO_1363 (O_1363,N_24124,N_24028);
and UO_1364 (O_1364,N_24492,N_24000);
nand UO_1365 (O_1365,N_24904,N_24217);
xnor UO_1366 (O_1366,N_24170,N_24235);
nor UO_1367 (O_1367,N_24819,N_24457);
nand UO_1368 (O_1368,N_24621,N_24931);
nand UO_1369 (O_1369,N_24454,N_24457);
nor UO_1370 (O_1370,N_24240,N_24470);
or UO_1371 (O_1371,N_24172,N_24823);
and UO_1372 (O_1372,N_24470,N_24048);
and UO_1373 (O_1373,N_24968,N_24353);
nor UO_1374 (O_1374,N_24397,N_24871);
nor UO_1375 (O_1375,N_24865,N_24754);
or UO_1376 (O_1376,N_24267,N_24395);
and UO_1377 (O_1377,N_24665,N_24631);
or UO_1378 (O_1378,N_24672,N_24400);
xnor UO_1379 (O_1379,N_24548,N_24558);
xor UO_1380 (O_1380,N_24627,N_24335);
xor UO_1381 (O_1381,N_24138,N_24252);
or UO_1382 (O_1382,N_24625,N_24644);
and UO_1383 (O_1383,N_24321,N_24675);
xor UO_1384 (O_1384,N_24482,N_24410);
or UO_1385 (O_1385,N_24177,N_24422);
nand UO_1386 (O_1386,N_24565,N_24891);
nor UO_1387 (O_1387,N_24420,N_24294);
xor UO_1388 (O_1388,N_24988,N_24029);
nand UO_1389 (O_1389,N_24762,N_24370);
nor UO_1390 (O_1390,N_24966,N_24095);
and UO_1391 (O_1391,N_24307,N_24580);
xor UO_1392 (O_1392,N_24303,N_24558);
nor UO_1393 (O_1393,N_24852,N_24960);
and UO_1394 (O_1394,N_24919,N_24606);
and UO_1395 (O_1395,N_24785,N_24216);
and UO_1396 (O_1396,N_24628,N_24466);
and UO_1397 (O_1397,N_24332,N_24067);
nand UO_1398 (O_1398,N_24369,N_24955);
nor UO_1399 (O_1399,N_24745,N_24108);
xor UO_1400 (O_1400,N_24143,N_24587);
xnor UO_1401 (O_1401,N_24763,N_24778);
nand UO_1402 (O_1402,N_24514,N_24589);
nand UO_1403 (O_1403,N_24729,N_24792);
nor UO_1404 (O_1404,N_24815,N_24661);
and UO_1405 (O_1405,N_24439,N_24065);
xnor UO_1406 (O_1406,N_24627,N_24574);
and UO_1407 (O_1407,N_24370,N_24358);
nand UO_1408 (O_1408,N_24815,N_24543);
nand UO_1409 (O_1409,N_24431,N_24642);
xnor UO_1410 (O_1410,N_24498,N_24278);
or UO_1411 (O_1411,N_24901,N_24203);
nor UO_1412 (O_1412,N_24175,N_24250);
or UO_1413 (O_1413,N_24962,N_24548);
or UO_1414 (O_1414,N_24539,N_24798);
xor UO_1415 (O_1415,N_24679,N_24449);
and UO_1416 (O_1416,N_24150,N_24562);
or UO_1417 (O_1417,N_24039,N_24855);
xnor UO_1418 (O_1418,N_24484,N_24241);
or UO_1419 (O_1419,N_24848,N_24067);
or UO_1420 (O_1420,N_24015,N_24334);
xnor UO_1421 (O_1421,N_24029,N_24587);
nor UO_1422 (O_1422,N_24185,N_24128);
nand UO_1423 (O_1423,N_24769,N_24947);
and UO_1424 (O_1424,N_24087,N_24739);
and UO_1425 (O_1425,N_24158,N_24273);
or UO_1426 (O_1426,N_24750,N_24695);
xnor UO_1427 (O_1427,N_24136,N_24403);
xnor UO_1428 (O_1428,N_24198,N_24874);
xnor UO_1429 (O_1429,N_24850,N_24904);
or UO_1430 (O_1430,N_24220,N_24335);
xnor UO_1431 (O_1431,N_24780,N_24156);
and UO_1432 (O_1432,N_24330,N_24814);
nor UO_1433 (O_1433,N_24563,N_24807);
xnor UO_1434 (O_1434,N_24959,N_24902);
or UO_1435 (O_1435,N_24864,N_24395);
xor UO_1436 (O_1436,N_24997,N_24061);
and UO_1437 (O_1437,N_24352,N_24302);
xnor UO_1438 (O_1438,N_24770,N_24840);
nor UO_1439 (O_1439,N_24652,N_24507);
nand UO_1440 (O_1440,N_24648,N_24862);
xor UO_1441 (O_1441,N_24320,N_24130);
nor UO_1442 (O_1442,N_24763,N_24620);
or UO_1443 (O_1443,N_24433,N_24861);
and UO_1444 (O_1444,N_24932,N_24942);
nand UO_1445 (O_1445,N_24459,N_24171);
nand UO_1446 (O_1446,N_24202,N_24964);
nor UO_1447 (O_1447,N_24255,N_24351);
xnor UO_1448 (O_1448,N_24507,N_24342);
xnor UO_1449 (O_1449,N_24874,N_24748);
nor UO_1450 (O_1450,N_24918,N_24322);
and UO_1451 (O_1451,N_24633,N_24163);
xnor UO_1452 (O_1452,N_24242,N_24622);
nand UO_1453 (O_1453,N_24567,N_24636);
nor UO_1454 (O_1454,N_24957,N_24653);
or UO_1455 (O_1455,N_24012,N_24487);
nand UO_1456 (O_1456,N_24563,N_24156);
or UO_1457 (O_1457,N_24504,N_24402);
and UO_1458 (O_1458,N_24793,N_24755);
xor UO_1459 (O_1459,N_24629,N_24823);
and UO_1460 (O_1460,N_24885,N_24701);
nor UO_1461 (O_1461,N_24084,N_24697);
or UO_1462 (O_1462,N_24824,N_24436);
nand UO_1463 (O_1463,N_24836,N_24646);
xor UO_1464 (O_1464,N_24120,N_24123);
nand UO_1465 (O_1465,N_24901,N_24404);
nand UO_1466 (O_1466,N_24688,N_24530);
xnor UO_1467 (O_1467,N_24018,N_24806);
nand UO_1468 (O_1468,N_24817,N_24112);
nand UO_1469 (O_1469,N_24022,N_24551);
nor UO_1470 (O_1470,N_24812,N_24136);
xnor UO_1471 (O_1471,N_24660,N_24090);
nand UO_1472 (O_1472,N_24728,N_24862);
nand UO_1473 (O_1473,N_24947,N_24119);
nor UO_1474 (O_1474,N_24253,N_24755);
nor UO_1475 (O_1475,N_24153,N_24144);
nor UO_1476 (O_1476,N_24857,N_24162);
nor UO_1477 (O_1477,N_24401,N_24860);
nor UO_1478 (O_1478,N_24514,N_24876);
or UO_1479 (O_1479,N_24634,N_24917);
and UO_1480 (O_1480,N_24023,N_24583);
or UO_1481 (O_1481,N_24284,N_24955);
nand UO_1482 (O_1482,N_24642,N_24556);
xnor UO_1483 (O_1483,N_24721,N_24367);
or UO_1484 (O_1484,N_24547,N_24749);
xor UO_1485 (O_1485,N_24914,N_24364);
nand UO_1486 (O_1486,N_24805,N_24608);
and UO_1487 (O_1487,N_24394,N_24301);
nand UO_1488 (O_1488,N_24265,N_24292);
nand UO_1489 (O_1489,N_24804,N_24683);
or UO_1490 (O_1490,N_24256,N_24913);
nor UO_1491 (O_1491,N_24221,N_24280);
nand UO_1492 (O_1492,N_24047,N_24232);
or UO_1493 (O_1493,N_24689,N_24031);
nand UO_1494 (O_1494,N_24159,N_24075);
xnor UO_1495 (O_1495,N_24465,N_24394);
nand UO_1496 (O_1496,N_24532,N_24515);
xnor UO_1497 (O_1497,N_24538,N_24773);
and UO_1498 (O_1498,N_24140,N_24573);
xor UO_1499 (O_1499,N_24509,N_24668);
nand UO_1500 (O_1500,N_24046,N_24301);
nor UO_1501 (O_1501,N_24553,N_24654);
or UO_1502 (O_1502,N_24752,N_24727);
or UO_1503 (O_1503,N_24466,N_24652);
or UO_1504 (O_1504,N_24368,N_24794);
xnor UO_1505 (O_1505,N_24429,N_24757);
nand UO_1506 (O_1506,N_24255,N_24124);
and UO_1507 (O_1507,N_24663,N_24440);
xnor UO_1508 (O_1508,N_24761,N_24054);
xnor UO_1509 (O_1509,N_24309,N_24125);
or UO_1510 (O_1510,N_24124,N_24681);
and UO_1511 (O_1511,N_24561,N_24238);
nor UO_1512 (O_1512,N_24627,N_24546);
nor UO_1513 (O_1513,N_24309,N_24531);
nor UO_1514 (O_1514,N_24945,N_24004);
and UO_1515 (O_1515,N_24736,N_24065);
nor UO_1516 (O_1516,N_24662,N_24389);
nand UO_1517 (O_1517,N_24839,N_24026);
or UO_1518 (O_1518,N_24693,N_24119);
nand UO_1519 (O_1519,N_24519,N_24875);
xor UO_1520 (O_1520,N_24768,N_24633);
xor UO_1521 (O_1521,N_24861,N_24120);
and UO_1522 (O_1522,N_24833,N_24882);
nor UO_1523 (O_1523,N_24622,N_24135);
nand UO_1524 (O_1524,N_24492,N_24375);
nor UO_1525 (O_1525,N_24605,N_24456);
nor UO_1526 (O_1526,N_24899,N_24044);
nor UO_1527 (O_1527,N_24412,N_24953);
xnor UO_1528 (O_1528,N_24122,N_24474);
xnor UO_1529 (O_1529,N_24408,N_24862);
and UO_1530 (O_1530,N_24622,N_24401);
and UO_1531 (O_1531,N_24436,N_24173);
or UO_1532 (O_1532,N_24783,N_24619);
xnor UO_1533 (O_1533,N_24256,N_24156);
and UO_1534 (O_1534,N_24543,N_24822);
and UO_1535 (O_1535,N_24644,N_24780);
nand UO_1536 (O_1536,N_24892,N_24665);
nor UO_1537 (O_1537,N_24310,N_24125);
nor UO_1538 (O_1538,N_24808,N_24335);
and UO_1539 (O_1539,N_24691,N_24452);
xor UO_1540 (O_1540,N_24960,N_24856);
and UO_1541 (O_1541,N_24864,N_24453);
xor UO_1542 (O_1542,N_24107,N_24738);
and UO_1543 (O_1543,N_24063,N_24318);
and UO_1544 (O_1544,N_24482,N_24131);
or UO_1545 (O_1545,N_24153,N_24502);
or UO_1546 (O_1546,N_24561,N_24417);
or UO_1547 (O_1547,N_24483,N_24419);
and UO_1548 (O_1548,N_24956,N_24363);
nor UO_1549 (O_1549,N_24544,N_24687);
or UO_1550 (O_1550,N_24460,N_24566);
nor UO_1551 (O_1551,N_24924,N_24494);
and UO_1552 (O_1552,N_24984,N_24364);
nand UO_1553 (O_1553,N_24760,N_24943);
xnor UO_1554 (O_1554,N_24943,N_24210);
nor UO_1555 (O_1555,N_24439,N_24081);
nand UO_1556 (O_1556,N_24779,N_24518);
xnor UO_1557 (O_1557,N_24036,N_24702);
or UO_1558 (O_1558,N_24290,N_24509);
or UO_1559 (O_1559,N_24900,N_24162);
or UO_1560 (O_1560,N_24839,N_24377);
nand UO_1561 (O_1561,N_24292,N_24258);
or UO_1562 (O_1562,N_24757,N_24130);
or UO_1563 (O_1563,N_24980,N_24592);
or UO_1564 (O_1564,N_24692,N_24392);
xnor UO_1565 (O_1565,N_24923,N_24311);
nand UO_1566 (O_1566,N_24703,N_24951);
and UO_1567 (O_1567,N_24945,N_24322);
and UO_1568 (O_1568,N_24218,N_24015);
nand UO_1569 (O_1569,N_24757,N_24789);
and UO_1570 (O_1570,N_24505,N_24436);
and UO_1571 (O_1571,N_24020,N_24769);
xnor UO_1572 (O_1572,N_24059,N_24273);
or UO_1573 (O_1573,N_24732,N_24539);
nor UO_1574 (O_1574,N_24732,N_24467);
xnor UO_1575 (O_1575,N_24784,N_24783);
nand UO_1576 (O_1576,N_24867,N_24326);
nor UO_1577 (O_1577,N_24108,N_24683);
nand UO_1578 (O_1578,N_24858,N_24554);
nor UO_1579 (O_1579,N_24308,N_24778);
xor UO_1580 (O_1580,N_24040,N_24002);
xor UO_1581 (O_1581,N_24751,N_24974);
or UO_1582 (O_1582,N_24548,N_24034);
nor UO_1583 (O_1583,N_24248,N_24361);
xnor UO_1584 (O_1584,N_24864,N_24675);
nor UO_1585 (O_1585,N_24767,N_24117);
or UO_1586 (O_1586,N_24747,N_24318);
nand UO_1587 (O_1587,N_24112,N_24363);
nor UO_1588 (O_1588,N_24471,N_24746);
xor UO_1589 (O_1589,N_24988,N_24360);
and UO_1590 (O_1590,N_24508,N_24562);
and UO_1591 (O_1591,N_24618,N_24871);
nand UO_1592 (O_1592,N_24130,N_24768);
nand UO_1593 (O_1593,N_24377,N_24754);
xnor UO_1594 (O_1594,N_24745,N_24867);
xor UO_1595 (O_1595,N_24068,N_24176);
xor UO_1596 (O_1596,N_24041,N_24793);
or UO_1597 (O_1597,N_24476,N_24822);
and UO_1598 (O_1598,N_24432,N_24080);
nand UO_1599 (O_1599,N_24381,N_24864);
nor UO_1600 (O_1600,N_24931,N_24450);
xor UO_1601 (O_1601,N_24355,N_24174);
or UO_1602 (O_1602,N_24871,N_24310);
and UO_1603 (O_1603,N_24330,N_24361);
nor UO_1604 (O_1604,N_24196,N_24488);
or UO_1605 (O_1605,N_24656,N_24725);
or UO_1606 (O_1606,N_24166,N_24485);
and UO_1607 (O_1607,N_24958,N_24396);
or UO_1608 (O_1608,N_24869,N_24986);
or UO_1609 (O_1609,N_24515,N_24651);
nor UO_1610 (O_1610,N_24513,N_24271);
nor UO_1611 (O_1611,N_24017,N_24209);
xor UO_1612 (O_1612,N_24338,N_24380);
xor UO_1613 (O_1613,N_24374,N_24880);
xnor UO_1614 (O_1614,N_24768,N_24756);
nor UO_1615 (O_1615,N_24766,N_24232);
or UO_1616 (O_1616,N_24109,N_24102);
and UO_1617 (O_1617,N_24349,N_24831);
nand UO_1618 (O_1618,N_24427,N_24170);
nor UO_1619 (O_1619,N_24295,N_24577);
and UO_1620 (O_1620,N_24415,N_24437);
nor UO_1621 (O_1621,N_24822,N_24854);
and UO_1622 (O_1622,N_24591,N_24193);
xor UO_1623 (O_1623,N_24711,N_24076);
and UO_1624 (O_1624,N_24952,N_24857);
or UO_1625 (O_1625,N_24581,N_24039);
xnor UO_1626 (O_1626,N_24509,N_24995);
nand UO_1627 (O_1627,N_24690,N_24130);
or UO_1628 (O_1628,N_24925,N_24966);
nor UO_1629 (O_1629,N_24499,N_24820);
nor UO_1630 (O_1630,N_24097,N_24603);
nor UO_1631 (O_1631,N_24732,N_24567);
and UO_1632 (O_1632,N_24225,N_24313);
nor UO_1633 (O_1633,N_24072,N_24995);
nor UO_1634 (O_1634,N_24625,N_24216);
xor UO_1635 (O_1635,N_24384,N_24742);
xnor UO_1636 (O_1636,N_24696,N_24068);
or UO_1637 (O_1637,N_24680,N_24726);
nor UO_1638 (O_1638,N_24775,N_24070);
or UO_1639 (O_1639,N_24027,N_24427);
nand UO_1640 (O_1640,N_24955,N_24275);
or UO_1641 (O_1641,N_24279,N_24604);
nor UO_1642 (O_1642,N_24351,N_24799);
xnor UO_1643 (O_1643,N_24106,N_24320);
nand UO_1644 (O_1644,N_24838,N_24032);
xnor UO_1645 (O_1645,N_24333,N_24032);
or UO_1646 (O_1646,N_24116,N_24411);
nor UO_1647 (O_1647,N_24575,N_24678);
xor UO_1648 (O_1648,N_24135,N_24169);
and UO_1649 (O_1649,N_24895,N_24683);
nor UO_1650 (O_1650,N_24080,N_24542);
or UO_1651 (O_1651,N_24460,N_24860);
xnor UO_1652 (O_1652,N_24725,N_24697);
xnor UO_1653 (O_1653,N_24588,N_24532);
or UO_1654 (O_1654,N_24891,N_24685);
or UO_1655 (O_1655,N_24862,N_24525);
nand UO_1656 (O_1656,N_24374,N_24338);
and UO_1657 (O_1657,N_24264,N_24889);
nand UO_1658 (O_1658,N_24635,N_24571);
and UO_1659 (O_1659,N_24565,N_24748);
and UO_1660 (O_1660,N_24470,N_24870);
nor UO_1661 (O_1661,N_24244,N_24821);
nand UO_1662 (O_1662,N_24313,N_24503);
or UO_1663 (O_1663,N_24715,N_24250);
nor UO_1664 (O_1664,N_24568,N_24087);
nand UO_1665 (O_1665,N_24663,N_24169);
nor UO_1666 (O_1666,N_24363,N_24003);
xnor UO_1667 (O_1667,N_24335,N_24886);
xnor UO_1668 (O_1668,N_24448,N_24856);
nand UO_1669 (O_1669,N_24585,N_24276);
nor UO_1670 (O_1670,N_24177,N_24159);
or UO_1671 (O_1671,N_24023,N_24774);
nand UO_1672 (O_1672,N_24379,N_24094);
nand UO_1673 (O_1673,N_24188,N_24348);
or UO_1674 (O_1674,N_24008,N_24880);
nor UO_1675 (O_1675,N_24103,N_24367);
nor UO_1676 (O_1676,N_24136,N_24486);
nand UO_1677 (O_1677,N_24185,N_24987);
nor UO_1678 (O_1678,N_24749,N_24284);
or UO_1679 (O_1679,N_24732,N_24379);
nor UO_1680 (O_1680,N_24978,N_24480);
xnor UO_1681 (O_1681,N_24830,N_24139);
nor UO_1682 (O_1682,N_24893,N_24440);
nor UO_1683 (O_1683,N_24031,N_24759);
or UO_1684 (O_1684,N_24010,N_24333);
and UO_1685 (O_1685,N_24039,N_24905);
xor UO_1686 (O_1686,N_24338,N_24671);
xor UO_1687 (O_1687,N_24488,N_24711);
nor UO_1688 (O_1688,N_24282,N_24747);
nand UO_1689 (O_1689,N_24475,N_24030);
and UO_1690 (O_1690,N_24316,N_24211);
nor UO_1691 (O_1691,N_24569,N_24958);
nand UO_1692 (O_1692,N_24748,N_24080);
xor UO_1693 (O_1693,N_24803,N_24357);
or UO_1694 (O_1694,N_24467,N_24949);
or UO_1695 (O_1695,N_24837,N_24498);
nand UO_1696 (O_1696,N_24985,N_24671);
nor UO_1697 (O_1697,N_24629,N_24292);
or UO_1698 (O_1698,N_24749,N_24353);
or UO_1699 (O_1699,N_24922,N_24924);
xnor UO_1700 (O_1700,N_24699,N_24638);
xnor UO_1701 (O_1701,N_24104,N_24625);
xor UO_1702 (O_1702,N_24282,N_24550);
or UO_1703 (O_1703,N_24967,N_24277);
xnor UO_1704 (O_1704,N_24425,N_24737);
nand UO_1705 (O_1705,N_24288,N_24910);
nor UO_1706 (O_1706,N_24862,N_24673);
xnor UO_1707 (O_1707,N_24534,N_24188);
nand UO_1708 (O_1708,N_24161,N_24124);
xnor UO_1709 (O_1709,N_24858,N_24482);
nand UO_1710 (O_1710,N_24202,N_24394);
and UO_1711 (O_1711,N_24118,N_24646);
nor UO_1712 (O_1712,N_24567,N_24589);
and UO_1713 (O_1713,N_24597,N_24504);
nand UO_1714 (O_1714,N_24947,N_24737);
nand UO_1715 (O_1715,N_24136,N_24453);
xnor UO_1716 (O_1716,N_24096,N_24565);
xnor UO_1717 (O_1717,N_24532,N_24391);
or UO_1718 (O_1718,N_24099,N_24695);
xor UO_1719 (O_1719,N_24466,N_24066);
nor UO_1720 (O_1720,N_24489,N_24996);
and UO_1721 (O_1721,N_24267,N_24579);
nor UO_1722 (O_1722,N_24045,N_24190);
and UO_1723 (O_1723,N_24982,N_24125);
xor UO_1724 (O_1724,N_24919,N_24163);
or UO_1725 (O_1725,N_24881,N_24033);
nand UO_1726 (O_1726,N_24000,N_24723);
or UO_1727 (O_1727,N_24392,N_24564);
xnor UO_1728 (O_1728,N_24515,N_24869);
or UO_1729 (O_1729,N_24052,N_24014);
nor UO_1730 (O_1730,N_24950,N_24538);
nor UO_1731 (O_1731,N_24882,N_24422);
and UO_1732 (O_1732,N_24779,N_24239);
nand UO_1733 (O_1733,N_24396,N_24870);
and UO_1734 (O_1734,N_24766,N_24806);
nor UO_1735 (O_1735,N_24350,N_24335);
nor UO_1736 (O_1736,N_24377,N_24647);
nor UO_1737 (O_1737,N_24337,N_24124);
and UO_1738 (O_1738,N_24170,N_24198);
and UO_1739 (O_1739,N_24762,N_24487);
xnor UO_1740 (O_1740,N_24781,N_24256);
nor UO_1741 (O_1741,N_24205,N_24798);
nand UO_1742 (O_1742,N_24888,N_24048);
xor UO_1743 (O_1743,N_24241,N_24842);
and UO_1744 (O_1744,N_24648,N_24186);
xor UO_1745 (O_1745,N_24465,N_24395);
or UO_1746 (O_1746,N_24613,N_24172);
xor UO_1747 (O_1747,N_24604,N_24999);
nor UO_1748 (O_1748,N_24706,N_24352);
nand UO_1749 (O_1749,N_24929,N_24805);
and UO_1750 (O_1750,N_24253,N_24269);
xor UO_1751 (O_1751,N_24747,N_24586);
or UO_1752 (O_1752,N_24833,N_24892);
and UO_1753 (O_1753,N_24887,N_24652);
nor UO_1754 (O_1754,N_24809,N_24921);
or UO_1755 (O_1755,N_24525,N_24796);
nor UO_1756 (O_1756,N_24897,N_24733);
or UO_1757 (O_1757,N_24928,N_24640);
or UO_1758 (O_1758,N_24386,N_24538);
or UO_1759 (O_1759,N_24380,N_24951);
nor UO_1760 (O_1760,N_24551,N_24617);
or UO_1761 (O_1761,N_24000,N_24162);
nand UO_1762 (O_1762,N_24115,N_24669);
nand UO_1763 (O_1763,N_24119,N_24641);
nor UO_1764 (O_1764,N_24998,N_24696);
nor UO_1765 (O_1765,N_24830,N_24157);
or UO_1766 (O_1766,N_24239,N_24068);
or UO_1767 (O_1767,N_24159,N_24540);
and UO_1768 (O_1768,N_24646,N_24026);
nor UO_1769 (O_1769,N_24176,N_24103);
xor UO_1770 (O_1770,N_24102,N_24098);
and UO_1771 (O_1771,N_24942,N_24944);
and UO_1772 (O_1772,N_24813,N_24668);
xnor UO_1773 (O_1773,N_24013,N_24669);
and UO_1774 (O_1774,N_24176,N_24804);
or UO_1775 (O_1775,N_24048,N_24933);
nor UO_1776 (O_1776,N_24297,N_24065);
or UO_1777 (O_1777,N_24046,N_24698);
xnor UO_1778 (O_1778,N_24543,N_24942);
nand UO_1779 (O_1779,N_24114,N_24084);
nor UO_1780 (O_1780,N_24827,N_24416);
or UO_1781 (O_1781,N_24831,N_24817);
nor UO_1782 (O_1782,N_24346,N_24642);
nand UO_1783 (O_1783,N_24202,N_24732);
nor UO_1784 (O_1784,N_24103,N_24720);
and UO_1785 (O_1785,N_24044,N_24448);
and UO_1786 (O_1786,N_24492,N_24771);
xnor UO_1787 (O_1787,N_24703,N_24984);
or UO_1788 (O_1788,N_24013,N_24055);
xnor UO_1789 (O_1789,N_24626,N_24540);
nand UO_1790 (O_1790,N_24755,N_24681);
xnor UO_1791 (O_1791,N_24755,N_24463);
nand UO_1792 (O_1792,N_24457,N_24635);
nor UO_1793 (O_1793,N_24840,N_24457);
nor UO_1794 (O_1794,N_24378,N_24567);
nand UO_1795 (O_1795,N_24411,N_24626);
xnor UO_1796 (O_1796,N_24741,N_24250);
xnor UO_1797 (O_1797,N_24708,N_24387);
nor UO_1798 (O_1798,N_24674,N_24286);
and UO_1799 (O_1799,N_24979,N_24980);
nor UO_1800 (O_1800,N_24459,N_24666);
and UO_1801 (O_1801,N_24177,N_24346);
nand UO_1802 (O_1802,N_24008,N_24011);
or UO_1803 (O_1803,N_24829,N_24713);
xor UO_1804 (O_1804,N_24922,N_24250);
nand UO_1805 (O_1805,N_24867,N_24236);
or UO_1806 (O_1806,N_24893,N_24663);
xnor UO_1807 (O_1807,N_24555,N_24812);
nand UO_1808 (O_1808,N_24594,N_24688);
nand UO_1809 (O_1809,N_24685,N_24644);
or UO_1810 (O_1810,N_24570,N_24412);
nand UO_1811 (O_1811,N_24367,N_24620);
or UO_1812 (O_1812,N_24184,N_24539);
nor UO_1813 (O_1813,N_24117,N_24035);
nor UO_1814 (O_1814,N_24047,N_24177);
and UO_1815 (O_1815,N_24333,N_24459);
xor UO_1816 (O_1816,N_24549,N_24525);
nand UO_1817 (O_1817,N_24229,N_24426);
and UO_1818 (O_1818,N_24973,N_24616);
and UO_1819 (O_1819,N_24761,N_24149);
and UO_1820 (O_1820,N_24385,N_24241);
nor UO_1821 (O_1821,N_24434,N_24492);
nand UO_1822 (O_1822,N_24476,N_24792);
and UO_1823 (O_1823,N_24865,N_24417);
nor UO_1824 (O_1824,N_24728,N_24791);
or UO_1825 (O_1825,N_24797,N_24845);
and UO_1826 (O_1826,N_24391,N_24673);
nor UO_1827 (O_1827,N_24996,N_24318);
nand UO_1828 (O_1828,N_24082,N_24770);
nor UO_1829 (O_1829,N_24798,N_24568);
and UO_1830 (O_1830,N_24872,N_24601);
nor UO_1831 (O_1831,N_24770,N_24526);
nor UO_1832 (O_1832,N_24870,N_24080);
or UO_1833 (O_1833,N_24250,N_24733);
or UO_1834 (O_1834,N_24488,N_24670);
or UO_1835 (O_1835,N_24388,N_24768);
and UO_1836 (O_1836,N_24458,N_24487);
or UO_1837 (O_1837,N_24329,N_24790);
or UO_1838 (O_1838,N_24524,N_24633);
nor UO_1839 (O_1839,N_24291,N_24325);
nor UO_1840 (O_1840,N_24627,N_24519);
nand UO_1841 (O_1841,N_24871,N_24677);
xor UO_1842 (O_1842,N_24841,N_24994);
xor UO_1843 (O_1843,N_24572,N_24295);
and UO_1844 (O_1844,N_24785,N_24310);
nand UO_1845 (O_1845,N_24712,N_24387);
xor UO_1846 (O_1846,N_24374,N_24442);
or UO_1847 (O_1847,N_24551,N_24392);
xnor UO_1848 (O_1848,N_24469,N_24979);
nor UO_1849 (O_1849,N_24823,N_24729);
or UO_1850 (O_1850,N_24002,N_24299);
and UO_1851 (O_1851,N_24218,N_24450);
nand UO_1852 (O_1852,N_24141,N_24777);
xor UO_1853 (O_1853,N_24724,N_24375);
and UO_1854 (O_1854,N_24150,N_24302);
or UO_1855 (O_1855,N_24644,N_24699);
and UO_1856 (O_1856,N_24611,N_24546);
nor UO_1857 (O_1857,N_24603,N_24302);
xor UO_1858 (O_1858,N_24332,N_24478);
or UO_1859 (O_1859,N_24180,N_24000);
nor UO_1860 (O_1860,N_24970,N_24087);
xor UO_1861 (O_1861,N_24632,N_24157);
nand UO_1862 (O_1862,N_24849,N_24355);
nor UO_1863 (O_1863,N_24108,N_24600);
and UO_1864 (O_1864,N_24720,N_24245);
or UO_1865 (O_1865,N_24984,N_24777);
or UO_1866 (O_1866,N_24592,N_24418);
xnor UO_1867 (O_1867,N_24393,N_24492);
nor UO_1868 (O_1868,N_24169,N_24868);
nand UO_1869 (O_1869,N_24750,N_24157);
nand UO_1870 (O_1870,N_24610,N_24196);
nor UO_1871 (O_1871,N_24135,N_24293);
or UO_1872 (O_1872,N_24876,N_24493);
xor UO_1873 (O_1873,N_24306,N_24155);
nor UO_1874 (O_1874,N_24913,N_24367);
nor UO_1875 (O_1875,N_24880,N_24277);
and UO_1876 (O_1876,N_24304,N_24604);
and UO_1877 (O_1877,N_24086,N_24673);
nor UO_1878 (O_1878,N_24779,N_24022);
xor UO_1879 (O_1879,N_24070,N_24742);
or UO_1880 (O_1880,N_24055,N_24363);
xnor UO_1881 (O_1881,N_24041,N_24179);
or UO_1882 (O_1882,N_24213,N_24944);
or UO_1883 (O_1883,N_24859,N_24350);
and UO_1884 (O_1884,N_24027,N_24058);
nor UO_1885 (O_1885,N_24092,N_24229);
nor UO_1886 (O_1886,N_24037,N_24689);
nand UO_1887 (O_1887,N_24064,N_24874);
xor UO_1888 (O_1888,N_24202,N_24997);
or UO_1889 (O_1889,N_24648,N_24501);
nor UO_1890 (O_1890,N_24025,N_24569);
and UO_1891 (O_1891,N_24538,N_24891);
nor UO_1892 (O_1892,N_24843,N_24367);
xnor UO_1893 (O_1893,N_24352,N_24140);
xor UO_1894 (O_1894,N_24641,N_24148);
or UO_1895 (O_1895,N_24125,N_24324);
and UO_1896 (O_1896,N_24788,N_24192);
or UO_1897 (O_1897,N_24115,N_24473);
and UO_1898 (O_1898,N_24350,N_24439);
nor UO_1899 (O_1899,N_24164,N_24973);
or UO_1900 (O_1900,N_24880,N_24509);
xor UO_1901 (O_1901,N_24071,N_24436);
nor UO_1902 (O_1902,N_24457,N_24563);
nor UO_1903 (O_1903,N_24133,N_24985);
nor UO_1904 (O_1904,N_24089,N_24011);
nand UO_1905 (O_1905,N_24961,N_24672);
nand UO_1906 (O_1906,N_24620,N_24577);
nand UO_1907 (O_1907,N_24021,N_24391);
nor UO_1908 (O_1908,N_24594,N_24709);
and UO_1909 (O_1909,N_24086,N_24026);
or UO_1910 (O_1910,N_24747,N_24579);
nand UO_1911 (O_1911,N_24879,N_24014);
nand UO_1912 (O_1912,N_24495,N_24383);
nor UO_1913 (O_1913,N_24528,N_24343);
nor UO_1914 (O_1914,N_24270,N_24011);
xnor UO_1915 (O_1915,N_24174,N_24235);
and UO_1916 (O_1916,N_24905,N_24543);
xor UO_1917 (O_1917,N_24630,N_24178);
and UO_1918 (O_1918,N_24246,N_24258);
xnor UO_1919 (O_1919,N_24477,N_24189);
nand UO_1920 (O_1920,N_24024,N_24428);
xor UO_1921 (O_1921,N_24060,N_24719);
nand UO_1922 (O_1922,N_24859,N_24675);
nor UO_1923 (O_1923,N_24939,N_24462);
xnor UO_1924 (O_1924,N_24358,N_24486);
or UO_1925 (O_1925,N_24420,N_24074);
or UO_1926 (O_1926,N_24009,N_24659);
xnor UO_1927 (O_1927,N_24916,N_24102);
and UO_1928 (O_1928,N_24181,N_24836);
xnor UO_1929 (O_1929,N_24732,N_24558);
xnor UO_1930 (O_1930,N_24834,N_24185);
nor UO_1931 (O_1931,N_24858,N_24010);
nand UO_1932 (O_1932,N_24043,N_24371);
nor UO_1933 (O_1933,N_24245,N_24498);
nand UO_1934 (O_1934,N_24766,N_24631);
and UO_1935 (O_1935,N_24158,N_24394);
and UO_1936 (O_1936,N_24330,N_24247);
and UO_1937 (O_1937,N_24102,N_24053);
nor UO_1938 (O_1938,N_24890,N_24009);
nand UO_1939 (O_1939,N_24630,N_24820);
and UO_1940 (O_1940,N_24356,N_24615);
nand UO_1941 (O_1941,N_24266,N_24093);
xnor UO_1942 (O_1942,N_24555,N_24040);
and UO_1943 (O_1943,N_24393,N_24239);
xor UO_1944 (O_1944,N_24333,N_24762);
nor UO_1945 (O_1945,N_24156,N_24434);
or UO_1946 (O_1946,N_24582,N_24426);
xnor UO_1947 (O_1947,N_24176,N_24169);
nand UO_1948 (O_1948,N_24185,N_24385);
or UO_1949 (O_1949,N_24056,N_24415);
nor UO_1950 (O_1950,N_24382,N_24539);
or UO_1951 (O_1951,N_24799,N_24156);
or UO_1952 (O_1952,N_24976,N_24138);
nand UO_1953 (O_1953,N_24702,N_24847);
nand UO_1954 (O_1954,N_24485,N_24081);
nor UO_1955 (O_1955,N_24752,N_24307);
nor UO_1956 (O_1956,N_24537,N_24057);
nor UO_1957 (O_1957,N_24362,N_24951);
and UO_1958 (O_1958,N_24507,N_24537);
and UO_1959 (O_1959,N_24313,N_24232);
xnor UO_1960 (O_1960,N_24170,N_24166);
nor UO_1961 (O_1961,N_24022,N_24009);
nor UO_1962 (O_1962,N_24574,N_24003);
or UO_1963 (O_1963,N_24123,N_24811);
or UO_1964 (O_1964,N_24967,N_24799);
or UO_1965 (O_1965,N_24225,N_24348);
or UO_1966 (O_1966,N_24630,N_24093);
xor UO_1967 (O_1967,N_24044,N_24414);
nor UO_1968 (O_1968,N_24819,N_24666);
and UO_1969 (O_1969,N_24214,N_24659);
or UO_1970 (O_1970,N_24723,N_24874);
xor UO_1971 (O_1971,N_24783,N_24844);
nor UO_1972 (O_1972,N_24180,N_24877);
or UO_1973 (O_1973,N_24053,N_24095);
xnor UO_1974 (O_1974,N_24509,N_24477);
or UO_1975 (O_1975,N_24641,N_24015);
or UO_1976 (O_1976,N_24268,N_24171);
nand UO_1977 (O_1977,N_24511,N_24026);
and UO_1978 (O_1978,N_24429,N_24681);
or UO_1979 (O_1979,N_24236,N_24287);
xnor UO_1980 (O_1980,N_24509,N_24230);
and UO_1981 (O_1981,N_24461,N_24467);
or UO_1982 (O_1982,N_24677,N_24709);
nand UO_1983 (O_1983,N_24729,N_24960);
or UO_1984 (O_1984,N_24659,N_24698);
or UO_1985 (O_1985,N_24656,N_24129);
xor UO_1986 (O_1986,N_24854,N_24488);
nor UO_1987 (O_1987,N_24712,N_24662);
xor UO_1988 (O_1988,N_24601,N_24459);
xnor UO_1989 (O_1989,N_24583,N_24548);
and UO_1990 (O_1990,N_24557,N_24736);
nor UO_1991 (O_1991,N_24082,N_24986);
and UO_1992 (O_1992,N_24531,N_24011);
and UO_1993 (O_1993,N_24631,N_24187);
or UO_1994 (O_1994,N_24331,N_24517);
xor UO_1995 (O_1995,N_24172,N_24911);
or UO_1996 (O_1996,N_24640,N_24200);
xor UO_1997 (O_1997,N_24344,N_24058);
nor UO_1998 (O_1998,N_24452,N_24300);
or UO_1999 (O_1999,N_24651,N_24330);
or UO_2000 (O_2000,N_24381,N_24240);
nor UO_2001 (O_2001,N_24398,N_24918);
nor UO_2002 (O_2002,N_24148,N_24674);
or UO_2003 (O_2003,N_24340,N_24033);
xor UO_2004 (O_2004,N_24304,N_24407);
nor UO_2005 (O_2005,N_24108,N_24492);
and UO_2006 (O_2006,N_24936,N_24692);
and UO_2007 (O_2007,N_24288,N_24550);
and UO_2008 (O_2008,N_24704,N_24013);
nor UO_2009 (O_2009,N_24629,N_24281);
nand UO_2010 (O_2010,N_24295,N_24705);
xnor UO_2011 (O_2011,N_24334,N_24375);
and UO_2012 (O_2012,N_24303,N_24281);
or UO_2013 (O_2013,N_24114,N_24971);
xnor UO_2014 (O_2014,N_24243,N_24701);
nand UO_2015 (O_2015,N_24440,N_24715);
nand UO_2016 (O_2016,N_24677,N_24049);
and UO_2017 (O_2017,N_24896,N_24475);
or UO_2018 (O_2018,N_24460,N_24163);
xor UO_2019 (O_2019,N_24988,N_24650);
and UO_2020 (O_2020,N_24779,N_24819);
xnor UO_2021 (O_2021,N_24047,N_24609);
nor UO_2022 (O_2022,N_24985,N_24254);
xor UO_2023 (O_2023,N_24375,N_24509);
and UO_2024 (O_2024,N_24929,N_24005);
and UO_2025 (O_2025,N_24048,N_24330);
and UO_2026 (O_2026,N_24668,N_24218);
or UO_2027 (O_2027,N_24850,N_24867);
nand UO_2028 (O_2028,N_24245,N_24430);
or UO_2029 (O_2029,N_24939,N_24077);
nor UO_2030 (O_2030,N_24975,N_24582);
nand UO_2031 (O_2031,N_24370,N_24036);
xnor UO_2032 (O_2032,N_24043,N_24224);
or UO_2033 (O_2033,N_24555,N_24417);
xor UO_2034 (O_2034,N_24552,N_24992);
and UO_2035 (O_2035,N_24077,N_24674);
xor UO_2036 (O_2036,N_24514,N_24153);
nand UO_2037 (O_2037,N_24109,N_24531);
or UO_2038 (O_2038,N_24281,N_24459);
and UO_2039 (O_2039,N_24071,N_24302);
and UO_2040 (O_2040,N_24726,N_24081);
nor UO_2041 (O_2041,N_24675,N_24389);
nand UO_2042 (O_2042,N_24811,N_24582);
nor UO_2043 (O_2043,N_24878,N_24969);
xor UO_2044 (O_2044,N_24059,N_24507);
and UO_2045 (O_2045,N_24287,N_24506);
or UO_2046 (O_2046,N_24979,N_24472);
nor UO_2047 (O_2047,N_24466,N_24052);
xor UO_2048 (O_2048,N_24157,N_24011);
nor UO_2049 (O_2049,N_24075,N_24821);
xor UO_2050 (O_2050,N_24630,N_24302);
nor UO_2051 (O_2051,N_24068,N_24762);
xor UO_2052 (O_2052,N_24213,N_24974);
nand UO_2053 (O_2053,N_24687,N_24032);
nor UO_2054 (O_2054,N_24174,N_24542);
and UO_2055 (O_2055,N_24440,N_24087);
and UO_2056 (O_2056,N_24959,N_24294);
or UO_2057 (O_2057,N_24380,N_24764);
nand UO_2058 (O_2058,N_24986,N_24430);
xnor UO_2059 (O_2059,N_24430,N_24802);
nand UO_2060 (O_2060,N_24325,N_24006);
nand UO_2061 (O_2061,N_24587,N_24198);
nor UO_2062 (O_2062,N_24266,N_24181);
or UO_2063 (O_2063,N_24010,N_24885);
xnor UO_2064 (O_2064,N_24998,N_24701);
xnor UO_2065 (O_2065,N_24483,N_24870);
or UO_2066 (O_2066,N_24802,N_24842);
and UO_2067 (O_2067,N_24650,N_24953);
xor UO_2068 (O_2068,N_24551,N_24584);
nor UO_2069 (O_2069,N_24561,N_24938);
nand UO_2070 (O_2070,N_24982,N_24615);
nor UO_2071 (O_2071,N_24265,N_24000);
nor UO_2072 (O_2072,N_24020,N_24718);
nor UO_2073 (O_2073,N_24019,N_24596);
or UO_2074 (O_2074,N_24846,N_24748);
xor UO_2075 (O_2075,N_24124,N_24269);
xnor UO_2076 (O_2076,N_24152,N_24113);
or UO_2077 (O_2077,N_24833,N_24815);
and UO_2078 (O_2078,N_24115,N_24118);
and UO_2079 (O_2079,N_24001,N_24244);
and UO_2080 (O_2080,N_24269,N_24656);
or UO_2081 (O_2081,N_24554,N_24093);
nor UO_2082 (O_2082,N_24654,N_24543);
nor UO_2083 (O_2083,N_24009,N_24861);
xor UO_2084 (O_2084,N_24618,N_24013);
and UO_2085 (O_2085,N_24845,N_24382);
nand UO_2086 (O_2086,N_24018,N_24222);
nand UO_2087 (O_2087,N_24942,N_24151);
and UO_2088 (O_2088,N_24290,N_24896);
nor UO_2089 (O_2089,N_24610,N_24684);
xnor UO_2090 (O_2090,N_24861,N_24295);
nand UO_2091 (O_2091,N_24676,N_24089);
nor UO_2092 (O_2092,N_24190,N_24927);
and UO_2093 (O_2093,N_24307,N_24291);
nand UO_2094 (O_2094,N_24875,N_24374);
or UO_2095 (O_2095,N_24732,N_24424);
or UO_2096 (O_2096,N_24995,N_24542);
xor UO_2097 (O_2097,N_24852,N_24580);
nor UO_2098 (O_2098,N_24329,N_24772);
and UO_2099 (O_2099,N_24229,N_24753);
nand UO_2100 (O_2100,N_24699,N_24058);
and UO_2101 (O_2101,N_24187,N_24605);
nor UO_2102 (O_2102,N_24831,N_24315);
or UO_2103 (O_2103,N_24927,N_24401);
or UO_2104 (O_2104,N_24818,N_24622);
or UO_2105 (O_2105,N_24094,N_24957);
nor UO_2106 (O_2106,N_24065,N_24762);
nor UO_2107 (O_2107,N_24776,N_24090);
nor UO_2108 (O_2108,N_24606,N_24774);
nor UO_2109 (O_2109,N_24666,N_24599);
or UO_2110 (O_2110,N_24120,N_24876);
or UO_2111 (O_2111,N_24986,N_24992);
nor UO_2112 (O_2112,N_24467,N_24544);
and UO_2113 (O_2113,N_24359,N_24252);
and UO_2114 (O_2114,N_24379,N_24408);
xnor UO_2115 (O_2115,N_24280,N_24665);
and UO_2116 (O_2116,N_24251,N_24234);
nand UO_2117 (O_2117,N_24561,N_24986);
nor UO_2118 (O_2118,N_24273,N_24869);
and UO_2119 (O_2119,N_24923,N_24110);
nand UO_2120 (O_2120,N_24825,N_24460);
and UO_2121 (O_2121,N_24007,N_24554);
nor UO_2122 (O_2122,N_24654,N_24500);
nand UO_2123 (O_2123,N_24457,N_24681);
nand UO_2124 (O_2124,N_24545,N_24980);
and UO_2125 (O_2125,N_24976,N_24656);
xnor UO_2126 (O_2126,N_24041,N_24811);
nand UO_2127 (O_2127,N_24456,N_24722);
nor UO_2128 (O_2128,N_24931,N_24640);
nor UO_2129 (O_2129,N_24871,N_24466);
and UO_2130 (O_2130,N_24778,N_24897);
xnor UO_2131 (O_2131,N_24294,N_24629);
nor UO_2132 (O_2132,N_24477,N_24539);
or UO_2133 (O_2133,N_24198,N_24506);
nor UO_2134 (O_2134,N_24847,N_24491);
and UO_2135 (O_2135,N_24394,N_24764);
nor UO_2136 (O_2136,N_24319,N_24810);
nand UO_2137 (O_2137,N_24679,N_24304);
and UO_2138 (O_2138,N_24806,N_24879);
and UO_2139 (O_2139,N_24278,N_24269);
or UO_2140 (O_2140,N_24170,N_24837);
xor UO_2141 (O_2141,N_24690,N_24907);
nand UO_2142 (O_2142,N_24163,N_24534);
nor UO_2143 (O_2143,N_24943,N_24196);
or UO_2144 (O_2144,N_24817,N_24661);
nor UO_2145 (O_2145,N_24029,N_24028);
nand UO_2146 (O_2146,N_24348,N_24030);
nand UO_2147 (O_2147,N_24356,N_24892);
or UO_2148 (O_2148,N_24281,N_24016);
and UO_2149 (O_2149,N_24864,N_24801);
and UO_2150 (O_2150,N_24499,N_24843);
or UO_2151 (O_2151,N_24574,N_24113);
or UO_2152 (O_2152,N_24759,N_24504);
or UO_2153 (O_2153,N_24218,N_24312);
and UO_2154 (O_2154,N_24408,N_24089);
and UO_2155 (O_2155,N_24259,N_24734);
xor UO_2156 (O_2156,N_24305,N_24832);
xnor UO_2157 (O_2157,N_24427,N_24674);
or UO_2158 (O_2158,N_24861,N_24844);
nor UO_2159 (O_2159,N_24483,N_24281);
and UO_2160 (O_2160,N_24964,N_24960);
and UO_2161 (O_2161,N_24312,N_24622);
nand UO_2162 (O_2162,N_24548,N_24449);
nand UO_2163 (O_2163,N_24985,N_24947);
nand UO_2164 (O_2164,N_24055,N_24828);
xor UO_2165 (O_2165,N_24834,N_24781);
nor UO_2166 (O_2166,N_24042,N_24683);
xor UO_2167 (O_2167,N_24435,N_24834);
or UO_2168 (O_2168,N_24637,N_24729);
nor UO_2169 (O_2169,N_24530,N_24902);
nor UO_2170 (O_2170,N_24151,N_24359);
nor UO_2171 (O_2171,N_24414,N_24791);
or UO_2172 (O_2172,N_24792,N_24796);
nand UO_2173 (O_2173,N_24470,N_24943);
and UO_2174 (O_2174,N_24569,N_24536);
nand UO_2175 (O_2175,N_24678,N_24751);
nand UO_2176 (O_2176,N_24011,N_24115);
nand UO_2177 (O_2177,N_24351,N_24033);
xnor UO_2178 (O_2178,N_24969,N_24766);
xor UO_2179 (O_2179,N_24899,N_24946);
xnor UO_2180 (O_2180,N_24954,N_24722);
xnor UO_2181 (O_2181,N_24612,N_24910);
xnor UO_2182 (O_2182,N_24700,N_24153);
nand UO_2183 (O_2183,N_24092,N_24866);
xor UO_2184 (O_2184,N_24261,N_24375);
nand UO_2185 (O_2185,N_24999,N_24590);
nand UO_2186 (O_2186,N_24220,N_24973);
nand UO_2187 (O_2187,N_24719,N_24473);
nand UO_2188 (O_2188,N_24633,N_24859);
nand UO_2189 (O_2189,N_24653,N_24487);
nand UO_2190 (O_2190,N_24548,N_24795);
nand UO_2191 (O_2191,N_24789,N_24085);
nor UO_2192 (O_2192,N_24341,N_24303);
and UO_2193 (O_2193,N_24317,N_24882);
nor UO_2194 (O_2194,N_24105,N_24856);
xnor UO_2195 (O_2195,N_24532,N_24417);
or UO_2196 (O_2196,N_24528,N_24583);
xnor UO_2197 (O_2197,N_24310,N_24740);
and UO_2198 (O_2198,N_24790,N_24611);
nand UO_2199 (O_2199,N_24284,N_24570);
and UO_2200 (O_2200,N_24687,N_24202);
xnor UO_2201 (O_2201,N_24807,N_24794);
xnor UO_2202 (O_2202,N_24405,N_24442);
xor UO_2203 (O_2203,N_24703,N_24401);
nor UO_2204 (O_2204,N_24357,N_24262);
and UO_2205 (O_2205,N_24031,N_24841);
nand UO_2206 (O_2206,N_24144,N_24296);
or UO_2207 (O_2207,N_24227,N_24035);
xor UO_2208 (O_2208,N_24454,N_24803);
and UO_2209 (O_2209,N_24986,N_24410);
nor UO_2210 (O_2210,N_24667,N_24234);
nand UO_2211 (O_2211,N_24888,N_24789);
nor UO_2212 (O_2212,N_24386,N_24911);
nor UO_2213 (O_2213,N_24731,N_24867);
xor UO_2214 (O_2214,N_24413,N_24609);
xor UO_2215 (O_2215,N_24487,N_24972);
and UO_2216 (O_2216,N_24582,N_24626);
nand UO_2217 (O_2217,N_24146,N_24789);
or UO_2218 (O_2218,N_24220,N_24859);
nor UO_2219 (O_2219,N_24032,N_24845);
nand UO_2220 (O_2220,N_24929,N_24443);
xnor UO_2221 (O_2221,N_24412,N_24498);
nor UO_2222 (O_2222,N_24392,N_24636);
or UO_2223 (O_2223,N_24032,N_24575);
or UO_2224 (O_2224,N_24652,N_24660);
nor UO_2225 (O_2225,N_24205,N_24496);
or UO_2226 (O_2226,N_24345,N_24229);
nand UO_2227 (O_2227,N_24430,N_24476);
nor UO_2228 (O_2228,N_24575,N_24329);
or UO_2229 (O_2229,N_24697,N_24985);
xnor UO_2230 (O_2230,N_24591,N_24539);
and UO_2231 (O_2231,N_24589,N_24691);
or UO_2232 (O_2232,N_24073,N_24400);
or UO_2233 (O_2233,N_24889,N_24721);
and UO_2234 (O_2234,N_24446,N_24253);
nand UO_2235 (O_2235,N_24897,N_24091);
nand UO_2236 (O_2236,N_24441,N_24865);
and UO_2237 (O_2237,N_24813,N_24726);
xor UO_2238 (O_2238,N_24215,N_24444);
nor UO_2239 (O_2239,N_24636,N_24488);
and UO_2240 (O_2240,N_24256,N_24293);
or UO_2241 (O_2241,N_24300,N_24423);
and UO_2242 (O_2242,N_24322,N_24187);
and UO_2243 (O_2243,N_24021,N_24703);
xor UO_2244 (O_2244,N_24583,N_24616);
nor UO_2245 (O_2245,N_24966,N_24165);
or UO_2246 (O_2246,N_24522,N_24236);
and UO_2247 (O_2247,N_24556,N_24203);
xnor UO_2248 (O_2248,N_24888,N_24029);
nor UO_2249 (O_2249,N_24232,N_24133);
and UO_2250 (O_2250,N_24148,N_24196);
nand UO_2251 (O_2251,N_24093,N_24927);
or UO_2252 (O_2252,N_24148,N_24661);
xnor UO_2253 (O_2253,N_24510,N_24597);
nand UO_2254 (O_2254,N_24763,N_24154);
or UO_2255 (O_2255,N_24487,N_24744);
or UO_2256 (O_2256,N_24311,N_24041);
xnor UO_2257 (O_2257,N_24510,N_24739);
xor UO_2258 (O_2258,N_24972,N_24787);
and UO_2259 (O_2259,N_24777,N_24220);
or UO_2260 (O_2260,N_24410,N_24675);
nand UO_2261 (O_2261,N_24775,N_24268);
and UO_2262 (O_2262,N_24037,N_24096);
xor UO_2263 (O_2263,N_24594,N_24171);
or UO_2264 (O_2264,N_24987,N_24568);
xnor UO_2265 (O_2265,N_24249,N_24804);
and UO_2266 (O_2266,N_24388,N_24362);
and UO_2267 (O_2267,N_24737,N_24879);
and UO_2268 (O_2268,N_24259,N_24513);
nand UO_2269 (O_2269,N_24947,N_24069);
xor UO_2270 (O_2270,N_24934,N_24644);
and UO_2271 (O_2271,N_24743,N_24486);
nand UO_2272 (O_2272,N_24363,N_24085);
nor UO_2273 (O_2273,N_24018,N_24116);
nand UO_2274 (O_2274,N_24627,N_24944);
nor UO_2275 (O_2275,N_24441,N_24772);
nand UO_2276 (O_2276,N_24760,N_24733);
or UO_2277 (O_2277,N_24696,N_24177);
or UO_2278 (O_2278,N_24643,N_24505);
or UO_2279 (O_2279,N_24752,N_24637);
xor UO_2280 (O_2280,N_24107,N_24737);
or UO_2281 (O_2281,N_24706,N_24443);
or UO_2282 (O_2282,N_24842,N_24485);
xor UO_2283 (O_2283,N_24022,N_24652);
nand UO_2284 (O_2284,N_24574,N_24453);
nor UO_2285 (O_2285,N_24326,N_24485);
or UO_2286 (O_2286,N_24496,N_24314);
nor UO_2287 (O_2287,N_24799,N_24620);
nor UO_2288 (O_2288,N_24965,N_24896);
nand UO_2289 (O_2289,N_24388,N_24259);
nand UO_2290 (O_2290,N_24734,N_24960);
nor UO_2291 (O_2291,N_24499,N_24802);
or UO_2292 (O_2292,N_24479,N_24299);
xor UO_2293 (O_2293,N_24319,N_24132);
nor UO_2294 (O_2294,N_24306,N_24315);
nor UO_2295 (O_2295,N_24164,N_24033);
or UO_2296 (O_2296,N_24042,N_24720);
nor UO_2297 (O_2297,N_24939,N_24192);
nor UO_2298 (O_2298,N_24028,N_24831);
nor UO_2299 (O_2299,N_24815,N_24514);
nor UO_2300 (O_2300,N_24836,N_24944);
or UO_2301 (O_2301,N_24606,N_24770);
or UO_2302 (O_2302,N_24959,N_24781);
and UO_2303 (O_2303,N_24848,N_24719);
nand UO_2304 (O_2304,N_24222,N_24313);
nor UO_2305 (O_2305,N_24847,N_24630);
nor UO_2306 (O_2306,N_24738,N_24301);
and UO_2307 (O_2307,N_24598,N_24221);
nor UO_2308 (O_2308,N_24428,N_24494);
nor UO_2309 (O_2309,N_24865,N_24540);
nand UO_2310 (O_2310,N_24441,N_24987);
nand UO_2311 (O_2311,N_24073,N_24913);
nand UO_2312 (O_2312,N_24423,N_24941);
nor UO_2313 (O_2313,N_24972,N_24893);
or UO_2314 (O_2314,N_24987,N_24215);
xnor UO_2315 (O_2315,N_24495,N_24892);
nor UO_2316 (O_2316,N_24936,N_24829);
or UO_2317 (O_2317,N_24601,N_24485);
xor UO_2318 (O_2318,N_24743,N_24525);
nand UO_2319 (O_2319,N_24554,N_24801);
nor UO_2320 (O_2320,N_24631,N_24386);
nand UO_2321 (O_2321,N_24031,N_24604);
and UO_2322 (O_2322,N_24110,N_24561);
nor UO_2323 (O_2323,N_24279,N_24905);
or UO_2324 (O_2324,N_24755,N_24268);
nand UO_2325 (O_2325,N_24917,N_24497);
xor UO_2326 (O_2326,N_24200,N_24074);
nor UO_2327 (O_2327,N_24765,N_24384);
nand UO_2328 (O_2328,N_24847,N_24753);
xnor UO_2329 (O_2329,N_24178,N_24326);
nand UO_2330 (O_2330,N_24932,N_24548);
nand UO_2331 (O_2331,N_24388,N_24370);
xor UO_2332 (O_2332,N_24697,N_24104);
nor UO_2333 (O_2333,N_24670,N_24940);
nor UO_2334 (O_2334,N_24424,N_24077);
or UO_2335 (O_2335,N_24686,N_24785);
nand UO_2336 (O_2336,N_24611,N_24477);
nor UO_2337 (O_2337,N_24830,N_24082);
or UO_2338 (O_2338,N_24504,N_24323);
nand UO_2339 (O_2339,N_24517,N_24896);
and UO_2340 (O_2340,N_24869,N_24731);
and UO_2341 (O_2341,N_24267,N_24958);
nor UO_2342 (O_2342,N_24207,N_24535);
xor UO_2343 (O_2343,N_24630,N_24871);
and UO_2344 (O_2344,N_24444,N_24358);
or UO_2345 (O_2345,N_24572,N_24802);
nor UO_2346 (O_2346,N_24371,N_24229);
nand UO_2347 (O_2347,N_24263,N_24629);
nand UO_2348 (O_2348,N_24118,N_24090);
nand UO_2349 (O_2349,N_24948,N_24162);
xor UO_2350 (O_2350,N_24975,N_24087);
nand UO_2351 (O_2351,N_24605,N_24320);
nand UO_2352 (O_2352,N_24990,N_24693);
and UO_2353 (O_2353,N_24699,N_24352);
nand UO_2354 (O_2354,N_24086,N_24455);
or UO_2355 (O_2355,N_24041,N_24429);
or UO_2356 (O_2356,N_24646,N_24334);
nand UO_2357 (O_2357,N_24572,N_24964);
nand UO_2358 (O_2358,N_24928,N_24748);
nand UO_2359 (O_2359,N_24133,N_24375);
nor UO_2360 (O_2360,N_24389,N_24908);
nand UO_2361 (O_2361,N_24865,N_24442);
and UO_2362 (O_2362,N_24674,N_24542);
nand UO_2363 (O_2363,N_24327,N_24668);
nand UO_2364 (O_2364,N_24828,N_24509);
and UO_2365 (O_2365,N_24765,N_24946);
xnor UO_2366 (O_2366,N_24191,N_24730);
nand UO_2367 (O_2367,N_24729,N_24714);
xor UO_2368 (O_2368,N_24675,N_24263);
or UO_2369 (O_2369,N_24895,N_24419);
nor UO_2370 (O_2370,N_24754,N_24752);
nand UO_2371 (O_2371,N_24903,N_24055);
nand UO_2372 (O_2372,N_24403,N_24970);
and UO_2373 (O_2373,N_24050,N_24943);
and UO_2374 (O_2374,N_24219,N_24064);
and UO_2375 (O_2375,N_24005,N_24989);
nand UO_2376 (O_2376,N_24711,N_24032);
nand UO_2377 (O_2377,N_24455,N_24471);
and UO_2378 (O_2378,N_24857,N_24141);
or UO_2379 (O_2379,N_24982,N_24599);
xnor UO_2380 (O_2380,N_24651,N_24288);
nor UO_2381 (O_2381,N_24072,N_24220);
nor UO_2382 (O_2382,N_24530,N_24367);
xor UO_2383 (O_2383,N_24735,N_24850);
xor UO_2384 (O_2384,N_24702,N_24145);
nand UO_2385 (O_2385,N_24224,N_24187);
nand UO_2386 (O_2386,N_24557,N_24658);
xor UO_2387 (O_2387,N_24492,N_24793);
nand UO_2388 (O_2388,N_24142,N_24055);
nor UO_2389 (O_2389,N_24647,N_24445);
and UO_2390 (O_2390,N_24093,N_24776);
xnor UO_2391 (O_2391,N_24998,N_24541);
xor UO_2392 (O_2392,N_24013,N_24104);
nor UO_2393 (O_2393,N_24074,N_24000);
xnor UO_2394 (O_2394,N_24266,N_24448);
or UO_2395 (O_2395,N_24874,N_24251);
or UO_2396 (O_2396,N_24012,N_24523);
nor UO_2397 (O_2397,N_24512,N_24202);
or UO_2398 (O_2398,N_24127,N_24371);
or UO_2399 (O_2399,N_24436,N_24853);
and UO_2400 (O_2400,N_24607,N_24386);
or UO_2401 (O_2401,N_24904,N_24466);
nand UO_2402 (O_2402,N_24801,N_24419);
or UO_2403 (O_2403,N_24810,N_24579);
and UO_2404 (O_2404,N_24810,N_24112);
or UO_2405 (O_2405,N_24824,N_24859);
xor UO_2406 (O_2406,N_24046,N_24786);
nor UO_2407 (O_2407,N_24380,N_24150);
nor UO_2408 (O_2408,N_24000,N_24867);
nand UO_2409 (O_2409,N_24268,N_24911);
nand UO_2410 (O_2410,N_24595,N_24489);
nor UO_2411 (O_2411,N_24403,N_24270);
or UO_2412 (O_2412,N_24559,N_24310);
and UO_2413 (O_2413,N_24037,N_24486);
xor UO_2414 (O_2414,N_24346,N_24460);
and UO_2415 (O_2415,N_24752,N_24282);
or UO_2416 (O_2416,N_24809,N_24331);
or UO_2417 (O_2417,N_24650,N_24850);
xor UO_2418 (O_2418,N_24636,N_24165);
or UO_2419 (O_2419,N_24211,N_24213);
xnor UO_2420 (O_2420,N_24776,N_24396);
nand UO_2421 (O_2421,N_24195,N_24709);
or UO_2422 (O_2422,N_24293,N_24399);
nor UO_2423 (O_2423,N_24871,N_24125);
xor UO_2424 (O_2424,N_24974,N_24513);
nand UO_2425 (O_2425,N_24154,N_24127);
or UO_2426 (O_2426,N_24583,N_24153);
and UO_2427 (O_2427,N_24800,N_24310);
or UO_2428 (O_2428,N_24056,N_24767);
nand UO_2429 (O_2429,N_24077,N_24877);
nand UO_2430 (O_2430,N_24982,N_24100);
or UO_2431 (O_2431,N_24310,N_24917);
or UO_2432 (O_2432,N_24562,N_24864);
and UO_2433 (O_2433,N_24281,N_24751);
nor UO_2434 (O_2434,N_24853,N_24323);
nor UO_2435 (O_2435,N_24354,N_24992);
or UO_2436 (O_2436,N_24153,N_24426);
or UO_2437 (O_2437,N_24566,N_24284);
and UO_2438 (O_2438,N_24915,N_24961);
or UO_2439 (O_2439,N_24588,N_24478);
and UO_2440 (O_2440,N_24001,N_24324);
xnor UO_2441 (O_2441,N_24203,N_24545);
or UO_2442 (O_2442,N_24616,N_24016);
nand UO_2443 (O_2443,N_24471,N_24765);
or UO_2444 (O_2444,N_24658,N_24483);
nand UO_2445 (O_2445,N_24733,N_24966);
xor UO_2446 (O_2446,N_24173,N_24583);
nand UO_2447 (O_2447,N_24150,N_24630);
and UO_2448 (O_2448,N_24734,N_24427);
xnor UO_2449 (O_2449,N_24479,N_24276);
or UO_2450 (O_2450,N_24699,N_24428);
xnor UO_2451 (O_2451,N_24469,N_24581);
and UO_2452 (O_2452,N_24110,N_24664);
nor UO_2453 (O_2453,N_24320,N_24323);
xor UO_2454 (O_2454,N_24184,N_24604);
xnor UO_2455 (O_2455,N_24236,N_24074);
or UO_2456 (O_2456,N_24040,N_24580);
xnor UO_2457 (O_2457,N_24619,N_24110);
and UO_2458 (O_2458,N_24099,N_24682);
or UO_2459 (O_2459,N_24959,N_24714);
or UO_2460 (O_2460,N_24311,N_24673);
or UO_2461 (O_2461,N_24581,N_24730);
xor UO_2462 (O_2462,N_24352,N_24238);
and UO_2463 (O_2463,N_24695,N_24755);
and UO_2464 (O_2464,N_24641,N_24429);
xnor UO_2465 (O_2465,N_24348,N_24759);
xor UO_2466 (O_2466,N_24334,N_24064);
or UO_2467 (O_2467,N_24984,N_24834);
nand UO_2468 (O_2468,N_24248,N_24040);
nor UO_2469 (O_2469,N_24221,N_24251);
or UO_2470 (O_2470,N_24636,N_24931);
and UO_2471 (O_2471,N_24399,N_24448);
nor UO_2472 (O_2472,N_24152,N_24326);
and UO_2473 (O_2473,N_24344,N_24190);
or UO_2474 (O_2474,N_24538,N_24273);
or UO_2475 (O_2475,N_24591,N_24041);
xnor UO_2476 (O_2476,N_24504,N_24397);
nand UO_2477 (O_2477,N_24625,N_24056);
or UO_2478 (O_2478,N_24409,N_24076);
or UO_2479 (O_2479,N_24331,N_24733);
or UO_2480 (O_2480,N_24762,N_24659);
and UO_2481 (O_2481,N_24513,N_24232);
or UO_2482 (O_2482,N_24727,N_24764);
and UO_2483 (O_2483,N_24277,N_24723);
nand UO_2484 (O_2484,N_24134,N_24029);
or UO_2485 (O_2485,N_24329,N_24031);
xnor UO_2486 (O_2486,N_24454,N_24836);
nand UO_2487 (O_2487,N_24889,N_24494);
and UO_2488 (O_2488,N_24973,N_24551);
nand UO_2489 (O_2489,N_24533,N_24170);
nand UO_2490 (O_2490,N_24560,N_24974);
nor UO_2491 (O_2491,N_24625,N_24276);
nor UO_2492 (O_2492,N_24625,N_24087);
xnor UO_2493 (O_2493,N_24413,N_24758);
nor UO_2494 (O_2494,N_24983,N_24724);
and UO_2495 (O_2495,N_24430,N_24738);
nor UO_2496 (O_2496,N_24783,N_24334);
and UO_2497 (O_2497,N_24441,N_24960);
nand UO_2498 (O_2498,N_24842,N_24985);
or UO_2499 (O_2499,N_24127,N_24517);
nand UO_2500 (O_2500,N_24029,N_24515);
nand UO_2501 (O_2501,N_24055,N_24876);
or UO_2502 (O_2502,N_24621,N_24150);
or UO_2503 (O_2503,N_24579,N_24134);
nand UO_2504 (O_2504,N_24887,N_24975);
nand UO_2505 (O_2505,N_24519,N_24136);
and UO_2506 (O_2506,N_24764,N_24955);
nand UO_2507 (O_2507,N_24991,N_24159);
xor UO_2508 (O_2508,N_24023,N_24210);
nand UO_2509 (O_2509,N_24943,N_24401);
xor UO_2510 (O_2510,N_24335,N_24895);
nor UO_2511 (O_2511,N_24577,N_24630);
xor UO_2512 (O_2512,N_24141,N_24217);
xor UO_2513 (O_2513,N_24169,N_24240);
nor UO_2514 (O_2514,N_24927,N_24972);
xnor UO_2515 (O_2515,N_24019,N_24020);
or UO_2516 (O_2516,N_24606,N_24033);
nand UO_2517 (O_2517,N_24157,N_24385);
and UO_2518 (O_2518,N_24955,N_24982);
nor UO_2519 (O_2519,N_24651,N_24096);
nor UO_2520 (O_2520,N_24717,N_24273);
or UO_2521 (O_2521,N_24302,N_24601);
or UO_2522 (O_2522,N_24729,N_24607);
or UO_2523 (O_2523,N_24766,N_24228);
nor UO_2524 (O_2524,N_24437,N_24601);
nor UO_2525 (O_2525,N_24460,N_24424);
and UO_2526 (O_2526,N_24233,N_24205);
or UO_2527 (O_2527,N_24261,N_24769);
and UO_2528 (O_2528,N_24847,N_24613);
and UO_2529 (O_2529,N_24212,N_24625);
nor UO_2530 (O_2530,N_24948,N_24128);
and UO_2531 (O_2531,N_24526,N_24034);
xor UO_2532 (O_2532,N_24474,N_24107);
nand UO_2533 (O_2533,N_24900,N_24865);
nand UO_2534 (O_2534,N_24022,N_24110);
and UO_2535 (O_2535,N_24425,N_24982);
nand UO_2536 (O_2536,N_24239,N_24500);
nand UO_2537 (O_2537,N_24263,N_24513);
nor UO_2538 (O_2538,N_24197,N_24563);
xor UO_2539 (O_2539,N_24293,N_24547);
and UO_2540 (O_2540,N_24319,N_24586);
or UO_2541 (O_2541,N_24452,N_24591);
nor UO_2542 (O_2542,N_24019,N_24333);
nand UO_2543 (O_2543,N_24937,N_24177);
xor UO_2544 (O_2544,N_24527,N_24760);
xnor UO_2545 (O_2545,N_24476,N_24587);
xor UO_2546 (O_2546,N_24833,N_24896);
or UO_2547 (O_2547,N_24311,N_24322);
nand UO_2548 (O_2548,N_24483,N_24156);
nand UO_2549 (O_2549,N_24888,N_24257);
nand UO_2550 (O_2550,N_24253,N_24358);
xor UO_2551 (O_2551,N_24194,N_24534);
nand UO_2552 (O_2552,N_24608,N_24899);
nor UO_2553 (O_2553,N_24709,N_24548);
xnor UO_2554 (O_2554,N_24175,N_24058);
nor UO_2555 (O_2555,N_24578,N_24443);
and UO_2556 (O_2556,N_24456,N_24598);
nor UO_2557 (O_2557,N_24916,N_24340);
and UO_2558 (O_2558,N_24515,N_24284);
nand UO_2559 (O_2559,N_24179,N_24188);
nor UO_2560 (O_2560,N_24486,N_24979);
xor UO_2561 (O_2561,N_24015,N_24312);
nor UO_2562 (O_2562,N_24235,N_24654);
or UO_2563 (O_2563,N_24447,N_24885);
nor UO_2564 (O_2564,N_24800,N_24449);
nor UO_2565 (O_2565,N_24022,N_24397);
or UO_2566 (O_2566,N_24876,N_24596);
or UO_2567 (O_2567,N_24489,N_24855);
nand UO_2568 (O_2568,N_24100,N_24010);
nand UO_2569 (O_2569,N_24051,N_24386);
xor UO_2570 (O_2570,N_24820,N_24958);
nand UO_2571 (O_2571,N_24211,N_24941);
or UO_2572 (O_2572,N_24152,N_24532);
or UO_2573 (O_2573,N_24412,N_24523);
and UO_2574 (O_2574,N_24753,N_24240);
xnor UO_2575 (O_2575,N_24366,N_24964);
or UO_2576 (O_2576,N_24520,N_24010);
xnor UO_2577 (O_2577,N_24025,N_24980);
nor UO_2578 (O_2578,N_24032,N_24882);
nand UO_2579 (O_2579,N_24495,N_24510);
or UO_2580 (O_2580,N_24867,N_24069);
and UO_2581 (O_2581,N_24984,N_24733);
nand UO_2582 (O_2582,N_24470,N_24166);
or UO_2583 (O_2583,N_24003,N_24900);
or UO_2584 (O_2584,N_24482,N_24873);
nor UO_2585 (O_2585,N_24737,N_24528);
xor UO_2586 (O_2586,N_24863,N_24154);
xnor UO_2587 (O_2587,N_24560,N_24342);
or UO_2588 (O_2588,N_24837,N_24597);
xor UO_2589 (O_2589,N_24765,N_24825);
and UO_2590 (O_2590,N_24641,N_24345);
or UO_2591 (O_2591,N_24226,N_24732);
nor UO_2592 (O_2592,N_24915,N_24422);
nor UO_2593 (O_2593,N_24459,N_24431);
xnor UO_2594 (O_2594,N_24457,N_24043);
and UO_2595 (O_2595,N_24426,N_24880);
nand UO_2596 (O_2596,N_24566,N_24322);
xor UO_2597 (O_2597,N_24011,N_24084);
nand UO_2598 (O_2598,N_24193,N_24365);
nor UO_2599 (O_2599,N_24677,N_24459);
xor UO_2600 (O_2600,N_24928,N_24385);
and UO_2601 (O_2601,N_24418,N_24282);
and UO_2602 (O_2602,N_24748,N_24613);
xor UO_2603 (O_2603,N_24601,N_24950);
nor UO_2604 (O_2604,N_24339,N_24221);
nand UO_2605 (O_2605,N_24655,N_24243);
and UO_2606 (O_2606,N_24333,N_24726);
nand UO_2607 (O_2607,N_24741,N_24713);
or UO_2608 (O_2608,N_24043,N_24435);
or UO_2609 (O_2609,N_24884,N_24343);
nand UO_2610 (O_2610,N_24898,N_24741);
or UO_2611 (O_2611,N_24777,N_24967);
or UO_2612 (O_2612,N_24979,N_24890);
or UO_2613 (O_2613,N_24641,N_24218);
nor UO_2614 (O_2614,N_24801,N_24013);
or UO_2615 (O_2615,N_24363,N_24497);
or UO_2616 (O_2616,N_24839,N_24798);
xor UO_2617 (O_2617,N_24771,N_24333);
nand UO_2618 (O_2618,N_24861,N_24767);
xor UO_2619 (O_2619,N_24655,N_24384);
nor UO_2620 (O_2620,N_24576,N_24315);
nor UO_2621 (O_2621,N_24323,N_24890);
and UO_2622 (O_2622,N_24446,N_24117);
or UO_2623 (O_2623,N_24607,N_24763);
nor UO_2624 (O_2624,N_24214,N_24814);
nor UO_2625 (O_2625,N_24865,N_24392);
or UO_2626 (O_2626,N_24576,N_24096);
nor UO_2627 (O_2627,N_24278,N_24990);
nor UO_2628 (O_2628,N_24966,N_24342);
xnor UO_2629 (O_2629,N_24983,N_24567);
or UO_2630 (O_2630,N_24284,N_24901);
nand UO_2631 (O_2631,N_24334,N_24734);
or UO_2632 (O_2632,N_24781,N_24324);
or UO_2633 (O_2633,N_24466,N_24927);
or UO_2634 (O_2634,N_24531,N_24537);
xnor UO_2635 (O_2635,N_24920,N_24359);
nor UO_2636 (O_2636,N_24109,N_24402);
and UO_2637 (O_2637,N_24842,N_24523);
or UO_2638 (O_2638,N_24351,N_24677);
xnor UO_2639 (O_2639,N_24963,N_24200);
xnor UO_2640 (O_2640,N_24698,N_24237);
xor UO_2641 (O_2641,N_24856,N_24254);
nand UO_2642 (O_2642,N_24661,N_24702);
nand UO_2643 (O_2643,N_24003,N_24974);
and UO_2644 (O_2644,N_24878,N_24317);
or UO_2645 (O_2645,N_24252,N_24324);
xnor UO_2646 (O_2646,N_24309,N_24922);
nand UO_2647 (O_2647,N_24295,N_24226);
or UO_2648 (O_2648,N_24375,N_24328);
xnor UO_2649 (O_2649,N_24449,N_24872);
and UO_2650 (O_2650,N_24528,N_24905);
nor UO_2651 (O_2651,N_24451,N_24486);
or UO_2652 (O_2652,N_24196,N_24175);
nand UO_2653 (O_2653,N_24051,N_24408);
or UO_2654 (O_2654,N_24057,N_24591);
nor UO_2655 (O_2655,N_24846,N_24254);
and UO_2656 (O_2656,N_24439,N_24064);
xnor UO_2657 (O_2657,N_24883,N_24278);
or UO_2658 (O_2658,N_24420,N_24320);
nand UO_2659 (O_2659,N_24982,N_24148);
and UO_2660 (O_2660,N_24151,N_24866);
nor UO_2661 (O_2661,N_24224,N_24039);
nand UO_2662 (O_2662,N_24794,N_24387);
or UO_2663 (O_2663,N_24480,N_24416);
nand UO_2664 (O_2664,N_24321,N_24714);
nand UO_2665 (O_2665,N_24433,N_24749);
nor UO_2666 (O_2666,N_24628,N_24546);
or UO_2667 (O_2667,N_24234,N_24337);
nand UO_2668 (O_2668,N_24637,N_24748);
xnor UO_2669 (O_2669,N_24909,N_24733);
nand UO_2670 (O_2670,N_24218,N_24887);
nor UO_2671 (O_2671,N_24934,N_24483);
nor UO_2672 (O_2672,N_24697,N_24135);
xnor UO_2673 (O_2673,N_24227,N_24073);
or UO_2674 (O_2674,N_24364,N_24436);
nand UO_2675 (O_2675,N_24785,N_24148);
xor UO_2676 (O_2676,N_24598,N_24591);
nor UO_2677 (O_2677,N_24765,N_24373);
nand UO_2678 (O_2678,N_24770,N_24938);
xnor UO_2679 (O_2679,N_24945,N_24689);
and UO_2680 (O_2680,N_24453,N_24288);
nand UO_2681 (O_2681,N_24978,N_24512);
and UO_2682 (O_2682,N_24936,N_24604);
or UO_2683 (O_2683,N_24163,N_24995);
or UO_2684 (O_2684,N_24083,N_24316);
xnor UO_2685 (O_2685,N_24442,N_24299);
nand UO_2686 (O_2686,N_24125,N_24070);
xnor UO_2687 (O_2687,N_24672,N_24025);
or UO_2688 (O_2688,N_24559,N_24650);
or UO_2689 (O_2689,N_24891,N_24008);
or UO_2690 (O_2690,N_24392,N_24190);
xor UO_2691 (O_2691,N_24060,N_24519);
xor UO_2692 (O_2692,N_24930,N_24195);
nor UO_2693 (O_2693,N_24885,N_24431);
xor UO_2694 (O_2694,N_24717,N_24615);
nand UO_2695 (O_2695,N_24926,N_24062);
or UO_2696 (O_2696,N_24306,N_24794);
xnor UO_2697 (O_2697,N_24673,N_24919);
or UO_2698 (O_2698,N_24020,N_24578);
and UO_2699 (O_2699,N_24421,N_24420);
xnor UO_2700 (O_2700,N_24250,N_24507);
nand UO_2701 (O_2701,N_24168,N_24197);
nor UO_2702 (O_2702,N_24249,N_24746);
xor UO_2703 (O_2703,N_24611,N_24773);
xor UO_2704 (O_2704,N_24085,N_24102);
and UO_2705 (O_2705,N_24545,N_24947);
nand UO_2706 (O_2706,N_24926,N_24223);
nand UO_2707 (O_2707,N_24907,N_24736);
nor UO_2708 (O_2708,N_24773,N_24130);
or UO_2709 (O_2709,N_24959,N_24639);
or UO_2710 (O_2710,N_24372,N_24206);
and UO_2711 (O_2711,N_24687,N_24551);
nor UO_2712 (O_2712,N_24200,N_24855);
nor UO_2713 (O_2713,N_24250,N_24959);
nor UO_2714 (O_2714,N_24974,N_24082);
or UO_2715 (O_2715,N_24822,N_24232);
xor UO_2716 (O_2716,N_24440,N_24384);
nand UO_2717 (O_2717,N_24191,N_24496);
nor UO_2718 (O_2718,N_24384,N_24233);
nor UO_2719 (O_2719,N_24129,N_24171);
nand UO_2720 (O_2720,N_24374,N_24945);
or UO_2721 (O_2721,N_24687,N_24117);
or UO_2722 (O_2722,N_24523,N_24755);
xnor UO_2723 (O_2723,N_24828,N_24425);
nand UO_2724 (O_2724,N_24670,N_24315);
or UO_2725 (O_2725,N_24905,N_24560);
nand UO_2726 (O_2726,N_24955,N_24894);
nand UO_2727 (O_2727,N_24504,N_24184);
or UO_2728 (O_2728,N_24747,N_24498);
xnor UO_2729 (O_2729,N_24922,N_24696);
nand UO_2730 (O_2730,N_24257,N_24724);
nand UO_2731 (O_2731,N_24641,N_24193);
nand UO_2732 (O_2732,N_24497,N_24418);
nand UO_2733 (O_2733,N_24076,N_24595);
or UO_2734 (O_2734,N_24395,N_24962);
xnor UO_2735 (O_2735,N_24613,N_24468);
nor UO_2736 (O_2736,N_24250,N_24711);
or UO_2737 (O_2737,N_24665,N_24909);
nor UO_2738 (O_2738,N_24548,N_24500);
and UO_2739 (O_2739,N_24970,N_24564);
nor UO_2740 (O_2740,N_24107,N_24597);
nor UO_2741 (O_2741,N_24800,N_24127);
and UO_2742 (O_2742,N_24960,N_24858);
and UO_2743 (O_2743,N_24266,N_24296);
nand UO_2744 (O_2744,N_24996,N_24060);
or UO_2745 (O_2745,N_24823,N_24628);
nand UO_2746 (O_2746,N_24532,N_24136);
and UO_2747 (O_2747,N_24169,N_24179);
or UO_2748 (O_2748,N_24185,N_24856);
nand UO_2749 (O_2749,N_24260,N_24509);
xnor UO_2750 (O_2750,N_24287,N_24645);
nor UO_2751 (O_2751,N_24884,N_24579);
and UO_2752 (O_2752,N_24973,N_24155);
nand UO_2753 (O_2753,N_24862,N_24797);
nand UO_2754 (O_2754,N_24420,N_24126);
nand UO_2755 (O_2755,N_24906,N_24582);
nor UO_2756 (O_2756,N_24155,N_24840);
nor UO_2757 (O_2757,N_24939,N_24867);
xnor UO_2758 (O_2758,N_24141,N_24367);
or UO_2759 (O_2759,N_24083,N_24016);
xnor UO_2760 (O_2760,N_24157,N_24930);
nor UO_2761 (O_2761,N_24313,N_24835);
or UO_2762 (O_2762,N_24791,N_24713);
xnor UO_2763 (O_2763,N_24584,N_24638);
nand UO_2764 (O_2764,N_24742,N_24573);
and UO_2765 (O_2765,N_24543,N_24620);
xor UO_2766 (O_2766,N_24947,N_24676);
nand UO_2767 (O_2767,N_24124,N_24512);
or UO_2768 (O_2768,N_24372,N_24418);
and UO_2769 (O_2769,N_24860,N_24369);
or UO_2770 (O_2770,N_24839,N_24780);
and UO_2771 (O_2771,N_24266,N_24651);
nor UO_2772 (O_2772,N_24657,N_24766);
or UO_2773 (O_2773,N_24904,N_24132);
nand UO_2774 (O_2774,N_24378,N_24377);
or UO_2775 (O_2775,N_24807,N_24129);
xor UO_2776 (O_2776,N_24799,N_24137);
or UO_2777 (O_2777,N_24519,N_24850);
or UO_2778 (O_2778,N_24689,N_24770);
xnor UO_2779 (O_2779,N_24705,N_24174);
or UO_2780 (O_2780,N_24416,N_24241);
and UO_2781 (O_2781,N_24496,N_24556);
and UO_2782 (O_2782,N_24752,N_24566);
nor UO_2783 (O_2783,N_24884,N_24832);
xor UO_2784 (O_2784,N_24572,N_24620);
xnor UO_2785 (O_2785,N_24795,N_24895);
xnor UO_2786 (O_2786,N_24102,N_24562);
or UO_2787 (O_2787,N_24857,N_24740);
and UO_2788 (O_2788,N_24565,N_24716);
nand UO_2789 (O_2789,N_24894,N_24730);
and UO_2790 (O_2790,N_24989,N_24967);
nand UO_2791 (O_2791,N_24432,N_24510);
and UO_2792 (O_2792,N_24960,N_24000);
nand UO_2793 (O_2793,N_24472,N_24961);
and UO_2794 (O_2794,N_24242,N_24464);
or UO_2795 (O_2795,N_24355,N_24594);
nand UO_2796 (O_2796,N_24695,N_24108);
nor UO_2797 (O_2797,N_24320,N_24343);
nor UO_2798 (O_2798,N_24852,N_24103);
nor UO_2799 (O_2799,N_24710,N_24533);
or UO_2800 (O_2800,N_24958,N_24792);
xor UO_2801 (O_2801,N_24418,N_24018);
or UO_2802 (O_2802,N_24746,N_24828);
and UO_2803 (O_2803,N_24121,N_24864);
and UO_2804 (O_2804,N_24094,N_24315);
nand UO_2805 (O_2805,N_24482,N_24870);
or UO_2806 (O_2806,N_24397,N_24583);
nand UO_2807 (O_2807,N_24859,N_24679);
xor UO_2808 (O_2808,N_24368,N_24723);
or UO_2809 (O_2809,N_24212,N_24531);
nand UO_2810 (O_2810,N_24971,N_24719);
xor UO_2811 (O_2811,N_24110,N_24554);
or UO_2812 (O_2812,N_24716,N_24440);
and UO_2813 (O_2813,N_24615,N_24358);
or UO_2814 (O_2814,N_24893,N_24945);
or UO_2815 (O_2815,N_24809,N_24823);
and UO_2816 (O_2816,N_24697,N_24278);
and UO_2817 (O_2817,N_24912,N_24639);
xnor UO_2818 (O_2818,N_24162,N_24203);
xor UO_2819 (O_2819,N_24171,N_24992);
xnor UO_2820 (O_2820,N_24767,N_24302);
and UO_2821 (O_2821,N_24351,N_24725);
and UO_2822 (O_2822,N_24696,N_24228);
or UO_2823 (O_2823,N_24632,N_24512);
nand UO_2824 (O_2824,N_24010,N_24926);
xnor UO_2825 (O_2825,N_24535,N_24374);
xor UO_2826 (O_2826,N_24776,N_24693);
xnor UO_2827 (O_2827,N_24133,N_24909);
and UO_2828 (O_2828,N_24269,N_24093);
and UO_2829 (O_2829,N_24915,N_24471);
or UO_2830 (O_2830,N_24490,N_24602);
xnor UO_2831 (O_2831,N_24252,N_24852);
nand UO_2832 (O_2832,N_24892,N_24084);
nand UO_2833 (O_2833,N_24352,N_24588);
xor UO_2834 (O_2834,N_24663,N_24141);
or UO_2835 (O_2835,N_24409,N_24652);
nor UO_2836 (O_2836,N_24997,N_24534);
or UO_2837 (O_2837,N_24625,N_24724);
nand UO_2838 (O_2838,N_24065,N_24200);
nor UO_2839 (O_2839,N_24812,N_24421);
or UO_2840 (O_2840,N_24118,N_24296);
xnor UO_2841 (O_2841,N_24425,N_24741);
and UO_2842 (O_2842,N_24964,N_24905);
and UO_2843 (O_2843,N_24126,N_24656);
xor UO_2844 (O_2844,N_24996,N_24279);
and UO_2845 (O_2845,N_24069,N_24852);
nand UO_2846 (O_2846,N_24879,N_24795);
nand UO_2847 (O_2847,N_24513,N_24337);
nand UO_2848 (O_2848,N_24634,N_24222);
nand UO_2849 (O_2849,N_24232,N_24095);
nand UO_2850 (O_2850,N_24821,N_24670);
xnor UO_2851 (O_2851,N_24987,N_24901);
nor UO_2852 (O_2852,N_24258,N_24268);
and UO_2853 (O_2853,N_24571,N_24813);
nand UO_2854 (O_2854,N_24442,N_24451);
and UO_2855 (O_2855,N_24023,N_24977);
nand UO_2856 (O_2856,N_24435,N_24503);
nor UO_2857 (O_2857,N_24998,N_24348);
nand UO_2858 (O_2858,N_24935,N_24516);
or UO_2859 (O_2859,N_24238,N_24167);
xor UO_2860 (O_2860,N_24160,N_24430);
nor UO_2861 (O_2861,N_24586,N_24429);
and UO_2862 (O_2862,N_24865,N_24509);
and UO_2863 (O_2863,N_24153,N_24511);
and UO_2864 (O_2864,N_24359,N_24972);
nand UO_2865 (O_2865,N_24548,N_24242);
nor UO_2866 (O_2866,N_24489,N_24794);
or UO_2867 (O_2867,N_24417,N_24670);
and UO_2868 (O_2868,N_24595,N_24074);
nand UO_2869 (O_2869,N_24820,N_24321);
or UO_2870 (O_2870,N_24090,N_24945);
nor UO_2871 (O_2871,N_24657,N_24501);
or UO_2872 (O_2872,N_24811,N_24338);
and UO_2873 (O_2873,N_24411,N_24624);
xnor UO_2874 (O_2874,N_24596,N_24312);
nor UO_2875 (O_2875,N_24958,N_24928);
and UO_2876 (O_2876,N_24045,N_24816);
nor UO_2877 (O_2877,N_24932,N_24558);
nor UO_2878 (O_2878,N_24705,N_24145);
nor UO_2879 (O_2879,N_24508,N_24576);
nor UO_2880 (O_2880,N_24356,N_24853);
nor UO_2881 (O_2881,N_24680,N_24686);
and UO_2882 (O_2882,N_24579,N_24745);
nand UO_2883 (O_2883,N_24033,N_24739);
nand UO_2884 (O_2884,N_24895,N_24573);
nor UO_2885 (O_2885,N_24640,N_24590);
or UO_2886 (O_2886,N_24444,N_24398);
xor UO_2887 (O_2887,N_24029,N_24395);
or UO_2888 (O_2888,N_24998,N_24553);
nor UO_2889 (O_2889,N_24645,N_24440);
or UO_2890 (O_2890,N_24669,N_24685);
xnor UO_2891 (O_2891,N_24187,N_24366);
xor UO_2892 (O_2892,N_24902,N_24074);
xnor UO_2893 (O_2893,N_24372,N_24343);
and UO_2894 (O_2894,N_24795,N_24776);
nand UO_2895 (O_2895,N_24734,N_24615);
xor UO_2896 (O_2896,N_24482,N_24115);
and UO_2897 (O_2897,N_24396,N_24219);
nor UO_2898 (O_2898,N_24609,N_24469);
and UO_2899 (O_2899,N_24104,N_24420);
xnor UO_2900 (O_2900,N_24755,N_24322);
xnor UO_2901 (O_2901,N_24161,N_24584);
or UO_2902 (O_2902,N_24081,N_24999);
and UO_2903 (O_2903,N_24186,N_24815);
nor UO_2904 (O_2904,N_24040,N_24009);
nand UO_2905 (O_2905,N_24627,N_24761);
and UO_2906 (O_2906,N_24879,N_24352);
nor UO_2907 (O_2907,N_24047,N_24498);
and UO_2908 (O_2908,N_24654,N_24332);
and UO_2909 (O_2909,N_24016,N_24825);
nand UO_2910 (O_2910,N_24353,N_24298);
and UO_2911 (O_2911,N_24379,N_24928);
xnor UO_2912 (O_2912,N_24469,N_24043);
nor UO_2913 (O_2913,N_24351,N_24170);
and UO_2914 (O_2914,N_24564,N_24026);
xnor UO_2915 (O_2915,N_24836,N_24024);
nor UO_2916 (O_2916,N_24409,N_24294);
xor UO_2917 (O_2917,N_24761,N_24372);
and UO_2918 (O_2918,N_24788,N_24310);
nand UO_2919 (O_2919,N_24171,N_24862);
and UO_2920 (O_2920,N_24714,N_24157);
nor UO_2921 (O_2921,N_24966,N_24954);
or UO_2922 (O_2922,N_24893,N_24407);
xor UO_2923 (O_2923,N_24879,N_24208);
nand UO_2924 (O_2924,N_24466,N_24855);
or UO_2925 (O_2925,N_24855,N_24893);
nand UO_2926 (O_2926,N_24383,N_24235);
nor UO_2927 (O_2927,N_24592,N_24168);
nor UO_2928 (O_2928,N_24595,N_24320);
nor UO_2929 (O_2929,N_24862,N_24383);
or UO_2930 (O_2930,N_24982,N_24896);
nor UO_2931 (O_2931,N_24412,N_24356);
and UO_2932 (O_2932,N_24464,N_24924);
and UO_2933 (O_2933,N_24566,N_24860);
nand UO_2934 (O_2934,N_24367,N_24735);
xnor UO_2935 (O_2935,N_24274,N_24535);
or UO_2936 (O_2936,N_24801,N_24062);
nor UO_2937 (O_2937,N_24351,N_24722);
nor UO_2938 (O_2938,N_24926,N_24044);
or UO_2939 (O_2939,N_24730,N_24648);
xor UO_2940 (O_2940,N_24711,N_24661);
and UO_2941 (O_2941,N_24074,N_24204);
nor UO_2942 (O_2942,N_24552,N_24730);
nor UO_2943 (O_2943,N_24069,N_24822);
xor UO_2944 (O_2944,N_24715,N_24919);
and UO_2945 (O_2945,N_24996,N_24138);
and UO_2946 (O_2946,N_24672,N_24423);
and UO_2947 (O_2947,N_24779,N_24200);
or UO_2948 (O_2948,N_24926,N_24032);
xor UO_2949 (O_2949,N_24329,N_24668);
nor UO_2950 (O_2950,N_24714,N_24834);
xor UO_2951 (O_2951,N_24765,N_24596);
nand UO_2952 (O_2952,N_24738,N_24457);
xor UO_2953 (O_2953,N_24957,N_24711);
and UO_2954 (O_2954,N_24276,N_24093);
and UO_2955 (O_2955,N_24722,N_24882);
and UO_2956 (O_2956,N_24865,N_24316);
or UO_2957 (O_2957,N_24632,N_24282);
or UO_2958 (O_2958,N_24790,N_24591);
nand UO_2959 (O_2959,N_24275,N_24388);
or UO_2960 (O_2960,N_24976,N_24122);
or UO_2961 (O_2961,N_24457,N_24834);
nand UO_2962 (O_2962,N_24376,N_24685);
xnor UO_2963 (O_2963,N_24603,N_24562);
xor UO_2964 (O_2964,N_24326,N_24965);
or UO_2965 (O_2965,N_24961,N_24633);
xnor UO_2966 (O_2966,N_24765,N_24443);
or UO_2967 (O_2967,N_24618,N_24850);
or UO_2968 (O_2968,N_24085,N_24747);
xnor UO_2969 (O_2969,N_24675,N_24594);
and UO_2970 (O_2970,N_24713,N_24809);
xnor UO_2971 (O_2971,N_24355,N_24194);
nor UO_2972 (O_2972,N_24123,N_24597);
nor UO_2973 (O_2973,N_24800,N_24677);
xor UO_2974 (O_2974,N_24411,N_24801);
xor UO_2975 (O_2975,N_24016,N_24368);
and UO_2976 (O_2976,N_24037,N_24651);
nand UO_2977 (O_2977,N_24944,N_24953);
or UO_2978 (O_2978,N_24399,N_24684);
or UO_2979 (O_2979,N_24288,N_24191);
or UO_2980 (O_2980,N_24948,N_24589);
nor UO_2981 (O_2981,N_24084,N_24376);
xnor UO_2982 (O_2982,N_24549,N_24140);
nor UO_2983 (O_2983,N_24763,N_24186);
nand UO_2984 (O_2984,N_24142,N_24376);
nor UO_2985 (O_2985,N_24451,N_24848);
or UO_2986 (O_2986,N_24557,N_24715);
xor UO_2987 (O_2987,N_24683,N_24877);
nor UO_2988 (O_2988,N_24371,N_24754);
and UO_2989 (O_2989,N_24240,N_24410);
nor UO_2990 (O_2990,N_24558,N_24215);
nor UO_2991 (O_2991,N_24168,N_24343);
nand UO_2992 (O_2992,N_24812,N_24573);
and UO_2993 (O_2993,N_24203,N_24774);
nand UO_2994 (O_2994,N_24346,N_24196);
and UO_2995 (O_2995,N_24026,N_24265);
or UO_2996 (O_2996,N_24091,N_24808);
and UO_2997 (O_2997,N_24453,N_24646);
nand UO_2998 (O_2998,N_24706,N_24205);
nor UO_2999 (O_2999,N_24333,N_24129);
endmodule